// Generator : SpinalHDL v1.4.2    git head : d65b8c01ad060f0c2a8c80ed1b1e9da6e6240532
// Component : SInt64fixTo63_0_ROUNDTOINF
// Git hash  : d151d69c0adb8fba5bc1372ea3c015e94de78c79
// Date      : 20/07/2020, 11:11:11
// Designer	: Zhengpeng Liao



module SInt64fixTo63_0_ROUNDTOINF (
  input      [63:0]   din,
  output     [63:0]   dout
);

  assign dout = din;

endmodule
