// Generator : SpinalHDL v1.4.0    git head : ecb5a80b713566f417ea3ea061f9969e73770a7f
// Date      : 21/05/2020, 11:11:29
// Component : ImpLoadUnit



module ImpLoadUnit (
  input               axi4_aw_valid,
  output              axi4_aw_ready,
  input      [31:0]   axi4_aw_payload_addr,
  input      [3:0]    axi4_aw_payload_id,
  input      [7:0]    axi4_aw_payload_len,
  input      [2:0]    axi4_aw_payload_size,
  input      [1:0]    axi4_aw_payload_burst,
  input               axi4_w_valid,
  output              axi4_w_ready,
  input      [31:0]   axi4_w_payload_data,
  input      [3:0]    axi4_w_payload_strb,
  input               axi4_w_payload_last,
  output              axi4_b_valid,
  input               axi4_b_ready,
  output     [3:0]    axi4_b_payload_id,
  output     [1:0]    axi4_b_payload_resp,
  output              io_impulse_out_valid,
  output     [15:0]   io_impulse_out_payload_0_0_real,
  output     [15:0]   io_impulse_out_payload_0_0_imag,
  output     [15:0]   io_impulse_out_payload_0_1_real,
  output     [15:0]   io_impulse_out_payload_0_1_imag,
  output     [15:0]   io_impulse_out_payload_1_0_real,
  output     [15:0]   io_impulse_out_payload_1_0_imag,
  output     [15:0]   io_impulse_out_payload_1_1_real,
  output     [15:0]   io_impulse_out_payload_1_1_imag,
  output     [15:0]   io_impulse_out_payload_2_0_real,
  output     [15:0]   io_impulse_out_payload_2_0_imag,
  output     [15:0]   io_impulse_out_payload_2_1_real,
  output     [15:0]   io_impulse_out_payload_2_1_imag,
  output     [15:0]   io_impulse_out_payload_3_0_real,
  output     [15:0]   io_impulse_out_payload_3_0_imag,
  output     [15:0]   io_impulse_out_payload_3_1_real,
  output     [15:0]   io_impulse_out_payload_3_1_imag,
  output     [15:0]   io_impulse_out_payload_4_0_real,
  output     [15:0]   io_impulse_out_payload_4_0_imag,
  output     [15:0]   io_impulse_out_payload_4_1_real,
  output     [15:0]   io_impulse_out_payload_4_1_imag,
  output     [15:0]   io_impulse_out_payload_5_0_real,
  output     [15:0]   io_impulse_out_payload_5_0_imag,
  output     [15:0]   io_impulse_out_payload_5_1_real,
  output     [15:0]   io_impulse_out_payload_5_1_imag,
  output     [15:0]   io_impulse_out_payload_6_0_real,
  output     [15:0]   io_impulse_out_payload_6_0_imag,
  output     [15:0]   io_impulse_out_payload_6_1_real,
  output     [15:0]   io_impulse_out_payload_6_1_imag,
  output     [15:0]   io_impulse_out_payload_7_0_real,
  output     [15:0]   io_impulse_out_payload_7_0_imag,
  output     [15:0]   io_impulse_out_payload_7_1_real,
  output     [15:0]   io_impulse_out_payload_7_1_imag,
  output     [15:0]   io_impulse_out_payload_8_0_real,
  output     [15:0]   io_impulse_out_payload_8_0_imag,
  output     [15:0]   io_impulse_out_payload_8_1_real,
  output     [15:0]   io_impulse_out_payload_8_1_imag,
  output     [15:0]   io_impulse_out_payload_9_0_real,
  output     [15:0]   io_impulse_out_payload_9_0_imag,
  output     [15:0]   io_impulse_out_payload_9_1_real,
  output     [15:0]   io_impulse_out_payload_9_1_imag,
  output     [15:0]   io_impulse_out_payload_10_0_real,
  output     [15:0]   io_impulse_out_payload_10_0_imag,
  output     [15:0]   io_impulse_out_payload_10_1_real,
  output     [15:0]   io_impulse_out_payload_10_1_imag,
  output     [15:0]   io_impulse_out_payload_11_0_real,
  output     [15:0]   io_impulse_out_payload_11_0_imag,
  output     [15:0]   io_impulse_out_payload_11_1_real,
  output     [15:0]   io_impulse_out_payload_11_1_imag,
  output     [15:0]   io_impulse_out_payload_12_0_real,
  output     [15:0]   io_impulse_out_payload_12_0_imag,
  output     [15:0]   io_impulse_out_payload_12_1_real,
  output     [15:0]   io_impulse_out_payload_12_1_imag,
  output     [15:0]   io_impulse_out_payload_13_0_real,
  output     [15:0]   io_impulse_out_payload_13_0_imag,
  output     [15:0]   io_impulse_out_payload_13_1_real,
  output     [15:0]   io_impulse_out_payload_13_1_imag,
  output     [15:0]   io_impulse_out_payload_14_0_real,
  output     [15:0]   io_impulse_out_payload_14_0_imag,
  output     [15:0]   io_impulse_out_payload_14_1_real,
  output     [15:0]   io_impulse_out_payload_14_1_imag,
  output     [15:0]   io_impulse_out_payload_15_0_real,
  output     [15:0]   io_impulse_out_payload_15_0_imag,
  output     [15:0]   io_impulse_out_payload_15_1_real,
  output     [15:0]   io_impulse_out_payload_15_1_imag,
  output     [15:0]   io_impulse_out_payload_16_0_real,
  output     [15:0]   io_impulse_out_payload_16_0_imag,
  output     [15:0]   io_impulse_out_payload_16_1_real,
  output     [15:0]   io_impulse_out_payload_16_1_imag,
  output     [15:0]   io_impulse_out_payload_17_0_real,
  output     [15:0]   io_impulse_out_payload_17_0_imag,
  output     [15:0]   io_impulse_out_payload_17_1_real,
  output     [15:0]   io_impulse_out_payload_17_1_imag,
  output     [15:0]   io_impulse_out_payload_18_0_real,
  output     [15:0]   io_impulse_out_payload_18_0_imag,
  output     [15:0]   io_impulse_out_payload_18_1_real,
  output     [15:0]   io_impulse_out_payload_18_1_imag,
  output     [15:0]   io_impulse_out_payload_19_0_real,
  output     [15:0]   io_impulse_out_payload_19_0_imag,
  output     [15:0]   io_impulse_out_payload_19_1_real,
  output     [15:0]   io_impulse_out_payload_19_1_imag,
  output     [15:0]   io_impulse_out_payload_20_0_real,
  output     [15:0]   io_impulse_out_payload_20_0_imag,
  output     [15:0]   io_impulse_out_payload_20_1_real,
  output     [15:0]   io_impulse_out_payload_20_1_imag,
  output     [15:0]   io_impulse_out_payload_21_0_real,
  output     [15:0]   io_impulse_out_payload_21_0_imag,
  output     [15:0]   io_impulse_out_payload_21_1_real,
  output     [15:0]   io_impulse_out_payload_21_1_imag,
  output     [15:0]   io_impulse_out_payload_22_0_real,
  output     [15:0]   io_impulse_out_payload_22_0_imag,
  output     [15:0]   io_impulse_out_payload_22_1_real,
  output     [15:0]   io_impulse_out_payload_22_1_imag,
  output     [15:0]   io_impulse_out_payload_23_0_real,
  output     [15:0]   io_impulse_out_payload_23_0_imag,
  output     [15:0]   io_impulse_out_payload_23_1_real,
  output     [15:0]   io_impulse_out_payload_23_1_imag,
  output     [15:0]   io_impulse_out_payload_24_0_real,
  output     [15:0]   io_impulse_out_payload_24_0_imag,
  output     [15:0]   io_impulse_out_payload_24_1_real,
  output     [15:0]   io_impulse_out_payload_24_1_imag,
  output     [15:0]   io_impulse_out_payload_25_0_real,
  output     [15:0]   io_impulse_out_payload_25_0_imag,
  output     [15:0]   io_impulse_out_payload_25_1_real,
  output     [15:0]   io_impulse_out_payload_25_1_imag,
  output     [15:0]   io_impulse_out_payload_26_0_real,
  output     [15:0]   io_impulse_out_payload_26_0_imag,
  output     [15:0]   io_impulse_out_payload_26_1_real,
  output     [15:0]   io_impulse_out_payload_26_1_imag,
  output     [15:0]   io_impulse_out_payload_27_0_real,
  output     [15:0]   io_impulse_out_payload_27_0_imag,
  output     [15:0]   io_impulse_out_payload_27_1_real,
  output     [15:0]   io_impulse_out_payload_27_1_imag,
  output     [15:0]   io_impulse_out_payload_28_0_real,
  output     [15:0]   io_impulse_out_payload_28_0_imag,
  output     [15:0]   io_impulse_out_payload_28_1_real,
  output     [15:0]   io_impulse_out_payload_28_1_imag,
  output     [15:0]   io_impulse_out_payload_29_0_real,
  output     [15:0]   io_impulse_out_payload_29_0_imag,
  output     [15:0]   io_impulse_out_payload_29_1_real,
  output     [15:0]   io_impulse_out_payload_29_1_imag,
  output     [15:0]   io_impulse_out_payload_30_0_real,
  output     [15:0]   io_impulse_out_payload_30_0_imag,
  output     [15:0]   io_impulse_out_payload_30_1_real,
  output     [15:0]   io_impulse_out_payload_30_1_imag,
  output     [15:0]   io_impulse_out_payload_31_0_real,
  output     [15:0]   io_impulse_out_payload_31_0_imag,
  output     [15:0]   io_impulse_out_payload_31_1_real,
  output     [15:0]   io_impulse_out_payload_31_1_imag,
  output     [15:0]   io_impulse_out_payload_32_0_real,
  output     [15:0]   io_impulse_out_payload_32_0_imag,
  output     [15:0]   io_impulse_out_payload_32_1_real,
  output     [15:0]   io_impulse_out_payload_32_1_imag,
  output     [15:0]   io_impulse_out_payload_33_0_real,
  output     [15:0]   io_impulse_out_payload_33_0_imag,
  output     [15:0]   io_impulse_out_payload_33_1_real,
  output     [15:0]   io_impulse_out_payload_33_1_imag,
  output     [15:0]   io_impulse_out_payload_34_0_real,
  output     [15:0]   io_impulse_out_payload_34_0_imag,
  output     [15:0]   io_impulse_out_payload_34_1_real,
  output     [15:0]   io_impulse_out_payload_34_1_imag,
  output     [15:0]   io_impulse_out_payload_35_0_real,
  output     [15:0]   io_impulse_out_payload_35_0_imag,
  output     [15:0]   io_impulse_out_payload_35_1_real,
  output     [15:0]   io_impulse_out_payload_35_1_imag,
  output     [15:0]   io_impulse_out_payload_36_0_real,
  output     [15:0]   io_impulse_out_payload_36_0_imag,
  output     [15:0]   io_impulse_out_payload_36_1_real,
  output     [15:0]   io_impulse_out_payload_36_1_imag,
  output     [15:0]   io_impulse_out_payload_37_0_real,
  output     [15:0]   io_impulse_out_payload_37_0_imag,
  output     [15:0]   io_impulse_out_payload_37_1_real,
  output     [15:0]   io_impulse_out_payload_37_1_imag,
  output     [15:0]   io_impulse_out_payload_38_0_real,
  output     [15:0]   io_impulse_out_payload_38_0_imag,
  output     [15:0]   io_impulse_out_payload_38_1_real,
  output     [15:0]   io_impulse_out_payload_38_1_imag,
  output     [15:0]   io_impulse_out_payload_39_0_real,
  output     [15:0]   io_impulse_out_payload_39_0_imag,
  output     [15:0]   io_impulse_out_payload_39_1_real,
  output     [15:0]   io_impulse_out_payload_39_1_imag,
  output     [15:0]   io_impulse_out_payload_40_0_real,
  output     [15:0]   io_impulse_out_payload_40_0_imag,
  output     [15:0]   io_impulse_out_payload_40_1_real,
  output     [15:0]   io_impulse_out_payload_40_1_imag,
  output     [15:0]   io_impulse_out_payload_41_0_real,
  output     [15:0]   io_impulse_out_payload_41_0_imag,
  output     [15:0]   io_impulse_out_payload_41_1_real,
  output     [15:0]   io_impulse_out_payload_41_1_imag,
  output     [15:0]   io_impulse_out_payload_42_0_real,
  output     [15:0]   io_impulse_out_payload_42_0_imag,
  output     [15:0]   io_impulse_out_payload_42_1_real,
  output     [15:0]   io_impulse_out_payload_42_1_imag,
  output     [15:0]   io_impulse_out_payload_43_0_real,
  output     [15:0]   io_impulse_out_payload_43_0_imag,
  output     [15:0]   io_impulse_out_payload_43_1_real,
  output     [15:0]   io_impulse_out_payload_43_1_imag,
  output     [15:0]   io_impulse_out_payload_44_0_real,
  output     [15:0]   io_impulse_out_payload_44_0_imag,
  output     [15:0]   io_impulse_out_payload_44_1_real,
  output     [15:0]   io_impulse_out_payload_44_1_imag,
  output     [15:0]   io_impulse_out_payload_45_0_real,
  output     [15:0]   io_impulse_out_payload_45_0_imag,
  output     [15:0]   io_impulse_out_payload_45_1_real,
  output     [15:0]   io_impulse_out_payload_45_1_imag,
  output     [15:0]   io_impulse_out_payload_46_0_real,
  output     [15:0]   io_impulse_out_payload_46_0_imag,
  output     [15:0]   io_impulse_out_payload_46_1_real,
  output     [15:0]   io_impulse_out_payload_46_1_imag,
  output     [15:0]   io_impulse_out_payload_47_0_real,
  output     [15:0]   io_impulse_out_payload_47_0_imag,
  output     [15:0]   io_impulse_out_payload_47_1_real,
  output     [15:0]   io_impulse_out_payload_47_1_imag,
  output     [15:0]   io_impulse_out_payload_48_0_real,
  output     [15:0]   io_impulse_out_payload_48_0_imag,
  output     [15:0]   io_impulse_out_payload_48_1_real,
  output     [15:0]   io_impulse_out_payload_48_1_imag,
  output     [15:0]   io_impulse_out_payload_49_0_real,
  output     [15:0]   io_impulse_out_payload_49_0_imag,
  output     [15:0]   io_impulse_out_payload_49_1_real,
  output     [15:0]   io_impulse_out_payload_49_1_imag,
  input               clk,
  input               reset 
);
  wire       [31:0]   _zz_203_;
  wire       [31:0]   _zz_204_;
  wire       [31:0]   _zz_205_;
  wire       [31:0]   _zz_206_;
  wire       [31:0]   _zz_207_;
  wire       [31:0]   _zz_208_;
  wire       [31:0]   _zz_209_;
  wire       [31:0]   _zz_210_;
  wire       [31:0]   _zz_211_;
  wire       [31:0]   _zz_212_;
  wire       [31:0]   _zz_213_;
  wire       [31:0]   _zz_214_;
  wire       [31:0]   _zz_215_;
  wire       [31:0]   _zz_216_;
  wire       [31:0]   _zz_217_;
  wire       [31:0]   _zz_218_;
  wire       [31:0]   _zz_219_;
  wire       [31:0]   _zz_220_;
  wire       [31:0]   _zz_221_;
  wire       [31:0]   _zz_222_;
  wire       [31:0]   _zz_223_;
  wire       [31:0]   _zz_224_;
  wire       [31:0]   _zz_225_;
  wire       [31:0]   _zz_226_;
  wire       [31:0]   _zz_227_;
  wire       [31:0]   _zz_228_;
  wire       [31:0]   _zz_229_;
  wire       [31:0]   _zz_230_;
  wire       [31:0]   _zz_231_;
  wire       [31:0]   _zz_232_;
  wire       [31:0]   _zz_233_;
  wire       [31:0]   _zz_234_;
  wire       [31:0]   _zz_235_;
  wire       [31:0]   _zz_236_;
  wire       [31:0]   _zz_237_;
  wire       [31:0]   _zz_238_;
  wire       [31:0]   _zz_239_;
  wire       [31:0]   _zz_240_;
  wire       [31:0]   _zz_241_;
  wire       [31:0]   _zz_242_;
  wire       [31:0]   _zz_243_;
  wire       [31:0]   _zz_244_;
  wire       [31:0]   _zz_245_;
  wire       [31:0]   _zz_246_;
  wire       [31:0]   _zz_247_;
  wire       [31:0]   _zz_248_;
  wire       [31:0]   _zz_249_;
  wire       [31:0]   _zz_250_;
  wire       [31:0]   _zz_251_;
  wire       [31:0]   _zz_252_;
  wire       [31:0]   _zz_253_;
  wire       [31:0]   _zz_254_;
  wire       [31:0]   _zz_255_;
  wire       [31:0]   _zz_256_;
  wire       [31:0]   _zz_257_;
  wire       [31:0]   _zz_258_;
  wire       [31:0]   _zz_259_;
  wire       [31:0]   _zz_260_;
  wire       [31:0]   _zz_261_;
  wire       [31:0]   _zz_262_;
  wire       [31:0]   _zz_263_;
  wire       [31:0]   _zz_264_;
  wire       [31:0]   _zz_265_;
  wire       [31:0]   _zz_266_;
  wire       [31:0]   _zz_267_;
  wire       [31:0]   _zz_268_;
  wire       [31:0]   _zz_269_;
  wire       [31:0]   _zz_270_;
  wire       [31:0]   _zz_271_;
  wire       [31:0]   _zz_272_;
  wire       [31:0]   _zz_273_;
  wire       [31:0]   _zz_274_;
  wire       [31:0]   _zz_275_;
  wire       [31:0]   _zz_276_;
  wire       [31:0]   _zz_277_;
  wire       [31:0]   _zz_278_;
  wire       [31:0]   _zz_279_;
  wire       [31:0]   _zz_280_;
  wire       [31:0]   _zz_281_;
  wire       [31:0]   _zz_282_;
  wire       [31:0]   _zz_283_;
  wire       [31:0]   _zz_284_;
  wire       [31:0]   _zz_285_;
  wire       [31:0]   _zz_286_;
  wire       [31:0]   _zz_287_;
  wire       [31:0]   _zz_288_;
  wire       [31:0]   _zz_289_;
  wire       [31:0]   _zz_290_;
  wire       [31:0]   _zz_291_;
  wire       [31:0]   _zz_292_;
  wire       [31:0]   _zz_293_;
  wire       [31:0]   _zz_294_;
  wire       [31:0]   _zz_295_;
  wire       [31:0]   _zz_296_;
  wire       [31:0]   _zz_297_;
  wire       [31:0]   _zz_298_;
  wire       [31:0]   _zz_299_;
  wire       [31:0]   _zz_300_;
  wire       [31:0]   _zz_301_;
  wire       [31:0]   _zz_302_;
  reg        [11:0]   _zz_303_;
  wire       [11:0]   _zz_304_;
  wire       [11:0]   _zz_305_;
  wire       [11:0]   _zz_306_;
  wire       [0:0]    _zz_307_;
  wire       [31:0]   _zz_308_;
  wire       [5:0]    _zz_309_;
  wire       [31:0]   _zz_310_;
  wire       [5:0]    _zz_311_;
  wire       [31:0]   _zz_312_;
  wire       [5:0]    _zz_313_;
  wire       [31:0]   _zz_314_;
  wire       [5:0]    _zz_315_;
  wire       [31:0]   _zz_316_;
  wire       [5:0]    _zz_317_;
  wire       [31:0]   _zz_318_;
  wire       [5:0]    _zz_319_;
  wire       [31:0]   _zz_320_;
  wire       [5:0]    _zz_321_;
  wire       [31:0]   _zz_322_;
  wire       [5:0]    _zz_323_;
  wire       [31:0]   _zz_324_;
  wire       [5:0]    _zz_325_;
  wire       [31:0]   _zz_326_;
  wire       [5:0]    _zz_327_;
  wire       [31:0]   _zz_328_;
  wire       [5:0]    _zz_329_;
  wire       [31:0]   _zz_330_;
  wire       [5:0]    _zz_331_;
  wire       [31:0]   _zz_332_;
  wire       [5:0]    _zz_333_;
  wire       [31:0]   _zz_334_;
  wire       [5:0]    _zz_335_;
  wire       [31:0]   _zz_336_;
  wire       [5:0]    _zz_337_;
  wire       [31:0]   _zz_338_;
  wire       [5:0]    _zz_339_;
  wire       [31:0]   _zz_340_;
  wire       [5:0]    _zz_341_;
  wire       [31:0]   _zz_342_;
  wire       [5:0]    _zz_343_;
  wire       [31:0]   _zz_344_;
  wire       [5:0]    _zz_345_;
  wire       [31:0]   _zz_346_;
  wire       [5:0]    _zz_347_;
  wire       [31:0]   _zz_348_;
  wire       [5:0]    _zz_349_;
  wire       [31:0]   _zz_350_;
  wire       [5:0]    _zz_351_;
  wire       [31:0]   _zz_352_;
  wire       [5:0]    _zz_353_;
  wire       [31:0]   _zz_354_;
  wire       [5:0]    _zz_355_;
  wire       [31:0]   _zz_356_;
  wire       [5:0]    _zz_357_;
  wire       [31:0]   _zz_358_;
  wire       [5:0]    _zz_359_;
  wire       [31:0]   _zz_360_;
  wire       [5:0]    _zz_361_;
  wire       [31:0]   _zz_362_;
  wire       [5:0]    _zz_363_;
  wire       [31:0]   _zz_364_;
  wire       [5:0]    _zz_365_;
  wire       [31:0]   _zz_366_;
  wire       [5:0]    _zz_367_;
  wire       [31:0]   _zz_368_;
  wire       [5:0]    _zz_369_;
  wire       [31:0]   _zz_370_;
  wire       [5:0]    _zz_371_;
  wire       [31:0]   _zz_372_;
  wire       [5:0]    _zz_373_;
  wire       [31:0]   _zz_374_;
  wire       [5:0]    _zz_375_;
  wire       [31:0]   _zz_376_;
  wire       [5:0]    _zz_377_;
  wire       [31:0]   _zz_378_;
  wire       [5:0]    _zz_379_;
  wire       [31:0]   _zz_380_;
  wire       [5:0]    _zz_381_;
  wire       [31:0]   _zz_382_;
  wire       [5:0]    _zz_383_;
  wire       [31:0]   _zz_384_;
  wire       [5:0]    _zz_385_;
  wire       [31:0]   _zz_386_;
  wire       [5:0]    _zz_387_;
  wire       [31:0]   _zz_388_;
  wire       [5:0]    _zz_389_;
  wire       [31:0]   _zz_390_;
  wire       [5:0]    _zz_391_;
  wire       [31:0]   _zz_392_;
  wire       [5:0]    _zz_393_;
  wire       [31:0]   _zz_394_;
  wire       [5:0]    _zz_395_;
  wire       [31:0]   _zz_396_;
  wire       [5:0]    _zz_397_;
  wire       [31:0]   _zz_398_;
  wire       [5:0]    _zz_399_;
  wire       [31:0]   _zz_400_;
  wire       [5:0]    _zz_401_;
  wire       [31:0]   _zz_402_;
  wire       [5:0]    _zz_403_;
  wire       [31:0]   _zz_404_;
  wire       [5:0]    _zz_405_;
  wire       [31:0]   _zz_406_;
  wire       [5:0]    _zz_407_;
  wire       [0:0]    _zz_408_;
  wire       [13:0]   _zz_409_;
  wire       [5:0]    _zz_410_;
  wire       [5:0]    _zz_411_;
  wire       [5:0]    _zz_412_;
  wire       [5:0]    _zz_413_;
  wire       [5:0]    _zz_414_;
  wire       [5:0]    _zz_415_;
  wire       [5:0]    _zz_416_;
  wire       [5:0]    _zz_417_;
  wire       [5:0]    _zz_418_;
  wire       [5:0]    _zz_419_;
  wire       [5:0]    _zz_420_;
  wire       [5:0]    _zz_421_;
  wire       [5:0]    _zz_422_;
  wire       [5:0]    _zz_423_;
  wire       [5:0]    _zz_424_;
  wire       [5:0]    _zz_425_;
  wire       [5:0]    _zz_426_;
  wire       [5:0]    _zz_427_;
  wire       [5:0]    _zz_428_;
  wire       [5:0]    _zz_429_;
  wire       [5:0]    _zz_430_;
  wire       [5:0]    _zz_431_;
  wire       [5:0]    _zz_432_;
  wire       [5:0]    _zz_433_;
  wire       [5:0]    _zz_434_;
  wire       [5:0]    _zz_435_;
  wire       [5:0]    _zz_436_;
  wire       [5:0]    _zz_437_;
  wire       [5:0]    _zz_438_;
  wire       [5:0]    _zz_439_;
  wire       [5:0]    _zz_440_;
  wire       [5:0]    _zz_441_;
  wire       [5:0]    _zz_442_;
  wire       [5:0]    _zz_443_;
  wire       [5:0]    _zz_444_;
  wire       [5:0]    _zz_445_;
  wire       [5:0]    _zz_446_;
  wire       [5:0]    _zz_447_;
  wire       [5:0]    _zz_448_;
  wire       [5:0]    _zz_449_;
  wire       [5:0]    _zz_450_;
  wire       [5:0]    _zz_451_;
  wire       [5:0]    _zz_452_;
  wire       [5:0]    _zz_453_;
  wire       [5:0]    _zz_454_;
  wire       [5:0]    _zz_455_;
  wire       [5:0]    _zz_456_;
  wire       [5:0]    _zz_457_;
  wire       [5:0]    _zz_458_;
  wire       [5:0]    _zz_459_;
  wire       [5:0]    _zz_460_;
  wire       [5:0]    _zz_461_;
  wire       [5:0]    _zz_462_;
  wire       [5:0]    _zz_463_;
  wire       [5:0]    _zz_464_;
  wire       [5:0]    _zz_465_;
  wire       [5:0]    _zz_466_;
  wire       [5:0]    _zz_467_;
  wire       [5:0]    _zz_468_;
  wire       [5:0]    _zz_469_;
  wire       [5:0]    _zz_470_;
  wire       [5:0]    _zz_471_;
  wire       [5:0]    _zz_472_;
  wire       [5:0]    _zz_473_;
  wire       [5:0]    _zz_474_;
  wire       [5:0]    _zz_475_;
  wire       [5:0]    _zz_476_;
  wire       [5:0]    _zz_477_;
  wire       [5:0]    _zz_478_;
  wire       [5:0]    _zz_479_;
  wire       [5:0]    _zz_480_;
  wire       [5:0]    _zz_481_;
  wire       [5:0]    _zz_482_;
  wire       [5:0]    _zz_483_;
  wire       [5:0]    _zz_484_;
  wire       [5:0]    _zz_485_;
  wire       [5:0]    _zz_486_;
  wire       [5:0]    _zz_487_;
  wire       [5:0]    _zz_488_;
  wire       [5:0]    _zz_489_;
  wire       [5:0]    _zz_490_;
  wire       [5:0]    _zz_491_;
  wire       [5:0]    _zz_492_;
  wire       [5:0]    _zz_493_;
  wire       [5:0]    _zz_494_;
  wire       [5:0]    _zz_495_;
  wire       [5:0]    _zz_496_;
  wire       [5:0]    _zz_497_;
  wire       [5:0]    _zz_498_;
  wire       [5:0]    _zz_499_;
  wire       [5:0]    _zz_500_;
  wire       [5:0]    _zz_501_;
  wire       [5:0]    _zz_502_;
  wire       [5:0]    _zz_503_;
  wire       [5:0]    _zz_504_;
  wire       [5:0]    _zz_505_;
  wire       [5:0]    _zz_506_;
  wire       [5:0]    _zz_507_;
  wire       [5:0]    _zz_508_;
  wire       [5:0]    _zz_509_;
  wire                _zz_510_;
  wire                _zz_511_;
  wire                _zz_512_;
  wire                _zz_513_;
  wire                _zz_514_;
  wire                _zz_515_;
  wire                _zz_516_;
  wire                _zz_517_;
  wire                _zz_518_;
  wire                _zz_519_;
  wire                _zz_520_;
  wire                _zz_521_;
  wire                _zz_522_;
  wire                _zz_523_;
  wire                _zz_524_;
  wire                _zz_525_;
  wire                _zz_526_;
  wire                _zz_527_;
  wire                _zz_528_;
  wire                _zz_529_;
  wire                _zz_530_;
  wire                _zz_531_;
  wire                _zz_532_;
  wire                _zz_533_;
  wire                _zz_534_;
  wire                _zz_535_;
  wire                _zz_536_;
  wire                _zz_537_;
  wire                _zz_538_;
  wire                _zz_539_;
  wire                _zz_540_;
  wire                _zz_541_;
  wire                _zz_542_;
  wire                _zz_543_;
  wire                _zz_544_;
  wire                _zz_545_;
  wire                _zz_546_;
  wire                _zz_547_;
  wire                _zz_548_;
  wire                _zz_549_;
  wire                _zz_550_;
  wire                _zz_551_;
  wire                _zz_552_;
  wire                _zz_553_;
  wire                _zz_554_;
  wire                _zz_555_;
  wire                _zz_556_;
  wire                _zz_557_;
  wire                _zz_558_;
  wire                _zz_559_;
  reg        [31:0]   aw_area_awaddr_r;
  reg        [7:0]    aw_area_awlen_r;
  reg        [2:0]    aw_area_awsize_r;
  reg        [3:0]    aw_area_awid_r;
  wire                transfer_done;
  reg                 transfer_done_1_;
  reg        [31:0]   load_data_area_current_addr;
  reg        [31:0]   Axi4Incr_result;
  wire       [19:0]   Axi4Incr_highCat;
  wire       [0:0]    Axi4Incr_sizeValue;
  wire       [11:0]   Axi4Incr_alignMask;
  wire       [11:0]   Axi4Incr_base;
  wire       [11:0]   Axi4Incr_baseIncr;
  reg        [1:0]    _zz_1_;
  wire       [1:0]    Axi4Incr_wrapCase;
  reg        [31:0]   axi4_w_payload_data_regNext;
  reg                 current_mem_addr_willIncrement;
  wire                current_mem_addr_willClear;
  reg        [13:0]   current_mem_addr_valueNext;
  reg        [13:0]   current_mem_addr_value;
  wire                current_mem_addr_willOverflowIfInc;
  wire                current_mem_addr_willOverflow;
  reg                 _zz_2_;
  wire       [13:0]   _zz_3_;
  wire       [31:0]   _zz_4_;
  wire       [13:0]   _zz_5_;
  wire       [31:0]   _zz_6_;
  wire       [13:0]   _zz_7_;
  wire       [31:0]   _zz_8_;
  wire       [13:0]   _zz_9_;
  wire       [31:0]   _zz_10_;
  wire       [13:0]   _zz_11_;
  wire       [31:0]   _zz_12_;
  wire       [13:0]   _zz_13_;
  wire       [31:0]   _zz_14_;
  wire       [13:0]   _zz_15_;
  wire       [31:0]   _zz_16_;
  wire       [13:0]   _zz_17_;
  wire       [31:0]   _zz_18_;
  wire       [13:0]   _zz_19_;
  wire       [31:0]   _zz_20_;
  wire       [13:0]   _zz_21_;
  wire       [31:0]   _zz_22_;
  wire       [13:0]   _zz_23_;
  wire       [31:0]   _zz_24_;
  wire       [13:0]   _zz_25_;
  wire       [31:0]   _zz_26_;
  wire       [13:0]   _zz_27_;
  wire       [31:0]   _zz_28_;
  wire       [13:0]   _zz_29_;
  wire       [31:0]   _zz_30_;
  wire       [13:0]   _zz_31_;
  wire       [31:0]   _zz_32_;
  wire       [13:0]   _zz_33_;
  wire       [31:0]   _zz_34_;
  wire       [13:0]   _zz_35_;
  wire       [31:0]   _zz_36_;
  wire       [13:0]   _zz_37_;
  wire       [31:0]   _zz_38_;
  wire       [13:0]   _zz_39_;
  wire       [31:0]   _zz_40_;
  wire       [13:0]   _zz_41_;
  wire       [31:0]   _zz_42_;
  wire       [13:0]   _zz_43_;
  wire       [31:0]   _zz_44_;
  wire       [13:0]   _zz_45_;
  wire       [31:0]   _zz_46_;
  wire       [13:0]   _zz_47_;
  wire       [31:0]   _zz_48_;
  wire       [13:0]   _zz_49_;
  wire       [31:0]   _zz_50_;
  wire       [13:0]   _zz_51_;
  wire       [31:0]   _zz_52_;
  wire       [13:0]   _zz_53_;
  wire       [31:0]   _zz_54_;
  wire       [13:0]   _zz_55_;
  wire       [31:0]   _zz_56_;
  wire       [13:0]   _zz_57_;
  wire       [31:0]   _zz_58_;
  wire       [13:0]   _zz_59_;
  wire       [31:0]   _zz_60_;
  wire       [13:0]   _zz_61_;
  wire       [31:0]   _zz_62_;
  wire       [13:0]   _zz_63_;
  wire       [31:0]   _zz_64_;
  wire       [13:0]   _zz_65_;
  wire       [31:0]   _zz_66_;
  wire       [13:0]   _zz_67_;
  wire       [31:0]   _zz_68_;
  wire       [13:0]   _zz_69_;
  wire       [31:0]   _zz_70_;
  wire       [13:0]   _zz_71_;
  wire       [31:0]   _zz_72_;
  wire       [13:0]   _zz_73_;
  wire       [31:0]   _zz_74_;
  wire       [13:0]   _zz_75_;
  wire       [31:0]   _zz_76_;
  wire       [13:0]   _zz_77_;
  wire       [31:0]   _zz_78_;
  wire       [13:0]   _zz_79_;
  wire       [31:0]   _zz_80_;
  wire       [13:0]   _zz_81_;
  wire       [31:0]   _zz_82_;
  wire       [13:0]   _zz_83_;
  wire       [31:0]   _zz_84_;
  wire       [13:0]   _zz_85_;
  wire       [31:0]   _zz_86_;
  wire       [13:0]   _zz_87_;
  wire       [31:0]   _zz_88_;
  wire       [13:0]   _zz_89_;
  wire       [31:0]   _zz_90_;
  wire       [13:0]   _zz_91_;
  wire       [31:0]   _zz_92_;
  wire       [13:0]   _zz_93_;
  wire       [31:0]   _zz_94_;
  wire       [13:0]   _zz_95_;
  wire       [31:0]   _zz_96_;
  wire       [13:0]   _zz_97_;
  wire       [31:0]   _zz_98_;
  wire       [13:0]   _zz_99_;
  wire       [31:0]   _zz_100_;
  wire       [13:0]   _zz_101_;
  wire       [31:0]   _zz_102_;
  wire       [13:0]   _zz_103_;
  wire       [31:0]   _zz_104_;
  wire       [13:0]   _zz_105_;
  wire       [31:0]   _zz_106_;
  wire       [13:0]   _zz_107_;
  wire       [31:0]   _zz_108_;
  wire       [13:0]   _zz_109_;
  wire       [31:0]   _zz_110_;
  wire       [13:0]   _zz_111_;
  wire       [31:0]   _zz_112_;
  wire       [13:0]   _zz_113_;
  wire       [31:0]   _zz_114_;
  wire       [13:0]   _zz_115_;
  wire       [31:0]   _zz_116_;
  wire       [13:0]   _zz_117_;
  wire       [31:0]   _zz_118_;
  wire       [13:0]   _zz_119_;
  wire       [31:0]   _zz_120_;
  wire       [13:0]   _zz_121_;
  wire       [31:0]   _zz_122_;
  wire       [13:0]   _zz_123_;
  wire       [31:0]   _zz_124_;
  wire       [13:0]   _zz_125_;
  wire       [31:0]   _zz_126_;
  wire       [13:0]   _zz_127_;
  wire       [31:0]   _zz_128_;
  wire       [13:0]   _zz_129_;
  wire       [31:0]   _zz_130_;
  wire       [13:0]   _zz_131_;
  wire       [31:0]   _zz_132_;
  wire       [13:0]   _zz_133_;
  wire       [31:0]   _zz_134_;
  wire       [13:0]   _zz_135_;
  wire       [31:0]   _zz_136_;
  wire       [13:0]   _zz_137_;
  wire       [31:0]   _zz_138_;
  wire       [13:0]   _zz_139_;
  wire       [31:0]   _zz_140_;
  wire       [13:0]   _zz_141_;
  wire       [31:0]   _zz_142_;
  wire       [13:0]   _zz_143_;
  wire       [31:0]   _zz_144_;
  wire       [13:0]   _zz_145_;
  wire       [31:0]   _zz_146_;
  wire       [13:0]   _zz_147_;
  wire       [31:0]   _zz_148_;
  wire       [13:0]   _zz_149_;
  wire       [31:0]   _zz_150_;
  wire       [13:0]   _zz_151_;
  wire       [31:0]   _zz_152_;
  wire       [13:0]   _zz_153_;
  wire       [31:0]   _zz_154_;
  wire       [13:0]   _zz_155_;
  wire       [31:0]   _zz_156_;
  wire       [13:0]   _zz_157_;
  wire       [31:0]   _zz_158_;
  wire       [13:0]   _zz_159_;
  wire       [31:0]   _zz_160_;
  wire       [13:0]   _zz_161_;
  wire       [31:0]   _zz_162_;
  wire       [13:0]   _zz_163_;
  wire       [31:0]   _zz_164_;
  wire       [13:0]   _zz_165_;
  wire       [31:0]   _zz_166_;
  wire       [13:0]   _zz_167_;
  wire       [31:0]   _zz_168_;
  wire       [13:0]   _zz_169_;
  wire       [31:0]   _zz_170_;
  wire       [13:0]   _zz_171_;
  wire       [31:0]   _zz_172_;
  wire       [13:0]   _zz_173_;
  wire       [31:0]   _zz_174_;
  wire       [13:0]   _zz_175_;
  wire       [31:0]   _zz_176_;
  wire       [13:0]   _zz_177_;
  wire       [31:0]   _zz_178_;
  wire       [13:0]   _zz_179_;
  wire       [31:0]   _zz_180_;
  wire       [13:0]   _zz_181_;
  wire       [31:0]   _zz_182_;
  wire       [13:0]   _zz_183_;
  wire       [31:0]   _zz_184_;
  wire       [13:0]   _zz_185_;
  wire       [31:0]   _zz_186_;
  wire       [13:0]   _zz_187_;
  wire       [31:0]   _zz_188_;
  wire       [13:0]   _zz_189_;
  wire       [31:0]   _zz_190_;
  wire       [13:0]   _zz_191_;
  wire       [31:0]   _zz_192_;
  wire       [13:0]   _zz_193_;
  wire       [31:0]   _zz_194_;
  wire       [13:0]   _zz_195_;
  wire       [31:0]   _zz_196_;
  wire       [13:0]   _zz_197_;
  wire       [31:0]   _zz_198_;
  wire       [13:0]   _zz_199_;
  wire       [31:0]   _zz_200_;
  wire       [13:0]   _zz_201_;
  wire       [31:0]   _zz_202_;
  reg [31:0] int_ram_array_0 [0:63];
  reg [31:0] int_ram_array_1 [0:63];
  reg [31:0] int_ram_array_2 [0:63];
  reg [31:0] int_ram_array_3 [0:63];
  reg [31:0] int_ram_array_4 [0:63];
  reg [31:0] int_ram_array_5 [0:63];
  reg [31:0] int_ram_array_6 [0:63];
  reg [31:0] int_ram_array_7 [0:63];
  reg [31:0] int_ram_array_8 [0:63];
  reg [31:0] int_ram_array_9 [0:63];
  reg [31:0] int_ram_array_10 [0:63];
  reg [31:0] int_ram_array_11 [0:63];
  reg [31:0] int_ram_array_12 [0:63];
  reg [31:0] int_ram_array_13 [0:63];
  reg [31:0] int_ram_array_14 [0:63];
  reg [31:0] int_ram_array_15 [0:63];
  reg [31:0] int_ram_array_16 [0:63];
  reg [31:0] int_ram_array_17 [0:63];
  reg [31:0] int_ram_array_18 [0:63];
  reg [31:0] int_ram_array_19 [0:63];
  reg [31:0] int_ram_array_20 [0:63];
  reg [31:0] int_ram_array_21 [0:63];
  reg [31:0] int_ram_array_22 [0:63];
  reg [31:0] int_ram_array_23 [0:63];
  reg [31:0] int_ram_array_24 [0:63];
  reg [31:0] int_ram_array_25 [0:63];
  reg [31:0] int_ram_array_26 [0:63];
  reg [31:0] int_ram_array_27 [0:63];
  reg [31:0] int_ram_array_28 [0:63];
  reg [31:0] int_ram_array_29 [0:63];
  reg [31:0] int_ram_array_30 [0:63];
  reg [31:0] int_ram_array_31 [0:63];
  reg [31:0] int_ram_array_32 [0:63];
  reg [31:0] int_ram_array_33 [0:63];
  reg [31:0] int_ram_array_34 [0:63];
  reg [31:0] int_ram_array_35 [0:63];
  reg [31:0] int_ram_array_36 [0:63];
  reg [31:0] int_ram_array_37 [0:63];
  reg [31:0] int_ram_array_38 [0:63];
  reg [31:0] int_ram_array_39 [0:63];
  reg [31:0] int_ram_array_40 [0:63];
  reg [31:0] int_ram_array_41 [0:63];
  reg [31:0] int_ram_array_42 [0:63];
  reg [31:0] int_ram_array_43 [0:63];
  reg [31:0] int_ram_array_44 [0:63];
  reg [31:0] int_ram_array_45 [0:63];
  reg [31:0] int_ram_array_46 [0:63];
  reg [31:0] int_ram_array_47 [0:63];
  reg [31:0] int_ram_array_48 [0:63];
  reg [31:0] int_ram_array_49 [0:63];

  assign _zz_304_ = aw_area_awaddr_r[11 : 0];
  assign _zz_305_ = _zz_304_;
  assign _zz_306_ = {11'd0, Axi4Incr_sizeValue};
  assign _zz_307_ = transfer_done_1_;
  assign _zz_308_ = (load_data_area_current_addr - 32'h0);
  assign _zz_309_ = _zz_308_[5:0];
  assign _zz_310_ = (load_data_area_current_addr - 32'h00000040);
  assign _zz_311_ = _zz_310_[5:0];
  assign _zz_312_ = (load_data_area_current_addr - 32'h00000080);
  assign _zz_313_ = _zz_312_[5:0];
  assign _zz_314_ = (load_data_area_current_addr - 32'h000000c0);
  assign _zz_315_ = _zz_314_[5:0];
  assign _zz_316_ = (load_data_area_current_addr - 32'h00000100);
  assign _zz_317_ = _zz_316_[5:0];
  assign _zz_318_ = (load_data_area_current_addr - 32'h00000140);
  assign _zz_319_ = _zz_318_[5:0];
  assign _zz_320_ = (load_data_area_current_addr - 32'h00000180);
  assign _zz_321_ = _zz_320_[5:0];
  assign _zz_322_ = (load_data_area_current_addr - 32'h000001c0);
  assign _zz_323_ = _zz_322_[5:0];
  assign _zz_324_ = (load_data_area_current_addr - 32'h00000200);
  assign _zz_325_ = _zz_324_[5:0];
  assign _zz_326_ = (load_data_area_current_addr - 32'h00000240);
  assign _zz_327_ = _zz_326_[5:0];
  assign _zz_328_ = (load_data_area_current_addr - 32'h00000280);
  assign _zz_329_ = _zz_328_[5:0];
  assign _zz_330_ = (load_data_area_current_addr - 32'h000002c0);
  assign _zz_331_ = _zz_330_[5:0];
  assign _zz_332_ = (load_data_area_current_addr - 32'h00000300);
  assign _zz_333_ = _zz_332_[5:0];
  assign _zz_334_ = (load_data_area_current_addr - 32'h00000340);
  assign _zz_335_ = _zz_334_[5:0];
  assign _zz_336_ = (load_data_area_current_addr - 32'h00000380);
  assign _zz_337_ = _zz_336_[5:0];
  assign _zz_338_ = (load_data_area_current_addr - 32'h000003c0);
  assign _zz_339_ = _zz_338_[5:0];
  assign _zz_340_ = (load_data_area_current_addr - 32'h00000400);
  assign _zz_341_ = _zz_340_[5:0];
  assign _zz_342_ = (load_data_area_current_addr - 32'h00000440);
  assign _zz_343_ = _zz_342_[5:0];
  assign _zz_344_ = (load_data_area_current_addr - 32'h00000480);
  assign _zz_345_ = _zz_344_[5:0];
  assign _zz_346_ = (load_data_area_current_addr - 32'h000004c0);
  assign _zz_347_ = _zz_346_[5:0];
  assign _zz_348_ = (load_data_area_current_addr - 32'h00000500);
  assign _zz_349_ = _zz_348_[5:0];
  assign _zz_350_ = (load_data_area_current_addr - 32'h00000540);
  assign _zz_351_ = _zz_350_[5:0];
  assign _zz_352_ = (load_data_area_current_addr - 32'h00000580);
  assign _zz_353_ = _zz_352_[5:0];
  assign _zz_354_ = (load_data_area_current_addr - 32'h000005c0);
  assign _zz_355_ = _zz_354_[5:0];
  assign _zz_356_ = (load_data_area_current_addr - 32'h00000600);
  assign _zz_357_ = _zz_356_[5:0];
  assign _zz_358_ = (load_data_area_current_addr - 32'h00000640);
  assign _zz_359_ = _zz_358_[5:0];
  assign _zz_360_ = (load_data_area_current_addr - 32'h00000680);
  assign _zz_361_ = _zz_360_[5:0];
  assign _zz_362_ = (load_data_area_current_addr - 32'h000006c0);
  assign _zz_363_ = _zz_362_[5:0];
  assign _zz_364_ = (load_data_area_current_addr - 32'h00000700);
  assign _zz_365_ = _zz_364_[5:0];
  assign _zz_366_ = (load_data_area_current_addr - 32'h00000740);
  assign _zz_367_ = _zz_366_[5:0];
  assign _zz_368_ = (load_data_area_current_addr - 32'h00000780);
  assign _zz_369_ = _zz_368_[5:0];
  assign _zz_370_ = (load_data_area_current_addr - 32'h000007c0);
  assign _zz_371_ = _zz_370_[5:0];
  assign _zz_372_ = (load_data_area_current_addr - 32'h00000800);
  assign _zz_373_ = _zz_372_[5:0];
  assign _zz_374_ = (load_data_area_current_addr - 32'h00000840);
  assign _zz_375_ = _zz_374_[5:0];
  assign _zz_376_ = (load_data_area_current_addr - 32'h00000880);
  assign _zz_377_ = _zz_376_[5:0];
  assign _zz_378_ = (load_data_area_current_addr - 32'h000008c0);
  assign _zz_379_ = _zz_378_[5:0];
  assign _zz_380_ = (load_data_area_current_addr - 32'h00000900);
  assign _zz_381_ = _zz_380_[5:0];
  assign _zz_382_ = (load_data_area_current_addr - 32'h00000940);
  assign _zz_383_ = _zz_382_[5:0];
  assign _zz_384_ = (load_data_area_current_addr - 32'h00000980);
  assign _zz_385_ = _zz_384_[5:0];
  assign _zz_386_ = (load_data_area_current_addr - 32'h000009c0);
  assign _zz_387_ = _zz_386_[5:0];
  assign _zz_388_ = (load_data_area_current_addr - 32'h00000a00);
  assign _zz_389_ = _zz_388_[5:0];
  assign _zz_390_ = (load_data_area_current_addr - 32'h00000a40);
  assign _zz_391_ = _zz_390_[5:0];
  assign _zz_392_ = (load_data_area_current_addr - 32'h00000a80);
  assign _zz_393_ = _zz_392_[5:0];
  assign _zz_394_ = (load_data_area_current_addr - 32'h00000ac0);
  assign _zz_395_ = _zz_394_[5:0];
  assign _zz_396_ = (load_data_area_current_addr - 32'h00000b00);
  assign _zz_397_ = _zz_396_[5:0];
  assign _zz_398_ = (load_data_area_current_addr - 32'h00000b40);
  assign _zz_399_ = _zz_398_[5:0];
  assign _zz_400_ = (load_data_area_current_addr - 32'h00000b80);
  assign _zz_401_ = _zz_400_[5:0];
  assign _zz_402_ = (load_data_area_current_addr - 32'h00000bc0);
  assign _zz_403_ = _zz_402_[5:0];
  assign _zz_404_ = (load_data_area_current_addr - 32'h00000c00);
  assign _zz_405_ = _zz_404_[5:0];
  assign _zz_406_ = (load_data_area_current_addr - 32'h00000c40);
  assign _zz_407_ = _zz_406_[5:0];
  assign _zz_408_ = current_mem_addr_willIncrement;
  assign _zz_409_ = {13'd0, _zz_408_};
  assign _zz_410_ = _zz_3_[5:0];
  assign _zz_411_ = _zz_5_[5:0];
  assign _zz_412_ = _zz_7_[5:0];
  assign _zz_413_ = _zz_9_[5:0];
  assign _zz_414_ = _zz_11_[5:0];
  assign _zz_415_ = _zz_13_[5:0];
  assign _zz_416_ = _zz_15_[5:0];
  assign _zz_417_ = _zz_17_[5:0];
  assign _zz_418_ = _zz_19_[5:0];
  assign _zz_419_ = _zz_21_[5:0];
  assign _zz_420_ = _zz_23_[5:0];
  assign _zz_421_ = _zz_25_[5:0];
  assign _zz_422_ = _zz_27_[5:0];
  assign _zz_423_ = _zz_29_[5:0];
  assign _zz_424_ = _zz_31_[5:0];
  assign _zz_425_ = _zz_33_[5:0];
  assign _zz_426_ = _zz_35_[5:0];
  assign _zz_427_ = _zz_37_[5:0];
  assign _zz_428_ = _zz_39_[5:0];
  assign _zz_429_ = _zz_41_[5:0];
  assign _zz_430_ = _zz_43_[5:0];
  assign _zz_431_ = _zz_45_[5:0];
  assign _zz_432_ = _zz_47_[5:0];
  assign _zz_433_ = _zz_49_[5:0];
  assign _zz_434_ = _zz_51_[5:0];
  assign _zz_435_ = _zz_53_[5:0];
  assign _zz_436_ = _zz_55_[5:0];
  assign _zz_437_ = _zz_57_[5:0];
  assign _zz_438_ = _zz_59_[5:0];
  assign _zz_439_ = _zz_61_[5:0];
  assign _zz_440_ = _zz_63_[5:0];
  assign _zz_441_ = _zz_65_[5:0];
  assign _zz_442_ = _zz_67_[5:0];
  assign _zz_443_ = _zz_69_[5:0];
  assign _zz_444_ = _zz_71_[5:0];
  assign _zz_445_ = _zz_73_[5:0];
  assign _zz_446_ = _zz_75_[5:0];
  assign _zz_447_ = _zz_77_[5:0];
  assign _zz_448_ = _zz_79_[5:0];
  assign _zz_449_ = _zz_81_[5:0];
  assign _zz_450_ = _zz_83_[5:0];
  assign _zz_451_ = _zz_85_[5:0];
  assign _zz_452_ = _zz_87_[5:0];
  assign _zz_453_ = _zz_89_[5:0];
  assign _zz_454_ = _zz_91_[5:0];
  assign _zz_455_ = _zz_93_[5:0];
  assign _zz_456_ = _zz_95_[5:0];
  assign _zz_457_ = _zz_97_[5:0];
  assign _zz_458_ = _zz_99_[5:0];
  assign _zz_459_ = _zz_101_[5:0];
  assign _zz_460_ = _zz_103_[5:0];
  assign _zz_461_ = _zz_105_[5:0];
  assign _zz_462_ = _zz_107_[5:0];
  assign _zz_463_ = _zz_109_[5:0];
  assign _zz_464_ = _zz_111_[5:0];
  assign _zz_465_ = _zz_113_[5:0];
  assign _zz_466_ = _zz_115_[5:0];
  assign _zz_467_ = _zz_117_[5:0];
  assign _zz_468_ = _zz_119_[5:0];
  assign _zz_469_ = _zz_121_[5:0];
  assign _zz_470_ = _zz_123_[5:0];
  assign _zz_471_ = _zz_125_[5:0];
  assign _zz_472_ = _zz_127_[5:0];
  assign _zz_473_ = _zz_129_[5:0];
  assign _zz_474_ = _zz_131_[5:0];
  assign _zz_475_ = _zz_133_[5:0];
  assign _zz_476_ = _zz_135_[5:0];
  assign _zz_477_ = _zz_137_[5:0];
  assign _zz_478_ = _zz_139_[5:0];
  assign _zz_479_ = _zz_141_[5:0];
  assign _zz_480_ = _zz_143_[5:0];
  assign _zz_481_ = _zz_145_[5:0];
  assign _zz_482_ = _zz_147_[5:0];
  assign _zz_483_ = _zz_149_[5:0];
  assign _zz_484_ = _zz_151_[5:0];
  assign _zz_485_ = _zz_153_[5:0];
  assign _zz_486_ = _zz_155_[5:0];
  assign _zz_487_ = _zz_157_[5:0];
  assign _zz_488_ = _zz_159_[5:0];
  assign _zz_489_ = _zz_161_[5:0];
  assign _zz_490_ = _zz_163_[5:0];
  assign _zz_491_ = _zz_165_[5:0];
  assign _zz_492_ = _zz_167_[5:0];
  assign _zz_493_ = _zz_169_[5:0];
  assign _zz_494_ = _zz_171_[5:0];
  assign _zz_495_ = _zz_173_[5:0];
  assign _zz_496_ = _zz_175_[5:0];
  assign _zz_497_ = _zz_177_[5:0];
  assign _zz_498_ = _zz_179_[5:0];
  assign _zz_499_ = _zz_181_[5:0];
  assign _zz_500_ = _zz_183_[5:0];
  assign _zz_501_ = _zz_185_[5:0];
  assign _zz_502_ = _zz_187_[5:0];
  assign _zz_503_ = _zz_189_[5:0];
  assign _zz_504_ = _zz_191_[5:0];
  assign _zz_505_ = _zz_193_[5:0];
  assign _zz_506_ = _zz_195_[5:0];
  assign _zz_507_ = _zz_197_[5:0];
  assign _zz_508_ = _zz_199_[5:0];
  assign _zz_509_ = _zz_201_[5:0];
  assign _zz_510_ = ((32'h0 <= load_data_area_current_addr) && (load_data_area_current_addr < 32'h0000003f));
  assign _zz_511_ = ((32'h00000040 <= load_data_area_current_addr) && (load_data_area_current_addr < 32'h0000007f));
  assign _zz_512_ = ((32'h00000080 <= load_data_area_current_addr) && (load_data_area_current_addr < 32'h000000bf));
  assign _zz_513_ = ((32'h000000c0 <= load_data_area_current_addr) && (load_data_area_current_addr < 32'h000000ff));
  assign _zz_514_ = ((32'h00000100 <= load_data_area_current_addr) && (load_data_area_current_addr < 32'h0000013f));
  assign _zz_515_ = ((32'h00000140 <= load_data_area_current_addr) && (load_data_area_current_addr < 32'h0000017f));
  assign _zz_516_ = ((32'h00000180 <= load_data_area_current_addr) && (load_data_area_current_addr < 32'h000001bf));
  assign _zz_517_ = ((32'h000001c0 <= load_data_area_current_addr) && (load_data_area_current_addr < 32'h000001ff));
  assign _zz_518_ = ((32'h00000200 <= load_data_area_current_addr) && (load_data_area_current_addr < 32'h0000023f));
  assign _zz_519_ = ((32'h00000240 <= load_data_area_current_addr) && (load_data_area_current_addr < 32'h0000027f));
  assign _zz_520_ = ((32'h00000280 <= load_data_area_current_addr) && (load_data_area_current_addr < 32'h000002bf));
  assign _zz_521_ = ((32'h000002c0 <= load_data_area_current_addr) && (load_data_area_current_addr < 32'h000002ff));
  assign _zz_522_ = ((32'h00000300 <= load_data_area_current_addr) && (load_data_area_current_addr < 32'h0000033f));
  assign _zz_523_ = ((32'h00000340 <= load_data_area_current_addr) && (load_data_area_current_addr < 32'h0000037f));
  assign _zz_524_ = ((32'h00000380 <= load_data_area_current_addr) && (load_data_area_current_addr < 32'h000003bf));
  assign _zz_525_ = ((32'h000003c0 <= load_data_area_current_addr) && (load_data_area_current_addr < 32'h000003ff));
  assign _zz_526_ = ((32'h00000400 <= load_data_area_current_addr) && (load_data_area_current_addr < 32'h0000043f));
  assign _zz_527_ = ((32'h00000440 <= load_data_area_current_addr) && (load_data_area_current_addr < 32'h0000047f));
  assign _zz_528_ = ((32'h00000480 <= load_data_area_current_addr) && (load_data_area_current_addr < 32'h000004bf));
  assign _zz_529_ = ((32'h000004c0 <= load_data_area_current_addr) && (load_data_area_current_addr < 32'h000004ff));
  assign _zz_530_ = ((32'h00000500 <= load_data_area_current_addr) && (load_data_area_current_addr < 32'h0000053f));
  assign _zz_531_ = ((32'h00000540 <= load_data_area_current_addr) && (load_data_area_current_addr < 32'h0000057f));
  assign _zz_532_ = ((32'h00000580 <= load_data_area_current_addr) && (load_data_area_current_addr < 32'h000005bf));
  assign _zz_533_ = ((32'h000005c0 <= load_data_area_current_addr) && (load_data_area_current_addr < 32'h000005ff));
  assign _zz_534_ = ((32'h00000600 <= load_data_area_current_addr) && (load_data_area_current_addr < 32'h0000063f));
  assign _zz_535_ = ((32'h00000640 <= load_data_area_current_addr) && (load_data_area_current_addr < 32'h0000067f));
  assign _zz_536_ = ((32'h00000680 <= load_data_area_current_addr) && (load_data_area_current_addr < 32'h000006bf));
  assign _zz_537_ = ((32'h000006c0 <= load_data_area_current_addr) && (load_data_area_current_addr < 32'h000006ff));
  assign _zz_538_ = ((32'h00000700 <= load_data_area_current_addr) && (load_data_area_current_addr < 32'h0000073f));
  assign _zz_539_ = ((32'h00000740 <= load_data_area_current_addr) && (load_data_area_current_addr < 32'h0000077f));
  assign _zz_540_ = ((32'h00000780 <= load_data_area_current_addr) && (load_data_area_current_addr < 32'h000007bf));
  assign _zz_541_ = ((32'h000007c0 <= load_data_area_current_addr) && (load_data_area_current_addr < 32'h000007ff));
  assign _zz_542_ = ((32'h00000800 <= load_data_area_current_addr) && (load_data_area_current_addr < 32'h0000083f));
  assign _zz_543_ = ((32'h00000840 <= load_data_area_current_addr) && (load_data_area_current_addr < 32'h0000087f));
  assign _zz_544_ = ((32'h00000880 <= load_data_area_current_addr) && (load_data_area_current_addr < 32'h000008bf));
  assign _zz_545_ = ((32'h000008c0 <= load_data_area_current_addr) && (load_data_area_current_addr < 32'h000008ff));
  assign _zz_546_ = ((32'h00000900 <= load_data_area_current_addr) && (load_data_area_current_addr < 32'h0000093f));
  assign _zz_547_ = ((32'h00000940 <= load_data_area_current_addr) && (load_data_area_current_addr < 32'h0000097f));
  assign _zz_548_ = ((32'h00000980 <= load_data_area_current_addr) && (load_data_area_current_addr < 32'h000009bf));
  assign _zz_549_ = ((32'h000009c0 <= load_data_area_current_addr) && (load_data_area_current_addr < 32'h000009ff));
  assign _zz_550_ = ((32'h00000a00 <= load_data_area_current_addr) && (load_data_area_current_addr < 32'h00000a3f));
  assign _zz_551_ = ((32'h00000a40 <= load_data_area_current_addr) && (load_data_area_current_addr < 32'h00000a7f));
  assign _zz_552_ = ((32'h00000a80 <= load_data_area_current_addr) && (load_data_area_current_addr < 32'h00000abf));
  assign _zz_553_ = ((32'h00000ac0 <= load_data_area_current_addr) && (load_data_area_current_addr < 32'h00000aff));
  assign _zz_554_ = ((32'h00000b00 <= load_data_area_current_addr) && (load_data_area_current_addr < 32'h00000b3f));
  assign _zz_555_ = ((32'h00000b40 <= load_data_area_current_addr) && (load_data_area_current_addr < 32'h00000b7f));
  assign _zz_556_ = ((32'h00000b80 <= load_data_area_current_addr) && (load_data_area_current_addr < 32'h00000bbf));
  assign _zz_557_ = ((32'h00000bc0 <= load_data_area_current_addr) && (load_data_area_current_addr < 32'h00000bff));
  assign _zz_558_ = ((32'h00000c00 <= load_data_area_current_addr) && (load_data_area_current_addr < 32'h00000c3f));
  assign _zz_559_ = ((32'h00000c40 <= load_data_area_current_addr) && (load_data_area_current_addr < 32'h00000c7f));
  always @ (posedge clk) begin
    if(_zz_510_) begin
      int_ram_array_0[_zz_309_] <= axi4_w_payload_data;
    end
  end

  assign _zz_203_ = int_ram_array_0[_zz_410_];
  assign _zz_204_ = int_ram_array_0[_zz_411_];
  always @ (posedge clk) begin
    if(_zz_511_) begin
      int_ram_array_1[_zz_311_] <= axi4_w_payload_data;
    end
  end

  assign _zz_205_ = int_ram_array_1[_zz_412_];
  assign _zz_206_ = int_ram_array_1[_zz_413_];
  always @ (posedge clk) begin
    if(_zz_512_) begin
      int_ram_array_2[_zz_313_] <= axi4_w_payload_data;
    end
  end

  assign _zz_207_ = int_ram_array_2[_zz_414_];
  assign _zz_208_ = int_ram_array_2[_zz_415_];
  always @ (posedge clk) begin
    if(_zz_513_) begin
      int_ram_array_3[_zz_315_] <= axi4_w_payload_data;
    end
  end

  assign _zz_209_ = int_ram_array_3[_zz_416_];
  assign _zz_210_ = int_ram_array_3[_zz_417_];
  always @ (posedge clk) begin
    if(_zz_514_) begin
      int_ram_array_4[_zz_317_] <= axi4_w_payload_data;
    end
  end

  assign _zz_211_ = int_ram_array_4[_zz_418_];
  assign _zz_212_ = int_ram_array_4[_zz_419_];
  always @ (posedge clk) begin
    if(_zz_515_) begin
      int_ram_array_5[_zz_319_] <= axi4_w_payload_data;
    end
  end

  assign _zz_213_ = int_ram_array_5[_zz_420_];
  assign _zz_214_ = int_ram_array_5[_zz_421_];
  always @ (posedge clk) begin
    if(_zz_516_) begin
      int_ram_array_6[_zz_321_] <= axi4_w_payload_data;
    end
  end

  assign _zz_215_ = int_ram_array_6[_zz_422_];
  assign _zz_216_ = int_ram_array_6[_zz_423_];
  always @ (posedge clk) begin
    if(_zz_517_) begin
      int_ram_array_7[_zz_323_] <= axi4_w_payload_data;
    end
  end

  assign _zz_217_ = int_ram_array_7[_zz_424_];
  assign _zz_218_ = int_ram_array_7[_zz_425_];
  always @ (posedge clk) begin
    if(_zz_518_) begin
      int_ram_array_8[_zz_325_] <= axi4_w_payload_data;
    end
  end

  assign _zz_219_ = int_ram_array_8[_zz_426_];
  assign _zz_220_ = int_ram_array_8[_zz_427_];
  always @ (posedge clk) begin
    if(_zz_519_) begin
      int_ram_array_9[_zz_327_] <= axi4_w_payload_data;
    end
  end

  assign _zz_221_ = int_ram_array_9[_zz_428_];
  assign _zz_222_ = int_ram_array_9[_zz_429_];
  always @ (posedge clk) begin
    if(_zz_520_) begin
      int_ram_array_10[_zz_329_] <= axi4_w_payload_data;
    end
  end

  assign _zz_223_ = int_ram_array_10[_zz_430_];
  assign _zz_224_ = int_ram_array_10[_zz_431_];
  always @ (posedge clk) begin
    if(_zz_521_) begin
      int_ram_array_11[_zz_331_] <= axi4_w_payload_data;
    end
  end

  assign _zz_225_ = int_ram_array_11[_zz_432_];
  assign _zz_226_ = int_ram_array_11[_zz_433_];
  always @ (posedge clk) begin
    if(_zz_522_) begin
      int_ram_array_12[_zz_333_] <= axi4_w_payload_data;
    end
  end

  assign _zz_227_ = int_ram_array_12[_zz_434_];
  assign _zz_228_ = int_ram_array_12[_zz_435_];
  always @ (posedge clk) begin
    if(_zz_523_) begin
      int_ram_array_13[_zz_335_] <= axi4_w_payload_data;
    end
  end

  assign _zz_229_ = int_ram_array_13[_zz_436_];
  assign _zz_230_ = int_ram_array_13[_zz_437_];
  always @ (posedge clk) begin
    if(_zz_524_) begin
      int_ram_array_14[_zz_337_] <= axi4_w_payload_data;
    end
  end

  assign _zz_231_ = int_ram_array_14[_zz_438_];
  assign _zz_232_ = int_ram_array_14[_zz_439_];
  always @ (posedge clk) begin
    if(_zz_525_) begin
      int_ram_array_15[_zz_339_] <= axi4_w_payload_data;
    end
  end

  assign _zz_233_ = int_ram_array_15[_zz_440_];
  assign _zz_234_ = int_ram_array_15[_zz_441_];
  always @ (posedge clk) begin
    if(_zz_526_) begin
      int_ram_array_16[_zz_341_] <= axi4_w_payload_data;
    end
  end

  assign _zz_235_ = int_ram_array_16[_zz_442_];
  assign _zz_236_ = int_ram_array_16[_zz_443_];
  always @ (posedge clk) begin
    if(_zz_527_) begin
      int_ram_array_17[_zz_343_] <= axi4_w_payload_data;
    end
  end

  assign _zz_237_ = int_ram_array_17[_zz_444_];
  assign _zz_238_ = int_ram_array_17[_zz_445_];
  always @ (posedge clk) begin
    if(_zz_528_) begin
      int_ram_array_18[_zz_345_] <= axi4_w_payload_data;
    end
  end

  assign _zz_239_ = int_ram_array_18[_zz_446_];
  assign _zz_240_ = int_ram_array_18[_zz_447_];
  always @ (posedge clk) begin
    if(_zz_529_) begin
      int_ram_array_19[_zz_347_] <= axi4_w_payload_data;
    end
  end

  assign _zz_241_ = int_ram_array_19[_zz_448_];
  assign _zz_242_ = int_ram_array_19[_zz_449_];
  always @ (posedge clk) begin
    if(_zz_530_) begin
      int_ram_array_20[_zz_349_] <= axi4_w_payload_data;
    end
  end

  assign _zz_243_ = int_ram_array_20[_zz_450_];
  assign _zz_244_ = int_ram_array_20[_zz_451_];
  always @ (posedge clk) begin
    if(_zz_531_) begin
      int_ram_array_21[_zz_351_] <= axi4_w_payload_data;
    end
  end

  assign _zz_245_ = int_ram_array_21[_zz_452_];
  assign _zz_246_ = int_ram_array_21[_zz_453_];
  always @ (posedge clk) begin
    if(_zz_532_) begin
      int_ram_array_22[_zz_353_] <= axi4_w_payload_data;
    end
  end

  assign _zz_247_ = int_ram_array_22[_zz_454_];
  assign _zz_248_ = int_ram_array_22[_zz_455_];
  always @ (posedge clk) begin
    if(_zz_533_) begin
      int_ram_array_23[_zz_355_] <= axi4_w_payload_data;
    end
  end

  assign _zz_249_ = int_ram_array_23[_zz_456_];
  assign _zz_250_ = int_ram_array_23[_zz_457_];
  always @ (posedge clk) begin
    if(_zz_534_) begin
      int_ram_array_24[_zz_357_] <= axi4_w_payload_data;
    end
  end

  assign _zz_251_ = int_ram_array_24[_zz_458_];
  assign _zz_252_ = int_ram_array_24[_zz_459_];
  always @ (posedge clk) begin
    if(_zz_535_) begin
      int_ram_array_25[_zz_359_] <= axi4_w_payload_data;
    end
  end

  assign _zz_253_ = int_ram_array_25[_zz_460_];
  assign _zz_254_ = int_ram_array_25[_zz_461_];
  always @ (posedge clk) begin
    if(_zz_536_) begin
      int_ram_array_26[_zz_361_] <= axi4_w_payload_data;
    end
  end

  assign _zz_255_ = int_ram_array_26[_zz_462_];
  assign _zz_256_ = int_ram_array_26[_zz_463_];
  always @ (posedge clk) begin
    if(_zz_537_) begin
      int_ram_array_27[_zz_363_] <= axi4_w_payload_data;
    end
  end

  assign _zz_257_ = int_ram_array_27[_zz_464_];
  assign _zz_258_ = int_ram_array_27[_zz_465_];
  always @ (posedge clk) begin
    if(_zz_538_) begin
      int_ram_array_28[_zz_365_] <= axi4_w_payload_data;
    end
  end

  assign _zz_259_ = int_ram_array_28[_zz_466_];
  assign _zz_260_ = int_ram_array_28[_zz_467_];
  always @ (posedge clk) begin
    if(_zz_539_) begin
      int_ram_array_29[_zz_367_] <= axi4_w_payload_data;
    end
  end

  assign _zz_261_ = int_ram_array_29[_zz_468_];
  assign _zz_262_ = int_ram_array_29[_zz_469_];
  always @ (posedge clk) begin
    if(_zz_540_) begin
      int_ram_array_30[_zz_369_] <= axi4_w_payload_data;
    end
  end

  assign _zz_263_ = int_ram_array_30[_zz_470_];
  assign _zz_264_ = int_ram_array_30[_zz_471_];
  always @ (posedge clk) begin
    if(_zz_541_) begin
      int_ram_array_31[_zz_371_] <= axi4_w_payload_data;
    end
  end

  assign _zz_265_ = int_ram_array_31[_zz_472_];
  assign _zz_266_ = int_ram_array_31[_zz_473_];
  always @ (posedge clk) begin
    if(_zz_542_) begin
      int_ram_array_32[_zz_373_] <= axi4_w_payload_data;
    end
  end

  assign _zz_267_ = int_ram_array_32[_zz_474_];
  assign _zz_268_ = int_ram_array_32[_zz_475_];
  always @ (posedge clk) begin
    if(_zz_543_) begin
      int_ram_array_33[_zz_375_] <= axi4_w_payload_data;
    end
  end

  assign _zz_269_ = int_ram_array_33[_zz_476_];
  assign _zz_270_ = int_ram_array_33[_zz_477_];
  always @ (posedge clk) begin
    if(_zz_544_) begin
      int_ram_array_34[_zz_377_] <= axi4_w_payload_data;
    end
  end

  assign _zz_271_ = int_ram_array_34[_zz_478_];
  assign _zz_272_ = int_ram_array_34[_zz_479_];
  always @ (posedge clk) begin
    if(_zz_545_) begin
      int_ram_array_35[_zz_379_] <= axi4_w_payload_data;
    end
  end

  assign _zz_273_ = int_ram_array_35[_zz_480_];
  assign _zz_274_ = int_ram_array_35[_zz_481_];
  always @ (posedge clk) begin
    if(_zz_546_) begin
      int_ram_array_36[_zz_381_] <= axi4_w_payload_data;
    end
  end

  assign _zz_275_ = int_ram_array_36[_zz_482_];
  assign _zz_276_ = int_ram_array_36[_zz_483_];
  always @ (posedge clk) begin
    if(_zz_547_) begin
      int_ram_array_37[_zz_383_] <= axi4_w_payload_data;
    end
  end

  assign _zz_277_ = int_ram_array_37[_zz_484_];
  assign _zz_278_ = int_ram_array_37[_zz_485_];
  always @ (posedge clk) begin
    if(_zz_548_) begin
      int_ram_array_38[_zz_385_] <= axi4_w_payload_data;
    end
  end

  assign _zz_279_ = int_ram_array_38[_zz_486_];
  assign _zz_280_ = int_ram_array_38[_zz_487_];
  always @ (posedge clk) begin
    if(_zz_549_) begin
      int_ram_array_39[_zz_387_] <= axi4_w_payload_data;
    end
  end

  assign _zz_281_ = int_ram_array_39[_zz_488_];
  assign _zz_282_ = int_ram_array_39[_zz_489_];
  always @ (posedge clk) begin
    if(_zz_550_) begin
      int_ram_array_40[_zz_389_] <= axi4_w_payload_data;
    end
  end

  assign _zz_283_ = int_ram_array_40[_zz_490_];
  assign _zz_284_ = int_ram_array_40[_zz_491_];
  always @ (posedge clk) begin
    if(_zz_551_) begin
      int_ram_array_41[_zz_391_] <= axi4_w_payload_data;
    end
  end

  assign _zz_285_ = int_ram_array_41[_zz_492_];
  assign _zz_286_ = int_ram_array_41[_zz_493_];
  always @ (posedge clk) begin
    if(_zz_552_) begin
      int_ram_array_42[_zz_393_] <= axi4_w_payload_data;
    end
  end

  assign _zz_287_ = int_ram_array_42[_zz_494_];
  assign _zz_288_ = int_ram_array_42[_zz_495_];
  always @ (posedge clk) begin
    if(_zz_553_) begin
      int_ram_array_43[_zz_395_] <= axi4_w_payload_data;
    end
  end

  assign _zz_289_ = int_ram_array_43[_zz_496_];
  assign _zz_290_ = int_ram_array_43[_zz_497_];
  always @ (posedge clk) begin
    if(_zz_554_) begin
      int_ram_array_44[_zz_397_] <= axi4_w_payload_data;
    end
  end

  assign _zz_291_ = int_ram_array_44[_zz_498_];
  assign _zz_292_ = int_ram_array_44[_zz_499_];
  always @ (posedge clk) begin
    if(_zz_555_) begin
      int_ram_array_45[_zz_399_] <= axi4_w_payload_data;
    end
  end

  assign _zz_293_ = int_ram_array_45[_zz_500_];
  assign _zz_294_ = int_ram_array_45[_zz_501_];
  always @ (posedge clk) begin
    if(_zz_556_) begin
      int_ram_array_46[_zz_401_] <= axi4_w_payload_data;
    end
  end

  assign _zz_295_ = int_ram_array_46[_zz_502_];
  assign _zz_296_ = int_ram_array_46[_zz_503_];
  always @ (posedge clk) begin
    if(_zz_557_) begin
      int_ram_array_47[_zz_403_] <= axi4_w_payload_data;
    end
  end

  assign _zz_297_ = int_ram_array_47[_zz_504_];
  assign _zz_298_ = int_ram_array_47[_zz_505_];
  always @ (posedge clk) begin
    if(_zz_558_) begin
      int_ram_array_48[_zz_405_] <= axi4_w_payload_data;
    end
  end

  assign _zz_299_ = int_ram_array_48[_zz_506_];
  assign _zz_300_ = int_ram_array_48[_zz_507_];
  always @ (posedge clk) begin
    if(_zz_559_) begin
      int_ram_array_49[_zz_407_] <= axi4_w_payload_data;
    end
  end

  assign _zz_301_ = int_ram_array_49[_zz_508_];
  assign _zz_302_ = int_ram_array_49[_zz_509_];
  always @(*) begin
    case(Axi4Incr_wrapCase)
      2'b00 : begin
        _zz_303_ = {Axi4Incr_base[11 : 1],Axi4Incr_baseIncr[0 : 0]};
      end
      2'b01 : begin
        _zz_303_ = {Axi4Incr_base[11 : 2],Axi4Incr_baseIncr[1 : 0]};
      end
      2'b10 : begin
        _zz_303_ = {Axi4Incr_base[11 : 3],Axi4Incr_baseIncr[2 : 0]};
      end
      default : begin
        _zz_303_ = {Axi4Incr_base[11 : 4],Axi4Incr_baseIncr[3 : 0]};
      end
    endcase
  end

  assign axi4_b_valid = axi4_w_valid;
  assign axi4_b_payload_id = aw_area_awid_r;
  assign axi4_b_payload_resp = (2'b00);
  assign axi4_aw_ready = 1'b1;
  assign axi4_w_ready = 1'b1;
  assign Axi4Incr_highCat = aw_area_awaddr_r[31 : 12];
  assign Axi4Incr_sizeValue = 1'b1;
  assign Axi4Incr_alignMask = 12'h0;
  assign Axi4Incr_base = (_zz_305_ & (~ Axi4Incr_alignMask));
  assign Axi4Incr_baseIncr = (Axi4Incr_base + _zz_306_);
  always @ (*) begin
    if((((aw_area_awlen_r & 8'h08) == 8'h08))) begin
        _zz_1_ = (2'b11);
    end else if((((aw_area_awlen_r & 8'h04) == 8'h04))) begin
        _zz_1_ = (2'b10);
    end else if((((aw_area_awlen_r & 8'h02) == 8'h02))) begin
        _zz_1_ = (2'b01);
    end else begin
        _zz_1_ = (2'b00);
    end
  end

  assign Axi4Incr_wrapCase = ((2'b00) + _zz_1_);
  always @ (*) begin
    case(axi4_aw_payload_burst)
      2'b00 : begin
        Axi4Incr_result = aw_area_awaddr_r;
      end
      2'b10 : begin
        Axi4Incr_result = {Axi4Incr_highCat,_zz_303_};
      end
      default : begin
        Axi4Incr_result = {Axi4Incr_highCat,Axi4Incr_baseIncr};
      end
    endcase
  end

  assign io_impulse_out_valid = transfer_done_1_;
  always @ (*) begin
    current_mem_addr_willIncrement = 1'b0;
    if((transfer_done_1_ || _zz_2_))begin
      current_mem_addr_willIncrement = 1'b1;
      current_mem_addr_willIncrement = 1'b1;
    end
  end

  assign current_mem_addr_willClear = 1'b0;
  assign current_mem_addr_willOverflowIfInc = (current_mem_addr_value == 14'h3fff);
  assign current_mem_addr_willOverflow = (current_mem_addr_willOverflowIfInc && current_mem_addr_willIncrement);
  always @ (*) begin
    current_mem_addr_valueNext = (current_mem_addr_value + _zz_409_);
    if(current_mem_addr_willClear)begin
      current_mem_addr_valueNext = 14'h0;
    end
  end

  assign _zz_3_ = (current_mem_addr_value + 14'h0);
  assign _zz_4_ = _zz_203_;
  assign io_impulse_out_payload_0_0_real = _zz_4_[15 : 0];
  assign io_impulse_out_payload_0_0_imag = _zz_4_[31 : 16];
  assign _zz_5_ = (current_mem_addr_value + 14'h0001);
  assign _zz_6_ = _zz_204_;
  assign io_impulse_out_payload_0_1_real = _zz_6_[15 : 0];
  assign io_impulse_out_payload_0_1_imag = _zz_6_[31 : 16];
  assign _zz_7_ = (current_mem_addr_value + 14'h0);
  assign _zz_8_ = _zz_205_;
  assign io_impulse_out_payload_1_0_real = _zz_8_[15 : 0];
  assign io_impulse_out_payload_1_0_imag = _zz_8_[31 : 16];
  assign _zz_9_ = (current_mem_addr_value + 14'h0001);
  assign _zz_10_ = _zz_206_;
  assign io_impulse_out_payload_1_1_real = _zz_10_[15 : 0];
  assign io_impulse_out_payload_1_1_imag = _zz_10_[31 : 16];
  assign _zz_11_ = (current_mem_addr_value + 14'h0);
  assign _zz_12_ = _zz_207_;
  assign io_impulse_out_payload_2_0_real = _zz_12_[15 : 0];
  assign io_impulse_out_payload_2_0_imag = _zz_12_[31 : 16];
  assign _zz_13_ = (current_mem_addr_value + 14'h0001);
  assign _zz_14_ = _zz_208_;
  assign io_impulse_out_payload_2_1_real = _zz_14_[15 : 0];
  assign io_impulse_out_payload_2_1_imag = _zz_14_[31 : 16];
  assign _zz_15_ = (current_mem_addr_value + 14'h0);
  assign _zz_16_ = _zz_209_;
  assign io_impulse_out_payload_3_0_real = _zz_16_[15 : 0];
  assign io_impulse_out_payload_3_0_imag = _zz_16_[31 : 16];
  assign _zz_17_ = (current_mem_addr_value + 14'h0001);
  assign _zz_18_ = _zz_210_;
  assign io_impulse_out_payload_3_1_real = _zz_18_[15 : 0];
  assign io_impulse_out_payload_3_1_imag = _zz_18_[31 : 16];
  assign _zz_19_ = (current_mem_addr_value + 14'h0);
  assign _zz_20_ = _zz_211_;
  assign io_impulse_out_payload_4_0_real = _zz_20_[15 : 0];
  assign io_impulse_out_payload_4_0_imag = _zz_20_[31 : 16];
  assign _zz_21_ = (current_mem_addr_value + 14'h0001);
  assign _zz_22_ = _zz_212_;
  assign io_impulse_out_payload_4_1_real = _zz_22_[15 : 0];
  assign io_impulse_out_payload_4_1_imag = _zz_22_[31 : 16];
  assign _zz_23_ = (current_mem_addr_value + 14'h0);
  assign _zz_24_ = _zz_213_;
  assign io_impulse_out_payload_5_0_real = _zz_24_[15 : 0];
  assign io_impulse_out_payload_5_0_imag = _zz_24_[31 : 16];
  assign _zz_25_ = (current_mem_addr_value + 14'h0001);
  assign _zz_26_ = _zz_214_;
  assign io_impulse_out_payload_5_1_real = _zz_26_[15 : 0];
  assign io_impulse_out_payload_5_1_imag = _zz_26_[31 : 16];
  assign _zz_27_ = (current_mem_addr_value + 14'h0);
  assign _zz_28_ = _zz_215_;
  assign io_impulse_out_payload_6_0_real = _zz_28_[15 : 0];
  assign io_impulse_out_payload_6_0_imag = _zz_28_[31 : 16];
  assign _zz_29_ = (current_mem_addr_value + 14'h0001);
  assign _zz_30_ = _zz_216_;
  assign io_impulse_out_payload_6_1_real = _zz_30_[15 : 0];
  assign io_impulse_out_payload_6_1_imag = _zz_30_[31 : 16];
  assign _zz_31_ = (current_mem_addr_value + 14'h0);
  assign _zz_32_ = _zz_217_;
  assign io_impulse_out_payload_7_0_real = _zz_32_[15 : 0];
  assign io_impulse_out_payload_7_0_imag = _zz_32_[31 : 16];
  assign _zz_33_ = (current_mem_addr_value + 14'h0001);
  assign _zz_34_ = _zz_218_;
  assign io_impulse_out_payload_7_1_real = _zz_34_[15 : 0];
  assign io_impulse_out_payload_7_1_imag = _zz_34_[31 : 16];
  assign _zz_35_ = (current_mem_addr_value + 14'h0);
  assign _zz_36_ = _zz_219_;
  assign io_impulse_out_payload_8_0_real = _zz_36_[15 : 0];
  assign io_impulse_out_payload_8_0_imag = _zz_36_[31 : 16];
  assign _zz_37_ = (current_mem_addr_value + 14'h0001);
  assign _zz_38_ = _zz_220_;
  assign io_impulse_out_payload_8_1_real = _zz_38_[15 : 0];
  assign io_impulse_out_payload_8_1_imag = _zz_38_[31 : 16];
  assign _zz_39_ = (current_mem_addr_value + 14'h0);
  assign _zz_40_ = _zz_221_;
  assign io_impulse_out_payload_9_0_real = _zz_40_[15 : 0];
  assign io_impulse_out_payload_9_0_imag = _zz_40_[31 : 16];
  assign _zz_41_ = (current_mem_addr_value + 14'h0001);
  assign _zz_42_ = _zz_222_;
  assign io_impulse_out_payload_9_1_real = _zz_42_[15 : 0];
  assign io_impulse_out_payload_9_1_imag = _zz_42_[31 : 16];
  assign _zz_43_ = (current_mem_addr_value + 14'h0);
  assign _zz_44_ = _zz_223_;
  assign io_impulse_out_payload_10_0_real = _zz_44_[15 : 0];
  assign io_impulse_out_payload_10_0_imag = _zz_44_[31 : 16];
  assign _zz_45_ = (current_mem_addr_value + 14'h0001);
  assign _zz_46_ = _zz_224_;
  assign io_impulse_out_payload_10_1_real = _zz_46_[15 : 0];
  assign io_impulse_out_payload_10_1_imag = _zz_46_[31 : 16];
  assign _zz_47_ = (current_mem_addr_value + 14'h0);
  assign _zz_48_ = _zz_225_;
  assign io_impulse_out_payload_11_0_real = _zz_48_[15 : 0];
  assign io_impulse_out_payload_11_0_imag = _zz_48_[31 : 16];
  assign _zz_49_ = (current_mem_addr_value + 14'h0001);
  assign _zz_50_ = _zz_226_;
  assign io_impulse_out_payload_11_1_real = _zz_50_[15 : 0];
  assign io_impulse_out_payload_11_1_imag = _zz_50_[31 : 16];
  assign _zz_51_ = (current_mem_addr_value + 14'h0);
  assign _zz_52_ = _zz_227_;
  assign io_impulse_out_payload_12_0_real = _zz_52_[15 : 0];
  assign io_impulse_out_payload_12_0_imag = _zz_52_[31 : 16];
  assign _zz_53_ = (current_mem_addr_value + 14'h0001);
  assign _zz_54_ = _zz_228_;
  assign io_impulse_out_payload_12_1_real = _zz_54_[15 : 0];
  assign io_impulse_out_payload_12_1_imag = _zz_54_[31 : 16];
  assign _zz_55_ = (current_mem_addr_value + 14'h0);
  assign _zz_56_ = _zz_229_;
  assign io_impulse_out_payload_13_0_real = _zz_56_[15 : 0];
  assign io_impulse_out_payload_13_0_imag = _zz_56_[31 : 16];
  assign _zz_57_ = (current_mem_addr_value + 14'h0001);
  assign _zz_58_ = _zz_230_;
  assign io_impulse_out_payload_13_1_real = _zz_58_[15 : 0];
  assign io_impulse_out_payload_13_1_imag = _zz_58_[31 : 16];
  assign _zz_59_ = (current_mem_addr_value + 14'h0);
  assign _zz_60_ = _zz_231_;
  assign io_impulse_out_payload_14_0_real = _zz_60_[15 : 0];
  assign io_impulse_out_payload_14_0_imag = _zz_60_[31 : 16];
  assign _zz_61_ = (current_mem_addr_value + 14'h0001);
  assign _zz_62_ = _zz_232_;
  assign io_impulse_out_payload_14_1_real = _zz_62_[15 : 0];
  assign io_impulse_out_payload_14_1_imag = _zz_62_[31 : 16];
  assign _zz_63_ = (current_mem_addr_value + 14'h0);
  assign _zz_64_ = _zz_233_;
  assign io_impulse_out_payload_15_0_real = _zz_64_[15 : 0];
  assign io_impulse_out_payload_15_0_imag = _zz_64_[31 : 16];
  assign _zz_65_ = (current_mem_addr_value + 14'h0001);
  assign _zz_66_ = _zz_234_;
  assign io_impulse_out_payload_15_1_real = _zz_66_[15 : 0];
  assign io_impulse_out_payload_15_1_imag = _zz_66_[31 : 16];
  assign _zz_67_ = (current_mem_addr_value + 14'h0);
  assign _zz_68_ = _zz_235_;
  assign io_impulse_out_payload_16_0_real = _zz_68_[15 : 0];
  assign io_impulse_out_payload_16_0_imag = _zz_68_[31 : 16];
  assign _zz_69_ = (current_mem_addr_value + 14'h0001);
  assign _zz_70_ = _zz_236_;
  assign io_impulse_out_payload_16_1_real = _zz_70_[15 : 0];
  assign io_impulse_out_payload_16_1_imag = _zz_70_[31 : 16];
  assign _zz_71_ = (current_mem_addr_value + 14'h0);
  assign _zz_72_ = _zz_237_;
  assign io_impulse_out_payload_17_0_real = _zz_72_[15 : 0];
  assign io_impulse_out_payload_17_0_imag = _zz_72_[31 : 16];
  assign _zz_73_ = (current_mem_addr_value + 14'h0001);
  assign _zz_74_ = _zz_238_;
  assign io_impulse_out_payload_17_1_real = _zz_74_[15 : 0];
  assign io_impulse_out_payload_17_1_imag = _zz_74_[31 : 16];
  assign _zz_75_ = (current_mem_addr_value + 14'h0);
  assign _zz_76_ = _zz_239_;
  assign io_impulse_out_payload_18_0_real = _zz_76_[15 : 0];
  assign io_impulse_out_payload_18_0_imag = _zz_76_[31 : 16];
  assign _zz_77_ = (current_mem_addr_value + 14'h0001);
  assign _zz_78_ = _zz_240_;
  assign io_impulse_out_payload_18_1_real = _zz_78_[15 : 0];
  assign io_impulse_out_payload_18_1_imag = _zz_78_[31 : 16];
  assign _zz_79_ = (current_mem_addr_value + 14'h0);
  assign _zz_80_ = _zz_241_;
  assign io_impulse_out_payload_19_0_real = _zz_80_[15 : 0];
  assign io_impulse_out_payload_19_0_imag = _zz_80_[31 : 16];
  assign _zz_81_ = (current_mem_addr_value + 14'h0001);
  assign _zz_82_ = _zz_242_;
  assign io_impulse_out_payload_19_1_real = _zz_82_[15 : 0];
  assign io_impulse_out_payload_19_1_imag = _zz_82_[31 : 16];
  assign _zz_83_ = (current_mem_addr_value + 14'h0);
  assign _zz_84_ = _zz_243_;
  assign io_impulse_out_payload_20_0_real = _zz_84_[15 : 0];
  assign io_impulse_out_payload_20_0_imag = _zz_84_[31 : 16];
  assign _zz_85_ = (current_mem_addr_value + 14'h0001);
  assign _zz_86_ = _zz_244_;
  assign io_impulse_out_payload_20_1_real = _zz_86_[15 : 0];
  assign io_impulse_out_payload_20_1_imag = _zz_86_[31 : 16];
  assign _zz_87_ = (current_mem_addr_value + 14'h0);
  assign _zz_88_ = _zz_245_;
  assign io_impulse_out_payload_21_0_real = _zz_88_[15 : 0];
  assign io_impulse_out_payload_21_0_imag = _zz_88_[31 : 16];
  assign _zz_89_ = (current_mem_addr_value + 14'h0001);
  assign _zz_90_ = _zz_246_;
  assign io_impulse_out_payload_21_1_real = _zz_90_[15 : 0];
  assign io_impulse_out_payload_21_1_imag = _zz_90_[31 : 16];
  assign _zz_91_ = (current_mem_addr_value + 14'h0);
  assign _zz_92_ = _zz_247_;
  assign io_impulse_out_payload_22_0_real = _zz_92_[15 : 0];
  assign io_impulse_out_payload_22_0_imag = _zz_92_[31 : 16];
  assign _zz_93_ = (current_mem_addr_value + 14'h0001);
  assign _zz_94_ = _zz_248_;
  assign io_impulse_out_payload_22_1_real = _zz_94_[15 : 0];
  assign io_impulse_out_payload_22_1_imag = _zz_94_[31 : 16];
  assign _zz_95_ = (current_mem_addr_value + 14'h0);
  assign _zz_96_ = _zz_249_;
  assign io_impulse_out_payload_23_0_real = _zz_96_[15 : 0];
  assign io_impulse_out_payload_23_0_imag = _zz_96_[31 : 16];
  assign _zz_97_ = (current_mem_addr_value + 14'h0001);
  assign _zz_98_ = _zz_250_;
  assign io_impulse_out_payload_23_1_real = _zz_98_[15 : 0];
  assign io_impulse_out_payload_23_1_imag = _zz_98_[31 : 16];
  assign _zz_99_ = (current_mem_addr_value + 14'h0);
  assign _zz_100_ = _zz_251_;
  assign io_impulse_out_payload_24_0_real = _zz_100_[15 : 0];
  assign io_impulse_out_payload_24_0_imag = _zz_100_[31 : 16];
  assign _zz_101_ = (current_mem_addr_value + 14'h0001);
  assign _zz_102_ = _zz_252_;
  assign io_impulse_out_payload_24_1_real = _zz_102_[15 : 0];
  assign io_impulse_out_payload_24_1_imag = _zz_102_[31 : 16];
  assign _zz_103_ = (current_mem_addr_value + 14'h0);
  assign _zz_104_ = _zz_253_;
  assign io_impulse_out_payload_25_0_real = _zz_104_[15 : 0];
  assign io_impulse_out_payload_25_0_imag = _zz_104_[31 : 16];
  assign _zz_105_ = (current_mem_addr_value + 14'h0001);
  assign _zz_106_ = _zz_254_;
  assign io_impulse_out_payload_25_1_real = _zz_106_[15 : 0];
  assign io_impulse_out_payload_25_1_imag = _zz_106_[31 : 16];
  assign _zz_107_ = (current_mem_addr_value + 14'h0);
  assign _zz_108_ = _zz_255_;
  assign io_impulse_out_payload_26_0_real = _zz_108_[15 : 0];
  assign io_impulse_out_payload_26_0_imag = _zz_108_[31 : 16];
  assign _zz_109_ = (current_mem_addr_value + 14'h0001);
  assign _zz_110_ = _zz_256_;
  assign io_impulse_out_payload_26_1_real = _zz_110_[15 : 0];
  assign io_impulse_out_payload_26_1_imag = _zz_110_[31 : 16];
  assign _zz_111_ = (current_mem_addr_value + 14'h0);
  assign _zz_112_ = _zz_257_;
  assign io_impulse_out_payload_27_0_real = _zz_112_[15 : 0];
  assign io_impulse_out_payload_27_0_imag = _zz_112_[31 : 16];
  assign _zz_113_ = (current_mem_addr_value + 14'h0001);
  assign _zz_114_ = _zz_258_;
  assign io_impulse_out_payload_27_1_real = _zz_114_[15 : 0];
  assign io_impulse_out_payload_27_1_imag = _zz_114_[31 : 16];
  assign _zz_115_ = (current_mem_addr_value + 14'h0);
  assign _zz_116_ = _zz_259_;
  assign io_impulse_out_payload_28_0_real = _zz_116_[15 : 0];
  assign io_impulse_out_payload_28_0_imag = _zz_116_[31 : 16];
  assign _zz_117_ = (current_mem_addr_value + 14'h0001);
  assign _zz_118_ = _zz_260_;
  assign io_impulse_out_payload_28_1_real = _zz_118_[15 : 0];
  assign io_impulse_out_payload_28_1_imag = _zz_118_[31 : 16];
  assign _zz_119_ = (current_mem_addr_value + 14'h0);
  assign _zz_120_ = _zz_261_;
  assign io_impulse_out_payload_29_0_real = _zz_120_[15 : 0];
  assign io_impulse_out_payload_29_0_imag = _zz_120_[31 : 16];
  assign _zz_121_ = (current_mem_addr_value + 14'h0001);
  assign _zz_122_ = _zz_262_;
  assign io_impulse_out_payload_29_1_real = _zz_122_[15 : 0];
  assign io_impulse_out_payload_29_1_imag = _zz_122_[31 : 16];
  assign _zz_123_ = (current_mem_addr_value + 14'h0);
  assign _zz_124_ = _zz_263_;
  assign io_impulse_out_payload_30_0_real = _zz_124_[15 : 0];
  assign io_impulse_out_payload_30_0_imag = _zz_124_[31 : 16];
  assign _zz_125_ = (current_mem_addr_value + 14'h0001);
  assign _zz_126_ = _zz_264_;
  assign io_impulse_out_payload_30_1_real = _zz_126_[15 : 0];
  assign io_impulse_out_payload_30_1_imag = _zz_126_[31 : 16];
  assign _zz_127_ = (current_mem_addr_value + 14'h0);
  assign _zz_128_ = _zz_265_;
  assign io_impulse_out_payload_31_0_real = _zz_128_[15 : 0];
  assign io_impulse_out_payload_31_0_imag = _zz_128_[31 : 16];
  assign _zz_129_ = (current_mem_addr_value + 14'h0001);
  assign _zz_130_ = _zz_266_;
  assign io_impulse_out_payload_31_1_real = _zz_130_[15 : 0];
  assign io_impulse_out_payload_31_1_imag = _zz_130_[31 : 16];
  assign _zz_131_ = (current_mem_addr_value + 14'h0);
  assign _zz_132_ = _zz_267_;
  assign io_impulse_out_payload_32_0_real = _zz_132_[15 : 0];
  assign io_impulse_out_payload_32_0_imag = _zz_132_[31 : 16];
  assign _zz_133_ = (current_mem_addr_value + 14'h0001);
  assign _zz_134_ = _zz_268_;
  assign io_impulse_out_payload_32_1_real = _zz_134_[15 : 0];
  assign io_impulse_out_payload_32_1_imag = _zz_134_[31 : 16];
  assign _zz_135_ = (current_mem_addr_value + 14'h0);
  assign _zz_136_ = _zz_269_;
  assign io_impulse_out_payload_33_0_real = _zz_136_[15 : 0];
  assign io_impulse_out_payload_33_0_imag = _zz_136_[31 : 16];
  assign _zz_137_ = (current_mem_addr_value + 14'h0001);
  assign _zz_138_ = _zz_270_;
  assign io_impulse_out_payload_33_1_real = _zz_138_[15 : 0];
  assign io_impulse_out_payload_33_1_imag = _zz_138_[31 : 16];
  assign _zz_139_ = (current_mem_addr_value + 14'h0);
  assign _zz_140_ = _zz_271_;
  assign io_impulse_out_payload_34_0_real = _zz_140_[15 : 0];
  assign io_impulse_out_payload_34_0_imag = _zz_140_[31 : 16];
  assign _zz_141_ = (current_mem_addr_value + 14'h0001);
  assign _zz_142_ = _zz_272_;
  assign io_impulse_out_payload_34_1_real = _zz_142_[15 : 0];
  assign io_impulse_out_payload_34_1_imag = _zz_142_[31 : 16];
  assign _zz_143_ = (current_mem_addr_value + 14'h0);
  assign _zz_144_ = _zz_273_;
  assign io_impulse_out_payload_35_0_real = _zz_144_[15 : 0];
  assign io_impulse_out_payload_35_0_imag = _zz_144_[31 : 16];
  assign _zz_145_ = (current_mem_addr_value + 14'h0001);
  assign _zz_146_ = _zz_274_;
  assign io_impulse_out_payload_35_1_real = _zz_146_[15 : 0];
  assign io_impulse_out_payload_35_1_imag = _zz_146_[31 : 16];
  assign _zz_147_ = (current_mem_addr_value + 14'h0);
  assign _zz_148_ = _zz_275_;
  assign io_impulse_out_payload_36_0_real = _zz_148_[15 : 0];
  assign io_impulse_out_payload_36_0_imag = _zz_148_[31 : 16];
  assign _zz_149_ = (current_mem_addr_value + 14'h0001);
  assign _zz_150_ = _zz_276_;
  assign io_impulse_out_payload_36_1_real = _zz_150_[15 : 0];
  assign io_impulse_out_payload_36_1_imag = _zz_150_[31 : 16];
  assign _zz_151_ = (current_mem_addr_value + 14'h0);
  assign _zz_152_ = _zz_277_;
  assign io_impulse_out_payload_37_0_real = _zz_152_[15 : 0];
  assign io_impulse_out_payload_37_0_imag = _zz_152_[31 : 16];
  assign _zz_153_ = (current_mem_addr_value + 14'h0001);
  assign _zz_154_ = _zz_278_;
  assign io_impulse_out_payload_37_1_real = _zz_154_[15 : 0];
  assign io_impulse_out_payload_37_1_imag = _zz_154_[31 : 16];
  assign _zz_155_ = (current_mem_addr_value + 14'h0);
  assign _zz_156_ = _zz_279_;
  assign io_impulse_out_payload_38_0_real = _zz_156_[15 : 0];
  assign io_impulse_out_payload_38_0_imag = _zz_156_[31 : 16];
  assign _zz_157_ = (current_mem_addr_value + 14'h0001);
  assign _zz_158_ = _zz_280_;
  assign io_impulse_out_payload_38_1_real = _zz_158_[15 : 0];
  assign io_impulse_out_payload_38_1_imag = _zz_158_[31 : 16];
  assign _zz_159_ = (current_mem_addr_value + 14'h0);
  assign _zz_160_ = _zz_281_;
  assign io_impulse_out_payload_39_0_real = _zz_160_[15 : 0];
  assign io_impulse_out_payload_39_0_imag = _zz_160_[31 : 16];
  assign _zz_161_ = (current_mem_addr_value + 14'h0001);
  assign _zz_162_ = _zz_282_;
  assign io_impulse_out_payload_39_1_real = _zz_162_[15 : 0];
  assign io_impulse_out_payload_39_1_imag = _zz_162_[31 : 16];
  assign _zz_163_ = (current_mem_addr_value + 14'h0);
  assign _zz_164_ = _zz_283_;
  assign io_impulse_out_payload_40_0_real = _zz_164_[15 : 0];
  assign io_impulse_out_payload_40_0_imag = _zz_164_[31 : 16];
  assign _zz_165_ = (current_mem_addr_value + 14'h0001);
  assign _zz_166_ = _zz_284_;
  assign io_impulse_out_payload_40_1_real = _zz_166_[15 : 0];
  assign io_impulse_out_payload_40_1_imag = _zz_166_[31 : 16];
  assign _zz_167_ = (current_mem_addr_value + 14'h0);
  assign _zz_168_ = _zz_285_;
  assign io_impulse_out_payload_41_0_real = _zz_168_[15 : 0];
  assign io_impulse_out_payload_41_0_imag = _zz_168_[31 : 16];
  assign _zz_169_ = (current_mem_addr_value + 14'h0001);
  assign _zz_170_ = _zz_286_;
  assign io_impulse_out_payload_41_1_real = _zz_170_[15 : 0];
  assign io_impulse_out_payload_41_1_imag = _zz_170_[31 : 16];
  assign _zz_171_ = (current_mem_addr_value + 14'h0);
  assign _zz_172_ = _zz_287_;
  assign io_impulse_out_payload_42_0_real = _zz_172_[15 : 0];
  assign io_impulse_out_payload_42_0_imag = _zz_172_[31 : 16];
  assign _zz_173_ = (current_mem_addr_value + 14'h0001);
  assign _zz_174_ = _zz_288_;
  assign io_impulse_out_payload_42_1_real = _zz_174_[15 : 0];
  assign io_impulse_out_payload_42_1_imag = _zz_174_[31 : 16];
  assign _zz_175_ = (current_mem_addr_value + 14'h0);
  assign _zz_176_ = _zz_289_;
  assign io_impulse_out_payload_43_0_real = _zz_176_[15 : 0];
  assign io_impulse_out_payload_43_0_imag = _zz_176_[31 : 16];
  assign _zz_177_ = (current_mem_addr_value + 14'h0001);
  assign _zz_178_ = _zz_290_;
  assign io_impulse_out_payload_43_1_real = _zz_178_[15 : 0];
  assign io_impulse_out_payload_43_1_imag = _zz_178_[31 : 16];
  assign _zz_179_ = (current_mem_addr_value + 14'h0);
  assign _zz_180_ = _zz_291_;
  assign io_impulse_out_payload_44_0_real = _zz_180_[15 : 0];
  assign io_impulse_out_payload_44_0_imag = _zz_180_[31 : 16];
  assign _zz_181_ = (current_mem_addr_value + 14'h0001);
  assign _zz_182_ = _zz_292_;
  assign io_impulse_out_payload_44_1_real = _zz_182_[15 : 0];
  assign io_impulse_out_payload_44_1_imag = _zz_182_[31 : 16];
  assign _zz_183_ = (current_mem_addr_value + 14'h0);
  assign _zz_184_ = _zz_293_;
  assign io_impulse_out_payload_45_0_real = _zz_184_[15 : 0];
  assign io_impulse_out_payload_45_0_imag = _zz_184_[31 : 16];
  assign _zz_185_ = (current_mem_addr_value + 14'h0001);
  assign _zz_186_ = _zz_294_;
  assign io_impulse_out_payload_45_1_real = _zz_186_[15 : 0];
  assign io_impulse_out_payload_45_1_imag = _zz_186_[31 : 16];
  assign _zz_187_ = (current_mem_addr_value + 14'h0);
  assign _zz_188_ = _zz_295_;
  assign io_impulse_out_payload_46_0_real = _zz_188_[15 : 0];
  assign io_impulse_out_payload_46_0_imag = _zz_188_[31 : 16];
  assign _zz_189_ = (current_mem_addr_value + 14'h0001);
  assign _zz_190_ = _zz_296_;
  assign io_impulse_out_payload_46_1_real = _zz_190_[15 : 0];
  assign io_impulse_out_payload_46_1_imag = _zz_190_[31 : 16];
  assign _zz_191_ = (current_mem_addr_value + 14'h0);
  assign _zz_192_ = _zz_297_;
  assign io_impulse_out_payload_47_0_real = _zz_192_[15 : 0];
  assign io_impulse_out_payload_47_0_imag = _zz_192_[31 : 16];
  assign _zz_193_ = (current_mem_addr_value + 14'h0001);
  assign _zz_194_ = _zz_298_;
  assign io_impulse_out_payload_47_1_real = _zz_194_[15 : 0];
  assign io_impulse_out_payload_47_1_imag = _zz_194_[31 : 16];
  assign _zz_195_ = (current_mem_addr_value + 14'h0);
  assign _zz_196_ = _zz_299_;
  assign io_impulse_out_payload_48_0_real = _zz_196_[15 : 0];
  assign io_impulse_out_payload_48_0_imag = _zz_196_[31 : 16];
  assign _zz_197_ = (current_mem_addr_value + 14'h0001);
  assign _zz_198_ = _zz_300_;
  assign io_impulse_out_payload_48_1_real = _zz_198_[15 : 0];
  assign io_impulse_out_payload_48_1_imag = _zz_198_[31 : 16];
  assign _zz_199_ = (current_mem_addr_value + 14'h0);
  assign _zz_200_ = _zz_301_;
  assign io_impulse_out_payload_49_0_real = _zz_200_[15 : 0];
  assign io_impulse_out_payload_49_0_imag = _zz_200_[31 : 16];
  assign _zz_201_ = (current_mem_addr_value + 14'h0001);
  assign _zz_202_ = _zz_302_;
  assign io_impulse_out_payload_49_1_real = _zz_202_[15 : 0];
  assign io_impulse_out_payload_49_1_imag = _zz_202_[31 : 16];
  always @ (posedge clk) begin
    if(axi4_aw_valid)begin
      aw_area_awaddr_r <= axi4_aw_payload_addr;
      aw_area_awlen_r <= axi4_aw_payload_len;
      aw_area_awsize_r <= axi4_aw_payload_size;
      aw_area_awid_r <= axi4_aw_payload_id;
    end
    if(axi4_w_valid)begin
      transfer_done_1_ <= (((32'h00000c80 <= load_data_area_current_addr) && (load_data_area_current_addr < 32'h00000c80)) ? axi4_w_payload_data_regNext[0] : _zz_307_[0]);
    end
  end

  always @ (posedge clk or posedge reset) begin
    if (reset) begin
      load_data_area_current_addr <= 32'h0;
      current_mem_addr_value <= 14'h0;
      _zz_2_ <= 1'b0;
    end else begin
      if(axi4_w_valid)begin
        load_data_area_current_addr <= Axi4Incr_result;
      end
      current_mem_addr_value <= current_mem_addr_valueNext;
      if(transfer_done_1_)begin
        _zz_2_ <= 1'b1;
      end else begin
        if(current_mem_addr_willOverflow)begin
          _zz_2_ <= 1'b0;
        end
      end
    end
  end

  always @ (posedge clk) begin
    axi4_w_payload_data_regNext <= axi4_w_payload_data;
  end


endmodule
