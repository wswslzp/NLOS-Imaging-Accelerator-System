// Generator : SpinalHDL v1.4.1    git head : 99d6d471af204b6d7d9f63fae58757e9d3c7b944
// Component : MyFFT
// Git hash  : 2a34fe18f42a28946060dbf37f9913e1060dc674



module MyFFT (
  input               io_data_in_valid,
  input      [15:0]   io_data_in_payload_0_real,
  input      [15:0]   io_data_in_payload_0_imag,
  input      [15:0]   io_data_in_payload_1_real,
  input      [15:0]   io_data_in_payload_1_imag,
  input      [15:0]   io_data_in_payload_2_real,
  input      [15:0]   io_data_in_payload_2_imag,
  input      [15:0]   io_data_in_payload_3_real,
  input      [15:0]   io_data_in_payload_3_imag,
  input      [15:0]   io_data_in_payload_4_real,
  input      [15:0]   io_data_in_payload_4_imag,
  input      [15:0]   io_data_in_payload_5_real,
  input      [15:0]   io_data_in_payload_5_imag,
  input      [15:0]   io_data_in_payload_6_real,
  input      [15:0]   io_data_in_payload_6_imag,
  input      [15:0]   io_data_in_payload_7_real,
  input      [15:0]   io_data_in_payload_7_imag,
  input      [15:0]   io_data_in_payload_8_real,
  input      [15:0]   io_data_in_payload_8_imag,
  input      [15:0]   io_data_in_payload_9_real,
  input      [15:0]   io_data_in_payload_9_imag,
  input      [15:0]   io_data_in_payload_10_real,
  input      [15:0]   io_data_in_payload_10_imag,
  input      [15:0]   io_data_in_payload_11_real,
  input      [15:0]   io_data_in_payload_11_imag,
  input      [15:0]   io_data_in_payload_12_real,
  input      [15:0]   io_data_in_payload_12_imag,
  input      [15:0]   io_data_in_payload_13_real,
  input      [15:0]   io_data_in_payload_13_imag,
  input      [15:0]   io_data_in_payload_14_real,
  input      [15:0]   io_data_in_payload_14_imag,
  input      [15:0]   io_data_in_payload_15_real,
  input      [15:0]   io_data_in_payload_15_imag,
  input      [15:0]   io_data_in_payload_16_real,
  input      [15:0]   io_data_in_payload_16_imag,
  input      [15:0]   io_data_in_payload_17_real,
  input      [15:0]   io_data_in_payload_17_imag,
  input      [15:0]   io_data_in_payload_18_real,
  input      [15:0]   io_data_in_payload_18_imag,
  input      [15:0]   io_data_in_payload_19_real,
  input      [15:0]   io_data_in_payload_19_imag,
  input      [15:0]   io_data_in_payload_20_real,
  input      [15:0]   io_data_in_payload_20_imag,
  input      [15:0]   io_data_in_payload_21_real,
  input      [15:0]   io_data_in_payload_21_imag,
  input      [15:0]   io_data_in_payload_22_real,
  input      [15:0]   io_data_in_payload_22_imag,
  input      [15:0]   io_data_in_payload_23_real,
  input      [15:0]   io_data_in_payload_23_imag,
  input      [15:0]   io_data_in_payload_24_real,
  input      [15:0]   io_data_in_payload_24_imag,
  input      [15:0]   io_data_in_payload_25_real,
  input      [15:0]   io_data_in_payload_25_imag,
  input      [15:0]   io_data_in_payload_26_real,
  input      [15:0]   io_data_in_payload_26_imag,
  input      [15:0]   io_data_in_payload_27_real,
  input      [15:0]   io_data_in_payload_27_imag,
  input      [15:0]   io_data_in_payload_28_real,
  input      [15:0]   io_data_in_payload_28_imag,
  input      [15:0]   io_data_in_payload_29_real,
  input      [15:0]   io_data_in_payload_29_imag,
  input      [15:0]   io_data_in_payload_30_real,
  input      [15:0]   io_data_in_payload_30_imag,
  input      [15:0]   io_data_in_payload_31_real,
  input      [15:0]   io_data_in_payload_31_imag,
  input      [15:0]   io_data_in_payload_32_real,
  input      [15:0]   io_data_in_payload_32_imag,
  input      [15:0]   io_data_in_payload_33_real,
  input      [15:0]   io_data_in_payload_33_imag,
  input      [15:0]   io_data_in_payload_34_real,
  input      [15:0]   io_data_in_payload_34_imag,
  input      [15:0]   io_data_in_payload_35_real,
  input      [15:0]   io_data_in_payload_35_imag,
  input      [15:0]   io_data_in_payload_36_real,
  input      [15:0]   io_data_in_payload_36_imag,
  input      [15:0]   io_data_in_payload_37_real,
  input      [15:0]   io_data_in_payload_37_imag,
  input      [15:0]   io_data_in_payload_38_real,
  input      [15:0]   io_data_in_payload_38_imag,
  input      [15:0]   io_data_in_payload_39_real,
  input      [15:0]   io_data_in_payload_39_imag,
  input      [15:0]   io_data_in_payload_40_real,
  input      [15:0]   io_data_in_payload_40_imag,
  input      [15:0]   io_data_in_payload_41_real,
  input      [15:0]   io_data_in_payload_41_imag,
  input      [15:0]   io_data_in_payload_42_real,
  input      [15:0]   io_data_in_payload_42_imag,
  input      [15:0]   io_data_in_payload_43_real,
  input      [15:0]   io_data_in_payload_43_imag,
  input      [15:0]   io_data_in_payload_44_real,
  input      [15:0]   io_data_in_payload_44_imag,
  input      [15:0]   io_data_in_payload_45_real,
  input      [15:0]   io_data_in_payload_45_imag,
  input      [15:0]   io_data_in_payload_46_real,
  input      [15:0]   io_data_in_payload_46_imag,
  input      [15:0]   io_data_in_payload_47_real,
  input      [15:0]   io_data_in_payload_47_imag,
  input      [15:0]   io_data_in_payload_48_real,
  input      [15:0]   io_data_in_payload_48_imag,
  input      [15:0]   io_data_in_payload_49_real,
  input      [15:0]   io_data_in_payload_49_imag,
  input      [15:0]   io_data_in_payload_50_real,
  input      [15:0]   io_data_in_payload_50_imag,
  input      [15:0]   io_data_in_payload_51_real,
  input      [15:0]   io_data_in_payload_51_imag,
  input      [15:0]   io_data_in_payload_52_real,
  input      [15:0]   io_data_in_payload_52_imag,
  input      [15:0]   io_data_in_payload_53_real,
  input      [15:0]   io_data_in_payload_53_imag,
  input      [15:0]   io_data_in_payload_54_real,
  input      [15:0]   io_data_in_payload_54_imag,
  input      [15:0]   io_data_in_payload_55_real,
  input      [15:0]   io_data_in_payload_55_imag,
  input      [15:0]   io_data_in_payload_56_real,
  input      [15:0]   io_data_in_payload_56_imag,
  input      [15:0]   io_data_in_payload_57_real,
  input      [15:0]   io_data_in_payload_57_imag,
  input      [15:0]   io_data_in_payload_58_real,
  input      [15:0]   io_data_in_payload_58_imag,
  input      [15:0]   io_data_in_payload_59_real,
  input      [15:0]   io_data_in_payload_59_imag,
  input      [15:0]   io_data_in_payload_60_real,
  input      [15:0]   io_data_in_payload_60_imag,
  input      [15:0]   io_data_in_payload_61_real,
  input      [15:0]   io_data_in_payload_61_imag,
  input      [15:0]   io_data_in_payload_62_real,
  input      [15:0]   io_data_in_payload_62_imag,
  input      [15:0]   io_data_in_payload_63_real,
  input      [15:0]   io_data_in_payload_63_imag,
  input      [15:0]   io_data_in_payload_64_real,
  input      [15:0]   io_data_in_payload_64_imag,
  input      [15:0]   io_data_in_payload_65_real,
  input      [15:0]   io_data_in_payload_65_imag,
  input      [15:0]   io_data_in_payload_66_real,
  input      [15:0]   io_data_in_payload_66_imag,
  input      [15:0]   io_data_in_payload_67_real,
  input      [15:0]   io_data_in_payload_67_imag,
  input      [15:0]   io_data_in_payload_68_real,
  input      [15:0]   io_data_in_payload_68_imag,
  input      [15:0]   io_data_in_payload_69_real,
  input      [15:0]   io_data_in_payload_69_imag,
  input      [15:0]   io_data_in_payload_70_real,
  input      [15:0]   io_data_in_payload_70_imag,
  input      [15:0]   io_data_in_payload_71_real,
  input      [15:0]   io_data_in_payload_71_imag,
  input      [15:0]   io_data_in_payload_72_real,
  input      [15:0]   io_data_in_payload_72_imag,
  input      [15:0]   io_data_in_payload_73_real,
  input      [15:0]   io_data_in_payload_73_imag,
  input      [15:0]   io_data_in_payload_74_real,
  input      [15:0]   io_data_in_payload_74_imag,
  input      [15:0]   io_data_in_payload_75_real,
  input      [15:0]   io_data_in_payload_75_imag,
  input      [15:0]   io_data_in_payload_76_real,
  input      [15:0]   io_data_in_payload_76_imag,
  input      [15:0]   io_data_in_payload_77_real,
  input      [15:0]   io_data_in_payload_77_imag,
  input      [15:0]   io_data_in_payload_78_real,
  input      [15:0]   io_data_in_payload_78_imag,
  input      [15:0]   io_data_in_payload_79_real,
  input      [15:0]   io_data_in_payload_79_imag,
  input      [15:0]   io_data_in_payload_80_real,
  input      [15:0]   io_data_in_payload_80_imag,
  input      [15:0]   io_data_in_payload_81_real,
  input      [15:0]   io_data_in_payload_81_imag,
  input      [15:0]   io_data_in_payload_82_real,
  input      [15:0]   io_data_in_payload_82_imag,
  input      [15:0]   io_data_in_payload_83_real,
  input      [15:0]   io_data_in_payload_83_imag,
  input      [15:0]   io_data_in_payload_84_real,
  input      [15:0]   io_data_in_payload_84_imag,
  input      [15:0]   io_data_in_payload_85_real,
  input      [15:0]   io_data_in_payload_85_imag,
  input      [15:0]   io_data_in_payload_86_real,
  input      [15:0]   io_data_in_payload_86_imag,
  input      [15:0]   io_data_in_payload_87_real,
  input      [15:0]   io_data_in_payload_87_imag,
  input      [15:0]   io_data_in_payload_88_real,
  input      [15:0]   io_data_in_payload_88_imag,
  input      [15:0]   io_data_in_payload_89_real,
  input      [15:0]   io_data_in_payload_89_imag,
  input      [15:0]   io_data_in_payload_90_real,
  input      [15:0]   io_data_in_payload_90_imag,
  input      [15:0]   io_data_in_payload_91_real,
  input      [15:0]   io_data_in_payload_91_imag,
  input      [15:0]   io_data_in_payload_92_real,
  input      [15:0]   io_data_in_payload_92_imag,
  input      [15:0]   io_data_in_payload_93_real,
  input      [15:0]   io_data_in_payload_93_imag,
  input      [15:0]   io_data_in_payload_94_real,
  input      [15:0]   io_data_in_payload_94_imag,
  input      [15:0]   io_data_in_payload_95_real,
  input      [15:0]   io_data_in_payload_95_imag,
  input      [15:0]   io_data_in_payload_96_real,
  input      [15:0]   io_data_in_payload_96_imag,
  input      [15:0]   io_data_in_payload_97_real,
  input      [15:0]   io_data_in_payload_97_imag,
  input      [15:0]   io_data_in_payload_98_real,
  input      [15:0]   io_data_in_payload_98_imag,
  input      [15:0]   io_data_in_payload_99_real,
  input      [15:0]   io_data_in_payload_99_imag,
  input      [15:0]   io_data_in_payload_100_real,
  input      [15:0]   io_data_in_payload_100_imag,
  input      [15:0]   io_data_in_payload_101_real,
  input      [15:0]   io_data_in_payload_101_imag,
  input      [15:0]   io_data_in_payload_102_real,
  input      [15:0]   io_data_in_payload_102_imag,
  input      [15:0]   io_data_in_payload_103_real,
  input      [15:0]   io_data_in_payload_103_imag,
  input      [15:0]   io_data_in_payload_104_real,
  input      [15:0]   io_data_in_payload_104_imag,
  input      [15:0]   io_data_in_payload_105_real,
  input      [15:0]   io_data_in_payload_105_imag,
  input      [15:0]   io_data_in_payload_106_real,
  input      [15:0]   io_data_in_payload_106_imag,
  input      [15:0]   io_data_in_payload_107_real,
  input      [15:0]   io_data_in_payload_107_imag,
  input      [15:0]   io_data_in_payload_108_real,
  input      [15:0]   io_data_in_payload_108_imag,
  input      [15:0]   io_data_in_payload_109_real,
  input      [15:0]   io_data_in_payload_109_imag,
  input      [15:0]   io_data_in_payload_110_real,
  input      [15:0]   io_data_in_payload_110_imag,
  input      [15:0]   io_data_in_payload_111_real,
  input      [15:0]   io_data_in_payload_111_imag,
  input      [15:0]   io_data_in_payload_112_real,
  input      [15:0]   io_data_in_payload_112_imag,
  input      [15:0]   io_data_in_payload_113_real,
  input      [15:0]   io_data_in_payload_113_imag,
  input      [15:0]   io_data_in_payload_114_real,
  input      [15:0]   io_data_in_payload_114_imag,
  input      [15:0]   io_data_in_payload_115_real,
  input      [15:0]   io_data_in_payload_115_imag,
  input      [15:0]   io_data_in_payload_116_real,
  input      [15:0]   io_data_in_payload_116_imag,
  input      [15:0]   io_data_in_payload_117_real,
  input      [15:0]   io_data_in_payload_117_imag,
  input      [15:0]   io_data_in_payload_118_real,
  input      [15:0]   io_data_in_payload_118_imag,
  input      [15:0]   io_data_in_payload_119_real,
  input      [15:0]   io_data_in_payload_119_imag,
  input      [15:0]   io_data_in_payload_120_real,
  input      [15:0]   io_data_in_payload_120_imag,
  input      [15:0]   io_data_in_payload_121_real,
  input      [15:0]   io_data_in_payload_121_imag,
  input      [15:0]   io_data_in_payload_122_real,
  input      [15:0]   io_data_in_payload_122_imag,
  input      [15:0]   io_data_in_payload_123_real,
  input      [15:0]   io_data_in_payload_123_imag,
  input      [15:0]   io_data_in_payload_124_real,
  input      [15:0]   io_data_in_payload_124_imag,
  input      [15:0]   io_data_in_payload_125_real,
  input      [15:0]   io_data_in_payload_125_imag,
  input      [15:0]   io_data_in_payload_126_real,
  input      [15:0]   io_data_in_payload_126_imag,
  input      [15:0]   io_data_in_payload_127_real,
  input      [15:0]   io_data_in_payload_127_imag,
  output              io_data_out_valid,
  output     [15:0]   io_data_out_payload_0_real,
  output     [15:0]   io_data_out_payload_0_imag,
  output     [15:0]   io_data_out_payload_1_real,
  output     [15:0]   io_data_out_payload_1_imag,
  output     [15:0]   io_data_out_payload_2_real,
  output     [15:0]   io_data_out_payload_2_imag,
  output     [15:0]   io_data_out_payload_3_real,
  output     [15:0]   io_data_out_payload_3_imag,
  output     [15:0]   io_data_out_payload_4_real,
  output     [15:0]   io_data_out_payload_4_imag,
  output     [15:0]   io_data_out_payload_5_real,
  output     [15:0]   io_data_out_payload_5_imag,
  output     [15:0]   io_data_out_payload_6_real,
  output     [15:0]   io_data_out_payload_6_imag,
  output     [15:0]   io_data_out_payload_7_real,
  output     [15:0]   io_data_out_payload_7_imag,
  output     [15:0]   io_data_out_payload_8_real,
  output     [15:0]   io_data_out_payload_8_imag,
  output     [15:0]   io_data_out_payload_9_real,
  output     [15:0]   io_data_out_payload_9_imag,
  output     [15:0]   io_data_out_payload_10_real,
  output     [15:0]   io_data_out_payload_10_imag,
  output     [15:0]   io_data_out_payload_11_real,
  output     [15:0]   io_data_out_payload_11_imag,
  output     [15:0]   io_data_out_payload_12_real,
  output     [15:0]   io_data_out_payload_12_imag,
  output     [15:0]   io_data_out_payload_13_real,
  output     [15:0]   io_data_out_payload_13_imag,
  output     [15:0]   io_data_out_payload_14_real,
  output     [15:0]   io_data_out_payload_14_imag,
  output     [15:0]   io_data_out_payload_15_real,
  output     [15:0]   io_data_out_payload_15_imag,
  output     [15:0]   io_data_out_payload_16_real,
  output     [15:0]   io_data_out_payload_16_imag,
  output     [15:0]   io_data_out_payload_17_real,
  output     [15:0]   io_data_out_payload_17_imag,
  output     [15:0]   io_data_out_payload_18_real,
  output     [15:0]   io_data_out_payload_18_imag,
  output     [15:0]   io_data_out_payload_19_real,
  output     [15:0]   io_data_out_payload_19_imag,
  output     [15:0]   io_data_out_payload_20_real,
  output     [15:0]   io_data_out_payload_20_imag,
  output     [15:0]   io_data_out_payload_21_real,
  output     [15:0]   io_data_out_payload_21_imag,
  output     [15:0]   io_data_out_payload_22_real,
  output     [15:0]   io_data_out_payload_22_imag,
  output     [15:0]   io_data_out_payload_23_real,
  output     [15:0]   io_data_out_payload_23_imag,
  output     [15:0]   io_data_out_payload_24_real,
  output     [15:0]   io_data_out_payload_24_imag,
  output     [15:0]   io_data_out_payload_25_real,
  output     [15:0]   io_data_out_payload_25_imag,
  output     [15:0]   io_data_out_payload_26_real,
  output     [15:0]   io_data_out_payload_26_imag,
  output     [15:0]   io_data_out_payload_27_real,
  output     [15:0]   io_data_out_payload_27_imag,
  output     [15:0]   io_data_out_payload_28_real,
  output     [15:0]   io_data_out_payload_28_imag,
  output     [15:0]   io_data_out_payload_29_real,
  output     [15:0]   io_data_out_payload_29_imag,
  output     [15:0]   io_data_out_payload_30_real,
  output     [15:0]   io_data_out_payload_30_imag,
  output     [15:0]   io_data_out_payload_31_real,
  output     [15:0]   io_data_out_payload_31_imag,
  output     [15:0]   io_data_out_payload_32_real,
  output     [15:0]   io_data_out_payload_32_imag,
  output     [15:0]   io_data_out_payload_33_real,
  output     [15:0]   io_data_out_payload_33_imag,
  output     [15:0]   io_data_out_payload_34_real,
  output     [15:0]   io_data_out_payload_34_imag,
  output     [15:0]   io_data_out_payload_35_real,
  output     [15:0]   io_data_out_payload_35_imag,
  output     [15:0]   io_data_out_payload_36_real,
  output     [15:0]   io_data_out_payload_36_imag,
  output     [15:0]   io_data_out_payload_37_real,
  output     [15:0]   io_data_out_payload_37_imag,
  output     [15:0]   io_data_out_payload_38_real,
  output     [15:0]   io_data_out_payload_38_imag,
  output     [15:0]   io_data_out_payload_39_real,
  output     [15:0]   io_data_out_payload_39_imag,
  output     [15:0]   io_data_out_payload_40_real,
  output     [15:0]   io_data_out_payload_40_imag,
  output     [15:0]   io_data_out_payload_41_real,
  output     [15:0]   io_data_out_payload_41_imag,
  output     [15:0]   io_data_out_payload_42_real,
  output     [15:0]   io_data_out_payload_42_imag,
  output     [15:0]   io_data_out_payload_43_real,
  output     [15:0]   io_data_out_payload_43_imag,
  output     [15:0]   io_data_out_payload_44_real,
  output     [15:0]   io_data_out_payload_44_imag,
  output     [15:0]   io_data_out_payload_45_real,
  output     [15:0]   io_data_out_payload_45_imag,
  output     [15:0]   io_data_out_payload_46_real,
  output     [15:0]   io_data_out_payload_46_imag,
  output     [15:0]   io_data_out_payload_47_real,
  output     [15:0]   io_data_out_payload_47_imag,
  output     [15:0]   io_data_out_payload_48_real,
  output     [15:0]   io_data_out_payload_48_imag,
  output     [15:0]   io_data_out_payload_49_real,
  output     [15:0]   io_data_out_payload_49_imag,
  output     [15:0]   io_data_out_payload_50_real,
  output     [15:0]   io_data_out_payload_50_imag,
  output     [15:0]   io_data_out_payload_51_real,
  output     [15:0]   io_data_out_payload_51_imag,
  output     [15:0]   io_data_out_payload_52_real,
  output     [15:0]   io_data_out_payload_52_imag,
  output     [15:0]   io_data_out_payload_53_real,
  output     [15:0]   io_data_out_payload_53_imag,
  output     [15:0]   io_data_out_payload_54_real,
  output     [15:0]   io_data_out_payload_54_imag,
  output     [15:0]   io_data_out_payload_55_real,
  output     [15:0]   io_data_out_payload_55_imag,
  output     [15:0]   io_data_out_payload_56_real,
  output     [15:0]   io_data_out_payload_56_imag,
  output     [15:0]   io_data_out_payload_57_real,
  output     [15:0]   io_data_out_payload_57_imag,
  output     [15:0]   io_data_out_payload_58_real,
  output     [15:0]   io_data_out_payload_58_imag,
  output     [15:0]   io_data_out_payload_59_real,
  output     [15:0]   io_data_out_payload_59_imag,
  output     [15:0]   io_data_out_payload_60_real,
  output     [15:0]   io_data_out_payload_60_imag,
  output     [15:0]   io_data_out_payload_61_real,
  output     [15:0]   io_data_out_payload_61_imag,
  output     [15:0]   io_data_out_payload_62_real,
  output     [15:0]   io_data_out_payload_62_imag,
  output     [15:0]   io_data_out_payload_63_real,
  output     [15:0]   io_data_out_payload_63_imag,
  output     [15:0]   io_data_out_payload_64_real,
  output     [15:0]   io_data_out_payload_64_imag,
  output     [15:0]   io_data_out_payload_65_real,
  output     [15:0]   io_data_out_payload_65_imag,
  output     [15:0]   io_data_out_payload_66_real,
  output     [15:0]   io_data_out_payload_66_imag,
  output     [15:0]   io_data_out_payload_67_real,
  output     [15:0]   io_data_out_payload_67_imag,
  output     [15:0]   io_data_out_payload_68_real,
  output     [15:0]   io_data_out_payload_68_imag,
  output     [15:0]   io_data_out_payload_69_real,
  output     [15:0]   io_data_out_payload_69_imag,
  output     [15:0]   io_data_out_payload_70_real,
  output     [15:0]   io_data_out_payload_70_imag,
  output     [15:0]   io_data_out_payload_71_real,
  output     [15:0]   io_data_out_payload_71_imag,
  output     [15:0]   io_data_out_payload_72_real,
  output     [15:0]   io_data_out_payload_72_imag,
  output     [15:0]   io_data_out_payload_73_real,
  output     [15:0]   io_data_out_payload_73_imag,
  output     [15:0]   io_data_out_payload_74_real,
  output     [15:0]   io_data_out_payload_74_imag,
  output     [15:0]   io_data_out_payload_75_real,
  output     [15:0]   io_data_out_payload_75_imag,
  output     [15:0]   io_data_out_payload_76_real,
  output     [15:0]   io_data_out_payload_76_imag,
  output     [15:0]   io_data_out_payload_77_real,
  output     [15:0]   io_data_out_payload_77_imag,
  output     [15:0]   io_data_out_payload_78_real,
  output     [15:0]   io_data_out_payload_78_imag,
  output     [15:0]   io_data_out_payload_79_real,
  output     [15:0]   io_data_out_payload_79_imag,
  output     [15:0]   io_data_out_payload_80_real,
  output     [15:0]   io_data_out_payload_80_imag,
  output     [15:0]   io_data_out_payload_81_real,
  output     [15:0]   io_data_out_payload_81_imag,
  output     [15:0]   io_data_out_payload_82_real,
  output     [15:0]   io_data_out_payload_82_imag,
  output     [15:0]   io_data_out_payload_83_real,
  output     [15:0]   io_data_out_payload_83_imag,
  output     [15:0]   io_data_out_payload_84_real,
  output     [15:0]   io_data_out_payload_84_imag,
  output     [15:0]   io_data_out_payload_85_real,
  output     [15:0]   io_data_out_payload_85_imag,
  output     [15:0]   io_data_out_payload_86_real,
  output     [15:0]   io_data_out_payload_86_imag,
  output     [15:0]   io_data_out_payload_87_real,
  output     [15:0]   io_data_out_payload_87_imag,
  output     [15:0]   io_data_out_payload_88_real,
  output     [15:0]   io_data_out_payload_88_imag,
  output     [15:0]   io_data_out_payload_89_real,
  output     [15:0]   io_data_out_payload_89_imag,
  output     [15:0]   io_data_out_payload_90_real,
  output     [15:0]   io_data_out_payload_90_imag,
  output     [15:0]   io_data_out_payload_91_real,
  output     [15:0]   io_data_out_payload_91_imag,
  output     [15:0]   io_data_out_payload_92_real,
  output     [15:0]   io_data_out_payload_92_imag,
  output     [15:0]   io_data_out_payload_93_real,
  output     [15:0]   io_data_out_payload_93_imag,
  output     [15:0]   io_data_out_payload_94_real,
  output     [15:0]   io_data_out_payload_94_imag,
  output     [15:0]   io_data_out_payload_95_real,
  output     [15:0]   io_data_out_payload_95_imag,
  output     [15:0]   io_data_out_payload_96_real,
  output     [15:0]   io_data_out_payload_96_imag,
  output     [15:0]   io_data_out_payload_97_real,
  output     [15:0]   io_data_out_payload_97_imag,
  output     [15:0]   io_data_out_payload_98_real,
  output     [15:0]   io_data_out_payload_98_imag,
  output     [15:0]   io_data_out_payload_99_real,
  output     [15:0]   io_data_out_payload_99_imag,
  output     [15:0]   io_data_out_payload_100_real,
  output     [15:0]   io_data_out_payload_100_imag,
  output     [15:0]   io_data_out_payload_101_real,
  output     [15:0]   io_data_out_payload_101_imag,
  output     [15:0]   io_data_out_payload_102_real,
  output     [15:0]   io_data_out_payload_102_imag,
  output     [15:0]   io_data_out_payload_103_real,
  output     [15:0]   io_data_out_payload_103_imag,
  output     [15:0]   io_data_out_payload_104_real,
  output     [15:0]   io_data_out_payload_104_imag,
  output     [15:0]   io_data_out_payload_105_real,
  output     [15:0]   io_data_out_payload_105_imag,
  output     [15:0]   io_data_out_payload_106_real,
  output     [15:0]   io_data_out_payload_106_imag,
  output     [15:0]   io_data_out_payload_107_real,
  output     [15:0]   io_data_out_payload_107_imag,
  output     [15:0]   io_data_out_payload_108_real,
  output     [15:0]   io_data_out_payload_108_imag,
  output     [15:0]   io_data_out_payload_109_real,
  output     [15:0]   io_data_out_payload_109_imag,
  output     [15:0]   io_data_out_payload_110_real,
  output     [15:0]   io_data_out_payload_110_imag,
  output     [15:0]   io_data_out_payload_111_real,
  output     [15:0]   io_data_out_payload_111_imag,
  output     [15:0]   io_data_out_payload_112_real,
  output     [15:0]   io_data_out_payload_112_imag,
  output     [15:0]   io_data_out_payload_113_real,
  output     [15:0]   io_data_out_payload_113_imag,
  output     [15:0]   io_data_out_payload_114_real,
  output     [15:0]   io_data_out_payload_114_imag,
  output     [15:0]   io_data_out_payload_115_real,
  output     [15:0]   io_data_out_payload_115_imag,
  output     [15:0]   io_data_out_payload_116_real,
  output     [15:0]   io_data_out_payload_116_imag,
  output     [15:0]   io_data_out_payload_117_real,
  output     [15:0]   io_data_out_payload_117_imag,
  output     [15:0]   io_data_out_payload_118_real,
  output     [15:0]   io_data_out_payload_118_imag,
  output     [15:0]   io_data_out_payload_119_real,
  output     [15:0]   io_data_out_payload_119_imag,
  output     [15:0]   io_data_out_payload_120_real,
  output     [15:0]   io_data_out_payload_120_imag,
  output     [15:0]   io_data_out_payload_121_real,
  output     [15:0]   io_data_out_payload_121_imag,
  output     [15:0]   io_data_out_payload_122_real,
  output     [15:0]   io_data_out_payload_122_imag,
  output     [15:0]   io_data_out_payload_123_real,
  output     [15:0]   io_data_out_payload_123_imag,
  output     [15:0]   io_data_out_payload_124_real,
  output     [15:0]   io_data_out_payload_124_imag,
  output     [15:0]   io_data_out_payload_125_real,
  output     [15:0]   io_data_out_payload_125_imag,
  output     [15:0]   io_data_out_payload_126_real,
  output     [15:0]   io_data_out_payload_126_imag,
  output     [15:0]   io_data_out_payload_127_real,
  output     [15:0]   io_data_out_payload_127_imag,
  input               clk,
  input               reset
);
  wire       [31:0]   _zz_4039;
  wire       [31:0]   _zz_4040;
  wire       [31:0]   _zz_4041;
  wire       [31:0]   _zz_4042;
  wire       [31:0]   _zz_4043;
  wire       [31:0]   _zz_4044;
  wire       [31:0]   _zz_4045;
  wire       [31:0]   _zz_4046;
  wire       [31:0]   _zz_4047;
  wire       [31:0]   _zz_4048;
  wire       [31:0]   _zz_4049;
  wire       [31:0]   _zz_4050;
  wire       [31:0]   _zz_4051;
  wire       [31:0]   _zz_4052;
  wire       [31:0]   _zz_4053;
  wire       [31:0]   _zz_4054;
  wire       [31:0]   _zz_4055;
  wire       [31:0]   _zz_4056;
  wire       [31:0]   _zz_4057;
  wire       [31:0]   _zz_4058;
  wire       [31:0]   _zz_4059;
  wire       [31:0]   _zz_4060;
  wire       [31:0]   _zz_4061;
  wire       [31:0]   _zz_4062;
  wire       [31:0]   _zz_4063;
  wire       [31:0]   _zz_4064;
  wire       [31:0]   _zz_4065;
  wire       [31:0]   _zz_4066;
  wire       [31:0]   _zz_4067;
  wire       [31:0]   _zz_4068;
  wire       [31:0]   _zz_4069;
  wire       [31:0]   _zz_4070;
  wire       [31:0]   _zz_4071;
  wire       [31:0]   _zz_4072;
  wire       [31:0]   _zz_4073;
  wire       [31:0]   _zz_4074;
  wire       [31:0]   _zz_4075;
  wire       [31:0]   _zz_4076;
  wire       [31:0]   _zz_4077;
  wire       [31:0]   _zz_4078;
  wire       [31:0]   _zz_4079;
  wire       [31:0]   _zz_4080;
  wire       [31:0]   _zz_4081;
  wire       [31:0]   _zz_4082;
  wire       [31:0]   _zz_4083;
  wire       [31:0]   _zz_4084;
  wire       [31:0]   _zz_4085;
  wire       [31:0]   _zz_4086;
  wire       [31:0]   _zz_4087;
  wire       [31:0]   _zz_4088;
  wire       [31:0]   _zz_4089;
  wire       [31:0]   _zz_4090;
  wire       [31:0]   _zz_4091;
  wire       [31:0]   _zz_4092;
  wire       [31:0]   _zz_4093;
  wire       [31:0]   _zz_4094;
  wire       [31:0]   _zz_4095;
  wire       [31:0]   _zz_4096;
  wire       [31:0]   _zz_4097;
  wire       [31:0]   _zz_4098;
  wire       [31:0]   _zz_4099;
  wire       [31:0]   _zz_4100;
  wire       [31:0]   _zz_4101;
  wire       [31:0]   _zz_4102;
  wire       [31:0]   _zz_4103;
  wire       [31:0]   _zz_4104;
  wire       [31:0]   _zz_4105;
  wire       [31:0]   _zz_4106;
  wire       [31:0]   _zz_4107;
  wire       [31:0]   _zz_4108;
  wire       [31:0]   _zz_4109;
  wire       [31:0]   _zz_4110;
  wire       [31:0]   _zz_4111;
  wire       [31:0]   _zz_4112;
  wire       [31:0]   _zz_4113;
  wire       [31:0]   _zz_4114;
  wire       [31:0]   _zz_4115;
  wire       [31:0]   _zz_4116;
  wire       [31:0]   _zz_4117;
  wire       [31:0]   _zz_4118;
  wire       [31:0]   _zz_4119;
  wire       [31:0]   _zz_4120;
  wire       [31:0]   _zz_4121;
  wire       [31:0]   _zz_4122;
  wire       [31:0]   _zz_4123;
  wire       [31:0]   _zz_4124;
  wire       [31:0]   _zz_4125;
  wire       [31:0]   _zz_4126;
  wire       [31:0]   _zz_4127;
  wire       [31:0]   _zz_4128;
  wire       [31:0]   _zz_4129;
  wire       [31:0]   _zz_4130;
  wire       [31:0]   _zz_4131;
  wire       [31:0]   _zz_4132;
  wire       [31:0]   _zz_4133;
  wire       [31:0]   _zz_4134;
  wire       [31:0]   _zz_4135;
  wire       [31:0]   _zz_4136;
  wire       [31:0]   _zz_4137;
  wire       [31:0]   _zz_4138;
  wire       [31:0]   _zz_4139;
  wire       [31:0]   _zz_4140;
  wire       [31:0]   _zz_4141;
  wire       [31:0]   _zz_4142;
  wire       [31:0]   _zz_4143;
  wire       [31:0]   _zz_4144;
  wire       [31:0]   _zz_4145;
  wire       [31:0]   _zz_4146;
  wire       [31:0]   _zz_4147;
  wire       [31:0]   _zz_4148;
  wire       [31:0]   _zz_4149;
  wire       [31:0]   _zz_4150;
  wire       [31:0]   _zz_4151;
  wire       [31:0]   _zz_4152;
  wire       [31:0]   _zz_4153;
  wire       [31:0]   _zz_4154;
  wire       [31:0]   _zz_4155;
  wire       [31:0]   _zz_4156;
  wire       [31:0]   _zz_4157;
  wire       [31:0]   _zz_4158;
  wire       [31:0]   _zz_4159;
  wire       [31:0]   _zz_4160;
  wire       [31:0]   _zz_4161;
  wire       [31:0]   _zz_4162;
  wire       [31:0]   _zz_4163;
  wire       [31:0]   _zz_4164;
  wire       [31:0]   _zz_4165;
  wire       [31:0]   _zz_4166;
  wire       [31:0]   _zz_4167;
  wire       [31:0]   _zz_4168;
  wire       [31:0]   _zz_4169;
  wire       [31:0]   _zz_4170;
  wire       [31:0]   _zz_4171;
  wire       [31:0]   _zz_4172;
  wire       [31:0]   _zz_4173;
  wire       [31:0]   _zz_4174;
  wire       [31:0]   _zz_4175;
  wire       [31:0]   _zz_4176;
  wire       [31:0]   _zz_4177;
  wire       [31:0]   _zz_4178;
  wire       [31:0]   _zz_4179;
  wire       [31:0]   _zz_4180;
  wire       [31:0]   _zz_4181;
  wire       [31:0]   _zz_4182;
  wire       [31:0]   _zz_4183;
  wire       [31:0]   _zz_4184;
  wire       [31:0]   _zz_4185;
  wire       [31:0]   _zz_4186;
  wire       [31:0]   _zz_4187;
  wire       [31:0]   _zz_4188;
  wire       [31:0]   _zz_4189;
  wire       [31:0]   _zz_4190;
  wire       [31:0]   _zz_4191;
  wire       [31:0]   _zz_4192;
  wire       [31:0]   _zz_4193;
  wire       [31:0]   _zz_4194;
  wire       [31:0]   _zz_4195;
  wire       [31:0]   _zz_4196;
  wire       [31:0]   _zz_4197;
  wire       [31:0]   _zz_4198;
  wire       [31:0]   _zz_4199;
  wire       [31:0]   _zz_4200;
  wire       [31:0]   _zz_4201;
  wire       [31:0]   _zz_4202;
  wire       [31:0]   _zz_4203;
  wire       [31:0]   _zz_4204;
  wire       [31:0]   _zz_4205;
  wire       [31:0]   _zz_4206;
  wire       [31:0]   _zz_4207;
  wire       [31:0]   _zz_4208;
  wire       [31:0]   _zz_4209;
  wire       [31:0]   _zz_4210;
  wire       [31:0]   _zz_4211;
  wire       [31:0]   _zz_4212;
  wire       [31:0]   _zz_4213;
  wire       [31:0]   _zz_4214;
  wire       [31:0]   _zz_4215;
  wire       [31:0]   _zz_4216;
  wire       [31:0]   _zz_4217;
  wire       [31:0]   _zz_4218;
  wire       [31:0]   _zz_4219;
  wire       [31:0]   _zz_4220;
  wire       [31:0]   _zz_4221;
  wire       [31:0]   _zz_4222;
  wire       [31:0]   _zz_4223;
  wire       [31:0]   _zz_4224;
  wire       [31:0]   _zz_4225;
  wire       [31:0]   _zz_4226;
  wire       [31:0]   _zz_4227;
  wire       [31:0]   _zz_4228;
  wire       [31:0]   _zz_4229;
  wire       [31:0]   _zz_4230;
  wire       [31:0]   _zz_4231;
  wire       [31:0]   _zz_4232;
  wire       [31:0]   _zz_4233;
  wire       [31:0]   _zz_4234;
  wire       [31:0]   _zz_4235;
  wire       [31:0]   _zz_4236;
  wire       [31:0]   _zz_4237;
  wire       [31:0]   _zz_4238;
  wire       [31:0]   _zz_4239;
  wire       [31:0]   _zz_4240;
  wire       [31:0]   _zz_4241;
  wire       [31:0]   _zz_4242;
  wire       [31:0]   _zz_4243;
  wire       [31:0]   _zz_4244;
  wire       [31:0]   _zz_4245;
  wire       [31:0]   _zz_4246;
  wire       [31:0]   _zz_4247;
  wire       [31:0]   _zz_4248;
  wire       [31:0]   _zz_4249;
  wire       [31:0]   _zz_4250;
  wire       [31:0]   _zz_4251;
  wire       [31:0]   _zz_4252;
  wire       [31:0]   _zz_4253;
  wire       [31:0]   _zz_4254;
  wire       [31:0]   _zz_4255;
  wire       [31:0]   _zz_4256;
  wire       [31:0]   _zz_4257;
  wire       [31:0]   _zz_4258;
  wire       [31:0]   _zz_4259;
  wire       [31:0]   _zz_4260;
  wire       [31:0]   _zz_4261;
  wire       [31:0]   _zz_4262;
  wire       [31:0]   _zz_4263;
  wire       [31:0]   _zz_4264;
  wire       [31:0]   _zz_4265;
  wire       [31:0]   _zz_4266;
  wire       [31:0]   _zz_4267;
  wire       [31:0]   _zz_4268;
  wire       [31:0]   _zz_4269;
  wire       [31:0]   _zz_4270;
  wire       [31:0]   _zz_4271;
  wire       [31:0]   _zz_4272;
  wire       [31:0]   _zz_4273;
  wire       [31:0]   _zz_4274;
  wire       [31:0]   _zz_4275;
  wire       [31:0]   _zz_4276;
  wire       [31:0]   _zz_4277;
  wire       [31:0]   _zz_4278;
  wire       [31:0]   _zz_4279;
  wire       [31:0]   _zz_4280;
  wire       [31:0]   _zz_4281;
  wire       [31:0]   _zz_4282;
  wire       [31:0]   _zz_4283;
  wire       [31:0]   _zz_4284;
  wire       [31:0]   _zz_4285;
  wire       [31:0]   _zz_4286;
  wire       [31:0]   _zz_4287;
  wire       [31:0]   _zz_4288;
  wire       [31:0]   _zz_4289;
  wire       [31:0]   _zz_4290;
  wire       [31:0]   _zz_4291;
  wire       [31:0]   _zz_4292;
  wire       [31:0]   _zz_4293;
  wire       [31:0]   _zz_4294;
  wire       [31:0]   _zz_4295;
  wire       [31:0]   _zz_4296;
  wire       [31:0]   _zz_4297;
  wire       [31:0]   _zz_4298;
  wire       [31:0]   _zz_4299;
  wire       [31:0]   _zz_4300;
  wire       [31:0]   _zz_4301;
  wire       [31:0]   _zz_4302;
  wire       [31:0]   _zz_4303;
  wire       [31:0]   _zz_4304;
  wire       [31:0]   _zz_4305;
  wire       [31:0]   _zz_4306;
  wire       [31:0]   _zz_4307;
  wire       [31:0]   _zz_4308;
  wire       [31:0]   _zz_4309;
  wire       [31:0]   _zz_4310;
  wire       [31:0]   _zz_4311;
  wire       [31:0]   _zz_4312;
  wire       [31:0]   _zz_4313;
  wire       [31:0]   _zz_4314;
  wire       [31:0]   _zz_4315;
  wire       [31:0]   _zz_4316;
  wire       [31:0]   _zz_4317;
  wire       [31:0]   _zz_4318;
  wire       [31:0]   _zz_4319;
  wire       [31:0]   _zz_4320;
  wire       [31:0]   _zz_4321;
  wire       [31:0]   _zz_4322;
  wire       [31:0]   _zz_4323;
  wire       [31:0]   _zz_4324;
  wire       [31:0]   _zz_4325;
  wire       [31:0]   _zz_4326;
  wire       [31:0]   _zz_4327;
  wire       [31:0]   _zz_4328;
  wire       [31:0]   _zz_4329;
  wire       [31:0]   _zz_4330;
  wire       [31:0]   _zz_4331;
  wire       [31:0]   _zz_4332;
  wire       [31:0]   _zz_4333;
  wire       [31:0]   _zz_4334;
  wire       [31:0]   _zz_4335;
  wire       [31:0]   _zz_4336;
  wire       [31:0]   _zz_4337;
  wire       [31:0]   _zz_4338;
  wire       [31:0]   _zz_4339;
  wire       [31:0]   _zz_4340;
  wire       [31:0]   _zz_4341;
  wire       [31:0]   _zz_4342;
  wire       [31:0]   _zz_4343;
  wire       [31:0]   _zz_4344;
  wire       [31:0]   _zz_4345;
  wire       [31:0]   _zz_4346;
  wire       [31:0]   _zz_4347;
  wire       [31:0]   _zz_4348;
  wire       [31:0]   _zz_4349;
  wire       [31:0]   _zz_4350;
  wire       [31:0]   _zz_4351;
  wire       [31:0]   _zz_4352;
  wire       [31:0]   _zz_4353;
  wire       [31:0]   _zz_4354;
  wire       [31:0]   _zz_4355;
  wire       [31:0]   _zz_4356;
  wire       [31:0]   _zz_4357;
  wire       [31:0]   _zz_4358;
  wire       [31:0]   _zz_4359;
  wire       [31:0]   _zz_4360;
  wire       [31:0]   _zz_4361;
  wire       [31:0]   _zz_4362;
  wire       [31:0]   _zz_4363;
  wire       [31:0]   _zz_4364;
  wire       [31:0]   _zz_4365;
  wire       [31:0]   _zz_4366;
  wire       [31:0]   _zz_4367;
  wire       [31:0]   _zz_4368;
  wire       [31:0]   _zz_4369;
  wire       [31:0]   _zz_4370;
  wire       [31:0]   _zz_4371;
  wire       [31:0]   _zz_4372;
  wire       [31:0]   _zz_4373;
  wire       [31:0]   _zz_4374;
  wire       [31:0]   _zz_4375;
  wire       [31:0]   _zz_4376;
  wire       [31:0]   _zz_4377;
  wire       [31:0]   _zz_4378;
  wire       [31:0]   _zz_4379;
  wire       [31:0]   _zz_4380;
  wire       [31:0]   _zz_4381;
  wire       [31:0]   _zz_4382;
  wire       [31:0]   _zz_4383;
  wire       [31:0]   _zz_4384;
  wire       [31:0]   _zz_4385;
  wire       [31:0]   _zz_4386;
  wire       [31:0]   _zz_4387;
  wire       [31:0]   _zz_4388;
  wire       [31:0]   _zz_4389;
  wire       [31:0]   _zz_4390;
  wire       [31:0]   _zz_4391;
  wire       [31:0]   _zz_4392;
  wire       [31:0]   _zz_4393;
  wire       [31:0]   _zz_4394;
  wire       [31:0]   _zz_4395;
  wire       [31:0]   _zz_4396;
  wire       [31:0]   _zz_4397;
  wire       [31:0]   _zz_4398;
  wire       [31:0]   _zz_4399;
  wire       [31:0]   _zz_4400;
  wire       [31:0]   _zz_4401;
  wire       [31:0]   _zz_4402;
  wire       [31:0]   _zz_4403;
  wire       [31:0]   _zz_4404;
  wire       [31:0]   _zz_4405;
  wire       [31:0]   _zz_4406;
  wire       [31:0]   _zz_4407;
  wire       [31:0]   _zz_4408;
  wire       [31:0]   _zz_4409;
  wire       [31:0]   _zz_4410;
  wire       [31:0]   _zz_4411;
  wire       [31:0]   _zz_4412;
  wire       [31:0]   _zz_4413;
  wire       [31:0]   _zz_4414;
  wire       [31:0]   _zz_4415;
  wire       [31:0]   _zz_4416;
  wire       [31:0]   _zz_4417;
  wire       [31:0]   _zz_4418;
  wire       [31:0]   _zz_4419;
  wire       [31:0]   _zz_4420;
  wire       [31:0]   _zz_4421;
  wire       [31:0]   _zz_4422;
  wire       [31:0]   _zz_4423;
  wire       [31:0]   _zz_4424;
  wire       [31:0]   _zz_4425;
  wire       [31:0]   _zz_4426;
  wire       [31:0]   _zz_4427;
  wire       [31:0]   _zz_4428;
  wire       [31:0]   _zz_4429;
  wire       [31:0]   _zz_4430;
  wire       [31:0]   _zz_4431;
  wire       [31:0]   _zz_4432;
  wire       [31:0]   _zz_4433;
  wire       [31:0]   _zz_4434;
  wire       [31:0]   _zz_4435;
  wire       [31:0]   _zz_4436;
  wire       [31:0]   _zz_4437;
  wire       [31:0]   _zz_4438;
  wire       [31:0]   _zz_4439;
  wire       [31:0]   _zz_4440;
  wire       [31:0]   _zz_4441;
  wire       [31:0]   _zz_4442;
  wire       [31:0]   _zz_4443;
  wire       [31:0]   _zz_4444;
  wire       [31:0]   _zz_4445;
  wire       [31:0]   _zz_4446;
  wire       [31:0]   _zz_4447;
  wire       [31:0]   _zz_4448;
  wire       [31:0]   _zz_4449;
  wire       [31:0]   _zz_4450;
  wire       [31:0]   _zz_4451;
  wire       [31:0]   _zz_4452;
  wire       [31:0]   _zz_4453;
  wire       [31:0]   _zz_4454;
  wire       [31:0]   _zz_4455;
  wire       [31:0]   _zz_4456;
  wire       [31:0]   _zz_4457;
  wire       [31:0]   _zz_4458;
  wire       [31:0]   _zz_4459;
  wire       [31:0]   _zz_4460;
  wire       [31:0]   _zz_4461;
  wire       [31:0]   _zz_4462;
  wire       [31:0]   _zz_4463;
  wire       [31:0]   _zz_4464;
  wire       [31:0]   _zz_4465;
  wire       [31:0]   _zz_4466;
  wire       [31:0]   _zz_4467;
  wire       [31:0]   _zz_4468;
  wire       [31:0]   _zz_4469;
  wire       [31:0]   _zz_4470;
  wire       [31:0]   _zz_4471;
  wire       [31:0]   _zz_4472;
  wire       [31:0]   _zz_4473;
  wire       [31:0]   _zz_4474;
  wire       [31:0]   _zz_4475;
  wire       [31:0]   _zz_4476;
  wire       [31:0]   _zz_4477;
  wire       [31:0]   _zz_4478;
  wire       [31:0]   _zz_4479;
  wire       [31:0]   _zz_4480;
  wire       [31:0]   _zz_4481;
  wire       [31:0]   _zz_4482;
  wire       [31:0]   _zz_4483;
  wire       [31:0]   _zz_4484;
  wire       [31:0]   _zz_4485;
  wire       [31:0]   _zz_4486;
  wire       [31:0]   _zz_4487;
  wire       [31:0]   _zz_4488;
  wire       [31:0]   _zz_4489;
  wire       [31:0]   _zz_4490;
  wire       [31:0]   _zz_4491;
  wire       [31:0]   _zz_4492;
  wire       [31:0]   _zz_4493;
  wire       [31:0]   _zz_4494;
  wire       [31:0]   _zz_4495;
  wire       [31:0]   _zz_4496;
  wire       [31:0]   _zz_4497;
  wire       [31:0]   _zz_4498;
  wire       [31:0]   _zz_4499;
  wire       [31:0]   _zz_4500;
  wire       [31:0]   _zz_4501;
  wire       [31:0]   _zz_4502;
  wire       [31:0]   _zz_4503;
  wire       [31:0]   _zz_4504;
  wire       [31:0]   _zz_4505;
  wire       [31:0]   _zz_4506;
  wire       [31:0]   _zz_4507;
  wire       [31:0]   _zz_4508;
  wire       [31:0]   _zz_4509;
  wire       [31:0]   _zz_4510;
  wire       [31:0]   _zz_4511;
  wire       [31:0]   _zz_4512;
  wire       [31:0]   _zz_4513;
  wire       [31:0]   _zz_4514;
  wire       [31:0]   _zz_4515;
  wire       [31:0]   _zz_4516;
  wire       [31:0]   _zz_4517;
  wire       [31:0]   _zz_4518;
  wire       [31:0]   _zz_4519;
  wire       [31:0]   _zz_4520;
  wire       [31:0]   _zz_4521;
  wire       [31:0]   _zz_4522;
  wire       [31:0]   _zz_4523;
  wire       [31:0]   _zz_4524;
  wire       [31:0]   _zz_4525;
  wire       [31:0]   _zz_4526;
  wire       [31:0]   _zz_4527;
  wire       [31:0]   _zz_4528;
  wire       [31:0]   _zz_4529;
  wire       [31:0]   _zz_4530;
  wire       [31:0]   _zz_4531;
  wire       [31:0]   _zz_4532;
  wire       [31:0]   _zz_4533;
  wire       [31:0]   _zz_4534;
  wire       [31:0]   _zz_4535;
  wire       [31:0]   _zz_4536;
  wire       [31:0]   _zz_4537;
  wire       [31:0]   _zz_4538;
  wire       [31:0]   _zz_4539;
  wire       [31:0]   _zz_4540;
  wire       [31:0]   _zz_4541;
  wire       [31:0]   _zz_4542;
  wire       [31:0]   _zz_4543;
  wire       [31:0]   _zz_4544;
  wire       [31:0]   _zz_4545;
  wire       [31:0]   _zz_4546;
  wire       [31:0]   _zz_4547;
  wire       [31:0]   _zz_4548;
  wire       [31:0]   _zz_4549;
  wire       [31:0]   _zz_4550;
  wire       [31:0]   _zz_4551;
  wire       [31:0]   _zz_4552;
  wire       [31:0]   _zz_4553;
  wire       [31:0]   _zz_4554;
  wire       [31:0]   _zz_4555;
  wire       [31:0]   _zz_4556;
  wire       [31:0]   _zz_4557;
  wire       [31:0]   _zz_4558;
  wire       [31:0]   _zz_4559;
  wire       [31:0]   _zz_4560;
  wire       [31:0]   _zz_4561;
  wire       [31:0]   _zz_4562;
  wire       [31:0]   _zz_4563;
  wire       [31:0]   _zz_4564;
  wire       [31:0]   _zz_4565;
  wire       [31:0]   _zz_4566;
  wire       [31:0]   _zz_4567;
  wire       [31:0]   _zz_4568;
  wire       [31:0]   _zz_4569;
  wire       [31:0]   _zz_4570;
  wire       [31:0]   _zz_4571;
  wire       [31:0]   _zz_4572;
  wire       [31:0]   _zz_4573;
  wire       [31:0]   _zz_4574;
  wire       [31:0]   _zz_4575;
  wire       [31:0]   _zz_4576;
  wire       [31:0]   _zz_4577;
  wire       [31:0]   _zz_4578;
  wire       [31:0]   _zz_4579;
  wire       [31:0]   _zz_4580;
  wire       [31:0]   _zz_4581;
  wire       [31:0]   _zz_4582;
  wire       [31:0]   _zz_4583;
  wire       [31:0]   _zz_4584;
  wire       [31:0]   _zz_4585;
  wire       [31:0]   _zz_4586;
  wire       [31:0]   _zz_4587;
  wire       [31:0]   _zz_4588;
  wire       [31:0]   _zz_4589;
  wire       [31:0]   _zz_4590;
  wire       [31:0]   _zz_4591;
  wire       [31:0]   _zz_4592;
  wire       [31:0]   _zz_4593;
  wire       [31:0]   _zz_4594;
  wire       [31:0]   _zz_4595;
  wire       [31:0]   _zz_4596;
  wire       [31:0]   _zz_4597;
  wire       [31:0]   _zz_4598;
  wire       [31:0]   _zz_4599;
  wire       [31:0]   _zz_4600;
  wire       [31:0]   _zz_4601;
  wire       [31:0]   _zz_4602;
  wire       [31:0]   _zz_4603;
  wire       [31:0]   _zz_4604;
  wire       [31:0]   _zz_4605;
  wire       [31:0]   _zz_4606;
  wire       [31:0]   _zz_4607;
  wire       [31:0]   _zz_4608;
  wire       [31:0]   _zz_4609;
  wire       [31:0]   _zz_4610;
  wire       [31:0]   _zz_4611;
  wire       [31:0]   _zz_4612;
  wire       [31:0]   _zz_4613;
  wire       [31:0]   _zz_4614;
  wire       [31:0]   _zz_4615;
  wire       [31:0]   _zz_4616;
  wire       [31:0]   _zz_4617;
  wire       [31:0]   _zz_4618;
  wire       [31:0]   _zz_4619;
  wire       [31:0]   _zz_4620;
  wire       [31:0]   _zz_4621;
  wire       [31:0]   _zz_4622;
  wire       [31:0]   _zz_4623;
  wire       [31:0]   _zz_4624;
  wire       [31:0]   _zz_4625;
  wire       [31:0]   _zz_4626;
  wire       [31:0]   _zz_4627;
  wire       [31:0]   _zz_4628;
  wire       [31:0]   _zz_4629;
  wire       [31:0]   _zz_4630;
  wire       [31:0]   _zz_4631;
  wire       [31:0]   _zz_4632;
  wire       [31:0]   _zz_4633;
  wire       [31:0]   _zz_4634;
  wire       [31:0]   _zz_4635;
  wire       [31:0]   _zz_4636;
  wire       [31:0]   _zz_4637;
  wire       [31:0]   _zz_4638;
  wire       [31:0]   _zz_4639;
  wire       [31:0]   _zz_4640;
  wire       [31:0]   _zz_4641;
  wire       [31:0]   _zz_4642;
  wire       [31:0]   _zz_4643;
  wire       [31:0]   _zz_4644;
  wire       [31:0]   _zz_4645;
  wire       [31:0]   _zz_4646;
  wire       [31:0]   _zz_4647;
  wire       [31:0]   _zz_4648;
  wire       [31:0]   _zz_4649;
  wire       [31:0]   _zz_4650;
  wire       [31:0]   _zz_4651;
  wire       [31:0]   _zz_4652;
  wire       [31:0]   _zz_4653;
  wire       [31:0]   _zz_4654;
  wire       [31:0]   _zz_4655;
  wire       [31:0]   _zz_4656;
  wire       [31:0]   _zz_4657;
  wire       [31:0]   _zz_4658;
  wire       [31:0]   _zz_4659;
  wire       [31:0]   _zz_4660;
  wire       [31:0]   _zz_4661;
  wire       [31:0]   _zz_4662;
  wire       [31:0]   _zz_4663;
  wire       [31:0]   _zz_4664;
  wire       [31:0]   _zz_4665;
  wire       [31:0]   _zz_4666;
  wire       [31:0]   _zz_4667;
  wire       [31:0]   _zz_4668;
  wire       [31:0]   _zz_4669;
  wire       [31:0]   _zz_4670;
  wire       [31:0]   _zz_4671;
  wire       [31:0]   _zz_4672;
  wire       [31:0]   _zz_4673;
  wire       [31:0]   _zz_4674;
  wire       [31:0]   _zz_4675;
  wire       [31:0]   _zz_4676;
  wire       [31:0]   _zz_4677;
  wire       [31:0]   _zz_4678;
  wire       [31:0]   _zz_4679;
  wire       [31:0]   _zz_4680;
  wire       [31:0]   _zz_4681;
  wire       [31:0]   _zz_4682;
  wire       [31:0]   _zz_4683;
  wire       [31:0]   _zz_4684;
  wire       [31:0]   _zz_4685;
  wire       [31:0]   _zz_4686;
  wire       [31:0]   _zz_4687;
  wire       [31:0]   _zz_4688;
  wire       [31:0]   _zz_4689;
  wire       [31:0]   _zz_4690;
  wire       [31:0]   _zz_4691;
  wire       [31:0]   _zz_4692;
  wire       [31:0]   _zz_4693;
  wire       [31:0]   _zz_4694;
  wire       [31:0]   _zz_4695;
  wire       [31:0]   _zz_4696;
  wire       [31:0]   _zz_4697;
  wire       [31:0]   _zz_4698;
  wire       [31:0]   _zz_4699;
  wire       [31:0]   _zz_4700;
  wire       [31:0]   _zz_4701;
  wire       [31:0]   _zz_4702;
  wire       [31:0]   _zz_4703;
  wire       [31:0]   _zz_4704;
  wire       [31:0]   _zz_4705;
  wire       [31:0]   _zz_4706;
  wire       [31:0]   _zz_4707;
  wire       [31:0]   _zz_4708;
  wire       [31:0]   _zz_4709;
  wire       [31:0]   _zz_4710;
  wire       [31:0]   _zz_4711;
  wire       [31:0]   _zz_4712;
  wire       [31:0]   _zz_4713;
  wire       [31:0]   _zz_4714;
  wire       [31:0]   _zz_4715;
  wire       [31:0]   _zz_4716;
  wire       [31:0]   _zz_4717;
  wire       [31:0]   _zz_4718;
  wire       [31:0]   _zz_4719;
  wire       [31:0]   _zz_4720;
  wire       [31:0]   _zz_4721;
  wire       [31:0]   _zz_4722;
  wire       [31:0]   _zz_4723;
  wire       [31:0]   _zz_4724;
  wire       [31:0]   _zz_4725;
  wire       [31:0]   _zz_4726;
  wire       [31:0]   _zz_4727;
  wire       [31:0]   _zz_4728;
  wire       [31:0]   _zz_4729;
  wire       [31:0]   _zz_4730;
  wire       [31:0]   _zz_4731;
  wire       [31:0]   _zz_4732;
  wire       [31:0]   _zz_4733;
  wire       [31:0]   _zz_4734;
  wire       [31:0]   _zz_4735;
  wire       [31:0]   _zz_4736;
  wire       [31:0]   _zz_4737;
  wire       [31:0]   _zz_4738;
  wire       [31:0]   _zz_4739;
  wire       [31:0]   _zz_4740;
  wire       [31:0]   _zz_4741;
  wire       [31:0]   _zz_4742;
  wire       [31:0]   _zz_4743;
  wire       [31:0]   _zz_4744;
  wire       [31:0]   _zz_4745;
  wire       [31:0]   _zz_4746;
  wire       [31:0]   _zz_4747;
  wire       [31:0]   _zz_4748;
  wire       [31:0]   _zz_4749;
  wire       [31:0]   _zz_4750;
  wire       [31:0]   _zz_4751;
  wire       [31:0]   _zz_4752;
  wire       [31:0]   _zz_4753;
  wire       [31:0]   _zz_4754;
  wire       [31:0]   _zz_4755;
  wire       [31:0]   _zz_4756;
  wire       [31:0]   _zz_4757;
  wire       [31:0]   _zz_4758;
  wire       [31:0]   _zz_4759;
  wire       [31:0]   _zz_4760;
  wire       [31:0]   _zz_4761;
  wire       [31:0]   _zz_4762;
  wire       [31:0]   _zz_4763;
  wire       [31:0]   _zz_4764;
  wire       [31:0]   _zz_4765;
  wire       [31:0]   _zz_4766;
  wire       [31:0]   _zz_4767;
  wire       [31:0]   _zz_4768;
  wire       [31:0]   _zz_4769;
  wire       [31:0]   _zz_4770;
  wire       [31:0]   _zz_4771;
  wire       [31:0]   _zz_4772;
  wire       [31:0]   _zz_4773;
  wire       [31:0]   _zz_4774;
  wire       [31:0]   _zz_4775;
  wire       [31:0]   _zz_4776;
  wire       [31:0]   _zz_4777;
  wire       [31:0]   _zz_4778;
  wire       [31:0]   _zz_4779;
  wire       [31:0]   _zz_4780;
  wire       [31:0]   _zz_4781;
  wire       [31:0]   _zz_4782;
  wire       [31:0]   _zz_4783;
  wire       [31:0]   _zz_4784;
  wire       [31:0]   _zz_4785;
  wire       [31:0]   _zz_4786;
  wire       [31:0]   _zz_4787;
  wire       [31:0]   _zz_4788;
  wire       [31:0]   _zz_4789;
  wire       [31:0]   _zz_4790;
  wire       [31:0]   _zz_4791;
  wire       [31:0]   _zz_4792;
  wire       [31:0]   _zz_4793;
  wire       [31:0]   _zz_4794;
  wire       [31:0]   _zz_4795;
  wire       [31:0]   _zz_4796;
  wire       [31:0]   _zz_4797;
  wire       [31:0]   _zz_4798;
  wire       [31:0]   _zz_4799;
  wire       [31:0]   _zz_4800;
  wire       [31:0]   _zz_4801;
  wire       [31:0]   _zz_4802;
  wire       [31:0]   _zz_4803;
  wire       [31:0]   _zz_4804;
  wire       [31:0]   _zz_4805;
  wire       [31:0]   _zz_4806;
  wire       [31:0]   _zz_4807;
  wire       [31:0]   _zz_4808;
  wire       [31:0]   _zz_4809;
  wire       [31:0]   _zz_4810;
  wire       [31:0]   _zz_4811;
  wire       [31:0]   _zz_4812;
  wire       [31:0]   _zz_4813;
  wire       [31:0]   _zz_4814;
  wire       [31:0]   _zz_4815;
  wire       [31:0]   _zz_4816;
  wire       [31:0]   _zz_4817;
  wire       [31:0]   _zz_4818;
  wire       [31:0]   _zz_4819;
  wire       [31:0]   _zz_4820;
  wire       [31:0]   _zz_4821;
  wire       [31:0]   _zz_4822;
  wire       [31:0]   _zz_4823;
  wire       [31:0]   _zz_4824;
  wire       [31:0]   _zz_4825;
  wire       [31:0]   _zz_4826;
  wire       [31:0]   _zz_4827;
  wire       [31:0]   _zz_4828;
  wire       [31:0]   _zz_4829;
  wire       [31:0]   _zz_4830;
  wire       [31:0]   _zz_4831;
  wire       [31:0]   _zz_4832;
  wire       [31:0]   _zz_4833;
  wire       [31:0]   _zz_4834;
  wire       [31:0]   _zz_4835;
  wire       [31:0]   _zz_4836;
  wire       [31:0]   _zz_4837;
  wire       [31:0]   _zz_4838;
  wire       [31:0]   _zz_4839;
  wire       [31:0]   _zz_4840;
  wire       [31:0]   _zz_4841;
  wire       [31:0]   _zz_4842;
  wire       [31:0]   _zz_4843;
  wire       [31:0]   _zz_4844;
  wire       [31:0]   _zz_4845;
  wire       [31:0]   _zz_4846;
  wire       [31:0]   _zz_4847;
  wire       [31:0]   _zz_4848;
  wire       [31:0]   _zz_4849;
  wire       [31:0]   _zz_4850;
  wire       [31:0]   _zz_4851;
  wire       [31:0]   _zz_4852;
  wire       [31:0]   _zz_4853;
  wire       [31:0]   _zz_4854;
  wire       [31:0]   _zz_4855;
  wire       [31:0]   _zz_4856;
  wire       [31:0]   _zz_4857;
  wire       [31:0]   _zz_4858;
  wire       [31:0]   _zz_4859;
  wire       [31:0]   _zz_4860;
  wire       [31:0]   _zz_4861;
  wire       [31:0]   _zz_4862;
  wire       [31:0]   _zz_4863;
  wire       [31:0]   _zz_4864;
  wire       [31:0]   _zz_4865;
  wire       [31:0]   _zz_4866;
  wire       [31:0]   _zz_4867;
  wire       [31:0]   _zz_4868;
  wire       [31:0]   _zz_4869;
  wire       [31:0]   _zz_4870;
  wire       [31:0]   _zz_4871;
  wire       [31:0]   _zz_4872;
  wire       [31:0]   _zz_4873;
  wire       [31:0]   _zz_4874;
  wire       [31:0]   _zz_4875;
  wire       [31:0]   _zz_4876;
  wire       [31:0]   _zz_4877;
  wire       [31:0]   _zz_4878;
  wire       [31:0]   _zz_4879;
  wire       [31:0]   _zz_4880;
  wire       [31:0]   _zz_4881;
  wire       [31:0]   _zz_4882;
  wire       [31:0]   _zz_4883;
  wire       [31:0]   _zz_4884;
  wire       [31:0]   _zz_4885;
  wire       [31:0]   _zz_4886;
  wire       [31:0]   _zz_4887;
  wire       [31:0]   _zz_4888;
  wire       [31:0]   _zz_4889;
  wire       [31:0]   _zz_4890;
  wire       [31:0]   _zz_4891;
  wire       [31:0]   _zz_4892;
  wire       [31:0]   _zz_4893;
  wire       [31:0]   _zz_4894;
  wire       [31:0]   _zz_4895;
  wire       [31:0]   _zz_4896;
  wire       [31:0]   _zz_4897;
  wire       [31:0]   _zz_4898;
  wire       [31:0]   _zz_4899;
  wire       [31:0]   _zz_4900;
  wire       [31:0]   _zz_4901;
  wire       [31:0]   _zz_4902;
  wire       [31:0]   _zz_4903;
  wire       [31:0]   _zz_4904;
  wire       [31:0]   _zz_4905;
  wire       [31:0]   _zz_4906;
  wire       [31:0]   _zz_4907;
  wire       [31:0]   _zz_4908;
  wire       [31:0]   _zz_4909;
  wire       [31:0]   _zz_4910;
  wire       [31:0]   _zz_4911;
  wire       [31:0]   _zz_4912;
  wire       [31:0]   _zz_4913;
  wire       [31:0]   _zz_4914;
  wire       [31:0]   _zz_4915;
  wire       [31:0]   _zz_4916;
  wire       [31:0]   _zz_4917;
  wire       [31:0]   _zz_4918;
  wire       [31:0]   _zz_4919;
  wire       [31:0]   _zz_4920;
  wire       [31:0]   _zz_4921;
  wire       [31:0]   _zz_4922;
  wire       [31:0]   _zz_4923;
  wire       [31:0]   _zz_4924;
  wire       [31:0]   _zz_4925;
  wire       [31:0]   _zz_4926;
  wire       [31:0]   _zz_4927;
  wire       [31:0]   _zz_4928;
  wire       [31:0]   _zz_4929;
  wire       [31:0]   _zz_4930;
  wire       [31:0]   _zz_4931;
  wire       [31:0]   _zz_4932;
  wire       [31:0]   _zz_4933;
  wire       [31:0]   _zz_4934;
  wire       [31:0]   _zz_4935;
  wire       [31:0]   _zz_4936;
  wire       [31:0]   _zz_4937;
  wire       [31:0]   _zz_4938;
  wire       [31:0]   _zz_4939;
  wire       [31:0]   _zz_4940;
  wire       [31:0]   _zz_4941;
  wire       [31:0]   _zz_4942;
  wire       [31:0]   _zz_4943;
  wire       [31:0]   _zz_4944;
  wire       [31:0]   _zz_4945;
  wire       [31:0]   _zz_4946;
  wire       [31:0]   _zz_4947;
  wire       [31:0]   _zz_4948;
  wire       [31:0]   _zz_4949;
  wire       [31:0]   _zz_4950;
  wire       [31:0]   _zz_4951;
  wire       [31:0]   _zz_4952;
  wire       [31:0]   _zz_4953;
  wire       [31:0]   _zz_4954;
  wire       [31:0]   _zz_4955;
  wire       [31:0]   _zz_4956;
  wire       [31:0]   _zz_4957;
  wire       [31:0]   _zz_4958;
  wire       [31:0]   _zz_4959;
  wire       [31:0]   _zz_4960;
  wire       [31:0]   _zz_4961;
  wire       [31:0]   _zz_4962;
  wire       [31:0]   _zz_4963;
  wire       [31:0]   _zz_4964;
  wire       [31:0]   _zz_4965;
  wire       [31:0]   _zz_4966;
  wire       [31:0]   _zz_4967;
  wire       [31:0]   _zz_4968;
  wire       [31:0]   _zz_4969;
  wire       [31:0]   _zz_4970;
  wire       [31:0]   _zz_4971;
  wire       [31:0]   _zz_4972;
  wire       [31:0]   _zz_4973;
  wire       [31:0]   _zz_4974;
  wire       [31:0]   _zz_4975;
  wire       [31:0]   _zz_4976;
  wire       [31:0]   _zz_4977;
  wire       [31:0]   _zz_4978;
  wire       [31:0]   _zz_4979;
  wire       [31:0]   _zz_4980;
  wire       [31:0]   _zz_4981;
  wire       [31:0]   _zz_4982;
  wire       [31:0]   _zz_4983;
  wire       [31:0]   _zz_4984;
  wire       [31:0]   _zz_4985;
  wire       [31:0]   _zz_4986;
  wire       [31:0]   _zz_4987;
  wire       [31:0]   _zz_4988;
  wire       [31:0]   _zz_4989;
  wire       [31:0]   _zz_4990;
  wire       [31:0]   _zz_4991;
  wire       [31:0]   _zz_4992;
  wire       [31:0]   _zz_4993;
  wire       [31:0]   _zz_4994;
  wire       [31:0]   _zz_4995;
  wire       [31:0]   _zz_4996;
  wire       [31:0]   _zz_4997;
  wire       [31:0]   _zz_4998;
  wire       [31:0]   _zz_4999;
  wire       [31:0]   _zz_5000;
  wire       [31:0]   _zz_5001;
  wire       [31:0]   _zz_5002;
  wire       [31:0]   _zz_5003;
  wire       [31:0]   _zz_5004;
  wire       [31:0]   _zz_5005;
  wire       [31:0]   _zz_5006;
  wire       [31:0]   _zz_5007;
  wire       [31:0]   _zz_5008;
  wire       [31:0]   _zz_5009;
  wire       [31:0]   _zz_5010;
  wire       [31:0]   _zz_5011;
  wire       [31:0]   _zz_5012;
  wire       [31:0]   _zz_5013;
  wire       [31:0]   _zz_5014;
  wire       [31:0]   _zz_5015;
  wire       [31:0]   _zz_5016;
  wire       [31:0]   _zz_5017;
  wire       [31:0]   _zz_5018;
  wire       [31:0]   _zz_5019;
  wire       [31:0]   _zz_5020;
  wire       [31:0]   _zz_5021;
  wire       [31:0]   _zz_5022;
  wire       [31:0]   _zz_5023;
  wire       [31:0]   _zz_5024;
  wire       [31:0]   _zz_5025;
  wire       [31:0]   _zz_5026;
  wire       [31:0]   _zz_5027;
  wire       [31:0]   _zz_5028;
  wire       [31:0]   _zz_5029;
  wire       [31:0]   _zz_5030;
  wire       [31:0]   _zz_5031;
  wire       [31:0]   _zz_5032;
  wire       [31:0]   _zz_5033;
  wire       [31:0]   _zz_5034;
  wire       [31:0]   _zz_5035;
  wire       [31:0]   _zz_5036;
  wire       [31:0]   _zz_5037;
  wire       [31:0]   _zz_5038;
  wire       [31:0]   _zz_5039;
  wire       [31:0]   _zz_5040;
  wire       [31:0]   _zz_5041;
  wire       [31:0]   _zz_5042;
  wire       [31:0]   _zz_5043;
  wire       [31:0]   _zz_5044;
  wire       [31:0]   _zz_5045;
  wire       [31:0]   _zz_5046;
  wire       [31:0]   _zz_5047;
  wire       [31:0]   _zz_5048;
  wire       [31:0]   _zz_5049;
  wire       [31:0]   _zz_5050;
  wire       [31:0]   _zz_5051;
  wire       [31:0]   _zz_5052;
  wire       [31:0]   _zz_5053;
  wire       [31:0]   _zz_5054;
  wire       [31:0]   _zz_5055;
  wire       [31:0]   _zz_5056;
  wire       [31:0]   _zz_5057;
  wire       [31:0]   _zz_5058;
  wire       [31:0]   _zz_5059;
  wire       [31:0]   _zz_5060;
  wire       [31:0]   _zz_5061;
  wire       [31:0]   _zz_5062;
  wire       [31:0]   _zz_5063;
  wire       [31:0]   _zz_5064;
  wire       [31:0]   _zz_5065;
  wire       [31:0]   _zz_5066;
  wire       [31:0]   _zz_5067;
  wire       [31:0]   _zz_5068;
  wire       [31:0]   _zz_5069;
  wire       [31:0]   _zz_5070;
  wire       [31:0]   _zz_5071;
  wire       [31:0]   _zz_5072;
  wire       [31:0]   _zz_5073;
  wire       [31:0]   _zz_5074;
  wire       [31:0]   _zz_5075;
  wire       [31:0]   _zz_5076;
  wire       [31:0]   _zz_5077;
  wire       [31:0]   _zz_5078;
  wire       [31:0]   _zz_5079;
  wire       [31:0]   _zz_5080;
  wire       [31:0]   _zz_5081;
  wire       [31:0]   _zz_5082;
  wire       [31:0]   _zz_5083;
  wire       [31:0]   _zz_5084;
  wire       [31:0]   _zz_5085;
  wire       [31:0]   _zz_5086;
  wire       [31:0]   _zz_5087;
  wire       [31:0]   _zz_5088;
  wire       [31:0]   _zz_5089;
  wire       [31:0]   _zz_5090;
  wire       [31:0]   _zz_5091;
  wire       [31:0]   _zz_5092;
  wire       [31:0]   _zz_5093;
  wire       [31:0]   _zz_5094;
  wire       [31:0]   _zz_5095;
  wire       [31:0]   _zz_5096;
  wire       [31:0]   _zz_5097;
  wire       [31:0]   _zz_5098;
  wire       [31:0]   _zz_5099;
  wire       [31:0]   _zz_5100;
  wire       [31:0]   _zz_5101;
  wire       [31:0]   _zz_5102;
  wire       [31:0]   _zz_5103;
  wire       [31:0]   _zz_5104;
  wire       [31:0]   _zz_5105;
  wire       [31:0]   _zz_5106;
  wire       [31:0]   _zz_5107;
  wire       [31:0]   _zz_5108;
  wire       [31:0]   _zz_5109;
  wire       [31:0]   _zz_5110;
  wire       [31:0]   _zz_5111;
  wire       [31:0]   _zz_5112;
  wire       [31:0]   _zz_5113;
  wire       [31:0]   _zz_5114;
  wire       [31:0]   _zz_5115;
  wire       [31:0]   _zz_5116;
  wire       [31:0]   _zz_5117;
  wire       [31:0]   _zz_5118;
  wire       [31:0]   _zz_5119;
  wire       [31:0]   _zz_5120;
  wire       [31:0]   _zz_5121;
  wire       [31:0]   _zz_5122;
  wire       [31:0]   _zz_5123;
  wire       [31:0]   _zz_5124;
  wire       [31:0]   _zz_5125;
  wire       [31:0]   _zz_5126;
  wire       [31:0]   _zz_5127;
  wire       [31:0]   _zz_5128;
  wire       [31:0]   _zz_5129;
  wire       [31:0]   _zz_5130;
  wire       [31:0]   _zz_5131;
  wire       [31:0]   _zz_5132;
  wire       [31:0]   _zz_5133;
  wire       [31:0]   _zz_5134;
  wire       [31:0]   _zz_5135;
  wire       [31:0]   _zz_5136;
  wire       [31:0]   _zz_5137;
  wire       [31:0]   _zz_5138;
  wire       [31:0]   _zz_5139;
  wire       [31:0]   _zz_5140;
  wire       [31:0]   _zz_5141;
  wire       [31:0]   _zz_5142;
  wire       [31:0]   _zz_5143;
  wire       [31:0]   _zz_5144;
  wire       [31:0]   _zz_5145;
  wire       [31:0]   _zz_5146;
  wire       [31:0]   _zz_5147;
  wire       [31:0]   _zz_5148;
  wire       [31:0]   _zz_5149;
  wire       [31:0]   _zz_5150;
  wire       [31:0]   _zz_5151;
  wire       [31:0]   _zz_5152;
  wire       [31:0]   _zz_5153;
  wire       [31:0]   _zz_5154;
  wire       [31:0]   _zz_5155;
  wire       [31:0]   _zz_5156;
  wire       [31:0]   _zz_5157;
  wire       [31:0]   _zz_5158;
  wire       [31:0]   _zz_5159;
  wire       [31:0]   _zz_5160;
  wire       [31:0]   _zz_5161;
  wire       [31:0]   _zz_5162;
  wire       [31:0]   _zz_5163;
  wire       [31:0]   _zz_5164;
  wire       [31:0]   _zz_5165;
  wire       [31:0]   _zz_5166;
  wire       [31:0]   _zz_5167;
  wire       [31:0]   _zz_5168;
  wire       [31:0]   _zz_5169;
  wire       [31:0]   _zz_5170;
  wire       [31:0]   _zz_5171;
  wire       [31:0]   _zz_5172;
  wire       [31:0]   _zz_5173;
  wire       [31:0]   _zz_5174;
  wire       [31:0]   _zz_5175;
  wire       [31:0]   _zz_5176;
  wire       [31:0]   _zz_5177;
  wire       [31:0]   _zz_5178;
  wire       [31:0]   _zz_5179;
  wire       [31:0]   _zz_5180;
  wire       [31:0]   _zz_5181;
  wire       [31:0]   _zz_5182;
  wire       [31:0]   _zz_5183;
  wire       [31:0]   _zz_5184;
  wire       [31:0]   _zz_5185;
  wire       [31:0]   _zz_5186;
  wire       [31:0]   _zz_5187;
  wire       [31:0]   _zz_5188;
  wire       [31:0]   _zz_5189;
  wire       [31:0]   _zz_5190;
  wire       [31:0]   _zz_5191;
  wire       [31:0]   _zz_5192;
  wire       [31:0]   _zz_5193;
  wire       [31:0]   _zz_5194;
  wire       [31:0]   _zz_5195;
  wire       [31:0]   _zz_5196;
  wire       [31:0]   _zz_5197;
  wire       [31:0]   _zz_5198;
  wire       [31:0]   _zz_5199;
  wire       [31:0]   _zz_5200;
  wire       [31:0]   _zz_5201;
  wire       [31:0]   _zz_5202;
  wire       [31:0]   _zz_5203;
  wire       [31:0]   _zz_5204;
  wire       [31:0]   _zz_5205;
  wire       [31:0]   _zz_5206;
  wire       [31:0]   _zz_5207;
  wire       [31:0]   _zz_5208;
  wire       [31:0]   _zz_5209;
  wire       [31:0]   _zz_5210;
  wire       [31:0]   _zz_5211;
  wire       [31:0]   _zz_5212;
  wire       [31:0]   _zz_5213;
  wire       [31:0]   _zz_5214;
  wire       [31:0]   _zz_5215;
  wire       [31:0]   _zz_5216;
  wire       [31:0]   _zz_5217;
  wire       [31:0]   _zz_5218;
  wire       [31:0]   _zz_5219;
  wire       [31:0]   _zz_5220;
  wire       [31:0]   _zz_5221;
  wire       [31:0]   _zz_5222;
  wire       [31:0]   _zz_5223;
  wire       [31:0]   _zz_5224;
  wire       [31:0]   _zz_5225;
  wire       [31:0]   _zz_5226;
  wire       [31:0]   _zz_5227;
  wire       [31:0]   _zz_5228;
  wire       [31:0]   _zz_5229;
  wire       [31:0]   _zz_5230;
  wire       [31:0]   _zz_5231;
  wire       [31:0]   _zz_5232;
  wire       [31:0]   _zz_5233;
  wire       [31:0]   _zz_5234;
  wire       [31:0]   _zz_5235;
  wire       [31:0]   _zz_5236;
  wire       [31:0]   _zz_5237;
  wire       [31:0]   _zz_5238;
  wire       [31:0]   _zz_5239;
  wire       [31:0]   _zz_5240;
  wire       [31:0]   _zz_5241;
  wire       [31:0]   _zz_5242;
  wire       [31:0]   _zz_5243;
  wire       [31:0]   _zz_5244;
  wire       [31:0]   _zz_5245;
  wire       [31:0]   _zz_5246;
  wire       [31:0]   _zz_5247;
  wire       [31:0]   _zz_5248;
  wire       [31:0]   _zz_5249;
  wire       [31:0]   _zz_5250;
  wire       [31:0]   _zz_5251;
  wire       [31:0]   _zz_5252;
  wire       [31:0]   _zz_5253;
  wire       [31:0]   _zz_5254;
  wire       [31:0]   _zz_5255;
  wire       [31:0]   _zz_5256;
  wire       [31:0]   _zz_5257;
  wire       [31:0]   _zz_5258;
  wire       [31:0]   _zz_5259;
  wire       [31:0]   _zz_5260;
  wire       [31:0]   _zz_5261;
  wire       [31:0]   _zz_5262;
  wire       [31:0]   _zz_5263;
  wire       [31:0]   _zz_5264;
  wire       [31:0]   _zz_5265;
  wire       [31:0]   _zz_5266;
  wire       [31:0]   _zz_5267;
  wire       [31:0]   _zz_5268;
  wire       [31:0]   _zz_5269;
  wire       [31:0]   _zz_5270;
  wire       [31:0]   _zz_5271;
  wire       [31:0]   _zz_5272;
  wire       [31:0]   _zz_5273;
  wire       [31:0]   _zz_5274;
  wire       [31:0]   _zz_5275;
  wire       [31:0]   _zz_5276;
  wire       [31:0]   _zz_5277;
  wire       [31:0]   _zz_5278;
  wire       [31:0]   _zz_5279;
  wire       [31:0]   _zz_5280;
  wire       [31:0]   _zz_5281;
  wire       [31:0]   _zz_5282;
  wire       [31:0]   _zz_5283;
  wire       [31:0]   _zz_5284;
  wire       [31:0]   _zz_5285;
  wire       [31:0]   _zz_5286;
  wire       [31:0]   _zz_5287;
  wire       [31:0]   _zz_5288;
  wire       [31:0]   _zz_5289;
  wire       [31:0]   _zz_5290;
  wire       [31:0]   _zz_5291;
  wire       [31:0]   _zz_5292;
  wire       [31:0]   _zz_5293;
  wire       [31:0]   _zz_5294;
  wire       [31:0]   _zz_5295;
  wire       [31:0]   _zz_5296;
  wire       [31:0]   _zz_5297;
  wire       [31:0]   _zz_5298;
  wire       [31:0]   _zz_5299;
  wire       [31:0]   _zz_5300;
  wire       [31:0]   _zz_5301;
  wire       [31:0]   _zz_5302;
  wire       [31:0]   _zz_5303;
  wire       [31:0]   _zz_5304;
  wire       [31:0]   _zz_5305;
  wire       [31:0]   _zz_5306;
  wire       [31:0]   _zz_5307;
  wire       [31:0]   _zz_5308;
  wire       [31:0]   _zz_5309;
  wire       [31:0]   _zz_5310;
  wire       [31:0]   _zz_5311;
  wire       [31:0]   _zz_5312;
  wire       [31:0]   _zz_5313;
  wire       [31:0]   _zz_5314;
  wire       [31:0]   _zz_5315;
  wire       [31:0]   _zz_5316;
  wire       [31:0]   _zz_5317;
  wire       [31:0]   _zz_5318;
  wire       [31:0]   _zz_5319;
  wire       [31:0]   _zz_5320;
  wire       [31:0]   _zz_5321;
  wire       [31:0]   _zz_5322;
  wire       [31:0]   _zz_5323;
  wire       [31:0]   _zz_5324;
  wire       [31:0]   _zz_5325;
  wire       [31:0]   _zz_5326;
  wire       [31:0]   _zz_5327;
  wire       [31:0]   _zz_5328;
  wire       [31:0]   _zz_5329;
  wire       [31:0]   _zz_5330;
  wire       [31:0]   _zz_5331;
  wire       [31:0]   _zz_5332;
  wire       [31:0]   _zz_5333;
  wire       [31:0]   _zz_5334;
  wire       [31:0]   _zz_5335;
  wire       [31:0]   _zz_5336;
  wire       [31:0]   _zz_5337;
  wire       [31:0]   _zz_5338;
  wire       [31:0]   _zz_5339;
  wire       [31:0]   _zz_5340;
  wire       [31:0]   _zz_5341;
  wire       [31:0]   _zz_5342;
  wire       [31:0]   _zz_5343;
  wire       [31:0]   _zz_5344;
  wire       [31:0]   _zz_5345;
  wire       [31:0]   _zz_5346;
  wire       [31:0]   _zz_5347;
  wire       [31:0]   _zz_5348;
  wire       [31:0]   _zz_5349;
  wire       [31:0]   _zz_5350;
  wire       [31:0]   _zz_5351;
  wire       [31:0]   _zz_5352;
  wire       [31:0]   _zz_5353;
  wire       [31:0]   _zz_5354;
  wire       [31:0]   _zz_5355;
  wire       [31:0]   _zz_5356;
  wire       [31:0]   _zz_5357;
  wire       [31:0]   _zz_5358;
  wire       [31:0]   _zz_5359;
  wire       [31:0]   _zz_5360;
  wire       [31:0]   _zz_5361;
  wire       [31:0]   _zz_5362;
  wire       [31:0]   _zz_5363;
  wire       [31:0]   _zz_5364;
  wire       [31:0]   _zz_5365;
  wire       [31:0]   _zz_5366;
  wire       [31:0]   _zz_5367;
  wire       [31:0]   _zz_5368;
  wire       [31:0]   _zz_5369;
  wire       [31:0]   _zz_5370;
  wire       [31:0]   _zz_5371;
  wire       [31:0]   _zz_5372;
  wire       [31:0]   _zz_5373;
  wire       [31:0]   _zz_5374;
  wire       [31:0]   _zz_5375;
  wire       [31:0]   _zz_5376;
  wire       [31:0]   _zz_5377;
  wire       [31:0]   _zz_5378;
  wire       [31:0]   _zz_5379;
  wire       [31:0]   _zz_5380;
  wire       [31:0]   _zz_5381;
  wire       [31:0]   _zz_5382;
  wire       [15:0]   fixTo_dout;
  wire       [15:0]   fixTo_1_dout;
  wire       [15:0]   fixTo_2_dout;
  wire       [15:0]   fixTo_3_dout;
  wire       [15:0]   fixTo_4_dout;
  wire       [15:0]   fixTo_5_dout;
  wire       [15:0]   fixTo_6_dout;
  wire       [15:0]   fixTo_7_dout;
  wire       [15:0]   fixTo_8_dout;
  wire       [15:0]   fixTo_9_dout;
  wire       [15:0]   fixTo_10_dout;
  wire       [15:0]   fixTo_11_dout;
  wire       [15:0]   fixTo_12_dout;
  wire       [15:0]   fixTo_13_dout;
  wire       [15:0]   fixTo_14_dout;
  wire       [15:0]   fixTo_15_dout;
  wire       [15:0]   fixTo_16_dout;
  wire       [15:0]   fixTo_17_dout;
  wire       [15:0]   fixTo_18_dout;
  wire       [15:0]   fixTo_19_dout;
  wire       [15:0]   fixTo_20_dout;
  wire       [15:0]   fixTo_21_dout;
  wire       [15:0]   fixTo_22_dout;
  wire       [15:0]   fixTo_23_dout;
  wire       [15:0]   fixTo_24_dout;
  wire       [15:0]   fixTo_25_dout;
  wire       [15:0]   fixTo_26_dout;
  wire       [15:0]   fixTo_27_dout;
  wire       [15:0]   fixTo_28_dout;
  wire       [15:0]   fixTo_29_dout;
  wire       [15:0]   fixTo_30_dout;
  wire       [15:0]   fixTo_31_dout;
  wire       [15:0]   fixTo_32_dout;
  wire       [15:0]   fixTo_33_dout;
  wire       [15:0]   fixTo_34_dout;
  wire       [15:0]   fixTo_35_dout;
  wire       [15:0]   fixTo_36_dout;
  wire       [15:0]   fixTo_37_dout;
  wire       [15:0]   fixTo_38_dout;
  wire       [15:0]   fixTo_39_dout;
  wire       [15:0]   fixTo_40_dout;
  wire       [15:0]   fixTo_41_dout;
  wire       [15:0]   fixTo_42_dout;
  wire       [15:0]   fixTo_43_dout;
  wire       [15:0]   fixTo_44_dout;
  wire       [15:0]   fixTo_45_dout;
  wire       [15:0]   fixTo_46_dout;
  wire       [15:0]   fixTo_47_dout;
  wire       [15:0]   fixTo_48_dout;
  wire       [15:0]   fixTo_49_dout;
  wire       [15:0]   fixTo_50_dout;
  wire       [15:0]   fixTo_51_dout;
  wire       [15:0]   fixTo_52_dout;
  wire       [15:0]   fixTo_53_dout;
  wire       [15:0]   fixTo_54_dout;
  wire       [15:0]   fixTo_55_dout;
  wire       [15:0]   fixTo_56_dout;
  wire       [15:0]   fixTo_57_dout;
  wire       [15:0]   fixTo_58_dout;
  wire       [15:0]   fixTo_59_dout;
  wire       [15:0]   fixTo_60_dout;
  wire       [15:0]   fixTo_61_dout;
  wire       [15:0]   fixTo_62_dout;
  wire       [15:0]   fixTo_63_dout;
  wire       [15:0]   fixTo_64_dout;
  wire       [15:0]   fixTo_65_dout;
  wire       [15:0]   fixTo_66_dout;
  wire       [15:0]   fixTo_67_dout;
  wire       [15:0]   fixTo_68_dout;
  wire       [15:0]   fixTo_69_dout;
  wire       [15:0]   fixTo_70_dout;
  wire       [15:0]   fixTo_71_dout;
  wire       [15:0]   fixTo_72_dout;
  wire       [15:0]   fixTo_73_dout;
  wire       [15:0]   fixTo_74_dout;
  wire       [15:0]   fixTo_75_dout;
  wire       [15:0]   fixTo_76_dout;
  wire       [15:0]   fixTo_77_dout;
  wire       [15:0]   fixTo_78_dout;
  wire       [15:0]   fixTo_79_dout;
  wire       [15:0]   fixTo_80_dout;
  wire       [15:0]   fixTo_81_dout;
  wire       [15:0]   fixTo_82_dout;
  wire       [15:0]   fixTo_83_dout;
  wire       [15:0]   fixTo_84_dout;
  wire       [15:0]   fixTo_85_dout;
  wire       [15:0]   fixTo_86_dout;
  wire       [15:0]   fixTo_87_dout;
  wire       [15:0]   fixTo_88_dout;
  wire       [15:0]   fixTo_89_dout;
  wire       [15:0]   fixTo_90_dout;
  wire       [15:0]   fixTo_91_dout;
  wire       [15:0]   fixTo_92_dout;
  wire       [15:0]   fixTo_93_dout;
  wire       [15:0]   fixTo_94_dout;
  wire       [15:0]   fixTo_95_dout;
  wire       [15:0]   fixTo_96_dout;
  wire       [15:0]   fixTo_97_dout;
  wire       [15:0]   fixTo_98_dout;
  wire       [15:0]   fixTo_99_dout;
  wire       [15:0]   fixTo_100_dout;
  wire       [15:0]   fixTo_101_dout;
  wire       [15:0]   fixTo_102_dout;
  wire       [15:0]   fixTo_103_dout;
  wire       [15:0]   fixTo_104_dout;
  wire       [15:0]   fixTo_105_dout;
  wire       [15:0]   fixTo_106_dout;
  wire       [15:0]   fixTo_107_dout;
  wire       [15:0]   fixTo_108_dout;
  wire       [15:0]   fixTo_109_dout;
  wire       [15:0]   fixTo_110_dout;
  wire       [15:0]   fixTo_111_dout;
  wire       [15:0]   fixTo_112_dout;
  wire       [15:0]   fixTo_113_dout;
  wire       [15:0]   fixTo_114_dout;
  wire       [15:0]   fixTo_115_dout;
  wire       [15:0]   fixTo_116_dout;
  wire       [15:0]   fixTo_117_dout;
  wire       [15:0]   fixTo_118_dout;
  wire       [15:0]   fixTo_119_dout;
  wire       [15:0]   fixTo_120_dout;
  wire       [15:0]   fixTo_121_dout;
  wire       [15:0]   fixTo_122_dout;
  wire       [15:0]   fixTo_123_dout;
  wire       [15:0]   fixTo_124_dout;
  wire       [15:0]   fixTo_125_dout;
  wire       [15:0]   fixTo_126_dout;
  wire       [15:0]   fixTo_127_dout;
  wire       [15:0]   fixTo_128_dout;
  wire       [15:0]   fixTo_129_dout;
  wire       [15:0]   fixTo_130_dout;
  wire       [15:0]   fixTo_131_dout;
  wire       [15:0]   fixTo_132_dout;
  wire       [15:0]   fixTo_133_dout;
  wire       [15:0]   fixTo_134_dout;
  wire       [15:0]   fixTo_135_dout;
  wire       [15:0]   fixTo_136_dout;
  wire       [15:0]   fixTo_137_dout;
  wire       [15:0]   fixTo_138_dout;
  wire       [15:0]   fixTo_139_dout;
  wire       [15:0]   fixTo_140_dout;
  wire       [15:0]   fixTo_141_dout;
  wire       [15:0]   fixTo_142_dout;
  wire       [15:0]   fixTo_143_dout;
  wire       [15:0]   fixTo_144_dout;
  wire       [15:0]   fixTo_145_dout;
  wire       [15:0]   fixTo_146_dout;
  wire       [15:0]   fixTo_147_dout;
  wire       [15:0]   fixTo_148_dout;
  wire       [15:0]   fixTo_149_dout;
  wire       [15:0]   fixTo_150_dout;
  wire       [15:0]   fixTo_151_dout;
  wire       [15:0]   fixTo_152_dout;
  wire       [15:0]   fixTo_153_dout;
  wire       [15:0]   fixTo_154_dout;
  wire       [15:0]   fixTo_155_dout;
  wire       [15:0]   fixTo_156_dout;
  wire       [15:0]   fixTo_157_dout;
  wire       [15:0]   fixTo_158_dout;
  wire       [15:0]   fixTo_159_dout;
  wire       [15:0]   fixTo_160_dout;
  wire       [15:0]   fixTo_161_dout;
  wire       [15:0]   fixTo_162_dout;
  wire       [15:0]   fixTo_163_dout;
  wire       [15:0]   fixTo_164_dout;
  wire       [15:0]   fixTo_165_dout;
  wire       [15:0]   fixTo_166_dout;
  wire       [15:0]   fixTo_167_dout;
  wire       [15:0]   fixTo_168_dout;
  wire       [15:0]   fixTo_169_dout;
  wire       [15:0]   fixTo_170_dout;
  wire       [15:0]   fixTo_171_dout;
  wire       [15:0]   fixTo_172_dout;
  wire       [15:0]   fixTo_173_dout;
  wire       [15:0]   fixTo_174_dout;
  wire       [15:0]   fixTo_175_dout;
  wire       [15:0]   fixTo_176_dout;
  wire       [15:0]   fixTo_177_dout;
  wire       [15:0]   fixTo_178_dout;
  wire       [15:0]   fixTo_179_dout;
  wire       [15:0]   fixTo_180_dout;
  wire       [15:0]   fixTo_181_dout;
  wire       [15:0]   fixTo_182_dout;
  wire       [15:0]   fixTo_183_dout;
  wire       [15:0]   fixTo_184_dout;
  wire       [15:0]   fixTo_185_dout;
  wire       [15:0]   fixTo_186_dout;
  wire       [15:0]   fixTo_187_dout;
  wire       [15:0]   fixTo_188_dout;
  wire       [15:0]   fixTo_189_dout;
  wire       [15:0]   fixTo_190_dout;
  wire       [15:0]   fixTo_191_dout;
  wire       [15:0]   fixTo_192_dout;
  wire       [15:0]   fixTo_193_dout;
  wire       [15:0]   fixTo_194_dout;
  wire       [15:0]   fixTo_195_dout;
  wire       [15:0]   fixTo_196_dout;
  wire       [15:0]   fixTo_197_dout;
  wire       [15:0]   fixTo_198_dout;
  wire       [15:0]   fixTo_199_dout;
  wire       [15:0]   fixTo_200_dout;
  wire       [15:0]   fixTo_201_dout;
  wire       [15:0]   fixTo_202_dout;
  wire       [15:0]   fixTo_203_dout;
  wire       [15:0]   fixTo_204_dout;
  wire       [15:0]   fixTo_205_dout;
  wire       [15:0]   fixTo_206_dout;
  wire       [15:0]   fixTo_207_dout;
  wire       [15:0]   fixTo_208_dout;
  wire       [15:0]   fixTo_209_dout;
  wire       [15:0]   fixTo_210_dout;
  wire       [15:0]   fixTo_211_dout;
  wire       [15:0]   fixTo_212_dout;
  wire       [15:0]   fixTo_213_dout;
  wire       [15:0]   fixTo_214_dout;
  wire       [15:0]   fixTo_215_dout;
  wire       [15:0]   fixTo_216_dout;
  wire       [15:0]   fixTo_217_dout;
  wire       [15:0]   fixTo_218_dout;
  wire       [15:0]   fixTo_219_dout;
  wire       [15:0]   fixTo_220_dout;
  wire       [15:0]   fixTo_221_dout;
  wire       [15:0]   fixTo_222_dout;
  wire       [15:0]   fixTo_223_dout;
  wire       [15:0]   fixTo_224_dout;
  wire       [15:0]   fixTo_225_dout;
  wire       [15:0]   fixTo_226_dout;
  wire       [15:0]   fixTo_227_dout;
  wire       [15:0]   fixTo_228_dout;
  wire       [15:0]   fixTo_229_dout;
  wire       [15:0]   fixTo_230_dout;
  wire       [15:0]   fixTo_231_dout;
  wire       [15:0]   fixTo_232_dout;
  wire       [15:0]   fixTo_233_dout;
  wire       [15:0]   fixTo_234_dout;
  wire       [15:0]   fixTo_235_dout;
  wire       [15:0]   fixTo_236_dout;
  wire       [15:0]   fixTo_237_dout;
  wire       [15:0]   fixTo_238_dout;
  wire       [15:0]   fixTo_239_dout;
  wire       [15:0]   fixTo_240_dout;
  wire       [15:0]   fixTo_241_dout;
  wire       [15:0]   fixTo_242_dout;
  wire       [15:0]   fixTo_243_dout;
  wire       [15:0]   fixTo_244_dout;
  wire       [15:0]   fixTo_245_dout;
  wire       [15:0]   fixTo_246_dout;
  wire       [15:0]   fixTo_247_dout;
  wire       [15:0]   fixTo_248_dout;
  wire       [15:0]   fixTo_249_dout;
  wire       [15:0]   fixTo_250_dout;
  wire       [15:0]   fixTo_251_dout;
  wire       [15:0]   fixTo_252_dout;
  wire       [15:0]   fixTo_253_dout;
  wire       [15:0]   fixTo_254_dout;
  wire       [15:0]   fixTo_255_dout;
  wire       [15:0]   fixTo_256_dout;
  wire       [15:0]   fixTo_257_dout;
  wire       [15:0]   fixTo_258_dout;
  wire       [15:0]   fixTo_259_dout;
  wire       [15:0]   fixTo_260_dout;
  wire       [15:0]   fixTo_261_dout;
  wire       [15:0]   fixTo_262_dout;
  wire       [15:0]   fixTo_263_dout;
  wire       [15:0]   fixTo_264_dout;
  wire       [15:0]   fixTo_265_dout;
  wire       [15:0]   fixTo_266_dout;
  wire       [15:0]   fixTo_267_dout;
  wire       [15:0]   fixTo_268_dout;
  wire       [15:0]   fixTo_269_dout;
  wire       [15:0]   fixTo_270_dout;
  wire       [15:0]   fixTo_271_dout;
  wire       [15:0]   fixTo_272_dout;
  wire       [15:0]   fixTo_273_dout;
  wire       [15:0]   fixTo_274_dout;
  wire       [15:0]   fixTo_275_dout;
  wire       [15:0]   fixTo_276_dout;
  wire       [15:0]   fixTo_277_dout;
  wire       [15:0]   fixTo_278_dout;
  wire       [15:0]   fixTo_279_dout;
  wire       [15:0]   fixTo_280_dout;
  wire       [15:0]   fixTo_281_dout;
  wire       [15:0]   fixTo_282_dout;
  wire       [15:0]   fixTo_283_dout;
  wire       [15:0]   fixTo_284_dout;
  wire       [15:0]   fixTo_285_dout;
  wire       [15:0]   fixTo_286_dout;
  wire       [15:0]   fixTo_287_dout;
  wire       [15:0]   fixTo_288_dout;
  wire       [15:0]   fixTo_289_dout;
  wire       [15:0]   fixTo_290_dout;
  wire       [15:0]   fixTo_291_dout;
  wire       [15:0]   fixTo_292_dout;
  wire       [15:0]   fixTo_293_dout;
  wire       [15:0]   fixTo_294_dout;
  wire       [15:0]   fixTo_295_dout;
  wire       [15:0]   fixTo_296_dout;
  wire       [15:0]   fixTo_297_dout;
  wire       [15:0]   fixTo_298_dout;
  wire       [15:0]   fixTo_299_dout;
  wire       [15:0]   fixTo_300_dout;
  wire       [15:0]   fixTo_301_dout;
  wire       [15:0]   fixTo_302_dout;
  wire       [15:0]   fixTo_303_dout;
  wire       [15:0]   fixTo_304_dout;
  wire       [15:0]   fixTo_305_dout;
  wire       [15:0]   fixTo_306_dout;
  wire       [15:0]   fixTo_307_dout;
  wire       [15:0]   fixTo_308_dout;
  wire       [15:0]   fixTo_309_dout;
  wire       [15:0]   fixTo_310_dout;
  wire       [15:0]   fixTo_311_dout;
  wire       [15:0]   fixTo_312_dout;
  wire       [15:0]   fixTo_313_dout;
  wire       [15:0]   fixTo_314_dout;
  wire       [15:0]   fixTo_315_dout;
  wire       [15:0]   fixTo_316_dout;
  wire       [15:0]   fixTo_317_dout;
  wire       [15:0]   fixTo_318_dout;
  wire       [15:0]   fixTo_319_dout;
  wire       [15:0]   fixTo_320_dout;
  wire       [15:0]   fixTo_321_dout;
  wire       [15:0]   fixTo_322_dout;
  wire       [15:0]   fixTo_323_dout;
  wire       [15:0]   fixTo_324_dout;
  wire       [15:0]   fixTo_325_dout;
  wire       [15:0]   fixTo_326_dout;
  wire       [15:0]   fixTo_327_dout;
  wire       [15:0]   fixTo_328_dout;
  wire       [15:0]   fixTo_329_dout;
  wire       [15:0]   fixTo_330_dout;
  wire       [15:0]   fixTo_331_dout;
  wire       [15:0]   fixTo_332_dout;
  wire       [15:0]   fixTo_333_dout;
  wire       [15:0]   fixTo_334_dout;
  wire       [15:0]   fixTo_335_dout;
  wire       [15:0]   fixTo_336_dout;
  wire       [15:0]   fixTo_337_dout;
  wire       [15:0]   fixTo_338_dout;
  wire       [15:0]   fixTo_339_dout;
  wire       [15:0]   fixTo_340_dout;
  wire       [15:0]   fixTo_341_dout;
  wire       [15:0]   fixTo_342_dout;
  wire       [15:0]   fixTo_343_dout;
  wire       [15:0]   fixTo_344_dout;
  wire       [15:0]   fixTo_345_dout;
  wire       [15:0]   fixTo_346_dout;
  wire       [15:0]   fixTo_347_dout;
  wire       [15:0]   fixTo_348_dout;
  wire       [15:0]   fixTo_349_dout;
  wire       [15:0]   fixTo_350_dout;
  wire       [15:0]   fixTo_351_dout;
  wire       [15:0]   fixTo_352_dout;
  wire       [15:0]   fixTo_353_dout;
  wire       [15:0]   fixTo_354_dout;
  wire       [15:0]   fixTo_355_dout;
  wire       [15:0]   fixTo_356_dout;
  wire       [15:0]   fixTo_357_dout;
  wire       [15:0]   fixTo_358_dout;
  wire       [15:0]   fixTo_359_dout;
  wire       [15:0]   fixTo_360_dout;
  wire       [15:0]   fixTo_361_dout;
  wire       [15:0]   fixTo_362_dout;
  wire       [15:0]   fixTo_363_dout;
  wire       [15:0]   fixTo_364_dout;
  wire       [15:0]   fixTo_365_dout;
  wire       [15:0]   fixTo_366_dout;
  wire       [15:0]   fixTo_367_dout;
  wire       [15:0]   fixTo_368_dout;
  wire       [15:0]   fixTo_369_dout;
  wire       [15:0]   fixTo_370_dout;
  wire       [15:0]   fixTo_371_dout;
  wire       [15:0]   fixTo_372_dout;
  wire       [15:0]   fixTo_373_dout;
  wire       [15:0]   fixTo_374_dout;
  wire       [15:0]   fixTo_375_dout;
  wire       [15:0]   fixTo_376_dout;
  wire       [15:0]   fixTo_377_dout;
  wire       [15:0]   fixTo_378_dout;
  wire       [15:0]   fixTo_379_dout;
  wire       [15:0]   fixTo_380_dout;
  wire       [15:0]   fixTo_381_dout;
  wire       [15:0]   fixTo_382_dout;
  wire       [15:0]   fixTo_383_dout;
  wire       [15:0]   fixTo_384_dout;
  wire       [15:0]   fixTo_385_dout;
  wire       [15:0]   fixTo_386_dout;
  wire       [15:0]   fixTo_387_dout;
  wire       [15:0]   fixTo_388_dout;
  wire       [15:0]   fixTo_389_dout;
  wire       [15:0]   fixTo_390_dout;
  wire       [15:0]   fixTo_391_dout;
  wire       [15:0]   fixTo_392_dout;
  wire       [15:0]   fixTo_393_dout;
  wire       [15:0]   fixTo_394_dout;
  wire       [15:0]   fixTo_395_dout;
  wire       [15:0]   fixTo_396_dout;
  wire       [15:0]   fixTo_397_dout;
  wire       [15:0]   fixTo_398_dout;
  wire       [15:0]   fixTo_399_dout;
  wire       [15:0]   fixTo_400_dout;
  wire       [15:0]   fixTo_401_dout;
  wire       [15:0]   fixTo_402_dout;
  wire       [15:0]   fixTo_403_dout;
  wire       [15:0]   fixTo_404_dout;
  wire       [15:0]   fixTo_405_dout;
  wire       [15:0]   fixTo_406_dout;
  wire       [15:0]   fixTo_407_dout;
  wire       [15:0]   fixTo_408_dout;
  wire       [15:0]   fixTo_409_dout;
  wire       [15:0]   fixTo_410_dout;
  wire       [15:0]   fixTo_411_dout;
  wire       [15:0]   fixTo_412_dout;
  wire       [15:0]   fixTo_413_dout;
  wire       [15:0]   fixTo_414_dout;
  wire       [15:0]   fixTo_415_dout;
  wire       [15:0]   fixTo_416_dout;
  wire       [15:0]   fixTo_417_dout;
  wire       [15:0]   fixTo_418_dout;
  wire       [15:0]   fixTo_419_dout;
  wire       [15:0]   fixTo_420_dout;
  wire       [15:0]   fixTo_421_dout;
  wire       [15:0]   fixTo_422_dout;
  wire       [15:0]   fixTo_423_dout;
  wire       [15:0]   fixTo_424_dout;
  wire       [15:0]   fixTo_425_dout;
  wire       [15:0]   fixTo_426_dout;
  wire       [15:0]   fixTo_427_dout;
  wire       [15:0]   fixTo_428_dout;
  wire       [15:0]   fixTo_429_dout;
  wire       [15:0]   fixTo_430_dout;
  wire       [15:0]   fixTo_431_dout;
  wire       [15:0]   fixTo_432_dout;
  wire       [15:0]   fixTo_433_dout;
  wire       [15:0]   fixTo_434_dout;
  wire       [15:0]   fixTo_435_dout;
  wire       [15:0]   fixTo_436_dout;
  wire       [15:0]   fixTo_437_dout;
  wire       [15:0]   fixTo_438_dout;
  wire       [15:0]   fixTo_439_dout;
  wire       [15:0]   fixTo_440_dout;
  wire       [15:0]   fixTo_441_dout;
  wire       [15:0]   fixTo_442_dout;
  wire       [15:0]   fixTo_443_dout;
  wire       [15:0]   fixTo_444_dout;
  wire       [15:0]   fixTo_445_dout;
  wire       [15:0]   fixTo_446_dout;
  wire       [15:0]   fixTo_447_dout;
  wire       [15:0]   fixTo_448_dout;
  wire       [15:0]   fixTo_449_dout;
  wire       [15:0]   fixTo_450_dout;
  wire       [15:0]   fixTo_451_dout;
  wire       [15:0]   fixTo_452_dout;
  wire       [15:0]   fixTo_453_dout;
  wire       [15:0]   fixTo_454_dout;
  wire       [15:0]   fixTo_455_dout;
  wire       [15:0]   fixTo_456_dout;
  wire       [15:0]   fixTo_457_dout;
  wire       [15:0]   fixTo_458_dout;
  wire       [15:0]   fixTo_459_dout;
  wire       [15:0]   fixTo_460_dout;
  wire       [15:0]   fixTo_461_dout;
  wire       [15:0]   fixTo_462_dout;
  wire       [15:0]   fixTo_463_dout;
  wire       [15:0]   fixTo_464_dout;
  wire       [15:0]   fixTo_465_dout;
  wire       [15:0]   fixTo_466_dout;
  wire       [15:0]   fixTo_467_dout;
  wire       [15:0]   fixTo_468_dout;
  wire       [15:0]   fixTo_469_dout;
  wire       [15:0]   fixTo_470_dout;
  wire       [15:0]   fixTo_471_dout;
  wire       [15:0]   fixTo_472_dout;
  wire       [15:0]   fixTo_473_dout;
  wire       [15:0]   fixTo_474_dout;
  wire       [15:0]   fixTo_475_dout;
  wire       [15:0]   fixTo_476_dout;
  wire       [15:0]   fixTo_477_dout;
  wire       [15:0]   fixTo_478_dout;
  wire       [15:0]   fixTo_479_dout;
  wire       [15:0]   fixTo_480_dout;
  wire       [15:0]   fixTo_481_dout;
  wire       [15:0]   fixTo_482_dout;
  wire       [15:0]   fixTo_483_dout;
  wire       [15:0]   fixTo_484_dout;
  wire       [15:0]   fixTo_485_dout;
  wire       [15:0]   fixTo_486_dout;
  wire       [15:0]   fixTo_487_dout;
  wire       [15:0]   fixTo_488_dout;
  wire       [15:0]   fixTo_489_dout;
  wire       [15:0]   fixTo_490_dout;
  wire       [15:0]   fixTo_491_dout;
  wire       [15:0]   fixTo_492_dout;
  wire       [15:0]   fixTo_493_dout;
  wire       [15:0]   fixTo_494_dout;
  wire       [15:0]   fixTo_495_dout;
  wire       [15:0]   fixTo_496_dout;
  wire       [15:0]   fixTo_497_dout;
  wire       [15:0]   fixTo_498_dout;
  wire       [15:0]   fixTo_499_dout;
  wire       [15:0]   fixTo_500_dout;
  wire       [15:0]   fixTo_501_dout;
  wire       [15:0]   fixTo_502_dout;
  wire       [15:0]   fixTo_503_dout;
  wire       [15:0]   fixTo_504_dout;
  wire       [15:0]   fixTo_505_dout;
  wire       [15:0]   fixTo_506_dout;
  wire       [15:0]   fixTo_507_dout;
  wire       [15:0]   fixTo_508_dout;
  wire       [15:0]   fixTo_509_dout;
  wire       [15:0]   fixTo_510_dout;
  wire       [15:0]   fixTo_511_dout;
  wire       [15:0]   fixTo_512_dout;
  wire       [15:0]   fixTo_513_dout;
  wire       [15:0]   fixTo_514_dout;
  wire       [15:0]   fixTo_515_dout;
  wire       [15:0]   fixTo_516_dout;
  wire       [15:0]   fixTo_517_dout;
  wire       [15:0]   fixTo_518_dout;
  wire       [15:0]   fixTo_519_dout;
  wire       [15:0]   fixTo_520_dout;
  wire       [15:0]   fixTo_521_dout;
  wire       [15:0]   fixTo_522_dout;
  wire       [15:0]   fixTo_523_dout;
  wire       [15:0]   fixTo_524_dout;
  wire       [15:0]   fixTo_525_dout;
  wire       [15:0]   fixTo_526_dout;
  wire       [15:0]   fixTo_527_dout;
  wire       [15:0]   fixTo_528_dout;
  wire       [15:0]   fixTo_529_dout;
  wire       [15:0]   fixTo_530_dout;
  wire       [15:0]   fixTo_531_dout;
  wire       [15:0]   fixTo_532_dout;
  wire       [15:0]   fixTo_533_dout;
  wire       [15:0]   fixTo_534_dout;
  wire       [15:0]   fixTo_535_dout;
  wire       [15:0]   fixTo_536_dout;
  wire       [15:0]   fixTo_537_dout;
  wire       [15:0]   fixTo_538_dout;
  wire       [15:0]   fixTo_539_dout;
  wire       [15:0]   fixTo_540_dout;
  wire       [15:0]   fixTo_541_dout;
  wire       [15:0]   fixTo_542_dout;
  wire       [15:0]   fixTo_543_dout;
  wire       [15:0]   fixTo_544_dout;
  wire       [15:0]   fixTo_545_dout;
  wire       [15:0]   fixTo_546_dout;
  wire       [15:0]   fixTo_547_dout;
  wire       [15:0]   fixTo_548_dout;
  wire       [15:0]   fixTo_549_dout;
  wire       [15:0]   fixTo_550_dout;
  wire       [15:0]   fixTo_551_dout;
  wire       [15:0]   fixTo_552_dout;
  wire       [15:0]   fixTo_553_dout;
  wire       [15:0]   fixTo_554_dout;
  wire       [15:0]   fixTo_555_dout;
  wire       [15:0]   fixTo_556_dout;
  wire       [15:0]   fixTo_557_dout;
  wire       [15:0]   fixTo_558_dout;
  wire       [15:0]   fixTo_559_dout;
  wire       [15:0]   fixTo_560_dout;
  wire       [15:0]   fixTo_561_dout;
  wire       [15:0]   fixTo_562_dout;
  wire       [15:0]   fixTo_563_dout;
  wire       [15:0]   fixTo_564_dout;
  wire       [15:0]   fixTo_565_dout;
  wire       [15:0]   fixTo_566_dout;
  wire       [15:0]   fixTo_567_dout;
  wire       [15:0]   fixTo_568_dout;
  wire       [15:0]   fixTo_569_dout;
  wire       [15:0]   fixTo_570_dout;
  wire       [15:0]   fixTo_571_dout;
  wire       [15:0]   fixTo_572_dout;
  wire       [15:0]   fixTo_573_dout;
  wire       [15:0]   fixTo_574_dout;
  wire       [15:0]   fixTo_575_dout;
  wire       [15:0]   fixTo_576_dout;
  wire       [15:0]   fixTo_577_dout;
  wire       [15:0]   fixTo_578_dout;
  wire       [15:0]   fixTo_579_dout;
  wire       [15:0]   fixTo_580_dout;
  wire       [15:0]   fixTo_581_dout;
  wire       [15:0]   fixTo_582_dout;
  wire       [15:0]   fixTo_583_dout;
  wire       [15:0]   fixTo_584_dout;
  wire       [15:0]   fixTo_585_dout;
  wire       [15:0]   fixTo_586_dout;
  wire       [15:0]   fixTo_587_dout;
  wire       [15:0]   fixTo_588_dout;
  wire       [15:0]   fixTo_589_dout;
  wire       [15:0]   fixTo_590_dout;
  wire       [15:0]   fixTo_591_dout;
  wire       [15:0]   fixTo_592_dout;
  wire       [15:0]   fixTo_593_dout;
  wire       [15:0]   fixTo_594_dout;
  wire       [15:0]   fixTo_595_dout;
  wire       [15:0]   fixTo_596_dout;
  wire       [15:0]   fixTo_597_dout;
  wire       [15:0]   fixTo_598_dout;
  wire       [15:0]   fixTo_599_dout;
  wire       [15:0]   fixTo_600_dout;
  wire       [15:0]   fixTo_601_dout;
  wire       [15:0]   fixTo_602_dout;
  wire       [15:0]   fixTo_603_dout;
  wire       [15:0]   fixTo_604_dout;
  wire       [15:0]   fixTo_605_dout;
  wire       [15:0]   fixTo_606_dout;
  wire       [15:0]   fixTo_607_dout;
  wire       [15:0]   fixTo_608_dout;
  wire       [15:0]   fixTo_609_dout;
  wire       [15:0]   fixTo_610_dout;
  wire       [15:0]   fixTo_611_dout;
  wire       [15:0]   fixTo_612_dout;
  wire       [15:0]   fixTo_613_dout;
  wire       [15:0]   fixTo_614_dout;
  wire       [15:0]   fixTo_615_dout;
  wire       [15:0]   fixTo_616_dout;
  wire       [15:0]   fixTo_617_dout;
  wire       [15:0]   fixTo_618_dout;
  wire       [15:0]   fixTo_619_dout;
  wire       [15:0]   fixTo_620_dout;
  wire       [15:0]   fixTo_621_dout;
  wire       [15:0]   fixTo_622_dout;
  wire       [15:0]   fixTo_623_dout;
  wire       [15:0]   fixTo_624_dout;
  wire       [15:0]   fixTo_625_dout;
  wire       [15:0]   fixTo_626_dout;
  wire       [15:0]   fixTo_627_dout;
  wire       [15:0]   fixTo_628_dout;
  wire       [15:0]   fixTo_629_dout;
  wire       [15:0]   fixTo_630_dout;
  wire       [15:0]   fixTo_631_dout;
  wire       [15:0]   fixTo_632_dout;
  wire       [15:0]   fixTo_633_dout;
  wire       [15:0]   fixTo_634_dout;
  wire       [15:0]   fixTo_635_dout;
  wire       [15:0]   fixTo_636_dout;
  wire       [15:0]   fixTo_637_dout;
  wire       [15:0]   fixTo_638_dout;
  wire       [15:0]   fixTo_639_dout;
  wire       [15:0]   fixTo_640_dout;
  wire       [15:0]   fixTo_641_dout;
  wire       [15:0]   fixTo_642_dout;
  wire       [15:0]   fixTo_643_dout;
  wire       [15:0]   fixTo_644_dout;
  wire       [15:0]   fixTo_645_dout;
  wire       [15:0]   fixTo_646_dout;
  wire       [15:0]   fixTo_647_dout;
  wire       [15:0]   fixTo_648_dout;
  wire       [15:0]   fixTo_649_dout;
  wire       [15:0]   fixTo_650_dout;
  wire       [15:0]   fixTo_651_dout;
  wire       [15:0]   fixTo_652_dout;
  wire       [15:0]   fixTo_653_dout;
  wire       [15:0]   fixTo_654_dout;
  wire       [15:0]   fixTo_655_dout;
  wire       [15:0]   fixTo_656_dout;
  wire       [15:0]   fixTo_657_dout;
  wire       [15:0]   fixTo_658_dout;
  wire       [15:0]   fixTo_659_dout;
  wire       [15:0]   fixTo_660_dout;
  wire       [15:0]   fixTo_661_dout;
  wire       [15:0]   fixTo_662_dout;
  wire       [15:0]   fixTo_663_dout;
  wire       [15:0]   fixTo_664_dout;
  wire       [15:0]   fixTo_665_dout;
  wire       [15:0]   fixTo_666_dout;
  wire       [15:0]   fixTo_667_dout;
  wire       [15:0]   fixTo_668_dout;
  wire       [15:0]   fixTo_669_dout;
  wire       [15:0]   fixTo_670_dout;
  wire       [15:0]   fixTo_671_dout;
  wire       [15:0]   fixTo_672_dout;
  wire       [15:0]   fixTo_673_dout;
  wire       [15:0]   fixTo_674_dout;
  wire       [15:0]   fixTo_675_dout;
  wire       [15:0]   fixTo_676_dout;
  wire       [15:0]   fixTo_677_dout;
  wire       [15:0]   fixTo_678_dout;
  wire       [15:0]   fixTo_679_dout;
  wire       [15:0]   fixTo_680_dout;
  wire       [15:0]   fixTo_681_dout;
  wire       [15:0]   fixTo_682_dout;
  wire       [15:0]   fixTo_683_dout;
  wire       [15:0]   fixTo_684_dout;
  wire       [15:0]   fixTo_685_dout;
  wire       [15:0]   fixTo_686_dout;
  wire       [15:0]   fixTo_687_dout;
  wire       [15:0]   fixTo_688_dout;
  wire       [15:0]   fixTo_689_dout;
  wire       [15:0]   fixTo_690_dout;
  wire       [15:0]   fixTo_691_dout;
  wire       [15:0]   fixTo_692_dout;
  wire       [15:0]   fixTo_693_dout;
  wire       [15:0]   fixTo_694_dout;
  wire       [15:0]   fixTo_695_dout;
  wire       [15:0]   fixTo_696_dout;
  wire       [15:0]   fixTo_697_dout;
  wire       [15:0]   fixTo_698_dout;
  wire       [15:0]   fixTo_699_dout;
  wire       [15:0]   fixTo_700_dout;
  wire       [15:0]   fixTo_701_dout;
  wire       [15:0]   fixTo_702_dout;
  wire       [15:0]   fixTo_703_dout;
  wire       [15:0]   fixTo_704_dout;
  wire       [15:0]   fixTo_705_dout;
  wire       [15:0]   fixTo_706_dout;
  wire       [15:0]   fixTo_707_dout;
  wire       [15:0]   fixTo_708_dout;
  wire       [15:0]   fixTo_709_dout;
  wire       [15:0]   fixTo_710_dout;
  wire       [15:0]   fixTo_711_dout;
  wire       [15:0]   fixTo_712_dout;
  wire       [15:0]   fixTo_713_dout;
  wire       [15:0]   fixTo_714_dout;
  wire       [15:0]   fixTo_715_dout;
  wire       [15:0]   fixTo_716_dout;
  wire       [15:0]   fixTo_717_dout;
  wire       [15:0]   fixTo_718_dout;
  wire       [15:0]   fixTo_719_dout;
  wire       [15:0]   fixTo_720_dout;
  wire       [15:0]   fixTo_721_dout;
  wire       [15:0]   fixTo_722_dout;
  wire       [15:0]   fixTo_723_dout;
  wire       [15:0]   fixTo_724_dout;
  wire       [15:0]   fixTo_725_dout;
  wire       [15:0]   fixTo_726_dout;
  wire       [15:0]   fixTo_727_dout;
  wire       [15:0]   fixTo_728_dout;
  wire       [15:0]   fixTo_729_dout;
  wire       [15:0]   fixTo_730_dout;
  wire       [15:0]   fixTo_731_dout;
  wire       [15:0]   fixTo_732_dout;
  wire       [15:0]   fixTo_733_dout;
  wire       [15:0]   fixTo_734_dout;
  wire       [15:0]   fixTo_735_dout;
  wire       [15:0]   fixTo_736_dout;
  wire       [15:0]   fixTo_737_dout;
  wire       [15:0]   fixTo_738_dout;
  wire       [15:0]   fixTo_739_dout;
  wire       [15:0]   fixTo_740_dout;
  wire       [15:0]   fixTo_741_dout;
  wire       [15:0]   fixTo_742_dout;
  wire       [15:0]   fixTo_743_dout;
  wire       [15:0]   fixTo_744_dout;
  wire       [15:0]   fixTo_745_dout;
  wire       [15:0]   fixTo_746_dout;
  wire       [15:0]   fixTo_747_dout;
  wire       [15:0]   fixTo_748_dout;
  wire       [15:0]   fixTo_749_dout;
  wire       [15:0]   fixTo_750_dout;
  wire       [15:0]   fixTo_751_dout;
  wire       [15:0]   fixTo_752_dout;
  wire       [15:0]   fixTo_753_dout;
  wire       [15:0]   fixTo_754_dout;
  wire       [15:0]   fixTo_755_dout;
  wire       [15:0]   fixTo_756_dout;
  wire       [15:0]   fixTo_757_dout;
  wire       [15:0]   fixTo_758_dout;
  wire       [15:0]   fixTo_759_dout;
  wire       [15:0]   fixTo_760_dout;
  wire       [15:0]   fixTo_761_dout;
  wire       [15:0]   fixTo_762_dout;
  wire       [15:0]   fixTo_763_dout;
  wire       [15:0]   fixTo_764_dout;
  wire       [15:0]   fixTo_765_dout;
  wire       [15:0]   fixTo_766_dout;
  wire       [15:0]   fixTo_767_dout;
  wire       [15:0]   fixTo_768_dout;
  wire       [15:0]   fixTo_769_dout;
  wire       [15:0]   fixTo_770_dout;
  wire       [15:0]   fixTo_771_dout;
  wire       [15:0]   fixTo_772_dout;
  wire       [15:0]   fixTo_773_dout;
  wire       [15:0]   fixTo_774_dout;
  wire       [15:0]   fixTo_775_dout;
  wire       [15:0]   fixTo_776_dout;
  wire       [15:0]   fixTo_777_dout;
  wire       [15:0]   fixTo_778_dout;
  wire       [15:0]   fixTo_779_dout;
  wire       [15:0]   fixTo_780_dout;
  wire       [15:0]   fixTo_781_dout;
  wire       [15:0]   fixTo_782_dout;
  wire       [15:0]   fixTo_783_dout;
  wire       [15:0]   fixTo_784_dout;
  wire       [15:0]   fixTo_785_dout;
  wire       [15:0]   fixTo_786_dout;
  wire       [15:0]   fixTo_787_dout;
  wire       [15:0]   fixTo_788_dout;
  wire       [15:0]   fixTo_789_dout;
  wire       [15:0]   fixTo_790_dout;
  wire       [15:0]   fixTo_791_dout;
  wire       [15:0]   fixTo_792_dout;
  wire       [15:0]   fixTo_793_dout;
  wire       [15:0]   fixTo_794_dout;
  wire       [15:0]   fixTo_795_dout;
  wire       [15:0]   fixTo_796_dout;
  wire       [15:0]   fixTo_797_dout;
  wire       [15:0]   fixTo_798_dout;
  wire       [15:0]   fixTo_799_dout;
  wire       [15:0]   fixTo_800_dout;
  wire       [15:0]   fixTo_801_dout;
  wire       [15:0]   fixTo_802_dout;
  wire       [15:0]   fixTo_803_dout;
  wire       [15:0]   fixTo_804_dout;
  wire       [15:0]   fixTo_805_dout;
  wire       [15:0]   fixTo_806_dout;
  wire       [15:0]   fixTo_807_dout;
  wire       [15:0]   fixTo_808_dout;
  wire       [15:0]   fixTo_809_dout;
  wire       [15:0]   fixTo_810_dout;
  wire       [15:0]   fixTo_811_dout;
  wire       [15:0]   fixTo_812_dout;
  wire       [15:0]   fixTo_813_dout;
  wire       [15:0]   fixTo_814_dout;
  wire       [15:0]   fixTo_815_dout;
  wire       [15:0]   fixTo_816_dout;
  wire       [15:0]   fixTo_817_dout;
  wire       [15:0]   fixTo_818_dout;
  wire       [15:0]   fixTo_819_dout;
  wire       [15:0]   fixTo_820_dout;
  wire       [15:0]   fixTo_821_dout;
  wire       [15:0]   fixTo_822_dout;
  wire       [15:0]   fixTo_823_dout;
  wire       [15:0]   fixTo_824_dout;
  wire       [15:0]   fixTo_825_dout;
  wire       [15:0]   fixTo_826_dout;
  wire       [15:0]   fixTo_827_dout;
  wire       [15:0]   fixTo_828_dout;
  wire       [15:0]   fixTo_829_dout;
  wire       [15:0]   fixTo_830_dout;
  wire       [15:0]   fixTo_831_dout;
  wire       [15:0]   fixTo_832_dout;
  wire       [15:0]   fixTo_833_dout;
  wire       [15:0]   fixTo_834_dout;
  wire       [15:0]   fixTo_835_dout;
  wire       [15:0]   fixTo_836_dout;
  wire       [15:0]   fixTo_837_dout;
  wire       [15:0]   fixTo_838_dout;
  wire       [15:0]   fixTo_839_dout;
  wire       [15:0]   fixTo_840_dout;
  wire       [15:0]   fixTo_841_dout;
  wire       [15:0]   fixTo_842_dout;
  wire       [15:0]   fixTo_843_dout;
  wire       [15:0]   fixTo_844_dout;
  wire       [15:0]   fixTo_845_dout;
  wire       [15:0]   fixTo_846_dout;
  wire       [15:0]   fixTo_847_dout;
  wire       [15:0]   fixTo_848_dout;
  wire       [15:0]   fixTo_849_dout;
  wire       [15:0]   fixTo_850_dout;
  wire       [15:0]   fixTo_851_dout;
  wire       [15:0]   fixTo_852_dout;
  wire       [15:0]   fixTo_853_dout;
  wire       [15:0]   fixTo_854_dout;
  wire       [15:0]   fixTo_855_dout;
  wire       [15:0]   fixTo_856_dout;
  wire       [15:0]   fixTo_857_dout;
  wire       [15:0]   fixTo_858_dout;
  wire       [15:0]   fixTo_859_dout;
  wire       [15:0]   fixTo_860_dout;
  wire       [15:0]   fixTo_861_dout;
  wire       [15:0]   fixTo_862_dout;
  wire       [15:0]   fixTo_863_dout;
  wire       [15:0]   fixTo_864_dout;
  wire       [15:0]   fixTo_865_dout;
  wire       [15:0]   fixTo_866_dout;
  wire       [15:0]   fixTo_867_dout;
  wire       [15:0]   fixTo_868_dout;
  wire       [15:0]   fixTo_869_dout;
  wire       [15:0]   fixTo_870_dout;
  wire       [15:0]   fixTo_871_dout;
  wire       [15:0]   fixTo_872_dout;
  wire       [15:0]   fixTo_873_dout;
  wire       [15:0]   fixTo_874_dout;
  wire       [15:0]   fixTo_875_dout;
  wire       [15:0]   fixTo_876_dout;
  wire       [15:0]   fixTo_877_dout;
  wire       [15:0]   fixTo_878_dout;
  wire       [15:0]   fixTo_879_dout;
  wire       [15:0]   fixTo_880_dout;
  wire       [15:0]   fixTo_881_dout;
  wire       [15:0]   fixTo_882_dout;
  wire       [15:0]   fixTo_883_dout;
  wire       [15:0]   fixTo_884_dout;
  wire       [15:0]   fixTo_885_dout;
  wire       [15:0]   fixTo_886_dout;
  wire       [15:0]   fixTo_887_dout;
  wire       [15:0]   fixTo_888_dout;
  wire       [15:0]   fixTo_889_dout;
  wire       [15:0]   fixTo_890_dout;
  wire       [15:0]   fixTo_891_dout;
  wire       [15:0]   fixTo_892_dout;
  wire       [15:0]   fixTo_893_dout;
  wire       [15:0]   fixTo_894_dout;
  wire       [15:0]   fixTo_895_dout;
  wire       [15:0]   fixTo_896_dout;
  wire       [15:0]   fixTo_897_dout;
  wire       [15:0]   fixTo_898_dout;
  wire       [15:0]   fixTo_899_dout;
  wire       [15:0]   fixTo_900_dout;
  wire       [15:0]   fixTo_901_dout;
  wire       [15:0]   fixTo_902_dout;
  wire       [15:0]   fixTo_903_dout;
  wire       [15:0]   fixTo_904_dout;
  wire       [15:0]   fixTo_905_dout;
  wire       [15:0]   fixTo_906_dout;
  wire       [15:0]   fixTo_907_dout;
  wire       [15:0]   fixTo_908_dout;
  wire       [15:0]   fixTo_909_dout;
  wire       [15:0]   fixTo_910_dout;
  wire       [15:0]   fixTo_911_dout;
  wire       [15:0]   fixTo_912_dout;
  wire       [15:0]   fixTo_913_dout;
  wire       [15:0]   fixTo_914_dout;
  wire       [15:0]   fixTo_915_dout;
  wire       [15:0]   fixTo_916_dout;
  wire       [15:0]   fixTo_917_dout;
  wire       [15:0]   fixTo_918_dout;
  wire       [15:0]   fixTo_919_dout;
  wire       [15:0]   fixTo_920_dout;
  wire       [15:0]   fixTo_921_dout;
  wire       [15:0]   fixTo_922_dout;
  wire       [15:0]   fixTo_923_dout;
  wire       [15:0]   fixTo_924_dout;
  wire       [15:0]   fixTo_925_dout;
  wire       [15:0]   fixTo_926_dout;
  wire       [15:0]   fixTo_927_dout;
  wire       [15:0]   fixTo_928_dout;
  wire       [15:0]   fixTo_929_dout;
  wire       [15:0]   fixTo_930_dout;
  wire       [15:0]   fixTo_931_dout;
  wire       [15:0]   fixTo_932_dout;
  wire       [15:0]   fixTo_933_dout;
  wire       [15:0]   fixTo_934_dout;
  wire       [15:0]   fixTo_935_dout;
  wire       [15:0]   fixTo_936_dout;
  wire       [15:0]   fixTo_937_dout;
  wire       [15:0]   fixTo_938_dout;
  wire       [15:0]   fixTo_939_dout;
  wire       [15:0]   fixTo_940_dout;
  wire       [15:0]   fixTo_941_dout;
  wire       [15:0]   fixTo_942_dout;
  wire       [15:0]   fixTo_943_dout;
  wire       [15:0]   fixTo_944_dout;
  wire       [15:0]   fixTo_945_dout;
  wire       [15:0]   fixTo_946_dout;
  wire       [15:0]   fixTo_947_dout;
  wire       [15:0]   fixTo_948_dout;
  wire       [15:0]   fixTo_949_dout;
  wire       [15:0]   fixTo_950_dout;
  wire       [15:0]   fixTo_951_dout;
  wire       [15:0]   fixTo_952_dout;
  wire       [15:0]   fixTo_953_dout;
  wire       [15:0]   fixTo_954_dout;
  wire       [15:0]   fixTo_955_dout;
  wire       [15:0]   fixTo_956_dout;
  wire       [15:0]   fixTo_957_dout;
  wire       [15:0]   fixTo_958_dout;
  wire       [15:0]   fixTo_959_dout;
  wire       [15:0]   fixTo_960_dout;
  wire       [15:0]   fixTo_961_dout;
  wire       [15:0]   fixTo_962_dout;
  wire       [15:0]   fixTo_963_dout;
  wire       [15:0]   fixTo_964_dout;
  wire       [15:0]   fixTo_965_dout;
  wire       [15:0]   fixTo_966_dout;
  wire       [15:0]   fixTo_967_dout;
  wire       [15:0]   fixTo_968_dout;
  wire       [15:0]   fixTo_969_dout;
  wire       [15:0]   fixTo_970_dout;
  wire       [15:0]   fixTo_971_dout;
  wire       [15:0]   fixTo_972_dout;
  wire       [15:0]   fixTo_973_dout;
  wire       [15:0]   fixTo_974_dout;
  wire       [15:0]   fixTo_975_dout;
  wire       [15:0]   fixTo_976_dout;
  wire       [15:0]   fixTo_977_dout;
  wire       [15:0]   fixTo_978_dout;
  wire       [15:0]   fixTo_979_dout;
  wire       [15:0]   fixTo_980_dout;
  wire       [15:0]   fixTo_981_dout;
  wire       [15:0]   fixTo_982_dout;
  wire       [15:0]   fixTo_983_dout;
  wire       [15:0]   fixTo_984_dout;
  wire       [15:0]   fixTo_985_dout;
  wire       [15:0]   fixTo_986_dout;
  wire       [15:0]   fixTo_987_dout;
  wire       [15:0]   fixTo_988_dout;
  wire       [15:0]   fixTo_989_dout;
  wire       [15:0]   fixTo_990_dout;
  wire       [15:0]   fixTo_991_dout;
  wire       [15:0]   fixTo_992_dout;
  wire       [15:0]   fixTo_993_dout;
  wire       [15:0]   fixTo_994_dout;
  wire       [15:0]   fixTo_995_dout;
  wire       [15:0]   fixTo_996_dout;
  wire       [15:0]   fixTo_997_dout;
  wire       [15:0]   fixTo_998_dout;
  wire       [15:0]   fixTo_999_dout;
  wire       [15:0]   fixTo_1000_dout;
  wire       [15:0]   fixTo_1001_dout;
  wire       [15:0]   fixTo_1002_dout;
  wire       [15:0]   fixTo_1003_dout;
  wire       [15:0]   fixTo_1004_dout;
  wire       [15:0]   fixTo_1005_dout;
  wire       [15:0]   fixTo_1006_dout;
  wire       [15:0]   fixTo_1007_dout;
  wire       [15:0]   fixTo_1008_dout;
  wire       [15:0]   fixTo_1009_dout;
  wire       [15:0]   fixTo_1010_dout;
  wire       [15:0]   fixTo_1011_dout;
  wire       [15:0]   fixTo_1012_dout;
  wire       [15:0]   fixTo_1013_dout;
  wire       [15:0]   fixTo_1014_dout;
  wire       [15:0]   fixTo_1015_dout;
  wire       [15:0]   fixTo_1016_dout;
  wire       [15:0]   fixTo_1017_dout;
  wire       [15:0]   fixTo_1018_dout;
  wire       [15:0]   fixTo_1019_dout;
  wire       [15:0]   fixTo_1020_dout;
  wire       [15:0]   fixTo_1021_dout;
  wire       [15:0]   fixTo_1022_dout;
  wire       [15:0]   fixTo_1023_dout;
  wire       [15:0]   fixTo_1024_dout;
  wire       [15:0]   fixTo_1025_dout;
  wire       [15:0]   fixTo_1026_dout;
  wire       [15:0]   fixTo_1027_dout;
  wire       [15:0]   fixTo_1028_dout;
  wire       [15:0]   fixTo_1029_dout;
  wire       [15:0]   fixTo_1030_dout;
  wire       [15:0]   fixTo_1031_dout;
  wire       [15:0]   fixTo_1032_dout;
  wire       [15:0]   fixTo_1033_dout;
  wire       [15:0]   fixTo_1034_dout;
  wire       [15:0]   fixTo_1035_dout;
  wire       [15:0]   fixTo_1036_dout;
  wire       [15:0]   fixTo_1037_dout;
  wire       [15:0]   fixTo_1038_dout;
  wire       [15:0]   fixTo_1039_dout;
  wire       [15:0]   fixTo_1040_dout;
  wire       [15:0]   fixTo_1041_dout;
  wire       [15:0]   fixTo_1042_dout;
  wire       [15:0]   fixTo_1043_dout;
  wire       [15:0]   fixTo_1044_dout;
  wire       [15:0]   fixTo_1045_dout;
  wire       [15:0]   fixTo_1046_dout;
  wire       [15:0]   fixTo_1047_dout;
  wire       [15:0]   fixTo_1048_dout;
  wire       [15:0]   fixTo_1049_dout;
  wire       [15:0]   fixTo_1050_dout;
  wire       [15:0]   fixTo_1051_dout;
  wire       [15:0]   fixTo_1052_dout;
  wire       [15:0]   fixTo_1053_dout;
  wire       [15:0]   fixTo_1054_dout;
  wire       [15:0]   fixTo_1055_dout;
  wire       [15:0]   fixTo_1056_dout;
  wire       [15:0]   fixTo_1057_dout;
  wire       [15:0]   fixTo_1058_dout;
  wire       [15:0]   fixTo_1059_dout;
  wire       [15:0]   fixTo_1060_dout;
  wire       [15:0]   fixTo_1061_dout;
  wire       [15:0]   fixTo_1062_dout;
  wire       [15:0]   fixTo_1063_dout;
  wire       [15:0]   fixTo_1064_dout;
  wire       [15:0]   fixTo_1065_dout;
  wire       [15:0]   fixTo_1066_dout;
  wire       [15:0]   fixTo_1067_dout;
  wire       [15:0]   fixTo_1068_dout;
  wire       [15:0]   fixTo_1069_dout;
  wire       [15:0]   fixTo_1070_dout;
  wire       [15:0]   fixTo_1071_dout;
  wire       [15:0]   fixTo_1072_dout;
  wire       [15:0]   fixTo_1073_dout;
  wire       [15:0]   fixTo_1074_dout;
  wire       [15:0]   fixTo_1075_dout;
  wire       [15:0]   fixTo_1076_dout;
  wire       [15:0]   fixTo_1077_dout;
  wire       [15:0]   fixTo_1078_dout;
  wire       [15:0]   fixTo_1079_dout;
  wire       [15:0]   fixTo_1080_dout;
  wire       [15:0]   fixTo_1081_dout;
  wire       [15:0]   fixTo_1082_dout;
  wire       [15:0]   fixTo_1083_dout;
  wire       [15:0]   fixTo_1084_dout;
  wire       [15:0]   fixTo_1085_dout;
  wire       [15:0]   fixTo_1086_dout;
  wire       [15:0]   fixTo_1087_dout;
  wire       [15:0]   fixTo_1088_dout;
  wire       [15:0]   fixTo_1089_dout;
  wire       [15:0]   fixTo_1090_dout;
  wire       [15:0]   fixTo_1091_dout;
  wire       [15:0]   fixTo_1092_dout;
  wire       [15:0]   fixTo_1093_dout;
  wire       [15:0]   fixTo_1094_dout;
  wire       [15:0]   fixTo_1095_dout;
  wire       [15:0]   fixTo_1096_dout;
  wire       [15:0]   fixTo_1097_dout;
  wire       [15:0]   fixTo_1098_dout;
  wire       [15:0]   fixTo_1099_dout;
  wire       [15:0]   fixTo_1100_dout;
  wire       [15:0]   fixTo_1101_dout;
  wire       [15:0]   fixTo_1102_dout;
  wire       [15:0]   fixTo_1103_dout;
  wire       [15:0]   fixTo_1104_dout;
  wire       [15:0]   fixTo_1105_dout;
  wire       [15:0]   fixTo_1106_dout;
  wire       [15:0]   fixTo_1107_dout;
  wire       [15:0]   fixTo_1108_dout;
  wire       [15:0]   fixTo_1109_dout;
  wire       [15:0]   fixTo_1110_dout;
  wire       [15:0]   fixTo_1111_dout;
  wire       [15:0]   fixTo_1112_dout;
  wire       [15:0]   fixTo_1113_dout;
  wire       [15:0]   fixTo_1114_dout;
  wire       [15:0]   fixTo_1115_dout;
  wire       [15:0]   fixTo_1116_dout;
  wire       [15:0]   fixTo_1117_dout;
  wire       [15:0]   fixTo_1118_dout;
  wire       [15:0]   fixTo_1119_dout;
  wire       [15:0]   fixTo_1120_dout;
  wire       [15:0]   fixTo_1121_dout;
  wire       [15:0]   fixTo_1122_dout;
  wire       [15:0]   fixTo_1123_dout;
  wire       [15:0]   fixTo_1124_dout;
  wire       [15:0]   fixTo_1125_dout;
  wire       [15:0]   fixTo_1126_dout;
  wire       [15:0]   fixTo_1127_dout;
  wire       [15:0]   fixTo_1128_dout;
  wire       [15:0]   fixTo_1129_dout;
  wire       [15:0]   fixTo_1130_dout;
  wire       [15:0]   fixTo_1131_dout;
  wire       [15:0]   fixTo_1132_dout;
  wire       [15:0]   fixTo_1133_dout;
  wire       [15:0]   fixTo_1134_dout;
  wire       [15:0]   fixTo_1135_dout;
  wire       [15:0]   fixTo_1136_dout;
  wire       [15:0]   fixTo_1137_dout;
  wire       [15:0]   fixTo_1138_dout;
  wire       [15:0]   fixTo_1139_dout;
  wire       [15:0]   fixTo_1140_dout;
  wire       [15:0]   fixTo_1141_dout;
  wire       [15:0]   fixTo_1142_dout;
  wire       [15:0]   fixTo_1143_dout;
  wire       [15:0]   fixTo_1144_dout;
  wire       [15:0]   fixTo_1145_dout;
  wire       [15:0]   fixTo_1146_dout;
  wire       [15:0]   fixTo_1147_dout;
  wire       [15:0]   fixTo_1148_dout;
  wire       [15:0]   fixTo_1149_dout;
  wire       [15:0]   fixTo_1150_dout;
  wire       [15:0]   fixTo_1151_dout;
  wire       [15:0]   fixTo_1152_dout;
  wire       [15:0]   fixTo_1153_dout;
  wire       [15:0]   fixTo_1154_dout;
  wire       [15:0]   fixTo_1155_dout;
  wire       [15:0]   fixTo_1156_dout;
  wire       [15:0]   fixTo_1157_dout;
  wire       [15:0]   fixTo_1158_dout;
  wire       [15:0]   fixTo_1159_dout;
  wire       [15:0]   fixTo_1160_dout;
  wire       [15:0]   fixTo_1161_dout;
  wire       [15:0]   fixTo_1162_dout;
  wire       [15:0]   fixTo_1163_dout;
  wire       [15:0]   fixTo_1164_dout;
  wire       [15:0]   fixTo_1165_dout;
  wire       [15:0]   fixTo_1166_dout;
  wire       [15:0]   fixTo_1167_dout;
  wire       [15:0]   fixTo_1168_dout;
  wire       [15:0]   fixTo_1169_dout;
  wire       [15:0]   fixTo_1170_dout;
  wire       [15:0]   fixTo_1171_dout;
  wire       [15:0]   fixTo_1172_dout;
  wire       [15:0]   fixTo_1173_dout;
  wire       [15:0]   fixTo_1174_dout;
  wire       [15:0]   fixTo_1175_dout;
  wire       [15:0]   fixTo_1176_dout;
  wire       [15:0]   fixTo_1177_dout;
  wire       [15:0]   fixTo_1178_dout;
  wire       [15:0]   fixTo_1179_dout;
  wire       [15:0]   fixTo_1180_dout;
  wire       [15:0]   fixTo_1181_dout;
  wire       [15:0]   fixTo_1182_dout;
  wire       [15:0]   fixTo_1183_dout;
  wire       [15:0]   fixTo_1184_dout;
  wire       [15:0]   fixTo_1185_dout;
  wire       [15:0]   fixTo_1186_dout;
  wire       [15:0]   fixTo_1187_dout;
  wire       [15:0]   fixTo_1188_dout;
  wire       [15:0]   fixTo_1189_dout;
  wire       [15:0]   fixTo_1190_dout;
  wire       [15:0]   fixTo_1191_dout;
  wire       [15:0]   fixTo_1192_dout;
  wire       [15:0]   fixTo_1193_dout;
  wire       [15:0]   fixTo_1194_dout;
  wire       [15:0]   fixTo_1195_dout;
  wire       [15:0]   fixTo_1196_dout;
  wire       [15:0]   fixTo_1197_dout;
  wire       [15:0]   fixTo_1198_dout;
  wire       [15:0]   fixTo_1199_dout;
  wire       [15:0]   fixTo_1200_dout;
  wire       [15:0]   fixTo_1201_dout;
  wire       [15:0]   fixTo_1202_dout;
  wire       [15:0]   fixTo_1203_dout;
  wire       [15:0]   fixTo_1204_dout;
  wire       [15:0]   fixTo_1205_dout;
  wire       [15:0]   fixTo_1206_dout;
  wire       [15:0]   fixTo_1207_dout;
  wire       [15:0]   fixTo_1208_dout;
  wire       [15:0]   fixTo_1209_dout;
  wire       [15:0]   fixTo_1210_dout;
  wire       [15:0]   fixTo_1211_dout;
  wire       [15:0]   fixTo_1212_dout;
  wire       [15:0]   fixTo_1213_dout;
  wire       [15:0]   fixTo_1214_dout;
  wire       [15:0]   fixTo_1215_dout;
  wire       [15:0]   fixTo_1216_dout;
  wire       [15:0]   fixTo_1217_dout;
  wire       [15:0]   fixTo_1218_dout;
  wire       [15:0]   fixTo_1219_dout;
  wire       [15:0]   fixTo_1220_dout;
  wire       [15:0]   fixTo_1221_dout;
  wire       [15:0]   fixTo_1222_dout;
  wire       [15:0]   fixTo_1223_dout;
  wire       [15:0]   fixTo_1224_dout;
  wire       [15:0]   fixTo_1225_dout;
  wire       [15:0]   fixTo_1226_dout;
  wire       [15:0]   fixTo_1227_dout;
  wire       [15:0]   fixTo_1228_dout;
  wire       [15:0]   fixTo_1229_dout;
  wire       [15:0]   fixTo_1230_dout;
  wire       [15:0]   fixTo_1231_dout;
  wire       [15:0]   fixTo_1232_dout;
  wire       [15:0]   fixTo_1233_dout;
  wire       [15:0]   fixTo_1234_dout;
  wire       [15:0]   fixTo_1235_dout;
  wire       [15:0]   fixTo_1236_dout;
  wire       [15:0]   fixTo_1237_dout;
  wire       [15:0]   fixTo_1238_dout;
  wire       [15:0]   fixTo_1239_dout;
  wire       [15:0]   fixTo_1240_dout;
  wire       [15:0]   fixTo_1241_dout;
  wire       [15:0]   fixTo_1242_dout;
  wire       [15:0]   fixTo_1243_dout;
  wire       [15:0]   fixTo_1244_dout;
  wire       [15:0]   fixTo_1245_dout;
  wire       [15:0]   fixTo_1246_dout;
  wire       [15:0]   fixTo_1247_dout;
  wire       [15:0]   fixTo_1248_dout;
  wire       [15:0]   fixTo_1249_dout;
  wire       [15:0]   fixTo_1250_dout;
  wire       [15:0]   fixTo_1251_dout;
  wire       [15:0]   fixTo_1252_dout;
  wire       [15:0]   fixTo_1253_dout;
  wire       [15:0]   fixTo_1254_dout;
  wire       [15:0]   fixTo_1255_dout;
  wire       [15:0]   fixTo_1256_dout;
  wire       [15:0]   fixTo_1257_dout;
  wire       [15:0]   fixTo_1258_dout;
  wire       [15:0]   fixTo_1259_dout;
  wire       [15:0]   fixTo_1260_dout;
  wire       [15:0]   fixTo_1261_dout;
  wire       [15:0]   fixTo_1262_dout;
  wire       [15:0]   fixTo_1263_dout;
  wire       [15:0]   fixTo_1264_dout;
  wire       [15:0]   fixTo_1265_dout;
  wire       [15:0]   fixTo_1266_dout;
  wire       [15:0]   fixTo_1267_dout;
  wire       [15:0]   fixTo_1268_dout;
  wire       [15:0]   fixTo_1269_dout;
  wire       [15:0]   fixTo_1270_dout;
  wire       [15:0]   fixTo_1271_dout;
  wire       [15:0]   fixTo_1272_dout;
  wire       [15:0]   fixTo_1273_dout;
  wire       [15:0]   fixTo_1274_dout;
  wire       [15:0]   fixTo_1275_dout;
  wire       [15:0]   fixTo_1276_dout;
  wire       [15:0]   fixTo_1277_dout;
  wire       [15:0]   fixTo_1278_dout;
  wire       [15:0]   fixTo_1279_dout;
  wire       [15:0]   fixTo_1280_dout;
  wire       [15:0]   fixTo_1281_dout;
  wire       [15:0]   fixTo_1282_dout;
  wire       [15:0]   fixTo_1283_dout;
  wire       [15:0]   fixTo_1284_dout;
  wire       [15:0]   fixTo_1285_dout;
  wire       [15:0]   fixTo_1286_dout;
  wire       [15:0]   fixTo_1287_dout;
  wire       [15:0]   fixTo_1288_dout;
  wire       [15:0]   fixTo_1289_dout;
  wire       [15:0]   fixTo_1290_dout;
  wire       [15:0]   fixTo_1291_dout;
  wire       [15:0]   fixTo_1292_dout;
  wire       [15:0]   fixTo_1293_dout;
  wire       [15:0]   fixTo_1294_dout;
  wire       [15:0]   fixTo_1295_dout;
  wire       [15:0]   fixTo_1296_dout;
  wire       [15:0]   fixTo_1297_dout;
  wire       [15:0]   fixTo_1298_dout;
  wire       [15:0]   fixTo_1299_dout;
  wire       [15:0]   fixTo_1300_dout;
  wire       [15:0]   fixTo_1301_dout;
  wire       [15:0]   fixTo_1302_dout;
  wire       [15:0]   fixTo_1303_dout;
  wire       [15:0]   fixTo_1304_dout;
  wire       [15:0]   fixTo_1305_dout;
  wire       [15:0]   fixTo_1306_dout;
  wire       [15:0]   fixTo_1307_dout;
  wire       [15:0]   fixTo_1308_dout;
  wire       [15:0]   fixTo_1309_dout;
  wire       [15:0]   fixTo_1310_dout;
  wire       [15:0]   fixTo_1311_dout;
  wire       [15:0]   fixTo_1312_dout;
  wire       [15:0]   fixTo_1313_dout;
  wire       [15:0]   fixTo_1314_dout;
  wire       [15:0]   fixTo_1315_dout;
  wire       [15:0]   fixTo_1316_dout;
  wire       [15:0]   fixTo_1317_dout;
  wire       [15:0]   fixTo_1318_dout;
  wire       [15:0]   fixTo_1319_dout;
  wire       [15:0]   fixTo_1320_dout;
  wire       [15:0]   fixTo_1321_dout;
  wire       [15:0]   fixTo_1322_dout;
  wire       [15:0]   fixTo_1323_dout;
  wire       [15:0]   fixTo_1324_dout;
  wire       [15:0]   fixTo_1325_dout;
  wire       [15:0]   fixTo_1326_dout;
  wire       [15:0]   fixTo_1327_dout;
  wire       [15:0]   fixTo_1328_dout;
  wire       [15:0]   fixTo_1329_dout;
  wire       [15:0]   fixTo_1330_dout;
  wire       [15:0]   fixTo_1331_dout;
  wire       [15:0]   fixTo_1332_dout;
  wire       [15:0]   fixTo_1333_dout;
  wire       [15:0]   fixTo_1334_dout;
  wire       [15:0]   fixTo_1335_dout;
  wire       [15:0]   fixTo_1336_dout;
  wire       [15:0]   fixTo_1337_dout;
  wire       [15:0]   fixTo_1338_dout;
  wire       [15:0]   fixTo_1339_dout;
  wire       [15:0]   fixTo_1340_dout;
  wire       [15:0]   fixTo_1341_dout;
  wire       [15:0]   fixTo_1342_dout;
  wire       [15:0]   fixTo_1343_dout;
  wire       [15:0]   _zz_5383;
  wire       [15:0]   _zz_5384;
  wire       [15:0]   _zz_5385;
  wire       [15:0]   _zz_5386;
  wire       [15:0]   _zz_5387;
  wire       [15:0]   _zz_5388;
  wire       [15:0]   _zz_5389;
  wire       [15:0]   _zz_5390;
  wire       [15:0]   _zz_5391;
  wire       [15:0]   _zz_5392;
  wire       [15:0]   _zz_5393;
  wire       [15:0]   _zz_5394;
  wire       [15:0]   _zz_5395;
  wire       [15:0]   _zz_5396;
  wire       [15:0]   _zz_5397;
  wire       [15:0]   _zz_5398;
  wire       [15:0]   _zz_5399;
  wire       [15:0]   _zz_5400;
  wire       [15:0]   _zz_5401;
  wire       [15:0]   _zz_5402;
  wire       [15:0]   _zz_5403;
  wire       [15:0]   _zz_5404;
  wire       [15:0]   _zz_5405;
  wire       [15:0]   _zz_5406;
  wire       [15:0]   _zz_5407;
  wire       [15:0]   _zz_5408;
  wire       [15:0]   _zz_5409;
  wire       [15:0]   _zz_5410;
  wire       [15:0]   _zz_5411;
  wire       [15:0]   _zz_5412;
  wire       [15:0]   _zz_5413;
  wire       [15:0]   _zz_5414;
  wire       [15:0]   _zz_5415;
  wire       [15:0]   _zz_5416;
  wire       [15:0]   _zz_5417;
  wire       [15:0]   _zz_5418;
  wire       [15:0]   _zz_5419;
  wire       [15:0]   _zz_5420;
  wire       [15:0]   _zz_5421;
  wire       [15:0]   _zz_5422;
  wire       [15:0]   _zz_5423;
  wire       [15:0]   _zz_5424;
  wire       [15:0]   _zz_5425;
  wire       [15:0]   _zz_5426;
  wire       [15:0]   _zz_5427;
  wire       [15:0]   _zz_5428;
  wire       [15:0]   _zz_5429;
  wire       [15:0]   _zz_5430;
  wire       [15:0]   _zz_5431;
  wire       [15:0]   _zz_5432;
  wire       [15:0]   _zz_5433;
  wire       [15:0]   _zz_5434;
  wire       [15:0]   _zz_5435;
  wire       [15:0]   _zz_5436;
  wire       [15:0]   _zz_5437;
  wire       [15:0]   _zz_5438;
  wire       [15:0]   _zz_5439;
  wire       [15:0]   _zz_5440;
  wire       [15:0]   _zz_5441;
  wire       [15:0]   _zz_5442;
  wire       [15:0]   _zz_5443;
  wire       [15:0]   _zz_5444;
  wire       [15:0]   _zz_5445;
  wire       [15:0]   _zz_5446;
  wire       [15:0]   _zz_5447;
  wire       [15:0]   _zz_5448;
  wire       [15:0]   _zz_5449;
  wire       [15:0]   _zz_5450;
  wire       [15:0]   _zz_5451;
  wire       [15:0]   _zz_5452;
  wire       [15:0]   _zz_5453;
  wire       [15:0]   _zz_5454;
  wire       [15:0]   _zz_5455;
  wire       [15:0]   _zz_5456;
  wire       [15:0]   _zz_5457;
  wire       [15:0]   _zz_5458;
  wire       [15:0]   _zz_5459;
  wire       [15:0]   _zz_5460;
  wire       [15:0]   _zz_5461;
  wire       [15:0]   _zz_5462;
  wire       [15:0]   _zz_5463;
  wire       [15:0]   _zz_5464;
  wire       [15:0]   _zz_5465;
  wire       [15:0]   _zz_5466;
  wire       [15:0]   _zz_5467;
  wire       [15:0]   _zz_5468;
  wire       [15:0]   _zz_5469;
  wire       [15:0]   _zz_5470;
  wire       [15:0]   _zz_5471;
  wire       [15:0]   _zz_5472;
  wire       [15:0]   _zz_5473;
  wire       [15:0]   _zz_5474;
  wire       [15:0]   _zz_5475;
  wire       [15:0]   _zz_5476;
  wire       [15:0]   _zz_5477;
  wire       [15:0]   _zz_5478;
  wire       [15:0]   _zz_5479;
  wire       [15:0]   _zz_5480;
  wire       [15:0]   _zz_5481;
  wire       [15:0]   _zz_5482;
  wire       [15:0]   _zz_5483;
  wire       [15:0]   _zz_5484;
  wire       [15:0]   _zz_5485;
  wire       [15:0]   _zz_5486;
  wire       [15:0]   _zz_5487;
  wire       [15:0]   _zz_5488;
  wire       [15:0]   _zz_5489;
  wire       [15:0]   _zz_5490;
  wire       [15:0]   _zz_5491;
  wire       [15:0]   _zz_5492;
  wire       [15:0]   _zz_5493;
  wire       [15:0]   _zz_5494;
  wire       [15:0]   _zz_5495;
  wire       [15:0]   _zz_5496;
  wire       [15:0]   _zz_5497;
  wire       [15:0]   _zz_5498;
  wire       [15:0]   _zz_5499;
  wire       [15:0]   _zz_5500;
  wire       [15:0]   _zz_5501;
  wire       [15:0]   _zz_5502;
  wire       [15:0]   _zz_5503;
  wire       [15:0]   _zz_5504;
  wire       [15:0]   _zz_5505;
  wire       [15:0]   _zz_5506;
  wire       [15:0]   _zz_5507;
  wire       [15:0]   _zz_5508;
  wire       [15:0]   _zz_5509;
  wire       [15:0]   _zz_5510;
  wire       [15:0]   _zz_5511;
  wire       [15:0]   _zz_5512;
  wire       [15:0]   _zz_5513;
  wire       [15:0]   _zz_5514;
  wire       [15:0]   _zz_5515;
  wire       [15:0]   _zz_5516;
  wire       [15:0]   _zz_5517;
  wire       [15:0]   _zz_5518;
  wire       [15:0]   _zz_5519;
  wire       [15:0]   _zz_5520;
  wire       [15:0]   _zz_5521;
  wire       [15:0]   _zz_5522;
  wire       [15:0]   _zz_5523;
  wire       [15:0]   _zz_5524;
  wire       [15:0]   _zz_5525;
  wire       [15:0]   _zz_5526;
  wire       [15:0]   _zz_5527;
  wire       [15:0]   _zz_5528;
  wire       [15:0]   _zz_5529;
  wire       [15:0]   _zz_5530;
  wire       [15:0]   _zz_5531;
  wire       [15:0]   _zz_5532;
  wire       [15:0]   _zz_5533;
  wire       [15:0]   _zz_5534;
  wire       [15:0]   _zz_5535;
  wire       [15:0]   _zz_5536;
  wire       [15:0]   _zz_5537;
  wire       [15:0]   _zz_5538;
  wire       [15:0]   _zz_5539;
  wire       [15:0]   _zz_5540;
  wire       [15:0]   _zz_5541;
  wire       [15:0]   _zz_5542;
  wire       [15:0]   _zz_5543;
  wire       [15:0]   _zz_5544;
  wire       [15:0]   _zz_5545;
  wire       [15:0]   _zz_5546;
  wire       [15:0]   _zz_5547;
  wire       [15:0]   _zz_5548;
  wire       [15:0]   _zz_5549;
  wire       [15:0]   _zz_5550;
  wire       [15:0]   _zz_5551;
  wire       [15:0]   _zz_5552;
  wire       [15:0]   _zz_5553;
  wire       [15:0]   _zz_5554;
  wire       [15:0]   _zz_5555;
  wire       [15:0]   _zz_5556;
  wire       [15:0]   _zz_5557;
  wire       [15:0]   _zz_5558;
  wire       [15:0]   _zz_5559;
  wire       [15:0]   _zz_5560;
  wire       [15:0]   _zz_5561;
  wire       [15:0]   _zz_5562;
  wire       [15:0]   _zz_5563;
  wire       [15:0]   _zz_5564;
  wire       [15:0]   _zz_5565;
  wire       [15:0]   _zz_5566;
  wire       [15:0]   _zz_5567;
  wire       [15:0]   _zz_5568;
  wire       [15:0]   _zz_5569;
  wire       [15:0]   _zz_5570;
  wire       [15:0]   _zz_5571;
  wire       [15:0]   _zz_5572;
  wire       [15:0]   _zz_5573;
  wire       [15:0]   _zz_5574;
  wire       [15:0]   _zz_5575;
  wire       [15:0]   _zz_5576;
  wire       [15:0]   _zz_5577;
  wire       [15:0]   _zz_5578;
  wire       [15:0]   _zz_5579;
  wire       [15:0]   _zz_5580;
  wire       [15:0]   _zz_5581;
  wire       [15:0]   _zz_5582;
  wire       [15:0]   _zz_5583;
  wire       [15:0]   _zz_5584;
  wire       [15:0]   _zz_5585;
  wire       [15:0]   _zz_5586;
  wire       [15:0]   _zz_5587;
  wire       [15:0]   _zz_5588;
  wire       [15:0]   _zz_5589;
  wire       [15:0]   _zz_5590;
  wire       [15:0]   _zz_5591;
  wire       [15:0]   _zz_5592;
  wire       [15:0]   _zz_5593;
  wire       [15:0]   _zz_5594;
  wire       [15:0]   _zz_5595;
  wire       [15:0]   _zz_5596;
  wire       [15:0]   _zz_5597;
  wire       [15:0]   _zz_5598;
  wire       [15:0]   _zz_5599;
  wire       [15:0]   _zz_5600;
  wire       [15:0]   _zz_5601;
  wire       [15:0]   _zz_5602;
  wire       [15:0]   _zz_5603;
  wire       [15:0]   _zz_5604;
  wire       [15:0]   _zz_5605;
  wire       [15:0]   _zz_5606;
  wire       [15:0]   _zz_5607;
  wire       [15:0]   _zz_5608;
  wire       [15:0]   _zz_5609;
  wire       [15:0]   _zz_5610;
  wire       [15:0]   _zz_5611;
  wire       [15:0]   _zz_5612;
  wire       [15:0]   _zz_5613;
  wire       [15:0]   _zz_5614;
  wire       [15:0]   _zz_5615;
  wire       [15:0]   _zz_5616;
  wire       [15:0]   _zz_5617;
  wire       [15:0]   _zz_5618;
  wire       [15:0]   _zz_5619;
  wire       [15:0]   _zz_5620;
  wire       [15:0]   _zz_5621;
  wire       [15:0]   _zz_5622;
  wire       [15:0]   _zz_5623;
  wire       [15:0]   _zz_5624;
  wire       [15:0]   _zz_5625;
  wire       [15:0]   _zz_5626;
  wire       [15:0]   _zz_5627;
  wire       [15:0]   _zz_5628;
  wire       [15:0]   _zz_5629;
  wire       [15:0]   _zz_5630;
  wire       [15:0]   _zz_5631;
  wire       [15:0]   _zz_5632;
  wire       [15:0]   _zz_5633;
  wire       [15:0]   _zz_5634;
  wire       [15:0]   _zz_5635;
  wire       [15:0]   _zz_5636;
  wire       [15:0]   _zz_5637;
  wire       [15:0]   _zz_5638;
  wire       [15:0]   _zz_5639;
  wire       [15:0]   _zz_5640;
  wire       [15:0]   _zz_5641;
  wire       [15:0]   _zz_5642;
  wire       [15:0]   _zz_5643;
  wire       [15:0]   _zz_5644;
  wire       [15:0]   _zz_5645;
  wire       [15:0]   _zz_5646;
  wire       [15:0]   _zz_5647;
  wire       [15:0]   _zz_5648;
  wire       [15:0]   _zz_5649;
  wire       [15:0]   _zz_5650;
  wire       [15:0]   _zz_5651;
  wire       [15:0]   _zz_5652;
  wire       [15:0]   _zz_5653;
  wire       [15:0]   _zz_5654;
  wire       [15:0]   _zz_5655;
  wire       [15:0]   _zz_5656;
  wire       [15:0]   _zz_5657;
  wire       [15:0]   _zz_5658;
  wire       [15:0]   _zz_5659;
  wire       [15:0]   _zz_5660;
  wire       [15:0]   _zz_5661;
  wire       [15:0]   _zz_5662;
  wire       [15:0]   _zz_5663;
  wire       [15:0]   _zz_5664;
  wire       [15:0]   _zz_5665;
  wire       [15:0]   _zz_5666;
  wire       [15:0]   _zz_5667;
  wire       [15:0]   _zz_5668;
  wire       [15:0]   _zz_5669;
  wire       [15:0]   _zz_5670;
  wire       [15:0]   _zz_5671;
  wire       [15:0]   _zz_5672;
  wire       [15:0]   _zz_5673;
  wire       [15:0]   _zz_5674;
  wire       [15:0]   _zz_5675;
  wire       [15:0]   _zz_5676;
  wire       [15:0]   _zz_5677;
  wire       [15:0]   _zz_5678;
  wire       [15:0]   _zz_5679;
  wire       [15:0]   _zz_5680;
  wire       [15:0]   _zz_5681;
  wire       [15:0]   _zz_5682;
  wire       [15:0]   _zz_5683;
  wire       [15:0]   _zz_5684;
  wire       [15:0]   _zz_5685;
  wire       [15:0]   _zz_5686;
  wire       [15:0]   _zz_5687;
  wire       [15:0]   _zz_5688;
  wire       [15:0]   _zz_5689;
  wire       [15:0]   _zz_5690;
  wire       [15:0]   _zz_5691;
  wire       [15:0]   _zz_5692;
  wire       [15:0]   _zz_5693;
  wire       [15:0]   _zz_5694;
  wire       [15:0]   _zz_5695;
  wire       [15:0]   _zz_5696;
  wire       [15:0]   _zz_5697;
  wire       [15:0]   _zz_5698;
  wire       [15:0]   _zz_5699;
  wire       [15:0]   _zz_5700;
  wire       [15:0]   _zz_5701;
  wire       [15:0]   _zz_5702;
  wire       [15:0]   _zz_5703;
  wire       [15:0]   _zz_5704;
  wire       [15:0]   _zz_5705;
  wire       [15:0]   _zz_5706;
  wire       [15:0]   _zz_5707;
  wire       [15:0]   _zz_5708;
  wire       [15:0]   _zz_5709;
  wire       [15:0]   _zz_5710;
  wire       [15:0]   _zz_5711;
  wire       [15:0]   _zz_5712;
  wire       [15:0]   _zz_5713;
  wire       [15:0]   _zz_5714;
  wire       [15:0]   _zz_5715;
  wire       [15:0]   _zz_5716;
  wire       [15:0]   _zz_5717;
  wire       [15:0]   _zz_5718;
  wire       [15:0]   _zz_5719;
  wire       [15:0]   _zz_5720;
  wire       [15:0]   _zz_5721;
  wire       [15:0]   _zz_5722;
  wire       [15:0]   _zz_5723;
  wire       [15:0]   _zz_5724;
  wire       [15:0]   _zz_5725;
  wire       [15:0]   _zz_5726;
  wire       [15:0]   _zz_5727;
  wire       [15:0]   _zz_5728;
  wire       [15:0]   _zz_5729;
  wire       [15:0]   _zz_5730;
  wire       [15:0]   _zz_5731;
  wire       [15:0]   _zz_5732;
  wire       [15:0]   _zz_5733;
  wire       [15:0]   _zz_5734;
  wire       [15:0]   _zz_5735;
  wire       [15:0]   _zz_5736;
  wire       [15:0]   _zz_5737;
  wire       [15:0]   _zz_5738;
  wire       [15:0]   _zz_5739;
  wire       [15:0]   _zz_5740;
  wire       [15:0]   _zz_5741;
  wire       [15:0]   _zz_5742;
  wire       [15:0]   _zz_5743;
  wire       [15:0]   _zz_5744;
  wire       [15:0]   _zz_5745;
  wire       [15:0]   _zz_5746;
  wire       [15:0]   _zz_5747;
  wire       [15:0]   _zz_5748;
  wire       [15:0]   _zz_5749;
  wire       [15:0]   _zz_5750;
  wire       [15:0]   _zz_5751;
  wire       [15:0]   _zz_5752;
  wire       [15:0]   _zz_5753;
  wire       [15:0]   _zz_5754;
  wire       [15:0]   _zz_5755;
  wire       [15:0]   _zz_5756;
  wire       [15:0]   _zz_5757;
  wire       [15:0]   _zz_5758;
  wire       [15:0]   _zz_5759;
  wire       [15:0]   _zz_5760;
  wire       [15:0]   _zz_5761;
  wire       [15:0]   _zz_5762;
  wire       [15:0]   _zz_5763;
  wire       [15:0]   _zz_5764;
  wire       [15:0]   _zz_5765;
  wire       [15:0]   _zz_5766;
  wire       [15:0]   _zz_5767;
  wire       [15:0]   _zz_5768;
  wire       [15:0]   _zz_5769;
  wire       [15:0]   _zz_5770;
  wire       [15:0]   _zz_5771;
  wire       [15:0]   _zz_5772;
  wire       [15:0]   _zz_5773;
  wire       [15:0]   _zz_5774;
  wire       [15:0]   _zz_5775;
  wire       [15:0]   _zz_5776;
  wire       [15:0]   _zz_5777;
  wire       [15:0]   _zz_5778;
  wire       [15:0]   _zz_5779;
  wire       [15:0]   _zz_5780;
  wire       [15:0]   _zz_5781;
  wire       [15:0]   _zz_5782;
  wire       [15:0]   _zz_5783;
  wire       [15:0]   _zz_5784;
  wire       [15:0]   _zz_5785;
  wire       [15:0]   _zz_5786;
  wire       [15:0]   _zz_5787;
  wire       [15:0]   _zz_5788;
  wire       [15:0]   _zz_5789;
  wire       [15:0]   _zz_5790;
  wire       [15:0]   _zz_5791;
  wire       [15:0]   _zz_5792;
  wire       [15:0]   _zz_5793;
  wire       [15:0]   _zz_5794;
  wire       [15:0]   _zz_5795;
  wire       [15:0]   _zz_5796;
  wire       [15:0]   _zz_5797;
  wire       [15:0]   _zz_5798;
  wire       [15:0]   _zz_5799;
  wire       [15:0]   _zz_5800;
  wire       [15:0]   _zz_5801;
  wire       [15:0]   _zz_5802;
  wire       [15:0]   _zz_5803;
  wire       [15:0]   _zz_5804;
  wire       [15:0]   _zz_5805;
  wire       [15:0]   _zz_5806;
  wire       [15:0]   _zz_5807;
  wire       [15:0]   _zz_5808;
  wire       [15:0]   _zz_5809;
  wire       [15:0]   _zz_5810;
  wire       [15:0]   _zz_5811;
  wire       [15:0]   _zz_5812;
  wire       [15:0]   _zz_5813;
  wire       [15:0]   _zz_5814;
  wire       [15:0]   _zz_5815;
  wire       [15:0]   _zz_5816;
  wire       [15:0]   _zz_5817;
  wire       [15:0]   _zz_5818;
  wire       [15:0]   _zz_5819;
  wire       [15:0]   _zz_5820;
  wire       [15:0]   _zz_5821;
  wire       [15:0]   _zz_5822;
  wire       [15:0]   _zz_5823;
  wire       [15:0]   _zz_5824;
  wire       [15:0]   _zz_5825;
  wire       [15:0]   _zz_5826;
  wire       [15:0]   _zz_5827;
  wire       [15:0]   _zz_5828;
  wire       [15:0]   _zz_5829;
  wire       [15:0]   _zz_5830;
  wire       [15:0]   _zz_5831;
  wire       [15:0]   _zz_5832;
  wire       [15:0]   _zz_5833;
  wire       [15:0]   _zz_5834;
  wire       [15:0]   _zz_5835;
  wire       [15:0]   _zz_5836;
  wire       [15:0]   _zz_5837;
  wire       [15:0]   _zz_5838;
  wire       [15:0]   _zz_5839;
  wire       [15:0]   _zz_5840;
  wire       [15:0]   _zz_5841;
  wire       [15:0]   _zz_5842;
  wire       [15:0]   _zz_5843;
  wire       [15:0]   _zz_5844;
  wire       [15:0]   _zz_5845;
  wire       [15:0]   _zz_5846;
  wire       [15:0]   _zz_5847;
  wire       [15:0]   _zz_5848;
  wire       [15:0]   _zz_5849;
  wire       [15:0]   _zz_5850;
  wire       [15:0]   _zz_5851;
  wire       [15:0]   _zz_5852;
  wire       [15:0]   _zz_5853;
  wire       [15:0]   _zz_5854;
  wire       [15:0]   _zz_5855;
  wire       [15:0]   _zz_5856;
  wire       [15:0]   _zz_5857;
  wire       [15:0]   _zz_5858;
  wire       [15:0]   _zz_5859;
  wire       [15:0]   _zz_5860;
  wire       [15:0]   _zz_5861;
  wire       [15:0]   _zz_5862;
  wire       [15:0]   _zz_5863;
  wire       [15:0]   _zz_5864;
  wire       [15:0]   _zz_5865;
  wire       [15:0]   _zz_5866;
  wire       [15:0]   _zz_5867;
  wire       [15:0]   _zz_5868;
  wire       [15:0]   _zz_5869;
  wire       [15:0]   _zz_5870;
  wire       [15:0]   _zz_5871;
  wire       [15:0]   _zz_5872;
  wire       [15:0]   _zz_5873;
  wire       [15:0]   _zz_5874;
  wire       [15:0]   _zz_5875;
  wire       [15:0]   _zz_5876;
  wire       [15:0]   _zz_5877;
  wire       [15:0]   _zz_5878;
  wire       [15:0]   _zz_5879;
  wire       [15:0]   _zz_5880;
  wire       [15:0]   _zz_5881;
  wire       [15:0]   _zz_5882;
  wire       [15:0]   _zz_5883;
  wire       [15:0]   _zz_5884;
  wire       [15:0]   _zz_5885;
  wire       [15:0]   _zz_5886;
  wire       [15:0]   _zz_5887;
  wire       [15:0]   _zz_5888;
  wire       [15:0]   _zz_5889;
  wire       [15:0]   _zz_5890;
  wire       [15:0]   _zz_5891;
  wire       [15:0]   _zz_5892;
  wire       [15:0]   _zz_5893;
  wire       [15:0]   _zz_5894;
  wire       [15:0]   _zz_5895;
  wire       [15:0]   _zz_5896;
  wire       [15:0]   _zz_5897;
  wire       [15:0]   _zz_5898;
  wire       [15:0]   _zz_5899;
  wire       [15:0]   _zz_5900;
  wire       [15:0]   _zz_5901;
  wire       [15:0]   _zz_5902;
  wire       [15:0]   _zz_5903;
  wire       [15:0]   _zz_5904;
  wire       [15:0]   _zz_5905;
  wire       [15:0]   _zz_5906;
  wire       [15:0]   _zz_5907;
  wire       [15:0]   _zz_5908;
  wire       [15:0]   _zz_5909;
  wire       [15:0]   _zz_5910;
  wire       [15:0]   _zz_5911;
  wire       [15:0]   _zz_5912;
  wire       [15:0]   _zz_5913;
  wire       [15:0]   _zz_5914;
  wire       [15:0]   _zz_5915;
  wire       [15:0]   _zz_5916;
  wire       [15:0]   _zz_5917;
  wire       [15:0]   _zz_5918;
  wire       [15:0]   _zz_5919;
  wire       [15:0]   _zz_5920;
  wire       [15:0]   _zz_5921;
  wire       [15:0]   _zz_5922;
  wire       [15:0]   _zz_5923;
  wire       [15:0]   _zz_5924;
  wire       [15:0]   _zz_5925;
  wire       [15:0]   _zz_5926;
  wire       [15:0]   _zz_5927;
  wire       [15:0]   _zz_5928;
  wire       [15:0]   _zz_5929;
  wire       [15:0]   _zz_5930;
  wire       [15:0]   _zz_5931;
  wire       [15:0]   _zz_5932;
  wire       [15:0]   _zz_5933;
  wire       [15:0]   _zz_5934;
  wire       [15:0]   _zz_5935;
  wire       [15:0]   _zz_5936;
  wire       [15:0]   _zz_5937;
  wire       [15:0]   _zz_5938;
  wire       [15:0]   _zz_5939;
  wire       [15:0]   _zz_5940;
  wire       [15:0]   _zz_5941;
  wire       [15:0]   _zz_5942;
  wire       [15:0]   _zz_5943;
  wire       [15:0]   _zz_5944;
  wire       [15:0]   _zz_5945;
  wire       [15:0]   _zz_5946;
  wire       [15:0]   _zz_5947;
  wire       [15:0]   _zz_5948;
  wire       [15:0]   _zz_5949;
  wire       [15:0]   _zz_5950;
  wire       [15:0]   _zz_5951;
  wire       [15:0]   _zz_5952;
  wire       [15:0]   _zz_5953;
  wire       [15:0]   _zz_5954;
  wire       [15:0]   _zz_5955;
  wire       [15:0]   _zz_5956;
  wire       [15:0]   _zz_5957;
  wire       [15:0]   _zz_5958;
  wire       [15:0]   _zz_5959;
  wire       [15:0]   _zz_5960;
  wire       [15:0]   _zz_5961;
  wire       [15:0]   _zz_5962;
  wire       [15:0]   _zz_5963;
  wire       [15:0]   _zz_5964;
  wire       [15:0]   _zz_5965;
  wire       [15:0]   _zz_5966;
  wire       [15:0]   _zz_5967;
  wire       [15:0]   _zz_5968;
  wire       [15:0]   _zz_5969;
  wire       [15:0]   _zz_5970;
  wire       [15:0]   _zz_5971;
  wire       [15:0]   _zz_5972;
  wire       [15:0]   _zz_5973;
  wire       [15:0]   _zz_5974;
  wire       [15:0]   _zz_5975;
  wire       [15:0]   _zz_5976;
  wire       [15:0]   _zz_5977;
  wire       [15:0]   _zz_5978;
  wire       [15:0]   _zz_5979;
  wire       [15:0]   _zz_5980;
  wire       [15:0]   _zz_5981;
  wire       [15:0]   _zz_5982;
  wire       [15:0]   _zz_5983;
  wire       [15:0]   _zz_5984;
  wire       [15:0]   _zz_5985;
  wire       [15:0]   _zz_5986;
  wire       [15:0]   _zz_5987;
  wire       [15:0]   _zz_5988;
  wire       [15:0]   _zz_5989;
  wire       [15:0]   _zz_5990;
  wire       [15:0]   _zz_5991;
  wire       [15:0]   _zz_5992;
  wire       [15:0]   _zz_5993;
  wire       [15:0]   _zz_5994;
  wire       [15:0]   _zz_5995;
  wire       [15:0]   _zz_5996;
  wire       [15:0]   _zz_5997;
  wire       [15:0]   _zz_5998;
  wire       [15:0]   _zz_5999;
  wire       [15:0]   _zz_6000;
  wire       [15:0]   _zz_6001;
  wire       [15:0]   _zz_6002;
  wire       [15:0]   _zz_6003;
  wire       [15:0]   _zz_6004;
  wire       [15:0]   _zz_6005;
  wire       [15:0]   _zz_6006;
  wire       [15:0]   _zz_6007;
  wire       [15:0]   _zz_6008;
  wire       [15:0]   _zz_6009;
  wire       [15:0]   _zz_6010;
  wire       [15:0]   _zz_6011;
  wire       [15:0]   _zz_6012;
  wire       [15:0]   _zz_6013;
  wire       [15:0]   _zz_6014;
  wire       [15:0]   _zz_6015;
  wire       [15:0]   _zz_6016;
  wire       [15:0]   _zz_6017;
  wire       [15:0]   _zz_6018;
  wire       [15:0]   _zz_6019;
  wire       [15:0]   _zz_6020;
  wire       [15:0]   _zz_6021;
  wire       [15:0]   _zz_6022;
  wire       [15:0]   _zz_6023;
  wire       [15:0]   _zz_6024;
  wire       [15:0]   _zz_6025;
  wire       [15:0]   _zz_6026;
  wire       [15:0]   _zz_6027;
  wire       [15:0]   _zz_6028;
  wire       [15:0]   _zz_6029;
  wire       [15:0]   _zz_6030;
  wire       [15:0]   _zz_6031;
  wire       [15:0]   _zz_6032;
  wire       [15:0]   _zz_6033;
  wire       [15:0]   _zz_6034;
  wire       [15:0]   _zz_6035;
  wire       [15:0]   _zz_6036;
  wire       [15:0]   _zz_6037;
  wire       [15:0]   _zz_6038;
  wire       [15:0]   _zz_6039;
  wire       [15:0]   _zz_6040;
  wire       [15:0]   _zz_6041;
  wire       [15:0]   _zz_6042;
  wire       [15:0]   _zz_6043;
  wire       [15:0]   _zz_6044;
  wire       [15:0]   _zz_6045;
  wire       [15:0]   _zz_6046;
  wire       [15:0]   _zz_6047;
  wire       [15:0]   _zz_6048;
  wire       [15:0]   _zz_6049;
  wire       [15:0]   _zz_6050;
  wire       [15:0]   _zz_6051;
  wire       [15:0]   _zz_6052;
  wire       [15:0]   _zz_6053;
  wire       [15:0]   _zz_6054;
  wire       [15:0]   _zz_6055;
  wire       [15:0]   _zz_6056;
  wire       [15:0]   _zz_6057;
  wire       [15:0]   _zz_6058;
  wire       [15:0]   _zz_6059;
  wire       [15:0]   _zz_6060;
  wire       [15:0]   _zz_6061;
  wire       [15:0]   _zz_6062;
  wire       [15:0]   _zz_6063;
  wire       [15:0]   _zz_6064;
  wire       [15:0]   _zz_6065;
  wire       [15:0]   _zz_6066;
  wire       [15:0]   _zz_6067;
  wire       [15:0]   _zz_6068;
  wire       [15:0]   _zz_6069;
  wire       [15:0]   _zz_6070;
  wire       [15:0]   _zz_6071;
  wire       [15:0]   _zz_6072;
  wire       [15:0]   _zz_6073;
  wire       [15:0]   _zz_6074;
  wire       [15:0]   _zz_6075;
  wire       [15:0]   _zz_6076;
  wire       [15:0]   _zz_6077;
  wire       [15:0]   _zz_6078;
  wire       [15:0]   _zz_6079;
  wire       [15:0]   _zz_6080;
  wire       [15:0]   _zz_6081;
  wire       [15:0]   _zz_6082;
  wire       [15:0]   _zz_6083;
  wire       [15:0]   _zz_6084;
  wire       [15:0]   _zz_6085;
  wire       [15:0]   _zz_6086;
  wire       [15:0]   _zz_6087;
  wire       [15:0]   _zz_6088;
  wire       [15:0]   _zz_6089;
  wire       [15:0]   _zz_6090;
  wire       [15:0]   _zz_6091;
  wire       [15:0]   _zz_6092;
  wire       [15:0]   _zz_6093;
  wire       [15:0]   _zz_6094;
  wire       [15:0]   _zz_6095;
  wire       [15:0]   _zz_6096;
  wire       [15:0]   _zz_6097;
  wire       [15:0]   _zz_6098;
  wire       [15:0]   _zz_6099;
  wire       [15:0]   _zz_6100;
  wire       [15:0]   _zz_6101;
  wire       [15:0]   _zz_6102;
  wire       [15:0]   _zz_6103;
  wire       [15:0]   _zz_6104;
  wire       [15:0]   _zz_6105;
  wire       [15:0]   _zz_6106;
  wire       [15:0]   _zz_6107;
  wire       [15:0]   _zz_6108;
  wire       [15:0]   _zz_6109;
  wire       [15:0]   _zz_6110;
  wire       [15:0]   _zz_6111;
  wire       [15:0]   _zz_6112;
  wire       [15:0]   _zz_6113;
  wire       [15:0]   _zz_6114;
  wire       [15:0]   _zz_6115;
  wire       [15:0]   _zz_6116;
  wire       [15:0]   _zz_6117;
  wire       [15:0]   _zz_6118;
  wire       [15:0]   _zz_6119;
  wire       [15:0]   _zz_6120;
  wire       [15:0]   _zz_6121;
  wire       [15:0]   _zz_6122;
  wire       [15:0]   _zz_6123;
  wire       [15:0]   _zz_6124;
  wire       [15:0]   _zz_6125;
  wire       [15:0]   _zz_6126;
  wire       [15:0]   _zz_6127;
  wire       [15:0]   _zz_6128;
  wire       [15:0]   _zz_6129;
  wire       [15:0]   _zz_6130;
  wire       [15:0]   _zz_6131;
  wire       [15:0]   _zz_6132;
  wire       [15:0]   _zz_6133;
  wire       [15:0]   _zz_6134;
  wire       [15:0]   _zz_6135;
  wire       [15:0]   _zz_6136;
  wire       [15:0]   _zz_6137;
  wire       [15:0]   _zz_6138;
  wire       [15:0]   _zz_6139;
  wire       [15:0]   _zz_6140;
  wire       [15:0]   _zz_6141;
  wire       [15:0]   _zz_6142;
  wire       [15:0]   _zz_6143;
  wire       [15:0]   _zz_6144;
  wire       [15:0]   _zz_6145;
  wire       [15:0]   _zz_6146;
  wire       [15:0]   _zz_6147;
  wire       [15:0]   _zz_6148;
  wire       [15:0]   _zz_6149;
  wire       [15:0]   _zz_6150;
  wire       [15:0]   _zz_6151;
  wire       [15:0]   _zz_6152;
  wire       [15:0]   _zz_6153;
  wire       [15:0]   _zz_6154;
  wire       [15:0]   _zz_6155;
  wire       [15:0]   _zz_6156;
  wire       [15:0]   _zz_6157;
  wire       [15:0]   _zz_6158;
  wire       [15:0]   _zz_6159;
  wire       [15:0]   _zz_6160;
  wire       [15:0]   _zz_6161;
  wire       [15:0]   _zz_6162;
  wire       [15:0]   _zz_6163;
  wire       [15:0]   _zz_6164;
  wire       [15:0]   _zz_6165;
  wire       [15:0]   _zz_6166;
  wire       [15:0]   _zz_6167;
  wire       [15:0]   _zz_6168;
  wire       [15:0]   _zz_6169;
  wire       [15:0]   _zz_6170;
  wire       [15:0]   _zz_6171;
  wire       [15:0]   _zz_6172;
  wire       [15:0]   _zz_6173;
  wire       [15:0]   _zz_6174;
  wire       [15:0]   _zz_6175;
  wire       [15:0]   _zz_6176;
  wire       [15:0]   _zz_6177;
  wire       [15:0]   _zz_6178;
  wire       [15:0]   _zz_6179;
  wire       [15:0]   _zz_6180;
  wire       [15:0]   _zz_6181;
  wire       [15:0]   _zz_6182;
  wire       [15:0]   _zz_6183;
  wire       [15:0]   _zz_6184;
  wire       [15:0]   _zz_6185;
  wire       [15:0]   _zz_6186;
  wire       [15:0]   _zz_6187;
  wire       [15:0]   _zz_6188;
  wire       [15:0]   _zz_6189;
  wire       [15:0]   _zz_6190;
  wire       [15:0]   _zz_6191;
  wire       [15:0]   _zz_6192;
  wire       [15:0]   _zz_6193;
  wire       [15:0]   _zz_6194;
  wire       [15:0]   _zz_6195;
  wire       [15:0]   _zz_6196;
  wire       [15:0]   _zz_6197;
  wire       [15:0]   _zz_6198;
  wire       [15:0]   _zz_6199;
  wire       [15:0]   _zz_6200;
  wire       [15:0]   _zz_6201;
  wire       [15:0]   _zz_6202;
  wire       [15:0]   _zz_6203;
  wire       [15:0]   _zz_6204;
  wire       [15:0]   _zz_6205;
  wire       [15:0]   _zz_6206;
  wire       [15:0]   _zz_6207;
  wire       [15:0]   _zz_6208;
  wire       [15:0]   _zz_6209;
  wire       [15:0]   _zz_6210;
  wire       [15:0]   _zz_6211;
  wire       [15:0]   _zz_6212;
  wire       [15:0]   _zz_6213;
  wire       [15:0]   _zz_6214;
  wire       [15:0]   _zz_6215;
  wire       [15:0]   _zz_6216;
  wire       [15:0]   _zz_6217;
  wire       [15:0]   _zz_6218;
  wire       [15:0]   _zz_6219;
  wire       [15:0]   _zz_6220;
  wire       [15:0]   _zz_6221;
  wire       [15:0]   _zz_6222;
  wire       [15:0]   _zz_6223;
  wire       [15:0]   _zz_6224;
  wire       [15:0]   _zz_6225;
  wire       [15:0]   _zz_6226;
  wire       [15:0]   _zz_6227;
  wire       [15:0]   _zz_6228;
  wire       [15:0]   _zz_6229;
  wire       [15:0]   _zz_6230;
  wire       [15:0]   _zz_6231;
  wire       [15:0]   _zz_6232;
  wire       [15:0]   _zz_6233;
  wire       [15:0]   _zz_6234;
  wire       [15:0]   _zz_6235;
  wire       [15:0]   _zz_6236;
  wire       [15:0]   _zz_6237;
  wire       [15:0]   _zz_6238;
  wire       [15:0]   _zz_6239;
  wire       [15:0]   _zz_6240;
  wire       [15:0]   _zz_6241;
  wire       [15:0]   _zz_6242;
  wire       [15:0]   _zz_6243;
  wire       [15:0]   _zz_6244;
  wire       [15:0]   _zz_6245;
  wire       [15:0]   _zz_6246;
  wire       [15:0]   _zz_6247;
  wire       [15:0]   _zz_6248;
  wire       [15:0]   _zz_6249;
  wire       [15:0]   _zz_6250;
  wire       [15:0]   _zz_6251;
  wire       [15:0]   _zz_6252;
  wire       [15:0]   _zz_6253;
  wire       [15:0]   _zz_6254;
  wire       [15:0]   _zz_6255;
  wire       [15:0]   _zz_6256;
  wire       [15:0]   _zz_6257;
  wire       [15:0]   _zz_6258;
  wire       [15:0]   _zz_6259;
  wire       [15:0]   _zz_6260;
  wire       [15:0]   _zz_6261;
  wire       [15:0]   _zz_6262;
  wire       [15:0]   _zz_6263;
  wire       [15:0]   _zz_6264;
  wire       [15:0]   _zz_6265;
  wire       [15:0]   _zz_6266;
  wire       [15:0]   _zz_6267;
  wire       [15:0]   _zz_6268;
  wire       [15:0]   _zz_6269;
  wire       [15:0]   _zz_6270;
  wire       [15:0]   _zz_6271;
  wire       [15:0]   _zz_6272;
  wire       [15:0]   _zz_6273;
  wire       [15:0]   _zz_6274;
  wire       [15:0]   _zz_6275;
  wire       [15:0]   _zz_6276;
  wire       [15:0]   _zz_6277;
  wire       [15:0]   _zz_6278;
  wire       [15:0]   _zz_6279;
  wire       [15:0]   _zz_6280;
  wire       [15:0]   _zz_6281;
  wire       [15:0]   _zz_6282;
  wire       [15:0]   _zz_6283;
  wire       [15:0]   _zz_6284;
  wire       [15:0]   _zz_6285;
  wire       [15:0]   _zz_6286;
  wire       [15:0]   _zz_6287;
  wire       [15:0]   _zz_6288;
  wire       [15:0]   _zz_6289;
  wire       [15:0]   _zz_6290;
  wire       [15:0]   _zz_6291;
  wire       [15:0]   _zz_6292;
  wire       [15:0]   _zz_6293;
  wire       [15:0]   _zz_6294;
  wire       [15:0]   _zz_6295;
  wire       [15:0]   _zz_6296;
  wire       [15:0]   _zz_6297;
  wire       [15:0]   _zz_6298;
  wire       [15:0]   _zz_6299;
  wire       [15:0]   _zz_6300;
  wire       [15:0]   _zz_6301;
  wire       [15:0]   _zz_6302;
  wire       [15:0]   _zz_6303;
  wire       [15:0]   _zz_6304;
  wire       [15:0]   _zz_6305;
  wire       [15:0]   _zz_6306;
  wire       [15:0]   _zz_6307;
  wire       [15:0]   _zz_6308;
  wire       [15:0]   _zz_6309;
  wire       [15:0]   _zz_6310;
  wire       [15:0]   _zz_6311;
  wire       [15:0]   _zz_6312;
  wire       [15:0]   _zz_6313;
  wire       [15:0]   _zz_6314;
  wire       [15:0]   _zz_6315;
  wire       [15:0]   _zz_6316;
  wire       [15:0]   _zz_6317;
  wire       [15:0]   _zz_6318;
  wire       [15:0]   _zz_6319;
  wire       [15:0]   _zz_6320;
  wire       [15:0]   _zz_6321;
  wire       [15:0]   _zz_6322;
  wire       [15:0]   _zz_6323;
  wire       [15:0]   _zz_6324;
  wire       [15:0]   _zz_6325;
  wire       [15:0]   _zz_6326;
  wire       [15:0]   _zz_6327;
  wire       [15:0]   _zz_6328;
  wire       [15:0]   _zz_6329;
  wire       [15:0]   _zz_6330;
  wire       [15:0]   _zz_6331;
  wire       [15:0]   _zz_6332;
  wire       [15:0]   _zz_6333;
  wire       [15:0]   _zz_6334;
  wire       [15:0]   _zz_6335;
  wire       [15:0]   _zz_6336;
  wire       [15:0]   _zz_6337;
  wire       [15:0]   _zz_6338;
  wire       [15:0]   _zz_6339;
  wire       [15:0]   _zz_6340;
  wire       [15:0]   _zz_6341;
  wire       [15:0]   _zz_6342;
  wire       [15:0]   _zz_6343;
  wire       [15:0]   _zz_6344;
  wire       [15:0]   _zz_6345;
  wire       [15:0]   _zz_6346;
  wire       [15:0]   _zz_6347;
  wire       [15:0]   _zz_6348;
  wire       [15:0]   _zz_6349;
  wire       [15:0]   _zz_6350;
  wire       [15:0]   _zz_6351;
  wire       [15:0]   _zz_6352;
  wire       [15:0]   _zz_6353;
  wire       [15:0]   _zz_6354;
  wire       [15:0]   _zz_6355;
  wire       [15:0]   _zz_6356;
  wire       [15:0]   _zz_6357;
  wire       [15:0]   _zz_6358;
  wire       [15:0]   _zz_6359;
  wire       [15:0]   _zz_6360;
  wire       [15:0]   _zz_6361;
  wire       [15:0]   _zz_6362;
  wire       [15:0]   _zz_6363;
  wire       [15:0]   _zz_6364;
  wire       [15:0]   _zz_6365;
  wire       [15:0]   _zz_6366;
  wire       [15:0]   _zz_6367;
  wire       [15:0]   _zz_6368;
  wire       [15:0]   _zz_6369;
  wire       [15:0]   _zz_6370;
  wire       [15:0]   _zz_6371;
  wire       [15:0]   _zz_6372;
  wire       [15:0]   _zz_6373;
  wire       [15:0]   _zz_6374;
  wire       [15:0]   _zz_6375;
  wire       [15:0]   _zz_6376;
  wire       [15:0]   _zz_6377;
  wire       [15:0]   _zz_6378;
  wire       [15:0]   _zz_6379;
  wire       [15:0]   _zz_6380;
  wire       [15:0]   _zz_6381;
  wire       [15:0]   _zz_6382;
  wire       [15:0]   _zz_6383;
  wire       [15:0]   _zz_6384;
  wire       [15:0]   _zz_6385;
  wire       [15:0]   _zz_6386;
  wire       [15:0]   _zz_6387;
  wire       [15:0]   _zz_6388;
  wire       [15:0]   _zz_6389;
  wire       [15:0]   _zz_6390;
  wire       [15:0]   _zz_6391;
  wire       [15:0]   _zz_6392;
  wire       [15:0]   _zz_6393;
  wire       [15:0]   _zz_6394;
  wire       [15:0]   _zz_6395;
  wire       [15:0]   _zz_6396;
  wire       [15:0]   _zz_6397;
  wire       [15:0]   _zz_6398;
  wire       [15:0]   _zz_6399;
  wire       [15:0]   _zz_6400;
  wire       [15:0]   _zz_6401;
  wire       [15:0]   _zz_6402;
  wire       [15:0]   _zz_6403;
  wire       [15:0]   _zz_6404;
  wire       [15:0]   _zz_6405;
  wire       [15:0]   _zz_6406;
  wire       [15:0]   _zz_6407;
  wire       [15:0]   _zz_6408;
  wire       [15:0]   _zz_6409;
  wire       [15:0]   _zz_6410;
  wire       [15:0]   _zz_6411;
  wire       [15:0]   _zz_6412;
  wire       [15:0]   _zz_6413;
  wire       [15:0]   _zz_6414;
  wire       [15:0]   _zz_6415;
  wire       [15:0]   _zz_6416;
  wire       [15:0]   _zz_6417;
  wire       [15:0]   _zz_6418;
  wire       [15:0]   _zz_6419;
  wire       [15:0]   _zz_6420;
  wire       [15:0]   _zz_6421;
  wire       [15:0]   _zz_6422;
  wire       [15:0]   _zz_6423;
  wire       [15:0]   _zz_6424;
  wire       [15:0]   _zz_6425;
  wire       [15:0]   _zz_6426;
  wire       [15:0]   _zz_6427;
  wire       [15:0]   _zz_6428;
  wire       [15:0]   _zz_6429;
  wire       [15:0]   _zz_6430;
  wire       [15:0]   _zz_6431;
  wire       [15:0]   _zz_6432;
  wire       [15:0]   _zz_6433;
  wire       [15:0]   _zz_6434;
  wire       [15:0]   _zz_6435;
  wire       [15:0]   _zz_6436;
  wire       [15:0]   _zz_6437;
  wire       [15:0]   _zz_6438;
  wire       [15:0]   _zz_6439;
  wire       [15:0]   _zz_6440;
  wire       [15:0]   _zz_6441;
  wire       [15:0]   _zz_6442;
  wire       [15:0]   _zz_6443;
  wire       [15:0]   _zz_6444;
  wire       [15:0]   _zz_6445;
  wire       [15:0]   _zz_6446;
  wire       [15:0]   _zz_6447;
  wire       [15:0]   _zz_6448;
  wire       [15:0]   _zz_6449;
  wire       [15:0]   _zz_6450;
  wire       [15:0]   _zz_6451;
  wire       [15:0]   _zz_6452;
  wire       [15:0]   _zz_6453;
  wire       [15:0]   _zz_6454;
  wire       [15:0]   _zz_6455;
  wire       [15:0]   _zz_6456;
  wire       [15:0]   _zz_6457;
  wire       [15:0]   _zz_6458;
  wire       [15:0]   _zz_6459;
  wire       [15:0]   _zz_6460;
  wire       [15:0]   _zz_6461;
  wire       [15:0]   _zz_6462;
  wire       [15:0]   _zz_6463;
  wire       [15:0]   _zz_6464;
  wire       [15:0]   _zz_6465;
  wire       [15:0]   _zz_6466;
  wire       [15:0]   _zz_6467;
  wire       [15:0]   _zz_6468;
  wire       [15:0]   _zz_6469;
  wire       [15:0]   _zz_6470;
  wire       [15:0]   _zz_6471;
  wire       [15:0]   _zz_6472;
  wire       [15:0]   _zz_6473;
  wire       [15:0]   _zz_6474;
  wire       [15:0]   _zz_6475;
  wire       [15:0]   _zz_6476;
  wire       [15:0]   _zz_6477;
  wire       [15:0]   _zz_6478;
  wire       [15:0]   _zz_6479;
  wire       [15:0]   _zz_6480;
  wire       [15:0]   _zz_6481;
  wire       [15:0]   _zz_6482;
  wire       [15:0]   _zz_6483;
  wire       [15:0]   _zz_6484;
  wire       [15:0]   _zz_6485;
  wire       [15:0]   _zz_6486;
  wire       [15:0]   _zz_6487;
  wire       [15:0]   _zz_6488;
  wire       [15:0]   _zz_6489;
  wire       [15:0]   _zz_6490;
  wire       [15:0]   _zz_6491;
  wire       [15:0]   _zz_6492;
  wire       [15:0]   _zz_6493;
  wire       [15:0]   _zz_6494;
  wire       [15:0]   _zz_6495;
  wire       [15:0]   _zz_6496;
  wire       [15:0]   _zz_6497;
  wire       [15:0]   _zz_6498;
  wire       [15:0]   _zz_6499;
  wire       [15:0]   _zz_6500;
  wire       [15:0]   _zz_6501;
  wire       [15:0]   _zz_6502;
  wire       [15:0]   _zz_6503;
  wire       [15:0]   _zz_6504;
  wire       [15:0]   _zz_6505;
  wire       [15:0]   _zz_6506;
  wire       [15:0]   _zz_6507;
  wire       [15:0]   _zz_6508;
  wire       [15:0]   _zz_6509;
  wire       [15:0]   _zz_6510;
  wire       [15:0]   _zz_6511;
  wire       [15:0]   _zz_6512;
  wire       [15:0]   _zz_6513;
  wire       [15:0]   _zz_6514;
  wire       [15:0]   _zz_6515;
  wire       [15:0]   _zz_6516;
  wire       [15:0]   _zz_6517;
  wire       [15:0]   _zz_6518;
  wire       [15:0]   _zz_6519;
  wire       [15:0]   _zz_6520;
  wire       [15:0]   _zz_6521;
  wire       [15:0]   _zz_6522;
  wire       [15:0]   _zz_6523;
  wire       [15:0]   _zz_6524;
  wire       [15:0]   _zz_6525;
  wire       [15:0]   _zz_6526;
  wire       [15:0]   _zz_6527;
  wire       [15:0]   _zz_6528;
  wire       [15:0]   _zz_6529;
  wire       [15:0]   _zz_6530;
  wire       [15:0]   _zz_6531;
  wire       [15:0]   _zz_6532;
  wire       [15:0]   _zz_6533;
  wire       [15:0]   _zz_6534;
  wire       [15:0]   _zz_6535;
  wire       [15:0]   _zz_6536;
  wire       [15:0]   _zz_6537;
  wire       [15:0]   _zz_6538;
  wire       [15:0]   _zz_6539;
  wire       [15:0]   _zz_6540;
  wire       [15:0]   _zz_6541;
  wire       [15:0]   _zz_6542;
  wire       [15:0]   _zz_6543;
  wire       [15:0]   _zz_6544;
  wire       [15:0]   _zz_6545;
  wire       [15:0]   _zz_6546;
  wire       [15:0]   _zz_6547;
  wire       [15:0]   _zz_6548;
  wire       [15:0]   _zz_6549;
  wire       [15:0]   _zz_6550;
  wire       [15:0]   _zz_6551;
  wire       [15:0]   _zz_6552;
  wire       [15:0]   _zz_6553;
  wire       [15:0]   _zz_6554;
  wire       [15:0]   _zz_6555;
  wire       [15:0]   _zz_6556;
  wire       [15:0]   _zz_6557;
  wire       [15:0]   _zz_6558;
  wire       [15:0]   _zz_6559;
  wire       [15:0]   _zz_6560;
  wire       [15:0]   _zz_6561;
  wire       [15:0]   _zz_6562;
  wire       [15:0]   _zz_6563;
  wire       [15:0]   _zz_6564;
  wire       [15:0]   _zz_6565;
  wire       [15:0]   _zz_6566;
  wire       [15:0]   _zz_6567;
  wire       [15:0]   _zz_6568;
  wire       [15:0]   _zz_6569;
  wire       [15:0]   _zz_6570;
  wire       [15:0]   _zz_6571;
  wire       [15:0]   _zz_6572;
  wire       [15:0]   _zz_6573;
  wire       [15:0]   _zz_6574;
  wire       [15:0]   _zz_6575;
  wire       [15:0]   _zz_6576;
  wire       [15:0]   _zz_6577;
  wire       [15:0]   _zz_6578;
  wire       [15:0]   _zz_6579;
  wire       [15:0]   _zz_6580;
  wire       [15:0]   _zz_6581;
  wire       [15:0]   _zz_6582;
  wire       [15:0]   _zz_6583;
  wire       [15:0]   _zz_6584;
  wire       [15:0]   _zz_6585;
  wire       [15:0]   _zz_6586;
  wire       [15:0]   _zz_6587;
  wire       [15:0]   _zz_6588;
  wire       [15:0]   _zz_6589;
  wire       [15:0]   _zz_6590;
  wire       [15:0]   _zz_6591;
  wire       [15:0]   _zz_6592;
  wire       [15:0]   _zz_6593;
  wire       [15:0]   _zz_6594;
  wire       [15:0]   _zz_6595;
  wire       [15:0]   _zz_6596;
  wire       [15:0]   _zz_6597;
  wire       [15:0]   _zz_6598;
  wire       [15:0]   _zz_6599;
  wire       [15:0]   _zz_6600;
  wire       [15:0]   _zz_6601;
  wire       [15:0]   _zz_6602;
  wire       [15:0]   _zz_6603;
  wire       [15:0]   _zz_6604;
  wire       [15:0]   _zz_6605;
  wire       [15:0]   _zz_6606;
  wire       [15:0]   _zz_6607;
  wire       [15:0]   _zz_6608;
  wire       [15:0]   _zz_6609;
  wire       [15:0]   _zz_6610;
  wire       [15:0]   _zz_6611;
  wire       [15:0]   _zz_6612;
  wire       [15:0]   _zz_6613;
  wire       [15:0]   _zz_6614;
  wire       [15:0]   _zz_6615;
  wire       [15:0]   _zz_6616;
  wire       [15:0]   _zz_6617;
  wire       [15:0]   _zz_6618;
  wire       [15:0]   _zz_6619;
  wire       [15:0]   _zz_6620;
  wire       [15:0]   _zz_6621;
  wire       [15:0]   _zz_6622;
  wire       [15:0]   _zz_6623;
  wire       [15:0]   _zz_6624;
  wire       [15:0]   _zz_6625;
  wire       [15:0]   _zz_6626;
  wire       [15:0]   _zz_6627;
  wire       [15:0]   _zz_6628;
  wire       [15:0]   _zz_6629;
  wire       [15:0]   _zz_6630;
  wire       [15:0]   _zz_6631;
  wire       [15:0]   _zz_6632;
  wire       [15:0]   _zz_6633;
  wire       [15:0]   _zz_6634;
  wire       [15:0]   _zz_6635;
  wire       [15:0]   _zz_6636;
  wire       [15:0]   _zz_6637;
  wire       [15:0]   _zz_6638;
  wire       [15:0]   _zz_6639;
  wire       [15:0]   _zz_6640;
  wire       [15:0]   _zz_6641;
  wire       [15:0]   _zz_6642;
  wire       [15:0]   _zz_6643;
  wire       [15:0]   _zz_6644;
  wire       [15:0]   _zz_6645;
  wire       [15:0]   _zz_6646;
  wire       [15:0]   _zz_6647;
  wire       [15:0]   _zz_6648;
  wire       [15:0]   _zz_6649;
  wire       [15:0]   _zz_6650;
  wire       [15:0]   _zz_6651;
  wire       [15:0]   _zz_6652;
  wire       [15:0]   _zz_6653;
  wire       [15:0]   _zz_6654;
  wire       [15:0]   _zz_6655;
  wire       [15:0]   _zz_6656;
  wire       [15:0]   _zz_6657;
  wire       [15:0]   _zz_6658;
  wire       [15:0]   _zz_6659;
  wire       [15:0]   _zz_6660;
  wire       [15:0]   _zz_6661;
  wire       [15:0]   _zz_6662;
  wire       [15:0]   _zz_6663;
  wire       [15:0]   _zz_6664;
  wire       [15:0]   _zz_6665;
  wire       [15:0]   _zz_6666;
  wire       [15:0]   _zz_6667;
  wire       [15:0]   _zz_6668;
  wire       [15:0]   _zz_6669;
  wire       [15:0]   _zz_6670;
  wire       [15:0]   _zz_6671;
  wire       [15:0]   _zz_6672;
  wire       [15:0]   _zz_6673;
  wire       [15:0]   _zz_6674;
  wire       [15:0]   _zz_6675;
  wire       [15:0]   _zz_6676;
  wire       [15:0]   _zz_6677;
  wire       [15:0]   _zz_6678;
  wire       [15:0]   _zz_6679;
  wire       [15:0]   _zz_6680;
  wire       [15:0]   _zz_6681;
  wire       [15:0]   _zz_6682;
  wire       [15:0]   _zz_6683;
  wire       [15:0]   _zz_6684;
  wire       [15:0]   _zz_6685;
  wire       [15:0]   _zz_6686;
  wire       [15:0]   _zz_6687;
  wire       [15:0]   _zz_6688;
  wire       [15:0]   _zz_6689;
  wire       [15:0]   _zz_6690;
  wire       [15:0]   _zz_6691;
  wire       [15:0]   _zz_6692;
  wire       [15:0]   _zz_6693;
  wire       [15:0]   _zz_6694;
  wire       [15:0]   _zz_6695;
  wire       [15:0]   _zz_6696;
  wire       [15:0]   _zz_6697;
  wire       [15:0]   _zz_6698;
  wire       [15:0]   _zz_6699;
  wire       [15:0]   _zz_6700;
  wire       [15:0]   _zz_6701;
  wire       [15:0]   _zz_6702;
  wire       [15:0]   _zz_6703;
  wire       [15:0]   _zz_6704;
  wire       [15:0]   _zz_6705;
  wire       [15:0]   _zz_6706;
  wire       [15:0]   _zz_6707;
  wire       [15:0]   _zz_6708;
  wire       [15:0]   _zz_6709;
  wire       [15:0]   _zz_6710;
  wire       [15:0]   _zz_6711;
  wire       [15:0]   _zz_6712;
  wire       [15:0]   _zz_6713;
  wire       [15:0]   _zz_6714;
  wire       [15:0]   _zz_6715;
  wire       [15:0]   _zz_6716;
  wire       [15:0]   _zz_6717;
  wire       [15:0]   _zz_6718;
  wire       [15:0]   _zz_6719;
  wire       [15:0]   _zz_6720;
  wire       [15:0]   _zz_6721;
  wire       [15:0]   _zz_6722;
  wire       [15:0]   _zz_6723;
  wire       [15:0]   _zz_6724;
  wire       [15:0]   _zz_6725;
  wire       [15:0]   _zz_6726;
  wire       [15:0]   _zz_6727;
  wire       [15:0]   _zz_6728;
  wire       [15:0]   _zz_6729;
  wire       [15:0]   _zz_6730;
  wire       [15:0]   _zz_6731;
  wire       [15:0]   _zz_6732;
  wire       [15:0]   _zz_6733;
  wire       [15:0]   _zz_6734;
  wire       [15:0]   _zz_6735;
  wire       [15:0]   _zz_6736;
  wire       [15:0]   _zz_6737;
  wire       [15:0]   _zz_6738;
  wire       [15:0]   _zz_6739;
  wire       [15:0]   _zz_6740;
  wire       [15:0]   _zz_6741;
  wire       [15:0]   _zz_6742;
  wire       [15:0]   _zz_6743;
  wire       [15:0]   _zz_6744;
  wire       [15:0]   _zz_6745;
  wire       [15:0]   _zz_6746;
  wire       [15:0]   _zz_6747;
  wire       [15:0]   _zz_6748;
  wire       [15:0]   _zz_6749;
  wire       [15:0]   _zz_6750;
  wire       [15:0]   _zz_6751;
  wire       [15:0]   _zz_6752;
  wire       [15:0]   _zz_6753;
  wire       [15:0]   _zz_6754;
  wire       [15:0]   _zz_6755;
  wire       [15:0]   _zz_6756;
  wire       [15:0]   _zz_6757;
  wire       [15:0]   _zz_6758;
  wire       [15:0]   _zz_6759;
  wire       [15:0]   _zz_6760;
  wire       [15:0]   _zz_6761;
  wire       [15:0]   _zz_6762;
  wire       [15:0]   _zz_6763;
  wire       [15:0]   _zz_6764;
  wire       [15:0]   _zz_6765;
  wire       [15:0]   _zz_6766;
  wire       [15:0]   _zz_6767;
  wire       [15:0]   _zz_6768;
  wire       [15:0]   _zz_6769;
  wire       [15:0]   _zz_6770;
  wire       [15:0]   _zz_6771;
  wire       [15:0]   _zz_6772;
  wire       [15:0]   _zz_6773;
  wire       [15:0]   _zz_6774;
  wire       [15:0]   _zz_6775;
  wire       [15:0]   _zz_6776;
  wire       [15:0]   _zz_6777;
  wire       [15:0]   _zz_6778;
  wire       [15:0]   _zz_6779;
  wire       [15:0]   _zz_6780;
  wire       [15:0]   _zz_6781;
  wire       [15:0]   _zz_6782;
  wire       [15:0]   _zz_6783;
  wire       [15:0]   _zz_6784;
  wire       [15:0]   _zz_6785;
  wire       [15:0]   _zz_6786;
  wire       [15:0]   _zz_6787;
  wire       [15:0]   _zz_6788;
  wire       [15:0]   _zz_6789;
  wire       [15:0]   _zz_6790;
  wire       [15:0]   _zz_6791;
  wire       [15:0]   _zz_6792;
  wire       [15:0]   _zz_6793;
  wire       [15:0]   _zz_6794;
  wire       [15:0]   _zz_6795;
  wire       [15:0]   _zz_6796;
  wire       [15:0]   _zz_6797;
  wire       [15:0]   _zz_6798;
  wire       [15:0]   _zz_6799;
  wire       [15:0]   _zz_6800;
  wire       [15:0]   _zz_6801;
  wire       [15:0]   _zz_6802;
  wire       [15:0]   _zz_6803;
  wire       [15:0]   _zz_6804;
  wire       [15:0]   _zz_6805;
  wire       [15:0]   _zz_6806;
  wire       [15:0]   _zz_6807;
  wire       [15:0]   _zz_6808;
  wire       [15:0]   _zz_6809;
  wire       [15:0]   _zz_6810;
  wire       [15:0]   _zz_6811;
  wire       [15:0]   _zz_6812;
  wire       [15:0]   _zz_6813;
  wire       [15:0]   _zz_6814;
  wire       [15:0]   _zz_6815;
  wire       [15:0]   _zz_6816;
  wire       [15:0]   _zz_6817;
  wire       [15:0]   _zz_6818;
  wire       [15:0]   _zz_6819;
  wire       [15:0]   _zz_6820;
  wire       [15:0]   _zz_6821;
  wire       [15:0]   _zz_6822;
  wire       [15:0]   _zz_6823;
  wire       [15:0]   _zz_6824;
  wire       [15:0]   _zz_6825;
  wire       [15:0]   _zz_6826;
  wire       [15:0]   _zz_6827;
  wire       [15:0]   _zz_6828;
  wire       [15:0]   _zz_6829;
  wire       [15:0]   _zz_6830;
  wire       [15:0]   _zz_6831;
  wire       [15:0]   _zz_6832;
  wire       [15:0]   _zz_6833;
  wire       [15:0]   _zz_6834;
  wire       [15:0]   _zz_6835;
  wire       [15:0]   _zz_6836;
  wire       [15:0]   _zz_6837;
  wire       [15:0]   _zz_6838;
  wire       [15:0]   _zz_6839;
  wire       [15:0]   _zz_6840;
  wire       [15:0]   _zz_6841;
  wire       [15:0]   _zz_6842;
  wire       [15:0]   _zz_6843;
  wire       [15:0]   _zz_6844;
  wire       [15:0]   _zz_6845;
  wire       [15:0]   _zz_6846;
  wire       [15:0]   _zz_6847;
  wire       [15:0]   _zz_6848;
  wire       [15:0]   _zz_6849;
  wire       [15:0]   _zz_6850;
  wire       [15:0]   _zz_6851;
  wire       [15:0]   _zz_6852;
  wire       [15:0]   _zz_6853;
  wire       [15:0]   _zz_6854;
  wire       [15:0]   _zz_6855;
  wire       [15:0]   _zz_6856;
  wire       [15:0]   _zz_6857;
  wire       [15:0]   _zz_6858;
  wire       [15:0]   _zz_6859;
  wire       [15:0]   _zz_6860;
  wire       [15:0]   _zz_6861;
  wire       [15:0]   _zz_6862;
  wire       [15:0]   _zz_6863;
  wire       [15:0]   _zz_6864;
  wire       [15:0]   _zz_6865;
  wire       [15:0]   _zz_6866;
  wire       [15:0]   _zz_6867;
  wire       [15:0]   _zz_6868;
  wire       [15:0]   _zz_6869;
  wire       [15:0]   _zz_6870;
  wire       [15:0]   _zz_6871;
  wire       [15:0]   _zz_6872;
  wire       [15:0]   _zz_6873;
  wire       [15:0]   _zz_6874;
  wire       [15:0]   _zz_6875;
  wire       [15:0]   _zz_6876;
  wire       [15:0]   _zz_6877;
  wire       [15:0]   _zz_6878;
  wire       [15:0]   _zz_6879;
  wire       [15:0]   _zz_6880;
  wire       [15:0]   _zz_6881;
  wire       [15:0]   _zz_6882;
  wire       [15:0]   _zz_6883;
  wire       [15:0]   _zz_6884;
  wire       [15:0]   _zz_6885;
  wire       [15:0]   _zz_6886;
  wire       [15:0]   _zz_6887;
  wire       [15:0]   _zz_6888;
  wire       [15:0]   _zz_6889;
  wire       [15:0]   _zz_6890;
  wire       [15:0]   _zz_6891;
  wire       [15:0]   _zz_6892;
  wire       [15:0]   _zz_6893;
  wire       [15:0]   _zz_6894;
  wire       [15:0]   _zz_6895;
  wire       [15:0]   _zz_6896;
  wire       [15:0]   _zz_6897;
  wire       [15:0]   _zz_6898;
  wire       [15:0]   _zz_6899;
  wire       [15:0]   _zz_6900;
  wire       [15:0]   _zz_6901;
  wire       [15:0]   _zz_6902;
  wire       [15:0]   _zz_6903;
  wire       [15:0]   _zz_6904;
  wire       [15:0]   _zz_6905;
  wire       [15:0]   _zz_6906;
  wire       [15:0]   _zz_6907;
  wire       [15:0]   _zz_6908;
  wire       [15:0]   _zz_6909;
  wire       [15:0]   _zz_6910;
  wire       [15:0]   _zz_6911;
  wire       [15:0]   _zz_6912;
  wire       [15:0]   _zz_6913;
  wire       [15:0]   _zz_6914;
  wire       [15:0]   _zz_6915;
  wire       [15:0]   _zz_6916;
  wire       [15:0]   _zz_6917;
  wire       [15:0]   _zz_6918;
  wire       [15:0]   _zz_6919;
  wire       [15:0]   _zz_6920;
  wire       [15:0]   _zz_6921;
  wire       [15:0]   _zz_6922;
  wire       [15:0]   _zz_6923;
  wire       [15:0]   _zz_6924;
  wire       [15:0]   _zz_6925;
  wire       [15:0]   _zz_6926;
  wire       [15:0]   _zz_6927;
  wire       [15:0]   _zz_6928;
  wire       [15:0]   _zz_6929;
  wire       [15:0]   _zz_6930;
  wire       [15:0]   _zz_6931;
  wire       [15:0]   _zz_6932;
  wire       [15:0]   _zz_6933;
  wire       [15:0]   _zz_6934;
  wire       [15:0]   _zz_6935;
  wire       [15:0]   _zz_6936;
  wire       [15:0]   _zz_6937;
  wire       [15:0]   _zz_6938;
  wire       [15:0]   _zz_6939;
  wire       [15:0]   _zz_6940;
  wire       [15:0]   _zz_6941;
  wire       [15:0]   _zz_6942;
  wire       [15:0]   _zz_6943;
  wire       [15:0]   _zz_6944;
  wire       [15:0]   _zz_6945;
  wire       [15:0]   _zz_6946;
  wire       [15:0]   _zz_6947;
  wire       [15:0]   _zz_6948;
  wire       [15:0]   _zz_6949;
  wire       [15:0]   _zz_6950;
  wire       [15:0]   _zz_6951;
  wire       [15:0]   _zz_6952;
  wire       [15:0]   _zz_6953;
  wire       [15:0]   _zz_6954;
  wire       [15:0]   _zz_6955;
  wire       [15:0]   _zz_6956;
  wire       [15:0]   _zz_6957;
  wire       [15:0]   _zz_6958;
  wire       [15:0]   _zz_6959;
  wire       [15:0]   _zz_6960;
  wire       [15:0]   _zz_6961;
  wire       [15:0]   _zz_6962;
  wire       [15:0]   _zz_6963;
  wire       [15:0]   _zz_6964;
  wire       [15:0]   _zz_6965;
  wire       [15:0]   _zz_6966;
  wire       [15:0]   _zz_6967;
  wire       [15:0]   _zz_6968;
  wire       [15:0]   _zz_6969;
  wire       [15:0]   _zz_6970;
  wire       [15:0]   _zz_6971;
  wire       [15:0]   _zz_6972;
  wire       [15:0]   _zz_6973;
  wire       [15:0]   _zz_6974;
  wire       [15:0]   _zz_6975;
  wire       [15:0]   _zz_6976;
  wire       [15:0]   _zz_6977;
  wire       [15:0]   _zz_6978;
  wire       [15:0]   _zz_6979;
  wire       [15:0]   _zz_6980;
  wire       [15:0]   _zz_6981;
  wire       [15:0]   _zz_6982;
  wire       [15:0]   _zz_6983;
  wire       [15:0]   _zz_6984;
  wire       [15:0]   _zz_6985;
  wire       [15:0]   _zz_6986;
  wire       [15:0]   _zz_6987;
  wire       [15:0]   _zz_6988;
  wire       [15:0]   _zz_6989;
  wire       [15:0]   _zz_6990;
  wire       [15:0]   _zz_6991;
  wire       [15:0]   _zz_6992;
  wire       [15:0]   _zz_6993;
  wire       [15:0]   _zz_6994;
  wire       [15:0]   _zz_6995;
  wire       [15:0]   _zz_6996;
  wire       [15:0]   _zz_6997;
  wire       [15:0]   _zz_6998;
  wire       [15:0]   _zz_6999;
  wire       [15:0]   _zz_7000;
  wire       [15:0]   _zz_7001;
  wire       [15:0]   _zz_7002;
  wire       [15:0]   _zz_7003;
  wire       [15:0]   _zz_7004;
  wire       [15:0]   _zz_7005;
  wire       [15:0]   _zz_7006;
  wire       [15:0]   _zz_7007;
  wire       [15:0]   _zz_7008;
  wire       [15:0]   _zz_7009;
  wire       [15:0]   _zz_7010;
  wire       [15:0]   _zz_7011;
  wire       [15:0]   _zz_7012;
  wire       [15:0]   _zz_7013;
  wire       [15:0]   _zz_7014;
  wire       [15:0]   _zz_7015;
  wire       [15:0]   _zz_7016;
  wire       [15:0]   _zz_7017;
  wire       [15:0]   _zz_7018;
  wire       [15:0]   _zz_7019;
  wire       [15:0]   _zz_7020;
  wire       [15:0]   _zz_7021;
  wire       [15:0]   _zz_7022;
  wire       [15:0]   _zz_7023;
  wire       [15:0]   _zz_7024;
  wire       [15:0]   _zz_7025;
  wire       [15:0]   _zz_7026;
  wire       [15:0]   _zz_7027;
  wire       [15:0]   _zz_7028;
  wire       [15:0]   _zz_7029;
  wire       [15:0]   _zz_7030;
  wire       [15:0]   _zz_7031;
  wire       [15:0]   _zz_7032;
  wire       [15:0]   _zz_7033;
  wire       [15:0]   _zz_7034;
  wire       [15:0]   _zz_7035;
  wire       [15:0]   _zz_7036;
  wire       [15:0]   _zz_7037;
  wire       [15:0]   _zz_7038;
  wire       [15:0]   _zz_7039;
  wire       [15:0]   _zz_7040;
  wire       [15:0]   _zz_7041;
  wire       [15:0]   _zz_7042;
  wire       [15:0]   _zz_7043;
  wire       [15:0]   _zz_7044;
  wire       [15:0]   _zz_7045;
  wire       [15:0]   _zz_7046;
  wire       [15:0]   _zz_7047;
  wire       [15:0]   _zz_7048;
  wire       [15:0]   _zz_7049;
  wire       [15:0]   _zz_7050;
  wire       [15:0]   _zz_7051;
  wire       [15:0]   _zz_7052;
  wire       [15:0]   _zz_7053;
  wire       [15:0]   _zz_7054;
  wire       [15:0]   _zz_7055;
  wire       [15:0]   _zz_7056;
  wire       [15:0]   _zz_7057;
  wire       [15:0]   _zz_7058;
  wire       [15:0]   _zz_7059;
  wire       [15:0]   _zz_7060;
  wire       [15:0]   _zz_7061;
  wire       [15:0]   _zz_7062;
  wire       [15:0]   _zz_7063;
  wire       [15:0]   _zz_7064;
  wire       [15:0]   _zz_7065;
  wire       [15:0]   _zz_7066;
  wire       [15:0]   _zz_7067;
  wire       [15:0]   _zz_7068;
  wire       [15:0]   _zz_7069;
  wire       [15:0]   _zz_7070;
  wire       [15:0]   _zz_7071;
  wire       [15:0]   _zz_7072;
  wire       [15:0]   _zz_7073;
  wire       [15:0]   _zz_7074;
  wire       [15:0]   _zz_7075;
  wire       [15:0]   _zz_7076;
  wire       [15:0]   _zz_7077;
  wire       [15:0]   _zz_7078;
  wire       [15:0]   _zz_7079;
  wire       [15:0]   _zz_7080;
  wire       [15:0]   _zz_7081;
  wire       [15:0]   _zz_7082;
  wire       [15:0]   _zz_7083;
  wire       [15:0]   _zz_7084;
  wire       [15:0]   _zz_7085;
  wire       [15:0]   _zz_7086;
  wire       [15:0]   _zz_7087;
  wire       [15:0]   _zz_7088;
  wire       [15:0]   _zz_7089;
  wire       [15:0]   _zz_7090;
  wire       [15:0]   _zz_7091;
  wire       [15:0]   _zz_7092;
  wire       [15:0]   _zz_7093;
  wire       [15:0]   _zz_7094;
  wire       [15:0]   _zz_7095;
  wire       [15:0]   _zz_7096;
  wire       [15:0]   _zz_7097;
  wire       [15:0]   _zz_7098;
  wire       [15:0]   _zz_7099;
  wire       [15:0]   _zz_7100;
  wire       [15:0]   _zz_7101;
  wire       [15:0]   _zz_7102;
  wire       [15:0]   _zz_7103;
  wire       [15:0]   _zz_7104;
  wire       [15:0]   _zz_7105;
  wire       [15:0]   _zz_7106;
  wire       [15:0]   _zz_7107;
  wire       [15:0]   _zz_7108;
  wire       [15:0]   _zz_7109;
  wire       [15:0]   _zz_7110;
  wire       [15:0]   _zz_7111;
  wire       [15:0]   _zz_7112;
  wire       [15:0]   _zz_7113;
  wire       [15:0]   _zz_7114;
  wire       [15:0]   _zz_7115;
  wire       [15:0]   _zz_7116;
  wire       [15:0]   _zz_7117;
  wire       [15:0]   _zz_7118;
  wire       [15:0]   _zz_7119;
  wire       [15:0]   _zz_7120;
  wire       [15:0]   _zz_7121;
  wire       [15:0]   _zz_7122;
  wire       [15:0]   _zz_7123;
  wire       [15:0]   _zz_7124;
  wire       [15:0]   _zz_7125;
  wire       [15:0]   _zz_7126;
  wire       [15:0]   _zz_7127;
  wire       [15:0]   _zz_7128;
  wire       [15:0]   _zz_7129;
  wire       [15:0]   _zz_7130;
  wire       [15:0]   _zz_7131;
  wire       [15:0]   _zz_7132;
  wire       [15:0]   _zz_7133;
  wire       [15:0]   _zz_7134;
  wire       [15:0]   _zz_7135;
  wire       [15:0]   _zz_7136;
  wire       [15:0]   _zz_7137;
  wire       [15:0]   _zz_7138;
  wire       [15:0]   _zz_7139;
  wire       [15:0]   _zz_7140;
  wire       [15:0]   _zz_7141;
  wire       [15:0]   _zz_7142;
  wire       [15:0]   _zz_7143;
  wire       [15:0]   _zz_7144;
  wire       [15:0]   _zz_7145;
  wire       [15:0]   _zz_7146;
  wire       [15:0]   _zz_7147;
  wire       [15:0]   _zz_7148;
  wire       [15:0]   _zz_7149;
  wire       [15:0]   _zz_7150;
  wire       [15:0]   _zz_7151;
  wire       [15:0]   _zz_7152;
  wire       [15:0]   _zz_7153;
  wire       [15:0]   _zz_7154;
  wire       [15:0]   _zz_7155;
  wire       [15:0]   _zz_7156;
  wire       [15:0]   _zz_7157;
  wire       [15:0]   _zz_7158;
  wire       [15:0]   _zz_7159;
  wire       [15:0]   _zz_7160;
  wire       [15:0]   _zz_7161;
  wire       [15:0]   _zz_7162;
  wire       [15:0]   _zz_7163;
  wire       [15:0]   _zz_7164;
  wire       [15:0]   _zz_7165;
  wire       [15:0]   _zz_7166;
  wire       [15:0]   _zz_7167;
  wire       [15:0]   _zz_7168;
  wire       [15:0]   _zz_7169;
  wire       [15:0]   _zz_7170;
  wire       [15:0]   _zz_7171;
  wire       [15:0]   _zz_7172;
  wire       [15:0]   _zz_7173;
  wire       [15:0]   _zz_7174;
  wire       [15:0]   _zz_7175;
  wire       [15:0]   _zz_7176;
  wire       [15:0]   _zz_7177;
  wire       [15:0]   _zz_7178;
  wire       [15:0]   _zz_7179;
  wire       [15:0]   _zz_7180;
  wire       [15:0]   _zz_7181;
  wire       [15:0]   _zz_7182;
  wire       [15:0]   _zz_7183;
  wire       [15:0]   _zz_7184;
  wire       [15:0]   _zz_7185;
  wire       [15:0]   _zz_7186;
  wire       [15:0]   _zz_7187;
  wire       [15:0]   _zz_7188;
  wire       [15:0]   _zz_7189;
  wire       [15:0]   _zz_7190;
  wire       [15:0]   _zz_7191;
  wire       [15:0]   _zz_7192;
  wire       [15:0]   _zz_7193;
  wire       [15:0]   _zz_7194;
  wire       [15:0]   _zz_7195;
  wire       [15:0]   _zz_7196;
  wire       [15:0]   _zz_7197;
  wire       [15:0]   _zz_7198;
  wire       [15:0]   _zz_7199;
  wire       [15:0]   _zz_7200;
  wire       [15:0]   _zz_7201;
  wire       [15:0]   _zz_7202;
  wire       [15:0]   _zz_7203;
  wire       [15:0]   _zz_7204;
  wire       [15:0]   _zz_7205;
  wire       [15:0]   _zz_7206;
  wire       [15:0]   _zz_7207;
  wire       [15:0]   _zz_7208;
  wire       [15:0]   _zz_7209;
  wire       [15:0]   _zz_7210;
  wire       [15:0]   _zz_7211;
  wire       [15:0]   _zz_7212;
  wire       [15:0]   _zz_7213;
  wire       [15:0]   _zz_7214;
  wire       [15:0]   _zz_7215;
  wire       [15:0]   _zz_7216;
  wire       [15:0]   _zz_7217;
  wire       [15:0]   _zz_7218;
  wire       [15:0]   _zz_7219;
  wire       [15:0]   _zz_7220;
  wire       [15:0]   _zz_7221;
  wire       [15:0]   _zz_7222;
  wire       [15:0]   _zz_7223;
  wire       [15:0]   _zz_7224;
  wire       [15:0]   _zz_7225;
  wire       [15:0]   _zz_7226;
  wire       [15:0]   _zz_7227;
  wire       [15:0]   _zz_7228;
  wire       [15:0]   _zz_7229;
  wire       [15:0]   _zz_7230;
  wire       [15:0]   _zz_7231;
  wire       [15:0]   _zz_7232;
  wire       [15:0]   _zz_7233;
  wire       [15:0]   _zz_7234;
  wire       [15:0]   _zz_7235;
  wire       [15:0]   _zz_7236;
  wire       [15:0]   _zz_7237;
  wire       [15:0]   _zz_7238;
  wire       [15:0]   _zz_7239;
  wire       [15:0]   _zz_7240;
  wire       [15:0]   _zz_7241;
  wire       [15:0]   _zz_7242;
  wire       [15:0]   _zz_7243;
  wire       [15:0]   _zz_7244;
  wire       [15:0]   _zz_7245;
  wire       [15:0]   _zz_7246;
  wire       [15:0]   _zz_7247;
  wire       [15:0]   _zz_7248;
  wire       [15:0]   _zz_7249;
  wire       [15:0]   _zz_7250;
  wire       [15:0]   _zz_7251;
  wire       [15:0]   _zz_7252;
  wire       [15:0]   _zz_7253;
  wire       [15:0]   _zz_7254;
  wire       [15:0]   _zz_7255;
  wire       [15:0]   _zz_7256;
  wire       [15:0]   _zz_7257;
  wire       [15:0]   _zz_7258;
  wire       [15:0]   _zz_7259;
  wire       [15:0]   _zz_7260;
  wire       [15:0]   _zz_7261;
  wire       [15:0]   _zz_7262;
  wire       [15:0]   _zz_7263;
  wire       [15:0]   _zz_7264;
  wire       [15:0]   _zz_7265;
  wire       [15:0]   _zz_7266;
  wire       [15:0]   _zz_7267;
  wire       [15:0]   _zz_7268;
  wire       [15:0]   _zz_7269;
  wire       [15:0]   _zz_7270;
  wire       [15:0]   _zz_7271;
  wire       [15:0]   _zz_7272;
  wire       [15:0]   _zz_7273;
  wire       [15:0]   _zz_7274;
  wire       [15:0]   _zz_7275;
  wire       [15:0]   _zz_7276;
  wire       [15:0]   _zz_7277;
  wire       [15:0]   _zz_7278;
  wire       [15:0]   _zz_7279;
  wire       [15:0]   _zz_7280;
  wire       [15:0]   _zz_7281;
  wire       [15:0]   _zz_7282;
  wire       [15:0]   _zz_7283;
  wire       [15:0]   _zz_7284;
  wire       [15:0]   _zz_7285;
  wire       [15:0]   _zz_7286;
  wire       [15:0]   _zz_7287;
  wire       [15:0]   _zz_7288;
  wire       [15:0]   _zz_7289;
  wire       [15:0]   _zz_7290;
  wire       [15:0]   _zz_7291;
  wire       [15:0]   _zz_7292;
  wire       [15:0]   _zz_7293;
  wire       [15:0]   _zz_7294;
  wire       [15:0]   _zz_7295;
  wire       [15:0]   _zz_7296;
  wire       [15:0]   _zz_7297;
  wire       [15:0]   _zz_7298;
  wire       [15:0]   _zz_7299;
  wire       [15:0]   _zz_7300;
  wire       [15:0]   _zz_7301;
  wire       [15:0]   _zz_7302;
  wire       [15:0]   _zz_7303;
  wire       [15:0]   _zz_7304;
  wire       [15:0]   _zz_7305;
  wire       [15:0]   _zz_7306;
  wire       [15:0]   _zz_7307;
  wire       [15:0]   _zz_7308;
  wire       [15:0]   _zz_7309;
  wire       [15:0]   _zz_7310;
  wire       [15:0]   _zz_7311;
  wire       [15:0]   _zz_7312;
  wire       [15:0]   _zz_7313;
  wire       [15:0]   _zz_7314;
  wire       [15:0]   _zz_7315;
  wire       [15:0]   _zz_7316;
  wire       [15:0]   _zz_7317;
  wire       [15:0]   _zz_7318;
  wire       [15:0]   _zz_7319;
  wire       [15:0]   _zz_7320;
  wire       [15:0]   _zz_7321;
  wire       [15:0]   _zz_7322;
  wire       [15:0]   _zz_7323;
  wire       [15:0]   _zz_7324;
  wire       [15:0]   _zz_7325;
  wire       [15:0]   _zz_7326;
  wire       [15:0]   _zz_7327;
  wire       [15:0]   _zz_7328;
  wire       [15:0]   _zz_7329;
  wire       [15:0]   _zz_7330;
  wire       [15:0]   _zz_7331;
  wire       [15:0]   _zz_7332;
  wire       [15:0]   _zz_7333;
  wire       [15:0]   _zz_7334;
  wire       [15:0]   _zz_7335;
  wire       [15:0]   _zz_7336;
  wire       [15:0]   _zz_7337;
  wire       [15:0]   _zz_7338;
  wire       [15:0]   _zz_7339;
  wire       [15:0]   _zz_7340;
  wire       [15:0]   _zz_7341;
  wire       [15:0]   _zz_7342;
  wire       [15:0]   _zz_7343;
  wire       [15:0]   _zz_7344;
  wire       [15:0]   _zz_7345;
  wire       [15:0]   _zz_7346;
  wire       [15:0]   _zz_7347;
  wire       [15:0]   _zz_7348;
  wire       [15:0]   _zz_7349;
  wire       [15:0]   _zz_7350;
  wire       [15:0]   _zz_7351;
  wire       [15:0]   _zz_7352;
  wire       [15:0]   _zz_7353;
  wire       [15:0]   _zz_7354;
  wire       [15:0]   _zz_7355;
  wire       [15:0]   _zz_7356;
  wire       [15:0]   _zz_7357;
  wire       [15:0]   _zz_7358;
  wire       [15:0]   _zz_7359;
  wire       [15:0]   _zz_7360;
  wire       [15:0]   _zz_7361;
  wire       [15:0]   _zz_7362;
  wire       [15:0]   _zz_7363;
  wire       [15:0]   _zz_7364;
  wire       [15:0]   _zz_7365;
  wire       [15:0]   _zz_7366;
  wire       [15:0]   _zz_7367;
  wire       [15:0]   _zz_7368;
  wire       [15:0]   _zz_7369;
  wire       [15:0]   _zz_7370;
  wire       [15:0]   _zz_7371;
  wire       [15:0]   _zz_7372;
  wire       [15:0]   _zz_7373;
  wire       [15:0]   _zz_7374;
  wire       [15:0]   _zz_7375;
  wire       [15:0]   _zz_7376;
  wire       [15:0]   _zz_7377;
  wire       [15:0]   _zz_7378;
  wire       [15:0]   _zz_7379;
  wire       [15:0]   _zz_7380;
  wire       [15:0]   _zz_7381;
  wire       [15:0]   _zz_7382;
  wire       [15:0]   _zz_7383;
  wire       [15:0]   _zz_7384;
  wire       [15:0]   _zz_7385;
  wire       [15:0]   _zz_7386;
  wire       [15:0]   _zz_7387;
  wire       [15:0]   _zz_7388;
  wire       [15:0]   _zz_7389;
  wire       [15:0]   _zz_7390;
  wire       [15:0]   _zz_7391;
  wire       [15:0]   _zz_7392;
  wire       [15:0]   _zz_7393;
  wire       [15:0]   _zz_7394;
  wire       [15:0]   _zz_7395;
  wire       [15:0]   _zz_7396;
  wire       [15:0]   _zz_7397;
  wire       [15:0]   _zz_7398;
  wire       [15:0]   _zz_7399;
  wire       [15:0]   _zz_7400;
  wire       [15:0]   _zz_7401;
  wire       [15:0]   _zz_7402;
  wire       [15:0]   _zz_7403;
  wire       [15:0]   _zz_7404;
  wire       [15:0]   _zz_7405;
  wire       [15:0]   _zz_7406;
  wire       [15:0]   _zz_7407;
  wire       [15:0]   _zz_7408;
  wire       [15:0]   _zz_7409;
  wire       [15:0]   _zz_7410;
  wire       [15:0]   _zz_7411;
  wire       [15:0]   _zz_7412;
  wire       [15:0]   _zz_7413;
  wire       [15:0]   _zz_7414;
  wire       [15:0]   _zz_7415;
  wire       [15:0]   _zz_7416;
  wire       [15:0]   _zz_7417;
  wire       [15:0]   _zz_7418;
  wire       [15:0]   _zz_7419;
  wire       [15:0]   _zz_7420;
  wire       [15:0]   _zz_7421;
  wire       [15:0]   _zz_7422;
  wire       [15:0]   _zz_7423;
  wire       [15:0]   _zz_7424;
  wire       [15:0]   _zz_7425;
  wire       [15:0]   _zz_7426;
  wire       [15:0]   _zz_7427;
  wire       [15:0]   _zz_7428;
  wire       [15:0]   _zz_7429;
  wire       [15:0]   _zz_7430;
  wire       [15:0]   _zz_7431;
  wire       [15:0]   _zz_7432;
  wire       [15:0]   _zz_7433;
  wire       [15:0]   _zz_7434;
  wire       [15:0]   _zz_7435;
  wire       [15:0]   _zz_7436;
  wire       [15:0]   _zz_7437;
  wire       [15:0]   _zz_7438;
  wire       [15:0]   _zz_7439;
  wire       [15:0]   _zz_7440;
  wire       [15:0]   _zz_7441;
  wire       [15:0]   _zz_7442;
  wire       [15:0]   _zz_7443;
  wire       [15:0]   _zz_7444;
  wire       [15:0]   _zz_7445;
  wire       [15:0]   _zz_7446;
  wire       [15:0]   _zz_7447;
  wire       [15:0]   _zz_7448;
  wire       [15:0]   _zz_7449;
  wire       [15:0]   _zz_7450;
  wire       [15:0]   _zz_7451;
  wire       [15:0]   _zz_7452;
  wire       [15:0]   _zz_7453;
  wire       [15:0]   _zz_7454;
  wire       [15:0]   _zz_7455;
  wire       [15:0]   _zz_7456;
  wire       [15:0]   _zz_7457;
  wire       [15:0]   _zz_7458;
  wire       [15:0]   _zz_7459;
  wire       [15:0]   _zz_7460;
  wire       [15:0]   _zz_7461;
  wire       [15:0]   _zz_7462;
  wire       [15:0]   _zz_7463;
  wire       [15:0]   _zz_7464;
  wire       [15:0]   _zz_7465;
  wire       [15:0]   _zz_7466;
  wire       [15:0]   _zz_7467;
  wire       [15:0]   _zz_7468;
  wire       [15:0]   _zz_7469;
  wire       [15:0]   _zz_7470;
  wire       [15:0]   _zz_7471;
  wire       [15:0]   _zz_7472;
  wire       [15:0]   _zz_7473;
  wire       [15:0]   _zz_7474;
  wire       [15:0]   _zz_7475;
  wire       [15:0]   _zz_7476;
  wire       [15:0]   _zz_7477;
  wire       [15:0]   _zz_7478;
  wire       [15:0]   _zz_7479;
  wire       [15:0]   _zz_7480;
  wire       [15:0]   _zz_7481;
  wire       [15:0]   _zz_7482;
  wire       [15:0]   _zz_7483;
  wire       [15:0]   _zz_7484;
  wire       [15:0]   _zz_7485;
  wire       [15:0]   _zz_7486;
  wire       [15:0]   _zz_7487;
  wire       [15:0]   _zz_7488;
  wire       [15:0]   _zz_7489;
  wire       [15:0]   _zz_7490;
  wire       [15:0]   _zz_7491;
  wire       [15:0]   _zz_7492;
  wire       [15:0]   _zz_7493;
  wire       [15:0]   _zz_7494;
  wire       [15:0]   _zz_7495;
  wire       [15:0]   _zz_7496;
  wire       [15:0]   _zz_7497;
  wire       [15:0]   _zz_7498;
  wire       [15:0]   _zz_7499;
  wire       [15:0]   _zz_7500;
  wire       [15:0]   _zz_7501;
  wire       [15:0]   _zz_7502;
  wire       [15:0]   _zz_7503;
  wire       [15:0]   _zz_7504;
  wire       [15:0]   _zz_7505;
  wire       [15:0]   _zz_7506;
  wire       [15:0]   _zz_7507;
  wire       [15:0]   _zz_7508;
  wire       [15:0]   _zz_7509;
  wire       [15:0]   _zz_7510;
  wire       [15:0]   _zz_7511;
  wire       [15:0]   _zz_7512;
  wire       [15:0]   _zz_7513;
  wire       [15:0]   _zz_7514;
  wire       [15:0]   _zz_7515;
  wire       [15:0]   _zz_7516;
  wire       [15:0]   _zz_7517;
  wire       [15:0]   _zz_7518;
  wire       [15:0]   _zz_7519;
  wire       [15:0]   _zz_7520;
  wire       [15:0]   _zz_7521;
  wire       [15:0]   _zz_7522;
  wire       [15:0]   _zz_7523;
  wire       [15:0]   _zz_7524;
  wire       [15:0]   _zz_7525;
  wire       [15:0]   _zz_7526;
  wire       [15:0]   _zz_7527;
  wire       [15:0]   _zz_7528;
  wire       [15:0]   _zz_7529;
  wire       [15:0]   _zz_7530;
  wire       [15:0]   _zz_7531;
  wire       [15:0]   _zz_7532;
  wire       [15:0]   _zz_7533;
  wire       [15:0]   _zz_7534;
  wire       [15:0]   _zz_7535;
  wire       [15:0]   _zz_7536;
  wire       [15:0]   _zz_7537;
  wire       [15:0]   _zz_7538;
  wire       [15:0]   _zz_7539;
  wire       [15:0]   _zz_7540;
  wire       [15:0]   _zz_7541;
  wire       [15:0]   _zz_7542;
  wire       [15:0]   _zz_7543;
  wire       [15:0]   _zz_7544;
  wire       [15:0]   _zz_7545;
  wire       [15:0]   _zz_7546;
  wire       [15:0]   _zz_7547;
  wire       [15:0]   _zz_7548;
  wire       [15:0]   _zz_7549;
  wire       [15:0]   _zz_7550;
  wire       [15:0]   _zz_7551;
  wire       [15:0]   _zz_7552;
  wire       [15:0]   _zz_7553;
  wire       [15:0]   _zz_7554;
  wire       [15:0]   _zz_7555;
  wire       [15:0]   _zz_7556;
  wire       [15:0]   _zz_7557;
  wire       [15:0]   _zz_7558;
  wire       [15:0]   _zz_7559;
  wire       [15:0]   _zz_7560;
  wire       [15:0]   _zz_7561;
  wire       [15:0]   _zz_7562;
  wire       [15:0]   _zz_7563;
  wire       [15:0]   _zz_7564;
  wire       [15:0]   _zz_7565;
  wire       [15:0]   _zz_7566;
  wire       [15:0]   _zz_7567;
  wire       [15:0]   _zz_7568;
  wire       [15:0]   _zz_7569;
  wire       [15:0]   _zz_7570;
  wire       [15:0]   _zz_7571;
  wire       [15:0]   _zz_7572;
  wire       [15:0]   _zz_7573;
  wire       [15:0]   _zz_7574;
  wire       [15:0]   _zz_7575;
  wire       [15:0]   _zz_7576;
  wire       [15:0]   _zz_7577;
  wire       [15:0]   _zz_7578;
  wire       [15:0]   _zz_7579;
  wire       [15:0]   _zz_7580;
  wire       [15:0]   _zz_7581;
  wire       [15:0]   _zz_7582;
  wire       [15:0]   _zz_7583;
  wire       [15:0]   _zz_7584;
  wire       [15:0]   _zz_7585;
  wire       [15:0]   _zz_7586;
  wire       [15:0]   _zz_7587;
  wire       [15:0]   _zz_7588;
  wire       [15:0]   _zz_7589;
  wire       [15:0]   _zz_7590;
  wire       [15:0]   _zz_7591;
  wire       [15:0]   _zz_7592;
  wire       [15:0]   _zz_7593;
  wire       [15:0]   _zz_7594;
  wire       [15:0]   _zz_7595;
  wire       [15:0]   _zz_7596;
  wire       [15:0]   _zz_7597;
  wire       [15:0]   _zz_7598;
  wire       [15:0]   _zz_7599;
  wire       [15:0]   _zz_7600;
  wire       [15:0]   _zz_7601;
  wire       [15:0]   _zz_7602;
  wire       [15:0]   _zz_7603;
  wire       [15:0]   _zz_7604;
  wire       [15:0]   _zz_7605;
  wire       [15:0]   _zz_7606;
  wire       [15:0]   _zz_7607;
  wire       [15:0]   _zz_7608;
  wire       [15:0]   _zz_7609;
  wire       [15:0]   _zz_7610;
  wire       [15:0]   _zz_7611;
  wire       [15:0]   _zz_7612;
  wire       [15:0]   _zz_7613;
  wire       [15:0]   _zz_7614;
  wire       [15:0]   _zz_7615;
  wire       [15:0]   _zz_7616;
  wire       [15:0]   _zz_7617;
  wire       [15:0]   _zz_7618;
  wire       [15:0]   _zz_7619;
  wire       [15:0]   _zz_7620;
  wire       [15:0]   _zz_7621;
  wire       [15:0]   _zz_7622;
  wire       [15:0]   _zz_7623;
  wire       [15:0]   _zz_7624;
  wire       [15:0]   _zz_7625;
  wire       [15:0]   _zz_7626;
  wire       [15:0]   _zz_7627;
  wire       [15:0]   _zz_7628;
  wire       [15:0]   _zz_7629;
  wire       [15:0]   _zz_7630;
  wire       [15:0]   _zz_7631;
  wire       [15:0]   _zz_7632;
  wire       [15:0]   _zz_7633;
  wire       [15:0]   _zz_7634;
  wire       [15:0]   _zz_7635;
  wire       [15:0]   _zz_7636;
  wire       [15:0]   _zz_7637;
  wire       [15:0]   _zz_7638;
  wire       [15:0]   _zz_7639;
  wire       [15:0]   _zz_7640;
  wire       [15:0]   _zz_7641;
  wire       [15:0]   _zz_7642;
  wire       [15:0]   _zz_7643;
  wire       [15:0]   _zz_7644;
  wire       [15:0]   _zz_7645;
  wire       [15:0]   _zz_7646;
  wire       [15:0]   _zz_7647;
  wire       [15:0]   _zz_7648;
  wire       [15:0]   _zz_7649;
  wire       [15:0]   _zz_7650;
  wire       [15:0]   _zz_7651;
  wire       [15:0]   _zz_7652;
  wire       [15:0]   _zz_7653;
  wire       [15:0]   _zz_7654;
  wire       [15:0]   _zz_7655;
  wire       [15:0]   _zz_7656;
  wire       [15:0]   _zz_7657;
  wire       [15:0]   _zz_7658;
  wire       [15:0]   _zz_7659;
  wire       [15:0]   _zz_7660;
  wire       [15:0]   _zz_7661;
  wire       [15:0]   _zz_7662;
  wire       [15:0]   _zz_7663;
  wire       [15:0]   _zz_7664;
  wire       [15:0]   _zz_7665;
  wire       [15:0]   _zz_7666;
  wire       [15:0]   _zz_7667;
  wire       [15:0]   _zz_7668;
  wire       [15:0]   _zz_7669;
  wire       [15:0]   _zz_7670;
  wire       [15:0]   _zz_7671;
  wire       [15:0]   _zz_7672;
  wire       [15:0]   _zz_7673;
  wire       [15:0]   _zz_7674;
  wire       [15:0]   _zz_7675;
  wire       [15:0]   _zz_7676;
  wire       [15:0]   _zz_7677;
  wire       [15:0]   _zz_7678;
  wire       [15:0]   _zz_7679;
  wire       [15:0]   _zz_7680;
  wire       [15:0]   _zz_7681;
  wire       [15:0]   _zz_7682;
  wire       [15:0]   _zz_7683;
  wire       [15:0]   _zz_7684;
  wire       [15:0]   _zz_7685;
  wire       [15:0]   _zz_7686;
  wire       [15:0]   _zz_7687;
  wire       [15:0]   _zz_7688;
  wire       [15:0]   _zz_7689;
  wire       [15:0]   _zz_7690;
  wire       [15:0]   _zz_7691;
  wire       [15:0]   _zz_7692;
  wire       [15:0]   _zz_7693;
  wire       [15:0]   _zz_7694;
  wire       [15:0]   _zz_7695;
  wire       [15:0]   _zz_7696;
  wire       [15:0]   _zz_7697;
  wire       [15:0]   _zz_7698;
  wire       [15:0]   _zz_7699;
  wire       [15:0]   _zz_7700;
  wire       [15:0]   _zz_7701;
  wire       [15:0]   _zz_7702;
  wire       [15:0]   _zz_7703;
  wire       [15:0]   _zz_7704;
  wire       [15:0]   _zz_7705;
  wire       [15:0]   _zz_7706;
  wire       [15:0]   _zz_7707;
  wire       [15:0]   _zz_7708;
  wire       [15:0]   _zz_7709;
  wire       [15:0]   _zz_7710;
  wire       [15:0]   _zz_7711;
  wire       [15:0]   _zz_7712;
  wire       [15:0]   _zz_7713;
  wire       [15:0]   _zz_7714;
  wire       [15:0]   _zz_7715;
  wire       [15:0]   _zz_7716;
  wire       [15:0]   _zz_7717;
  wire       [15:0]   _zz_7718;
  wire       [15:0]   _zz_7719;
  wire       [15:0]   _zz_7720;
  wire       [15:0]   _zz_7721;
  wire       [15:0]   _zz_7722;
  wire       [15:0]   _zz_7723;
  wire       [15:0]   _zz_7724;
  wire       [15:0]   _zz_7725;
  wire       [15:0]   _zz_7726;
  wire       [15:0]   _zz_7727;
  wire       [15:0]   _zz_7728;
  wire       [15:0]   _zz_7729;
  wire       [15:0]   _zz_7730;
  wire       [15:0]   _zz_7731;
  wire       [15:0]   _zz_7732;
  wire       [15:0]   _zz_7733;
  wire       [15:0]   _zz_7734;
  wire       [15:0]   _zz_7735;
  wire       [15:0]   _zz_7736;
  wire       [15:0]   _zz_7737;
  wire       [15:0]   _zz_7738;
  wire       [15:0]   _zz_7739;
  wire       [15:0]   _zz_7740;
  wire       [15:0]   _zz_7741;
  wire       [15:0]   _zz_7742;
  wire       [15:0]   _zz_7743;
  wire       [15:0]   _zz_7744;
  wire       [15:0]   _zz_7745;
  wire       [15:0]   _zz_7746;
  wire       [15:0]   _zz_7747;
  wire       [15:0]   _zz_7748;
  wire       [15:0]   _zz_7749;
  wire       [15:0]   _zz_7750;
  wire       [15:0]   _zz_7751;
  wire       [15:0]   _zz_7752;
  wire       [15:0]   _zz_7753;
  wire       [15:0]   _zz_7754;
  wire       [15:0]   _zz_7755;
  wire       [15:0]   _zz_7756;
  wire       [15:0]   _zz_7757;
  wire       [15:0]   _zz_7758;
  wire       [15:0]   _zz_7759;
  wire       [15:0]   _zz_7760;
  wire       [15:0]   _zz_7761;
  wire       [15:0]   _zz_7762;
  wire       [15:0]   _zz_7763;
  wire       [15:0]   _zz_7764;
  wire       [15:0]   _zz_7765;
  wire       [15:0]   _zz_7766;
  wire       [15:0]   _zz_7767;
  wire       [15:0]   _zz_7768;
  wire       [15:0]   _zz_7769;
  wire       [15:0]   _zz_7770;
  wire       [15:0]   _zz_7771;
  wire       [15:0]   _zz_7772;
  wire       [15:0]   _zz_7773;
  wire       [15:0]   _zz_7774;
  wire       [15:0]   _zz_7775;
  wire       [15:0]   _zz_7776;
  wire       [15:0]   _zz_7777;
  wire       [15:0]   _zz_7778;
  wire       [15:0]   _zz_7779;
  wire       [15:0]   _zz_7780;
  wire       [15:0]   _zz_7781;
  wire       [15:0]   _zz_7782;
  wire       [15:0]   _zz_7783;
  wire       [15:0]   _zz_7784;
  wire       [15:0]   _zz_7785;
  wire       [15:0]   _zz_7786;
  wire       [15:0]   _zz_7787;
  wire       [15:0]   _zz_7788;
  wire       [15:0]   _zz_7789;
  wire       [15:0]   _zz_7790;
  wire       [15:0]   _zz_7791;
  wire       [15:0]   _zz_7792;
  wire       [15:0]   _zz_7793;
  wire       [15:0]   _zz_7794;
  wire       [15:0]   _zz_7795;
  wire       [15:0]   _zz_7796;
  wire       [15:0]   _zz_7797;
  wire       [15:0]   _zz_7798;
  wire       [15:0]   _zz_7799;
  wire       [15:0]   _zz_7800;
  wire       [15:0]   _zz_7801;
  wire       [15:0]   _zz_7802;
  wire       [15:0]   _zz_7803;
  wire       [15:0]   _zz_7804;
  wire       [15:0]   _zz_7805;
  wire       [15:0]   _zz_7806;
  wire       [15:0]   _zz_7807;
  wire       [15:0]   _zz_7808;
  wire       [15:0]   _zz_7809;
  wire       [15:0]   _zz_7810;
  wire       [15:0]   _zz_7811;
  wire       [15:0]   _zz_7812;
  wire       [15:0]   _zz_7813;
  wire       [15:0]   _zz_7814;
  wire       [15:0]   _zz_7815;
  wire       [15:0]   _zz_7816;
  wire       [15:0]   _zz_7817;
  wire       [15:0]   _zz_7818;
  wire       [15:0]   _zz_7819;
  wire       [15:0]   _zz_7820;
  wire       [15:0]   _zz_7821;
  wire       [15:0]   _zz_7822;
  wire       [15:0]   _zz_7823;
  wire       [15:0]   _zz_7824;
  wire       [15:0]   _zz_7825;
  wire       [15:0]   _zz_7826;
  wire       [15:0]   _zz_7827;
  wire       [15:0]   _zz_7828;
  wire       [15:0]   _zz_7829;
  wire       [15:0]   _zz_7830;
  wire       [15:0]   _zz_7831;
  wire       [15:0]   _zz_7832;
  wire       [15:0]   _zz_7833;
  wire       [15:0]   _zz_7834;
  wire       [15:0]   _zz_7835;
  wire       [15:0]   _zz_7836;
  wire       [15:0]   _zz_7837;
  wire       [15:0]   _zz_7838;
  wire       [15:0]   _zz_7839;
  wire       [15:0]   _zz_7840;
  wire       [15:0]   _zz_7841;
  wire       [15:0]   _zz_7842;
  wire       [15:0]   _zz_7843;
  wire       [15:0]   _zz_7844;
  wire       [15:0]   _zz_7845;
  wire       [15:0]   _zz_7846;
  wire       [15:0]   _zz_7847;
  wire       [15:0]   _zz_7848;
  wire       [15:0]   _zz_7849;
  wire       [15:0]   _zz_7850;
  wire       [15:0]   _zz_7851;
  wire       [15:0]   _zz_7852;
  wire       [15:0]   _zz_7853;
  wire       [15:0]   _zz_7854;
  wire       [15:0]   _zz_7855;
  wire       [15:0]   _zz_7856;
  wire       [15:0]   _zz_7857;
  wire       [15:0]   _zz_7858;
  wire       [15:0]   _zz_7859;
  wire       [15:0]   _zz_7860;
  wire       [15:0]   _zz_7861;
  wire       [15:0]   _zz_7862;
  wire       [15:0]   _zz_7863;
  wire       [15:0]   _zz_7864;
  wire       [15:0]   _zz_7865;
  wire       [15:0]   _zz_7866;
  wire       [15:0]   _zz_7867;
  wire       [15:0]   _zz_7868;
  wire       [15:0]   _zz_7869;
  wire       [15:0]   _zz_7870;
  wire       [15:0]   _zz_7871;
  wire       [15:0]   _zz_7872;
  wire       [15:0]   _zz_7873;
  wire       [15:0]   _zz_7874;
  wire       [15:0]   _zz_7875;
  wire       [15:0]   _zz_7876;
  wire       [15:0]   _zz_7877;
  wire       [15:0]   _zz_7878;
  wire       [15:0]   _zz_7879;
  wire       [15:0]   _zz_7880;
  wire       [15:0]   _zz_7881;
  wire       [15:0]   _zz_7882;
  wire       [15:0]   _zz_7883;
  wire       [15:0]   _zz_7884;
  wire       [15:0]   _zz_7885;
  wire       [15:0]   _zz_7886;
  wire       [15:0]   _zz_7887;
  wire       [15:0]   _zz_7888;
  wire       [15:0]   _zz_7889;
  wire       [15:0]   _zz_7890;
  wire       [15:0]   _zz_7891;
  wire       [15:0]   _zz_7892;
  wire       [15:0]   _zz_7893;
  wire       [15:0]   _zz_7894;
  wire       [15:0]   _zz_7895;
  wire       [15:0]   _zz_7896;
  wire       [15:0]   _zz_7897;
  wire       [15:0]   _zz_7898;
  wire       [15:0]   _zz_7899;
  wire       [15:0]   _zz_7900;
  wire       [15:0]   _zz_7901;
  wire       [15:0]   _zz_7902;
  wire       [15:0]   _zz_7903;
  wire       [15:0]   _zz_7904;
  wire       [15:0]   _zz_7905;
  wire       [15:0]   _zz_7906;
  wire       [15:0]   _zz_7907;
  wire       [15:0]   _zz_7908;
  wire       [15:0]   _zz_7909;
  wire       [15:0]   _zz_7910;
  wire       [15:0]   _zz_7911;
  wire       [15:0]   _zz_7912;
  wire       [15:0]   _zz_7913;
  wire       [15:0]   _zz_7914;
  wire       [15:0]   _zz_7915;
  wire       [15:0]   _zz_7916;
  wire       [15:0]   _zz_7917;
  wire       [15:0]   _zz_7918;
  wire       [15:0]   _zz_7919;
  wire       [15:0]   _zz_7920;
  wire       [15:0]   _zz_7921;
  wire       [15:0]   _zz_7922;
  wire       [15:0]   _zz_7923;
  wire       [15:0]   _zz_7924;
  wire       [15:0]   _zz_7925;
  wire       [15:0]   _zz_7926;
  wire       [15:0]   _zz_7927;
  wire       [15:0]   _zz_7928;
  wire       [15:0]   _zz_7929;
  wire       [15:0]   _zz_7930;
  wire       [15:0]   _zz_7931;
  wire       [15:0]   _zz_7932;
  wire       [15:0]   _zz_7933;
  wire       [15:0]   _zz_7934;
  wire       [15:0]   _zz_7935;
  wire       [15:0]   _zz_7936;
  wire       [15:0]   _zz_7937;
  wire       [15:0]   _zz_7938;
  wire       [15:0]   _zz_7939;
  wire       [15:0]   _zz_7940;
  wire       [15:0]   _zz_7941;
  wire       [15:0]   _zz_7942;
  wire       [15:0]   _zz_7943;
  wire       [15:0]   _zz_7944;
  wire       [15:0]   _zz_7945;
  wire       [15:0]   _zz_7946;
  wire       [15:0]   _zz_7947;
  wire       [15:0]   _zz_7948;
  wire       [15:0]   _zz_7949;
  wire       [15:0]   _zz_7950;
  wire       [15:0]   _zz_7951;
  wire       [15:0]   _zz_7952;
  wire       [15:0]   _zz_7953;
  wire       [15:0]   _zz_7954;
  wire       [15:0]   _zz_7955;
  wire       [15:0]   _zz_7956;
  wire       [15:0]   _zz_7957;
  wire       [15:0]   _zz_7958;
  wire       [15:0]   _zz_7959;
  wire       [15:0]   _zz_7960;
  wire       [15:0]   _zz_7961;
  wire       [15:0]   _zz_7962;
  wire       [15:0]   _zz_7963;
  wire       [15:0]   _zz_7964;
  wire       [15:0]   _zz_7965;
  wire       [15:0]   _zz_7966;
  wire       [15:0]   _zz_7967;
  wire       [15:0]   _zz_7968;
  wire       [15:0]   _zz_7969;
  wire       [15:0]   _zz_7970;
  wire       [15:0]   _zz_7971;
  wire       [15:0]   _zz_7972;
  wire       [15:0]   _zz_7973;
  wire       [15:0]   _zz_7974;
  wire       [15:0]   _zz_7975;
  wire       [15:0]   _zz_7976;
  wire       [15:0]   _zz_7977;
  wire       [15:0]   _zz_7978;
  wire       [15:0]   _zz_7979;
  wire       [15:0]   _zz_7980;
  wire       [15:0]   _zz_7981;
  wire       [15:0]   _zz_7982;
  wire       [15:0]   _zz_7983;
  wire       [15:0]   _zz_7984;
  wire       [15:0]   _zz_7985;
  wire       [15:0]   _zz_7986;
  wire       [15:0]   _zz_7987;
  wire       [15:0]   _zz_7988;
  wire       [15:0]   _zz_7989;
  wire       [15:0]   _zz_7990;
  wire       [15:0]   _zz_7991;
  wire       [15:0]   _zz_7992;
  wire       [15:0]   _zz_7993;
  wire       [15:0]   _zz_7994;
  wire       [15:0]   _zz_7995;
  wire       [15:0]   _zz_7996;
  wire       [15:0]   _zz_7997;
  wire       [15:0]   _zz_7998;
  wire       [15:0]   _zz_7999;
  wire       [15:0]   _zz_8000;
  wire       [15:0]   _zz_8001;
  wire       [15:0]   _zz_8002;
  wire       [15:0]   _zz_8003;
  wire       [15:0]   _zz_8004;
  wire       [15:0]   _zz_8005;
  wire       [15:0]   _zz_8006;
  wire       [15:0]   _zz_8007;
  wire       [15:0]   _zz_8008;
  wire       [15:0]   _zz_8009;
  wire       [15:0]   _zz_8010;
  wire       [15:0]   _zz_8011;
  wire       [15:0]   _zz_8012;
  wire       [15:0]   _zz_8013;
  wire       [15:0]   _zz_8014;
  wire       [15:0]   _zz_8015;
  wire       [15:0]   _zz_8016;
  wire       [15:0]   _zz_8017;
  wire       [15:0]   _zz_8018;
  wire       [15:0]   _zz_8019;
  wire       [15:0]   _zz_8020;
  wire       [15:0]   _zz_8021;
  wire       [15:0]   _zz_8022;
  wire       [15:0]   _zz_8023;
  wire       [15:0]   _zz_8024;
  wire       [15:0]   _zz_8025;
  wire       [15:0]   _zz_8026;
  wire       [15:0]   _zz_8027;
  wire       [15:0]   _zz_8028;
  wire       [15:0]   _zz_8029;
  wire       [15:0]   _zz_8030;
  wire       [15:0]   _zz_8031;
  wire       [15:0]   _zz_8032;
  wire       [15:0]   _zz_8033;
  wire       [15:0]   _zz_8034;
  wire       [15:0]   _zz_8035;
  wire       [15:0]   _zz_8036;
  wire       [15:0]   _zz_8037;
  wire       [15:0]   _zz_8038;
  wire       [15:0]   _zz_8039;
  wire       [15:0]   _zz_8040;
  wire       [15:0]   _zz_8041;
  wire       [15:0]   _zz_8042;
  wire       [15:0]   _zz_8043;
  wire       [15:0]   _zz_8044;
  wire       [15:0]   _zz_8045;
  wire       [15:0]   _zz_8046;
  wire       [15:0]   _zz_8047;
  wire       [15:0]   _zz_8048;
  wire       [15:0]   _zz_8049;
  wire       [15:0]   _zz_8050;
  wire       [15:0]   _zz_8051;
  wire       [15:0]   _zz_8052;
  wire       [15:0]   _zz_8053;
  wire       [15:0]   _zz_8054;
  wire       [15:0]   _zz_8055;
  wire       [15:0]   _zz_8056;
  wire       [15:0]   _zz_8057;
  wire       [15:0]   _zz_8058;
  wire       [15:0]   _zz_8059;
  wire       [15:0]   _zz_8060;
  wire       [15:0]   _zz_8061;
  wire       [15:0]   _zz_8062;
  wire       [15:0]   _zz_8063;
  wire       [15:0]   _zz_8064;
  wire       [15:0]   _zz_8065;
  wire       [15:0]   _zz_8066;
  wire       [15:0]   _zz_8067;
  wire       [15:0]   _zz_8068;
  wire       [15:0]   _zz_8069;
  wire       [15:0]   _zz_8070;
  wire       [15:0]   _zz_8071;
  wire       [15:0]   _zz_8072;
  wire       [15:0]   _zz_8073;
  wire       [15:0]   _zz_8074;
  wire       [15:0]   _zz_8075;
  wire       [15:0]   _zz_8076;
  wire       [15:0]   _zz_8077;
  wire       [15:0]   _zz_8078;
  wire       [15:0]   _zz_8079;
  wire       [15:0]   _zz_8080;
  wire       [15:0]   _zz_8081;
  wire       [15:0]   _zz_8082;
  wire       [15:0]   _zz_8083;
  wire       [15:0]   _zz_8084;
  wire       [15:0]   _zz_8085;
  wire       [15:0]   _zz_8086;
  wire       [15:0]   _zz_8087;
  wire       [15:0]   _zz_8088;
  wire       [15:0]   _zz_8089;
  wire       [15:0]   _zz_8090;
  wire       [15:0]   _zz_8091;
  wire       [15:0]   _zz_8092;
  wire       [15:0]   _zz_8093;
  wire       [15:0]   _zz_8094;
  wire       [15:0]   _zz_8095;
  wire       [15:0]   _zz_8096;
  wire       [15:0]   _zz_8097;
  wire       [15:0]   _zz_8098;
  wire       [15:0]   _zz_8099;
  wire       [15:0]   _zz_8100;
  wire       [15:0]   _zz_8101;
  wire       [15:0]   _zz_8102;
  wire       [15:0]   _zz_8103;
  wire       [15:0]   _zz_8104;
  wire       [15:0]   _zz_8105;
  wire       [15:0]   _zz_8106;
  wire       [15:0]   _zz_8107;
  wire       [15:0]   _zz_8108;
  wire       [15:0]   _zz_8109;
  wire       [15:0]   _zz_8110;
  wire       [15:0]   _zz_8111;
  wire       [15:0]   _zz_8112;
  wire       [15:0]   _zz_8113;
  wire       [15:0]   _zz_8114;
  wire       [15:0]   _zz_8115;
  wire       [15:0]   _zz_8116;
  wire       [15:0]   _zz_8117;
  wire       [15:0]   _zz_8118;
  wire       [15:0]   _zz_8119;
  wire       [15:0]   _zz_8120;
  wire       [15:0]   _zz_8121;
  wire       [15:0]   _zz_8122;
  wire       [15:0]   _zz_8123;
  wire       [15:0]   _zz_8124;
  wire       [15:0]   _zz_8125;
  wire       [15:0]   _zz_8126;
  wire       [15:0]   _zz_8127;
  wire       [15:0]   _zz_8128;
  wire       [15:0]   _zz_8129;
  wire       [15:0]   _zz_8130;
  wire       [15:0]   _zz_8131;
  wire       [15:0]   _zz_8132;
  wire       [15:0]   _zz_8133;
  wire       [15:0]   _zz_8134;
  wire       [15:0]   _zz_8135;
  wire       [15:0]   _zz_8136;
  wire       [15:0]   _zz_8137;
  wire       [15:0]   _zz_8138;
  wire       [15:0]   _zz_8139;
  wire       [15:0]   _zz_8140;
  wire       [15:0]   _zz_8141;
  wire       [15:0]   _zz_8142;
  wire       [15:0]   _zz_8143;
  wire       [15:0]   _zz_8144;
  wire       [15:0]   _zz_8145;
  wire       [15:0]   _zz_8146;
  wire       [15:0]   _zz_8147;
  wire       [15:0]   _zz_8148;
  wire       [15:0]   _zz_8149;
  wire       [15:0]   _zz_8150;
  wire       [15:0]   _zz_8151;
  wire       [15:0]   _zz_8152;
  wire       [15:0]   _zz_8153;
  wire       [15:0]   _zz_8154;
  wire       [15:0]   _zz_8155;
  wire       [15:0]   _zz_8156;
  wire       [15:0]   _zz_8157;
  wire       [15:0]   _zz_8158;
  wire       [15:0]   _zz_8159;
  wire       [15:0]   _zz_8160;
  wire       [15:0]   _zz_8161;
  wire       [15:0]   _zz_8162;
  wire       [15:0]   _zz_8163;
  wire       [15:0]   _zz_8164;
  wire       [15:0]   _zz_8165;
  wire       [15:0]   _zz_8166;
  wire       [15:0]   _zz_8167;
  wire       [15:0]   _zz_8168;
  wire       [15:0]   _zz_8169;
  wire       [15:0]   _zz_8170;
  wire       [15:0]   _zz_8171;
  wire       [15:0]   _zz_8172;
  wire       [15:0]   _zz_8173;
  wire       [15:0]   _zz_8174;
  wire       [15:0]   _zz_8175;
  wire       [15:0]   _zz_8176;
  wire       [15:0]   _zz_8177;
  wire       [15:0]   _zz_8178;
  wire       [15:0]   _zz_8179;
  wire       [15:0]   _zz_8180;
  wire       [15:0]   _zz_8181;
  wire       [15:0]   _zz_8182;
  wire       [15:0]   _zz_8183;
  wire       [15:0]   _zz_8184;
  wire       [15:0]   _zz_8185;
  wire       [15:0]   _zz_8186;
  wire       [15:0]   _zz_8187;
  wire       [15:0]   _zz_8188;
  wire       [15:0]   _zz_8189;
  wire       [15:0]   _zz_8190;
  wire       [15:0]   _zz_8191;
  wire       [15:0]   _zz_8192;
  wire       [15:0]   _zz_8193;
  wire       [15:0]   _zz_8194;
  wire       [15:0]   _zz_8195;
  wire       [15:0]   _zz_8196;
  wire       [15:0]   _zz_8197;
  wire       [15:0]   _zz_8198;
  wire       [15:0]   _zz_8199;
  wire       [15:0]   _zz_8200;
  wire       [15:0]   _zz_8201;
  wire       [15:0]   _zz_8202;
  wire       [15:0]   _zz_8203;
  wire       [15:0]   _zz_8204;
  wire       [15:0]   _zz_8205;
  wire       [15:0]   _zz_8206;
  wire       [15:0]   _zz_8207;
  wire       [15:0]   _zz_8208;
  wire       [15:0]   _zz_8209;
  wire       [15:0]   _zz_8210;
  wire       [15:0]   _zz_8211;
  wire       [15:0]   _zz_8212;
  wire       [15:0]   _zz_8213;
  wire       [15:0]   _zz_8214;
  wire       [15:0]   _zz_8215;
  wire       [15:0]   _zz_8216;
  wire       [15:0]   _zz_8217;
  wire       [15:0]   _zz_8218;
  wire       [15:0]   _zz_8219;
  wire       [15:0]   _zz_8220;
  wire       [15:0]   _zz_8221;
  wire       [15:0]   _zz_8222;
  wire       [15:0]   _zz_8223;
  wire       [15:0]   _zz_8224;
  wire       [15:0]   _zz_8225;
  wire       [15:0]   _zz_8226;
  wire       [15:0]   _zz_8227;
  wire       [15:0]   _zz_8228;
  wire       [15:0]   _zz_8229;
  wire       [15:0]   _zz_8230;
  wire       [15:0]   _zz_8231;
  wire       [15:0]   _zz_8232;
  wire       [15:0]   _zz_8233;
  wire       [15:0]   _zz_8234;
  wire       [15:0]   _zz_8235;
  wire       [15:0]   _zz_8236;
  wire       [15:0]   _zz_8237;
  wire       [15:0]   _zz_8238;
  wire       [15:0]   _zz_8239;
  wire       [15:0]   _zz_8240;
  wire       [15:0]   _zz_8241;
  wire       [15:0]   _zz_8242;
  wire       [15:0]   _zz_8243;
  wire       [15:0]   _zz_8244;
  wire       [15:0]   _zz_8245;
  wire       [15:0]   _zz_8246;
  wire       [15:0]   _zz_8247;
  wire       [15:0]   _zz_8248;
  wire       [15:0]   _zz_8249;
  wire       [15:0]   _zz_8250;
  wire       [15:0]   _zz_8251;
  wire       [15:0]   _zz_8252;
  wire       [15:0]   _zz_8253;
  wire       [15:0]   _zz_8254;
  wire       [15:0]   _zz_8255;
  wire       [15:0]   _zz_8256;
  wire       [15:0]   _zz_8257;
  wire       [15:0]   _zz_8258;
  wire       [15:0]   _zz_8259;
  wire       [15:0]   _zz_8260;
  wire       [15:0]   _zz_8261;
  wire       [15:0]   _zz_8262;
  wire       [15:0]   _zz_8263;
  wire       [15:0]   _zz_8264;
  wire       [15:0]   _zz_8265;
  wire       [15:0]   _zz_8266;
  wire       [15:0]   _zz_8267;
  wire       [15:0]   _zz_8268;
  wire       [15:0]   _zz_8269;
  wire       [15:0]   _zz_8270;
  wire       [15:0]   _zz_8271;
  wire       [15:0]   _zz_8272;
  wire       [15:0]   _zz_8273;
  wire       [15:0]   _zz_8274;
  wire       [15:0]   _zz_8275;
  wire       [15:0]   _zz_8276;
  wire       [15:0]   _zz_8277;
  wire       [15:0]   _zz_8278;
  wire       [15:0]   _zz_8279;
  wire       [15:0]   _zz_8280;
  wire       [15:0]   _zz_8281;
  wire       [15:0]   _zz_8282;
  wire       [15:0]   _zz_8283;
  wire       [15:0]   _zz_8284;
  wire       [15:0]   _zz_8285;
  wire       [15:0]   _zz_8286;
  wire       [15:0]   _zz_8287;
  wire       [15:0]   _zz_8288;
  wire       [15:0]   _zz_8289;
  wire       [15:0]   _zz_8290;
  wire       [15:0]   _zz_8291;
  wire       [15:0]   _zz_8292;
  wire       [15:0]   _zz_8293;
  wire       [15:0]   _zz_8294;
  wire       [15:0]   _zz_8295;
  wire       [15:0]   _zz_8296;
  wire       [15:0]   _zz_8297;
  wire       [15:0]   _zz_8298;
  wire       [15:0]   _zz_8299;
  wire       [15:0]   _zz_8300;
  wire       [15:0]   _zz_8301;
  wire       [15:0]   _zz_8302;
  wire       [15:0]   _zz_8303;
  wire       [15:0]   _zz_8304;
  wire       [15:0]   _zz_8305;
  wire       [15:0]   _zz_8306;
  wire       [15:0]   _zz_8307;
  wire       [15:0]   _zz_8308;
  wire       [15:0]   _zz_8309;
  wire       [15:0]   _zz_8310;
  wire       [15:0]   _zz_8311;
  wire       [15:0]   _zz_8312;
  wire       [15:0]   _zz_8313;
  wire       [15:0]   _zz_8314;
  wire       [15:0]   _zz_8315;
  wire       [15:0]   _zz_8316;
  wire       [15:0]   _zz_8317;
  wire       [15:0]   _zz_8318;
  wire       [15:0]   _zz_8319;
  wire       [15:0]   _zz_8320;
  wire       [15:0]   _zz_8321;
  wire       [15:0]   _zz_8322;
  wire       [15:0]   _zz_8323;
  wire       [15:0]   _zz_8324;
  wire       [15:0]   _zz_8325;
  wire       [15:0]   _zz_8326;
  wire       [15:0]   _zz_8327;
  wire       [15:0]   _zz_8328;
  wire       [15:0]   _zz_8329;
  wire       [15:0]   _zz_8330;
  wire       [15:0]   _zz_8331;
  wire       [15:0]   _zz_8332;
  wire       [15:0]   _zz_8333;
  wire       [15:0]   _zz_8334;
  wire       [15:0]   _zz_8335;
  wire       [15:0]   _zz_8336;
  wire       [15:0]   _zz_8337;
  wire       [15:0]   _zz_8338;
  wire       [15:0]   _zz_8339;
  wire       [15:0]   _zz_8340;
  wire       [15:0]   _zz_8341;
  wire       [15:0]   _zz_8342;
  wire       [15:0]   _zz_8343;
  wire       [15:0]   _zz_8344;
  wire       [15:0]   _zz_8345;
  wire       [15:0]   _zz_8346;
  wire       [15:0]   _zz_8347;
  wire       [15:0]   _zz_8348;
  wire       [15:0]   _zz_8349;
  wire       [15:0]   _zz_8350;
  wire       [15:0]   _zz_8351;
  wire       [15:0]   _zz_8352;
  wire       [15:0]   _zz_8353;
  wire       [15:0]   _zz_8354;
  wire       [15:0]   _zz_8355;
  wire       [15:0]   _zz_8356;
  wire       [15:0]   _zz_8357;
  wire       [15:0]   _zz_8358;
  wire       [15:0]   _zz_8359;
  wire       [15:0]   _zz_8360;
  wire       [15:0]   _zz_8361;
  wire       [15:0]   _zz_8362;
  wire       [15:0]   _zz_8363;
  wire       [15:0]   _zz_8364;
  wire       [15:0]   _zz_8365;
  wire       [15:0]   _zz_8366;
  wire       [15:0]   _zz_8367;
  wire       [15:0]   _zz_8368;
  wire       [15:0]   _zz_8369;
  wire       [15:0]   _zz_8370;
  wire       [15:0]   _zz_8371;
  wire       [15:0]   _zz_8372;
  wire       [15:0]   _zz_8373;
  wire       [15:0]   _zz_8374;
  wire       [15:0]   _zz_8375;
  wire       [15:0]   _zz_8376;
  wire       [15:0]   _zz_8377;
  wire       [15:0]   _zz_8378;
  wire       [15:0]   _zz_8379;
  wire       [15:0]   _zz_8380;
  wire       [15:0]   _zz_8381;
  wire       [15:0]   _zz_8382;
  wire       [15:0]   _zz_8383;
  wire       [15:0]   _zz_8384;
  wire       [15:0]   _zz_8385;
  wire       [15:0]   _zz_8386;
  wire       [15:0]   _zz_8387;
  wire       [15:0]   _zz_8388;
  wire       [15:0]   _zz_8389;
  wire       [15:0]   _zz_8390;
  wire       [15:0]   _zz_8391;
  wire       [15:0]   _zz_8392;
  wire       [15:0]   _zz_8393;
  wire       [15:0]   _zz_8394;
  wire       [15:0]   _zz_8395;
  wire       [15:0]   _zz_8396;
  wire       [15:0]   _zz_8397;
  wire       [15:0]   _zz_8398;
  wire       [15:0]   _zz_8399;
  wire       [15:0]   _zz_8400;
  wire       [15:0]   _zz_8401;
  wire       [15:0]   _zz_8402;
  wire       [15:0]   _zz_8403;
  wire       [15:0]   _zz_8404;
  wire       [15:0]   _zz_8405;
  wire       [15:0]   _zz_8406;
  wire       [15:0]   _zz_8407;
  wire       [15:0]   _zz_8408;
  wire       [15:0]   _zz_8409;
  wire       [15:0]   _zz_8410;
  wire       [15:0]   _zz_8411;
  wire       [15:0]   _zz_8412;
  wire       [15:0]   _zz_8413;
  wire       [15:0]   _zz_8414;
  wire       [15:0]   _zz_8415;
  wire       [15:0]   _zz_8416;
  wire       [15:0]   _zz_8417;
  wire       [15:0]   _zz_8418;
  wire       [15:0]   _zz_8419;
  wire       [15:0]   _zz_8420;
  wire       [15:0]   _zz_8421;
  wire       [15:0]   _zz_8422;
  wire       [15:0]   _zz_8423;
  wire       [15:0]   _zz_8424;
  wire       [15:0]   _zz_8425;
  wire       [15:0]   _zz_8426;
  wire       [15:0]   _zz_8427;
  wire       [15:0]   _zz_8428;
  wire       [15:0]   _zz_8429;
  wire       [15:0]   _zz_8430;
  wire       [15:0]   _zz_8431;
  wire       [15:0]   _zz_8432;
  wire       [15:0]   _zz_8433;
  wire       [15:0]   _zz_8434;
  wire       [15:0]   _zz_8435;
  wire       [15:0]   _zz_8436;
  wire       [15:0]   _zz_8437;
  wire       [15:0]   _zz_8438;
  wire       [15:0]   _zz_8439;
  wire       [15:0]   _zz_8440;
  wire       [15:0]   _zz_8441;
  wire       [15:0]   _zz_8442;
  wire       [15:0]   _zz_8443;
  wire       [15:0]   _zz_8444;
  wire       [15:0]   _zz_8445;
  wire       [15:0]   _zz_8446;
  wire       [15:0]   _zz_8447;
  wire       [15:0]   _zz_8448;
  wire       [15:0]   _zz_8449;
  wire       [15:0]   _zz_8450;
  wire       [15:0]   _zz_8451;
  wire       [15:0]   _zz_8452;
  wire       [15:0]   _zz_8453;
  wire       [15:0]   _zz_8454;
  wire       [15:0]   _zz_8455;
  wire       [15:0]   _zz_8456;
  wire       [15:0]   _zz_8457;
  wire       [15:0]   _zz_8458;
  wire       [15:0]   _zz_8459;
  wire       [15:0]   _zz_8460;
  wire       [15:0]   _zz_8461;
  wire       [15:0]   _zz_8462;
  wire       [15:0]   _zz_8463;
  wire       [15:0]   _zz_8464;
  wire       [15:0]   _zz_8465;
  wire       [15:0]   _zz_8466;
  wire       [15:0]   _zz_8467;
  wire       [15:0]   _zz_8468;
  wire       [15:0]   _zz_8469;
  wire       [15:0]   _zz_8470;
  wire       [15:0]   _zz_8471;
  wire       [15:0]   _zz_8472;
  wire       [15:0]   _zz_8473;
  wire       [15:0]   _zz_8474;
  wire       [15:0]   _zz_8475;
  wire       [15:0]   _zz_8476;
  wire       [15:0]   _zz_8477;
  wire       [15:0]   _zz_8478;
  wire       [15:0]   _zz_8479;
  wire       [15:0]   _zz_8480;
  wire       [15:0]   _zz_8481;
  wire       [15:0]   _zz_8482;
  wire       [15:0]   _zz_8483;
  wire       [15:0]   _zz_8484;
  wire       [15:0]   _zz_8485;
  wire       [15:0]   _zz_8486;
  wire       [15:0]   _zz_8487;
  wire       [15:0]   _zz_8488;
  wire       [15:0]   _zz_8489;
  wire       [15:0]   _zz_8490;
  wire       [15:0]   _zz_8491;
  wire       [15:0]   _zz_8492;
  wire       [15:0]   _zz_8493;
  wire       [15:0]   _zz_8494;
  wire       [15:0]   _zz_8495;
  wire       [15:0]   _zz_8496;
  wire       [15:0]   _zz_8497;
  wire       [15:0]   _zz_8498;
  wire       [15:0]   _zz_8499;
  wire       [15:0]   _zz_8500;
  wire       [15:0]   _zz_8501;
  wire       [15:0]   _zz_8502;
  wire       [15:0]   _zz_8503;
  wire       [15:0]   _zz_8504;
  wire       [15:0]   _zz_8505;
  wire       [15:0]   _zz_8506;
  wire       [15:0]   _zz_8507;
  wire       [15:0]   _zz_8508;
  wire       [15:0]   _zz_8509;
  wire       [15:0]   _zz_8510;
  wire       [15:0]   _zz_8511;
  wire       [15:0]   _zz_8512;
  wire       [15:0]   _zz_8513;
  wire       [15:0]   _zz_8514;
  wire       [15:0]   _zz_8515;
  wire       [15:0]   _zz_8516;
  wire       [15:0]   _zz_8517;
  wire       [15:0]   _zz_8518;
  wire       [15:0]   _zz_8519;
  wire       [15:0]   _zz_8520;
  wire       [15:0]   _zz_8521;
  wire       [15:0]   _zz_8522;
  wire       [15:0]   _zz_8523;
  wire       [15:0]   _zz_8524;
  wire       [15:0]   _zz_8525;
  wire       [15:0]   _zz_8526;
  wire       [15:0]   _zz_8527;
  wire       [15:0]   _zz_8528;
  wire       [15:0]   _zz_8529;
  wire       [15:0]   _zz_8530;
  wire       [15:0]   _zz_8531;
  wire       [15:0]   _zz_8532;
  wire       [15:0]   _zz_8533;
  wire       [15:0]   _zz_8534;
  wire       [15:0]   _zz_8535;
  wire       [15:0]   _zz_8536;
  wire       [15:0]   _zz_8537;
  wire       [15:0]   _zz_8538;
  wire       [15:0]   _zz_8539;
  wire       [15:0]   _zz_8540;
  wire       [15:0]   _zz_8541;
  wire       [15:0]   _zz_8542;
  wire       [15:0]   _zz_8543;
  wire       [15:0]   _zz_8544;
  wire       [15:0]   _zz_8545;
  wire       [15:0]   _zz_8546;
  wire       [15:0]   _zz_8547;
  wire       [15:0]   _zz_8548;
  wire       [15:0]   _zz_8549;
  wire       [15:0]   _zz_8550;
  wire       [15:0]   _zz_8551;
  wire       [15:0]   _zz_8552;
  wire       [15:0]   _zz_8553;
  wire       [15:0]   _zz_8554;
  wire       [15:0]   _zz_8555;
  wire       [15:0]   _zz_8556;
  wire       [15:0]   _zz_8557;
  wire       [15:0]   _zz_8558;
  wire       [15:0]   _zz_8559;
  wire       [15:0]   _zz_8560;
  wire       [15:0]   _zz_8561;
  wire       [15:0]   _zz_8562;
  wire       [15:0]   _zz_8563;
  wire       [15:0]   _zz_8564;
  wire       [15:0]   _zz_8565;
  wire       [15:0]   _zz_8566;
  wire       [15:0]   _zz_8567;
  wire       [15:0]   _zz_8568;
  wire       [15:0]   _zz_8569;
  wire       [15:0]   _zz_8570;
  wire       [15:0]   _zz_8571;
  wire       [15:0]   _zz_8572;
  wire       [15:0]   _zz_8573;
  wire       [15:0]   _zz_8574;
  wire       [15:0]   _zz_8575;
  wire       [15:0]   _zz_8576;
  wire       [15:0]   _zz_8577;
  wire       [15:0]   _zz_8578;
  wire       [15:0]   _zz_8579;
  wire       [15:0]   _zz_8580;
  wire       [15:0]   _zz_8581;
  wire       [15:0]   _zz_8582;
  wire       [15:0]   _zz_8583;
  wire       [15:0]   _zz_8584;
  wire       [15:0]   _zz_8585;
  wire       [15:0]   _zz_8586;
  wire       [15:0]   _zz_8587;
  wire       [15:0]   _zz_8588;
  wire       [15:0]   _zz_8589;
  wire       [15:0]   _zz_8590;
  wire       [15:0]   _zz_8591;
  wire       [15:0]   _zz_8592;
  wire       [15:0]   _zz_8593;
  wire       [15:0]   _zz_8594;
  wire       [15:0]   _zz_8595;
  wire       [15:0]   _zz_8596;
  wire       [15:0]   _zz_8597;
  wire       [15:0]   _zz_8598;
  wire       [15:0]   _zz_8599;
  wire       [15:0]   _zz_8600;
  wire       [15:0]   _zz_8601;
  wire       [15:0]   _zz_8602;
  wire       [15:0]   _zz_8603;
  wire       [15:0]   _zz_8604;
  wire       [15:0]   _zz_8605;
  wire       [15:0]   _zz_8606;
  wire       [15:0]   _zz_8607;
  wire       [15:0]   _zz_8608;
  wire       [15:0]   _zz_8609;
  wire       [15:0]   _zz_8610;
  wire       [15:0]   _zz_8611;
  wire       [15:0]   _zz_8612;
  wire       [15:0]   _zz_8613;
  wire       [15:0]   _zz_8614;
  wire       [15:0]   _zz_8615;
  wire       [15:0]   _zz_8616;
  wire       [15:0]   _zz_8617;
  wire       [15:0]   _zz_8618;
  wire       [15:0]   _zz_8619;
  wire       [15:0]   _zz_8620;
  wire       [15:0]   _zz_8621;
  wire       [15:0]   _zz_8622;
  wire       [15:0]   _zz_8623;
  wire       [15:0]   _zz_8624;
  wire       [15:0]   _zz_8625;
  wire       [15:0]   _zz_8626;
  wire       [15:0]   _zz_8627;
  wire       [15:0]   _zz_8628;
  wire       [15:0]   _zz_8629;
  wire       [15:0]   _zz_8630;
  wire       [15:0]   _zz_8631;
  wire       [15:0]   _zz_8632;
  wire       [15:0]   _zz_8633;
  wire       [15:0]   _zz_8634;
  wire       [15:0]   _zz_8635;
  wire       [15:0]   _zz_8636;
  wire       [15:0]   _zz_8637;
  wire       [15:0]   _zz_8638;
  wire       [15:0]   _zz_8639;
  wire       [15:0]   _zz_8640;
  wire       [15:0]   _zz_8641;
  wire       [15:0]   _zz_8642;
  wire       [15:0]   _zz_8643;
  wire       [15:0]   _zz_8644;
  wire       [15:0]   _zz_8645;
  wire       [15:0]   _zz_8646;
  wire       [15:0]   _zz_8647;
  wire       [15:0]   _zz_8648;
  wire       [15:0]   _zz_8649;
  wire       [15:0]   _zz_8650;
  wire       [15:0]   _zz_8651;
  wire       [15:0]   _zz_8652;
  wire       [15:0]   _zz_8653;
  wire       [15:0]   _zz_8654;
  wire       [15:0]   _zz_8655;
  wire       [15:0]   _zz_8656;
  wire       [15:0]   _zz_8657;
  wire       [15:0]   _zz_8658;
  wire       [15:0]   _zz_8659;
  wire       [15:0]   _zz_8660;
  wire       [15:0]   _zz_8661;
  wire       [15:0]   _zz_8662;
  wire       [15:0]   _zz_8663;
  wire       [15:0]   _zz_8664;
  wire       [15:0]   _zz_8665;
  wire       [15:0]   _zz_8666;
  wire       [15:0]   _zz_8667;
  wire       [15:0]   _zz_8668;
  wire       [15:0]   _zz_8669;
  wire       [15:0]   _zz_8670;
  wire       [15:0]   _zz_8671;
  wire       [15:0]   _zz_8672;
  wire       [15:0]   _zz_8673;
  wire       [15:0]   _zz_8674;
  wire       [15:0]   _zz_8675;
  wire       [15:0]   _zz_8676;
  wire       [15:0]   _zz_8677;
  wire       [15:0]   _zz_8678;
  wire       [15:0]   _zz_8679;
  wire       [15:0]   _zz_8680;
  wire       [15:0]   _zz_8681;
  wire       [15:0]   _zz_8682;
  wire       [15:0]   _zz_8683;
  wire       [15:0]   _zz_8684;
  wire       [15:0]   _zz_8685;
  wire       [15:0]   _zz_8686;
  wire       [15:0]   _zz_8687;
  wire       [15:0]   _zz_8688;
  wire       [15:0]   _zz_8689;
  wire       [15:0]   _zz_8690;
  wire       [15:0]   _zz_8691;
  wire       [15:0]   _zz_8692;
  wire       [15:0]   _zz_8693;
  wire       [15:0]   _zz_8694;
  wire       [15:0]   _zz_8695;
  wire       [15:0]   _zz_8696;
  wire       [15:0]   _zz_8697;
  wire       [15:0]   _zz_8698;
  wire       [15:0]   _zz_8699;
  wire       [15:0]   _zz_8700;
  wire       [15:0]   _zz_8701;
  wire       [15:0]   _zz_8702;
  wire       [15:0]   _zz_8703;
  wire       [15:0]   _zz_8704;
  wire       [15:0]   _zz_8705;
  wire       [15:0]   _zz_8706;
  wire       [15:0]   _zz_8707;
  wire       [15:0]   _zz_8708;
  wire       [15:0]   _zz_8709;
  wire       [15:0]   _zz_8710;
  wire       [15:0]   _zz_8711;
  wire       [15:0]   _zz_8712;
  wire       [15:0]   _zz_8713;
  wire       [15:0]   _zz_8714;
  wire       [15:0]   _zz_8715;
  wire       [15:0]   _zz_8716;
  wire       [15:0]   _zz_8717;
  wire       [15:0]   _zz_8718;
  wire       [15:0]   _zz_8719;
  wire       [15:0]   _zz_8720;
  wire       [15:0]   _zz_8721;
  wire       [15:0]   _zz_8722;
  wire       [15:0]   _zz_8723;
  wire       [15:0]   _zz_8724;
  wire       [15:0]   _zz_8725;
  wire       [15:0]   _zz_8726;
  wire       [15:0]   _zz_8727;
  wire       [15:0]   _zz_8728;
  wire       [15:0]   _zz_8729;
  wire       [15:0]   _zz_8730;
  wire       [15:0]   _zz_8731;
  wire       [15:0]   _zz_8732;
  wire       [15:0]   _zz_8733;
  wire       [15:0]   _zz_8734;
  wire       [15:0]   _zz_8735;
  wire       [15:0]   _zz_8736;
  wire       [15:0]   _zz_8737;
  wire       [15:0]   _zz_8738;
  wire       [15:0]   _zz_8739;
  wire       [15:0]   _zz_8740;
  wire       [15:0]   _zz_8741;
  wire       [15:0]   _zz_8742;
  wire       [15:0]   _zz_8743;
  wire       [15:0]   _zz_8744;
  wire       [15:0]   _zz_8745;
  wire       [15:0]   _zz_8746;
  wire       [15:0]   _zz_8747;
  wire       [15:0]   _zz_8748;
  wire       [15:0]   _zz_8749;
  wire       [15:0]   _zz_8750;
  wire       [15:0]   _zz_8751;
  wire       [15:0]   _zz_8752;
  wire       [15:0]   _zz_8753;
  wire       [15:0]   _zz_8754;
  wire       [15:0]   _zz_8755;
  wire       [15:0]   _zz_8756;
  wire       [15:0]   _zz_8757;
  wire       [15:0]   _zz_8758;
  wire       [15:0]   _zz_8759;
  wire       [15:0]   _zz_8760;
  wire       [15:0]   _zz_8761;
  wire       [15:0]   _zz_8762;
  wire       [15:0]   _zz_8763;
  wire       [15:0]   _zz_8764;
  wire       [15:0]   _zz_8765;
  wire       [15:0]   _zz_8766;
  wire       [15:0]   _zz_8767;
  wire       [15:0]   _zz_8768;
  wire       [15:0]   _zz_8769;
  wire       [15:0]   _zz_8770;
  wire       [15:0]   _zz_8771;
  wire       [15:0]   _zz_8772;
  wire       [15:0]   _zz_8773;
  wire       [15:0]   _zz_8774;
  wire       [15:0]   _zz_8775;
  wire       [15:0]   _zz_8776;
  wire       [15:0]   _zz_8777;
  wire       [15:0]   _zz_8778;
  wire       [15:0]   _zz_8779;
  wire       [15:0]   _zz_8780;
  wire       [15:0]   _zz_8781;
  wire       [15:0]   _zz_8782;
  wire       [15:0]   _zz_8783;
  wire       [15:0]   _zz_8784;
  wire       [15:0]   _zz_8785;
  wire       [15:0]   _zz_8786;
  wire       [15:0]   _zz_8787;
  wire       [15:0]   _zz_8788;
  wire       [15:0]   _zz_8789;
  wire       [15:0]   _zz_8790;
  wire       [15:0]   _zz_8791;
  wire       [15:0]   _zz_8792;
  wire       [15:0]   _zz_8793;
  wire       [15:0]   _zz_8794;
  wire       [15:0]   _zz_8795;
  wire       [15:0]   _zz_8796;
  wire       [15:0]   _zz_8797;
  wire       [15:0]   _zz_8798;
  wire       [15:0]   _zz_8799;
  wire       [15:0]   _zz_8800;
  wire       [15:0]   _zz_8801;
  wire       [15:0]   _zz_8802;
  wire       [15:0]   _zz_8803;
  wire       [15:0]   _zz_8804;
  wire       [15:0]   _zz_8805;
  wire       [15:0]   _zz_8806;
  wire       [15:0]   _zz_8807;
  wire       [15:0]   _zz_8808;
  wire       [15:0]   _zz_8809;
  wire       [15:0]   _zz_8810;
  wire       [15:0]   _zz_8811;
  wire       [15:0]   _zz_8812;
  wire       [15:0]   _zz_8813;
  wire       [15:0]   _zz_8814;
  wire       [15:0]   _zz_8815;
  wire       [15:0]   _zz_8816;
  wire       [15:0]   _zz_8817;
  wire       [15:0]   _zz_8818;
  wire       [15:0]   _zz_8819;
  wire       [15:0]   _zz_8820;
  wire       [15:0]   _zz_8821;
  wire       [15:0]   _zz_8822;
  wire       [15:0]   _zz_8823;
  wire       [15:0]   _zz_8824;
  wire       [15:0]   _zz_8825;
  wire       [15:0]   _zz_8826;
  wire       [15:0]   _zz_8827;
  wire       [15:0]   _zz_8828;
  wire       [15:0]   _zz_8829;
  wire       [15:0]   _zz_8830;
  wire       [15:0]   _zz_8831;
  wire       [15:0]   _zz_8832;
  wire       [15:0]   _zz_8833;
  wire       [15:0]   _zz_8834;
  wire       [15:0]   _zz_8835;
  wire       [15:0]   _zz_8836;
  wire       [15:0]   _zz_8837;
  wire       [15:0]   _zz_8838;
  wire       [15:0]   _zz_8839;
  wire       [15:0]   _zz_8840;
  wire       [15:0]   _zz_8841;
  wire       [15:0]   _zz_8842;
  wire       [15:0]   _zz_8843;
  wire       [15:0]   _zz_8844;
  wire       [15:0]   _zz_8845;
  wire       [15:0]   _zz_8846;
  wire       [15:0]   _zz_8847;
  wire       [15:0]   _zz_8848;
  wire       [15:0]   _zz_8849;
  wire       [15:0]   _zz_8850;
  wire       [15:0]   _zz_8851;
  wire       [15:0]   _zz_8852;
  wire       [15:0]   _zz_8853;
  wire       [15:0]   _zz_8854;
  wire       [15:0]   _zz_8855;
  wire       [15:0]   _zz_8856;
  wire       [15:0]   _zz_8857;
  wire       [15:0]   _zz_8858;
  wire       [15:0]   _zz_8859;
  wire       [15:0]   _zz_8860;
  wire       [15:0]   _zz_8861;
  wire       [15:0]   _zz_8862;
  wire       [15:0]   _zz_8863;
  wire       [15:0]   _zz_8864;
  wire       [15:0]   _zz_8865;
  wire       [15:0]   _zz_8866;
  wire       [15:0]   _zz_8867;
  wire       [15:0]   _zz_8868;
  wire       [15:0]   _zz_8869;
  wire       [15:0]   _zz_8870;
  wire       [15:0]   _zz_8871;
  wire       [15:0]   _zz_8872;
  wire       [15:0]   _zz_8873;
  wire       [15:0]   _zz_8874;
  wire       [15:0]   _zz_8875;
  wire       [15:0]   _zz_8876;
  wire       [15:0]   _zz_8877;
  wire       [15:0]   _zz_8878;
  wire       [15:0]   _zz_8879;
  wire       [15:0]   _zz_8880;
  wire       [15:0]   _zz_8881;
  wire       [15:0]   _zz_8882;
  wire       [15:0]   _zz_8883;
  wire       [15:0]   _zz_8884;
  wire       [15:0]   _zz_8885;
  wire       [15:0]   _zz_8886;
  wire       [15:0]   _zz_8887;
  wire       [15:0]   _zz_8888;
  wire       [15:0]   _zz_8889;
  wire       [15:0]   _zz_8890;
  wire       [15:0]   _zz_8891;
  wire       [15:0]   _zz_8892;
  wire       [15:0]   _zz_8893;
  wire       [15:0]   _zz_8894;
  wire       [15:0]   _zz_8895;
  wire       [15:0]   _zz_8896;
  wire       [15:0]   _zz_8897;
  wire       [15:0]   _zz_8898;
  wire       [15:0]   _zz_8899;
  wire       [15:0]   _zz_8900;
  wire       [15:0]   _zz_8901;
  wire       [15:0]   _zz_8902;
  wire       [15:0]   _zz_8903;
  wire       [15:0]   _zz_8904;
  wire       [15:0]   _zz_8905;
  wire       [15:0]   _zz_8906;
  wire       [15:0]   _zz_8907;
  wire       [15:0]   _zz_8908;
  wire       [15:0]   _zz_8909;
  wire       [15:0]   _zz_8910;
  wire       [15:0]   _zz_8911;
  wire       [15:0]   _zz_8912;
  wire       [15:0]   _zz_8913;
  wire       [15:0]   _zz_8914;
  wire       [15:0]   _zz_8915;
  wire       [15:0]   _zz_8916;
  wire       [15:0]   _zz_8917;
  wire       [15:0]   _zz_8918;
  wire       [15:0]   _zz_8919;
  wire       [15:0]   _zz_8920;
  wire       [15:0]   _zz_8921;
  wire       [15:0]   _zz_8922;
  wire       [15:0]   _zz_8923;
  wire       [15:0]   _zz_8924;
  wire       [15:0]   _zz_8925;
  wire       [15:0]   _zz_8926;
  wire       [15:0]   _zz_8927;
  wire       [15:0]   _zz_8928;
  wire       [15:0]   _zz_8929;
  wire       [15:0]   _zz_8930;
  wire       [15:0]   _zz_8931;
  wire       [15:0]   _zz_8932;
  wire       [15:0]   _zz_8933;
  wire       [15:0]   _zz_8934;
  wire       [15:0]   _zz_8935;
  wire       [15:0]   _zz_8936;
  wire       [15:0]   _zz_8937;
  wire       [15:0]   _zz_8938;
  wire       [15:0]   _zz_8939;
  wire       [15:0]   _zz_8940;
  wire       [15:0]   _zz_8941;
  wire       [15:0]   _zz_8942;
  wire       [15:0]   _zz_8943;
  wire       [15:0]   _zz_8944;
  wire       [15:0]   _zz_8945;
  wire       [15:0]   _zz_8946;
  wire       [15:0]   _zz_8947;
  wire       [15:0]   _zz_8948;
  wire       [15:0]   _zz_8949;
  wire       [15:0]   _zz_8950;
  wire       [15:0]   _zz_8951;
  wire       [15:0]   _zz_8952;
  wire       [15:0]   _zz_8953;
  wire       [15:0]   _zz_8954;
  wire       [15:0]   _zz_8955;
  wire       [15:0]   _zz_8956;
  wire       [15:0]   _zz_8957;
  wire       [15:0]   _zz_8958;
  wire       [15:0]   _zz_8959;
  wire       [15:0]   _zz_8960;
  wire       [15:0]   _zz_8961;
  wire       [15:0]   _zz_8962;
  wire       [15:0]   _zz_8963;
  wire       [15:0]   _zz_8964;
  wire       [15:0]   _zz_8965;
  wire       [15:0]   _zz_8966;
  wire       [15:0]   _zz_8967;
  wire       [15:0]   _zz_8968;
  wire       [15:0]   _zz_8969;
  wire       [15:0]   _zz_8970;
  wire       [15:0]   _zz_8971;
  wire       [15:0]   _zz_8972;
  wire       [15:0]   _zz_8973;
  wire       [15:0]   _zz_8974;
  wire       [15:0]   _zz_8975;
  wire       [15:0]   _zz_8976;
  wire       [15:0]   _zz_8977;
  wire       [15:0]   _zz_8978;
  wire       [15:0]   _zz_8979;
  wire       [15:0]   _zz_8980;
  wire       [15:0]   _zz_8981;
  wire       [15:0]   _zz_8982;
  wire       [15:0]   _zz_8983;
  wire       [15:0]   _zz_8984;
  wire       [15:0]   _zz_8985;
  wire       [15:0]   _zz_8986;
  wire       [15:0]   _zz_8987;
  wire       [15:0]   _zz_8988;
  wire       [15:0]   _zz_8989;
  wire       [15:0]   _zz_8990;
  wire       [15:0]   _zz_8991;
  wire       [15:0]   _zz_8992;
  wire       [15:0]   _zz_8993;
  wire       [15:0]   _zz_8994;
  wire       [15:0]   _zz_8995;
  wire       [15:0]   _zz_8996;
  wire       [15:0]   _zz_8997;
  wire       [15:0]   _zz_8998;
  wire       [15:0]   _zz_8999;
  wire       [15:0]   _zz_9000;
  wire       [15:0]   _zz_9001;
  wire       [15:0]   _zz_9002;
  wire       [15:0]   _zz_9003;
  wire       [15:0]   _zz_9004;
  wire       [15:0]   _zz_9005;
  wire       [15:0]   _zz_9006;
  wire       [15:0]   _zz_9007;
  wire       [15:0]   _zz_9008;
  wire       [15:0]   _zz_9009;
  wire       [15:0]   _zz_9010;
  wire       [15:0]   _zz_9011;
  wire       [15:0]   _zz_9012;
  wire       [15:0]   _zz_9013;
  wire       [15:0]   _zz_9014;
  wire       [15:0]   _zz_9015;
  wire       [15:0]   _zz_9016;
  wire       [15:0]   _zz_9017;
  wire       [15:0]   _zz_9018;
  wire       [15:0]   _zz_9019;
  wire       [15:0]   _zz_9020;
  wire       [15:0]   _zz_9021;
  wire       [15:0]   _zz_9022;
  wire       [15:0]   _zz_9023;
  wire       [15:0]   _zz_9024;
  wire       [15:0]   _zz_9025;
  wire       [15:0]   _zz_9026;
  wire       [15:0]   _zz_9027;
  wire       [15:0]   _zz_9028;
  wire       [15:0]   _zz_9029;
  wire       [15:0]   _zz_9030;
  wire       [15:0]   _zz_9031;
  wire       [15:0]   _zz_9032;
  wire       [15:0]   _zz_9033;
  wire       [15:0]   _zz_9034;
  wire       [15:0]   _zz_9035;
  wire       [15:0]   _zz_9036;
  wire       [15:0]   _zz_9037;
  wire       [15:0]   _zz_9038;
  wire       [15:0]   _zz_9039;
  wire       [15:0]   _zz_9040;
  wire       [15:0]   _zz_9041;
  wire       [15:0]   _zz_9042;
  wire       [15:0]   _zz_9043;
  wire       [15:0]   _zz_9044;
  wire       [15:0]   _zz_9045;
  wire       [15:0]   _zz_9046;
  wire       [15:0]   _zz_9047;
  wire       [15:0]   _zz_9048;
  wire       [15:0]   _zz_9049;
  wire       [15:0]   _zz_9050;
  wire       [15:0]   _zz_9051;
  wire       [15:0]   _zz_9052;
  wire       [15:0]   _zz_9053;
  wire       [15:0]   _zz_9054;
  wire       [15:0]   _zz_9055;
  wire       [15:0]   _zz_9056;
  wire       [15:0]   _zz_9057;
  wire       [15:0]   _zz_9058;
  wire       [15:0]   _zz_9059;
  wire       [15:0]   _zz_9060;
  wire       [15:0]   _zz_9061;
  wire       [15:0]   _zz_9062;
  wire       [15:0]   _zz_9063;
  wire       [15:0]   _zz_9064;
  wire       [15:0]   _zz_9065;
  wire       [15:0]   _zz_9066;
  wire       [15:0]   _zz_9067;
  wire       [15:0]   _zz_9068;
  wire       [15:0]   _zz_9069;
  wire       [15:0]   _zz_9070;
  wire       [15:0]   _zz_9071;
  wire       [15:0]   _zz_9072;
  wire       [15:0]   _zz_9073;
  wire       [15:0]   _zz_9074;
  wire       [15:0]   _zz_9075;
  wire       [15:0]   _zz_9076;
  wire       [15:0]   _zz_9077;
  wire       [15:0]   _zz_9078;
  wire       [15:0]   _zz_9079;
  wire       [15:0]   _zz_9080;
  wire       [15:0]   _zz_9081;
  wire       [15:0]   _zz_9082;
  wire       [15:0]   _zz_9083;
  wire       [15:0]   _zz_9084;
  wire       [15:0]   _zz_9085;
  wire       [15:0]   _zz_9086;
  wire       [15:0]   _zz_9087;
  wire       [15:0]   _zz_9088;
  wire       [15:0]   _zz_9089;
  wire       [15:0]   _zz_9090;
  wire       [15:0]   _zz_9091;
  wire       [15:0]   _zz_9092;
  wire       [15:0]   _zz_9093;
  wire       [15:0]   _zz_9094;
  wire       [15:0]   _zz_9095;
  wire       [15:0]   _zz_9096;
  wire       [15:0]   _zz_9097;
  wire       [15:0]   _zz_9098;
  wire       [15:0]   _zz_9099;
  wire       [15:0]   _zz_9100;
  wire       [15:0]   _zz_9101;
  wire       [15:0]   _zz_9102;
  wire       [15:0]   _zz_9103;
  wire       [15:0]   _zz_9104;
  wire       [15:0]   _zz_9105;
  wire       [15:0]   _zz_9106;
  wire       [15:0]   _zz_9107;
  wire       [15:0]   _zz_9108;
  wire       [15:0]   _zz_9109;
  wire       [15:0]   _zz_9110;
  wire       [15:0]   _zz_9111;
  wire       [15:0]   _zz_9112;
  wire       [15:0]   _zz_9113;
  wire       [15:0]   _zz_9114;
  wire       [15:0]   _zz_9115;
  wire       [15:0]   _zz_9116;
  wire       [15:0]   _zz_9117;
  wire       [15:0]   _zz_9118;
  wire       [15:0]   _zz_9119;
  wire       [15:0]   _zz_9120;
  wire       [15:0]   _zz_9121;
  wire       [15:0]   _zz_9122;
  wire       [15:0]   _zz_9123;
  wire       [15:0]   _zz_9124;
  wire       [15:0]   _zz_9125;
  wire       [15:0]   _zz_9126;
  wire       [15:0]   _zz_9127;
  wire       [15:0]   _zz_9128;
  wire       [15:0]   _zz_9129;
  wire       [15:0]   _zz_9130;
  wire       [15:0]   _zz_9131;
  wire       [15:0]   _zz_9132;
  wire       [15:0]   _zz_9133;
  wire       [15:0]   _zz_9134;
  wire       [15:0]   _zz_9135;
  wire       [15:0]   _zz_9136;
  wire       [15:0]   _zz_9137;
  wire       [15:0]   _zz_9138;
  wire       [15:0]   _zz_9139;
  wire       [15:0]   _zz_9140;
  wire       [15:0]   _zz_9141;
  wire       [15:0]   _zz_9142;
  wire       [15:0]   _zz_9143;
  wire       [15:0]   _zz_9144;
  wire       [15:0]   _zz_9145;
  wire       [15:0]   _zz_9146;
  wire       [15:0]   _zz_9147;
  wire       [15:0]   _zz_9148;
  wire       [15:0]   _zz_9149;
  wire       [15:0]   _zz_9150;
  wire       [15:0]   _zz_9151;
  wire       [15:0]   _zz_9152;
  wire       [15:0]   _zz_9153;
  wire       [15:0]   _zz_9154;
  wire       [15:0]   _zz_9155;
  wire       [15:0]   _zz_9156;
  wire       [15:0]   _zz_9157;
  wire       [15:0]   _zz_9158;
  wire       [15:0]   _zz_9159;
  wire       [15:0]   _zz_9160;
  wire       [15:0]   _zz_9161;
  wire       [15:0]   _zz_9162;
  wire       [15:0]   _zz_9163;
  wire       [15:0]   _zz_9164;
  wire       [15:0]   _zz_9165;
  wire       [15:0]   _zz_9166;
  wire       [15:0]   _zz_9167;
  wire       [15:0]   _zz_9168;
  wire       [15:0]   _zz_9169;
  wire       [15:0]   _zz_9170;
  wire       [15:0]   _zz_9171;
  wire       [15:0]   _zz_9172;
  wire       [15:0]   _zz_9173;
  wire       [15:0]   _zz_9174;
  wire       [15:0]   _zz_9175;
  wire       [15:0]   _zz_9176;
  wire       [15:0]   _zz_9177;
  wire       [15:0]   _zz_9178;
  wire       [15:0]   _zz_9179;
  wire       [15:0]   _zz_9180;
  wire       [15:0]   _zz_9181;
  wire       [15:0]   _zz_9182;
  wire       [15:0]   _zz_9183;
  wire       [15:0]   _zz_9184;
  wire       [15:0]   _zz_9185;
  wire       [15:0]   _zz_9186;
  wire       [15:0]   _zz_9187;
  wire       [15:0]   _zz_9188;
  wire       [15:0]   _zz_9189;
  wire       [15:0]   _zz_9190;
  wire       [15:0]   _zz_9191;
  wire       [15:0]   _zz_9192;
  wire       [15:0]   _zz_9193;
  wire       [15:0]   _zz_9194;
  wire       [15:0]   _zz_9195;
  wire       [15:0]   _zz_9196;
  wire       [15:0]   _zz_9197;
  wire       [15:0]   _zz_9198;
  wire       [15:0]   _zz_9199;
  wire       [15:0]   _zz_9200;
  wire       [15:0]   _zz_9201;
  wire       [15:0]   _zz_9202;
  wire       [15:0]   _zz_9203;
  wire       [15:0]   _zz_9204;
  wire       [15:0]   _zz_9205;
  wire       [15:0]   _zz_9206;
  wire       [15:0]   _zz_9207;
  wire       [15:0]   _zz_9208;
  wire       [15:0]   _zz_9209;
  wire       [15:0]   _zz_9210;
  wire       [15:0]   _zz_9211;
  wire       [15:0]   _zz_9212;
  wire       [15:0]   _zz_9213;
  wire       [15:0]   _zz_9214;
  wire       [15:0]   _zz_9215;
  wire       [15:0]   _zz_9216;
  wire       [15:0]   _zz_9217;
  wire       [15:0]   _zz_9218;
  wire       [15:0]   _zz_9219;
  wire       [15:0]   _zz_9220;
  wire       [15:0]   _zz_9221;
  wire       [15:0]   _zz_9222;
  wire       [15:0]   _zz_9223;
  wire       [15:0]   _zz_9224;
  wire       [15:0]   _zz_9225;
  wire       [15:0]   _zz_9226;
  wire       [15:0]   _zz_9227;
  wire       [15:0]   _zz_9228;
  wire       [15:0]   _zz_9229;
  wire       [15:0]   _zz_9230;
  wire       [15:0]   _zz_9231;
  wire       [15:0]   _zz_9232;
  wire       [15:0]   _zz_9233;
  wire       [15:0]   _zz_9234;
  wire       [15:0]   _zz_9235;
  wire       [15:0]   _zz_9236;
  wire       [15:0]   _zz_9237;
  wire       [15:0]   _zz_9238;
  wire       [15:0]   _zz_9239;
  wire       [15:0]   _zz_9240;
  wire       [15:0]   _zz_9241;
  wire       [15:0]   _zz_9242;
  wire       [15:0]   _zz_9243;
  wire       [15:0]   _zz_9244;
  wire       [15:0]   _zz_9245;
  wire       [15:0]   _zz_9246;
  wire       [15:0]   _zz_9247;
  wire       [15:0]   _zz_9248;
  wire       [15:0]   _zz_9249;
  wire       [15:0]   _zz_9250;
  wire       [15:0]   _zz_9251;
  wire       [15:0]   _zz_9252;
  wire       [15:0]   _zz_9253;
  wire       [15:0]   _zz_9254;
  wire       [15:0]   _zz_9255;
  wire       [15:0]   _zz_9256;
  wire       [15:0]   _zz_9257;
  wire       [15:0]   _zz_9258;
  wire       [15:0]   _zz_9259;
  wire       [15:0]   _zz_9260;
  wire       [15:0]   _zz_9261;
  wire       [15:0]   _zz_9262;
  wire       [15:0]   _zz_9263;
  wire       [15:0]   _zz_9264;
  wire       [15:0]   _zz_9265;
  wire       [15:0]   _zz_9266;
  wire       [15:0]   _zz_9267;
  wire       [15:0]   _zz_9268;
  wire       [15:0]   _zz_9269;
  wire       [15:0]   _zz_9270;
  wire       [15:0]   _zz_9271;
  wire       [15:0]   _zz_9272;
  wire       [15:0]   _zz_9273;
  wire       [15:0]   _zz_9274;
  wire       [15:0]   _zz_9275;
  wire       [15:0]   _zz_9276;
  wire       [15:0]   _zz_9277;
  wire       [15:0]   _zz_9278;
  wire       [15:0]   _zz_9279;
  wire       [15:0]   _zz_9280;
  wire       [15:0]   _zz_9281;
  wire       [15:0]   _zz_9282;
  wire       [15:0]   _zz_9283;
  wire       [15:0]   _zz_9284;
  wire       [15:0]   _zz_9285;
  wire       [15:0]   _zz_9286;
  wire       [15:0]   _zz_9287;
  wire       [15:0]   _zz_9288;
  wire       [15:0]   _zz_9289;
  wire       [15:0]   _zz_9290;
  wire       [15:0]   _zz_9291;
  wire       [15:0]   _zz_9292;
  wire       [15:0]   _zz_9293;
  wire       [15:0]   _zz_9294;
  wire       [15:0]   _zz_9295;
  wire       [15:0]   _zz_9296;
  wire       [15:0]   _zz_9297;
  wire       [15:0]   _zz_9298;
  wire       [15:0]   _zz_9299;
  wire       [15:0]   _zz_9300;
  wire       [15:0]   _zz_9301;
  wire       [15:0]   _zz_9302;
  wire       [15:0]   _zz_9303;
  wire       [15:0]   _zz_9304;
  wire       [15:0]   _zz_9305;
  wire       [15:0]   _zz_9306;
  wire       [15:0]   _zz_9307;
  wire       [15:0]   _zz_9308;
  wire       [15:0]   _zz_9309;
  wire       [15:0]   _zz_9310;
  wire       [15:0]   _zz_9311;
  wire       [15:0]   _zz_9312;
  wire       [15:0]   _zz_9313;
  wire       [15:0]   _zz_9314;
  wire       [15:0]   _zz_9315;
  wire       [15:0]   _zz_9316;
  wire       [15:0]   _zz_9317;
  wire       [15:0]   _zz_9318;
  wire       [15:0]   _zz_9319;
  wire       [15:0]   _zz_9320;
  wire       [15:0]   _zz_9321;
  wire       [15:0]   _zz_9322;
  wire       [15:0]   _zz_9323;
  wire       [15:0]   _zz_9324;
  wire       [15:0]   _zz_9325;
  wire       [15:0]   _zz_9326;
  wire       [15:0]   _zz_9327;
  wire       [15:0]   _zz_9328;
  wire       [15:0]   _zz_9329;
  wire       [15:0]   _zz_9330;
  wire       [15:0]   _zz_9331;
  wire       [15:0]   _zz_9332;
  wire       [15:0]   _zz_9333;
  wire       [15:0]   _zz_9334;
  wire       [15:0]   _zz_9335;
  wire       [15:0]   _zz_9336;
  wire       [15:0]   _zz_9337;
  wire       [15:0]   _zz_9338;
  wire       [15:0]   _zz_9339;
  wire       [15:0]   _zz_9340;
  wire       [15:0]   _zz_9341;
  wire       [15:0]   _zz_9342;
  wire       [15:0]   _zz_9343;
  wire       [15:0]   _zz_9344;
  wire       [15:0]   _zz_9345;
  wire       [15:0]   _zz_9346;
  wire       [15:0]   _zz_9347;
  wire       [15:0]   _zz_9348;
  wire       [15:0]   _zz_9349;
  wire       [15:0]   _zz_9350;
  wire       [15:0]   _zz_9351;
  wire       [15:0]   _zz_9352;
  wire       [15:0]   _zz_9353;
  wire       [15:0]   _zz_9354;
  wire       [15:0]   _zz_9355;
  wire       [15:0]   _zz_9356;
  wire       [15:0]   _zz_9357;
  wire       [15:0]   _zz_9358;
  wire       [15:0]   _zz_9359;
  wire       [15:0]   _zz_9360;
  wire       [15:0]   _zz_9361;
  wire       [15:0]   _zz_9362;
  wire       [15:0]   _zz_9363;
  wire       [15:0]   _zz_9364;
  wire       [15:0]   _zz_9365;
  wire       [15:0]   _zz_9366;
  wire       [15:0]   _zz_9367;
  wire       [15:0]   _zz_9368;
  wire       [15:0]   _zz_9369;
  wire       [15:0]   _zz_9370;
  wire       [15:0]   _zz_9371;
  wire       [15:0]   _zz_9372;
  wire       [15:0]   _zz_9373;
  wire       [15:0]   _zz_9374;
  wire       [15:0]   _zz_9375;
  wire       [15:0]   _zz_9376;
  wire       [15:0]   _zz_9377;
  wire       [15:0]   _zz_9378;
  wire       [15:0]   _zz_9379;
  wire       [15:0]   _zz_9380;
  wire       [15:0]   _zz_9381;
  wire       [15:0]   _zz_9382;
  wire       [15:0]   _zz_9383;
  wire       [15:0]   _zz_9384;
  wire       [15:0]   _zz_9385;
  wire       [15:0]   _zz_9386;
  wire       [15:0]   _zz_9387;
  wire       [15:0]   _zz_9388;
  wire       [15:0]   _zz_9389;
  wire       [15:0]   _zz_9390;
  wire       [15:0]   _zz_9391;
  wire       [15:0]   _zz_9392;
  wire       [15:0]   _zz_9393;
  wire       [15:0]   _zz_9394;
  wire       [15:0]   _zz_9395;
  wire       [15:0]   _zz_9396;
  wire       [15:0]   _zz_9397;
  wire       [15:0]   _zz_9398;
  wire       [15:0]   _zz_9399;
  wire       [15:0]   _zz_9400;
  wire       [15:0]   _zz_9401;
  wire       [15:0]   _zz_9402;
  wire       [15:0]   _zz_9403;
  wire       [15:0]   _zz_9404;
  wire       [15:0]   _zz_9405;
  wire       [15:0]   _zz_9406;
  wire       [15:0]   _zz_9407;
  wire       [15:0]   _zz_9408;
  wire       [15:0]   _zz_9409;
  wire       [15:0]   _zz_9410;
  wire       [15:0]   _zz_9411;
  wire       [15:0]   _zz_9412;
  wire       [15:0]   _zz_9413;
  wire       [15:0]   _zz_9414;
  wire       [15:0]   _zz_9415;
  wire       [15:0]   _zz_9416;
  wire       [15:0]   _zz_9417;
  wire       [15:0]   _zz_9418;
  wire       [15:0]   _zz_9419;
  wire       [15:0]   _zz_9420;
  wire       [15:0]   _zz_9421;
  wire       [15:0]   _zz_9422;
  wire       [15:0]   _zz_9423;
  wire       [15:0]   _zz_9424;
  wire       [15:0]   _zz_9425;
  wire       [15:0]   _zz_9426;
  wire       [15:0]   _zz_9427;
  wire       [15:0]   _zz_9428;
  wire       [15:0]   _zz_9429;
  wire       [15:0]   _zz_9430;
  wire       [15:0]   _zz_9431;
  wire       [15:0]   _zz_9432;
  wire       [15:0]   _zz_9433;
  wire       [15:0]   _zz_9434;
  wire       [15:0]   _zz_9435;
  wire       [15:0]   _zz_9436;
  wire       [15:0]   _zz_9437;
  wire       [15:0]   _zz_9438;
  wire       [15:0]   _zz_9439;
  wire       [15:0]   _zz_9440;
  wire       [15:0]   _zz_9441;
  wire       [15:0]   _zz_9442;
  wire       [15:0]   _zz_9443;
  wire       [15:0]   _zz_9444;
  wire       [15:0]   _zz_9445;
  wire       [15:0]   _zz_9446;
  wire       [15:0]   _zz_9447;
  wire       [15:0]   _zz_9448;
  wire       [15:0]   _zz_9449;
  wire       [15:0]   _zz_9450;
  wire       [15:0]   _zz_9451;
  wire       [15:0]   _zz_9452;
  wire       [15:0]   _zz_9453;
  wire       [15:0]   _zz_9454;
  wire       [15:0]   _zz_9455;
  wire       [15:0]   _zz_9456;
  wire       [15:0]   _zz_9457;
  wire       [15:0]   _zz_9458;
  wire       [15:0]   _zz_9459;
  wire       [15:0]   _zz_9460;
  wire       [15:0]   _zz_9461;
  wire       [15:0]   _zz_9462;
  wire       [15:0]   _zz_9463;
  wire       [15:0]   _zz_9464;
  wire       [15:0]   _zz_9465;
  wire       [15:0]   _zz_9466;
  wire       [15:0]   _zz_9467;
  wire       [15:0]   _zz_9468;
  wire       [15:0]   _zz_9469;
  wire       [15:0]   _zz_9470;
  wire       [15:0]   _zz_9471;
  wire       [15:0]   _zz_9472;
  wire       [15:0]   _zz_9473;
  wire       [15:0]   _zz_9474;
  wire       [15:0]   _zz_9475;
  wire       [15:0]   _zz_9476;
  wire       [15:0]   _zz_9477;
  wire       [15:0]   _zz_9478;
  wire       [15:0]   _zz_9479;
  wire       [15:0]   _zz_9480;
  wire       [15:0]   _zz_9481;
  wire       [15:0]   _zz_9482;
  wire       [15:0]   _zz_9483;
  wire       [15:0]   _zz_9484;
  wire       [15:0]   _zz_9485;
  wire       [15:0]   _zz_9486;
  wire       [15:0]   _zz_9487;
  wire       [15:0]   _zz_9488;
  wire       [15:0]   _zz_9489;
  wire       [15:0]   _zz_9490;
  wire       [15:0]   _zz_9491;
  wire       [15:0]   _zz_9492;
  wire       [15:0]   _zz_9493;
  wire       [15:0]   _zz_9494;
  wire       [15:0]   _zz_9495;
  wire       [15:0]   _zz_9496;
  wire       [15:0]   _zz_9497;
  wire       [15:0]   _zz_9498;
  wire       [15:0]   _zz_9499;
  wire       [15:0]   _zz_9500;
  wire       [15:0]   _zz_9501;
  wire       [15:0]   _zz_9502;
  wire       [15:0]   _zz_9503;
  wire       [15:0]   _zz_9504;
  wire       [15:0]   _zz_9505;
  wire       [15:0]   _zz_9506;
  wire       [15:0]   _zz_9507;
  wire       [15:0]   _zz_9508;
  wire       [15:0]   _zz_9509;
  wire       [15:0]   _zz_9510;
  wire       [15:0]   _zz_9511;
  wire       [15:0]   _zz_9512;
  wire       [15:0]   _zz_9513;
  wire       [15:0]   _zz_9514;
  wire       [15:0]   _zz_9515;
  wire       [15:0]   _zz_9516;
  wire       [15:0]   _zz_9517;
  wire       [15:0]   _zz_9518;
  wire       [15:0]   _zz_9519;
  wire       [15:0]   _zz_9520;
  wire       [15:0]   _zz_9521;
  wire       [15:0]   _zz_9522;
  wire       [15:0]   _zz_9523;
  wire       [15:0]   _zz_9524;
  wire       [15:0]   _zz_9525;
  wire       [15:0]   _zz_9526;
  wire       [15:0]   _zz_9527;
  wire       [15:0]   _zz_9528;
  wire       [15:0]   _zz_9529;
  wire       [15:0]   _zz_9530;
  wire       [15:0]   _zz_9531;
  wire       [15:0]   _zz_9532;
  wire       [15:0]   _zz_9533;
  wire       [15:0]   _zz_9534;
  wire       [15:0]   _zz_9535;
  wire       [15:0]   _zz_9536;
  wire       [15:0]   _zz_9537;
  wire       [15:0]   _zz_9538;
  wire       [15:0]   _zz_9539;
  wire       [15:0]   _zz_9540;
  wire       [15:0]   _zz_9541;
  wire       [15:0]   _zz_9542;
  wire       [15:0]   _zz_9543;
  wire       [15:0]   _zz_9544;
  wire       [15:0]   _zz_9545;
  wire       [15:0]   _zz_9546;
  wire       [15:0]   _zz_9547;
  wire       [15:0]   _zz_9548;
  wire       [15:0]   _zz_9549;
  wire       [15:0]   _zz_9550;
  wire       [15:0]   _zz_9551;
  wire       [15:0]   _zz_9552;
  wire       [15:0]   _zz_9553;
  wire       [15:0]   _zz_9554;
  wire       [15:0]   _zz_9555;
  wire       [15:0]   _zz_9556;
  wire       [15:0]   _zz_9557;
  wire       [15:0]   _zz_9558;
  wire       [15:0]   _zz_9559;
  wire       [15:0]   _zz_9560;
  wire       [15:0]   _zz_9561;
  wire       [15:0]   _zz_9562;
  wire       [15:0]   _zz_9563;
  wire       [15:0]   _zz_9564;
  wire       [15:0]   _zz_9565;
  wire       [15:0]   _zz_9566;
  wire       [15:0]   _zz_9567;
  wire       [15:0]   _zz_9568;
  wire       [15:0]   _zz_9569;
  wire       [15:0]   _zz_9570;
  wire       [15:0]   _zz_9571;
  wire       [15:0]   _zz_9572;
  wire       [15:0]   _zz_9573;
  wire       [15:0]   _zz_9574;
  wire       [15:0]   _zz_9575;
  wire       [15:0]   _zz_9576;
  wire       [15:0]   _zz_9577;
  wire       [15:0]   _zz_9578;
  wire       [15:0]   _zz_9579;
  wire       [15:0]   _zz_9580;
  wire       [15:0]   _zz_9581;
  wire       [15:0]   _zz_9582;
  wire       [15:0]   _zz_9583;
  wire       [15:0]   _zz_9584;
  wire       [15:0]   _zz_9585;
  wire       [15:0]   _zz_9586;
  wire       [15:0]   _zz_9587;
  wire       [15:0]   _zz_9588;
  wire       [15:0]   _zz_9589;
  wire       [15:0]   _zz_9590;
  wire       [15:0]   _zz_9591;
  wire       [15:0]   _zz_9592;
  wire       [15:0]   _zz_9593;
  wire       [15:0]   _zz_9594;
  wire       [15:0]   _zz_9595;
  wire       [15:0]   _zz_9596;
  wire       [15:0]   _zz_9597;
  wire       [15:0]   _zz_9598;
  wire       [15:0]   _zz_9599;
  wire       [15:0]   _zz_9600;
  wire       [15:0]   _zz_9601;
  wire       [15:0]   _zz_9602;
  wire       [15:0]   _zz_9603;
  wire       [15:0]   _zz_9604;
  wire       [15:0]   _zz_9605;
  wire       [15:0]   _zz_9606;
  wire       [15:0]   _zz_9607;
  wire       [15:0]   _zz_9608;
  wire       [15:0]   _zz_9609;
  wire       [15:0]   _zz_9610;
  wire       [15:0]   _zz_9611;
  wire       [15:0]   _zz_9612;
  wire       [15:0]   _zz_9613;
  wire       [15:0]   _zz_9614;
  wire       [15:0]   _zz_9615;
  wire       [15:0]   _zz_9616;
  wire       [15:0]   _zz_9617;
  wire       [15:0]   _zz_9618;
  wire       [15:0]   _zz_9619;
  wire       [15:0]   _zz_9620;
  wire       [15:0]   _zz_9621;
  wire       [15:0]   _zz_9622;
  wire       [15:0]   _zz_9623;
  wire       [15:0]   _zz_9624;
  wire       [15:0]   _zz_9625;
  wire       [15:0]   _zz_9626;
  wire       [15:0]   _zz_9627;
  wire       [15:0]   _zz_9628;
  wire       [15:0]   _zz_9629;
  wire       [15:0]   _zz_9630;
  wire       [15:0]   _zz_9631;
  wire       [15:0]   _zz_9632;
  wire       [15:0]   _zz_9633;
  wire       [15:0]   _zz_9634;
  wire       [15:0]   _zz_9635;
  wire       [15:0]   _zz_9636;
  wire       [15:0]   _zz_9637;
  wire       [15:0]   _zz_9638;
  wire       [15:0]   _zz_9639;
  wire       [15:0]   _zz_9640;
  wire       [15:0]   _zz_9641;
  wire       [15:0]   _zz_9642;
  wire       [15:0]   _zz_9643;
  wire       [15:0]   _zz_9644;
  wire       [15:0]   _zz_9645;
  wire       [15:0]   _zz_9646;
  wire       [15:0]   _zz_9647;
  wire       [15:0]   _zz_9648;
  wire       [15:0]   _zz_9649;
  wire       [15:0]   _zz_9650;
  wire       [15:0]   _zz_9651;
  wire       [15:0]   _zz_9652;
  wire       [15:0]   _zz_9653;
  wire       [15:0]   _zz_9654;
  wire       [15:0]   _zz_9655;
  wire       [15:0]   _zz_9656;
  wire       [15:0]   _zz_9657;
  wire       [15:0]   _zz_9658;
  wire       [15:0]   _zz_9659;
  wire       [15:0]   _zz_9660;
  wire       [15:0]   _zz_9661;
  wire       [15:0]   _zz_9662;
  wire       [15:0]   _zz_9663;
  wire       [15:0]   _zz_9664;
  wire       [15:0]   _zz_9665;
  wire       [15:0]   _zz_9666;
  wire       [15:0]   _zz_9667;
  wire       [15:0]   _zz_9668;
  wire       [15:0]   _zz_9669;
  wire       [15:0]   _zz_9670;
  wire       [15:0]   _zz_9671;
  wire       [15:0]   _zz_9672;
  wire       [15:0]   _zz_9673;
  wire       [15:0]   _zz_9674;
  wire       [15:0]   _zz_9675;
  wire       [15:0]   _zz_9676;
  wire       [15:0]   _zz_9677;
  wire       [15:0]   _zz_9678;
  wire       [15:0]   _zz_9679;
  wire       [15:0]   _zz_9680;
  wire       [15:0]   _zz_9681;
  wire       [15:0]   _zz_9682;
  wire       [15:0]   _zz_9683;
  wire       [15:0]   _zz_9684;
  wire       [15:0]   _zz_9685;
  wire       [15:0]   _zz_9686;
  wire       [15:0]   _zz_9687;
  wire       [15:0]   _zz_9688;
  wire       [15:0]   _zz_9689;
  wire       [15:0]   _zz_9690;
  wire       [15:0]   _zz_9691;
  wire       [15:0]   _zz_9692;
  wire       [15:0]   _zz_9693;
  wire       [15:0]   _zz_9694;
  wire       [15:0]   _zz_9695;
  wire       [15:0]   _zz_9696;
  wire       [15:0]   _zz_9697;
  wire       [15:0]   _zz_9698;
  wire       [15:0]   _zz_9699;
  wire       [15:0]   _zz_9700;
  wire       [15:0]   _zz_9701;
  wire       [15:0]   _zz_9702;
  wire       [15:0]   _zz_9703;
  wire       [15:0]   _zz_9704;
  wire       [15:0]   _zz_9705;
  wire       [15:0]   _zz_9706;
  wire       [15:0]   _zz_9707;
  wire       [15:0]   _zz_9708;
  wire       [15:0]   _zz_9709;
  wire       [15:0]   _zz_9710;
  wire       [15:0]   _zz_9711;
  wire       [15:0]   _zz_9712;
  wire       [15:0]   _zz_9713;
  wire       [15:0]   _zz_9714;
  wire       [15:0]   _zz_9715;
  wire       [15:0]   _zz_9716;
  wire       [15:0]   _zz_9717;
  wire       [15:0]   _zz_9718;
  wire       [15:0]   _zz_9719;
  wire       [15:0]   _zz_9720;
  wire       [15:0]   _zz_9721;
  wire       [15:0]   _zz_9722;
  wire       [15:0]   _zz_9723;
  wire       [15:0]   _zz_9724;
  wire       [15:0]   _zz_9725;
  wire       [15:0]   _zz_9726;
  wire       [15:0]   _zz_9727;
  wire       [15:0]   _zz_9728;
  wire       [15:0]   _zz_9729;
  wire       [15:0]   _zz_9730;
  wire       [15:0]   _zz_9731;
  wire       [15:0]   _zz_9732;
  wire       [15:0]   _zz_9733;
  wire       [15:0]   _zz_9734;
  wire       [15:0]   _zz_9735;
  wire       [15:0]   _zz_9736;
  wire       [15:0]   _zz_9737;
  wire       [15:0]   _zz_9738;
  wire       [15:0]   _zz_9739;
  wire       [15:0]   _zz_9740;
  wire       [15:0]   _zz_9741;
  wire       [15:0]   _zz_9742;
  wire       [15:0]   _zz_9743;
  wire       [15:0]   _zz_9744;
  wire       [15:0]   _zz_9745;
  wire       [15:0]   _zz_9746;
  wire       [15:0]   _zz_9747;
  wire       [15:0]   _zz_9748;
  wire       [15:0]   _zz_9749;
  wire       [15:0]   _zz_9750;
  wire       [15:0]   _zz_9751;
  wire       [15:0]   _zz_9752;
  wire       [15:0]   _zz_9753;
  wire       [15:0]   _zz_9754;
  wire       [15:0]   _zz_9755;
  wire       [15:0]   _zz_9756;
  wire       [15:0]   _zz_9757;
  wire       [15:0]   _zz_9758;
  wire       [15:0]   _zz_9759;
  wire       [15:0]   _zz_9760;
  wire       [15:0]   _zz_9761;
  wire       [15:0]   _zz_9762;
  wire       [15:0]   _zz_9763;
  wire       [15:0]   _zz_9764;
  wire       [15:0]   _zz_9765;
  wire       [15:0]   _zz_9766;
  wire       [15:0]   _zz_9767;
  wire       [15:0]   _zz_9768;
  wire       [15:0]   _zz_9769;
  wire       [15:0]   _zz_9770;
  wire       [15:0]   _zz_9771;
  wire       [15:0]   _zz_9772;
  wire       [15:0]   _zz_9773;
  wire       [15:0]   _zz_9774;
  wire       [15:0]   _zz_9775;
  wire       [15:0]   _zz_9776;
  wire       [15:0]   _zz_9777;
  wire       [15:0]   _zz_9778;
  wire       [15:0]   _zz_9779;
  wire       [15:0]   _zz_9780;
  wire       [15:0]   _zz_9781;
  wire       [15:0]   _zz_9782;
  wire       [15:0]   _zz_9783;
  wire       [15:0]   _zz_9784;
  wire       [15:0]   _zz_9785;
  wire       [15:0]   _zz_9786;
  wire       [15:0]   _zz_9787;
  wire       [15:0]   _zz_9788;
  wire       [15:0]   _zz_9789;
  wire       [15:0]   _zz_9790;
  wire       [15:0]   _zz_9791;
  wire       [15:0]   _zz_9792;
  wire       [15:0]   _zz_9793;
  wire       [15:0]   _zz_9794;
  wire       [15:0]   _zz_9795;
  wire       [15:0]   _zz_9796;
  wire       [15:0]   _zz_9797;
  wire       [15:0]   _zz_9798;
  wire       [15:0]   _zz_9799;
  wire       [15:0]   _zz_9800;
  wire       [15:0]   _zz_9801;
  wire       [15:0]   _zz_9802;
  wire       [15:0]   _zz_9803;
  wire       [15:0]   _zz_9804;
  wire       [15:0]   _zz_9805;
  wire       [15:0]   _zz_9806;
  wire       [15:0]   _zz_9807;
  wire       [15:0]   _zz_9808;
  wire       [15:0]   _zz_9809;
  wire       [15:0]   _zz_9810;
  wire       [15:0]   _zz_9811;
  wire       [15:0]   _zz_9812;
  wire       [15:0]   _zz_9813;
  wire       [15:0]   _zz_9814;
  wire       [15:0]   _zz_9815;
  wire       [15:0]   _zz_9816;
  wire       [15:0]   _zz_9817;
  wire       [15:0]   _zz_9818;
  wire       [15:0]   _zz_9819;
  wire       [15:0]   _zz_9820;
  wire       [15:0]   _zz_9821;
  wire       [15:0]   _zz_9822;
  wire       [15:0]   _zz_9823;
  wire       [15:0]   _zz_9824;
  wire       [15:0]   _zz_9825;
  wire       [15:0]   _zz_9826;
  wire       [15:0]   _zz_9827;
  wire       [15:0]   _zz_9828;
  wire       [15:0]   _zz_9829;
  wire       [15:0]   _zz_9830;
  wire       [15:0]   _zz_9831;
  wire       [15:0]   _zz_9832;
  wire       [15:0]   _zz_9833;
  wire       [15:0]   _zz_9834;
  wire       [15:0]   _zz_9835;
  wire       [15:0]   _zz_9836;
  wire       [15:0]   _zz_9837;
  wire       [15:0]   _zz_9838;
  wire       [15:0]   _zz_9839;
  wire       [15:0]   _zz_9840;
  wire       [15:0]   _zz_9841;
  wire       [15:0]   _zz_9842;
  wire       [15:0]   _zz_9843;
  wire       [15:0]   _zz_9844;
  wire       [15:0]   _zz_9845;
  wire       [15:0]   _zz_9846;
  wire       [15:0]   _zz_9847;
  wire       [15:0]   _zz_9848;
  wire       [15:0]   _zz_9849;
  wire       [15:0]   _zz_9850;
  wire       [15:0]   _zz_9851;
  wire       [15:0]   _zz_9852;
  wire       [15:0]   _zz_9853;
  wire       [15:0]   _zz_9854;
  wire       [15:0]   _zz_9855;
  wire       [15:0]   _zz_9856;
  wire       [15:0]   _zz_9857;
  wire       [15:0]   _zz_9858;
  wire       [15:0]   _zz_9859;
  wire       [15:0]   _zz_9860;
  wire       [15:0]   _zz_9861;
  wire       [15:0]   _zz_9862;
  wire       [15:0]   _zz_9863;
  wire       [15:0]   _zz_9864;
  wire       [15:0]   _zz_9865;
  wire       [15:0]   _zz_9866;
  wire       [15:0]   _zz_9867;
  wire       [15:0]   _zz_9868;
  wire       [15:0]   _zz_9869;
  wire       [15:0]   _zz_9870;
  wire       [15:0]   _zz_9871;
  wire       [15:0]   _zz_9872;
  wire       [15:0]   _zz_9873;
  wire       [15:0]   _zz_9874;
  wire       [15:0]   _zz_9875;
  wire       [15:0]   _zz_9876;
  wire       [15:0]   _zz_9877;
  wire       [15:0]   _zz_9878;
  wire       [15:0]   _zz_9879;
  wire       [15:0]   _zz_9880;
  wire       [15:0]   _zz_9881;
  wire       [15:0]   _zz_9882;
  wire       [15:0]   _zz_9883;
  wire       [15:0]   _zz_9884;
  wire       [15:0]   _zz_9885;
  wire       [15:0]   _zz_9886;
  wire       [15:0]   _zz_9887;
  wire       [15:0]   _zz_9888;
  wire       [15:0]   _zz_9889;
  wire       [15:0]   _zz_9890;
  wire       [15:0]   _zz_9891;
  wire       [15:0]   _zz_9892;
  wire       [15:0]   _zz_9893;
  wire       [15:0]   _zz_9894;
  wire       [15:0]   _zz_9895;
  wire       [15:0]   _zz_9896;
  wire       [15:0]   _zz_9897;
  wire       [15:0]   _zz_9898;
  wire       [15:0]   _zz_9899;
  wire       [15:0]   _zz_9900;
  wire       [15:0]   _zz_9901;
  wire       [15:0]   _zz_9902;
  wire       [15:0]   _zz_9903;
  wire       [15:0]   _zz_9904;
  wire       [15:0]   _zz_9905;
  wire       [15:0]   _zz_9906;
  wire       [15:0]   _zz_9907;
  wire       [15:0]   _zz_9908;
  wire       [15:0]   _zz_9909;
  wire       [15:0]   _zz_9910;
  wire       [15:0]   _zz_9911;
  wire       [15:0]   _zz_9912;
  wire       [15:0]   _zz_9913;
  wire       [15:0]   _zz_9914;
  wire       [15:0]   _zz_9915;
  wire       [15:0]   _zz_9916;
  wire       [15:0]   _zz_9917;
  wire       [15:0]   _zz_9918;
  wire       [15:0]   _zz_9919;
  wire       [15:0]   _zz_9920;
  wire       [15:0]   _zz_9921;
  wire       [15:0]   _zz_9922;
  wire       [15:0]   _zz_9923;
  wire       [15:0]   _zz_9924;
  wire       [15:0]   _zz_9925;
  wire       [15:0]   _zz_9926;
  wire       [15:0]   _zz_9927;
  wire       [15:0]   _zz_9928;
  wire       [15:0]   _zz_9929;
  wire       [15:0]   _zz_9930;
  wire       [15:0]   _zz_9931;
  wire       [15:0]   _zz_9932;
  wire       [15:0]   _zz_9933;
  wire       [15:0]   _zz_9934;
  wire       [15:0]   _zz_9935;
  wire       [15:0]   _zz_9936;
  wire       [15:0]   _zz_9937;
  wire       [15:0]   _zz_9938;
  wire       [15:0]   _zz_9939;
  wire       [15:0]   _zz_9940;
  wire       [15:0]   _zz_9941;
  wire       [15:0]   _zz_9942;
  wire       [15:0]   _zz_9943;
  wire       [15:0]   _zz_9944;
  wire       [15:0]   _zz_9945;
  wire       [15:0]   _zz_9946;
  wire       [15:0]   _zz_9947;
  wire       [15:0]   _zz_9948;
  wire       [15:0]   _zz_9949;
  wire       [15:0]   _zz_9950;
  wire       [15:0]   _zz_9951;
  wire       [15:0]   _zz_9952;
  wire       [15:0]   _zz_9953;
  wire       [15:0]   _zz_9954;
  wire       [15:0]   _zz_9955;
  wire       [15:0]   _zz_9956;
  wire       [15:0]   _zz_9957;
  wire       [15:0]   _zz_9958;
  wire       [15:0]   _zz_9959;
  wire       [15:0]   _zz_9960;
  wire       [15:0]   _zz_9961;
  wire       [15:0]   _zz_9962;
  wire       [15:0]   _zz_9963;
  wire       [15:0]   _zz_9964;
  wire       [15:0]   _zz_9965;
  wire       [15:0]   _zz_9966;
  wire       [15:0]   _zz_9967;
  wire       [15:0]   _zz_9968;
  wire       [15:0]   _zz_9969;
  wire       [15:0]   _zz_9970;
  wire       [15:0]   _zz_9971;
  wire       [15:0]   _zz_9972;
  wire       [15:0]   _zz_9973;
  wire       [15:0]   _zz_9974;
  wire       [15:0]   _zz_9975;
  wire       [15:0]   _zz_9976;
  wire       [15:0]   _zz_9977;
  wire       [15:0]   _zz_9978;
  wire       [15:0]   _zz_9979;
  wire       [15:0]   _zz_9980;
  wire       [15:0]   _zz_9981;
  wire       [15:0]   _zz_9982;
  wire       [15:0]   _zz_9983;
  wire       [15:0]   _zz_9984;
  wire       [15:0]   _zz_9985;
  wire       [15:0]   _zz_9986;
  wire       [15:0]   _zz_9987;
  wire       [15:0]   _zz_9988;
  wire       [15:0]   _zz_9989;
  wire       [15:0]   _zz_9990;
  wire       [15:0]   _zz_9991;
  wire       [15:0]   _zz_9992;
  wire       [15:0]   _zz_9993;
  wire       [15:0]   _zz_9994;
  wire       [15:0]   _zz_9995;
  wire       [15:0]   _zz_9996;
  wire       [15:0]   _zz_9997;
  wire       [15:0]   _zz_9998;
  wire       [15:0]   _zz_9999;
  wire       [15:0]   _zz_10000;
  wire       [15:0]   _zz_10001;
  wire       [15:0]   _zz_10002;
  wire       [15:0]   _zz_10003;
  wire       [15:0]   _zz_10004;
  wire       [15:0]   _zz_10005;
  wire       [15:0]   _zz_10006;
  wire       [15:0]   _zz_10007;
  wire       [15:0]   _zz_10008;
  wire       [15:0]   _zz_10009;
  wire       [15:0]   _zz_10010;
  wire       [15:0]   _zz_10011;
  wire       [15:0]   _zz_10012;
  wire       [15:0]   _zz_10013;
  wire       [15:0]   _zz_10014;
  wire       [15:0]   _zz_10015;
  wire       [15:0]   _zz_10016;
  wire       [15:0]   _zz_10017;
  wire       [15:0]   _zz_10018;
  wire       [15:0]   _zz_10019;
  wire       [15:0]   _zz_10020;
  wire       [15:0]   _zz_10021;
  wire       [15:0]   _zz_10022;
  wire       [15:0]   _zz_10023;
  wire       [15:0]   _zz_10024;
  wire       [15:0]   _zz_10025;
  wire       [15:0]   _zz_10026;
  wire       [15:0]   _zz_10027;
  wire       [15:0]   _zz_10028;
  wire       [15:0]   _zz_10029;
  wire       [15:0]   _zz_10030;
  wire       [15:0]   _zz_10031;
  wire       [15:0]   _zz_10032;
  wire       [15:0]   _zz_10033;
  wire       [15:0]   _zz_10034;
  wire       [15:0]   _zz_10035;
  wire       [15:0]   _zz_10036;
  wire       [15:0]   _zz_10037;
  wire       [15:0]   _zz_10038;
  wire       [15:0]   _zz_10039;
  wire       [15:0]   _zz_10040;
  wire       [15:0]   _zz_10041;
  wire       [15:0]   _zz_10042;
  wire       [15:0]   _zz_10043;
  wire       [15:0]   _zz_10044;
  wire       [15:0]   _zz_10045;
  wire       [15:0]   _zz_10046;
  wire       [15:0]   _zz_10047;
  wire       [15:0]   _zz_10048;
  wire       [15:0]   _zz_10049;
  wire       [15:0]   _zz_10050;
  wire       [15:0]   _zz_10051;
  wire       [15:0]   _zz_10052;
  wire       [15:0]   _zz_10053;
  wire       [15:0]   _zz_10054;
  wire       [15:0]   _zz_10055;
  wire       [15:0]   _zz_10056;
  wire       [15:0]   _zz_10057;
  wire       [15:0]   _zz_10058;
  wire       [15:0]   _zz_10059;
  wire       [15:0]   _zz_10060;
  wire       [15:0]   _zz_10061;
  wire       [15:0]   _zz_10062;
  wire       [15:0]   _zz_10063;
  wire       [15:0]   _zz_10064;
  wire       [15:0]   _zz_10065;
  wire       [15:0]   _zz_10066;
  wire       [15:0]   _zz_10067;
  wire       [15:0]   _zz_10068;
  wire       [15:0]   _zz_10069;
  wire       [15:0]   _zz_10070;
  wire       [15:0]   _zz_10071;
  wire       [15:0]   _zz_10072;
  wire       [15:0]   _zz_10073;
  wire       [15:0]   _zz_10074;
  wire       [15:0]   _zz_10075;
  wire       [15:0]   _zz_10076;
  wire       [15:0]   _zz_10077;
  wire       [15:0]   _zz_10078;
  wire       [15:0]   _zz_10079;
  wire       [15:0]   _zz_10080;
  wire       [15:0]   _zz_10081;
  wire       [15:0]   _zz_10082;
  wire       [15:0]   _zz_10083;
  wire       [15:0]   _zz_10084;
  wire       [15:0]   _zz_10085;
  wire       [15:0]   _zz_10086;
  wire       [15:0]   _zz_10087;
  wire       [15:0]   _zz_10088;
  wire       [15:0]   _zz_10089;
  wire       [15:0]   _zz_10090;
  wire       [15:0]   _zz_10091;
  wire       [15:0]   _zz_10092;
  wire       [15:0]   _zz_10093;
  wire       [15:0]   _zz_10094;
  wire       [15:0]   _zz_10095;
  wire       [15:0]   _zz_10096;
  wire       [15:0]   _zz_10097;
  wire       [15:0]   _zz_10098;
  wire       [15:0]   _zz_10099;
  wire       [15:0]   _zz_10100;
  wire       [15:0]   _zz_10101;
  wire       [15:0]   _zz_10102;
  wire       [15:0]   _zz_10103;
  wire       [15:0]   _zz_10104;
  wire       [15:0]   _zz_10105;
  wire       [15:0]   _zz_10106;
  wire       [15:0]   _zz_10107;
  wire       [15:0]   _zz_10108;
  wire       [15:0]   _zz_10109;
  wire       [15:0]   _zz_10110;
  wire       [15:0]   _zz_10111;
  wire       [15:0]   _zz_10112;
  wire       [15:0]   _zz_10113;
  wire       [15:0]   _zz_10114;
  wire       [15:0]   _zz_10115;
  wire       [15:0]   _zz_10116;
  wire       [15:0]   _zz_10117;
  wire       [15:0]   _zz_10118;
  wire       [15:0]   _zz_10119;
  wire       [15:0]   _zz_10120;
  wire       [15:0]   _zz_10121;
  wire       [15:0]   _zz_10122;
  wire       [15:0]   _zz_10123;
  wire       [15:0]   _zz_10124;
  wire       [15:0]   _zz_10125;
  wire       [15:0]   _zz_10126;
  wire       [15:0]   _zz_10127;
  wire       [15:0]   _zz_10128;
  wire       [15:0]   _zz_10129;
  wire       [15:0]   _zz_10130;
  wire       [15:0]   _zz_10131;
  wire       [15:0]   _zz_10132;
  wire       [15:0]   _zz_10133;
  wire       [15:0]   _zz_10134;
  wire       [15:0]   _zz_10135;
  wire       [15:0]   _zz_10136;
  wire       [15:0]   _zz_10137;
  wire       [15:0]   _zz_10138;
  wire       [15:0]   _zz_10139;
  wire       [15:0]   _zz_10140;
  wire       [15:0]   _zz_10141;
  wire       [15:0]   _zz_10142;
  wire       [15:0]   _zz_10143;
  wire       [15:0]   _zz_10144;
  wire       [15:0]   _zz_10145;
  wire       [15:0]   _zz_10146;
  wire       [15:0]   _zz_10147;
  wire       [15:0]   _zz_10148;
  wire       [15:0]   _zz_10149;
  wire       [15:0]   _zz_10150;
  wire       [15:0]   _zz_10151;
  wire       [15:0]   _zz_10152;
  wire       [15:0]   _zz_10153;
  wire       [15:0]   _zz_10154;
  wire       [15:0]   _zz_10155;
  wire       [15:0]   _zz_10156;
  wire       [15:0]   _zz_10157;
  wire       [15:0]   _zz_10158;
  wire       [15:0]   _zz_10159;
  wire       [15:0]   _zz_10160;
  wire       [15:0]   _zz_10161;
  wire       [15:0]   _zz_10162;
  wire       [15:0]   _zz_10163;
  wire       [15:0]   _zz_10164;
  wire       [15:0]   _zz_10165;
  wire       [15:0]   _zz_10166;
  wire       [15:0]   _zz_10167;
  wire       [15:0]   _zz_10168;
  wire       [15:0]   _zz_10169;
  wire       [15:0]   _zz_10170;
  wire       [15:0]   _zz_10171;
  wire       [15:0]   _zz_10172;
  wire       [15:0]   _zz_10173;
  wire       [15:0]   _zz_10174;
  wire       [15:0]   _zz_10175;
  wire       [15:0]   _zz_10176;
  wire       [15:0]   _zz_10177;
  wire       [15:0]   _zz_10178;
  wire       [15:0]   _zz_10179;
  wire       [15:0]   _zz_10180;
  wire       [15:0]   _zz_10181;
  wire       [15:0]   _zz_10182;
  wire       [15:0]   _zz_10183;
  wire       [15:0]   _zz_10184;
  wire       [15:0]   _zz_10185;
  wire       [15:0]   _zz_10186;
  wire       [15:0]   _zz_10187;
  wire       [15:0]   _zz_10188;
  wire       [15:0]   _zz_10189;
  wire       [15:0]   _zz_10190;
  wire       [15:0]   _zz_10191;
  wire       [15:0]   _zz_10192;
  wire       [15:0]   _zz_10193;
  wire       [15:0]   _zz_10194;
  wire       [15:0]   _zz_10195;
  wire       [15:0]   _zz_10196;
  wire       [15:0]   _zz_10197;
  wire       [15:0]   _zz_10198;
  wire       [15:0]   _zz_10199;
  wire       [15:0]   _zz_10200;
  wire       [15:0]   _zz_10201;
  wire       [15:0]   _zz_10202;
  wire       [15:0]   _zz_10203;
  wire       [15:0]   _zz_10204;
  wire       [15:0]   _zz_10205;
  wire       [15:0]   _zz_10206;
  wire       [15:0]   _zz_10207;
  wire       [15:0]   _zz_10208;
  wire       [15:0]   _zz_10209;
  wire       [15:0]   _zz_10210;
  wire       [15:0]   _zz_10211;
  wire       [15:0]   _zz_10212;
  wire       [15:0]   _zz_10213;
  wire       [15:0]   _zz_10214;
  wire       [15:0]   _zz_10215;
  wire       [15:0]   _zz_10216;
  wire       [15:0]   _zz_10217;
  wire       [15:0]   _zz_10218;
  wire       [15:0]   _zz_10219;
  wire       [15:0]   _zz_10220;
  wire       [15:0]   _zz_10221;
  wire       [15:0]   _zz_10222;
  wire       [15:0]   _zz_10223;
  wire       [15:0]   _zz_10224;
  wire       [15:0]   _zz_10225;
  wire       [15:0]   _zz_10226;
  wire       [15:0]   _zz_10227;
  wire       [15:0]   _zz_10228;
  wire       [15:0]   _zz_10229;
  wire       [15:0]   _zz_10230;
  wire       [15:0]   _zz_10231;
  wire       [15:0]   _zz_10232;
  wire       [15:0]   _zz_10233;
  wire       [15:0]   _zz_10234;
  wire       [15:0]   _zz_10235;
  wire       [15:0]   _zz_10236;
  wire       [15:0]   _zz_10237;
  wire       [15:0]   _zz_10238;
  wire       [15:0]   _zz_10239;
  wire       [15:0]   _zz_10240;
  wire       [15:0]   _zz_10241;
  wire       [15:0]   _zz_10242;
  wire       [15:0]   _zz_10243;
  wire       [15:0]   _zz_10244;
  wire       [15:0]   _zz_10245;
  wire       [15:0]   _zz_10246;
  wire       [15:0]   _zz_10247;
  wire       [15:0]   _zz_10248;
  wire       [15:0]   _zz_10249;
  wire       [15:0]   _zz_10250;
  wire       [15:0]   _zz_10251;
  wire       [15:0]   _zz_10252;
  wire       [15:0]   _zz_10253;
  wire       [15:0]   _zz_10254;
  wire       [15:0]   _zz_10255;
  wire       [15:0]   _zz_10256;
  wire       [15:0]   _zz_10257;
  wire       [15:0]   _zz_10258;
  wire       [15:0]   _zz_10259;
  wire       [15:0]   _zz_10260;
  wire       [15:0]   _zz_10261;
  wire       [15:0]   _zz_10262;
  wire       [15:0]   _zz_10263;
  wire       [15:0]   _zz_10264;
  wire       [15:0]   _zz_10265;
  wire       [15:0]   _zz_10266;
  wire       [15:0]   _zz_10267;
  wire       [15:0]   _zz_10268;
  wire       [15:0]   _zz_10269;
  wire       [15:0]   _zz_10270;
  wire       [15:0]   _zz_10271;
  wire       [15:0]   _zz_10272;
  wire       [15:0]   _zz_10273;
  wire       [15:0]   _zz_10274;
  wire       [15:0]   _zz_10275;
  wire       [15:0]   _zz_10276;
  wire       [15:0]   _zz_10277;
  wire       [15:0]   _zz_10278;
  wire       [15:0]   _zz_10279;
  wire       [15:0]   _zz_10280;
  wire       [15:0]   _zz_10281;
  wire       [15:0]   _zz_10282;
  wire       [15:0]   _zz_10283;
  wire       [15:0]   _zz_10284;
  wire       [15:0]   _zz_10285;
  wire       [15:0]   _zz_10286;
  wire       [15:0]   _zz_10287;
  wire       [15:0]   _zz_10288;
  wire       [15:0]   _zz_10289;
  wire       [15:0]   _zz_10290;
  wire       [15:0]   _zz_10291;
  wire       [15:0]   _zz_10292;
  wire       [15:0]   _zz_10293;
  wire       [15:0]   _zz_10294;
  wire       [15:0]   _zz_10295;
  wire       [15:0]   _zz_10296;
  wire       [15:0]   _zz_10297;
  wire       [15:0]   _zz_10298;
  wire       [15:0]   _zz_10299;
  wire       [15:0]   _zz_10300;
  wire       [15:0]   _zz_10301;
  wire       [15:0]   _zz_10302;
  wire       [15:0]   _zz_10303;
  wire       [15:0]   _zz_10304;
  wire       [15:0]   _zz_10305;
  wire       [15:0]   _zz_10306;
  wire       [15:0]   _zz_10307;
  wire       [15:0]   _zz_10308;
  wire       [15:0]   _zz_10309;
  wire       [15:0]   _zz_10310;
  wire       [15:0]   _zz_10311;
  wire       [15:0]   _zz_10312;
  wire       [15:0]   _zz_10313;
  wire       [15:0]   _zz_10314;
  wire       [15:0]   _zz_10315;
  wire       [15:0]   _zz_10316;
  wire       [15:0]   _zz_10317;
  wire       [15:0]   _zz_10318;
  wire       [15:0]   _zz_10319;
  wire       [15:0]   _zz_10320;
  wire       [15:0]   _zz_10321;
  wire       [15:0]   _zz_10322;
  wire       [15:0]   _zz_10323;
  wire       [15:0]   _zz_10324;
  wire       [15:0]   _zz_10325;
  wire       [15:0]   _zz_10326;
  wire       [15:0]   _zz_10327;
  wire       [15:0]   _zz_10328;
  wire       [15:0]   _zz_10329;
  wire       [15:0]   _zz_10330;
  wire       [15:0]   _zz_10331;
  wire       [15:0]   _zz_10332;
  wire       [15:0]   _zz_10333;
  wire       [15:0]   _zz_10334;
  wire       [15:0]   _zz_10335;
  wire       [15:0]   _zz_10336;
  wire       [15:0]   _zz_10337;
  wire       [15:0]   _zz_10338;
  wire       [15:0]   _zz_10339;
  wire       [15:0]   _zz_10340;
  wire       [15:0]   _zz_10341;
  wire       [15:0]   _zz_10342;
  wire       [15:0]   _zz_10343;
  wire       [15:0]   _zz_10344;
  wire       [15:0]   _zz_10345;
  wire       [15:0]   _zz_10346;
  wire       [15:0]   _zz_10347;
  wire       [15:0]   _zz_10348;
  wire       [15:0]   _zz_10349;
  wire       [15:0]   _zz_10350;
  wire       [15:0]   _zz_10351;
  wire       [15:0]   _zz_10352;
  wire       [15:0]   _zz_10353;
  wire       [15:0]   _zz_10354;
  wire       [15:0]   _zz_10355;
  wire       [15:0]   _zz_10356;
  wire       [15:0]   _zz_10357;
  wire       [15:0]   _zz_10358;
  wire       [15:0]   _zz_10359;
  wire       [15:0]   _zz_10360;
  wire       [15:0]   _zz_10361;
  wire       [15:0]   _zz_10362;
  wire       [15:0]   _zz_10363;
  wire       [15:0]   _zz_10364;
  wire       [15:0]   _zz_10365;
  wire       [15:0]   _zz_10366;
  wire       [15:0]   _zz_10367;
  wire       [15:0]   _zz_10368;
  wire       [15:0]   _zz_10369;
  wire       [15:0]   _zz_10370;
  wire       [15:0]   _zz_10371;
  wire       [15:0]   _zz_10372;
  wire       [15:0]   _zz_10373;
  wire       [15:0]   _zz_10374;
  wire       [15:0]   _zz_10375;
  wire       [15:0]   _zz_10376;
  wire       [15:0]   _zz_10377;
  wire       [15:0]   _zz_10378;
  wire       [15:0]   _zz_10379;
  wire       [15:0]   _zz_10380;
  wire       [15:0]   _zz_10381;
  wire       [15:0]   _zz_10382;
  wire       [15:0]   _zz_10383;
  wire       [15:0]   _zz_10384;
  wire       [15:0]   _zz_10385;
  wire       [15:0]   _zz_10386;
  wire       [15:0]   _zz_10387;
  wire       [15:0]   _zz_10388;
  wire       [15:0]   _zz_10389;
  wire       [15:0]   _zz_10390;
  wire       [15:0]   _zz_10391;
  wire       [15:0]   _zz_10392;
  wire       [15:0]   _zz_10393;
  wire       [15:0]   _zz_10394;
  wire       [15:0]   _zz_10395;
  wire       [15:0]   _zz_10396;
  wire       [15:0]   _zz_10397;
  wire       [15:0]   _zz_10398;
  wire       [15:0]   _zz_10399;
  wire       [15:0]   _zz_10400;
  wire       [15:0]   _zz_10401;
  wire       [15:0]   _zz_10402;
  wire       [15:0]   _zz_10403;
  wire       [15:0]   _zz_10404;
  wire       [15:0]   _zz_10405;
  wire       [15:0]   _zz_10406;
  wire       [15:0]   _zz_10407;
  wire       [15:0]   _zz_10408;
  wire       [15:0]   _zz_10409;
  wire       [15:0]   _zz_10410;
  wire       [15:0]   _zz_10411;
  wire       [15:0]   _zz_10412;
  wire       [15:0]   _zz_10413;
  wire       [15:0]   _zz_10414;
  wire       [15:0]   _zz_10415;
  wire       [15:0]   _zz_10416;
  wire       [15:0]   _zz_10417;
  wire       [15:0]   _zz_10418;
  wire       [15:0]   _zz_10419;
  wire       [15:0]   _zz_10420;
  wire       [15:0]   _zz_10421;
  wire       [15:0]   _zz_10422;
  wire       [15:0]   _zz_10423;
  wire       [15:0]   _zz_10424;
  wire       [15:0]   _zz_10425;
  wire       [15:0]   _zz_10426;
  wire       [15:0]   _zz_10427;
  wire       [15:0]   _zz_10428;
  wire       [15:0]   _zz_10429;
  wire       [15:0]   _zz_10430;
  wire       [15:0]   _zz_10431;
  wire       [15:0]   _zz_10432;
  wire       [15:0]   _zz_10433;
  wire       [15:0]   _zz_10434;
  wire       [15:0]   _zz_10435;
  wire       [15:0]   _zz_10436;
  wire       [15:0]   _zz_10437;
  wire       [15:0]   _zz_10438;
  wire       [15:0]   _zz_10439;
  wire       [15:0]   _zz_10440;
  wire       [15:0]   _zz_10441;
  wire       [15:0]   _zz_10442;
  wire       [15:0]   _zz_10443;
  wire       [15:0]   _zz_10444;
  wire       [15:0]   _zz_10445;
  wire       [15:0]   _zz_10446;
  wire       [15:0]   _zz_10447;
  wire       [15:0]   _zz_10448;
  wire       [15:0]   _zz_10449;
  wire       [15:0]   _zz_10450;
  wire       [15:0]   _zz_10451;
  wire       [15:0]   _zz_10452;
  wire       [15:0]   _zz_10453;
  wire       [15:0]   _zz_10454;
  wire       [15:0]   _zz_10455;
  wire       [15:0]   _zz_10456;
  wire       [15:0]   _zz_10457;
  wire       [15:0]   _zz_10458;
  wire       [15:0]   _zz_10459;
  wire       [15:0]   _zz_10460;
  wire       [15:0]   _zz_10461;
  wire       [15:0]   _zz_10462;
  wire       [15:0]   _zz_10463;
  wire       [15:0]   _zz_10464;
  wire       [15:0]   _zz_10465;
  wire       [15:0]   _zz_10466;
  wire       [15:0]   _zz_10467;
  wire       [15:0]   _zz_10468;
  wire       [15:0]   _zz_10469;
  wire       [15:0]   _zz_10470;
  wire       [15:0]   _zz_10471;
  wire       [15:0]   _zz_10472;
  wire       [15:0]   _zz_10473;
  wire       [15:0]   _zz_10474;
  wire       [15:0]   _zz_10475;
  wire       [15:0]   _zz_10476;
  wire       [15:0]   _zz_10477;
  wire       [15:0]   _zz_10478;
  wire       [15:0]   _zz_10479;
  wire       [15:0]   _zz_10480;
  wire       [15:0]   _zz_10481;
  wire       [15:0]   _zz_10482;
  wire       [15:0]   _zz_10483;
  wire       [15:0]   _zz_10484;
  wire       [15:0]   _zz_10485;
  wire       [15:0]   _zz_10486;
  wire       [15:0]   _zz_10487;
  wire       [15:0]   _zz_10488;
  wire       [15:0]   _zz_10489;
  wire       [15:0]   _zz_10490;
  wire       [15:0]   _zz_10491;
  wire       [15:0]   _zz_10492;
  wire       [15:0]   _zz_10493;
  wire       [15:0]   _zz_10494;
  wire       [15:0]   _zz_10495;
  wire       [15:0]   _zz_10496;
  wire       [15:0]   _zz_10497;
  wire       [15:0]   _zz_10498;
  wire       [15:0]   _zz_10499;
  wire       [15:0]   _zz_10500;
  wire       [15:0]   _zz_10501;
  wire       [15:0]   _zz_10502;
  wire       [15:0]   _zz_10503;
  wire       [15:0]   _zz_10504;
  wire       [15:0]   _zz_10505;
  wire       [15:0]   _zz_10506;
  wire       [15:0]   _zz_10507;
  wire       [15:0]   _zz_10508;
  wire       [15:0]   _zz_10509;
  wire       [15:0]   _zz_10510;
  wire       [15:0]   _zz_10511;
  wire       [15:0]   _zz_10512;
  wire       [15:0]   _zz_10513;
  wire       [15:0]   _zz_10514;
  wire       [15:0]   _zz_10515;
  wire       [15:0]   _zz_10516;
  wire       [15:0]   _zz_10517;
  wire       [15:0]   _zz_10518;
  wire       [15:0]   _zz_10519;
  wire       [15:0]   _zz_10520;
  wire       [15:0]   _zz_10521;
  wire       [15:0]   _zz_10522;
  wire       [15:0]   _zz_10523;
  wire       [15:0]   _zz_10524;
  wire       [15:0]   _zz_10525;
  wire       [15:0]   _zz_10526;
  wire       [15:0]   _zz_10527;
  wire       [15:0]   _zz_10528;
  wire       [15:0]   _zz_10529;
  wire       [15:0]   _zz_10530;
  wire       [15:0]   _zz_10531;
  wire       [15:0]   _zz_10532;
  wire       [15:0]   _zz_10533;
  wire       [15:0]   _zz_10534;
  wire       [15:0]   _zz_10535;
  wire       [15:0]   _zz_10536;
  wire       [15:0]   _zz_10537;
  wire       [15:0]   _zz_10538;
  wire       [15:0]   _zz_10539;
  wire       [15:0]   _zz_10540;
  wire       [15:0]   _zz_10541;
  wire       [15:0]   _zz_10542;
  wire       [15:0]   _zz_10543;
  wire       [15:0]   _zz_10544;
  wire       [15:0]   _zz_10545;
  wire       [15:0]   _zz_10546;
  wire       [15:0]   _zz_10547;
  wire       [15:0]   _zz_10548;
  wire       [15:0]   _zz_10549;
  wire       [15:0]   _zz_10550;
  wire       [15:0]   _zz_10551;
  wire       [15:0]   _zz_10552;
  wire       [15:0]   _zz_10553;
  wire       [15:0]   _zz_10554;
  wire       [15:0]   _zz_10555;
  wire       [15:0]   _zz_10556;
  wire       [15:0]   _zz_10557;
  wire       [15:0]   _zz_10558;
  wire       [15:0]   _zz_10559;
  wire       [15:0]   _zz_10560;
  wire       [15:0]   _zz_10561;
  wire       [15:0]   _zz_10562;
  wire       [15:0]   _zz_10563;
  wire       [15:0]   _zz_10564;
  wire       [15:0]   _zz_10565;
  wire       [15:0]   _zz_10566;
  wire       [15:0]   _zz_10567;
  wire       [15:0]   _zz_10568;
  wire       [15:0]   _zz_10569;
  wire       [15:0]   _zz_10570;
  wire       [15:0]   _zz_10571;
  wire       [15:0]   _zz_10572;
  wire       [15:0]   _zz_10573;
  wire       [15:0]   _zz_10574;
  wire       [15:0]   _zz_10575;
  wire       [15:0]   _zz_10576;
  wire       [15:0]   _zz_10577;
  wire       [15:0]   _zz_10578;
  wire       [15:0]   _zz_10579;
  wire       [15:0]   _zz_10580;
  wire       [15:0]   _zz_10581;
  wire       [15:0]   _zz_10582;
  wire       [15:0]   _zz_10583;
  wire       [15:0]   _zz_10584;
  wire       [15:0]   _zz_10585;
  wire       [15:0]   _zz_10586;
  wire       [15:0]   _zz_10587;
  wire       [15:0]   _zz_10588;
  wire       [15:0]   _zz_10589;
  wire       [15:0]   _zz_10590;
  wire       [15:0]   _zz_10591;
  wire       [15:0]   _zz_10592;
  wire       [15:0]   _zz_10593;
  wire       [15:0]   _zz_10594;
  wire       [15:0]   _zz_10595;
  wire       [15:0]   _zz_10596;
  wire       [15:0]   _zz_10597;
  wire       [15:0]   _zz_10598;
  wire       [15:0]   _zz_10599;
  wire       [15:0]   _zz_10600;
  wire       [15:0]   _zz_10601;
  wire       [15:0]   _zz_10602;
  wire       [15:0]   _zz_10603;
  wire       [15:0]   _zz_10604;
  wire       [15:0]   _zz_10605;
  wire       [15:0]   _zz_10606;
  wire       [15:0]   _zz_10607;
  wire       [15:0]   _zz_10608;
  wire       [15:0]   _zz_10609;
  wire       [15:0]   _zz_10610;
  wire       [15:0]   _zz_10611;
  wire       [15:0]   _zz_10612;
  wire       [15:0]   _zz_10613;
  wire       [15:0]   _zz_10614;
  wire       [15:0]   _zz_10615;
  wire       [15:0]   _zz_10616;
  wire       [15:0]   _zz_10617;
  wire       [15:0]   _zz_10618;
  wire       [15:0]   _zz_10619;
  wire       [15:0]   _zz_10620;
  wire       [15:0]   _zz_10621;
  wire       [15:0]   _zz_10622;
  wire       [15:0]   _zz_10623;
  wire       [15:0]   _zz_10624;
  wire       [15:0]   _zz_10625;
  wire       [15:0]   _zz_10626;
  wire       [15:0]   _zz_10627;
  wire       [15:0]   _zz_10628;
  wire       [15:0]   _zz_10629;
  wire       [15:0]   _zz_10630;
  wire       [15:0]   _zz_10631;
  wire       [15:0]   _zz_10632;
  wire       [15:0]   _zz_10633;
  wire       [15:0]   _zz_10634;
  wire       [15:0]   _zz_10635;
  wire       [15:0]   _zz_10636;
  wire       [15:0]   _zz_10637;
  wire       [15:0]   _zz_10638;
  wire       [15:0]   _zz_10639;
  wire       [15:0]   _zz_10640;
  wire       [15:0]   _zz_10641;
  wire       [15:0]   _zz_10642;
  wire       [15:0]   _zz_10643;
  wire       [15:0]   _zz_10644;
  wire       [15:0]   _zz_10645;
  wire       [15:0]   _zz_10646;
  wire       [15:0]   _zz_10647;
  wire       [15:0]   _zz_10648;
  wire       [15:0]   _zz_10649;
  wire       [15:0]   _zz_10650;
  wire       [15:0]   _zz_10651;
  wire       [15:0]   _zz_10652;
  wire       [15:0]   _zz_10653;
  wire       [15:0]   _zz_10654;
  wire       [15:0]   _zz_10655;
  wire       [15:0]   _zz_10656;
  wire       [15:0]   _zz_10657;
  wire       [15:0]   _zz_10658;
  wire       [15:0]   _zz_10659;
  wire       [15:0]   _zz_10660;
  wire       [15:0]   _zz_10661;
  wire       [15:0]   _zz_10662;
  wire       [15:0]   _zz_10663;
  wire       [15:0]   _zz_10664;
  wire       [15:0]   _zz_10665;
  wire       [15:0]   _zz_10666;
  wire       [15:0]   _zz_10667;
  wire       [15:0]   _zz_10668;
  wire       [15:0]   _zz_10669;
  wire       [15:0]   _zz_10670;
  wire       [15:0]   _zz_10671;
  wire       [15:0]   _zz_10672;
  wire       [15:0]   _zz_10673;
  wire       [15:0]   _zz_10674;
  wire       [15:0]   _zz_10675;
  wire       [15:0]   _zz_10676;
  wire       [15:0]   _zz_10677;
  wire       [15:0]   _zz_10678;
  wire       [15:0]   _zz_10679;
  wire       [15:0]   _zz_10680;
  wire       [15:0]   _zz_10681;
  wire       [15:0]   _zz_10682;
  wire       [15:0]   _zz_10683;
  wire       [15:0]   _zz_10684;
  wire       [15:0]   _zz_10685;
  wire       [15:0]   _zz_10686;
  wire       [15:0]   _zz_10687;
  wire       [15:0]   _zz_10688;
  wire       [15:0]   _zz_10689;
  wire       [15:0]   _zz_10690;
  wire       [15:0]   _zz_10691;
  wire       [15:0]   _zz_10692;
  wire       [15:0]   _zz_10693;
  wire       [15:0]   _zz_10694;
  wire       [15:0]   _zz_10695;
  wire       [15:0]   _zz_10696;
  wire       [15:0]   _zz_10697;
  wire       [15:0]   _zz_10698;
  wire       [15:0]   _zz_10699;
  wire       [15:0]   _zz_10700;
  wire       [15:0]   _zz_10701;
  wire       [15:0]   _zz_10702;
  wire       [15:0]   _zz_10703;
  wire       [15:0]   _zz_10704;
  wire       [15:0]   _zz_10705;
  wire       [15:0]   _zz_10706;
  wire       [15:0]   _zz_10707;
  wire       [15:0]   _zz_10708;
  wire       [15:0]   _zz_10709;
  wire       [15:0]   _zz_10710;
  wire       [15:0]   _zz_10711;
  wire       [15:0]   _zz_10712;
  wire       [15:0]   _zz_10713;
  wire       [15:0]   _zz_10714;
  wire       [15:0]   _zz_10715;
  wire       [15:0]   _zz_10716;
  wire       [15:0]   _zz_10717;
  wire       [15:0]   _zz_10718;
  wire       [15:0]   _zz_10719;
  wire       [15:0]   _zz_10720;
  wire       [15:0]   _zz_10721;
  wire       [15:0]   _zz_10722;
  wire       [15:0]   _zz_10723;
  wire       [15:0]   _zz_10724;
  wire       [15:0]   _zz_10725;
  wire       [15:0]   _zz_10726;
  wire       [15:0]   _zz_10727;
  wire       [15:0]   _zz_10728;
  wire       [15:0]   _zz_10729;
  wire       [15:0]   _zz_10730;
  wire       [15:0]   _zz_10731;
  wire       [15:0]   _zz_10732;
  wire       [15:0]   _zz_10733;
  wire       [15:0]   _zz_10734;
  wire       [15:0]   _zz_10735;
  wire       [15:0]   _zz_10736;
  wire       [15:0]   _zz_10737;
  wire       [15:0]   _zz_10738;
  wire       [15:0]   _zz_10739;
  wire       [15:0]   _zz_10740;
  wire       [15:0]   _zz_10741;
  wire       [15:0]   _zz_10742;
  wire       [15:0]   _zz_10743;
  wire       [15:0]   _zz_10744;
  wire       [15:0]   _zz_10745;
  wire       [15:0]   _zz_10746;
  wire       [15:0]   _zz_10747;
  wire       [15:0]   _zz_10748;
  wire       [15:0]   _zz_10749;
  wire       [15:0]   _zz_10750;
  wire       [15:0]   _zz_10751;
  wire       [15:0]   _zz_10752;
  wire       [15:0]   _zz_10753;
  wire       [15:0]   _zz_10754;
  wire       [15:0]   _zz_10755;
  wire       [15:0]   _zz_10756;
  wire       [15:0]   _zz_10757;
  wire       [15:0]   _zz_10758;
  wire       [15:0]   _zz_10759;
  wire       [15:0]   _zz_10760;
  wire       [15:0]   _zz_10761;
  wire       [15:0]   _zz_10762;
  wire       [15:0]   _zz_10763;
  wire       [15:0]   _zz_10764;
  wire       [15:0]   _zz_10765;
  wire       [15:0]   _zz_10766;
  wire       [15:0]   _zz_10767;
  wire       [15:0]   _zz_10768;
  wire       [15:0]   _zz_10769;
  wire       [15:0]   _zz_10770;
  wire       [15:0]   _zz_10771;
  wire       [15:0]   _zz_10772;
  wire       [15:0]   _zz_10773;
  wire       [15:0]   _zz_10774;
  wire       [15:0]   _zz_10775;
  wire       [15:0]   _zz_10776;
  wire       [15:0]   _zz_10777;
  wire       [15:0]   _zz_10778;
  wire       [15:0]   _zz_10779;
  wire       [15:0]   _zz_10780;
  wire       [15:0]   _zz_10781;
  wire       [15:0]   _zz_10782;
  wire       [15:0]   _zz_10783;
  wire       [15:0]   _zz_10784;
  wire       [15:0]   _zz_10785;
  wire       [15:0]   _zz_10786;
  wire       [15:0]   _zz_10787;
  wire       [15:0]   _zz_10788;
  wire       [15:0]   _zz_10789;
  wire       [15:0]   _zz_10790;
  wire       [15:0]   _zz_10791;
  wire       [15:0]   _zz_10792;
  wire       [15:0]   _zz_10793;
  wire       [15:0]   _zz_10794;
  wire       [15:0]   _zz_10795;
  wire       [15:0]   _zz_10796;
  wire       [15:0]   _zz_10797;
  wire       [15:0]   _zz_10798;
  wire       [15:0]   _zz_10799;
  wire       [15:0]   _zz_10800;
  wire       [15:0]   _zz_10801;
  wire       [15:0]   _zz_10802;
  wire       [15:0]   _zz_10803;
  wire       [15:0]   _zz_10804;
  wire       [15:0]   _zz_10805;
  wire       [15:0]   _zz_10806;
  wire       [15:0]   _zz_10807;
  wire       [15:0]   _zz_10808;
  wire       [15:0]   _zz_10809;
  wire       [15:0]   _zz_10810;
  wire       [15:0]   _zz_10811;
  wire       [15:0]   _zz_10812;
  wire       [15:0]   _zz_10813;
  wire       [15:0]   _zz_10814;
  wire       [15:0]   _zz_10815;
  wire       [15:0]   _zz_10816;
  wire       [15:0]   _zz_10817;
  wire       [15:0]   _zz_10818;
  wire       [15:0]   _zz_10819;
  wire       [15:0]   _zz_10820;
  wire       [15:0]   _zz_10821;
  wire       [15:0]   _zz_10822;
  wire       [15:0]   _zz_10823;
  wire       [15:0]   _zz_10824;
  wire       [15:0]   _zz_10825;
  wire       [15:0]   _zz_10826;
  wire       [15:0]   _zz_10827;
  wire       [15:0]   _zz_10828;
  wire       [15:0]   _zz_10829;
  wire       [15:0]   _zz_10830;
  wire       [15:0]   _zz_10831;
  wire       [15:0]   _zz_10832;
  wire       [15:0]   _zz_10833;
  wire       [15:0]   _zz_10834;
  wire       [15:0]   _zz_10835;
  wire       [15:0]   _zz_10836;
  wire       [15:0]   _zz_10837;
  wire       [15:0]   _zz_10838;
  wire       [15:0]   _zz_10839;
  wire       [15:0]   _zz_10840;
  wire       [15:0]   _zz_10841;
  wire       [15:0]   _zz_10842;
  wire       [15:0]   _zz_10843;
  wire       [15:0]   _zz_10844;
  wire       [15:0]   _zz_10845;
  wire       [15:0]   _zz_10846;
  wire       [15:0]   _zz_10847;
  wire       [15:0]   _zz_10848;
  wire       [15:0]   _zz_10849;
  wire       [15:0]   _zz_10850;
  wire       [15:0]   _zz_10851;
  wire       [15:0]   _zz_10852;
  wire       [15:0]   _zz_10853;
  wire       [15:0]   _zz_10854;
  wire       [15:0]   _zz_10855;
  wire       [15:0]   _zz_10856;
  wire       [15:0]   _zz_10857;
  wire       [15:0]   _zz_10858;
  wire       [15:0]   _zz_10859;
  wire       [15:0]   _zz_10860;
  wire       [15:0]   _zz_10861;
  wire       [15:0]   _zz_10862;
  wire       [15:0]   _zz_10863;
  wire       [15:0]   _zz_10864;
  wire       [15:0]   _zz_10865;
  wire       [15:0]   _zz_10866;
  wire       [15:0]   _zz_10867;
  wire       [15:0]   _zz_10868;
  wire       [15:0]   _zz_10869;
  wire       [15:0]   _zz_10870;
  wire       [15:0]   _zz_10871;
  wire       [15:0]   _zz_10872;
  wire       [15:0]   _zz_10873;
  wire       [15:0]   _zz_10874;
  wire       [15:0]   _zz_10875;
  wire       [15:0]   _zz_10876;
  wire       [15:0]   _zz_10877;
  wire       [15:0]   _zz_10878;
  wire       [15:0]   _zz_10879;
  wire       [15:0]   _zz_10880;
  wire       [15:0]   _zz_10881;
  wire       [15:0]   _zz_10882;
  wire       [15:0]   _zz_10883;
  wire       [15:0]   _zz_10884;
  wire       [15:0]   _zz_10885;
  wire       [15:0]   _zz_10886;
  wire       [15:0]   _zz_10887;
  wire       [15:0]   _zz_10888;
  wire       [15:0]   _zz_10889;
  wire       [15:0]   _zz_10890;
  wire       [15:0]   _zz_10891;
  wire       [15:0]   _zz_10892;
  wire       [15:0]   _zz_10893;
  wire       [15:0]   _zz_10894;
  wire       [15:0]   _zz_10895;
  wire       [15:0]   _zz_10896;
  wire       [15:0]   _zz_10897;
  wire       [15:0]   _zz_10898;
  wire       [15:0]   _zz_10899;
  wire       [15:0]   _zz_10900;
  wire       [15:0]   _zz_10901;
  wire       [15:0]   _zz_10902;
  wire       [15:0]   _zz_10903;
  wire       [15:0]   _zz_10904;
  wire       [15:0]   _zz_10905;
  wire       [15:0]   _zz_10906;
  wire       [15:0]   _zz_10907;
  wire       [15:0]   _zz_10908;
  wire       [15:0]   _zz_10909;
  wire       [15:0]   _zz_10910;
  wire       [15:0]   _zz_10911;
  wire       [15:0]   _zz_10912;
  wire       [15:0]   _zz_10913;
  wire       [15:0]   _zz_10914;
  wire       [15:0]   _zz_10915;
  wire       [15:0]   _zz_10916;
  wire       [15:0]   _zz_10917;
  wire       [15:0]   _zz_10918;
  wire       [15:0]   _zz_10919;
  wire       [15:0]   _zz_10920;
  wire       [15:0]   _zz_10921;
  wire       [15:0]   _zz_10922;
  wire       [15:0]   _zz_10923;
  wire       [15:0]   _zz_10924;
  wire       [15:0]   _zz_10925;
  wire       [15:0]   _zz_10926;
  wire       [15:0]   _zz_10927;
  wire       [15:0]   _zz_10928;
  wire       [15:0]   _zz_10929;
  wire       [15:0]   _zz_10930;
  wire       [15:0]   _zz_10931;
  wire       [15:0]   _zz_10932;
  wire       [15:0]   _zz_10933;
  wire       [15:0]   _zz_10934;
  wire       [15:0]   _zz_10935;
  wire       [15:0]   _zz_10936;
  wire       [15:0]   _zz_10937;
  wire       [15:0]   _zz_10938;
  wire       [15:0]   _zz_10939;
  wire       [15:0]   _zz_10940;
  wire       [15:0]   _zz_10941;
  wire       [15:0]   _zz_10942;
  wire       [15:0]   _zz_10943;
  wire       [15:0]   _zz_10944;
  wire       [15:0]   _zz_10945;
  wire       [15:0]   _zz_10946;
  wire       [15:0]   _zz_10947;
  wire       [15:0]   _zz_10948;
  wire       [15:0]   _zz_10949;
  wire       [15:0]   _zz_10950;
  wire       [15:0]   _zz_10951;
  wire       [15:0]   _zz_10952;
  wire       [15:0]   _zz_10953;
  wire       [15:0]   _zz_10954;
  wire       [15:0]   _zz_10955;
  wire       [15:0]   _zz_10956;
  wire       [15:0]   _zz_10957;
  wire       [15:0]   _zz_10958;
  wire       [15:0]   _zz_10959;
  wire       [15:0]   _zz_10960;
  wire       [15:0]   _zz_10961;
  wire       [15:0]   _zz_10962;
  wire       [15:0]   _zz_10963;
  wire       [15:0]   _zz_10964;
  wire       [15:0]   _zz_10965;
  wire       [15:0]   _zz_10966;
  wire       [15:0]   _zz_10967;
  wire       [15:0]   _zz_10968;
  wire       [15:0]   _zz_10969;
  wire       [15:0]   _zz_10970;
  wire       [15:0]   _zz_10971;
  wire       [15:0]   _zz_10972;
  wire       [15:0]   _zz_10973;
  wire       [15:0]   _zz_10974;
  wire       [15:0]   _zz_10975;
  wire       [15:0]   _zz_10976;
  wire       [15:0]   _zz_10977;
  wire       [15:0]   _zz_10978;
  wire       [15:0]   _zz_10979;
  wire       [15:0]   _zz_10980;
  wire       [15:0]   _zz_10981;
  wire       [15:0]   _zz_10982;
  wire       [15:0]   _zz_10983;
  wire       [15:0]   _zz_10984;
  wire       [15:0]   _zz_10985;
  wire       [15:0]   _zz_10986;
  wire       [15:0]   _zz_10987;
  wire       [15:0]   _zz_10988;
  wire       [15:0]   _zz_10989;
  wire       [15:0]   _zz_10990;
  wire       [15:0]   _zz_10991;
  wire       [15:0]   _zz_10992;
  wire       [15:0]   _zz_10993;
  wire       [15:0]   _zz_10994;
  wire       [15:0]   _zz_10995;
  wire       [15:0]   _zz_10996;
  wire       [15:0]   _zz_10997;
  wire       [15:0]   _zz_10998;
  wire       [15:0]   _zz_10999;
  wire       [15:0]   _zz_11000;
  wire       [15:0]   _zz_11001;
  wire       [15:0]   _zz_11002;
  wire       [15:0]   _zz_11003;
  wire       [15:0]   _zz_11004;
  wire       [15:0]   _zz_11005;
  wire       [15:0]   _zz_11006;
  wire       [15:0]   _zz_11007;
  wire       [15:0]   _zz_11008;
  wire       [15:0]   _zz_11009;
  wire       [15:0]   _zz_11010;
  wire       [15:0]   _zz_11011;
  wire       [15:0]   _zz_11012;
  wire       [15:0]   _zz_11013;
  wire       [15:0]   _zz_11014;
  wire       [15:0]   _zz_11015;
  wire       [15:0]   _zz_11016;
  wire       [15:0]   _zz_11017;
  wire       [15:0]   _zz_11018;
  wire       [15:0]   _zz_11019;
  wire       [15:0]   _zz_11020;
  wire       [15:0]   _zz_11021;
  wire       [15:0]   _zz_11022;
  wire       [15:0]   _zz_11023;
  wire       [15:0]   _zz_11024;
  wire       [15:0]   _zz_11025;
  wire       [15:0]   _zz_11026;
  wire       [15:0]   _zz_11027;
  wire       [15:0]   _zz_11028;
  wire       [15:0]   _zz_11029;
  wire       [15:0]   _zz_11030;
  wire       [15:0]   _zz_11031;
  wire       [15:0]   _zz_11032;
  wire       [15:0]   _zz_11033;
  wire       [15:0]   _zz_11034;
  wire       [15:0]   _zz_11035;
  wire       [15:0]   _zz_11036;
  wire       [15:0]   _zz_11037;
  wire       [15:0]   _zz_11038;
  wire       [15:0]   _zz_11039;
  wire       [15:0]   _zz_11040;
  wire       [15:0]   _zz_11041;
  wire       [15:0]   _zz_11042;
  wire       [15:0]   _zz_11043;
  wire       [15:0]   _zz_11044;
  wire       [15:0]   _zz_11045;
  wire       [15:0]   _zz_11046;
  wire       [15:0]   _zz_11047;
  wire       [15:0]   _zz_11048;
  wire       [15:0]   _zz_11049;
  wire       [15:0]   _zz_11050;
  wire       [15:0]   _zz_11051;
  wire       [15:0]   _zz_11052;
  wire       [15:0]   _zz_11053;
  wire       [15:0]   _zz_11054;
  wire       [15:0]   _zz_11055;
  wire       [15:0]   _zz_11056;
  wire       [15:0]   _zz_11057;
  wire       [15:0]   _zz_11058;
  wire       [15:0]   _zz_11059;
  wire       [15:0]   _zz_11060;
  wire       [15:0]   _zz_11061;
  wire       [15:0]   _zz_11062;
  wire       [15:0]   _zz_11063;
  wire       [15:0]   _zz_11064;
  wire       [15:0]   _zz_11065;
  wire       [15:0]   _zz_11066;
  wire       [15:0]   _zz_11067;
  wire       [15:0]   _zz_11068;
  wire       [15:0]   _zz_11069;
  wire       [15:0]   _zz_11070;
  wire       [15:0]   _zz_11071;
  wire       [15:0]   _zz_11072;
  wire       [15:0]   _zz_11073;
  wire       [15:0]   _zz_11074;
  wire       [15:0]   _zz_11075;
  wire       [15:0]   _zz_11076;
  wire       [15:0]   _zz_11077;
  wire       [15:0]   _zz_11078;
  wire       [15:0]   _zz_11079;
  wire       [15:0]   _zz_11080;
  wire       [15:0]   _zz_11081;
  wire       [15:0]   _zz_11082;
  wire       [15:0]   _zz_11083;
  wire       [15:0]   _zz_11084;
  wire       [15:0]   _zz_11085;
  wire       [15:0]   _zz_11086;
  wire       [15:0]   _zz_11087;
  wire       [15:0]   _zz_11088;
  wire       [15:0]   _zz_11089;
  wire       [15:0]   _zz_11090;
  wire       [15:0]   _zz_11091;
  wire       [15:0]   _zz_11092;
  wire       [15:0]   _zz_11093;
  wire       [15:0]   _zz_11094;
  wire       [15:0]   _zz_11095;
  wire       [15:0]   _zz_11096;
  wire       [15:0]   _zz_11097;
  wire       [15:0]   _zz_11098;
  wire       [15:0]   _zz_11099;
  wire       [15:0]   _zz_11100;
  wire       [15:0]   _zz_11101;
  wire       [15:0]   _zz_11102;
  wire       [15:0]   _zz_11103;
  wire       [15:0]   _zz_11104;
  wire       [15:0]   _zz_11105;
  wire       [15:0]   _zz_11106;
  wire       [15:0]   _zz_11107;
  wire       [15:0]   _zz_11108;
  wire       [15:0]   _zz_11109;
  wire       [15:0]   _zz_11110;
  wire       [15:0]   _zz_11111;
  wire       [15:0]   _zz_11112;
  wire       [15:0]   _zz_11113;
  wire       [15:0]   _zz_11114;
  wire       [15:0]   _zz_11115;
  wire       [15:0]   _zz_11116;
  wire       [15:0]   _zz_11117;
  wire       [15:0]   _zz_11118;
  wire       [15:0]   _zz_11119;
  wire       [15:0]   _zz_11120;
  wire       [15:0]   _zz_11121;
  wire       [15:0]   _zz_11122;
  wire       [15:0]   _zz_11123;
  wire       [15:0]   _zz_11124;
  wire       [15:0]   _zz_11125;
  wire       [15:0]   _zz_11126;
  wire       [15:0]   _zz_11127;
  wire       [15:0]   _zz_11128;
  wire       [15:0]   _zz_11129;
  wire       [15:0]   _zz_11130;
  wire       [15:0]   _zz_11131;
  wire       [15:0]   _zz_11132;
  wire       [15:0]   _zz_11133;
  wire       [15:0]   _zz_11134;
  wire       [15:0]   _zz_11135;
  wire       [15:0]   _zz_11136;
  wire       [15:0]   _zz_11137;
  wire       [15:0]   _zz_11138;
  wire       [15:0]   _zz_11139;
  wire       [15:0]   _zz_11140;
  wire       [15:0]   _zz_11141;
  wire       [15:0]   _zz_11142;
  wire       [15:0]   _zz_11143;
  wire       [15:0]   _zz_11144;
  wire       [15:0]   _zz_11145;
  wire       [15:0]   _zz_11146;
  wire       [15:0]   _zz_11147;
  wire       [15:0]   _zz_11148;
  wire       [15:0]   _zz_11149;
  wire       [15:0]   _zz_11150;
  wire       [15:0]   _zz_11151;
  wire       [15:0]   _zz_11152;
  wire       [15:0]   _zz_11153;
  wire       [15:0]   _zz_11154;
  wire       [15:0]   _zz_11155;
  wire       [15:0]   _zz_11156;
  wire       [15:0]   _zz_11157;
  wire       [15:0]   _zz_11158;
  wire       [15:0]   _zz_11159;
  wire       [15:0]   _zz_11160;
  wire       [15:0]   _zz_11161;
  wire       [15:0]   _zz_11162;
  wire       [15:0]   _zz_11163;
  wire       [15:0]   _zz_11164;
  wire       [15:0]   _zz_11165;
  wire       [15:0]   _zz_11166;
  wire       [15:0]   _zz_11167;
  wire       [15:0]   _zz_11168;
  wire       [15:0]   _zz_11169;
  wire       [15:0]   _zz_11170;
  wire       [15:0]   _zz_11171;
  wire       [15:0]   _zz_11172;
  wire       [15:0]   _zz_11173;
  wire       [15:0]   _zz_11174;
  wire       [15:0]   _zz_11175;
  wire       [15:0]   _zz_11176;
  wire       [15:0]   _zz_11177;
  wire       [15:0]   _zz_11178;
  wire       [15:0]   _zz_11179;
  wire       [15:0]   _zz_11180;
  wire       [15:0]   _zz_11181;
  wire       [15:0]   _zz_11182;
  wire       [15:0]   _zz_11183;
  wire       [15:0]   _zz_11184;
  wire       [15:0]   _zz_11185;
  wire       [15:0]   _zz_11186;
  wire       [15:0]   _zz_11187;
  wire       [15:0]   _zz_11188;
  wire       [15:0]   _zz_11189;
  wire       [15:0]   _zz_11190;
  wire       [15:0]   _zz_11191;
  wire       [15:0]   _zz_11192;
  wire       [15:0]   _zz_11193;
  wire       [15:0]   _zz_11194;
  wire       [15:0]   _zz_11195;
  wire       [15:0]   _zz_11196;
  wire       [15:0]   _zz_11197;
  wire       [15:0]   _zz_11198;
  wire       [15:0]   _zz_11199;
  wire       [15:0]   _zz_11200;
  wire       [15:0]   _zz_11201;
  wire       [15:0]   _zz_11202;
  wire       [15:0]   _zz_11203;
  wire       [15:0]   _zz_11204;
  wire       [15:0]   _zz_11205;
  wire       [15:0]   _zz_11206;
  wire       [15:0]   _zz_11207;
  wire       [15:0]   _zz_11208;
  wire       [15:0]   _zz_11209;
  wire       [15:0]   _zz_11210;
  wire       [15:0]   _zz_11211;
  wire       [15:0]   _zz_11212;
  wire       [15:0]   _zz_11213;
  wire       [15:0]   _zz_11214;
  wire       [15:0]   _zz_11215;
  wire       [15:0]   _zz_11216;
  wire       [15:0]   _zz_11217;
  wire       [15:0]   _zz_11218;
  wire       [15:0]   _zz_11219;
  wire       [15:0]   _zz_11220;
  wire       [15:0]   _zz_11221;
  wire       [15:0]   _zz_11222;
  wire       [15:0]   _zz_11223;
  wire       [15:0]   _zz_11224;
  wire       [15:0]   _zz_11225;
  wire       [15:0]   _zz_11226;
  wire       [15:0]   _zz_11227;
  wire       [15:0]   _zz_11228;
  wire       [15:0]   _zz_11229;
  wire       [15:0]   _zz_11230;
  wire       [15:0]   _zz_11231;
  wire       [15:0]   _zz_11232;
  wire       [15:0]   _zz_11233;
  wire       [15:0]   _zz_11234;
  wire       [15:0]   _zz_11235;
  wire       [15:0]   _zz_11236;
  wire       [15:0]   _zz_11237;
  wire       [15:0]   _zz_11238;
  wire       [15:0]   _zz_11239;
  wire       [15:0]   _zz_11240;
  wire       [15:0]   _zz_11241;
  wire       [15:0]   _zz_11242;
  wire       [15:0]   _zz_11243;
  wire       [15:0]   _zz_11244;
  wire       [15:0]   _zz_11245;
  wire       [15:0]   _zz_11246;
  wire       [15:0]   _zz_11247;
  wire       [15:0]   _zz_11248;
  wire       [15:0]   _zz_11249;
  wire       [15:0]   _zz_11250;
  wire       [15:0]   _zz_11251;
  wire       [15:0]   _zz_11252;
  wire       [15:0]   _zz_11253;
  wire       [15:0]   _zz_11254;
  wire       [15:0]   _zz_11255;
  wire       [15:0]   _zz_11256;
  wire       [15:0]   _zz_11257;
  wire       [15:0]   _zz_11258;
  wire       [15:0]   _zz_11259;
  wire       [15:0]   _zz_11260;
  wire       [15:0]   _zz_11261;
  wire       [15:0]   _zz_11262;
  wire       [15:0]   _zz_11263;
  wire       [15:0]   _zz_11264;
  wire       [15:0]   _zz_11265;
  wire       [15:0]   _zz_11266;
  wire       [15:0]   _zz_11267;
  wire       [15:0]   _zz_11268;
  wire       [15:0]   _zz_11269;
  wire       [15:0]   _zz_11270;
  wire       [15:0]   _zz_11271;
  wire       [15:0]   _zz_11272;
  wire       [15:0]   _zz_11273;
  wire       [15:0]   _zz_11274;
  wire       [15:0]   _zz_11275;
  wire       [15:0]   _zz_11276;
  wire       [15:0]   _zz_11277;
  wire       [15:0]   _zz_11278;
  wire       [15:0]   _zz_11279;
  wire       [15:0]   _zz_11280;
  wire       [15:0]   _zz_11281;
  wire       [15:0]   _zz_11282;
  wire       [15:0]   _zz_11283;
  wire       [15:0]   _zz_11284;
  wire       [15:0]   _zz_11285;
  wire       [15:0]   _zz_11286;
  wire       [15:0]   _zz_11287;
  wire       [15:0]   _zz_11288;
  wire       [15:0]   _zz_11289;
  wire       [15:0]   _zz_11290;
  wire       [15:0]   _zz_11291;
  wire       [15:0]   _zz_11292;
  wire       [15:0]   _zz_11293;
  wire       [15:0]   _zz_11294;
  wire       [15:0]   _zz_11295;
  wire       [15:0]   _zz_11296;
  wire       [15:0]   _zz_11297;
  wire       [15:0]   _zz_11298;
  wire       [15:0]   _zz_11299;
  wire       [15:0]   _zz_11300;
  wire       [15:0]   _zz_11301;
  wire       [15:0]   _zz_11302;
  wire       [15:0]   _zz_11303;
  wire       [15:0]   _zz_11304;
  wire       [15:0]   _zz_11305;
  wire       [15:0]   _zz_11306;
  wire       [15:0]   _zz_11307;
  wire       [15:0]   _zz_11308;
  wire       [15:0]   _zz_11309;
  wire       [15:0]   _zz_11310;
  wire       [15:0]   _zz_11311;
  wire       [15:0]   _zz_11312;
  wire       [15:0]   _zz_11313;
  wire       [15:0]   _zz_11314;
  wire       [15:0]   _zz_11315;
  wire       [15:0]   _zz_11316;
  wire       [15:0]   _zz_11317;
  wire       [15:0]   _zz_11318;
  wire       [15:0]   _zz_11319;
  wire       [15:0]   _zz_11320;
  wire       [15:0]   _zz_11321;
  wire       [15:0]   _zz_11322;
  wire       [15:0]   _zz_11323;
  wire       [15:0]   _zz_11324;
  wire       [15:0]   _zz_11325;
  wire       [15:0]   _zz_11326;
  wire       [15:0]   _zz_11327;
  wire       [15:0]   _zz_11328;
  wire       [15:0]   _zz_11329;
  wire       [15:0]   _zz_11330;
  wire       [15:0]   _zz_11331;
  wire       [15:0]   _zz_11332;
  wire       [15:0]   _zz_11333;
  wire       [15:0]   _zz_11334;
  wire       [15:0]   _zz_11335;
  wire       [15:0]   _zz_11336;
  wire       [15:0]   _zz_11337;
  wire       [15:0]   _zz_11338;
  wire       [15:0]   _zz_11339;
  wire       [15:0]   _zz_11340;
  wire       [15:0]   _zz_11341;
  wire       [15:0]   _zz_11342;
  wire       [15:0]   _zz_11343;
  wire       [15:0]   _zz_11344;
  wire       [15:0]   _zz_11345;
  wire       [15:0]   _zz_11346;
  wire       [15:0]   _zz_11347;
  wire       [15:0]   _zz_11348;
  wire       [15:0]   _zz_11349;
  wire       [15:0]   _zz_11350;
  wire       [15:0]   _zz_11351;
  wire       [15:0]   _zz_11352;
  wire       [15:0]   _zz_11353;
  wire       [15:0]   _zz_11354;
  wire       [15:0]   _zz_11355;
  wire       [15:0]   _zz_11356;
  wire       [15:0]   _zz_11357;
  wire       [15:0]   _zz_11358;
  wire       [15:0]   _zz_11359;
  wire       [15:0]   _zz_11360;
  wire       [15:0]   _zz_11361;
  wire       [15:0]   _zz_11362;
  wire       [15:0]   _zz_11363;
  wire       [15:0]   _zz_11364;
  wire       [15:0]   _zz_11365;
  wire       [15:0]   _zz_11366;
  wire       [15:0]   _zz_11367;
  wire       [15:0]   _zz_11368;
  wire       [15:0]   _zz_11369;
  wire       [15:0]   _zz_11370;
  wire       [15:0]   _zz_11371;
  wire       [15:0]   _zz_11372;
  wire       [15:0]   _zz_11373;
  wire       [15:0]   _zz_11374;
  wire       [15:0]   _zz_11375;
  wire       [15:0]   _zz_11376;
  wire       [15:0]   _zz_11377;
  wire       [15:0]   _zz_11378;
  wire       [15:0]   _zz_11379;
  wire       [15:0]   _zz_11380;
  wire       [15:0]   _zz_11381;
  wire       [15:0]   _zz_11382;
  wire       [15:0]   _zz_11383;
  wire       [15:0]   _zz_11384;
  wire       [15:0]   _zz_11385;
  wire       [15:0]   _zz_11386;
  wire       [15:0]   _zz_11387;
  wire       [15:0]   _zz_11388;
  wire       [15:0]   _zz_11389;
  wire       [15:0]   _zz_11390;
  wire       [15:0]   _zz_11391;
  wire       [15:0]   _zz_11392;
  wire       [15:0]   _zz_11393;
  wire       [15:0]   _zz_11394;
  wire       [15:0]   _zz_11395;
  wire       [15:0]   _zz_11396;
  wire       [15:0]   _zz_11397;
  wire       [15:0]   _zz_11398;
  wire       [15:0]   _zz_11399;
  wire       [15:0]   _zz_11400;
  wire       [15:0]   _zz_11401;
  wire       [15:0]   _zz_11402;
  wire       [15:0]   _zz_11403;
  wire       [15:0]   _zz_11404;
  wire       [15:0]   _zz_11405;
  wire       [15:0]   _zz_11406;
  wire       [15:0]   _zz_11407;
  wire       [15:0]   _zz_11408;
  wire       [15:0]   _zz_11409;
  wire       [15:0]   _zz_11410;
  wire       [15:0]   _zz_11411;
  wire       [15:0]   _zz_11412;
  wire       [15:0]   _zz_11413;
  wire       [15:0]   _zz_11414;
  wire       [15:0]   _zz_11415;
  wire       [15:0]   _zz_11416;
  wire       [15:0]   _zz_11417;
  wire       [15:0]   _zz_11418;
  wire       [15:0]   _zz_11419;
  wire       [15:0]   _zz_11420;
  wire       [15:0]   _zz_11421;
  wire       [15:0]   _zz_11422;
  wire       [15:0]   _zz_11423;
  wire       [15:0]   _zz_11424;
  wire       [15:0]   _zz_11425;
  wire       [15:0]   _zz_11426;
  wire       [15:0]   _zz_11427;
  wire       [15:0]   _zz_11428;
  wire       [15:0]   _zz_11429;
  wire       [15:0]   _zz_11430;
  wire       [15:0]   _zz_11431;
  wire       [15:0]   _zz_11432;
  wire       [15:0]   _zz_11433;
  wire       [15:0]   _zz_11434;
  wire       [15:0]   _zz_11435;
  wire       [15:0]   _zz_11436;
  wire       [15:0]   _zz_11437;
  wire       [15:0]   _zz_11438;
  wire       [15:0]   _zz_11439;
  wire       [15:0]   _zz_11440;
  wire       [15:0]   _zz_11441;
  wire       [15:0]   _zz_11442;
  wire       [15:0]   _zz_11443;
  wire       [15:0]   _zz_11444;
  wire       [15:0]   _zz_11445;
  wire       [15:0]   _zz_11446;
  wire       [15:0]   _zz_11447;
  wire       [15:0]   _zz_11448;
  wire       [15:0]   _zz_11449;
  wire       [15:0]   _zz_11450;
  wire       [15:0]   _zz_11451;
  wire       [15:0]   _zz_11452;
  wire       [15:0]   _zz_11453;
  wire       [15:0]   _zz_11454;
  wire       [15:0]   _zz_11455;
  wire       [15:0]   _zz_11456;
  wire       [15:0]   _zz_11457;
  wire       [15:0]   _zz_11458;
  wire       [15:0]   _zz_11459;
  wire       [15:0]   _zz_11460;
  wire       [15:0]   _zz_11461;
  wire       [15:0]   _zz_11462;
  wire       [15:0]   _zz_11463;
  wire       [15:0]   _zz_11464;
  wire       [15:0]   _zz_11465;
  wire       [15:0]   _zz_11466;
  wire       [15:0]   _zz_11467;
  wire       [15:0]   _zz_11468;
  wire       [15:0]   _zz_11469;
  wire       [15:0]   _zz_11470;
  wire       [15:0]   _zz_11471;
  wire       [15:0]   _zz_11472;
  wire       [15:0]   _zz_11473;
  wire       [15:0]   _zz_11474;
  wire       [15:0]   _zz_11475;
  wire       [15:0]   _zz_11476;
  wire       [15:0]   _zz_11477;
  wire       [15:0]   _zz_11478;
  wire       [15:0]   _zz_11479;
  wire       [15:0]   _zz_11480;
  wire       [15:0]   _zz_11481;
  wire       [15:0]   _zz_11482;
  wire       [15:0]   _zz_11483;
  wire       [15:0]   _zz_11484;
  wire       [15:0]   _zz_11485;
  wire       [15:0]   _zz_11486;
  wire       [15:0]   _zz_11487;
  wire       [15:0]   _zz_11488;
  wire       [15:0]   _zz_11489;
  wire       [15:0]   _zz_11490;
  wire       [15:0]   _zz_11491;
  wire       [15:0]   _zz_11492;
  wire       [15:0]   _zz_11493;
  wire       [15:0]   _zz_11494;
  wire       [15:0]   _zz_11495;
  wire       [15:0]   _zz_11496;
  wire       [15:0]   _zz_11497;
  wire       [15:0]   _zz_11498;
  wire       [15:0]   _zz_11499;
  wire       [15:0]   _zz_11500;
  wire       [15:0]   _zz_11501;
  wire       [15:0]   _zz_11502;
  wire       [15:0]   _zz_11503;
  wire       [15:0]   _zz_11504;
  wire       [15:0]   _zz_11505;
  wire       [15:0]   _zz_11506;
  wire       [15:0]   _zz_11507;
  wire       [15:0]   _zz_11508;
  wire       [15:0]   _zz_11509;
  wire       [15:0]   _zz_11510;
  wire       [15:0]   _zz_11511;
  wire       [15:0]   _zz_11512;
  wire       [15:0]   _zz_11513;
  wire       [15:0]   _zz_11514;
  wire       [15:0]   _zz_11515;
  wire       [15:0]   _zz_11516;
  wire       [15:0]   _zz_11517;
  wire       [15:0]   _zz_11518;
  wire       [15:0]   _zz_11519;
  wire       [15:0]   _zz_11520;
  wire       [15:0]   _zz_11521;
  wire       [15:0]   _zz_11522;
  wire       [15:0]   _zz_11523;
  wire       [15:0]   _zz_11524;
  wire       [15:0]   _zz_11525;
  wire       [15:0]   _zz_11526;
  wire       [15:0]   _zz_11527;
  wire       [15:0]   _zz_11528;
  wire       [15:0]   _zz_11529;
  wire       [15:0]   _zz_11530;
  wire       [15:0]   _zz_11531;
  wire       [15:0]   _zz_11532;
  wire       [15:0]   _zz_11533;
  wire       [15:0]   _zz_11534;
  wire       [15:0]   _zz_11535;
  wire       [15:0]   _zz_11536;
  wire       [15:0]   _zz_11537;
  wire       [15:0]   _zz_11538;
  wire       [15:0]   _zz_11539;
  wire       [15:0]   _zz_11540;
  wire       [15:0]   _zz_11541;
  wire       [15:0]   _zz_11542;
  wire       [15:0]   _zz_11543;
  wire       [15:0]   _zz_11544;
  wire       [15:0]   _zz_11545;
  wire       [15:0]   _zz_11546;
  wire       [15:0]   _zz_11547;
  wire       [15:0]   _zz_11548;
  wire       [15:0]   _zz_11549;
  wire       [15:0]   _zz_11550;
  wire       [15:0]   _zz_11551;
  wire       [15:0]   _zz_11552;
  wire       [15:0]   _zz_11553;
  wire       [15:0]   _zz_11554;
  wire       [15:0]   _zz_11555;
  wire       [15:0]   _zz_11556;
  wire       [15:0]   _zz_11557;
  wire       [15:0]   _zz_11558;
  wire       [15:0]   _zz_11559;
  wire       [15:0]   _zz_11560;
  wire       [15:0]   _zz_11561;
  wire       [15:0]   _zz_11562;
  wire       [15:0]   _zz_11563;
  wire       [15:0]   _zz_11564;
  wire       [15:0]   _zz_11565;
  wire       [15:0]   _zz_11566;
  wire       [15:0]   _zz_11567;
  wire       [15:0]   _zz_11568;
  wire       [15:0]   _zz_11569;
  wire       [15:0]   _zz_11570;
  wire       [15:0]   _zz_11571;
  wire       [15:0]   _zz_11572;
  wire       [15:0]   _zz_11573;
  wire       [15:0]   _zz_11574;
  wire       [15:0]   _zz_11575;
  wire       [15:0]   _zz_11576;
  wire       [15:0]   _zz_11577;
  wire       [15:0]   _zz_11578;
  wire       [15:0]   _zz_11579;
  wire       [15:0]   _zz_11580;
  wire       [15:0]   _zz_11581;
  wire       [15:0]   _zz_11582;
  wire       [15:0]   _zz_11583;
  wire       [15:0]   _zz_11584;
  wire       [15:0]   _zz_11585;
  wire       [15:0]   _zz_11586;
  wire       [15:0]   _zz_11587;
  wire       [15:0]   _zz_11588;
  wire       [15:0]   _zz_11589;
  wire       [15:0]   _zz_11590;
  wire       [15:0]   _zz_11591;
  wire       [15:0]   _zz_11592;
  wire       [15:0]   _zz_11593;
  wire       [15:0]   _zz_11594;
  wire       [15:0]   _zz_11595;
  wire       [15:0]   _zz_11596;
  wire       [15:0]   _zz_11597;
  wire       [15:0]   _zz_11598;
  wire       [15:0]   _zz_11599;
  wire       [15:0]   _zz_11600;
  wire       [15:0]   _zz_11601;
  wire       [15:0]   _zz_11602;
  wire       [15:0]   _zz_11603;
  wire       [15:0]   _zz_11604;
  wire       [15:0]   _zz_11605;
  wire       [15:0]   _zz_11606;
  wire       [15:0]   _zz_11607;
  wire       [15:0]   _zz_11608;
  wire       [15:0]   _zz_11609;
  wire       [15:0]   _zz_11610;
  wire       [15:0]   _zz_11611;
  wire       [15:0]   _zz_11612;
  wire       [15:0]   _zz_11613;
  wire       [15:0]   _zz_11614;
  wire       [15:0]   _zz_11615;
  wire       [15:0]   _zz_11616;
  wire       [15:0]   _zz_11617;
  wire       [15:0]   _zz_11618;
  wire       [15:0]   _zz_11619;
  wire       [15:0]   _zz_11620;
  wire       [15:0]   _zz_11621;
  wire       [15:0]   _zz_11622;
  wire       [15:0]   _zz_11623;
  wire       [15:0]   _zz_11624;
  wire       [15:0]   _zz_11625;
  wire       [15:0]   _zz_11626;
  wire       [15:0]   _zz_11627;
  wire       [15:0]   _zz_11628;
  wire       [15:0]   _zz_11629;
  wire       [15:0]   _zz_11630;
  wire       [15:0]   _zz_11631;
  wire       [15:0]   _zz_11632;
  wire       [15:0]   _zz_11633;
  wire       [15:0]   _zz_11634;
  wire       [15:0]   _zz_11635;
  wire       [15:0]   _zz_11636;
  wire       [15:0]   _zz_11637;
  wire       [15:0]   _zz_11638;
  wire       [15:0]   _zz_11639;
  wire       [15:0]   _zz_11640;
  wire       [15:0]   _zz_11641;
  wire       [15:0]   _zz_11642;
  wire       [15:0]   _zz_11643;
  wire       [15:0]   _zz_11644;
  wire       [15:0]   _zz_11645;
  wire       [15:0]   _zz_11646;
  wire       [15:0]   _zz_11647;
  wire       [15:0]   _zz_11648;
  wire       [15:0]   _zz_11649;
  wire       [15:0]   _zz_11650;
  wire       [15:0]   _zz_11651;
  wire       [15:0]   _zz_11652;
  wire       [15:0]   _zz_11653;
  wire       [15:0]   _zz_11654;
  wire       [15:0]   _zz_11655;
  wire       [15:0]   _zz_11656;
  wire       [15:0]   _zz_11657;
  wire       [15:0]   _zz_11658;
  wire       [15:0]   _zz_11659;
  wire       [15:0]   _zz_11660;
  wire       [15:0]   _zz_11661;
  wire       [15:0]   _zz_11662;
  wire       [15:0]   _zz_11663;
  wire       [15:0]   _zz_11664;
  wire       [15:0]   _zz_11665;
  wire       [15:0]   _zz_11666;
  wire       [15:0]   _zz_11667;
  wire       [15:0]   _zz_11668;
  wire       [15:0]   _zz_11669;
  wire       [15:0]   _zz_11670;
  wire       [15:0]   _zz_11671;
  wire       [15:0]   _zz_11672;
  wire       [15:0]   _zz_11673;
  wire       [15:0]   _zz_11674;
  wire       [15:0]   _zz_11675;
  wire       [15:0]   _zz_11676;
  wire       [15:0]   _zz_11677;
  wire       [15:0]   _zz_11678;
  wire       [15:0]   _zz_11679;
  wire       [15:0]   _zz_11680;
  wire       [15:0]   _zz_11681;
  wire       [15:0]   _zz_11682;
  wire       [15:0]   _zz_11683;
  wire       [15:0]   _zz_11684;
  wire       [15:0]   _zz_11685;
  wire       [15:0]   _zz_11686;
  wire       [15:0]   _zz_11687;
  wire       [15:0]   _zz_11688;
  wire       [15:0]   _zz_11689;
  wire       [15:0]   _zz_11690;
  wire       [15:0]   _zz_11691;
  wire       [15:0]   _zz_11692;
  wire       [15:0]   _zz_11693;
  wire       [15:0]   _zz_11694;
  wire       [15:0]   _zz_11695;
  wire       [15:0]   _zz_11696;
  wire       [15:0]   _zz_11697;
  wire       [15:0]   _zz_11698;
  wire       [15:0]   _zz_11699;
  wire       [15:0]   _zz_11700;
  wire       [15:0]   _zz_11701;
  wire       [15:0]   _zz_11702;
  wire       [15:0]   _zz_11703;
  wire       [15:0]   _zz_11704;
  wire       [15:0]   _zz_11705;
  wire       [15:0]   _zz_11706;
  wire       [15:0]   _zz_11707;
  wire       [15:0]   _zz_11708;
  wire       [15:0]   _zz_11709;
  wire       [15:0]   _zz_11710;
  wire       [15:0]   _zz_11711;
  wire       [15:0]   _zz_11712;
  wire       [15:0]   _zz_11713;
  wire       [15:0]   _zz_11714;
  wire       [15:0]   _zz_11715;
  wire       [15:0]   _zz_11716;
  wire       [15:0]   _zz_11717;
  wire       [15:0]   _zz_11718;
  wire       [15:0]   _zz_11719;
  wire       [15:0]   _zz_11720;
  wire       [15:0]   _zz_11721;
  wire       [15:0]   _zz_11722;
  wire       [15:0]   _zz_11723;
  wire       [15:0]   _zz_11724;
  wire       [15:0]   _zz_11725;
  wire       [15:0]   _zz_11726;
  wire       [15:0]   _zz_11727;
  wire       [15:0]   _zz_11728;
  wire       [15:0]   _zz_11729;
  wire       [15:0]   _zz_11730;
  wire       [15:0]   _zz_11731;
  wire       [15:0]   _zz_11732;
  wire       [15:0]   _zz_11733;
  wire       [15:0]   _zz_11734;
  wire       [15:0]   _zz_11735;
  wire       [15:0]   _zz_11736;
  wire       [15:0]   _zz_11737;
  wire       [15:0]   _zz_11738;
  wire       [15:0]   _zz_11739;
  wire       [15:0]   _zz_11740;
  wire       [15:0]   _zz_11741;
  wire       [15:0]   _zz_11742;
  wire       [15:0]   _zz_11743;
  wire       [15:0]   _zz_11744;
  wire       [15:0]   _zz_11745;
  wire       [15:0]   _zz_11746;
  wire       [15:0]   _zz_11747;
  wire       [15:0]   _zz_11748;
  wire       [15:0]   _zz_11749;
  wire       [15:0]   _zz_11750;
  wire       [15:0]   _zz_11751;
  wire       [15:0]   _zz_11752;
  wire       [15:0]   _zz_11753;
  wire       [15:0]   _zz_11754;
  wire       [15:0]   _zz_11755;
  wire       [15:0]   _zz_11756;
  wire       [15:0]   _zz_11757;
  wire       [15:0]   _zz_11758;
  wire       [15:0]   _zz_11759;
  wire       [15:0]   _zz_11760;
  wire       [15:0]   _zz_11761;
  wire       [15:0]   _zz_11762;
  wire       [15:0]   _zz_11763;
  wire       [15:0]   _zz_11764;
  wire       [15:0]   _zz_11765;
  wire       [15:0]   _zz_11766;
  wire       [15:0]   _zz_11767;
  wire       [15:0]   _zz_11768;
  wire       [15:0]   _zz_11769;
  wire       [15:0]   _zz_11770;
  wire       [15:0]   _zz_11771;
  wire       [15:0]   _zz_11772;
  wire       [15:0]   _zz_11773;
  wire       [15:0]   _zz_11774;
  wire       [15:0]   _zz_11775;
  wire       [15:0]   _zz_11776;
  wire       [15:0]   _zz_11777;
  wire       [15:0]   _zz_11778;
  wire       [15:0]   _zz_11779;
  wire       [15:0]   _zz_11780;
  wire       [15:0]   _zz_11781;
  wire       [15:0]   _zz_11782;
  wire       [15:0]   _zz_11783;
  wire       [15:0]   _zz_11784;
  wire       [15:0]   _zz_11785;
  wire       [15:0]   _zz_11786;
  wire       [15:0]   _zz_11787;
  wire       [15:0]   _zz_11788;
  wire       [15:0]   _zz_11789;
  wire       [15:0]   _zz_11790;
  wire       [15:0]   _zz_11791;
  wire       [15:0]   _zz_11792;
  wire       [15:0]   _zz_11793;
  wire       [15:0]   _zz_11794;
  wire       [15:0]   _zz_11795;
  wire       [15:0]   _zz_11796;
  wire       [15:0]   _zz_11797;
  wire       [15:0]   _zz_11798;
  wire       [15:0]   _zz_11799;
  wire       [15:0]   _zz_11800;
  wire       [15:0]   _zz_11801;
  wire       [15:0]   _zz_11802;
  wire       [15:0]   _zz_11803;
  wire       [15:0]   _zz_11804;
  wire       [15:0]   _zz_11805;
  wire       [15:0]   _zz_11806;
  wire       [15:0]   _zz_11807;
  wire       [15:0]   _zz_11808;
  wire       [15:0]   _zz_11809;
  wire       [15:0]   _zz_11810;
  wire       [15:0]   _zz_11811;
  wire       [15:0]   _zz_11812;
  wire       [15:0]   _zz_11813;
  wire       [15:0]   _zz_11814;
  wire       [15:0]   _zz_11815;
  wire       [15:0]   _zz_11816;
  wire       [15:0]   _zz_11817;
  wire       [15:0]   _zz_11818;
  wire       [15:0]   _zz_11819;
  wire       [15:0]   _zz_11820;
  wire       [15:0]   _zz_11821;
  wire       [15:0]   _zz_11822;
  wire       [15:0]   _zz_11823;
  wire       [15:0]   _zz_11824;
  wire       [15:0]   _zz_11825;
  wire       [15:0]   _zz_11826;
  wire       [15:0]   _zz_11827;
  wire       [15:0]   _zz_11828;
  wire       [15:0]   _zz_11829;
  wire       [15:0]   _zz_11830;
  wire       [15:0]   _zz_11831;
  wire       [15:0]   _zz_11832;
  wire       [15:0]   _zz_11833;
  wire       [15:0]   _zz_11834;
  wire       [15:0]   _zz_11835;
  wire       [15:0]   _zz_11836;
  wire       [15:0]   _zz_11837;
  wire       [15:0]   _zz_11838;
  wire       [15:0]   _zz_11839;
  wire       [15:0]   _zz_11840;
  wire       [15:0]   _zz_11841;
  wire       [15:0]   _zz_11842;
  wire       [15:0]   _zz_11843;
  wire       [15:0]   _zz_11844;
  wire       [15:0]   _zz_11845;
  wire       [15:0]   _zz_11846;
  wire       [15:0]   _zz_11847;
  wire       [15:0]   _zz_11848;
  wire       [15:0]   _zz_11849;
  wire       [15:0]   _zz_11850;
  wire       [15:0]   _zz_11851;
  wire       [15:0]   _zz_11852;
  wire       [15:0]   _zz_11853;
  wire       [15:0]   _zz_11854;
  wire       [15:0]   _zz_11855;
  wire       [15:0]   _zz_11856;
  wire       [15:0]   _zz_11857;
  wire       [15:0]   _zz_11858;
  wire       [15:0]   _zz_11859;
  wire       [15:0]   _zz_11860;
  wire       [15:0]   _zz_11861;
  wire       [15:0]   _zz_11862;
  wire       [15:0]   _zz_11863;
  wire       [15:0]   _zz_11864;
  wire       [15:0]   _zz_11865;
  wire       [15:0]   _zz_11866;
  wire       [15:0]   _zz_11867;
  wire       [15:0]   _zz_11868;
  wire       [15:0]   _zz_11869;
  wire       [15:0]   _zz_11870;
  wire       [15:0]   _zz_11871;
  wire       [15:0]   _zz_11872;
  wire       [15:0]   _zz_11873;
  wire       [15:0]   _zz_11874;
  wire       [15:0]   _zz_11875;
  wire       [15:0]   _zz_11876;
  wire       [15:0]   _zz_11877;
  wire       [15:0]   _zz_11878;
  wire       [15:0]   _zz_11879;
  wire       [15:0]   _zz_11880;
  wire       [15:0]   _zz_11881;
  wire       [15:0]   _zz_11882;
  wire       [15:0]   _zz_11883;
  wire       [15:0]   _zz_11884;
  wire       [15:0]   _zz_11885;
  wire       [15:0]   _zz_11886;
  wire       [15:0]   _zz_11887;
  wire       [15:0]   _zz_11888;
  wire       [15:0]   _zz_11889;
  wire       [15:0]   _zz_11890;
  wire       [15:0]   _zz_11891;
  wire       [15:0]   _zz_11892;
  wire       [15:0]   _zz_11893;
  wire       [15:0]   _zz_11894;
  wire       [15:0]   _zz_11895;
  wire       [15:0]   _zz_11896;
  wire       [15:0]   _zz_11897;
  wire       [15:0]   _zz_11898;
  wire       [15:0]   _zz_11899;
  wire       [15:0]   _zz_11900;
  wire       [15:0]   _zz_11901;
  wire       [15:0]   _zz_11902;
  wire       [15:0]   _zz_11903;
  wire       [15:0]   _zz_11904;
  wire       [15:0]   _zz_11905;
  wire       [15:0]   _zz_11906;
  wire       [15:0]   _zz_11907;
  wire       [15:0]   _zz_11908;
  wire       [15:0]   _zz_11909;
  wire       [15:0]   _zz_11910;
  wire       [15:0]   _zz_11911;
  wire       [15:0]   _zz_11912;
  wire       [15:0]   _zz_11913;
  wire       [15:0]   _zz_11914;
  wire       [15:0]   _zz_11915;
  wire       [15:0]   _zz_11916;
  wire       [15:0]   _zz_11917;
  wire       [15:0]   _zz_11918;
  wire       [15:0]   _zz_11919;
  wire       [15:0]   _zz_11920;
  wire       [15:0]   _zz_11921;
  wire       [15:0]   _zz_11922;
  wire       [15:0]   _zz_11923;
  wire       [15:0]   _zz_11924;
  wire       [15:0]   _zz_11925;
  wire       [15:0]   _zz_11926;
  wire       [15:0]   _zz_11927;
  wire       [15:0]   _zz_11928;
  wire       [15:0]   _zz_11929;
  wire       [15:0]   _zz_11930;
  wire       [15:0]   _zz_11931;
  wire       [15:0]   _zz_11932;
  wire       [15:0]   _zz_11933;
  wire       [15:0]   _zz_11934;
  wire       [15:0]   _zz_11935;
  wire       [15:0]   _zz_11936;
  wire       [15:0]   _zz_11937;
  wire       [15:0]   _zz_11938;
  wire       [15:0]   _zz_11939;
  wire       [15:0]   _zz_11940;
  wire       [15:0]   _zz_11941;
  wire       [15:0]   _zz_11942;
  wire       [15:0]   _zz_11943;
  wire       [15:0]   _zz_11944;
  wire       [15:0]   _zz_11945;
  wire       [15:0]   _zz_11946;
  wire       [15:0]   _zz_11947;
  wire       [15:0]   _zz_11948;
  wire       [15:0]   _zz_11949;
  wire       [15:0]   _zz_11950;
  wire       [15:0]   _zz_11951;
  wire       [15:0]   _zz_11952;
  wire       [15:0]   _zz_11953;
  wire       [15:0]   _zz_11954;
  wire       [15:0]   _zz_11955;
  wire       [15:0]   _zz_11956;
  wire       [15:0]   _zz_11957;
  wire       [15:0]   _zz_11958;
  wire       [15:0]   _zz_11959;
  wire       [15:0]   _zz_11960;
  wire       [15:0]   _zz_11961;
  wire       [15:0]   _zz_11962;
  wire       [15:0]   _zz_11963;
  wire       [15:0]   _zz_11964;
  wire       [15:0]   _zz_11965;
  wire       [15:0]   _zz_11966;
  wire       [15:0]   _zz_11967;
  wire       [15:0]   _zz_11968;
  wire       [15:0]   _zz_11969;
  wire       [15:0]   _zz_11970;
  wire       [15:0]   _zz_11971;
  wire       [15:0]   _zz_11972;
  wire       [15:0]   _zz_11973;
  wire       [15:0]   _zz_11974;
  wire       [15:0]   _zz_11975;
  wire       [15:0]   _zz_11976;
  wire       [15:0]   _zz_11977;
  wire       [15:0]   _zz_11978;
  wire       [15:0]   _zz_11979;
  wire       [15:0]   _zz_11980;
  wire       [15:0]   _zz_11981;
  wire       [15:0]   _zz_11982;
  wire       [15:0]   _zz_11983;
  wire       [15:0]   _zz_11984;
  wire       [15:0]   _zz_11985;
  wire       [15:0]   _zz_11986;
  wire       [15:0]   _zz_11987;
  wire       [15:0]   _zz_11988;
  wire       [15:0]   _zz_11989;
  wire       [15:0]   _zz_11990;
  wire       [15:0]   _zz_11991;
  wire       [15:0]   _zz_11992;
  wire       [15:0]   _zz_11993;
  wire       [15:0]   _zz_11994;
  wire       [15:0]   _zz_11995;
  wire       [15:0]   _zz_11996;
  wire       [15:0]   _zz_11997;
  wire       [15:0]   _zz_11998;
  wire       [15:0]   _zz_11999;
  wire       [15:0]   _zz_12000;
  wire       [15:0]   _zz_12001;
  wire       [15:0]   _zz_12002;
  wire       [15:0]   _zz_12003;
  wire       [15:0]   _zz_12004;
  wire       [15:0]   _zz_12005;
  wire       [15:0]   _zz_12006;
  wire       [15:0]   _zz_12007;
  wire       [15:0]   _zz_12008;
  wire       [15:0]   _zz_12009;
  wire       [15:0]   _zz_12010;
  wire       [15:0]   _zz_12011;
  wire       [15:0]   _zz_12012;
  wire       [15:0]   _zz_12013;
  wire       [15:0]   _zz_12014;
  wire       [15:0]   _zz_12015;
  wire       [15:0]   _zz_12016;
  wire       [15:0]   _zz_12017;
  wire       [15:0]   _zz_12018;
  wire       [15:0]   _zz_12019;
  wire       [15:0]   _zz_12020;
  wire       [15:0]   _zz_12021;
  wire       [15:0]   _zz_12022;
  wire       [15:0]   _zz_12023;
  wire       [15:0]   _zz_12024;
  wire       [15:0]   _zz_12025;
  wire       [15:0]   _zz_12026;
  wire       [15:0]   _zz_12027;
  wire       [15:0]   _zz_12028;
  wire       [15:0]   _zz_12029;
  wire       [15:0]   _zz_12030;
  wire       [15:0]   _zz_12031;
  wire       [15:0]   _zz_12032;
  wire       [15:0]   _zz_12033;
  wire       [15:0]   _zz_12034;
  wire       [15:0]   _zz_12035;
  wire       [15:0]   _zz_12036;
  wire       [15:0]   _zz_12037;
  wire       [15:0]   _zz_12038;
  wire       [15:0]   _zz_12039;
  wire       [15:0]   _zz_12040;
  wire       [15:0]   _zz_12041;
  wire       [15:0]   _zz_12042;
  wire       [15:0]   _zz_12043;
  wire       [15:0]   _zz_12044;
  wire       [15:0]   _zz_12045;
  wire       [15:0]   _zz_12046;
  wire       [15:0]   _zz_12047;
  wire       [15:0]   _zz_12048;
  wire       [15:0]   _zz_12049;
  wire       [15:0]   _zz_12050;
  wire       [15:0]   _zz_12051;
  wire       [15:0]   _zz_12052;
  wire       [15:0]   _zz_12053;
  wire       [15:0]   _zz_12054;
  wire       [15:0]   _zz_12055;
  wire       [15:0]   _zz_12056;
  wire       [15:0]   _zz_12057;
  wire       [15:0]   _zz_12058;
  wire       [15:0]   _zz_12059;
  wire       [15:0]   _zz_12060;
  wire       [15:0]   _zz_12061;
  wire       [15:0]   _zz_12062;
  wire       [15:0]   _zz_12063;
  wire       [15:0]   _zz_12064;
  wire       [15:0]   _zz_12065;
  wire       [15:0]   _zz_12066;
  wire       [15:0]   _zz_12067;
  wire       [15:0]   _zz_12068;
  wire       [15:0]   _zz_12069;
  wire       [15:0]   _zz_12070;
  wire       [15:0]   _zz_12071;
  wire       [15:0]   _zz_12072;
  wire       [15:0]   _zz_12073;
  wire       [15:0]   _zz_12074;
  wire       [15:0]   _zz_12075;
  wire       [15:0]   _zz_12076;
  wire       [15:0]   _zz_12077;
  wire       [15:0]   _zz_12078;
  wire       [15:0]   _zz_12079;
  wire       [15:0]   _zz_12080;
  wire       [15:0]   _zz_12081;
  wire       [15:0]   _zz_12082;
  wire       [15:0]   _zz_12083;
  wire       [15:0]   _zz_12084;
  wire       [15:0]   _zz_12085;
  wire       [15:0]   _zz_12086;
  wire       [15:0]   _zz_12087;
  wire       [15:0]   _zz_12088;
  wire       [15:0]   _zz_12089;
  wire       [15:0]   _zz_12090;
  wire       [15:0]   _zz_12091;
  wire       [15:0]   _zz_12092;
  wire       [15:0]   _zz_12093;
  wire       [15:0]   _zz_12094;
  wire       [15:0]   _zz_12095;
  wire       [15:0]   _zz_12096;
  wire       [15:0]   _zz_12097;
  wire       [15:0]   _zz_12098;
  wire       [15:0]   _zz_12099;
  wire       [15:0]   _zz_12100;
  wire       [15:0]   _zz_12101;
  wire       [15:0]   _zz_12102;
  wire       [15:0]   _zz_12103;
  wire       [15:0]   _zz_12104;
  wire       [15:0]   _zz_12105;
  wire       [15:0]   _zz_12106;
  wire       [15:0]   _zz_12107;
  wire       [15:0]   _zz_12108;
  wire       [15:0]   _zz_12109;
  wire       [15:0]   _zz_12110;
  wire       [15:0]   _zz_12111;
  wire       [15:0]   _zz_12112;
  wire       [15:0]   _zz_12113;
  wire       [15:0]   _zz_12114;
  wire       [15:0]   _zz_12115;
  wire       [15:0]   _zz_12116;
  wire       [15:0]   _zz_12117;
  wire       [15:0]   _zz_12118;
  wire       [15:0]   _zz_12119;
  wire       [15:0]   _zz_12120;
  wire       [15:0]   _zz_12121;
  wire       [15:0]   _zz_12122;
  wire       [15:0]   _zz_12123;
  wire       [15:0]   _zz_12124;
  wire       [15:0]   _zz_12125;
  wire       [15:0]   _zz_12126;
  wire       [15:0]   _zz_12127;
  wire       [15:0]   _zz_12128;
  wire       [15:0]   _zz_12129;
  wire       [15:0]   _zz_12130;
  wire       [15:0]   _zz_12131;
  wire       [15:0]   _zz_12132;
  wire       [15:0]   _zz_12133;
  wire       [15:0]   _zz_12134;
  wire       [15:0]   _zz_12135;
  wire       [15:0]   _zz_12136;
  wire       [15:0]   _zz_12137;
  wire       [15:0]   _zz_12138;
  wire       [15:0]   _zz_12139;
  wire       [15:0]   _zz_12140;
  wire       [15:0]   _zz_12141;
  wire       [15:0]   _zz_12142;
  wire       [15:0]   _zz_12143;
  wire       [15:0]   _zz_12144;
  wire       [15:0]   _zz_12145;
  wire       [15:0]   _zz_12146;
  wire       [15:0]   _zz_12147;
  wire       [15:0]   _zz_12148;
  wire       [15:0]   _zz_12149;
  wire       [15:0]   _zz_12150;
  wire       [15:0]   _zz_12151;
  wire       [15:0]   _zz_12152;
  wire       [15:0]   _zz_12153;
  wire       [15:0]   _zz_12154;
  wire       [15:0]   _zz_12155;
  wire       [15:0]   _zz_12156;
  wire       [15:0]   _zz_12157;
  wire       [15:0]   _zz_12158;
  wire       [15:0]   _zz_12159;
  wire       [15:0]   _zz_12160;
  wire       [15:0]   _zz_12161;
  wire       [15:0]   _zz_12162;
  wire       [15:0]   _zz_12163;
  wire       [15:0]   _zz_12164;
  wire       [15:0]   _zz_12165;
  wire       [15:0]   _zz_12166;
  wire       [15:0]   _zz_12167;
  wire       [15:0]   _zz_12168;
  wire       [15:0]   _zz_12169;
  wire       [15:0]   _zz_12170;
  wire       [15:0]   _zz_12171;
  wire       [15:0]   _zz_12172;
  wire       [15:0]   _zz_12173;
  wire       [15:0]   _zz_12174;
  wire       [15:0]   _zz_12175;
  wire       [15:0]   _zz_12176;
  wire       [15:0]   _zz_12177;
  wire       [15:0]   _zz_12178;
  wire       [15:0]   _zz_12179;
  wire       [15:0]   _zz_12180;
  wire       [15:0]   _zz_12181;
  wire       [15:0]   _zz_12182;
  wire       [15:0]   _zz_12183;
  wire       [15:0]   _zz_12184;
  wire       [15:0]   _zz_12185;
  wire       [15:0]   _zz_12186;
  wire       [15:0]   _zz_12187;
  wire       [15:0]   _zz_12188;
  wire       [15:0]   _zz_12189;
  wire       [15:0]   _zz_12190;
  wire       [15:0]   _zz_12191;
  wire       [15:0]   _zz_12192;
  wire       [15:0]   _zz_12193;
  wire       [15:0]   _zz_12194;
  wire       [15:0]   _zz_12195;
  wire       [15:0]   _zz_12196;
  wire       [15:0]   _zz_12197;
  wire       [15:0]   _zz_12198;
  wire       [15:0]   _zz_12199;
  wire       [15:0]   _zz_12200;
  wire       [15:0]   _zz_12201;
  wire       [15:0]   _zz_12202;
  wire       [15:0]   _zz_12203;
  wire       [15:0]   _zz_12204;
  wire       [15:0]   _zz_12205;
  wire       [15:0]   _zz_12206;
  wire       [15:0]   _zz_12207;
  wire       [15:0]   _zz_12208;
  wire       [15:0]   _zz_12209;
  wire       [15:0]   _zz_12210;
  wire       [15:0]   _zz_12211;
  wire       [15:0]   _zz_12212;
  wire       [15:0]   _zz_12213;
  wire       [15:0]   _zz_12214;
  wire       [15:0]   _zz_12215;
  wire       [15:0]   _zz_12216;
  wire       [15:0]   _zz_12217;
  wire       [15:0]   _zz_12218;
  wire       [15:0]   _zz_12219;
  wire       [15:0]   _zz_12220;
  wire       [15:0]   _zz_12221;
  wire       [15:0]   _zz_12222;
  wire       [15:0]   _zz_12223;
  wire       [15:0]   _zz_12224;
  wire       [15:0]   _zz_12225;
  wire       [15:0]   _zz_12226;
  wire       [15:0]   _zz_12227;
  wire       [15:0]   _zz_12228;
  wire       [15:0]   _zz_12229;
  wire       [15:0]   _zz_12230;
  wire       [15:0]   _zz_12231;
  wire       [15:0]   _zz_12232;
  wire       [15:0]   _zz_12233;
  wire       [15:0]   _zz_12234;
  wire       [15:0]   _zz_12235;
  wire       [15:0]   _zz_12236;
  wire       [15:0]   _zz_12237;
  wire       [15:0]   _zz_12238;
  wire       [15:0]   _zz_12239;
  wire       [15:0]   _zz_12240;
  wire       [15:0]   _zz_12241;
  wire       [15:0]   _zz_12242;
  wire       [15:0]   _zz_12243;
  wire       [15:0]   _zz_12244;
  wire       [15:0]   _zz_12245;
  wire       [15:0]   _zz_12246;
  wire       [15:0]   _zz_12247;
  wire       [15:0]   _zz_12248;
  wire       [15:0]   _zz_12249;
  wire       [15:0]   _zz_12250;
  wire       [15:0]   _zz_12251;
  wire       [15:0]   _zz_12252;
  wire       [15:0]   _zz_12253;
  wire       [15:0]   _zz_12254;
  wire       [15:0]   _zz_12255;
  wire       [15:0]   _zz_12256;
  wire       [15:0]   _zz_12257;
  wire       [15:0]   _zz_12258;
  wire       [15:0]   _zz_12259;
  wire       [15:0]   _zz_12260;
  wire       [15:0]   _zz_12261;
  wire       [15:0]   _zz_12262;
  wire       [15:0]   _zz_12263;
  wire       [15:0]   _zz_12264;
  wire       [15:0]   _zz_12265;
  wire       [15:0]   _zz_12266;
  wire       [15:0]   _zz_12267;
  wire       [15:0]   _zz_12268;
  wire       [15:0]   _zz_12269;
  wire       [15:0]   _zz_12270;
  wire       [15:0]   _zz_12271;
  wire       [15:0]   _zz_12272;
  wire       [15:0]   _zz_12273;
  wire       [15:0]   _zz_12274;
  wire       [15:0]   _zz_12275;
  wire       [15:0]   _zz_12276;
  wire       [15:0]   _zz_12277;
  wire       [15:0]   _zz_12278;
  wire       [15:0]   _zz_12279;
  wire       [15:0]   _zz_12280;
  wire       [15:0]   _zz_12281;
  wire       [15:0]   _zz_12282;
  wire       [15:0]   _zz_12283;
  wire       [15:0]   _zz_12284;
  wire       [15:0]   _zz_12285;
  wire       [15:0]   _zz_12286;
  wire       [15:0]   _zz_12287;
  wire       [15:0]   _zz_12288;
  wire       [15:0]   _zz_12289;
  wire       [15:0]   _zz_12290;
  wire       [15:0]   _zz_12291;
  wire       [15:0]   _zz_12292;
  wire       [15:0]   _zz_12293;
  wire       [15:0]   _zz_12294;
  wire       [15:0]   _zz_12295;
  wire       [15:0]   _zz_12296;
  wire       [15:0]   _zz_12297;
  wire       [15:0]   _zz_12298;
  wire       [15:0]   _zz_12299;
  wire       [15:0]   _zz_12300;
  wire       [15:0]   _zz_12301;
  wire       [15:0]   _zz_12302;
  wire       [15:0]   _zz_12303;
  wire       [15:0]   _zz_12304;
  wire       [15:0]   _zz_12305;
  wire       [15:0]   _zz_12306;
  wire       [15:0]   _zz_12307;
  wire       [15:0]   _zz_12308;
  wire       [15:0]   _zz_12309;
  wire       [15:0]   _zz_12310;
  wire       [15:0]   _zz_12311;
  wire       [15:0]   _zz_12312;
  wire       [15:0]   _zz_12313;
  wire       [15:0]   _zz_12314;
  wire       [15:0]   _zz_12315;
  wire       [15:0]   _zz_12316;
  wire       [15:0]   _zz_12317;
  wire       [15:0]   _zz_12318;
  wire       [15:0]   _zz_12319;
  wire       [15:0]   _zz_12320;
  wire       [15:0]   _zz_12321;
  wire       [15:0]   _zz_12322;
  wire       [15:0]   _zz_12323;
  wire       [15:0]   _zz_12324;
  wire       [15:0]   _zz_12325;
  wire       [15:0]   _zz_12326;
  wire       [15:0]   _zz_12327;
  wire       [15:0]   _zz_12328;
  wire       [15:0]   _zz_12329;
  wire       [15:0]   _zz_12330;
  wire       [15:0]   _zz_12331;
  wire       [15:0]   _zz_12332;
  wire       [15:0]   _zz_12333;
  wire       [15:0]   _zz_12334;
  wire       [15:0]   _zz_12335;
  wire       [15:0]   _zz_12336;
  wire       [15:0]   _zz_12337;
  wire       [15:0]   _zz_12338;
  wire       [15:0]   _zz_12339;
  wire       [15:0]   _zz_12340;
  wire       [15:0]   _zz_12341;
  wire       [15:0]   _zz_12342;
  wire       [15:0]   _zz_12343;
  wire       [15:0]   _zz_12344;
  wire       [15:0]   _zz_12345;
  wire       [15:0]   _zz_12346;
  wire       [15:0]   _zz_12347;
  wire       [15:0]   _zz_12348;
  wire       [15:0]   _zz_12349;
  wire       [15:0]   _zz_12350;
  wire       [15:0]   _zz_12351;
  wire       [15:0]   _zz_12352;
  wire       [15:0]   _zz_12353;
  wire       [15:0]   _zz_12354;
  wire       [15:0]   _zz_12355;
  wire       [15:0]   _zz_12356;
  wire       [15:0]   _zz_12357;
  wire       [15:0]   _zz_12358;
  wire       [15:0]   _zz_12359;
  wire       [15:0]   _zz_12360;
  wire       [15:0]   _zz_12361;
  wire       [15:0]   _zz_12362;
  wire       [15:0]   _zz_12363;
  wire       [15:0]   _zz_12364;
  wire       [15:0]   _zz_12365;
  wire       [15:0]   _zz_12366;
  wire       [15:0]   _zz_12367;
  wire       [15:0]   _zz_12368;
  wire       [15:0]   _zz_12369;
  wire       [15:0]   _zz_12370;
  wire       [15:0]   _zz_12371;
  wire       [15:0]   _zz_12372;
  wire       [15:0]   _zz_12373;
  wire       [15:0]   _zz_12374;
  wire       [15:0]   _zz_12375;
  wire       [15:0]   _zz_12376;
  wire       [15:0]   _zz_12377;
  wire       [15:0]   _zz_12378;
  wire       [15:0]   _zz_12379;
  wire       [15:0]   _zz_12380;
  wire       [15:0]   _zz_12381;
  wire       [15:0]   _zz_12382;
  wire       [15:0]   _zz_12383;
  wire       [15:0]   _zz_12384;
  wire       [15:0]   _zz_12385;
  wire       [15:0]   _zz_12386;
  wire       [15:0]   _zz_12387;
  wire       [15:0]   _zz_12388;
  wire       [15:0]   _zz_12389;
  wire       [15:0]   _zz_12390;
  wire       [15:0]   _zz_12391;
  wire       [15:0]   _zz_12392;
  wire       [15:0]   _zz_12393;
  wire       [15:0]   _zz_12394;
  wire       [15:0]   _zz_12395;
  wire       [15:0]   _zz_12396;
  wire       [15:0]   _zz_12397;
  wire       [15:0]   _zz_12398;
  wire       [15:0]   _zz_12399;
  wire       [15:0]   _zz_12400;
  wire       [15:0]   _zz_12401;
  wire       [15:0]   _zz_12402;
  wire       [15:0]   _zz_12403;
  wire       [15:0]   _zz_12404;
  wire       [15:0]   _zz_12405;
  wire       [15:0]   _zz_12406;
  wire       [15:0]   _zz_12407;
  wire       [15:0]   _zz_12408;
  wire       [15:0]   _zz_12409;
  wire       [15:0]   _zz_12410;
  wire       [15:0]   _zz_12411;
  wire       [15:0]   _zz_12412;
  wire       [15:0]   _zz_12413;
  wire       [15:0]   _zz_12414;
  wire       [15:0]   _zz_12415;
  wire       [15:0]   _zz_12416;
  wire       [15:0]   _zz_12417;
  wire       [15:0]   _zz_12418;
  wire       [15:0]   _zz_12419;
  wire       [15:0]   _zz_12420;
  wire       [15:0]   _zz_12421;
  wire       [15:0]   _zz_12422;
  wire       [15:0]   _zz_12423;
  wire       [15:0]   _zz_12424;
  wire       [15:0]   _zz_12425;
  wire       [15:0]   _zz_12426;
  wire       [15:0]   _zz_12427;
  wire       [15:0]   _zz_12428;
  wire       [15:0]   _zz_12429;
  wire       [15:0]   _zz_12430;
  wire       [15:0]   _zz_12431;
  wire       [15:0]   _zz_12432;
  wire       [15:0]   _zz_12433;
  wire       [15:0]   _zz_12434;
  wire       [15:0]   _zz_12435;
  wire       [15:0]   _zz_12436;
  wire       [15:0]   _zz_12437;
  wire       [15:0]   _zz_12438;
  wire       [15:0]   _zz_12439;
  wire       [15:0]   _zz_12440;
  wire       [15:0]   _zz_12441;
  wire       [15:0]   _zz_12442;
  wire       [15:0]   _zz_12443;
  wire       [15:0]   _zz_12444;
  wire       [15:0]   _zz_12445;
  wire       [15:0]   _zz_12446;
  wire       [15:0]   _zz_12447;
  wire       [15:0]   _zz_12448;
  wire       [15:0]   _zz_12449;
  wire       [15:0]   _zz_12450;
  wire       [15:0]   _zz_12451;
  wire       [15:0]   _zz_12452;
  wire       [15:0]   _zz_12453;
  wire       [15:0]   _zz_12454;
  wire       [15:0]   _zz_12455;
  wire       [15:0]   _zz_12456;
  wire       [15:0]   _zz_12457;
  wire       [15:0]   _zz_12458;
  wire       [15:0]   _zz_12459;
  wire       [15:0]   _zz_12460;
  wire       [15:0]   _zz_12461;
  wire       [15:0]   _zz_12462;
  wire       [15:0]   _zz_12463;
  wire       [15:0]   _zz_12464;
  wire       [15:0]   _zz_12465;
  wire       [15:0]   _zz_12466;
  wire       [15:0]   _zz_12467;
  wire       [15:0]   _zz_12468;
  wire       [15:0]   _zz_12469;
  wire       [15:0]   _zz_12470;
  wire       [15:0]   _zz_12471;
  wire       [15:0]   _zz_12472;
  wire       [15:0]   _zz_12473;
  wire       [15:0]   _zz_12474;
  wire       [15:0]   _zz_12475;
  wire       [15:0]   _zz_12476;
  wire       [15:0]   _zz_12477;
  wire       [15:0]   _zz_12478;
  wire       [15:0]   _zz_12479;
  wire       [15:0]   _zz_12480;
  wire       [15:0]   _zz_12481;
  wire       [15:0]   _zz_12482;
  wire       [15:0]   _zz_12483;
  wire       [15:0]   _zz_12484;
  wire       [15:0]   _zz_12485;
  wire       [15:0]   _zz_12486;
  wire       [15:0]   _zz_12487;
  wire       [15:0]   _zz_12488;
  wire       [15:0]   _zz_12489;
  wire       [15:0]   _zz_12490;
  wire       [15:0]   _zz_12491;
  wire       [15:0]   _zz_12492;
  wire       [15:0]   _zz_12493;
  wire       [15:0]   _zz_12494;
  wire       [15:0]   _zz_12495;
  wire       [15:0]   _zz_12496;
  wire       [15:0]   _zz_12497;
  wire       [15:0]   _zz_12498;
  wire       [15:0]   _zz_12499;
  wire       [15:0]   _zz_12500;
  wire       [15:0]   _zz_12501;
  wire       [15:0]   _zz_12502;
  wire       [15:0]   _zz_12503;
  wire       [15:0]   _zz_12504;
  wire       [15:0]   _zz_12505;
  wire       [15:0]   _zz_12506;
  wire       [15:0]   _zz_12507;
  wire       [15:0]   _zz_12508;
  wire       [15:0]   _zz_12509;
  wire       [15:0]   _zz_12510;
  wire       [15:0]   _zz_12511;
  wire       [15:0]   _zz_12512;
  wire       [15:0]   _zz_12513;
  wire       [15:0]   _zz_12514;
  wire       [15:0]   _zz_12515;
  wire       [15:0]   _zz_12516;
  wire       [15:0]   _zz_12517;
  wire       [15:0]   _zz_12518;
  wire       [15:0]   _zz_12519;
  wire       [15:0]   _zz_12520;
  wire       [15:0]   _zz_12521;
  wire       [15:0]   _zz_12522;
  wire       [15:0]   _zz_12523;
  wire       [15:0]   _zz_12524;
  wire       [15:0]   _zz_12525;
  wire       [15:0]   _zz_12526;
  wire       [15:0]   _zz_12527;
  wire       [15:0]   _zz_12528;
  wire       [15:0]   _zz_12529;
  wire       [15:0]   _zz_12530;
  wire       [15:0]   _zz_12531;
  wire       [15:0]   _zz_12532;
  wire       [15:0]   _zz_12533;
  wire       [15:0]   _zz_12534;
  wire       [15:0]   _zz_12535;
  wire       [15:0]   _zz_12536;
  wire       [15:0]   _zz_12537;
  wire       [15:0]   _zz_12538;
  wire       [15:0]   _zz_12539;
  wire       [15:0]   _zz_12540;
  wire       [15:0]   _zz_12541;
  wire       [15:0]   _zz_12542;
  wire       [15:0]   _zz_12543;
  wire       [15:0]   _zz_12544;
  wire       [15:0]   _zz_12545;
  wire       [15:0]   _zz_12546;
  wire       [15:0]   _zz_12547;
  wire       [15:0]   _zz_12548;
  wire       [15:0]   _zz_12549;
  wire       [15:0]   _zz_12550;
  wire       [15:0]   _zz_12551;
  wire       [15:0]   _zz_12552;
  wire       [15:0]   _zz_12553;
  wire       [15:0]   _zz_12554;
  wire       [15:0]   _zz_12555;
  wire       [15:0]   _zz_12556;
  wire       [15:0]   _zz_12557;
  wire       [15:0]   _zz_12558;
  wire       [15:0]   _zz_12559;
  wire       [15:0]   _zz_12560;
  wire       [15:0]   _zz_12561;
  wire       [15:0]   _zz_12562;
  wire       [15:0]   _zz_12563;
  wire       [15:0]   _zz_12564;
  wire       [15:0]   _zz_12565;
  wire       [15:0]   _zz_12566;
  wire       [15:0]   _zz_12567;
  wire       [15:0]   _zz_12568;
  wire       [15:0]   _zz_12569;
  wire       [15:0]   _zz_12570;
  wire       [15:0]   _zz_12571;
  wire       [15:0]   _zz_12572;
  wire       [15:0]   _zz_12573;
  wire       [15:0]   _zz_12574;
  wire       [15:0]   _zz_12575;
  wire       [15:0]   _zz_12576;
  wire       [15:0]   _zz_12577;
  wire       [15:0]   _zz_12578;
  wire       [15:0]   _zz_12579;
  wire       [15:0]   _zz_12580;
  wire       [15:0]   _zz_12581;
  wire       [15:0]   _zz_12582;
  wire       [15:0]   _zz_12583;
  wire       [15:0]   _zz_12584;
  wire       [15:0]   _zz_12585;
  wire       [15:0]   _zz_12586;
  wire       [15:0]   _zz_12587;
  wire       [15:0]   _zz_12588;
  wire       [15:0]   _zz_12589;
  wire       [15:0]   _zz_12590;
  wire       [15:0]   _zz_12591;
  wire       [15:0]   _zz_12592;
  wire       [15:0]   _zz_12593;
  wire       [15:0]   _zz_12594;
  wire       [15:0]   _zz_12595;
  wire       [15:0]   _zz_12596;
  wire       [15:0]   _zz_12597;
  wire       [15:0]   _zz_12598;
  wire       [15:0]   _zz_12599;
  wire       [15:0]   _zz_12600;
  wire       [15:0]   _zz_12601;
  wire       [15:0]   _zz_12602;
  wire       [15:0]   _zz_12603;
  wire       [15:0]   _zz_12604;
  wire       [15:0]   _zz_12605;
  wire       [15:0]   _zz_12606;
  wire       [15:0]   _zz_12607;
  wire       [15:0]   _zz_12608;
  wire       [15:0]   _zz_12609;
  wire       [15:0]   _zz_12610;
  wire       [15:0]   _zz_12611;
  wire       [15:0]   _zz_12612;
  wire       [15:0]   _zz_12613;
  wire       [15:0]   _zz_12614;
  wire       [15:0]   _zz_12615;
  wire       [15:0]   _zz_12616;
  wire       [15:0]   _zz_12617;
  wire       [15:0]   _zz_12618;
  wire       [15:0]   _zz_12619;
  wire       [15:0]   _zz_12620;
  wire       [15:0]   _zz_12621;
  wire       [15:0]   _zz_12622;
  wire       [15:0]   _zz_12623;
  wire       [15:0]   _zz_12624;
  wire       [15:0]   _zz_12625;
  wire       [15:0]   _zz_12626;
  wire       [15:0]   _zz_12627;
  wire       [15:0]   _zz_12628;
  wire       [15:0]   _zz_12629;
  wire       [15:0]   _zz_12630;
  wire       [15:0]   _zz_12631;
  wire       [15:0]   _zz_12632;
  wire       [15:0]   _zz_12633;
  wire       [15:0]   _zz_12634;
  wire       [15:0]   _zz_12635;
  wire       [15:0]   _zz_12636;
  wire       [15:0]   _zz_12637;
  wire       [15:0]   _zz_12638;
  wire       [15:0]   _zz_12639;
  wire       [15:0]   _zz_12640;
  wire       [15:0]   _zz_12641;
  wire       [15:0]   _zz_12642;
  wire       [15:0]   _zz_12643;
  wire       [15:0]   _zz_12644;
  wire       [15:0]   _zz_12645;
  wire       [15:0]   _zz_12646;
  wire       [15:0]   _zz_12647;
  wire       [15:0]   _zz_12648;
  wire       [15:0]   _zz_12649;
  wire       [15:0]   _zz_12650;
  wire       [15:0]   _zz_12651;
  wire       [15:0]   _zz_12652;
  wire       [15:0]   _zz_12653;
  wire       [15:0]   _zz_12654;
  wire       [15:0]   _zz_12655;
  wire       [15:0]   _zz_12656;
  wire       [15:0]   _zz_12657;
  wire       [15:0]   _zz_12658;
  wire       [15:0]   _zz_12659;
  wire       [15:0]   _zz_12660;
  wire       [15:0]   _zz_12661;
  wire       [15:0]   _zz_12662;
  wire       [15:0]   _zz_12663;
  wire       [15:0]   _zz_12664;
  wire       [15:0]   _zz_12665;
  wire       [15:0]   _zz_12666;
  wire       [15:0]   _zz_12667;
  wire       [15:0]   _zz_12668;
  wire       [15:0]   _zz_12669;
  wire       [15:0]   _zz_12670;
  wire       [15:0]   _zz_12671;
  wire       [15:0]   _zz_12672;
  wire       [15:0]   _zz_12673;
  wire       [15:0]   _zz_12674;
  wire       [15:0]   _zz_12675;
  wire       [15:0]   _zz_12676;
  wire       [15:0]   _zz_12677;
  wire       [15:0]   _zz_12678;
  wire       [15:0]   _zz_12679;
  wire       [15:0]   _zz_12680;
  wire       [15:0]   _zz_12681;
  wire       [15:0]   _zz_12682;
  wire       [15:0]   _zz_12683;
  wire       [15:0]   _zz_12684;
  wire       [15:0]   _zz_12685;
  wire       [15:0]   _zz_12686;
  wire       [15:0]   _zz_12687;
  wire       [15:0]   _zz_12688;
  wire       [15:0]   _zz_12689;
  wire       [15:0]   _zz_12690;
  wire       [15:0]   _zz_12691;
  wire       [15:0]   _zz_12692;
  wire       [15:0]   _zz_12693;
  wire       [15:0]   _zz_12694;
  wire       [15:0]   _zz_12695;
  wire       [15:0]   _zz_12696;
  wire       [15:0]   _zz_12697;
  wire       [15:0]   _zz_12698;
  wire       [15:0]   _zz_12699;
  wire       [15:0]   _zz_12700;
  wire       [15:0]   _zz_12701;
  wire       [15:0]   _zz_12702;
  wire       [15:0]   _zz_12703;
  wire       [15:0]   _zz_12704;
  wire       [15:0]   _zz_12705;
  wire       [15:0]   _zz_12706;
  wire       [15:0]   _zz_12707;
  wire       [15:0]   _zz_12708;
  wire       [15:0]   _zz_12709;
  wire       [15:0]   _zz_12710;
  wire       [15:0]   _zz_12711;
  wire       [15:0]   _zz_12712;
  wire       [15:0]   _zz_12713;
  wire       [15:0]   _zz_12714;
  wire       [15:0]   _zz_12715;
  wire       [15:0]   _zz_12716;
  wire       [15:0]   _zz_12717;
  wire       [15:0]   _zz_12718;
  wire       [15:0]   _zz_12719;
  wire       [15:0]   _zz_12720;
  wire       [15:0]   _zz_12721;
  wire       [15:0]   _zz_12722;
  wire       [15:0]   _zz_12723;
  wire       [15:0]   _zz_12724;
  wire       [15:0]   _zz_12725;
  wire       [15:0]   _zz_12726;
  wire       [15:0]   _zz_12727;
  wire       [15:0]   _zz_12728;
  wire       [15:0]   _zz_12729;
  wire       [15:0]   _zz_12730;
  wire       [15:0]   _zz_12731;
  wire       [15:0]   _zz_12732;
  wire       [15:0]   _zz_12733;
  wire       [15:0]   _zz_12734;
  wire       [15:0]   _zz_12735;
  wire       [15:0]   _zz_12736;
  wire       [15:0]   _zz_12737;
  wire       [15:0]   _zz_12738;
  wire       [15:0]   _zz_12739;
  wire       [15:0]   _zz_12740;
  wire       [15:0]   _zz_12741;
  wire       [15:0]   _zz_12742;
  wire       [15:0]   _zz_12743;
  wire       [15:0]   _zz_12744;
  wire       [15:0]   _zz_12745;
  wire       [15:0]   _zz_12746;
  wire       [15:0]   _zz_12747;
  wire       [15:0]   _zz_12748;
  wire       [15:0]   _zz_12749;
  wire       [15:0]   _zz_12750;
  wire       [15:0]   _zz_12751;
  wire       [15:0]   _zz_12752;
  wire       [15:0]   _zz_12753;
  wire       [15:0]   _zz_12754;
  wire       [15:0]   _zz_12755;
  wire       [15:0]   _zz_12756;
  wire       [15:0]   _zz_12757;
  wire       [15:0]   _zz_12758;
  wire       [15:0]   _zz_12759;
  wire       [15:0]   _zz_12760;
  wire       [15:0]   _zz_12761;
  wire       [15:0]   _zz_12762;
  wire       [15:0]   _zz_12763;
  wire       [15:0]   _zz_12764;
  wire       [15:0]   _zz_12765;
  wire       [15:0]   _zz_12766;
  wire       [15:0]   _zz_12767;
  wire       [15:0]   _zz_12768;
  wire       [15:0]   _zz_12769;
  wire       [15:0]   _zz_12770;
  wire       [15:0]   _zz_12771;
  wire       [15:0]   _zz_12772;
  wire       [15:0]   _zz_12773;
  wire       [15:0]   _zz_12774;
  wire       [15:0]   _zz_12775;
  wire       [15:0]   _zz_12776;
  wire       [15:0]   _zz_12777;
  wire       [15:0]   _zz_12778;
  wire       [15:0]   _zz_12779;
  wire       [15:0]   _zz_12780;
  wire       [15:0]   _zz_12781;
  wire       [15:0]   _zz_12782;
  wire       [15:0]   _zz_12783;
  wire       [15:0]   _zz_12784;
  wire       [15:0]   _zz_12785;
  wire       [15:0]   _zz_12786;
  wire       [15:0]   _zz_12787;
  wire       [15:0]   _zz_12788;
  wire       [15:0]   _zz_12789;
  wire       [15:0]   _zz_12790;
  wire       [15:0]   _zz_12791;
  wire       [15:0]   _zz_12792;
  wire       [15:0]   _zz_12793;
  wire       [15:0]   _zz_12794;
  wire       [15:0]   _zz_12795;
  wire       [15:0]   _zz_12796;
  wire       [15:0]   _zz_12797;
  wire       [15:0]   _zz_12798;
  wire       [15:0]   _zz_12799;
  wire       [15:0]   _zz_12800;
  wire       [15:0]   _zz_12801;
  wire       [15:0]   _zz_12802;
  wire       [15:0]   _zz_12803;
  wire       [15:0]   _zz_12804;
  wire       [15:0]   _zz_12805;
  wire       [15:0]   _zz_12806;
  wire       [15:0]   _zz_12807;
  wire       [15:0]   _zz_12808;
  wire       [15:0]   _zz_12809;
  wire       [15:0]   _zz_12810;
  wire       [15:0]   _zz_12811;
  wire       [15:0]   _zz_12812;
  wire       [15:0]   _zz_12813;
  wire       [15:0]   _zz_12814;
  wire       [15:0]   _zz_12815;
  wire       [15:0]   _zz_12816;
  wire       [15:0]   _zz_12817;
  wire       [15:0]   _zz_12818;
  wire       [15:0]   _zz_12819;
  wire       [15:0]   _zz_12820;
  wire       [15:0]   _zz_12821;
  wire       [15:0]   _zz_12822;
  wire       [15:0]   _zz_12823;
  wire       [15:0]   _zz_12824;
  wire       [15:0]   _zz_12825;
  wire       [15:0]   _zz_12826;
  wire       [15:0]   _zz_12827;
  wire       [15:0]   _zz_12828;
  wire       [15:0]   _zz_12829;
  wire       [15:0]   _zz_12830;
  wire       [15:0]   _zz_12831;
  wire       [15:0]   _zz_12832;
  wire       [15:0]   _zz_12833;
  wire       [15:0]   _zz_12834;
  wire       [15:0]   _zz_12835;
  wire       [15:0]   _zz_12836;
  wire       [15:0]   _zz_12837;
  wire       [15:0]   _zz_12838;
  wire       [15:0]   _zz_12839;
  wire       [15:0]   _zz_12840;
  wire       [15:0]   _zz_12841;
  wire       [15:0]   _zz_12842;
  wire       [15:0]   _zz_12843;
  wire       [15:0]   _zz_12844;
  wire       [15:0]   _zz_12845;
  wire       [15:0]   _zz_12846;
  wire       [15:0]   _zz_12847;
  wire       [15:0]   _zz_12848;
  wire       [15:0]   _zz_12849;
  wire       [15:0]   _zz_12850;
  wire       [15:0]   _zz_12851;
  wire       [15:0]   _zz_12852;
  wire       [15:0]   _zz_12853;
  wire       [15:0]   _zz_12854;
  wire       [15:0]   _zz_12855;
  wire       [15:0]   _zz_12856;
  wire       [15:0]   _zz_12857;
  wire       [15:0]   _zz_12858;
  wire       [15:0]   _zz_12859;
  wire       [15:0]   _zz_12860;
  wire       [15:0]   _zz_12861;
  wire       [15:0]   _zz_12862;
  wire       [15:0]   _zz_12863;
  wire       [15:0]   _zz_12864;
  wire       [15:0]   _zz_12865;
  wire       [15:0]   _zz_12866;
  wire       [15:0]   _zz_12867;
  wire       [15:0]   _zz_12868;
  wire       [15:0]   _zz_12869;
  wire       [15:0]   _zz_12870;
  wire       [15:0]   _zz_12871;
  wire       [15:0]   _zz_12872;
  wire       [15:0]   _zz_12873;
  wire       [15:0]   _zz_12874;
  wire       [15:0]   _zz_12875;
  wire       [15:0]   _zz_12876;
  wire       [15:0]   _zz_12877;
  wire       [15:0]   _zz_12878;
  wire       [15:0]   _zz_12879;
  wire       [15:0]   _zz_12880;
  wire       [15:0]   _zz_12881;
  wire       [15:0]   _zz_12882;
  wire       [15:0]   _zz_12883;
  wire       [15:0]   _zz_12884;
  wire       [15:0]   _zz_12885;
  wire       [15:0]   _zz_12886;
  wire       [15:0]   _zz_12887;
  wire       [15:0]   _zz_12888;
  wire       [15:0]   _zz_12889;
  wire       [15:0]   _zz_12890;
  wire       [15:0]   _zz_12891;
  wire       [15:0]   _zz_12892;
  wire       [15:0]   _zz_12893;
  wire       [15:0]   _zz_12894;
  wire       [15:0]   _zz_12895;
  wire       [15:0]   _zz_12896;
  wire       [15:0]   _zz_12897;
  wire       [15:0]   _zz_12898;
  wire       [15:0]   _zz_12899;
  wire       [15:0]   _zz_12900;
  wire       [15:0]   _zz_12901;
  wire       [15:0]   _zz_12902;
  wire       [15:0]   _zz_12903;
  wire       [15:0]   _zz_12904;
  wire       [15:0]   _zz_12905;
  wire       [15:0]   _zz_12906;
  wire       [15:0]   _zz_12907;
  wire       [15:0]   _zz_12908;
  wire       [15:0]   _zz_12909;
  wire       [15:0]   _zz_12910;
  wire       [15:0]   _zz_12911;
  wire       [15:0]   _zz_12912;
  wire       [15:0]   _zz_12913;
  wire       [15:0]   _zz_12914;
  wire       [15:0]   _zz_12915;
  wire       [15:0]   _zz_12916;
  wire       [15:0]   _zz_12917;
  wire       [15:0]   _zz_12918;
  wire       [15:0]   _zz_12919;
  wire       [15:0]   _zz_12920;
  wire       [15:0]   _zz_12921;
  wire       [15:0]   _zz_12922;
  wire       [15:0]   _zz_12923;
  wire       [15:0]   _zz_12924;
  wire       [15:0]   _zz_12925;
  wire       [15:0]   _zz_12926;
  wire       [15:0]   _zz_12927;
  wire       [15:0]   _zz_12928;
  wire       [15:0]   _zz_12929;
  wire       [15:0]   _zz_12930;
  wire       [15:0]   _zz_12931;
  wire       [15:0]   _zz_12932;
  wire       [15:0]   _zz_12933;
  wire       [15:0]   _zz_12934;
  wire       [15:0]   _zz_12935;
  wire       [15:0]   _zz_12936;
  wire       [15:0]   _zz_12937;
  wire       [15:0]   _zz_12938;
  wire       [15:0]   _zz_12939;
  wire       [15:0]   _zz_12940;
  wire       [15:0]   _zz_12941;
  wire       [15:0]   _zz_12942;
  wire       [15:0]   _zz_12943;
  wire       [15:0]   _zz_12944;
  wire       [15:0]   _zz_12945;
  wire       [15:0]   _zz_12946;
  wire       [15:0]   _zz_12947;
  wire       [15:0]   _zz_12948;
  wire       [15:0]   _zz_12949;
  wire       [15:0]   _zz_12950;
  wire       [15:0]   _zz_12951;
  wire       [15:0]   _zz_12952;
  wire       [15:0]   _zz_12953;
  wire       [15:0]   _zz_12954;
  wire       [15:0]   _zz_12955;
  wire       [15:0]   _zz_12956;
  wire       [15:0]   _zz_12957;
  wire       [15:0]   _zz_12958;
  wire       [15:0]   _zz_12959;
  wire       [15:0]   _zz_12960;
  wire       [15:0]   _zz_12961;
  wire       [15:0]   _zz_12962;
  wire       [15:0]   _zz_12963;
  wire       [15:0]   _zz_12964;
  wire       [15:0]   _zz_12965;
  wire       [15:0]   _zz_12966;
  wire       [15:0]   _zz_12967;
  wire       [15:0]   _zz_12968;
  wire       [15:0]   _zz_12969;
  wire       [15:0]   _zz_12970;
  wire       [15:0]   _zz_12971;
  wire       [15:0]   _zz_12972;
  wire       [15:0]   _zz_12973;
  wire       [15:0]   _zz_12974;
  wire       [15:0]   _zz_12975;
  wire       [15:0]   _zz_12976;
  wire       [15:0]   _zz_12977;
  wire       [15:0]   _zz_12978;
  wire       [15:0]   _zz_12979;
  wire       [15:0]   _zz_12980;
  wire       [15:0]   _zz_12981;
  wire       [15:0]   _zz_12982;
  wire       [15:0]   _zz_12983;
  wire       [15:0]   _zz_12984;
  wire       [15:0]   _zz_12985;
  wire       [15:0]   _zz_12986;
  wire       [15:0]   _zz_12987;
  wire       [15:0]   _zz_12988;
  wire       [15:0]   _zz_12989;
  wire       [15:0]   _zz_12990;
  wire       [15:0]   _zz_12991;
  wire       [15:0]   _zz_12992;
  wire       [15:0]   _zz_12993;
  wire       [15:0]   _zz_12994;
  wire       [15:0]   _zz_12995;
  wire       [15:0]   _zz_12996;
  wire       [15:0]   _zz_12997;
  wire       [15:0]   _zz_12998;
  wire       [15:0]   _zz_12999;
  wire       [15:0]   _zz_13000;
  wire       [15:0]   _zz_13001;
  wire       [15:0]   _zz_13002;
  wire       [15:0]   _zz_13003;
  wire       [15:0]   _zz_13004;
  wire       [15:0]   _zz_13005;
  wire       [15:0]   _zz_13006;
  wire       [15:0]   _zz_13007;
  wire       [15:0]   _zz_13008;
  wire       [15:0]   _zz_13009;
  wire       [15:0]   _zz_13010;
  wire       [15:0]   _zz_13011;
  wire       [15:0]   _zz_13012;
  wire       [15:0]   _zz_13013;
  wire       [15:0]   _zz_13014;
  wire       [15:0]   _zz_13015;
  wire       [15:0]   _zz_13016;
  wire       [15:0]   _zz_13017;
  wire       [15:0]   _zz_13018;
  wire       [15:0]   _zz_13019;
  wire       [15:0]   _zz_13020;
  wire       [15:0]   _zz_13021;
  wire       [15:0]   _zz_13022;
  wire       [15:0]   _zz_13023;
  wire       [15:0]   _zz_13024;
  wire       [15:0]   _zz_13025;
  wire       [15:0]   _zz_13026;
  wire       [15:0]   _zz_13027;
  wire       [15:0]   _zz_13028;
  wire       [15:0]   _zz_13029;
  wire       [15:0]   _zz_13030;
  wire       [15:0]   _zz_13031;
  wire       [15:0]   _zz_13032;
  wire       [15:0]   _zz_13033;
  wire       [15:0]   _zz_13034;
  wire       [15:0]   _zz_13035;
  wire       [15:0]   _zz_13036;
  wire       [15:0]   _zz_13037;
  wire       [15:0]   _zz_13038;
  wire       [15:0]   _zz_13039;
  wire       [15:0]   _zz_13040;
  wire       [15:0]   _zz_13041;
  wire       [15:0]   _zz_13042;
  wire       [15:0]   _zz_13043;
  wire       [15:0]   _zz_13044;
  wire       [15:0]   _zz_13045;
  wire       [15:0]   _zz_13046;
  wire       [15:0]   _zz_13047;
  wire       [15:0]   _zz_13048;
  wire       [15:0]   _zz_13049;
  wire       [15:0]   _zz_13050;
  wire       [15:0]   _zz_13051;
  wire       [15:0]   _zz_13052;
  wire       [15:0]   _zz_13053;
  wire       [15:0]   _zz_13054;
  wire       [15:0]   _zz_13055;
  wire       [15:0]   _zz_13056;
  wire       [15:0]   _zz_13057;
  wire       [15:0]   _zz_13058;
  wire       [15:0]   _zz_13059;
  wire       [15:0]   _zz_13060;
  wire       [15:0]   _zz_13061;
  wire       [15:0]   _zz_13062;
  wire       [15:0]   _zz_13063;
  wire       [15:0]   _zz_13064;
  wire       [15:0]   _zz_13065;
  wire       [15:0]   _zz_13066;
  wire       [15:0]   _zz_13067;
  wire       [15:0]   _zz_13068;
  wire       [15:0]   _zz_13069;
  wire       [15:0]   _zz_13070;
  wire       [15:0]   _zz_13071;
  wire       [15:0]   _zz_13072;
  wire       [15:0]   _zz_13073;
  wire       [15:0]   _zz_13074;
  wire       [15:0]   _zz_13075;
  wire       [15:0]   _zz_13076;
  wire       [15:0]   _zz_13077;
  wire       [15:0]   _zz_13078;
  wire       [15:0]   _zz_13079;
  wire       [15:0]   _zz_13080;
  wire       [15:0]   _zz_13081;
  wire       [15:0]   _zz_13082;
  wire       [15:0]   _zz_13083;
  wire       [15:0]   _zz_13084;
  wire       [15:0]   _zz_13085;
  wire       [15:0]   _zz_13086;
  wire       [15:0]   _zz_13087;
  wire       [15:0]   _zz_13088;
  wire       [15:0]   _zz_13089;
  wire       [15:0]   _zz_13090;
  wire       [15:0]   _zz_13091;
  wire       [15:0]   _zz_13092;
  wire       [15:0]   _zz_13093;
  wire       [15:0]   _zz_13094;
  wire       [15:0]   _zz_13095;
  wire       [15:0]   _zz_13096;
  wire       [15:0]   _zz_13097;
  wire       [15:0]   _zz_13098;
  wire       [15:0]   _zz_13099;
  wire       [15:0]   _zz_13100;
  wire       [15:0]   _zz_13101;
  wire       [15:0]   _zz_13102;
  wire       [15:0]   _zz_13103;
  wire       [15:0]   _zz_13104;
  wire       [15:0]   _zz_13105;
  wire       [15:0]   _zz_13106;
  wire       [15:0]   _zz_13107;
  wire       [15:0]   _zz_13108;
  wire       [15:0]   _zz_13109;
  wire       [15:0]   _zz_13110;
  wire       [15:0]   _zz_13111;
  wire       [15:0]   _zz_13112;
  wire       [15:0]   _zz_13113;
  wire       [15:0]   _zz_13114;
  wire       [15:0]   _zz_13115;
  wire       [15:0]   _zz_13116;
  wire       [15:0]   _zz_13117;
  wire       [15:0]   _zz_13118;
  wire       [15:0]   _zz_13119;
  wire       [15:0]   _zz_13120;
  wire       [15:0]   _zz_13121;
  wire       [15:0]   _zz_13122;
  wire       [15:0]   _zz_13123;
  wire       [15:0]   _zz_13124;
  wire       [15:0]   _zz_13125;
  wire       [15:0]   _zz_13126;
  wire       [15:0]   _zz_13127;
  wire       [15:0]   _zz_13128;
  wire       [15:0]   _zz_13129;
  wire       [15:0]   _zz_13130;
  wire       [15:0]   _zz_13131;
  wire       [15:0]   _zz_13132;
  wire       [15:0]   _zz_13133;
  wire       [15:0]   _zz_13134;
  wire       [15:0]   _zz_13135;
  wire       [15:0]   _zz_13136;
  wire       [15:0]   _zz_13137;
  wire       [15:0]   _zz_13138;
  wire       [15:0]   _zz_13139;
  wire       [15:0]   _zz_13140;
  wire       [15:0]   _zz_13141;
  wire       [15:0]   _zz_13142;
  wire       [15:0]   _zz_13143;
  wire       [15:0]   _zz_13144;
  wire       [15:0]   _zz_13145;
  wire       [15:0]   _zz_13146;
  wire       [15:0]   _zz_13147;
  wire       [15:0]   _zz_13148;
  wire       [15:0]   _zz_13149;
  wire       [15:0]   _zz_13150;
  wire       [15:0]   _zz_13151;
  wire       [15:0]   _zz_13152;
  wire       [15:0]   _zz_13153;
  wire       [15:0]   _zz_13154;
  wire       [15:0]   _zz_13155;
  wire       [15:0]   _zz_13156;
  wire       [15:0]   _zz_13157;
  wire       [15:0]   _zz_13158;
  wire       [15:0]   _zz_13159;
  wire       [15:0]   _zz_13160;
  wire       [15:0]   _zz_13161;
  wire       [15:0]   _zz_13162;
  wire       [15:0]   _zz_13163;
  wire       [15:0]   _zz_13164;
  wire       [15:0]   _zz_13165;
  wire       [15:0]   _zz_13166;
  wire       [15:0]   _zz_13167;
  wire       [15:0]   _zz_13168;
  wire       [15:0]   _zz_13169;
  wire       [15:0]   _zz_13170;
  wire       [15:0]   _zz_13171;
  wire       [15:0]   _zz_13172;
  wire       [15:0]   _zz_13173;
  wire       [15:0]   _zz_13174;
  wire       [15:0]   _zz_13175;
  wire       [15:0]   _zz_13176;
  wire       [15:0]   _zz_13177;
  wire       [15:0]   _zz_13178;
  wire       [15:0]   _zz_13179;
  wire       [15:0]   _zz_13180;
  wire       [15:0]   _zz_13181;
  wire       [15:0]   _zz_13182;
  wire       [15:0]   _zz_13183;
  wire       [15:0]   _zz_13184;
  wire       [15:0]   _zz_13185;
  wire       [15:0]   _zz_13186;
  wire       [15:0]   _zz_13187;
  wire       [15:0]   _zz_13188;
  wire       [15:0]   _zz_13189;
  wire       [15:0]   _zz_13190;
  wire       [15:0]   _zz_13191;
  wire       [15:0]   _zz_13192;
  wire       [15:0]   _zz_13193;
  wire       [15:0]   _zz_13194;
  wire       [15:0]   _zz_13195;
  wire       [15:0]   _zz_13196;
  wire       [15:0]   _zz_13197;
  wire       [15:0]   _zz_13198;
  wire       [15:0]   _zz_13199;
  wire       [15:0]   _zz_13200;
  wire       [15:0]   _zz_13201;
  wire       [15:0]   _zz_13202;
  wire       [15:0]   _zz_13203;
  wire       [15:0]   _zz_13204;
  wire       [15:0]   _zz_13205;
  wire       [15:0]   _zz_13206;
  wire       [15:0]   _zz_13207;
  wire       [15:0]   _zz_13208;
  wire       [15:0]   _zz_13209;
  wire       [15:0]   _zz_13210;
  wire       [15:0]   _zz_13211;
  wire       [15:0]   _zz_13212;
  wire       [15:0]   _zz_13213;
  wire       [15:0]   _zz_13214;
  wire       [15:0]   _zz_13215;
  wire       [15:0]   _zz_13216;
  wire       [15:0]   _zz_13217;
  wire       [15:0]   _zz_13218;
  wire       [15:0]   _zz_13219;
  wire       [15:0]   _zz_13220;
  wire       [15:0]   _zz_13221;
  wire       [15:0]   _zz_13222;
  wire       [15:0]   _zz_13223;
  wire       [15:0]   _zz_13224;
  wire       [15:0]   _zz_13225;
  wire       [15:0]   _zz_13226;
  wire       [15:0]   _zz_13227;
  wire       [15:0]   _zz_13228;
  wire       [15:0]   _zz_13229;
  wire       [15:0]   _zz_13230;
  wire       [15:0]   _zz_13231;
  wire       [15:0]   _zz_13232;
  wire       [15:0]   _zz_13233;
  wire       [15:0]   _zz_13234;
  wire       [15:0]   _zz_13235;
  wire       [15:0]   _zz_13236;
  wire       [15:0]   _zz_13237;
  wire       [15:0]   _zz_13238;
  wire       [15:0]   _zz_13239;
  wire       [15:0]   _zz_13240;
  wire       [15:0]   _zz_13241;
  wire       [15:0]   _zz_13242;
  wire       [15:0]   _zz_13243;
  wire       [15:0]   _zz_13244;
  wire       [15:0]   _zz_13245;
  wire       [15:0]   _zz_13246;
  wire       [15:0]   _zz_13247;
  wire       [15:0]   _zz_13248;
  wire       [15:0]   _zz_13249;
  wire       [15:0]   _zz_13250;
  wire       [15:0]   _zz_13251;
  wire       [15:0]   _zz_13252;
  wire       [15:0]   _zz_13253;
  wire       [15:0]   _zz_13254;
  wire       [15:0]   _zz_13255;
  wire       [15:0]   _zz_13256;
  wire       [15:0]   _zz_13257;
  wire       [15:0]   _zz_13258;
  wire       [15:0]   _zz_13259;
  wire       [15:0]   _zz_13260;
  wire       [15:0]   _zz_13261;
  wire       [15:0]   _zz_13262;
  wire       [15:0]   _zz_13263;
  wire       [15:0]   _zz_13264;
  wire       [15:0]   _zz_13265;
  wire       [15:0]   _zz_13266;
  wire       [15:0]   _zz_13267;
  wire       [15:0]   _zz_13268;
  wire       [15:0]   _zz_13269;
  wire       [15:0]   _zz_13270;
  wire       [15:0]   _zz_13271;
  wire       [15:0]   _zz_13272;
  wire       [15:0]   _zz_13273;
  wire       [15:0]   _zz_13274;
  wire       [15:0]   _zz_13275;
  wire       [15:0]   _zz_13276;
  wire       [15:0]   _zz_13277;
  wire       [15:0]   _zz_13278;
  wire       [15:0]   _zz_13279;
  wire       [15:0]   _zz_13280;
  wire       [15:0]   _zz_13281;
  wire       [15:0]   _zz_13282;
  wire       [15:0]   _zz_13283;
  wire       [15:0]   _zz_13284;
  wire       [15:0]   _zz_13285;
  wire       [15:0]   _zz_13286;
  wire       [15:0]   _zz_13287;
  wire       [15:0]   _zz_13288;
  wire       [15:0]   _zz_13289;
  wire       [15:0]   _zz_13290;
  wire       [15:0]   _zz_13291;
  wire       [15:0]   _zz_13292;
  wire       [15:0]   _zz_13293;
  wire       [15:0]   _zz_13294;
  wire       [15:0]   _zz_13295;
  wire       [15:0]   _zz_13296;
  wire       [15:0]   _zz_13297;
  wire       [15:0]   _zz_13298;
  wire       [15:0]   _zz_13299;
  wire       [15:0]   _zz_13300;
  wire       [15:0]   _zz_13301;
  wire       [15:0]   _zz_13302;
  wire       [15:0]   _zz_13303;
  wire       [15:0]   _zz_13304;
  wire       [15:0]   _zz_13305;
  wire       [15:0]   _zz_13306;
  wire       [15:0]   _zz_13307;
  wire       [15:0]   _zz_13308;
  wire       [15:0]   _zz_13309;
  wire       [15:0]   _zz_13310;
  wire       [15:0]   _zz_13311;
  wire       [15:0]   _zz_13312;
  wire       [15:0]   _zz_13313;
  wire       [15:0]   _zz_13314;
  wire       [15:0]   _zz_13315;
  wire       [15:0]   _zz_13316;
  wire       [15:0]   _zz_13317;
  wire       [15:0]   _zz_13318;
  wire       [15:0]   _zz_13319;
  wire       [15:0]   _zz_13320;
  wire       [15:0]   _zz_13321;
  wire       [15:0]   _zz_13322;
  wire       [15:0]   _zz_13323;
  wire       [15:0]   _zz_13324;
  wire       [15:0]   _zz_13325;
  wire       [15:0]   _zz_13326;
  wire       [15:0]   _zz_13327;
  wire       [15:0]   _zz_13328;
  wire       [15:0]   _zz_13329;
  wire       [15:0]   _zz_13330;
  wire       [15:0]   _zz_13331;
  wire       [15:0]   _zz_13332;
  wire       [15:0]   _zz_13333;
  wire       [15:0]   _zz_13334;
  wire       [15:0]   _zz_13335;
  wire       [15:0]   _zz_13336;
  wire       [15:0]   _zz_13337;
  wire       [15:0]   _zz_13338;
  wire       [15:0]   _zz_13339;
  wire       [15:0]   _zz_13340;
  wire       [15:0]   _zz_13341;
  wire       [15:0]   _zz_13342;
  wire       [15:0]   _zz_13343;
  wire       [15:0]   _zz_13344;
  wire       [15:0]   _zz_13345;
  wire       [15:0]   _zz_13346;
  wire       [15:0]   _zz_13347;
  wire       [15:0]   _zz_13348;
  wire       [15:0]   _zz_13349;
  wire       [15:0]   _zz_13350;
  wire       [15:0]   _zz_13351;
  wire       [15:0]   _zz_13352;
  wire       [15:0]   _zz_13353;
  wire       [15:0]   _zz_13354;
  wire       [15:0]   _zz_13355;
  wire       [15:0]   _zz_13356;
  wire       [15:0]   _zz_13357;
  wire       [15:0]   _zz_13358;
  wire       [15:0]   _zz_13359;
  wire       [15:0]   _zz_13360;
  wire       [15:0]   _zz_13361;
  wire       [15:0]   _zz_13362;
  wire       [15:0]   _zz_13363;
  wire       [15:0]   _zz_13364;
  wire       [15:0]   _zz_13365;
  wire       [15:0]   _zz_13366;
  wire       [15:0]   _zz_13367;
  wire       [15:0]   _zz_13368;
  wire       [15:0]   _zz_13369;
  wire       [15:0]   _zz_13370;
  wire       [15:0]   _zz_13371;
  wire       [15:0]   _zz_13372;
  wire       [15:0]   _zz_13373;
  wire       [15:0]   _zz_13374;
  wire       [15:0]   _zz_13375;
  wire       [15:0]   _zz_13376;
  wire       [15:0]   _zz_13377;
  wire       [15:0]   _zz_13378;
  wire       [15:0]   _zz_13379;
  wire       [15:0]   _zz_13380;
  wire       [15:0]   _zz_13381;
  wire       [15:0]   _zz_13382;
  wire       [15:0]   _zz_13383;
  wire       [15:0]   _zz_13384;
  wire       [15:0]   _zz_13385;
  wire       [15:0]   _zz_13386;
  wire       [15:0]   _zz_13387;
  wire       [15:0]   _zz_13388;
  wire       [15:0]   _zz_13389;
  wire       [15:0]   _zz_13390;
  wire       [15:0]   _zz_13391;
  wire       [15:0]   _zz_13392;
  wire       [15:0]   _zz_13393;
  wire       [15:0]   _zz_13394;
  wire       [15:0]   _zz_13395;
  wire       [15:0]   _zz_13396;
  wire       [15:0]   _zz_13397;
  wire       [15:0]   _zz_13398;
  wire       [15:0]   _zz_13399;
  wire       [15:0]   _zz_13400;
  wire       [15:0]   _zz_13401;
  wire       [15:0]   _zz_13402;
  wire       [15:0]   _zz_13403;
  wire       [15:0]   _zz_13404;
  wire       [15:0]   _zz_13405;
  wire       [15:0]   _zz_13406;
  wire       [15:0]   _zz_13407;
  wire       [15:0]   _zz_13408;
  wire       [15:0]   _zz_13409;
  wire       [15:0]   _zz_13410;
  wire       [15:0]   _zz_13411;
  wire       [15:0]   _zz_13412;
  wire       [15:0]   _zz_13413;
  wire       [15:0]   _zz_13414;
  wire       [15:0]   _zz_13415;
  wire       [15:0]   _zz_13416;
  wire       [15:0]   _zz_13417;
  wire       [15:0]   _zz_13418;
  wire       [15:0]   _zz_13419;
  wire       [15:0]   _zz_13420;
  wire       [15:0]   _zz_13421;
  wire       [15:0]   _zz_13422;
  wire       [15:0]   _zz_13423;
  wire       [15:0]   _zz_13424;
  wire       [15:0]   _zz_13425;
  wire       [15:0]   _zz_13426;
  wire       [15:0]   _zz_13427;
  wire       [15:0]   _zz_13428;
  wire       [15:0]   _zz_13429;
  wire       [15:0]   _zz_13430;
  wire       [15:0]   _zz_13431;
  wire       [15:0]   _zz_13432;
  wire       [15:0]   _zz_13433;
  wire       [15:0]   _zz_13434;
  wire       [15:0]   _zz_13435;
  wire       [15:0]   _zz_13436;
  wire       [15:0]   _zz_13437;
  wire       [15:0]   _zz_13438;
  wire       [15:0]   _zz_13439;
  wire       [15:0]   _zz_13440;
  wire       [15:0]   _zz_13441;
  wire       [15:0]   _zz_13442;
  wire       [15:0]   _zz_13443;
  wire       [15:0]   _zz_13444;
  wire       [15:0]   _zz_13445;
  wire       [15:0]   _zz_13446;
  wire       [15:0]   _zz_13447;
  wire       [15:0]   _zz_13448;
  wire       [15:0]   _zz_13449;
  wire       [15:0]   _zz_13450;
  wire       [15:0]   _zz_13451;
  wire       [15:0]   _zz_13452;
  wire       [15:0]   _zz_13453;
  wire       [15:0]   _zz_13454;
  wire       [15:0]   _zz_13455;
  wire       [15:0]   _zz_13456;
  wire       [15:0]   _zz_13457;
  wire       [15:0]   _zz_13458;
  wire       [15:0]   _zz_13459;
  wire       [15:0]   _zz_13460;
  wire       [15:0]   _zz_13461;
  wire       [15:0]   _zz_13462;
  wire       [15:0]   _zz_13463;
  wire       [15:0]   _zz_13464;
  wire       [15:0]   _zz_13465;
  wire       [15:0]   _zz_13466;
  wire       [15:0]   _zz_13467;
  wire       [15:0]   _zz_13468;
  wire       [15:0]   _zz_13469;
  wire       [15:0]   _zz_13470;
  wire       [15:0]   _zz_13471;
  wire       [15:0]   _zz_13472;
  wire       [15:0]   _zz_13473;
  wire       [15:0]   _zz_13474;
  wire       [15:0]   _zz_13475;
  wire       [15:0]   _zz_13476;
  wire       [15:0]   _zz_13477;
  wire       [15:0]   _zz_13478;
  wire       [15:0]   _zz_13479;
  wire       [15:0]   _zz_13480;
  wire       [15:0]   _zz_13481;
  wire       [15:0]   _zz_13482;
  wire       [15:0]   _zz_13483;
  wire       [15:0]   _zz_13484;
  wire       [15:0]   _zz_13485;
  wire       [15:0]   _zz_13486;
  wire       [15:0]   _zz_13487;
  wire       [15:0]   _zz_13488;
  wire       [15:0]   _zz_13489;
  wire       [15:0]   _zz_13490;
  wire       [15:0]   _zz_13491;
  wire       [15:0]   _zz_13492;
  wire       [15:0]   _zz_13493;
  wire       [15:0]   _zz_13494;
  wire       [15:0]   _zz_13495;
  wire       [15:0]   _zz_13496;
  wire       [15:0]   _zz_13497;
  wire       [15:0]   _zz_13498;
  wire       [15:0]   _zz_13499;
  wire       [15:0]   _zz_13500;
  wire       [15:0]   _zz_13501;
  wire       [15:0]   _zz_13502;
  wire       [15:0]   _zz_13503;
  wire       [15:0]   _zz_13504;
  wire       [15:0]   _zz_13505;
  wire       [15:0]   _zz_13506;
  wire       [15:0]   _zz_13507;
  wire       [15:0]   _zz_13508;
  wire       [15:0]   _zz_13509;
  wire       [15:0]   _zz_13510;
  wire       [15:0]   _zz_13511;
  wire       [15:0]   _zz_13512;
  wire       [15:0]   _zz_13513;
  wire       [15:0]   _zz_13514;
  wire       [15:0]   _zz_13515;
  wire       [15:0]   _zz_13516;
  wire       [15:0]   _zz_13517;
  wire       [15:0]   _zz_13518;
  wire       [15:0]   _zz_13519;
  wire       [15:0]   _zz_13520;
  wire       [15:0]   _zz_13521;
  wire       [15:0]   _zz_13522;
  wire       [15:0]   _zz_13523;
  wire       [15:0]   _zz_13524;
  wire       [15:0]   _zz_13525;
  wire       [15:0]   _zz_13526;
  wire       [15:0]   _zz_13527;
  wire       [15:0]   _zz_13528;
  wire       [15:0]   _zz_13529;
  wire       [15:0]   _zz_13530;
  wire       [15:0]   _zz_13531;
  wire       [15:0]   _zz_13532;
  wire       [15:0]   _zz_13533;
  wire       [15:0]   _zz_13534;
  wire       [15:0]   _zz_13535;
  wire       [15:0]   _zz_13536;
  wire       [15:0]   _zz_13537;
  wire       [15:0]   _zz_13538;
  wire       [15:0]   _zz_13539;
  wire       [15:0]   _zz_13540;
  wire       [15:0]   _zz_13541;
  wire       [15:0]   _zz_13542;
  wire       [15:0]   _zz_13543;
  wire       [15:0]   _zz_13544;
  wire       [15:0]   _zz_13545;
  wire       [15:0]   _zz_13546;
  wire       [15:0]   _zz_13547;
  wire       [15:0]   _zz_13548;
  wire       [15:0]   _zz_13549;
  wire       [15:0]   _zz_13550;
  wire       [15:0]   _zz_13551;
  wire       [15:0]   _zz_13552;
  wire       [15:0]   _zz_13553;
  wire       [15:0]   _zz_13554;
  wire       [15:0]   _zz_13555;
  wire       [15:0]   _zz_13556;
  wire       [15:0]   _zz_13557;
  wire       [15:0]   _zz_13558;
  wire       [15:0]   _zz_13559;
  wire       [15:0]   _zz_13560;
  wire       [15:0]   _zz_13561;
  wire       [15:0]   _zz_13562;
  wire       [15:0]   _zz_13563;
  wire       [15:0]   _zz_13564;
  wire       [15:0]   _zz_13565;
  wire       [15:0]   _zz_13566;
  wire       [15:0]   _zz_13567;
  wire       [15:0]   _zz_13568;
  wire       [15:0]   _zz_13569;
  wire       [15:0]   _zz_13570;
  wire       [15:0]   _zz_13571;
  wire       [15:0]   _zz_13572;
  wire       [15:0]   _zz_13573;
  wire       [15:0]   _zz_13574;
  wire       [15:0]   _zz_13575;
  wire       [15:0]   _zz_13576;
  wire       [15:0]   _zz_13577;
  wire       [15:0]   _zz_13578;
  wire       [15:0]   _zz_13579;
  wire       [15:0]   _zz_13580;
  wire       [15:0]   _zz_13581;
  wire       [15:0]   _zz_13582;
  wire       [15:0]   _zz_13583;
  wire       [15:0]   _zz_13584;
  wire       [15:0]   _zz_13585;
  wire       [15:0]   _zz_13586;
  wire       [15:0]   _zz_13587;
  wire       [15:0]   _zz_13588;
  wire       [15:0]   _zz_13589;
  wire       [15:0]   _zz_13590;
  wire       [15:0]   _zz_13591;
  wire       [15:0]   _zz_13592;
  wire       [15:0]   _zz_13593;
  wire       [15:0]   _zz_13594;
  wire       [15:0]   _zz_13595;
  wire       [15:0]   _zz_13596;
  wire       [15:0]   _zz_13597;
  wire       [15:0]   _zz_13598;
  wire       [15:0]   _zz_13599;
  wire       [15:0]   _zz_13600;
  wire       [15:0]   _zz_13601;
  wire       [15:0]   _zz_13602;
  wire       [15:0]   _zz_13603;
  wire       [15:0]   _zz_13604;
  wire       [15:0]   _zz_13605;
  wire       [15:0]   _zz_13606;
  wire       [15:0]   _zz_13607;
  wire       [15:0]   _zz_13608;
  wire       [15:0]   _zz_13609;
  wire       [15:0]   _zz_13610;
  wire       [15:0]   _zz_13611;
  wire       [15:0]   _zz_13612;
  wire       [15:0]   _zz_13613;
  wire       [15:0]   _zz_13614;
  wire       [15:0]   _zz_13615;
  wire       [15:0]   _zz_13616;
  wire       [15:0]   _zz_13617;
  wire       [15:0]   _zz_13618;
  wire       [15:0]   _zz_13619;
  wire       [15:0]   _zz_13620;
  wire       [15:0]   _zz_13621;
  wire       [15:0]   _zz_13622;
  wire       [15:0]   _zz_13623;
  wire       [15:0]   _zz_13624;
  wire       [15:0]   _zz_13625;
  wire       [15:0]   _zz_13626;
  wire       [15:0]   _zz_13627;
  wire       [15:0]   _zz_13628;
  wire       [15:0]   _zz_13629;
  wire       [15:0]   _zz_13630;
  wire       [15:0]   _zz_13631;
  wire       [15:0]   _zz_13632;
  wire       [15:0]   _zz_13633;
  wire       [15:0]   _zz_13634;
  wire       [15:0]   _zz_13635;
  wire       [15:0]   _zz_13636;
  wire       [15:0]   _zz_13637;
  wire       [15:0]   _zz_13638;
  wire       [15:0]   _zz_13639;
  wire       [15:0]   _zz_13640;
  wire       [15:0]   _zz_13641;
  wire       [15:0]   _zz_13642;
  wire       [15:0]   _zz_13643;
  wire       [15:0]   _zz_13644;
  wire       [15:0]   _zz_13645;
  wire       [15:0]   _zz_13646;
  wire       [15:0]   _zz_13647;
  wire       [15:0]   _zz_13648;
  wire       [15:0]   _zz_13649;
  wire       [15:0]   _zz_13650;
  wire       [15:0]   _zz_13651;
  wire       [15:0]   _zz_13652;
  wire       [15:0]   _zz_13653;
  wire       [15:0]   _zz_13654;
  wire       [15:0]   _zz_13655;
  wire       [15:0]   _zz_13656;
  wire       [15:0]   _zz_13657;
  wire       [15:0]   _zz_13658;
  wire       [15:0]   _zz_13659;
  wire       [15:0]   _zz_13660;
  wire       [15:0]   _zz_13661;
  wire       [15:0]   _zz_13662;
  wire       [15:0]   _zz_13663;
  wire       [15:0]   _zz_13664;
  wire       [15:0]   _zz_13665;
  wire       [15:0]   _zz_13666;
  wire       [15:0]   _zz_13667;
  wire       [15:0]   _zz_13668;
  wire       [15:0]   _zz_13669;
  wire       [15:0]   _zz_13670;
  wire       [15:0]   _zz_13671;
  wire       [15:0]   _zz_13672;
  wire       [15:0]   _zz_13673;
  wire       [15:0]   _zz_13674;
  wire       [15:0]   _zz_13675;
  wire       [15:0]   _zz_13676;
  wire       [15:0]   _zz_13677;
  wire       [15:0]   _zz_13678;
  wire       [15:0]   _zz_13679;
  wire       [15:0]   _zz_13680;
  wire       [15:0]   _zz_13681;
  wire       [15:0]   _zz_13682;
  wire       [15:0]   _zz_13683;
  wire       [15:0]   _zz_13684;
  wire       [15:0]   _zz_13685;
  wire       [15:0]   _zz_13686;
  wire       [15:0]   _zz_13687;
  wire       [15:0]   _zz_13688;
  wire       [15:0]   _zz_13689;
  wire       [15:0]   _zz_13690;
  wire       [15:0]   _zz_13691;
  wire       [15:0]   _zz_13692;
  wire       [15:0]   _zz_13693;
  wire       [15:0]   _zz_13694;
  wire       [15:0]   _zz_13695;
  wire       [15:0]   _zz_13696;
  wire       [15:0]   _zz_13697;
  wire       [15:0]   _zz_13698;
  wire       [15:0]   _zz_13699;
  wire       [15:0]   _zz_13700;
  wire       [15:0]   _zz_13701;
  wire       [15:0]   _zz_13702;
  wire       [15:0]   _zz_13703;
  wire       [15:0]   _zz_13704;
  wire       [15:0]   _zz_13705;
  wire       [15:0]   _zz_13706;
  wire       [15:0]   _zz_13707;
  wire       [15:0]   _zz_13708;
  wire       [15:0]   _zz_13709;
  wire       [15:0]   _zz_13710;
  wire       [15:0]   _zz_13711;
  wire       [15:0]   _zz_13712;
  wire       [15:0]   _zz_13713;
  wire       [15:0]   _zz_13714;
  wire       [15:0]   _zz_13715;
  wire       [15:0]   _zz_13716;
  wire       [15:0]   _zz_13717;
  wire       [15:0]   _zz_13718;
  wire       [15:0]   _zz_13719;
  wire       [15:0]   _zz_13720;
  wire       [15:0]   _zz_13721;
  wire       [15:0]   _zz_13722;
  wire       [15:0]   _zz_13723;
  wire       [15:0]   _zz_13724;
  wire       [15:0]   _zz_13725;
  wire       [15:0]   _zz_13726;
  wire       [15:0]   _zz_13727;
  wire       [15:0]   _zz_13728;
  wire       [15:0]   _zz_13729;
  wire       [15:0]   _zz_13730;
  wire       [15:0]   _zz_13731;
  wire       [15:0]   _zz_13732;
  wire       [15:0]   _zz_13733;
  wire       [15:0]   _zz_13734;
  wire       [15:0]   _zz_13735;
  wire       [15:0]   _zz_13736;
  wire       [15:0]   _zz_13737;
  wire       [15:0]   _zz_13738;
  wire       [15:0]   _zz_13739;
  wire       [15:0]   _zz_13740;
  wire       [15:0]   _zz_13741;
  wire       [15:0]   _zz_13742;
  wire       [15:0]   _zz_13743;
  wire       [15:0]   _zz_13744;
  wire       [15:0]   _zz_13745;
  wire       [15:0]   _zz_13746;
  wire       [15:0]   _zz_13747;
  wire       [15:0]   _zz_13748;
  wire       [15:0]   _zz_13749;
  wire       [15:0]   _zz_13750;
  wire       [15:0]   _zz_13751;
  wire       [15:0]   _zz_13752;
  wire       [15:0]   _zz_13753;
  wire       [15:0]   _zz_13754;
  wire       [15:0]   _zz_13755;
  wire       [15:0]   _zz_13756;
  wire       [15:0]   _zz_13757;
  wire       [15:0]   _zz_13758;
  wire       [15:0]   _zz_13759;
  wire       [15:0]   _zz_13760;
  wire       [15:0]   _zz_13761;
  wire       [15:0]   _zz_13762;
  wire       [15:0]   _zz_13763;
  wire       [15:0]   _zz_13764;
  wire       [15:0]   _zz_13765;
  wire       [15:0]   _zz_13766;
  wire       [15:0]   _zz_13767;
  wire       [15:0]   _zz_13768;
  wire       [15:0]   _zz_13769;
  wire       [15:0]   _zz_13770;
  wire       [15:0]   _zz_13771;
  wire       [15:0]   _zz_13772;
  wire       [15:0]   _zz_13773;
  wire       [15:0]   _zz_13774;
  wire       [15:0]   _zz_13775;
  wire       [15:0]   _zz_13776;
  wire       [15:0]   _zz_13777;
  wire       [15:0]   _zz_13778;
  wire       [15:0]   _zz_13779;
  wire       [15:0]   _zz_13780;
  wire       [15:0]   _zz_13781;
  wire       [15:0]   _zz_13782;
  wire       [15:0]   _zz_13783;
  wire       [15:0]   _zz_13784;
  wire       [15:0]   _zz_13785;
  wire       [15:0]   _zz_13786;
  wire       [15:0]   _zz_13787;
  wire       [15:0]   _zz_13788;
  wire       [15:0]   _zz_13789;
  wire       [15:0]   _zz_13790;
  wire       [15:0]   _zz_13791;
  wire       [15:0]   _zz_13792;
  wire       [15:0]   _zz_13793;
  wire       [15:0]   _zz_13794;
  wire       [15:0]   _zz_13795;
  wire       [15:0]   _zz_13796;
  wire       [15:0]   _zz_13797;
  wire       [15:0]   _zz_13798;
  wire       [15:0]   _zz_13799;
  wire       [15:0]   _zz_13800;
  wire       [15:0]   _zz_13801;
  wire       [15:0]   _zz_13802;
  wire       [15:0]   _zz_13803;
  wire       [15:0]   _zz_13804;
  wire       [15:0]   _zz_13805;
  wire       [15:0]   _zz_13806;
  wire       [15:0]   _zz_13807;
  wire       [15:0]   _zz_13808;
  wire       [15:0]   _zz_13809;
  wire       [15:0]   _zz_13810;
  wire       [15:0]   _zz_13811;
  wire       [15:0]   _zz_13812;
  wire       [15:0]   _zz_13813;
  wire       [15:0]   _zz_13814;
  wire       [15:0]   _zz_13815;
  wire       [15:0]   _zz_13816;
  wire       [15:0]   _zz_13817;
  wire       [15:0]   _zz_13818;
  wire       [15:0]   _zz_13819;
  wire       [15:0]   _zz_13820;
  wire       [15:0]   _zz_13821;
  wire       [15:0]   _zz_13822;
  wire       [15:0]   _zz_13823;
  wire       [15:0]   _zz_13824;
  wire       [15:0]   _zz_13825;
  wire       [15:0]   _zz_13826;
  wire       [15:0]   _zz_13827;
  wire       [15:0]   _zz_13828;
  wire       [15:0]   _zz_13829;
  wire       [15:0]   _zz_13830;
  wire       [15:0]   _zz_13831;
  wire       [15:0]   _zz_13832;
  wire       [15:0]   _zz_13833;
  wire       [15:0]   _zz_13834;
  wire       [15:0]   _zz_13835;
  wire       [15:0]   _zz_13836;
  wire       [15:0]   _zz_13837;
  wire       [15:0]   _zz_13838;
  wire       [15:0]   _zz_13839;
  wire       [15:0]   _zz_13840;
  wire       [15:0]   _zz_13841;
  wire       [15:0]   _zz_13842;
  wire       [15:0]   _zz_13843;
  wire       [15:0]   _zz_13844;
  wire       [15:0]   _zz_13845;
  wire       [15:0]   _zz_13846;
  wire       [15:0]   _zz_13847;
  wire       [15:0]   _zz_13848;
  wire       [15:0]   _zz_13849;
  wire       [15:0]   _zz_13850;
  wire       [15:0]   _zz_13851;
  wire       [15:0]   _zz_13852;
  wire       [15:0]   _zz_13853;
  wire       [15:0]   _zz_13854;
  wire       [15:0]   _zz_13855;
  wire       [15:0]   _zz_13856;
  wire       [15:0]   _zz_13857;
  wire       [15:0]   _zz_13858;
  wire       [15:0]   _zz_13859;
  wire       [15:0]   _zz_13860;
  wire       [15:0]   _zz_13861;
  wire       [15:0]   _zz_13862;
  wire       [15:0]   _zz_13863;
  wire       [15:0]   _zz_13864;
  wire       [15:0]   _zz_13865;
  wire       [15:0]   _zz_13866;
  wire       [15:0]   _zz_13867;
  wire       [15:0]   _zz_13868;
  wire       [15:0]   _zz_13869;
  wire       [15:0]   _zz_13870;
  wire       [15:0]   _zz_13871;
  wire       [15:0]   _zz_13872;
  wire       [15:0]   _zz_13873;
  wire       [15:0]   _zz_13874;
  wire       [15:0]   _zz_13875;
  wire       [15:0]   _zz_13876;
  wire       [15:0]   _zz_13877;
  wire       [15:0]   _zz_13878;
  wire       [15:0]   _zz_13879;
  wire       [15:0]   _zz_13880;
  wire       [15:0]   _zz_13881;
  wire       [15:0]   _zz_13882;
  wire       [15:0]   _zz_13883;
  wire       [15:0]   _zz_13884;
  wire       [15:0]   _zz_13885;
  wire       [15:0]   _zz_13886;
  wire       [15:0]   _zz_13887;
  wire       [15:0]   _zz_13888;
  wire       [15:0]   _zz_13889;
  wire       [15:0]   _zz_13890;
  wire       [15:0]   _zz_13891;
  wire       [15:0]   _zz_13892;
  wire       [15:0]   _zz_13893;
  wire       [15:0]   _zz_13894;
  wire       [15:0]   _zz_13895;
  wire       [15:0]   _zz_13896;
  wire       [15:0]   _zz_13897;
  wire       [15:0]   _zz_13898;
  wire       [15:0]   _zz_13899;
  wire       [15:0]   _zz_13900;
  wire       [15:0]   _zz_13901;
  wire       [15:0]   _zz_13902;
  wire       [15:0]   _zz_13903;
  wire       [15:0]   _zz_13904;
  wire       [15:0]   _zz_13905;
  wire       [15:0]   _zz_13906;
  wire       [15:0]   _zz_13907;
  wire       [15:0]   _zz_13908;
  wire       [15:0]   _zz_13909;
  wire       [15:0]   _zz_13910;
  wire       [15:0]   _zz_13911;
  wire       [15:0]   _zz_13912;
  wire       [15:0]   _zz_13913;
  wire       [15:0]   _zz_13914;
  wire       [15:0]   _zz_13915;
  wire       [15:0]   _zz_13916;
  wire       [15:0]   _zz_13917;
  wire       [15:0]   _zz_13918;
  wire       [15:0]   _zz_13919;
  wire       [15:0]   _zz_13920;
  wire       [15:0]   _zz_13921;
  wire       [15:0]   _zz_13922;
  wire       [15:0]   _zz_13923;
  wire       [15:0]   _zz_13924;
  wire       [15:0]   _zz_13925;
  wire       [15:0]   _zz_13926;
  wire       [15:0]   _zz_13927;
  wire       [15:0]   _zz_13928;
  wire       [15:0]   _zz_13929;
  wire       [15:0]   _zz_13930;
  wire       [15:0]   _zz_13931;
  wire       [15:0]   _zz_13932;
  wire       [15:0]   _zz_13933;
  wire       [15:0]   _zz_13934;
  wire       [15:0]   _zz_13935;
  wire       [15:0]   _zz_13936;
  wire       [15:0]   _zz_13937;
  wire       [15:0]   _zz_13938;
  wire       [15:0]   _zz_13939;
  wire       [15:0]   _zz_13940;
  wire       [15:0]   _zz_13941;
  wire       [15:0]   _zz_13942;
  wire       [15:0]   _zz_13943;
  wire       [15:0]   _zz_13944;
  wire       [15:0]   _zz_13945;
  wire       [15:0]   _zz_13946;
  wire       [15:0]   _zz_13947;
  wire       [15:0]   _zz_13948;
  wire       [15:0]   _zz_13949;
  wire       [15:0]   _zz_13950;
  wire       [15:0]   _zz_13951;
  wire       [15:0]   _zz_13952;
  wire       [15:0]   _zz_13953;
  wire       [15:0]   _zz_13954;
  wire       [15:0]   _zz_13955;
  wire       [15:0]   _zz_13956;
  wire       [15:0]   _zz_13957;
  wire       [15:0]   _zz_13958;
  wire       [15:0]   _zz_13959;
  wire       [15:0]   _zz_13960;
  wire       [15:0]   _zz_13961;
  wire       [15:0]   _zz_13962;
  wire       [15:0]   _zz_13963;
  wire       [15:0]   _zz_13964;
  wire       [15:0]   _zz_13965;
  wire       [15:0]   _zz_13966;
  wire       [15:0]   _zz_13967;
  wire       [15:0]   _zz_13968;
  wire       [15:0]   _zz_13969;
  wire       [15:0]   _zz_13970;
  wire       [15:0]   _zz_13971;
  wire       [15:0]   _zz_13972;
  wire       [15:0]   _zz_13973;
  wire       [15:0]   _zz_13974;
  wire       [15:0]   _zz_13975;
  wire       [15:0]   _zz_13976;
  wire       [15:0]   _zz_13977;
  wire       [15:0]   _zz_13978;
  wire       [15:0]   _zz_13979;
  wire       [15:0]   _zz_13980;
  wire       [15:0]   _zz_13981;
  wire       [15:0]   _zz_13982;
  wire       [15:0]   _zz_13983;
  wire       [15:0]   _zz_13984;
  wire       [15:0]   _zz_13985;
  wire       [15:0]   _zz_13986;
  wire       [15:0]   _zz_13987;
  wire       [15:0]   _zz_13988;
  wire       [15:0]   _zz_13989;
  wire       [15:0]   _zz_13990;
  wire       [15:0]   _zz_13991;
  wire       [15:0]   _zz_13992;
  wire       [15:0]   _zz_13993;
  wire       [15:0]   _zz_13994;
  wire       [15:0]   _zz_13995;
  wire       [15:0]   _zz_13996;
  wire       [15:0]   _zz_13997;
  wire       [15:0]   _zz_13998;
  wire       [15:0]   _zz_13999;
  wire       [15:0]   _zz_14000;
  wire       [15:0]   _zz_14001;
  wire       [15:0]   _zz_14002;
  wire       [15:0]   _zz_14003;
  wire       [15:0]   _zz_14004;
  wire       [15:0]   _zz_14005;
  wire       [15:0]   _zz_14006;
  wire       [15:0]   _zz_14007;
  wire       [15:0]   _zz_14008;
  wire       [15:0]   _zz_14009;
  wire       [15:0]   _zz_14010;
  wire       [15:0]   _zz_14011;
  wire       [15:0]   _zz_14012;
  wire       [15:0]   _zz_14013;
  wire       [15:0]   _zz_14014;
  wire       [15:0]   _zz_14015;
  wire       [15:0]   _zz_14016;
  wire       [15:0]   _zz_14017;
  wire       [15:0]   _zz_14018;
  wire       [15:0]   _zz_14019;
  wire       [15:0]   _zz_14020;
  wire       [15:0]   _zz_14021;
  wire       [15:0]   _zz_14022;
  wire       [15:0]   _zz_14023;
  wire       [15:0]   _zz_14024;
  wire       [15:0]   _zz_14025;
  wire       [15:0]   _zz_14026;
  wire       [15:0]   _zz_14027;
  wire       [15:0]   _zz_14028;
  wire       [15:0]   _zz_14029;
  wire       [15:0]   _zz_14030;
  wire       [15:0]   _zz_14031;
  wire       [15:0]   _zz_14032;
  wire       [15:0]   _zz_14033;
  wire       [15:0]   _zz_14034;
  wire       [15:0]   _zz_14035;
  wire       [15:0]   _zz_14036;
  wire       [15:0]   _zz_14037;
  wire       [15:0]   _zz_14038;
  wire       [15:0]   _zz_14039;
  wire       [15:0]   _zz_14040;
  wire       [15:0]   _zz_14041;
  wire       [15:0]   _zz_14042;
  wire       [15:0]   _zz_14043;
  wire       [15:0]   _zz_14044;
  wire       [15:0]   _zz_14045;
  wire       [15:0]   _zz_14046;
  wire       [15:0]   _zz_14047;
  wire       [15:0]   _zz_14048;
  wire       [15:0]   _zz_14049;
  wire       [15:0]   _zz_14050;
  wire       [15:0]   _zz_14051;
  wire       [15:0]   _zz_14052;
  wire       [15:0]   _zz_14053;
  wire       [15:0]   _zz_14054;
  wire       [15:0]   _zz_14055;
  wire       [15:0]   _zz_14056;
  wire       [15:0]   _zz_14057;
  wire       [15:0]   _zz_14058;
  wire       [15:0]   _zz_14059;
  wire       [15:0]   _zz_14060;
  wire       [15:0]   _zz_14061;
  wire       [15:0]   _zz_14062;
  wire       [15:0]   _zz_14063;
  wire       [15:0]   _zz_14064;
  wire       [15:0]   _zz_14065;
  wire       [15:0]   _zz_14066;
  wire       [15:0]   _zz_14067;
  wire       [15:0]   _zz_14068;
  wire       [15:0]   _zz_14069;
  wire       [15:0]   _zz_14070;
  wire       [15:0]   _zz_14071;
  wire       [15:0]   _zz_14072;
  wire       [15:0]   _zz_14073;
  wire       [15:0]   _zz_14074;
  wire       [15:0]   _zz_14075;
  wire       [15:0]   _zz_14076;
  wire       [15:0]   _zz_14077;
  wire       [15:0]   _zz_14078;
  wire       [15:0]   _zz_14079;
  wire       [15:0]   _zz_14080;
  wire       [15:0]   _zz_14081;
  wire       [15:0]   _zz_14082;
  wire       [15:0]   _zz_14083;
  wire       [15:0]   _zz_14084;
  wire       [15:0]   _zz_14085;
  wire       [15:0]   _zz_14086;
  wire       [15:0]   _zz_14087;
  wire       [15:0]   _zz_14088;
  wire       [15:0]   _zz_14089;
  wire       [15:0]   _zz_14090;
  wire       [15:0]   _zz_14091;
  wire       [15:0]   _zz_14092;
  wire       [15:0]   _zz_14093;
  wire       [15:0]   _zz_14094;
  wire       [15:0]   _zz_14095;
  wire       [15:0]   _zz_14096;
  wire       [15:0]   _zz_14097;
  wire       [15:0]   _zz_14098;
  wire       [15:0]   _zz_14099;
  wire       [15:0]   _zz_14100;
  wire       [15:0]   _zz_14101;
  wire       [15:0]   _zz_14102;
  wire       [15:0]   _zz_14103;
  wire       [15:0]   _zz_14104;
  wire       [15:0]   _zz_14105;
  wire       [15:0]   _zz_14106;
  wire       [15:0]   _zz_14107;
  wire       [15:0]   _zz_14108;
  wire       [15:0]   _zz_14109;
  wire       [15:0]   _zz_14110;
  wire       [15:0]   _zz_14111;
  wire       [15:0]   _zz_14112;
  wire       [15:0]   _zz_14113;
  wire       [15:0]   _zz_14114;
  wire       [15:0]   _zz_14115;
  wire       [15:0]   _zz_14116;
  wire       [15:0]   _zz_14117;
  wire       [15:0]   _zz_14118;
  wire       [15:0]   _zz_14119;
  wire       [15:0]   _zz_14120;
  wire       [15:0]   _zz_14121;
  wire       [15:0]   _zz_14122;
  wire       [15:0]   _zz_14123;
  wire       [15:0]   _zz_14124;
  wire       [15:0]   _zz_14125;
  wire       [15:0]   _zz_14126;
  wire       [15:0]   _zz_14127;
  wire       [15:0]   _zz_14128;
  wire       [15:0]   _zz_14129;
  wire       [15:0]   _zz_14130;
  wire       [15:0]   _zz_14131;
  wire       [15:0]   _zz_14132;
  wire       [15:0]   _zz_14133;
  wire       [15:0]   _zz_14134;
  wire       [15:0]   _zz_14135;
  wire       [15:0]   _zz_14136;
  wire       [15:0]   _zz_14137;
  wire       [15:0]   _zz_14138;
  wire       [15:0]   _zz_14139;
  wire       [15:0]   _zz_14140;
  wire       [15:0]   _zz_14141;
  wire       [15:0]   _zz_14142;
  wire       [15:0]   _zz_14143;
  wire       [15:0]   _zz_14144;
  wire       [15:0]   _zz_14145;
  wire       [15:0]   _zz_14146;
  wire       [15:0]   _zz_14147;
  wire       [15:0]   _zz_14148;
  wire       [15:0]   _zz_14149;
  wire       [15:0]   _zz_14150;
  wire       [15:0]   _zz_14151;
  wire       [15:0]   _zz_14152;
  wire       [15:0]   _zz_14153;
  wire       [15:0]   _zz_14154;
  wire       [15:0]   _zz_14155;
  wire       [15:0]   _zz_14156;
  wire       [15:0]   _zz_14157;
  wire       [15:0]   _zz_14158;
  wire       [15:0]   _zz_14159;
  wire       [15:0]   _zz_14160;
  wire       [15:0]   _zz_14161;
  wire       [15:0]   _zz_14162;
  wire       [15:0]   _zz_14163;
  wire       [15:0]   _zz_14164;
  wire       [15:0]   _zz_14165;
  wire       [15:0]   _zz_14166;
  wire       [15:0]   _zz_14167;
  wire       [15:0]   _zz_14168;
  wire       [15:0]   _zz_14169;
  wire       [15:0]   _zz_14170;
  wire       [15:0]   _zz_14171;
  wire       [15:0]   _zz_14172;
  wire       [15:0]   _zz_14173;
  wire       [15:0]   _zz_14174;
  wire       [15:0]   _zz_14175;
  wire       [15:0]   _zz_14176;
  wire       [15:0]   _zz_14177;
  wire       [15:0]   _zz_14178;
  wire       [15:0]   _zz_14179;
  wire       [15:0]   _zz_14180;
  wire       [15:0]   _zz_14181;
  wire       [15:0]   _zz_14182;
  wire       [15:0]   _zz_14183;
  wire       [15:0]   _zz_14184;
  wire       [15:0]   _zz_14185;
  wire       [15:0]   _zz_14186;
  wire       [15:0]   _zz_14187;
  wire       [15:0]   _zz_14188;
  wire       [15:0]   _zz_14189;
  wire       [15:0]   _zz_14190;
  wire       [15:0]   _zz_14191;
  wire       [15:0]   _zz_14192;
  wire       [15:0]   _zz_14193;
  wire       [15:0]   _zz_14194;
  wire       [15:0]   _zz_14195;
  wire       [15:0]   _zz_14196;
  wire       [15:0]   _zz_14197;
  wire       [15:0]   _zz_14198;
  wire       [15:0]   _zz_14199;
  wire       [15:0]   _zz_14200;
  wire       [15:0]   _zz_14201;
  wire       [15:0]   _zz_14202;
  wire       [15:0]   _zz_14203;
  wire       [15:0]   _zz_14204;
  wire       [15:0]   _zz_14205;
  wire       [15:0]   _zz_14206;
  wire       [15:0]   _zz_14207;
  wire       [15:0]   _zz_14208;
  wire       [15:0]   _zz_14209;
  wire       [15:0]   _zz_14210;
  wire       [15:0]   _zz_14211;
  wire       [15:0]   _zz_14212;
  wire       [15:0]   _zz_14213;
  wire       [15:0]   _zz_14214;
  wire       [15:0]   _zz_14215;
  wire       [15:0]   _zz_14216;
  wire       [15:0]   _zz_14217;
  wire       [15:0]   _zz_14218;
  wire       [15:0]   _zz_14219;
  wire       [15:0]   _zz_14220;
  wire       [15:0]   _zz_14221;
  wire       [15:0]   _zz_14222;
  wire       [15:0]   _zz_14223;
  wire       [15:0]   _zz_14224;
  wire       [15:0]   _zz_14225;
  wire       [15:0]   _zz_14226;
  wire       [15:0]   _zz_14227;
  wire       [15:0]   _zz_14228;
  wire       [15:0]   _zz_14229;
  wire       [15:0]   _zz_14230;
  wire       [15:0]   _zz_14231;
  wire       [15:0]   _zz_14232;
  wire       [15:0]   _zz_14233;
  wire       [15:0]   _zz_14234;
  wire       [15:0]   _zz_14235;
  wire       [15:0]   _zz_14236;
  wire       [15:0]   _zz_14237;
  wire       [15:0]   _zz_14238;
  wire       [15:0]   _zz_14239;
  wire       [15:0]   _zz_14240;
  wire       [15:0]   _zz_14241;
  wire       [15:0]   _zz_14242;
  wire       [15:0]   _zz_14243;
  wire       [15:0]   _zz_14244;
  wire       [15:0]   _zz_14245;
  wire       [15:0]   _zz_14246;
  wire       [15:0]   _zz_14247;
  wire       [15:0]   _zz_14248;
  wire       [15:0]   _zz_14249;
  wire       [15:0]   _zz_14250;
  wire       [15:0]   _zz_14251;
  wire       [15:0]   _zz_14252;
  wire       [15:0]   _zz_14253;
  wire       [15:0]   _zz_14254;
  wire       [15:0]   _zz_14255;
  wire       [15:0]   _zz_14256;
  wire       [15:0]   _zz_14257;
  wire       [15:0]   _zz_14258;
  wire       [15:0]   _zz_14259;
  wire       [15:0]   _zz_14260;
  wire       [15:0]   _zz_14261;
  wire       [15:0]   _zz_14262;
  wire       [15:0]   _zz_14263;
  wire       [15:0]   _zz_14264;
  wire       [15:0]   _zz_14265;
  wire       [15:0]   _zz_14266;
  wire       [15:0]   _zz_14267;
  wire       [15:0]   _zz_14268;
  wire       [15:0]   _zz_14269;
  wire       [15:0]   _zz_14270;
  wire       [15:0]   _zz_14271;
  wire       [15:0]   _zz_14272;
  wire       [15:0]   _zz_14273;
  wire       [15:0]   _zz_14274;
  wire       [15:0]   _zz_14275;
  wire       [15:0]   _zz_14276;
  wire       [15:0]   _zz_14277;
  wire       [15:0]   _zz_14278;
  wire       [15:0]   _zz_14279;
  wire       [15:0]   _zz_14280;
  wire       [15:0]   _zz_14281;
  wire       [15:0]   _zz_14282;
  wire       [15:0]   _zz_14283;
  wire       [15:0]   _zz_14284;
  wire       [15:0]   _zz_14285;
  wire       [15:0]   _zz_14286;
  wire       [15:0]   _zz_14287;
  wire       [15:0]   _zz_14288;
  wire       [15:0]   _zz_14289;
  wire       [15:0]   _zz_14290;
  wire       [15:0]   _zz_14291;
  wire       [15:0]   _zz_14292;
  wire       [15:0]   _zz_14293;
  wire       [15:0]   _zz_14294;
  wire       [15:0]   _zz_14295;
  wire       [15:0]   _zz_14296;
  wire       [15:0]   _zz_14297;
  wire       [15:0]   _zz_14298;
  wire       [15:0]   _zz_14299;
  wire       [15:0]   _zz_14300;
  wire       [15:0]   _zz_14301;
  wire       [15:0]   _zz_14302;
  wire       [15:0]   _zz_14303;
  wire       [15:0]   _zz_14304;
  wire       [15:0]   _zz_14305;
  wire       [15:0]   _zz_14306;
  wire       [15:0]   _zz_14307;
  wire       [15:0]   _zz_14308;
  wire       [15:0]   _zz_14309;
  wire       [15:0]   _zz_14310;
  wire       [15:0]   _zz_14311;
  wire       [15:0]   _zz_14312;
  wire       [15:0]   _zz_14313;
  wire       [15:0]   _zz_14314;
  wire       [15:0]   _zz_14315;
  wire       [15:0]   _zz_14316;
  wire       [15:0]   _zz_14317;
  wire       [15:0]   _zz_14318;
  wire       [15:0]   _zz_14319;
  wire       [15:0]   _zz_14320;
  wire       [15:0]   _zz_14321;
  wire       [15:0]   _zz_14322;
  wire       [15:0]   _zz_14323;
  wire       [15:0]   _zz_14324;
  wire       [15:0]   _zz_14325;
  wire       [15:0]   _zz_14326;
  wire       [15:0]   _zz_14327;
  wire       [15:0]   _zz_14328;
  wire       [15:0]   _zz_14329;
  wire       [15:0]   _zz_14330;
  wire       [15:0]   _zz_14331;
  wire       [15:0]   _zz_14332;
  wire       [15:0]   _zz_14333;
  wire       [15:0]   _zz_14334;
  wire       [15:0]   _zz_14335;
  wire       [15:0]   _zz_14336;
  wire       [15:0]   _zz_14337;
  wire       [15:0]   _zz_14338;
  wire       [15:0]   _zz_14339;
  wire       [15:0]   _zz_14340;
  wire       [15:0]   _zz_14341;
  wire       [15:0]   _zz_14342;
  wire       [15:0]   _zz_14343;
  wire       [15:0]   _zz_14344;
  wire       [15:0]   _zz_14345;
  wire       [15:0]   _zz_14346;
  wire       [15:0]   _zz_14347;
  wire       [15:0]   _zz_14348;
  wire       [15:0]   _zz_14349;
  wire       [15:0]   _zz_14350;
  wire       [15:0]   _zz_14351;
  wire       [15:0]   _zz_14352;
  wire       [15:0]   _zz_14353;
  wire       [15:0]   _zz_14354;
  wire       [15:0]   _zz_14355;
  wire       [15:0]   _zz_14356;
  wire       [15:0]   _zz_14357;
  wire       [15:0]   _zz_14358;
  wire       [15:0]   _zz_14359;
  wire       [15:0]   _zz_14360;
  wire       [15:0]   _zz_14361;
  wire       [15:0]   _zz_14362;
  wire       [15:0]   _zz_14363;
  wire       [15:0]   _zz_14364;
  wire       [15:0]   _zz_14365;
  wire       [15:0]   _zz_14366;
  wire       [15:0]   _zz_14367;
  wire       [15:0]   _zz_14368;
  wire       [15:0]   _zz_14369;
  wire       [15:0]   _zz_14370;
  wire       [15:0]   _zz_14371;
  wire       [15:0]   _zz_14372;
  wire       [15:0]   _zz_14373;
  wire       [15:0]   _zz_14374;
  wire       [15:0]   _zz_14375;
  wire       [15:0]   _zz_14376;
  wire       [15:0]   _zz_14377;
  wire       [15:0]   _zz_14378;
  wire       [15:0]   _zz_14379;
  wire       [15:0]   _zz_14380;
  wire       [15:0]   _zz_14381;
  wire       [15:0]   _zz_14382;
  wire       [15:0]   _zz_14383;
  wire       [15:0]   _zz_14384;
  wire       [15:0]   _zz_14385;
  wire       [15:0]   _zz_14386;
  wire       [15:0]   _zz_14387;
  wire       [15:0]   _zz_14388;
  wire       [15:0]   _zz_14389;
  wire       [15:0]   _zz_14390;
  wire       [15:0]   _zz_14391;
  wire       [15:0]   _zz_14392;
  wire       [15:0]   _zz_14393;
  wire       [15:0]   _zz_14394;
  wire       [15:0]   _zz_14395;
  wire       [15:0]   _zz_14396;
  wire       [15:0]   _zz_14397;
  wire       [15:0]   _zz_14398;
  wire       [15:0]   _zz_14399;
  wire       [15:0]   _zz_14400;
  wire       [15:0]   _zz_14401;
  wire       [15:0]   _zz_14402;
  wire       [15:0]   _zz_14403;
  wire       [15:0]   _zz_14404;
  wire       [15:0]   _zz_14405;
  wire       [15:0]   _zz_14406;
  wire       [15:0]   _zz_14407;
  wire       [15:0]   _zz_14408;
  wire       [15:0]   _zz_14409;
  wire       [15:0]   _zz_14410;
  wire       [15:0]   _zz_14411;
  wire       [15:0]   _zz_14412;
  wire       [15:0]   _zz_14413;
  wire       [15:0]   _zz_14414;
  wire       [15:0]   _zz_14415;
  wire       [15:0]   _zz_14416;
  wire       [15:0]   _zz_14417;
  wire       [15:0]   _zz_14418;
  wire       [15:0]   _zz_14419;
  wire       [15:0]   _zz_14420;
  wire       [15:0]   _zz_14421;
  wire       [15:0]   _zz_14422;
  wire       [15:0]   _zz_14423;
  wire       [15:0]   _zz_14424;
  wire       [15:0]   _zz_14425;
  wire       [15:0]   _zz_14426;
  wire       [15:0]   _zz_14427;
  wire       [15:0]   _zz_14428;
  wire       [15:0]   _zz_14429;
  wire       [15:0]   _zz_14430;
  wire       [15:0]   _zz_14431;
  wire       [15:0]   _zz_14432;
  wire       [15:0]   _zz_14433;
  wire       [15:0]   _zz_14434;
  wire       [15:0]   _zz_14435;
  wire       [15:0]   _zz_14436;
  wire       [15:0]   _zz_14437;
  wire       [15:0]   _zz_14438;
  wire       [15:0]   _zz_14439;
  wire       [15:0]   _zz_14440;
  wire       [15:0]   _zz_14441;
  wire       [15:0]   _zz_14442;
  wire       [15:0]   _zz_14443;
  wire       [15:0]   _zz_14444;
  wire       [15:0]   _zz_14445;
  wire       [15:0]   _zz_14446;
  wire       [15:0]   _zz_14447;
  wire       [15:0]   _zz_14448;
  wire       [15:0]   _zz_14449;
  wire       [15:0]   _zz_14450;
  wire       [15:0]   _zz_14451;
  wire       [15:0]   _zz_14452;
  wire       [15:0]   _zz_14453;
  wire       [15:0]   _zz_14454;
  wire       [15:0]   _zz_14455;
  wire       [15:0]   _zz_14456;
  wire       [15:0]   _zz_14457;
  wire       [15:0]   _zz_14458;
  wire       [15:0]   _zz_14459;
  wire       [15:0]   _zz_14460;
  wire       [15:0]   _zz_14461;
  wire       [15:0]   _zz_14462;
  wire       [15:0]   _zz_14463;
  wire       [15:0]   _zz_14464;
  wire       [15:0]   _zz_14465;
  wire       [15:0]   _zz_14466;
  wire       [15:0]   _zz_14467;
  wire       [15:0]   _zz_14468;
  wire       [15:0]   _zz_14469;
  wire       [15:0]   _zz_14470;
  wire       [15:0]   _zz_14471;
  wire       [15:0]   _zz_14472;
  wire       [15:0]   _zz_14473;
  wire       [15:0]   _zz_14474;
  wire       [15:0]   _zz_14475;
  wire       [15:0]   _zz_14476;
  wire       [15:0]   _zz_14477;
  wire       [15:0]   _zz_14478;
  wire       [15:0]   _zz_14479;
  wire       [15:0]   _zz_14480;
  wire       [15:0]   _zz_14481;
  wire       [15:0]   _zz_14482;
  wire       [15:0]   _zz_14483;
  wire       [15:0]   _zz_14484;
  wire       [15:0]   _zz_14485;
  wire       [15:0]   _zz_14486;
  wire       [15:0]   _zz_14487;
  wire       [15:0]   _zz_14488;
  wire       [15:0]   _zz_14489;
  wire       [15:0]   _zz_14490;
  wire       [15:0]   _zz_14491;
  wire       [15:0]   _zz_14492;
  wire       [15:0]   _zz_14493;
  wire       [15:0]   _zz_14494;
  wire       [15:0]   _zz_14495;
  wire       [15:0]   _zz_14496;
  wire       [15:0]   _zz_14497;
  wire       [15:0]   _zz_14498;
  wire       [15:0]   _zz_14499;
  wire       [15:0]   _zz_14500;
  wire       [15:0]   _zz_14501;
  wire       [15:0]   _zz_14502;
  wire       [15:0]   _zz_14503;
  wire       [15:0]   _zz_14504;
  wire       [15:0]   _zz_14505;
  wire       [15:0]   _zz_14506;
  wire       [15:0]   _zz_14507;
  wire       [15:0]   _zz_14508;
  wire       [15:0]   _zz_14509;
  wire       [15:0]   _zz_14510;
  wire       [15:0]   _zz_14511;
  wire       [15:0]   _zz_14512;
  wire       [15:0]   _zz_14513;
  wire       [15:0]   _zz_14514;
  wire       [15:0]   _zz_14515;
  wire       [15:0]   _zz_14516;
  wire       [15:0]   _zz_14517;
  wire       [15:0]   _zz_14518;
  wire       [15:0]   _zz_14519;
  wire       [15:0]   _zz_14520;
  wire       [15:0]   _zz_14521;
  wire       [15:0]   _zz_14522;
  wire       [15:0]   _zz_14523;
  wire       [15:0]   _zz_14524;
  wire       [15:0]   _zz_14525;
  wire       [15:0]   _zz_14526;
  wire       [15:0]   _zz_14527;
  wire       [15:0]   _zz_14528;
  wire       [15:0]   _zz_14529;
  wire       [15:0]   _zz_14530;
  wire       [15:0]   _zz_14531;
  wire       [15:0]   _zz_14532;
  wire       [15:0]   _zz_14533;
  wire       [15:0]   _zz_14534;
  wire       [15:0]   _zz_14535;
  wire       [15:0]   _zz_14536;
  wire       [15:0]   _zz_14537;
  wire       [15:0]   _zz_14538;
  wire       [15:0]   _zz_14539;
  wire       [15:0]   _zz_14540;
  wire       [15:0]   _zz_14541;
  wire       [15:0]   _zz_14542;
  wire       [15:0]   _zz_14543;
  wire       [15:0]   _zz_14544;
  wire       [15:0]   _zz_14545;
  wire       [15:0]   _zz_14546;
  wire       [15:0]   _zz_14547;
  wire       [15:0]   _zz_14548;
  wire       [15:0]   _zz_14549;
  wire       [15:0]   _zz_14550;
  wire       [15:0]   _zz_14551;
  wire       [15:0]   _zz_14552;
  wire       [15:0]   _zz_14553;
  wire       [15:0]   _zz_14554;
  wire       [15:0]   _zz_14555;
  wire       [15:0]   _zz_14556;
  wire       [15:0]   _zz_14557;
  wire       [15:0]   _zz_14558;
  wire       [15:0]   _zz_14559;
  wire       [15:0]   _zz_14560;
  wire       [15:0]   _zz_14561;
  wire       [15:0]   _zz_14562;
  wire       [15:0]   _zz_14563;
  wire       [15:0]   _zz_14564;
  wire       [15:0]   _zz_14565;
  wire       [15:0]   _zz_14566;
  wire       [15:0]   _zz_14567;
  wire       [15:0]   _zz_14568;
  wire       [15:0]   _zz_14569;
  wire       [15:0]   _zz_14570;
  wire       [15:0]   _zz_14571;
  wire       [15:0]   _zz_14572;
  wire       [15:0]   _zz_14573;
  wire       [15:0]   _zz_14574;
  wire       [15:0]   _zz_14575;
  wire       [15:0]   _zz_14576;
  wire       [15:0]   _zz_14577;
  wire       [15:0]   _zz_14578;
  wire       [15:0]   _zz_14579;
  wire       [15:0]   _zz_14580;
  wire       [15:0]   _zz_14581;
  wire       [15:0]   _zz_14582;
  wire       [15:0]   _zz_14583;
  wire       [15:0]   _zz_14584;
  wire       [15:0]   _zz_14585;
  wire       [15:0]   _zz_14586;
  wire       [15:0]   _zz_14587;
  wire       [15:0]   _zz_14588;
  wire       [15:0]   _zz_14589;
  wire       [15:0]   _zz_14590;
  wire       [15:0]   _zz_14591;
  wire       [15:0]   _zz_14592;
  wire       [15:0]   _zz_14593;
  wire       [15:0]   _zz_14594;
  wire       [15:0]   _zz_14595;
  wire       [15:0]   _zz_14596;
  wire       [15:0]   _zz_14597;
  wire       [15:0]   _zz_14598;
  wire       [15:0]   _zz_14599;
  wire       [15:0]   _zz_14600;
  wire       [15:0]   _zz_14601;
  wire       [15:0]   _zz_14602;
  wire       [15:0]   _zz_14603;
  wire       [15:0]   _zz_14604;
  wire       [15:0]   _zz_14605;
  wire       [15:0]   _zz_14606;
  wire       [15:0]   _zz_14607;
  wire       [15:0]   _zz_14608;
  wire       [15:0]   _zz_14609;
  wire       [15:0]   _zz_14610;
  wire       [15:0]   _zz_14611;
  wire       [15:0]   _zz_14612;
  wire       [15:0]   _zz_14613;
  wire       [15:0]   _zz_14614;
  wire       [15:0]   _zz_14615;
  wire       [15:0]   _zz_14616;
  wire       [15:0]   _zz_14617;
  wire       [15:0]   _zz_14618;
  wire       [15:0]   _zz_14619;
  wire       [15:0]   _zz_14620;
  wire       [15:0]   _zz_14621;
  wire       [15:0]   _zz_14622;
  wire       [15:0]   _zz_14623;
  wire       [15:0]   _zz_14624;
  wire       [15:0]   _zz_14625;
  wire       [15:0]   _zz_14626;
  wire       [15:0]   _zz_14627;
  wire       [15:0]   _zz_14628;
  wire       [15:0]   _zz_14629;
  wire       [15:0]   _zz_14630;
  wire       [15:0]   _zz_14631;
  wire       [15:0]   _zz_14632;
  wire       [15:0]   _zz_14633;
  wire       [15:0]   _zz_14634;
  wire       [15:0]   _zz_14635;
  wire       [15:0]   _zz_14636;
  wire       [15:0]   _zz_14637;
  wire       [15:0]   _zz_14638;
  wire       [15:0]   _zz_14639;
  wire       [15:0]   _zz_14640;
  wire       [15:0]   _zz_14641;
  wire       [15:0]   _zz_14642;
  wire       [15:0]   _zz_14643;
  wire       [15:0]   _zz_14644;
  wire       [15:0]   _zz_14645;
  wire       [15:0]   _zz_14646;
  wire       [15:0]   _zz_14647;
  wire       [15:0]   _zz_14648;
  wire       [15:0]   _zz_14649;
  wire       [15:0]   _zz_14650;
  wire       [15:0]   _zz_14651;
  wire       [15:0]   _zz_14652;
  wire       [15:0]   _zz_14653;
  wire       [15:0]   _zz_14654;
  wire       [15:0]   _zz_14655;
  wire       [15:0]   _zz_14656;
  wire       [15:0]   _zz_14657;
  wire       [15:0]   _zz_14658;
  wire       [15:0]   _zz_14659;
  wire       [15:0]   _zz_14660;
  wire       [15:0]   _zz_14661;
  wire       [15:0]   _zz_14662;
  wire       [15:0]   _zz_14663;
  wire       [15:0]   _zz_14664;
  wire       [15:0]   _zz_14665;
  wire       [15:0]   _zz_14666;
  wire       [15:0]   _zz_14667;
  wire       [15:0]   _zz_14668;
  wire       [15:0]   _zz_14669;
  wire       [15:0]   _zz_14670;
  wire       [15:0]   _zz_14671;
  wire       [15:0]   _zz_14672;
  wire       [15:0]   _zz_14673;
  wire       [15:0]   _zz_14674;
  wire       [15:0]   _zz_14675;
  wire       [15:0]   _zz_14676;
  wire       [15:0]   _zz_14677;
  wire       [15:0]   _zz_14678;
  wire       [15:0]   _zz_14679;
  wire       [15:0]   _zz_14680;
  wire       [15:0]   _zz_14681;
  wire       [15:0]   _zz_14682;
  wire       [15:0]   _zz_14683;
  wire       [15:0]   _zz_14684;
  wire       [15:0]   _zz_14685;
  wire       [15:0]   _zz_14686;
  wire       [15:0]   _zz_14687;
  wire       [15:0]   _zz_14688;
  wire       [15:0]   _zz_14689;
  wire       [15:0]   _zz_14690;
  wire       [15:0]   _zz_14691;
  wire       [15:0]   _zz_14692;
  wire       [15:0]   _zz_14693;
  wire       [15:0]   _zz_14694;
  wire       [15:0]   _zz_14695;
  wire       [15:0]   _zz_14696;
  wire       [15:0]   _zz_14697;
  wire       [15:0]   _zz_14698;
  wire       [15:0]   _zz_14699;
  wire       [15:0]   _zz_14700;
  wire       [15:0]   _zz_14701;
  wire       [15:0]   _zz_14702;
  wire       [15:0]   _zz_14703;
  wire       [15:0]   _zz_14704;
  wire       [15:0]   _zz_14705;
  wire       [15:0]   _zz_14706;
  wire       [15:0]   _zz_14707;
  wire       [15:0]   _zz_14708;
  wire       [15:0]   _zz_14709;
  wire       [15:0]   _zz_14710;
  wire       [15:0]   _zz_14711;
  wire       [15:0]   _zz_14712;
  wire       [15:0]   _zz_14713;
  wire       [15:0]   _zz_14714;
  wire       [15:0]   _zz_14715;
  wire       [15:0]   _zz_14716;
  wire       [15:0]   _zz_14717;
  wire       [15:0]   _zz_14718;
  wire       [15:0]   _zz_14719;
  wire       [15:0]   _zz_14720;
  wire       [15:0]   _zz_14721;
  wire       [15:0]   _zz_14722;
  wire       [15:0]   _zz_14723;
  wire       [15:0]   _zz_14724;
  wire       [15:0]   _zz_14725;
  wire       [15:0]   _zz_14726;
  wire       [15:0]   _zz_14727;
  wire       [15:0]   _zz_14728;
  wire       [15:0]   _zz_14729;
  wire       [15:0]   _zz_14730;
  wire       [15:0]   _zz_14731;
  wire       [15:0]   _zz_14732;
  wire       [15:0]   _zz_14733;
  wire       [15:0]   _zz_14734;
  wire       [15:0]   _zz_14735;
  wire       [15:0]   _zz_14736;
  wire       [15:0]   _zz_14737;
  wire       [15:0]   _zz_14738;
  wire       [15:0]   _zz_14739;
  wire       [15:0]   _zz_14740;
  wire       [15:0]   _zz_14741;
  wire       [15:0]   _zz_14742;
  wire       [15:0]   _zz_14743;
  wire       [15:0]   _zz_14744;
  wire       [15:0]   _zz_14745;
  wire       [15:0]   _zz_14746;
  wire       [15:0]   _zz_14747;
  wire       [15:0]   _zz_14748;
  wire       [15:0]   _zz_14749;
  wire       [15:0]   _zz_14750;
  wire       [15:0]   _zz_14751;
  wire       [15:0]   _zz_14752;
  wire       [15:0]   _zz_14753;
  wire       [15:0]   _zz_14754;
  wire       [15:0]   _zz_14755;
  wire       [15:0]   _zz_14756;
  wire       [15:0]   _zz_14757;
  wire       [15:0]   _zz_14758;
  wire       [15:0]   _zz_14759;
  wire       [15:0]   _zz_14760;
  wire       [15:0]   _zz_14761;
  wire       [15:0]   _zz_14762;
  wire       [15:0]   _zz_14763;
  wire       [15:0]   _zz_14764;
  wire       [15:0]   _zz_14765;
  wire       [15:0]   _zz_14766;
  wire       [15:0]   _zz_14767;
  wire       [15:0]   _zz_14768;
  wire       [15:0]   _zz_14769;
  wire       [15:0]   _zz_14770;
  wire       [15:0]   _zz_14771;
  wire       [15:0]   _zz_14772;
  wire       [15:0]   _zz_14773;
  wire       [15:0]   _zz_14774;
  wire       [15:0]   _zz_14775;
  wire       [15:0]   _zz_14776;
  wire       [15:0]   _zz_14777;
  wire       [15:0]   _zz_14778;
  wire       [15:0]   _zz_14779;
  wire       [15:0]   _zz_14780;
  wire       [15:0]   _zz_14781;
  wire       [15:0]   _zz_14782;
  wire       [15:0]   _zz_14783;
  wire       [15:0]   _zz_14784;
  wire       [15:0]   _zz_14785;
  wire       [15:0]   _zz_14786;
  wire       [15:0]   _zz_14787;
  wire       [15:0]   _zz_14788;
  wire       [15:0]   _zz_14789;
  wire       [15:0]   _zz_14790;
  wire       [15:0]   _zz_14791;
  wire       [15:0]   _zz_14792;
  wire       [15:0]   _zz_14793;
  wire       [15:0]   _zz_14794;
  wire       [15:0]   _zz_14795;
  wire       [15:0]   _zz_14796;
  wire       [15:0]   _zz_14797;
  wire       [15:0]   _zz_14798;
  wire       [15:0]   _zz_14799;
  wire       [15:0]   _zz_14800;
  wire       [15:0]   _zz_14801;
  wire       [15:0]   _zz_14802;
  wire       [15:0]   _zz_14803;
  wire       [15:0]   _zz_14804;
  wire       [15:0]   _zz_14805;
  wire       [15:0]   _zz_14806;
  wire       [15:0]   _zz_14807;
  wire       [15:0]   _zz_14808;
  wire       [15:0]   _zz_14809;
  wire       [15:0]   _zz_14810;
  wire       [15:0]   _zz_14811;
  wire       [15:0]   _zz_14812;
  wire       [15:0]   _zz_14813;
  wire       [15:0]   _zz_14814;
  wire       [15:0]   _zz_14815;
  wire       [15:0]   _zz_14816;
  wire       [15:0]   _zz_14817;
  wire       [15:0]   _zz_14818;
  wire       [15:0]   _zz_14819;
  wire       [15:0]   _zz_14820;
  wire       [15:0]   _zz_14821;
  wire       [15:0]   _zz_14822;
  wire       [15:0]   _zz_14823;
  wire       [15:0]   _zz_14824;
  wire       [15:0]   _zz_14825;
  wire       [15:0]   _zz_14826;
  wire       [15:0]   _zz_14827;
  wire       [15:0]   _zz_14828;
  wire       [15:0]   _zz_14829;
  wire       [15:0]   _zz_14830;
  wire       [15:0]   _zz_14831;
  wire       [15:0]   _zz_14832;
  wire       [15:0]   _zz_14833;
  wire       [15:0]   _zz_14834;
  wire       [15:0]   _zz_14835;
  wire       [15:0]   _zz_14836;
  wire       [15:0]   _zz_14837;
  wire       [15:0]   _zz_14838;
  wire       [15:0]   _zz_14839;
  wire       [15:0]   _zz_14840;
  wire       [15:0]   _zz_14841;
  wire       [15:0]   _zz_14842;
  wire       [15:0]   _zz_14843;
  wire       [15:0]   _zz_14844;
  wire       [15:0]   _zz_14845;
  wire       [15:0]   _zz_14846;
  wire       [15:0]   _zz_14847;
  wire       [15:0]   _zz_14848;
  wire       [15:0]   _zz_14849;
  wire       [15:0]   _zz_14850;
  wire       [15:0]   _zz_14851;
  wire       [15:0]   _zz_14852;
  wire       [15:0]   _zz_14853;
  wire       [15:0]   _zz_14854;
  wire       [15:0]   _zz_14855;
  wire       [15:0]   _zz_14856;
  wire       [15:0]   _zz_14857;
  wire       [15:0]   _zz_14858;
  wire       [15:0]   _zz_14859;
  wire       [15:0]   _zz_14860;
  wire       [15:0]   _zz_14861;
  wire       [15:0]   _zz_14862;
  wire       [15:0]   _zz_14863;
  wire       [15:0]   _zz_14864;
  wire       [15:0]   _zz_14865;
  wire       [15:0]   _zz_14866;
  wire       [15:0]   _zz_14867;
  wire       [15:0]   _zz_14868;
  wire       [15:0]   _zz_14869;
  wire       [15:0]   _zz_14870;
  wire       [15:0]   _zz_14871;
  wire       [15:0]   _zz_14872;
  wire       [15:0]   _zz_14873;
  wire       [15:0]   _zz_14874;
  wire       [15:0]   _zz_14875;
  wire       [15:0]   _zz_14876;
  wire       [15:0]   _zz_14877;
  wire       [15:0]   _zz_14878;
  wire       [15:0]   _zz_14879;
  wire       [15:0]   _zz_14880;
  wire       [15:0]   _zz_14881;
  wire       [15:0]   _zz_14882;
  wire       [15:0]   _zz_14883;
  wire       [15:0]   _zz_14884;
  wire       [15:0]   _zz_14885;
  wire       [15:0]   _zz_14886;
  wire       [15:0]   _zz_14887;
  wire       [15:0]   _zz_14888;
  wire       [15:0]   _zz_14889;
  wire       [15:0]   _zz_14890;
  wire       [15:0]   _zz_14891;
  wire       [15:0]   _zz_14892;
  wire       [15:0]   _zz_14893;
  wire       [15:0]   _zz_14894;
  wire       [15:0]   _zz_14895;
  wire       [15:0]   _zz_14896;
  wire       [15:0]   _zz_14897;
  wire       [15:0]   _zz_14898;
  wire       [15:0]   _zz_14899;
  wire       [15:0]   _zz_14900;
  wire       [15:0]   _zz_14901;
  wire       [15:0]   _zz_14902;
  wire       [15:0]   _zz_14903;
  wire       [15:0]   _zz_14904;
  wire       [15:0]   _zz_14905;
  wire       [15:0]   _zz_14906;
  wire       [15:0]   _zz_14907;
  wire       [15:0]   _zz_14908;
  wire       [15:0]   _zz_14909;
  wire       [15:0]   _zz_14910;
  wire       [15:0]   _zz_14911;
  wire       [15:0]   _zz_14912;
  wire       [15:0]   _zz_14913;
  wire       [15:0]   _zz_14914;
  wire       [15:0]   _zz_14915;
  wire       [15:0]   _zz_14916;
  wire       [15:0]   _zz_14917;
  wire       [15:0]   _zz_14918;
  wire       [15:0]   _zz_14919;
  wire       [15:0]   _zz_14920;
  wire       [15:0]   _zz_14921;
  wire       [15:0]   _zz_14922;
  wire       [15:0]   _zz_14923;
  wire       [15:0]   _zz_14924;
  wire       [15:0]   _zz_14925;
  wire       [15:0]   _zz_14926;
  wire       [15:0]   _zz_14927;
  wire       [15:0]   _zz_14928;
  wire       [15:0]   _zz_14929;
  wire       [15:0]   _zz_14930;
  wire       [15:0]   _zz_14931;
  wire       [15:0]   _zz_14932;
  wire       [15:0]   _zz_14933;
  wire       [15:0]   _zz_14934;
  wire       [15:0]   _zz_14935;
  wire       [15:0]   _zz_14936;
  wire       [15:0]   _zz_14937;
  wire       [15:0]   _zz_14938;
  wire       [15:0]   _zz_14939;
  wire       [15:0]   _zz_14940;
  wire       [15:0]   _zz_14941;
  wire       [15:0]   _zz_14942;
  wire       [15:0]   _zz_14943;
  wire       [15:0]   _zz_14944;
  wire       [15:0]   _zz_14945;
  wire       [15:0]   _zz_14946;
  wire       [15:0]   _zz_14947;
  wire       [15:0]   _zz_14948;
  wire       [15:0]   _zz_14949;
  wire       [15:0]   _zz_14950;
  wire       [15:0]   _zz_14951;
  wire       [15:0]   _zz_14952;
  wire       [15:0]   _zz_14953;
  wire       [15:0]   _zz_14954;
  wire       [15:0]   _zz_14955;
  wire       [15:0]   _zz_14956;
  wire       [15:0]   _zz_14957;
  wire       [15:0]   _zz_14958;
  wire       [15:0]   _zz_14959;
  wire       [15:0]   _zz_14960;
  wire       [15:0]   _zz_14961;
  wire       [15:0]   _zz_14962;
  wire       [15:0]   _zz_14963;
  wire       [15:0]   _zz_14964;
  wire       [15:0]   _zz_14965;
  wire       [15:0]   _zz_14966;
  wire       [15:0]   _zz_14967;
  wire       [15:0]   _zz_14968;
  wire       [15:0]   _zz_14969;
  wire       [15:0]   _zz_14970;
  wire       [15:0]   _zz_14971;
  wire       [15:0]   _zz_14972;
  wire       [15:0]   _zz_14973;
  wire       [15:0]   _zz_14974;
  wire       [15:0]   _zz_14975;
  wire       [15:0]   _zz_14976;
  wire       [15:0]   _zz_14977;
  wire       [15:0]   _zz_14978;
  wire       [15:0]   _zz_14979;
  wire       [15:0]   _zz_14980;
  wire       [15:0]   _zz_14981;
  wire       [15:0]   _zz_14982;
  wire       [15:0]   _zz_14983;
  wire       [15:0]   _zz_14984;
  wire       [15:0]   _zz_14985;
  wire       [15:0]   _zz_14986;
  wire       [15:0]   _zz_14987;
  wire       [15:0]   _zz_14988;
  wire       [15:0]   _zz_14989;
  wire       [15:0]   _zz_14990;
  wire       [15:0]   _zz_14991;
  wire       [15:0]   _zz_14992;
  wire       [15:0]   _zz_14993;
  wire       [15:0]   _zz_14994;
  wire       [15:0]   _zz_14995;
  wire       [15:0]   _zz_14996;
  wire       [15:0]   _zz_14997;
  wire       [15:0]   _zz_14998;
  wire       [15:0]   _zz_14999;
  wire       [15:0]   _zz_15000;
  wire       [15:0]   _zz_15001;
  wire       [15:0]   _zz_15002;
  wire       [15:0]   _zz_15003;
  wire       [15:0]   _zz_15004;
  wire       [15:0]   _zz_15005;
  wire       [15:0]   _zz_15006;
  wire       [15:0]   _zz_15007;
  wire       [15:0]   _zz_15008;
  wire       [15:0]   _zz_15009;
  wire       [15:0]   _zz_15010;
  wire       [15:0]   _zz_15011;
  wire       [15:0]   _zz_15012;
  wire       [15:0]   _zz_15013;
  wire       [15:0]   _zz_15014;
  wire       [15:0]   _zz_15015;
  wire       [15:0]   _zz_15016;
  wire       [15:0]   _zz_15017;
  wire       [15:0]   _zz_15018;
  wire       [15:0]   _zz_15019;
  wire       [15:0]   _zz_15020;
  wire       [15:0]   _zz_15021;
  wire       [15:0]   _zz_15022;
  wire       [15:0]   _zz_15023;
  wire       [15:0]   _zz_15024;
  wire       [15:0]   _zz_15025;
  wire       [15:0]   _zz_15026;
  wire       [15:0]   _zz_15027;
  wire       [15:0]   _zz_15028;
  wire       [15:0]   _zz_15029;
  wire       [15:0]   _zz_15030;
  wire       [15:0]   _zz_15031;
  wire       [15:0]   _zz_15032;
  wire       [15:0]   _zz_15033;
  wire       [15:0]   _zz_15034;
  wire       [15:0]   _zz_15035;
  wire       [15:0]   _zz_15036;
  wire       [15:0]   _zz_15037;
  wire       [15:0]   _zz_15038;
  wire       [15:0]   _zz_15039;
  wire       [15:0]   _zz_15040;
  wire       [15:0]   _zz_15041;
  wire       [15:0]   _zz_15042;
  wire       [15:0]   _zz_15043;
  wire       [15:0]   _zz_15044;
  wire       [15:0]   _zz_15045;
  wire       [15:0]   _zz_15046;
  wire       [15:0]   _zz_15047;
  wire       [15:0]   _zz_15048;
  wire       [15:0]   _zz_15049;
  wire       [15:0]   _zz_15050;
  wire       [15:0]   _zz_15051;
  wire       [15:0]   _zz_15052;
  wire       [15:0]   _zz_15053;
  wire       [15:0]   _zz_15054;
  wire       [15:0]   _zz_15055;
  wire       [15:0]   _zz_15056;
  wire       [15:0]   _zz_15057;
  wire       [15:0]   _zz_15058;
  wire       [15:0]   _zz_15059;
  wire       [15:0]   _zz_15060;
  wire       [15:0]   _zz_15061;
  wire       [15:0]   _zz_15062;
  wire       [15:0]   _zz_15063;
  wire       [15:0]   _zz_15064;
  wire       [15:0]   _zz_15065;
  wire       [15:0]   _zz_15066;
  wire       [15:0]   _zz_15067;
  wire       [15:0]   _zz_15068;
  wire       [15:0]   _zz_15069;
  wire       [15:0]   _zz_15070;
  wire       [15:0]   _zz_15071;
  wire       [15:0]   _zz_15072;
  wire       [15:0]   _zz_15073;
  wire       [15:0]   _zz_15074;
  wire       [15:0]   _zz_15075;
  wire       [15:0]   _zz_15076;
  wire       [15:0]   _zz_15077;
  wire       [15:0]   _zz_15078;
  wire       [15:0]   _zz_15079;
  wire       [15:0]   _zz_15080;
  wire       [15:0]   _zz_15081;
  wire       [15:0]   _zz_15082;
  wire       [15:0]   _zz_15083;
  wire       [15:0]   _zz_15084;
  wire       [15:0]   _zz_15085;
  wire       [15:0]   _zz_15086;
  wire       [15:0]   _zz_15087;
  wire       [15:0]   _zz_15088;
  wire       [15:0]   _zz_15089;
  wire       [15:0]   _zz_15090;
  wire       [15:0]   _zz_15091;
  wire       [15:0]   _zz_15092;
  wire       [15:0]   _zz_15093;
  wire       [15:0]   _zz_15094;
  wire       [15:0]   _zz_15095;
  wire       [15:0]   _zz_15096;
  wire       [15:0]   _zz_15097;
  wire       [15:0]   _zz_15098;
  wire       [15:0]   _zz_15099;
  wire       [15:0]   _zz_15100;
  wire       [15:0]   _zz_15101;
  wire       [15:0]   _zz_15102;
  wire       [15:0]   _zz_15103;
  wire       [15:0]   _zz_15104;
  wire       [15:0]   _zz_15105;
  wire       [15:0]   _zz_15106;
  wire       [15:0]   _zz_15107;
  wire       [15:0]   _zz_15108;
  wire       [15:0]   _zz_15109;
  wire       [15:0]   _zz_15110;
  wire       [15:0]   _zz_15111;
  wire       [15:0]   _zz_15112;
  wire       [15:0]   _zz_15113;
  wire       [15:0]   _zz_15114;
  wire       [15:0]   _zz_15115;
  wire       [15:0]   _zz_15116;
  wire       [15:0]   _zz_15117;
  wire       [15:0]   _zz_15118;
  wire       [15:0]   _zz_15119;
  wire       [15:0]   _zz_15120;
  wire       [15:0]   _zz_15121;
  wire       [15:0]   _zz_15122;
  wire       [15:0]   _zz_15123;
  wire       [15:0]   _zz_15124;
  wire       [15:0]   _zz_15125;
  wire       [15:0]   _zz_15126;
  wire       [15:0]   _zz_15127;
  wire       [15:0]   _zz_15128;
  wire       [15:0]   _zz_15129;
  wire       [15:0]   _zz_15130;
  wire       [15:0]   _zz_15131;
  wire       [15:0]   _zz_15132;
  wire       [15:0]   _zz_15133;
  wire       [15:0]   _zz_15134;
  wire       [15:0]   _zz_15135;
  wire       [15:0]   _zz_15136;
  wire       [15:0]   _zz_15137;
  wire       [15:0]   _zz_15138;
  wire       [15:0]   _zz_15139;
  wire       [15:0]   _zz_15140;
  wire       [15:0]   _zz_15141;
  wire       [15:0]   _zz_15142;
  wire       [15:0]   _zz_15143;
  wire       [15:0]   _zz_15144;
  wire       [15:0]   _zz_15145;
  wire       [15:0]   _zz_15146;
  wire       [15:0]   _zz_15147;
  wire       [15:0]   _zz_15148;
  wire       [15:0]   _zz_15149;
  wire       [15:0]   _zz_15150;
  wire       [15:0]   _zz_15151;
  wire       [15:0]   _zz_15152;
  wire       [15:0]   _zz_15153;
  wire       [15:0]   _zz_15154;
  wire       [15:0]   _zz_15155;
  wire       [15:0]   _zz_15156;
  wire       [15:0]   _zz_15157;
  wire       [15:0]   _zz_15158;
  wire       [15:0]   _zz_15159;
  wire       [15:0]   _zz_15160;
  wire       [15:0]   _zz_15161;
  wire       [15:0]   _zz_15162;
  wire       [15:0]   _zz_15163;
  wire       [15:0]   _zz_15164;
  wire       [15:0]   _zz_15165;
  wire       [15:0]   _zz_15166;
  wire       [15:0]   _zz_15167;
  wire       [15:0]   _zz_15168;
  wire       [15:0]   _zz_15169;
  wire       [15:0]   _zz_15170;
  wire       [15:0]   _zz_15171;
  wire       [15:0]   _zz_15172;
  wire       [15:0]   _zz_15173;
  wire       [15:0]   _zz_15174;
  wire       [15:0]   _zz_15175;
  wire       [15:0]   _zz_15176;
  wire       [15:0]   _zz_15177;
  wire       [15:0]   _zz_15178;
  wire       [15:0]   _zz_15179;
  wire       [15:0]   _zz_15180;
  wire       [15:0]   _zz_15181;
  wire       [15:0]   _zz_15182;
  wire       [15:0]   _zz_15183;
  wire       [15:0]   _zz_15184;
  wire       [15:0]   _zz_15185;
  wire       [15:0]   _zz_15186;
  wire       [15:0]   _zz_15187;
  wire       [15:0]   _zz_15188;
  wire       [15:0]   _zz_15189;
  wire       [15:0]   _zz_15190;
  wire       [15:0]   _zz_15191;
  wire       [15:0]   _zz_15192;
  wire       [15:0]   _zz_15193;
  wire       [15:0]   _zz_15194;
  wire       [15:0]   _zz_15195;
  wire       [15:0]   _zz_15196;
  wire       [15:0]   _zz_15197;
  wire       [15:0]   _zz_15198;
  wire       [15:0]   _zz_15199;
  wire       [15:0]   _zz_15200;
  wire       [15:0]   _zz_15201;
  wire       [15:0]   _zz_15202;
  wire       [15:0]   _zz_15203;
  wire       [15:0]   _zz_15204;
  wire       [15:0]   _zz_15205;
  wire       [15:0]   _zz_15206;
  wire       [15:0]   _zz_15207;
  wire       [15:0]   _zz_15208;
  wire       [15:0]   _zz_15209;
  wire       [15:0]   _zz_15210;
  wire       [15:0]   _zz_15211;
  wire       [15:0]   _zz_15212;
  wire       [15:0]   _zz_15213;
  wire       [15:0]   _zz_15214;
  wire       [15:0]   _zz_15215;
  wire       [15:0]   _zz_15216;
  wire       [15:0]   _zz_15217;
  wire       [15:0]   _zz_15218;
  wire       [15:0]   _zz_15219;
  wire       [15:0]   _zz_15220;
  wire       [15:0]   _zz_15221;
  wire       [15:0]   _zz_15222;
  wire       [15:0]   _zz_15223;
  wire       [15:0]   _zz_15224;
  wire       [15:0]   _zz_15225;
  wire       [15:0]   _zz_15226;
  wire       [15:0]   _zz_15227;
  wire       [15:0]   _zz_15228;
  wire       [15:0]   _zz_15229;
  wire       [15:0]   _zz_15230;
  wire       [15:0]   _zz_15231;
  wire       [15:0]   _zz_15232;
  wire       [15:0]   _zz_15233;
  wire       [15:0]   _zz_15234;
  wire       [15:0]   _zz_15235;
  wire       [15:0]   _zz_15236;
  wire       [15:0]   _zz_15237;
  wire       [15:0]   _zz_15238;
  wire       [15:0]   _zz_15239;
  wire       [15:0]   _zz_15240;
  wire       [15:0]   _zz_15241;
  wire       [15:0]   _zz_15242;
  wire       [15:0]   _zz_15243;
  wire       [15:0]   _zz_15244;
  wire       [15:0]   _zz_15245;
  wire       [15:0]   _zz_15246;
  wire       [15:0]   _zz_15247;
  wire       [15:0]   _zz_15248;
  wire       [15:0]   _zz_15249;
  wire       [15:0]   _zz_15250;
  wire       [15:0]   _zz_15251;
  wire       [15:0]   _zz_15252;
  wire       [15:0]   _zz_15253;
  wire       [15:0]   _zz_15254;
  wire       [15:0]   _zz_15255;
  wire       [15:0]   _zz_15256;
  wire       [15:0]   _zz_15257;
  wire       [15:0]   _zz_15258;
  wire       [15:0]   _zz_15259;
  wire       [15:0]   _zz_15260;
  wire       [15:0]   _zz_15261;
  wire       [15:0]   _zz_15262;
  wire       [15:0]   _zz_15263;
  wire       [15:0]   _zz_15264;
  wire       [15:0]   _zz_15265;
  wire       [15:0]   _zz_15266;
  wire       [15:0]   _zz_15267;
  wire       [15:0]   _zz_15268;
  wire       [15:0]   _zz_15269;
  wire       [15:0]   _zz_15270;
  wire       [15:0]   _zz_15271;
  wire       [15:0]   _zz_15272;
  wire       [15:0]   _zz_15273;
  wire       [15:0]   _zz_15274;
  wire       [15:0]   _zz_15275;
  wire       [15:0]   _zz_15276;
  wire       [15:0]   _zz_15277;
  wire       [15:0]   _zz_15278;
  wire       [15:0]   _zz_15279;
  wire       [15:0]   _zz_15280;
  wire       [15:0]   _zz_15281;
  wire       [15:0]   _zz_15282;
  wire       [15:0]   _zz_15283;
  wire       [15:0]   _zz_15284;
  wire       [15:0]   _zz_15285;
  wire       [15:0]   _zz_15286;
  wire       [15:0]   _zz_15287;
  wire       [15:0]   _zz_15288;
  wire       [15:0]   _zz_15289;
  wire       [15:0]   _zz_15290;
  wire       [15:0]   _zz_15291;
  wire       [15:0]   _zz_15292;
  wire       [15:0]   _zz_15293;
  wire       [15:0]   _zz_15294;
  wire       [15:0]   _zz_15295;
  wire       [15:0]   _zz_15296;
  wire       [15:0]   _zz_15297;
  wire       [15:0]   _zz_15298;
  wire       [15:0]   _zz_15299;
  wire       [15:0]   _zz_15300;
  wire       [15:0]   _zz_15301;
  wire       [15:0]   _zz_15302;
  wire       [15:0]   _zz_15303;
  wire       [15:0]   _zz_15304;
  wire       [15:0]   _zz_15305;
  wire       [15:0]   _zz_15306;
  wire       [15:0]   _zz_15307;
  wire       [15:0]   _zz_15308;
  wire       [15:0]   _zz_15309;
  wire       [15:0]   _zz_15310;
  wire       [15:0]   _zz_15311;
  wire       [15:0]   _zz_15312;
  wire       [15:0]   _zz_15313;
  wire       [15:0]   _zz_15314;
  wire       [15:0]   _zz_15315;
  wire       [15:0]   _zz_15316;
  wire       [15:0]   _zz_15317;
  wire       [15:0]   _zz_15318;
  wire       [15:0]   _zz_15319;
  wire       [15:0]   _zz_15320;
  wire       [15:0]   _zz_15321;
  wire       [15:0]   _zz_15322;
  wire       [15:0]   _zz_15323;
  wire       [15:0]   _zz_15324;
  wire       [15:0]   _zz_15325;
  wire       [15:0]   _zz_15326;
  wire       [15:0]   _zz_15327;
  wire       [15:0]   _zz_15328;
  wire       [15:0]   _zz_15329;
  wire       [15:0]   _zz_15330;
  wire       [15:0]   _zz_15331;
  wire       [15:0]   _zz_15332;
  wire       [15:0]   _zz_15333;
  wire       [15:0]   _zz_15334;
  wire       [15:0]   _zz_15335;
  wire       [15:0]   _zz_15336;
  wire       [15:0]   _zz_15337;
  wire       [15:0]   _zz_15338;
  wire       [15:0]   _zz_15339;
  wire       [15:0]   _zz_15340;
  wire       [15:0]   _zz_15341;
  wire       [15:0]   _zz_15342;
  wire       [15:0]   _zz_15343;
  wire       [15:0]   _zz_15344;
  wire       [15:0]   _zz_15345;
  wire       [15:0]   _zz_15346;
  wire       [15:0]   _zz_15347;
  wire       [15:0]   _zz_15348;
  wire       [15:0]   _zz_15349;
  wire       [15:0]   _zz_15350;
  wire       [15:0]   _zz_15351;
  wire       [15:0]   _zz_15352;
  wire       [15:0]   _zz_15353;
  wire       [15:0]   _zz_15354;
  wire       [15:0]   _zz_15355;
  wire       [15:0]   _zz_15356;
  wire       [15:0]   _zz_15357;
  wire       [15:0]   _zz_15358;
  wire       [15:0]   _zz_15359;
  wire       [15:0]   _zz_15360;
  wire       [15:0]   _zz_15361;
  wire       [15:0]   _zz_15362;
  wire       [15:0]   _zz_15363;
  wire       [15:0]   _zz_15364;
  wire       [15:0]   _zz_15365;
  wire       [15:0]   _zz_15366;
  wire       [15:0]   _zz_15367;
  wire       [15:0]   _zz_15368;
  wire       [15:0]   _zz_15369;
  wire       [15:0]   _zz_15370;
  wire       [15:0]   _zz_15371;
  wire       [15:0]   _zz_15372;
  wire       [15:0]   _zz_15373;
  wire       [15:0]   _zz_15374;
  wire       [15:0]   _zz_15375;
  wire       [15:0]   _zz_15376;
  wire       [15:0]   _zz_15377;
  wire       [15:0]   _zz_15378;
  wire       [15:0]   _zz_15379;
  wire       [15:0]   _zz_15380;
  wire       [15:0]   _zz_15381;
  wire       [15:0]   _zz_15382;
  wire       [15:0]   _zz_15383;
  wire       [15:0]   _zz_15384;
  wire       [15:0]   _zz_15385;
  wire       [15:0]   _zz_15386;
  wire       [15:0]   _zz_15387;
  wire       [15:0]   _zz_15388;
  wire       [15:0]   _zz_15389;
  wire       [15:0]   _zz_15390;
  wire       [15:0]   _zz_15391;
  wire       [15:0]   _zz_15392;
  wire       [15:0]   _zz_15393;
  wire       [15:0]   _zz_15394;
  wire       [15:0]   _zz_15395;
  wire       [15:0]   _zz_15396;
  wire       [15:0]   _zz_15397;
  wire       [15:0]   _zz_15398;
  wire       [15:0]   _zz_15399;
  wire       [15:0]   _zz_15400;
  wire       [15:0]   _zz_15401;
  wire       [15:0]   _zz_15402;
  wire       [15:0]   _zz_15403;
  wire       [15:0]   _zz_15404;
  wire       [15:0]   _zz_15405;
  wire       [15:0]   _zz_15406;
  wire       [15:0]   _zz_15407;
  wire       [15:0]   _zz_15408;
  wire       [15:0]   _zz_15409;
  wire       [15:0]   _zz_15410;
  wire       [15:0]   _zz_15411;
  wire       [15:0]   _zz_15412;
  wire       [15:0]   _zz_15413;
  wire       [15:0]   _zz_15414;
  wire       [15:0]   _zz_15415;
  wire       [15:0]   _zz_15416;
  wire       [15:0]   _zz_15417;
  wire       [15:0]   _zz_15418;
  wire       [15:0]   _zz_15419;
  wire       [15:0]   _zz_15420;
  wire       [15:0]   _zz_15421;
  wire       [15:0]   _zz_15422;
  wire       [15:0]   _zz_15423;
  wire       [15:0]   _zz_15424;
  wire       [15:0]   _zz_15425;
  wire       [15:0]   _zz_15426;
  wire       [15:0]   _zz_15427;
  wire       [15:0]   _zz_15428;
  wire       [15:0]   _zz_15429;
  wire       [15:0]   _zz_15430;
  wire       [15:0]   _zz_15431;
  wire       [15:0]   _zz_15432;
  wire       [15:0]   _zz_15433;
  wire       [15:0]   _zz_15434;
  wire       [15:0]   _zz_15435;
  wire       [15:0]   _zz_15436;
  wire       [15:0]   _zz_15437;
  wire       [15:0]   _zz_15438;
  wire       [15:0]   _zz_15439;
  wire       [15:0]   _zz_15440;
  wire       [15:0]   _zz_15441;
  wire       [15:0]   _zz_15442;
  wire       [15:0]   _zz_15443;
  wire       [15:0]   _zz_15444;
  wire       [15:0]   _zz_15445;
  wire       [15:0]   _zz_15446;
  wire       [15:0]   _zz_15447;
  wire       [15:0]   _zz_15448;
  wire       [15:0]   _zz_15449;
  wire       [15:0]   _zz_15450;
  wire       [15:0]   _zz_15451;
  wire       [15:0]   _zz_15452;
  wire       [15:0]   _zz_15453;
  wire       [15:0]   _zz_15454;
  wire       [15:0]   _zz_15455;
  wire       [15:0]   _zz_15456;
  wire       [15:0]   _zz_15457;
  wire       [15:0]   _zz_15458;
  wire       [15:0]   _zz_15459;
  wire       [15:0]   _zz_15460;
  wire       [15:0]   _zz_15461;
  wire       [15:0]   _zz_15462;
  wire       [15:0]   _zz_15463;
  wire       [15:0]   _zz_15464;
  wire       [15:0]   _zz_15465;
  wire       [15:0]   _zz_15466;
  wire       [15:0]   _zz_15467;
  wire       [15:0]   _zz_15468;
  wire       [15:0]   _zz_15469;
  wire       [15:0]   _zz_15470;
  wire       [15:0]   _zz_15471;
  wire       [15:0]   _zz_15472;
  wire       [15:0]   _zz_15473;
  wire       [15:0]   _zz_15474;
  wire       [15:0]   _zz_15475;
  wire       [15:0]   _zz_15476;
  wire       [15:0]   _zz_15477;
  wire       [15:0]   _zz_15478;
  wire       [15:0]   _zz_15479;
  wire       [15:0]   _zz_15480;
  wire       [15:0]   _zz_15481;
  wire       [15:0]   _zz_15482;
  wire       [15:0]   _zz_15483;
  wire       [15:0]   _zz_15484;
  wire       [15:0]   _zz_15485;
  wire       [15:0]   _zz_15486;
  wire       [15:0]   _zz_15487;
  wire       [15:0]   _zz_15488;
  wire       [15:0]   _zz_15489;
  wire       [15:0]   _zz_15490;
  wire       [15:0]   _zz_15491;
  wire       [15:0]   _zz_15492;
  wire       [15:0]   _zz_15493;
  wire       [15:0]   _zz_15494;
  wire       [15:0]   _zz_15495;
  wire       [15:0]   _zz_15496;
  wire       [15:0]   _zz_15497;
  wire       [15:0]   _zz_15498;
  wire       [15:0]   _zz_15499;
  wire       [15:0]   _zz_15500;
  wire       [15:0]   _zz_15501;
  wire       [15:0]   _zz_15502;
  wire       [15:0]   _zz_15503;
  wire       [15:0]   _zz_15504;
  wire       [15:0]   _zz_15505;
  wire       [15:0]   _zz_15506;
  wire       [15:0]   _zz_15507;
  wire       [15:0]   _zz_15508;
  wire       [15:0]   _zz_15509;
  wire       [15:0]   _zz_15510;
  wire       [15:0]   _zz_15511;
  wire       [15:0]   _zz_15512;
  wire       [15:0]   _zz_15513;
  wire       [15:0]   _zz_15514;
  wire       [15:0]   _zz_15515;
  wire       [15:0]   _zz_15516;
  wire       [15:0]   _zz_15517;
  wire       [15:0]   _zz_15518;
  wire       [15:0]   _zz_15519;
  wire       [15:0]   _zz_15520;
  wire       [15:0]   _zz_15521;
  wire       [15:0]   _zz_15522;
  wire       [15:0]   _zz_15523;
  wire       [15:0]   _zz_15524;
  wire       [15:0]   _zz_15525;
  wire       [15:0]   _zz_15526;
  wire       [15:0]   _zz_15527;
  wire       [15:0]   _zz_15528;
  wire       [15:0]   _zz_15529;
  wire       [15:0]   _zz_15530;
  wire       [15:0]   _zz_15531;
  wire       [15:0]   _zz_15532;
  wire       [15:0]   _zz_15533;
  wire       [15:0]   _zz_15534;
  wire       [15:0]   _zz_15535;
  wire       [15:0]   _zz_15536;
  wire       [15:0]   _zz_15537;
  wire       [15:0]   _zz_15538;
  wire       [15:0]   _zz_15539;
  wire       [15:0]   _zz_15540;
  wire       [15:0]   _zz_15541;
  wire       [15:0]   _zz_15542;
  wire       [15:0]   _zz_15543;
  wire       [15:0]   _zz_15544;
  wire       [15:0]   _zz_15545;
  wire       [15:0]   _zz_15546;
  wire       [15:0]   _zz_15547;
  wire       [15:0]   _zz_15548;
  wire       [15:0]   _zz_15549;
  wire       [15:0]   _zz_15550;
  wire       [15:0]   _zz_15551;
  wire       [15:0]   _zz_15552;
  wire       [15:0]   _zz_15553;
  wire       [15:0]   _zz_15554;
  wire       [15:0]   _zz_15555;
  wire       [15:0]   _zz_15556;
  wire       [15:0]   _zz_15557;
  wire       [15:0]   _zz_15558;
  wire       [15:0]   _zz_15559;
  wire       [15:0]   _zz_15560;
  wire       [15:0]   _zz_15561;
  wire       [15:0]   _zz_15562;
  wire       [15:0]   _zz_15563;
  wire       [15:0]   _zz_15564;
  wire       [15:0]   _zz_15565;
  wire       [15:0]   _zz_15566;
  wire       [15:0]   _zz_15567;
  wire       [15:0]   _zz_15568;
  wire       [15:0]   _zz_15569;
  wire       [15:0]   _zz_15570;
  wire       [15:0]   _zz_15571;
  wire       [15:0]   _zz_15572;
  wire       [15:0]   _zz_15573;
  wire       [15:0]   _zz_15574;
  wire       [15:0]   _zz_15575;
  wire       [15:0]   _zz_15576;
  wire       [15:0]   _zz_15577;
  wire       [15:0]   _zz_15578;
  wire       [15:0]   _zz_15579;
  wire       [15:0]   _zz_15580;
  wire       [15:0]   _zz_15581;
  wire       [15:0]   _zz_15582;
  wire       [15:0]   _zz_15583;
  wire       [15:0]   _zz_15584;
  wire       [15:0]   _zz_15585;
  wire       [15:0]   _zz_15586;
  wire       [15:0]   _zz_15587;
  wire       [15:0]   _zz_15588;
  wire       [15:0]   _zz_15589;
  wire       [15:0]   _zz_15590;
  wire       [15:0]   _zz_15591;
  wire       [15:0]   _zz_15592;
  wire       [15:0]   _zz_15593;
  wire       [15:0]   _zz_15594;
  wire       [15:0]   _zz_15595;
  wire       [15:0]   _zz_15596;
  wire       [15:0]   _zz_15597;
  wire       [15:0]   _zz_15598;
  wire       [15:0]   _zz_15599;
  wire       [15:0]   _zz_15600;
  wire       [15:0]   _zz_15601;
  wire       [15:0]   _zz_15602;
  wire       [15:0]   _zz_15603;
  wire       [15:0]   _zz_15604;
  wire       [15:0]   _zz_15605;
  wire       [15:0]   _zz_15606;
  wire       [15:0]   _zz_15607;
  wire       [15:0]   _zz_15608;
  wire       [15:0]   _zz_15609;
  wire       [15:0]   _zz_15610;
  wire       [15:0]   _zz_15611;
  wire       [15:0]   _zz_15612;
  wire       [15:0]   _zz_15613;
  wire       [15:0]   _zz_15614;
  wire       [15:0]   _zz_15615;
  wire       [15:0]   _zz_15616;
  wire       [15:0]   _zz_15617;
  wire       [15:0]   _zz_15618;
  wire       [15:0]   _zz_15619;
  wire       [15:0]   _zz_15620;
  wire       [15:0]   _zz_15621;
  wire       [15:0]   _zz_15622;
  wire       [15:0]   _zz_15623;
  wire       [15:0]   _zz_15624;
  wire       [15:0]   _zz_15625;
  wire       [15:0]   _zz_15626;
  wire       [15:0]   _zz_15627;
  wire       [15:0]   _zz_15628;
  wire       [15:0]   _zz_15629;
  wire       [15:0]   _zz_15630;
  wire       [15:0]   _zz_15631;
  wire       [15:0]   _zz_15632;
  wire       [15:0]   _zz_15633;
  wire       [15:0]   _zz_15634;
  wire       [15:0]   _zz_15635;
  wire       [15:0]   _zz_15636;
  wire       [15:0]   _zz_15637;
  wire       [15:0]   _zz_15638;
  wire       [15:0]   _zz_15639;
  wire       [15:0]   _zz_15640;
  wire       [15:0]   _zz_15641;
  wire       [15:0]   _zz_15642;
  wire       [15:0]   _zz_15643;
  wire       [15:0]   _zz_15644;
  wire       [15:0]   _zz_15645;
  wire       [15:0]   _zz_15646;
  wire       [15:0]   _zz_15647;
  wire       [15:0]   _zz_15648;
  wire       [15:0]   _zz_15649;
  wire       [15:0]   _zz_15650;
  wire       [15:0]   _zz_15651;
  wire       [15:0]   _zz_15652;
  wire       [15:0]   _zz_15653;
  wire       [15:0]   _zz_15654;
  wire       [15:0]   _zz_15655;
  wire       [15:0]   _zz_15656;
  wire       [15:0]   _zz_15657;
  wire       [15:0]   _zz_15658;
  wire       [15:0]   _zz_15659;
  wire       [15:0]   _zz_15660;
  wire       [15:0]   _zz_15661;
  wire       [15:0]   _zz_15662;
  wire       [15:0]   _zz_15663;
  wire       [15:0]   _zz_15664;
  wire       [15:0]   _zz_15665;
  wire       [15:0]   _zz_15666;
  wire       [15:0]   _zz_15667;
  wire       [15:0]   _zz_15668;
  wire       [15:0]   _zz_15669;
  wire       [15:0]   _zz_15670;
  wire       [15:0]   _zz_15671;
  wire       [15:0]   _zz_15672;
  wire       [15:0]   _zz_15673;
  wire       [15:0]   _zz_15674;
  wire       [15:0]   _zz_15675;
  wire       [15:0]   _zz_15676;
  wire       [15:0]   _zz_15677;
  wire       [15:0]   _zz_15678;
  wire       [15:0]   _zz_15679;
  wire       [15:0]   _zz_15680;
  wire       [15:0]   _zz_15681;
  wire       [15:0]   _zz_15682;
  wire       [15:0]   _zz_15683;
  wire       [15:0]   _zz_15684;
  wire       [15:0]   _zz_15685;
  wire       [15:0]   _zz_15686;
  wire       [15:0]   _zz_15687;
  wire       [15:0]   _zz_15688;
  wire       [15:0]   _zz_15689;
  wire       [15:0]   _zz_15690;
  wire       [15:0]   _zz_15691;
  wire       [15:0]   _zz_15692;
  wire       [15:0]   _zz_15693;
  wire       [15:0]   _zz_15694;
  wire       [15:0]   _zz_15695;
  wire       [15:0]   _zz_15696;
  wire       [15:0]   _zz_15697;
  wire       [15:0]   _zz_15698;
  wire       [15:0]   _zz_15699;
  wire       [15:0]   _zz_15700;
  wire       [15:0]   _zz_15701;
  wire       [15:0]   _zz_15702;
  wire       [15:0]   _zz_15703;
  wire       [15:0]   _zz_15704;
  wire       [15:0]   _zz_15705;
  wire       [15:0]   _zz_15706;
  wire       [15:0]   _zz_15707;
  wire       [15:0]   _zz_15708;
  wire       [15:0]   _zz_15709;
  wire       [15:0]   _zz_15710;
  wire       [15:0]   _zz_15711;
  wire       [15:0]   _zz_15712;
  wire       [15:0]   _zz_15713;
  wire       [15:0]   _zz_15714;
  wire       [15:0]   _zz_15715;
  wire       [15:0]   _zz_15716;
  wire       [15:0]   _zz_15717;
  wire       [15:0]   _zz_15718;
  wire       [15:0]   _zz_15719;
  wire       [15:0]   _zz_15720;
  wire       [15:0]   _zz_15721;
  wire       [15:0]   _zz_15722;
  wire       [15:0]   _zz_15723;
  wire       [15:0]   _zz_15724;
  wire       [15:0]   _zz_15725;
  wire       [15:0]   _zz_15726;
  wire       [15:0]   _zz_15727;
  wire       [15:0]   _zz_15728;
  wire       [15:0]   _zz_15729;
  wire       [15:0]   _zz_15730;
  wire       [15:0]   _zz_15731;
  wire       [15:0]   _zz_15732;
  wire       [15:0]   _zz_15733;
  wire       [15:0]   _zz_15734;
  wire       [15:0]   _zz_15735;
  wire       [15:0]   _zz_15736;
  wire       [15:0]   _zz_15737;
  wire       [15:0]   _zz_15738;
  wire       [15:0]   _zz_15739;
  wire       [15:0]   _zz_15740;
  wire       [15:0]   _zz_15741;
  wire       [15:0]   _zz_15742;
  wire       [15:0]   _zz_15743;
  wire       [15:0]   _zz_15744;
  wire       [15:0]   _zz_15745;
  wire       [15:0]   _zz_15746;
  wire       [15:0]   _zz_15747;
  wire       [15:0]   _zz_15748;
  wire       [15:0]   _zz_15749;
  wire       [15:0]   _zz_15750;
  wire       [15:0]   _zz_15751;
  wire       [15:0]   _zz_15752;
  wire       [15:0]   _zz_15753;
  wire       [15:0]   _zz_15754;
  wire       [15:0]   _zz_15755;
  wire       [15:0]   _zz_15756;
  wire       [15:0]   _zz_15757;
  wire       [15:0]   _zz_15758;
  wire       [15:0]   _zz_15759;
  wire       [15:0]   _zz_15760;
  wire       [15:0]   _zz_15761;
  wire       [15:0]   _zz_15762;
  wire       [15:0]   _zz_15763;
  wire       [15:0]   _zz_15764;
  wire       [15:0]   _zz_15765;
  wire       [15:0]   _zz_15766;
  wire       [15:0]   _zz_15767;
  wire       [15:0]   _zz_15768;
  wire       [15:0]   _zz_15769;
  wire       [15:0]   _zz_15770;
  wire       [15:0]   _zz_15771;
  wire       [15:0]   _zz_15772;
  wire       [15:0]   _zz_15773;
  wire       [15:0]   _zz_15774;
  wire       [15:0]   _zz_15775;
  wire       [15:0]   _zz_15776;
  wire       [15:0]   _zz_15777;
  wire       [15:0]   _zz_15778;
  wire       [15:0]   _zz_15779;
  wire       [15:0]   _zz_15780;
  wire       [15:0]   _zz_15781;
  wire       [15:0]   _zz_15782;
  wire       [15:0]   _zz_15783;
  wire       [15:0]   _zz_15784;
  wire       [15:0]   _zz_15785;
  wire       [15:0]   _zz_15786;
  wire       [15:0]   _zz_15787;
  wire       [15:0]   _zz_15788;
  wire       [15:0]   _zz_15789;
  wire       [15:0]   _zz_15790;
  wire       [15:0]   _zz_15791;
  wire       [15:0]   _zz_15792;
  wire       [15:0]   _zz_15793;
  wire       [15:0]   _zz_15794;
  wire       [15:0]   _zz_15795;
  wire       [15:0]   _zz_15796;
  wire       [15:0]   _zz_15797;
  wire       [15:0]   _zz_15798;
  wire       [15:0]   _zz_15799;
  wire       [15:0]   _zz_15800;
  wire       [15:0]   _zz_15801;
  wire       [15:0]   _zz_15802;
  wire       [15:0]   _zz_15803;
  wire       [15:0]   _zz_15804;
  wire       [15:0]   _zz_15805;
  wire       [15:0]   _zz_15806;
  wire       [15:0]   _zz_15807;
  wire       [15:0]   _zz_15808;
  wire       [15:0]   _zz_15809;
  wire       [15:0]   _zz_15810;
  wire       [15:0]   _zz_15811;
  wire       [15:0]   _zz_15812;
  wire       [15:0]   _zz_15813;
  wire       [15:0]   _zz_15814;
  wire       [15:0]   _zz_15815;
  wire       [15:0]   _zz_15816;
  wire       [15:0]   _zz_15817;
  wire       [15:0]   _zz_15818;
  wire       [15:0]   _zz_15819;
  wire       [15:0]   _zz_15820;
  wire       [15:0]   _zz_15821;
  wire       [15:0]   _zz_15822;
  wire       [15:0]   _zz_15823;
  wire       [15:0]   _zz_15824;
  wire       [15:0]   _zz_15825;
  wire       [15:0]   _zz_15826;
  wire       [15:0]   _zz_15827;
  wire       [15:0]   _zz_15828;
  wire       [15:0]   _zz_15829;
  wire       [15:0]   _zz_15830;
  wire       [15:0]   _zz_15831;
  wire       [15:0]   _zz_15832;
  wire       [15:0]   _zz_15833;
  wire       [15:0]   _zz_15834;
  wire       [15:0]   _zz_15835;
  wire       [15:0]   _zz_15836;
  wire       [15:0]   _zz_15837;
  wire       [15:0]   _zz_15838;
  wire       [15:0]   _zz_15839;
  wire       [15:0]   _zz_15840;
  wire       [15:0]   _zz_15841;
  wire       [15:0]   _zz_15842;
  wire       [15:0]   _zz_15843;
  wire       [15:0]   _zz_15844;
  wire       [15:0]   _zz_15845;
  wire       [15:0]   _zz_15846;
  wire       [15:0]   _zz_15847;
  wire       [15:0]   _zz_15848;
  wire       [15:0]   _zz_15849;
  wire       [15:0]   _zz_15850;
  wire       [15:0]   _zz_15851;
  wire       [15:0]   _zz_15852;
  wire       [15:0]   _zz_15853;
  wire       [15:0]   _zz_15854;
  wire       [15:0]   _zz_15855;
  wire       [15:0]   _zz_15856;
  wire       [15:0]   _zz_15857;
  wire       [15:0]   _zz_15858;
  wire       [15:0]   _zz_15859;
  wire       [15:0]   _zz_15860;
  wire       [15:0]   _zz_15861;
  wire       [15:0]   _zz_15862;
  wire       [15:0]   _zz_15863;
  wire       [15:0]   _zz_15864;
  wire       [15:0]   _zz_15865;
  wire       [15:0]   _zz_15866;
  wire       [15:0]   _zz_15867;
  wire       [15:0]   _zz_15868;
  wire       [15:0]   _zz_15869;
  wire       [15:0]   _zz_15870;
  wire       [15:0]   _zz_15871;
  wire       [15:0]   _zz_15872;
  wire       [15:0]   _zz_15873;
  wire       [15:0]   _zz_15874;
  wire       [15:0]   _zz_15875;
  wire       [15:0]   _zz_15876;
  wire       [15:0]   _zz_15877;
  wire       [15:0]   _zz_15878;
  wire       [15:0]   _zz_15879;
  wire       [15:0]   _zz_15880;
  wire       [15:0]   _zz_15881;
  wire       [15:0]   _zz_15882;
  wire       [15:0]   _zz_15883;
  wire       [15:0]   _zz_15884;
  wire       [15:0]   _zz_15885;
  wire       [15:0]   _zz_15886;
  wire       [15:0]   _zz_15887;
  wire       [15:0]   _zz_15888;
  wire       [15:0]   _zz_15889;
  wire       [15:0]   _zz_15890;
  wire       [15:0]   _zz_15891;
  wire       [15:0]   _zz_15892;
  wire       [15:0]   _zz_15893;
  wire       [15:0]   _zz_15894;
  wire       [15:0]   _zz_15895;
  wire       [15:0]   _zz_15896;
  wire       [15:0]   _zz_15897;
  wire       [15:0]   _zz_15898;
  wire       [15:0]   _zz_15899;
  wire       [15:0]   _zz_15900;
  wire       [15:0]   _zz_15901;
  wire       [15:0]   _zz_15902;
  wire       [15:0]   _zz_15903;
  wire       [15:0]   _zz_15904;
  wire       [15:0]   _zz_15905;
  wire       [15:0]   _zz_15906;
  wire       [15:0]   _zz_15907;
  wire       [15:0]   _zz_15908;
  wire       [15:0]   _zz_15909;
  wire       [15:0]   _zz_15910;
  wire       [15:0]   _zz_15911;
  wire       [15:0]   _zz_15912;
  wire       [15:0]   _zz_15913;
  wire       [15:0]   _zz_15914;
  wire       [15:0]   _zz_15915;
  wire       [15:0]   _zz_15916;
  wire       [15:0]   _zz_15917;
  wire       [15:0]   _zz_15918;
  wire       [15:0]   _zz_15919;
  wire       [15:0]   _zz_15920;
  wire       [15:0]   _zz_15921;
  wire       [15:0]   _zz_15922;
  wire       [15:0]   _zz_15923;
  wire       [15:0]   _zz_15924;
  wire       [15:0]   _zz_15925;
  wire       [15:0]   _zz_15926;
  wire       [15:0]   _zz_15927;
  wire       [15:0]   _zz_15928;
  wire       [15:0]   _zz_15929;
  wire       [15:0]   _zz_15930;
  wire       [15:0]   _zz_15931;
  wire       [15:0]   _zz_15932;
  wire       [15:0]   _zz_15933;
  wire       [15:0]   _zz_15934;
  wire       [15:0]   _zz_15935;
  wire       [15:0]   _zz_15936;
  wire       [15:0]   _zz_15937;
  wire       [15:0]   _zz_15938;
  wire       [15:0]   _zz_15939;
  wire       [15:0]   _zz_15940;
  wire       [15:0]   _zz_15941;
  wire       [15:0]   _zz_15942;
  wire       [15:0]   _zz_15943;
  wire       [15:0]   _zz_15944;
  wire       [15:0]   _zz_15945;
  wire       [15:0]   _zz_15946;
  wire       [15:0]   _zz_15947;
  wire       [15:0]   _zz_15948;
  wire       [15:0]   _zz_15949;
  wire       [15:0]   _zz_15950;
  wire       [15:0]   _zz_15951;
  wire       [15:0]   _zz_15952;
  wire       [15:0]   _zz_15953;
  wire       [15:0]   _zz_15954;
  wire       [15:0]   _zz_15955;
  wire       [15:0]   _zz_15956;
  wire       [15:0]   _zz_15957;
  wire       [15:0]   _zz_15958;
  wire       [15:0]   _zz_15959;
  wire       [15:0]   _zz_15960;
  wire       [15:0]   _zz_15961;
  wire       [15:0]   _zz_15962;
  wire       [15:0]   _zz_15963;
  wire       [15:0]   _zz_15964;
  wire       [15:0]   _zz_15965;
  wire       [15:0]   _zz_15966;
  wire       [15:0]   _zz_15967;
  wire       [15:0]   _zz_15968;
  wire       [15:0]   _zz_15969;
  wire       [15:0]   _zz_15970;
  wire       [15:0]   _zz_15971;
  wire       [15:0]   _zz_15972;
  wire       [15:0]   _zz_15973;
  wire       [15:0]   _zz_15974;
  wire       [15:0]   _zz_15975;
  wire       [15:0]   _zz_15976;
  wire       [15:0]   _zz_15977;
  wire       [15:0]   _zz_15978;
  wire       [15:0]   _zz_15979;
  wire       [15:0]   _zz_15980;
  wire       [15:0]   _zz_15981;
  wire       [15:0]   _zz_15982;
  wire       [15:0]   _zz_15983;
  wire       [15:0]   _zz_15984;
  wire       [15:0]   _zz_15985;
  wire       [15:0]   _zz_15986;
  wire       [15:0]   _zz_15987;
  wire       [15:0]   _zz_15988;
  wire       [15:0]   _zz_15989;
  wire       [15:0]   _zz_15990;
  wire       [15:0]   _zz_15991;
  wire       [15:0]   _zz_15992;
  wire       [15:0]   _zz_15993;
  wire       [15:0]   _zz_15994;
  wire       [15:0]   _zz_15995;
  wire       [15:0]   _zz_15996;
  wire       [15:0]   _zz_15997;
  wire       [15:0]   _zz_15998;
  wire       [15:0]   _zz_15999;
  wire       [15:0]   _zz_16000;
  wire       [15:0]   _zz_16001;
  wire       [15:0]   _zz_16002;
  wire       [15:0]   _zz_16003;
  wire       [15:0]   _zz_16004;
  wire       [15:0]   _zz_16005;
  wire       [15:0]   _zz_16006;
  wire       [15:0]   _zz_16007;
  wire       [15:0]   _zz_16008;
  wire       [15:0]   _zz_16009;
  wire       [15:0]   _zz_16010;
  wire       [15:0]   _zz_16011;
  wire       [15:0]   _zz_16012;
  wire       [15:0]   _zz_16013;
  wire       [15:0]   _zz_16014;
  wire       [15:0]   _zz_16015;
  wire       [15:0]   _zz_16016;
  wire       [15:0]   _zz_16017;
  wire       [15:0]   _zz_16018;
  wire       [15:0]   _zz_16019;
  wire       [15:0]   _zz_16020;
  wire       [15:0]   _zz_16021;
  wire       [15:0]   _zz_16022;
  wire       [15:0]   _zz_16023;
  wire       [15:0]   _zz_16024;
  wire       [15:0]   _zz_16025;
  wire       [15:0]   _zz_16026;
  wire       [15:0]   _zz_16027;
  wire       [15:0]   _zz_16028;
  wire       [15:0]   _zz_16029;
  wire       [15:0]   _zz_16030;
  wire       [15:0]   _zz_16031;
  wire       [15:0]   _zz_16032;
  wire       [15:0]   _zz_16033;
  wire       [15:0]   _zz_16034;
  wire       [15:0]   _zz_16035;
  wire       [15:0]   _zz_16036;
  wire       [15:0]   _zz_16037;
  wire       [15:0]   _zz_16038;
  wire       [15:0]   _zz_16039;
  wire       [15:0]   _zz_16040;
  wire       [15:0]   _zz_16041;
  wire       [15:0]   _zz_16042;
  wire       [15:0]   _zz_16043;
  wire       [15:0]   _zz_16044;
  wire       [15:0]   _zz_16045;
  wire       [15:0]   _zz_16046;
  wire       [15:0]   _zz_16047;
  wire       [15:0]   _zz_16048;
  wire       [15:0]   _zz_16049;
  wire       [15:0]   _zz_16050;
  wire       [15:0]   _zz_16051;
  wire       [15:0]   _zz_16052;
  wire       [15:0]   _zz_16053;
  wire       [15:0]   _zz_16054;
  wire       [15:0]   _zz_16055;
  wire       [15:0]   _zz_16056;
  wire       [15:0]   _zz_16057;
  wire       [15:0]   _zz_16058;
  wire       [15:0]   _zz_16059;
  wire       [15:0]   _zz_16060;
  wire       [15:0]   _zz_16061;
  wire       [15:0]   _zz_16062;
  wire       [15:0]   _zz_16063;
  wire       [15:0]   _zz_16064;
  wire       [15:0]   _zz_16065;
  wire       [15:0]   _zz_16066;
  wire       [15:0]   _zz_16067;
  wire       [15:0]   _zz_16068;
  wire       [15:0]   _zz_16069;
  wire       [15:0]   _zz_16070;
  wire       [15:0]   _zz_16071;
  wire       [15:0]   _zz_16072;
  wire       [15:0]   _zz_16073;
  wire       [15:0]   _zz_16074;
  wire       [15:0]   _zz_16075;
  wire       [15:0]   _zz_16076;
  wire       [15:0]   _zz_16077;
  wire       [15:0]   _zz_16078;
  wire       [15:0]   _zz_16079;
  wire       [15:0]   _zz_16080;
  wire       [15:0]   _zz_16081;
  wire       [15:0]   _zz_16082;
  wire       [15:0]   _zz_16083;
  wire       [15:0]   _zz_16084;
  wire       [15:0]   _zz_16085;
  wire       [15:0]   _zz_16086;
  wire       [15:0]   _zz_16087;
  wire       [15:0]   _zz_16088;
  wire       [15:0]   _zz_16089;
  wire       [15:0]   _zz_16090;
  wire       [15:0]   _zz_16091;
  wire       [15:0]   _zz_16092;
  wire       [15:0]   _zz_16093;
  wire       [15:0]   _zz_16094;
  wire       [15:0]   _zz_16095;
  wire       [15:0]   _zz_16096;
  wire       [15:0]   _zz_16097;
  wire       [15:0]   _zz_16098;
  wire       [15:0]   _zz_16099;
  wire       [15:0]   _zz_16100;
  wire       [15:0]   _zz_16101;
  wire       [15:0]   _zz_16102;
  wire       [15:0]   _zz_16103;
  wire       [15:0]   _zz_16104;
  wire       [15:0]   _zz_16105;
  wire       [15:0]   _zz_16106;
  wire       [15:0]   _zz_16107;
  wire       [15:0]   _zz_16108;
  wire       [15:0]   _zz_16109;
  wire       [15:0]   _zz_16110;
  wire       [15:0]   _zz_16111;
  wire       [15:0]   _zz_16112;
  wire       [15:0]   _zz_16113;
  wire       [15:0]   _zz_16114;
  wire       [15:0]   _zz_16115;
  wire       [15:0]   _zz_16116;
  wire       [15:0]   _zz_16117;
  wire       [15:0]   _zz_16118;
  wire       [15:0]   _zz_16119;
  wire       [15:0]   _zz_16120;
  wire       [15:0]   _zz_16121;
  wire       [15:0]   _zz_16122;
  wire       [15:0]   _zz_16123;
  wire       [15:0]   _zz_16124;
  wire       [15:0]   _zz_16125;
  wire       [15:0]   _zz_16126;
  wire       [15:0]   _zz_16127;
  wire       [15:0]   _zz_16128;
  wire       [15:0]   _zz_16129;
  wire       [15:0]   _zz_16130;
  wire       [15:0]   _zz_16131;
  wire       [15:0]   _zz_16132;
  wire       [15:0]   _zz_16133;
  wire       [15:0]   _zz_16134;
  wire       [0:0]    _zz_16135;
  wire       [3:0]    _zz_16136;
  reg        [15:0]   data_in_0_real;
  reg        [15:0]   data_in_0_imag;
  reg        [15:0]   data_in_1_real;
  reg        [15:0]   data_in_1_imag;
  reg        [15:0]   data_in_2_real;
  reg        [15:0]   data_in_2_imag;
  reg        [15:0]   data_in_3_real;
  reg        [15:0]   data_in_3_imag;
  reg        [15:0]   data_in_4_real;
  reg        [15:0]   data_in_4_imag;
  reg        [15:0]   data_in_5_real;
  reg        [15:0]   data_in_5_imag;
  reg        [15:0]   data_in_6_real;
  reg        [15:0]   data_in_6_imag;
  reg        [15:0]   data_in_7_real;
  reg        [15:0]   data_in_7_imag;
  reg        [15:0]   data_in_8_real;
  reg        [15:0]   data_in_8_imag;
  reg        [15:0]   data_in_9_real;
  reg        [15:0]   data_in_9_imag;
  reg        [15:0]   data_in_10_real;
  reg        [15:0]   data_in_10_imag;
  reg        [15:0]   data_in_11_real;
  reg        [15:0]   data_in_11_imag;
  reg        [15:0]   data_in_12_real;
  reg        [15:0]   data_in_12_imag;
  reg        [15:0]   data_in_13_real;
  reg        [15:0]   data_in_13_imag;
  reg        [15:0]   data_in_14_real;
  reg        [15:0]   data_in_14_imag;
  reg        [15:0]   data_in_15_real;
  reg        [15:0]   data_in_15_imag;
  reg        [15:0]   data_in_16_real;
  reg        [15:0]   data_in_16_imag;
  reg        [15:0]   data_in_17_real;
  reg        [15:0]   data_in_17_imag;
  reg        [15:0]   data_in_18_real;
  reg        [15:0]   data_in_18_imag;
  reg        [15:0]   data_in_19_real;
  reg        [15:0]   data_in_19_imag;
  reg        [15:0]   data_in_20_real;
  reg        [15:0]   data_in_20_imag;
  reg        [15:0]   data_in_21_real;
  reg        [15:0]   data_in_21_imag;
  reg        [15:0]   data_in_22_real;
  reg        [15:0]   data_in_22_imag;
  reg        [15:0]   data_in_23_real;
  reg        [15:0]   data_in_23_imag;
  reg        [15:0]   data_in_24_real;
  reg        [15:0]   data_in_24_imag;
  reg        [15:0]   data_in_25_real;
  reg        [15:0]   data_in_25_imag;
  reg        [15:0]   data_in_26_real;
  reg        [15:0]   data_in_26_imag;
  reg        [15:0]   data_in_27_real;
  reg        [15:0]   data_in_27_imag;
  reg        [15:0]   data_in_28_real;
  reg        [15:0]   data_in_28_imag;
  reg        [15:0]   data_in_29_real;
  reg        [15:0]   data_in_29_imag;
  reg        [15:0]   data_in_30_real;
  reg        [15:0]   data_in_30_imag;
  reg        [15:0]   data_in_31_real;
  reg        [15:0]   data_in_31_imag;
  reg        [15:0]   data_in_32_real;
  reg        [15:0]   data_in_32_imag;
  reg        [15:0]   data_in_33_real;
  reg        [15:0]   data_in_33_imag;
  reg        [15:0]   data_in_34_real;
  reg        [15:0]   data_in_34_imag;
  reg        [15:0]   data_in_35_real;
  reg        [15:0]   data_in_35_imag;
  reg        [15:0]   data_in_36_real;
  reg        [15:0]   data_in_36_imag;
  reg        [15:0]   data_in_37_real;
  reg        [15:0]   data_in_37_imag;
  reg        [15:0]   data_in_38_real;
  reg        [15:0]   data_in_38_imag;
  reg        [15:0]   data_in_39_real;
  reg        [15:0]   data_in_39_imag;
  reg        [15:0]   data_in_40_real;
  reg        [15:0]   data_in_40_imag;
  reg        [15:0]   data_in_41_real;
  reg        [15:0]   data_in_41_imag;
  reg        [15:0]   data_in_42_real;
  reg        [15:0]   data_in_42_imag;
  reg        [15:0]   data_in_43_real;
  reg        [15:0]   data_in_43_imag;
  reg        [15:0]   data_in_44_real;
  reg        [15:0]   data_in_44_imag;
  reg        [15:0]   data_in_45_real;
  reg        [15:0]   data_in_45_imag;
  reg        [15:0]   data_in_46_real;
  reg        [15:0]   data_in_46_imag;
  reg        [15:0]   data_in_47_real;
  reg        [15:0]   data_in_47_imag;
  reg        [15:0]   data_in_48_real;
  reg        [15:0]   data_in_48_imag;
  reg        [15:0]   data_in_49_real;
  reg        [15:0]   data_in_49_imag;
  reg        [15:0]   data_in_50_real;
  reg        [15:0]   data_in_50_imag;
  reg        [15:0]   data_in_51_real;
  reg        [15:0]   data_in_51_imag;
  reg        [15:0]   data_in_52_real;
  reg        [15:0]   data_in_52_imag;
  reg        [15:0]   data_in_53_real;
  reg        [15:0]   data_in_53_imag;
  reg        [15:0]   data_in_54_real;
  reg        [15:0]   data_in_54_imag;
  reg        [15:0]   data_in_55_real;
  reg        [15:0]   data_in_55_imag;
  reg        [15:0]   data_in_56_real;
  reg        [15:0]   data_in_56_imag;
  reg        [15:0]   data_in_57_real;
  reg        [15:0]   data_in_57_imag;
  reg        [15:0]   data_in_58_real;
  reg        [15:0]   data_in_58_imag;
  reg        [15:0]   data_in_59_real;
  reg        [15:0]   data_in_59_imag;
  reg        [15:0]   data_in_60_real;
  reg        [15:0]   data_in_60_imag;
  reg        [15:0]   data_in_61_real;
  reg        [15:0]   data_in_61_imag;
  reg        [15:0]   data_in_62_real;
  reg        [15:0]   data_in_62_imag;
  reg        [15:0]   data_in_63_real;
  reg        [15:0]   data_in_63_imag;
  reg        [15:0]   data_in_64_real;
  reg        [15:0]   data_in_64_imag;
  reg        [15:0]   data_in_65_real;
  reg        [15:0]   data_in_65_imag;
  reg        [15:0]   data_in_66_real;
  reg        [15:0]   data_in_66_imag;
  reg        [15:0]   data_in_67_real;
  reg        [15:0]   data_in_67_imag;
  reg        [15:0]   data_in_68_real;
  reg        [15:0]   data_in_68_imag;
  reg        [15:0]   data_in_69_real;
  reg        [15:0]   data_in_69_imag;
  reg        [15:0]   data_in_70_real;
  reg        [15:0]   data_in_70_imag;
  reg        [15:0]   data_in_71_real;
  reg        [15:0]   data_in_71_imag;
  reg        [15:0]   data_in_72_real;
  reg        [15:0]   data_in_72_imag;
  reg        [15:0]   data_in_73_real;
  reg        [15:0]   data_in_73_imag;
  reg        [15:0]   data_in_74_real;
  reg        [15:0]   data_in_74_imag;
  reg        [15:0]   data_in_75_real;
  reg        [15:0]   data_in_75_imag;
  reg        [15:0]   data_in_76_real;
  reg        [15:0]   data_in_76_imag;
  reg        [15:0]   data_in_77_real;
  reg        [15:0]   data_in_77_imag;
  reg        [15:0]   data_in_78_real;
  reg        [15:0]   data_in_78_imag;
  reg        [15:0]   data_in_79_real;
  reg        [15:0]   data_in_79_imag;
  reg        [15:0]   data_in_80_real;
  reg        [15:0]   data_in_80_imag;
  reg        [15:0]   data_in_81_real;
  reg        [15:0]   data_in_81_imag;
  reg        [15:0]   data_in_82_real;
  reg        [15:0]   data_in_82_imag;
  reg        [15:0]   data_in_83_real;
  reg        [15:0]   data_in_83_imag;
  reg        [15:0]   data_in_84_real;
  reg        [15:0]   data_in_84_imag;
  reg        [15:0]   data_in_85_real;
  reg        [15:0]   data_in_85_imag;
  reg        [15:0]   data_in_86_real;
  reg        [15:0]   data_in_86_imag;
  reg        [15:0]   data_in_87_real;
  reg        [15:0]   data_in_87_imag;
  reg        [15:0]   data_in_88_real;
  reg        [15:0]   data_in_88_imag;
  reg        [15:0]   data_in_89_real;
  reg        [15:0]   data_in_89_imag;
  reg        [15:0]   data_in_90_real;
  reg        [15:0]   data_in_90_imag;
  reg        [15:0]   data_in_91_real;
  reg        [15:0]   data_in_91_imag;
  reg        [15:0]   data_in_92_real;
  reg        [15:0]   data_in_92_imag;
  reg        [15:0]   data_in_93_real;
  reg        [15:0]   data_in_93_imag;
  reg        [15:0]   data_in_94_real;
  reg        [15:0]   data_in_94_imag;
  reg        [15:0]   data_in_95_real;
  reg        [15:0]   data_in_95_imag;
  reg        [15:0]   data_in_96_real;
  reg        [15:0]   data_in_96_imag;
  reg        [15:0]   data_in_97_real;
  reg        [15:0]   data_in_97_imag;
  reg        [15:0]   data_in_98_real;
  reg        [15:0]   data_in_98_imag;
  reg        [15:0]   data_in_99_real;
  reg        [15:0]   data_in_99_imag;
  reg        [15:0]   data_in_100_real;
  reg        [15:0]   data_in_100_imag;
  reg        [15:0]   data_in_101_real;
  reg        [15:0]   data_in_101_imag;
  reg        [15:0]   data_in_102_real;
  reg        [15:0]   data_in_102_imag;
  reg        [15:0]   data_in_103_real;
  reg        [15:0]   data_in_103_imag;
  reg        [15:0]   data_in_104_real;
  reg        [15:0]   data_in_104_imag;
  reg        [15:0]   data_in_105_real;
  reg        [15:0]   data_in_105_imag;
  reg        [15:0]   data_in_106_real;
  reg        [15:0]   data_in_106_imag;
  reg        [15:0]   data_in_107_real;
  reg        [15:0]   data_in_107_imag;
  reg        [15:0]   data_in_108_real;
  reg        [15:0]   data_in_108_imag;
  reg        [15:0]   data_in_109_real;
  reg        [15:0]   data_in_109_imag;
  reg        [15:0]   data_in_110_real;
  reg        [15:0]   data_in_110_imag;
  reg        [15:0]   data_in_111_real;
  reg        [15:0]   data_in_111_imag;
  reg        [15:0]   data_in_112_real;
  reg        [15:0]   data_in_112_imag;
  reg        [15:0]   data_in_113_real;
  reg        [15:0]   data_in_113_imag;
  reg        [15:0]   data_in_114_real;
  reg        [15:0]   data_in_114_imag;
  reg        [15:0]   data_in_115_real;
  reg        [15:0]   data_in_115_imag;
  reg        [15:0]   data_in_116_real;
  reg        [15:0]   data_in_116_imag;
  reg        [15:0]   data_in_117_real;
  reg        [15:0]   data_in_117_imag;
  reg        [15:0]   data_in_118_real;
  reg        [15:0]   data_in_118_imag;
  reg        [15:0]   data_in_119_real;
  reg        [15:0]   data_in_119_imag;
  reg        [15:0]   data_in_120_real;
  reg        [15:0]   data_in_120_imag;
  reg        [15:0]   data_in_121_real;
  reg        [15:0]   data_in_121_imag;
  reg        [15:0]   data_in_122_real;
  reg        [15:0]   data_in_122_imag;
  reg        [15:0]   data_in_123_real;
  reg        [15:0]   data_in_123_imag;
  reg        [15:0]   data_in_124_real;
  reg        [15:0]   data_in_124_imag;
  reg        [15:0]   data_in_125_real;
  reg        [15:0]   data_in_125_imag;
  reg        [15:0]   data_in_126_real;
  reg        [15:0]   data_in_126_imag;
  reg        [15:0]   data_in_127_real;
  reg        [15:0]   data_in_127_imag;
  wire       [15:0]   twiddle_factor_table_0_real;
  wire       [15:0]   twiddle_factor_table_0_imag;
  wire       [15:0]   twiddle_factor_table_1_real;
  wire       [15:0]   twiddle_factor_table_1_imag;
  wire       [15:0]   twiddle_factor_table_2_real;
  wire       [15:0]   twiddle_factor_table_2_imag;
  wire       [15:0]   twiddle_factor_table_3_real;
  wire       [15:0]   twiddle_factor_table_3_imag;
  wire       [15:0]   twiddle_factor_table_4_real;
  wire       [15:0]   twiddle_factor_table_4_imag;
  wire       [15:0]   twiddle_factor_table_5_real;
  wire       [15:0]   twiddle_factor_table_5_imag;
  wire       [15:0]   twiddle_factor_table_6_real;
  wire       [15:0]   twiddle_factor_table_6_imag;
  wire       [15:0]   twiddle_factor_table_7_real;
  wire       [15:0]   twiddle_factor_table_7_imag;
  wire       [15:0]   twiddle_factor_table_8_real;
  wire       [15:0]   twiddle_factor_table_8_imag;
  wire       [15:0]   twiddle_factor_table_9_real;
  wire       [15:0]   twiddle_factor_table_9_imag;
  wire       [15:0]   twiddle_factor_table_10_real;
  wire       [15:0]   twiddle_factor_table_10_imag;
  wire       [15:0]   twiddle_factor_table_11_real;
  wire       [15:0]   twiddle_factor_table_11_imag;
  wire       [15:0]   twiddle_factor_table_12_real;
  wire       [15:0]   twiddle_factor_table_12_imag;
  wire       [15:0]   twiddle_factor_table_13_real;
  wire       [15:0]   twiddle_factor_table_13_imag;
  wire       [15:0]   twiddle_factor_table_14_real;
  wire       [15:0]   twiddle_factor_table_14_imag;
  wire       [15:0]   twiddle_factor_table_15_real;
  wire       [15:0]   twiddle_factor_table_15_imag;
  wire       [15:0]   twiddle_factor_table_16_real;
  wire       [15:0]   twiddle_factor_table_16_imag;
  wire       [15:0]   twiddle_factor_table_17_real;
  wire       [15:0]   twiddle_factor_table_17_imag;
  wire       [15:0]   twiddle_factor_table_18_real;
  wire       [15:0]   twiddle_factor_table_18_imag;
  wire       [15:0]   twiddle_factor_table_19_real;
  wire       [15:0]   twiddle_factor_table_19_imag;
  wire       [15:0]   twiddle_factor_table_20_real;
  wire       [15:0]   twiddle_factor_table_20_imag;
  wire       [15:0]   twiddle_factor_table_21_real;
  wire       [15:0]   twiddle_factor_table_21_imag;
  wire       [15:0]   twiddle_factor_table_22_real;
  wire       [15:0]   twiddle_factor_table_22_imag;
  wire       [15:0]   twiddle_factor_table_23_real;
  wire       [15:0]   twiddle_factor_table_23_imag;
  wire       [15:0]   twiddle_factor_table_24_real;
  wire       [15:0]   twiddle_factor_table_24_imag;
  wire       [15:0]   twiddle_factor_table_25_real;
  wire       [15:0]   twiddle_factor_table_25_imag;
  wire       [15:0]   twiddle_factor_table_26_real;
  wire       [15:0]   twiddle_factor_table_26_imag;
  wire       [15:0]   twiddle_factor_table_27_real;
  wire       [15:0]   twiddle_factor_table_27_imag;
  wire       [15:0]   twiddle_factor_table_28_real;
  wire       [15:0]   twiddle_factor_table_28_imag;
  wire       [15:0]   twiddle_factor_table_29_real;
  wire       [15:0]   twiddle_factor_table_29_imag;
  wire       [15:0]   twiddle_factor_table_30_real;
  wire       [15:0]   twiddle_factor_table_30_imag;
  wire       [15:0]   twiddle_factor_table_31_real;
  wire       [15:0]   twiddle_factor_table_31_imag;
  wire       [15:0]   twiddle_factor_table_32_real;
  wire       [15:0]   twiddle_factor_table_32_imag;
  wire       [15:0]   twiddle_factor_table_33_real;
  wire       [15:0]   twiddle_factor_table_33_imag;
  wire       [15:0]   twiddle_factor_table_34_real;
  wire       [15:0]   twiddle_factor_table_34_imag;
  wire       [15:0]   twiddle_factor_table_35_real;
  wire       [15:0]   twiddle_factor_table_35_imag;
  wire       [15:0]   twiddle_factor_table_36_real;
  wire       [15:0]   twiddle_factor_table_36_imag;
  wire       [15:0]   twiddle_factor_table_37_real;
  wire       [15:0]   twiddle_factor_table_37_imag;
  wire       [15:0]   twiddle_factor_table_38_real;
  wire       [15:0]   twiddle_factor_table_38_imag;
  wire       [15:0]   twiddle_factor_table_39_real;
  wire       [15:0]   twiddle_factor_table_39_imag;
  wire       [15:0]   twiddle_factor_table_40_real;
  wire       [15:0]   twiddle_factor_table_40_imag;
  wire       [15:0]   twiddle_factor_table_41_real;
  wire       [15:0]   twiddle_factor_table_41_imag;
  wire       [15:0]   twiddle_factor_table_42_real;
  wire       [15:0]   twiddle_factor_table_42_imag;
  wire       [15:0]   twiddle_factor_table_43_real;
  wire       [15:0]   twiddle_factor_table_43_imag;
  wire       [15:0]   twiddle_factor_table_44_real;
  wire       [15:0]   twiddle_factor_table_44_imag;
  wire       [15:0]   twiddle_factor_table_45_real;
  wire       [15:0]   twiddle_factor_table_45_imag;
  wire       [15:0]   twiddle_factor_table_46_real;
  wire       [15:0]   twiddle_factor_table_46_imag;
  wire       [15:0]   twiddle_factor_table_47_real;
  wire       [15:0]   twiddle_factor_table_47_imag;
  wire       [15:0]   twiddle_factor_table_48_real;
  wire       [15:0]   twiddle_factor_table_48_imag;
  wire       [15:0]   twiddle_factor_table_49_real;
  wire       [15:0]   twiddle_factor_table_49_imag;
  wire       [15:0]   twiddle_factor_table_50_real;
  wire       [15:0]   twiddle_factor_table_50_imag;
  wire       [15:0]   twiddle_factor_table_51_real;
  wire       [15:0]   twiddle_factor_table_51_imag;
  wire       [15:0]   twiddle_factor_table_52_real;
  wire       [15:0]   twiddle_factor_table_52_imag;
  wire       [15:0]   twiddle_factor_table_53_real;
  wire       [15:0]   twiddle_factor_table_53_imag;
  wire       [15:0]   twiddle_factor_table_54_real;
  wire       [15:0]   twiddle_factor_table_54_imag;
  wire       [15:0]   twiddle_factor_table_55_real;
  wire       [15:0]   twiddle_factor_table_55_imag;
  wire       [15:0]   twiddle_factor_table_56_real;
  wire       [15:0]   twiddle_factor_table_56_imag;
  wire       [15:0]   twiddle_factor_table_57_real;
  wire       [15:0]   twiddle_factor_table_57_imag;
  wire       [15:0]   twiddle_factor_table_58_real;
  wire       [15:0]   twiddle_factor_table_58_imag;
  wire       [15:0]   twiddle_factor_table_59_real;
  wire       [15:0]   twiddle_factor_table_59_imag;
  wire       [15:0]   twiddle_factor_table_60_real;
  wire       [15:0]   twiddle_factor_table_60_imag;
  wire       [15:0]   twiddle_factor_table_61_real;
  wire       [15:0]   twiddle_factor_table_61_imag;
  wire       [15:0]   twiddle_factor_table_62_real;
  wire       [15:0]   twiddle_factor_table_62_imag;
  wire       [15:0]   twiddle_factor_table_63_real;
  wire       [15:0]   twiddle_factor_table_63_imag;
  wire       [15:0]   twiddle_factor_table_64_real;
  wire       [15:0]   twiddle_factor_table_64_imag;
  wire       [15:0]   twiddle_factor_table_65_real;
  wire       [15:0]   twiddle_factor_table_65_imag;
  wire       [15:0]   twiddle_factor_table_66_real;
  wire       [15:0]   twiddle_factor_table_66_imag;
  wire       [15:0]   twiddle_factor_table_67_real;
  wire       [15:0]   twiddle_factor_table_67_imag;
  wire       [15:0]   twiddle_factor_table_68_real;
  wire       [15:0]   twiddle_factor_table_68_imag;
  wire       [15:0]   twiddle_factor_table_69_real;
  wire       [15:0]   twiddle_factor_table_69_imag;
  wire       [15:0]   twiddle_factor_table_70_real;
  wire       [15:0]   twiddle_factor_table_70_imag;
  wire       [15:0]   twiddle_factor_table_71_real;
  wire       [15:0]   twiddle_factor_table_71_imag;
  wire       [15:0]   twiddle_factor_table_72_real;
  wire       [15:0]   twiddle_factor_table_72_imag;
  wire       [15:0]   twiddle_factor_table_73_real;
  wire       [15:0]   twiddle_factor_table_73_imag;
  wire       [15:0]   twiddle_factor_table_74_real;
  wire       [15:0]   twiddle_factor_table_74_imag;
  wire       [15:0]   twiddle_factor_table_75_real;
  wire       [15:0]   twiddle_factor_table_75_imag;
  wire       [15:0]   twiddle_factor_table_76_real;
  wire       [15:0]   twiddle_factor_table_76_imag;
  wire       [15:0]   twiddle_factor_table_77_real;
  wire       [15:0]   twiddle_factor_table_77_imag;
  wire       [15:0]   twiddle_factor_table_78_real;
  wire       [15:0]   twiddle_factor_table_78_imag;
  wire       [15:0]   twiddle_factor_table_79_real;
  wire       [15:0]   twiddle_factor_table_79_imag;
  wire       [15:0]   twiddle_factor_table_80_real;
  wire       [15:0]   twiddle_factor_table_80_imag;
  wire       [15:0]   twiddle_factor_table_81_real;
  wire       [15:0]   twiddle_factor_table_81_imag;
  wire       [15:0]   twiddle_factor_table_82_real;
  wire       [15:0]   twiddle_factor_table_82_imag;
  wire       [15:0]   twiddle_factor_table_83_real;
  wire       [15:0]   twiddle_factor_table_83_imag;
  wire       [15:0]   twiddle_factor_table_84_real;
  wire       [15:0]   twiddle_factor_table_84_imag;
  wire       [15:0]   twiddle_factor_table_85_real;
  wire       [15:0]   twiddle_factor_table_85_imag;
  wire       [15:0]   twiddle_factor_table_86_real;
  wire       [15:0]   twiddle_factor_table_86_imag;
  wire       [15:0]   twiddle_factor_table_87_real;
  wire       [15:0]   twiddle_factor_table_87_imag;
  wire       [15:0]   twiddle_factor_table_88_real;
  wire       [15:0]   twiddle_factor_table_88_imag;
  wire       [15:0]   twiddle_factor_table_89_real;
  wire       [15:0]   twiddle_factor_table_89_imag;
  wire       [15:0]   twiddle_factor_table_90_real;
  wire       [15:0]   twiddle_factor_table_90_imag;
  wire       [15:0]   twiddle_factor_table_91_real;
  wire       [15:0]   twiddle_factor_table_91_imag;
  wire       [15:0]   twiddle_factor_table_92_real;
  wire       [15:0]   twiddle_factor_table_92_imag;
  wire       [15:0]   twiddle_factor_table_93_real;
  wire       [15:0]   twiddle_factor_table_93_imag;
  wire       [15:0]   twiddle_factor_table_94_real;
  wire       [15:0]   twiddle_factor_table_94_imag;
  wire       [15:0]   twiddle_factor_table_95_real;
  wire       [15:0]   twiddle_factor_table_95_imag;
  wire       [15:0]   twiddle_factor_table_96_real;
  wire       [15:0]   twiddle_factor_table_96_imag;
  wire       [15:0]   twiddle_factor_table_97_real;
  wire       [15:0]   twiddle_factor_table_97_imag;
  wire       [15:0]   twiddle_factor_table_98_real;
  wire       [15:0]   twiddle_factor_table_98_imag;
  wire       [15:0]   twiddle_factor_table_99_real;
  wire       [15:0]   twiddle_factor_table_99_imag;
  wire       [15:0]   twiddle_factor_table_100_real;
  wire       [15:0]   twiddle_factor_table_100_imag;
  wire       [15:0]   twiddle_factor_table_101_real;
  wire       [15:0]   twiddle_factor_table_101_imag;
  wire       [15:0]   twiddle_factor_table_102_real;
  wire       [15:0]   twiddle_factor_table_102_imag;
  wire       [15:0]   twiddle_factor_table_103_real;
  wire       [15:0]   twiddle_factor_table_103_imag;
  wire       [15:0]   twiddle_factor_table_104_real;
  wire       [15:0]   twiddle_factor_table_104_imag;
  wire       [15:0]   twiddle_factor_table_105_real;
  wire       [15:0]   twiddle_factor_table_105_imag;
  wire       [15:0]   twiddle_factor_table_106_real;
  wire       [15:0]   twiddle_factor_table_106_imag;
  wire       [15:0]   twiddle_factor_table_107_real;
  wire       [15:0]   twiddle_factor_table_107_imag;
  wire       [15:0]   twiddle_factor_table_108_real;
  wire       [15:0]   twiddle_factor_table_108_imag;
  wire       [15:0]   twiddle_factor_table_109_real;
  wire       [15:0]   twiddle_factor_table_109_imag;
  wire       [15:0]   twiddle_factor_table_110_real;
  wire       [15:0]   twiddle_factor_table_110_imag;
  wire       [15:0]   twiddle_factor_table_111_real;
  wire       [15:0]   twiddle_factor_table_111_imag;
  wire       [15:0]   twiddle_factor_table_112_real;
  wire       [15:0]   twiddle_factor_table_112_imag;
  wire       [15:0]   twiddle_factor_table_113_real;
  wire       [15:0]   twiddle_factor_table_113_imag;
  wire       [15:0]   twiddle_factor_table_114_real;
  wire       [15:0]   twiddle_factor_table_114_imag;
  wire       [15:0]   twiddle_factor_table_115_real;
  wire       [15:0]   twiddle_factor_table_115_imag;
  wire       [15:0]   twiddle_factor_table_116_real;
  wire       [15:0]   twiddle_factor_table_116_imag;
  wire       [15:0]   twiddle_factor_table_117_real;
  wire       [15:0]   twiddle_factor_table_117_imag;
  wire       [15:0]   twiddle_factor_table_118_real;
  wire       [15:0]   twiddle_factor_table_118_imag;
  wire       [15:0]   twiddle_factor_table_119_real;
  wire       [15:0]   twiddle_factor_table_119_imag;
  wire       [15:0]   twiddle_factor_table_120_real;
  wire       [15:0]   twiddle_factor_table_120_imag;
  wire       [15:0]   twiddle_factor_table_121_real;
  wire       [15:0]   twiddle_factor_table_121_imag;
  wire       [15:0]   twiddle_factor_table_122_real;
  wire       [15:0]   twiddle_factor_table_122_imag;
  wire       [15:0]   twiddle_factor_table_123_real;
  wire       [15:0]   twiddle_factor_table_123_imag;
  wire       [15:0]   twiddle_factor_table_124_real;
  wire       [15:0]   twiddle_factor_table_124_imag;
  wire       [15:0]   twiddle_factor_table_125_real;
  wire       [15:0]   twiddle_factor_table_125_imag;
  wire       [15:0]   twiddle_factor_table_126_real;
  wire       [15:0]   twiddle_factor_table_126_imag;
  wire       [15:0]   data_reorder_0_real;
  wire       [15:0]   data_reorder_0_imag;
  wire       [15:0]   data_reorder_1_real;
  wire       [15:0]   data_reorder_1_imag;
  wire       [15:0]   data_reorder_2_real;
  wire       [15:0]   data_reorder_2_imag;
  wire       [15:0]   data_reorder_3_real;
  wire       [15:0]   data_reorder_3_imag;
  wire       [15:0]   data_reorder_4_real;
  wire       [15:0]   data_reorder_4_imag;
  wire       [15:0]   data_reorder_5_real;
  wire       [15:0]   data_reorder_5_imag;
  wire       [15:0]   data_reorder_6_real;
  wire       [15:0]   data_reorder_6_imag;
  wire       [15:0]   data_reorder_7_real;
  wire       [15:0]   data_reorder_7_imag;
  wire       [15:0]   data_reorder_8_real;
  wire       [15:0]   data_reorder_8_imag;
  wire       [15:0]   data_reorder_9_real;
  wire       [15:0]   data_reorder_9_imag;
  wire       [15:0]   data_reorder_10_real;
  wire       [15:0]   data_reorder_10_imag;
  wire       [15:0]   data_reorder_11_real;
  wire       [15:0]   data_reorder_11_imag;
  wire       [15:0]   data_reorder_12_real;
  wire       [15:0]   data_reorder_12_imag;
  wire       [15:0]   data_reorder_13_real;
  wire       [15:0]   data_reorder_13_imag;
  wire       [15:0]   data_reorder_14_real;
  wire       [15:0]   data_reorder_14_imag;
  wire       [15:0]   data_reorder_15_real;
  wire       [15:0]   data_reorder_15_imag;
  wire       [15:0]   data_reorder_16_real;
  wire       [15:0]   data_reorder_16_imag;
  wire       [15:0]   data_reorder_17_real;
  wire       [15:0]   data_reorder_17_imag;
  wire       [15:0]   data_reorder_18_real;
  wire       [15:0]   data_reorder_18_imag;
  wire       [15:0]   data_reorder_19_real;
  wire       [15:0]   data_reorder_19_imag;
  wire       [15:0]   data_reorder_20_real;
  wire       [15:0]   data_reorder_20_imag;
  wire       [15:0]   data_reorder_21_real;
  wire       [15:0]   data_reorder_21_imag;
  wire       [15:0]   data_reorder_22_real;
  wire       [15:0]   data_reorder_22_imag;
  wire       [15:0]   data_reorder_23_real;
  wire       [15:0]   data_reorder_23_imag;
  wire       [15:0]   data_reorder_24_real;
  wire       [15:0]   data_reorder_24_imag;
  wire       [15:0]   data_reorder_25_real;
  wire       [15:0]   data_reorder_25_imag;
  wire       [15:0]   data_reorder_26_real;
  wire       [15:0]   data_reorder_26_imag;
  wire       [15:0]   data_reorder_27_real;
  wire       [15:0]   data_reorder_27_imag;
  wire       [15:0]   data_reorder_28_real;
  wire       [15:0]   data_reorder_28_imag;
  wire       [15:0]   data_reorder_29_real;
  wire       [15:0]   data_reorder_29_imag;
  wire       [15:0]   data_reorder_30_real;
  wire       [15:0]   data_reorder_30_imag;
  wire       [15:0]   data_reorder_31_real;
  wire       [15:0]   data_reorder_31_imag;
  wire       [15:0]   data_reorder_32_real;
  wire       [15:0]   data_reorder_32_imag;
  wire       [15:0]   data_reorder_33_real;
  wire       [15:0]   data_reorder_33_imag;
  wire       [15:0]   data_reorder_34_real;
  wire       [15:0]   data_reorder_34_imag;
  wire       [15:0]   data_reorder_35_real;
  wire       [15:0]   data_reorder_35_imag;
  wire       [15:0]   data_reorder_36_real;
  wire       [15:0]   data_reorder_36_imag;
  wire       [15:0]   data_reorder_37_real;
  wire       [15:0]   data_reorder_37_imag;
  wire       [15:0]   data_reorder_38_real;
  wire       [15:0]   data_reorder_38_imag;
  wire       [15:0]   data_reorder_39_real;
  wire       [15:0]   data_reorder_39_imag;
  wire       [15:0]   data_reorder_40_real;
  wire       [15:0]   data_reorder_40_imag;
  wire       [15:0]   data_reorder_41_real;
  wire       [15:0]   data_reorder_41_imag;
  wire       [15:0]   data_reorder_42_real;
  wire       [15:0]   data_reorder_42_imag;
  wire       [15:0]   data_reorder_43_real;
  wire       [15:0]   data_reorder_43_imag;
  wire       [15:0]   data_reorder_44_real;
  wire       [15:0]   data_reorder_44_imag;
  wire       [15:0]   data_reorder_45_real;
  wire       [15:0]   data_reorder_45_imag;
  wire       [15:0]   data_reorder_46_real;
  wire       [15:0]   data_reorder_46_imag;
  wire       [15:0]   data_reorder_47_real;
  wire       [15:0]   data_reorder_47_imag;
  wire       [15:0]   data_reorder_48_real;
  wire       [15:0]   data_reorder_48_imag;
  wire       [15:0]   data_reorder_49_real;
  wire       [15:0]   data_reorder_49_imag;
  wire       [15:0]   data_reorder_50_real;
  wire       [15:0]   data_reorder_50_imag;
  wire       [15:0]   data_reorder_51_real;
  wire       [15:0]   data_reorder_51_imag;
  wire       [15:0]   data_reorder_52_real;
  wire       [15:0]   data_reorder_52_imag;
  wire       [15:0]   data_reorder_53_real;
  wire       [15:0]   data_reorder_53_imag;
  wire       [15:0]   data_reorder_54_real;
  wire       [15:0]   data_reorder_54_imag;
  wire       [15:0]   data_reorder_55_real;
  wire       [15:0]   data_reorder_55_imag;
  wire       [15:0]   data_reorder_56_real;
  wire       [15:0]   data_reorder_56_imag;
  wire       [15:0]   data_reorder_57_real;
  wire       [15:0]   data_reorder_57_imag;
  wire       [15:0]   data_reorder_58_real;
  wire       [15:0]   data_reorder_58_imag;
  wire       [15:0]   data_reorder_59_real;
  wire       [15:0]   data_reorder_59_imag;
  wire       [15:0]   data_reorder_60_real;
  wire       [15:0]   data_reorder_60_imag;
  wire       [15:0]   data_reorder_61_real;
  wire       [15:0]   data_reorder_61_imag;
  wire       [15:0]   data_reorder_62_real;
  wire       [15:0]   data_reorder_62_imag;
  wire       [15:0]   data_reorder_63_real;
  wire       [15:0]   data_reorder_63_imag;
  wire       [15:0]   data_reorder_64_real;
  wire       [15:0]   data_reorder_64_imag;
  wire       [15:0]   data_reorder_65_real;
  wire       [15:0]   data_reorder_65_imag;
  wire       [15:0]   data_reorder_66_real;
  wire       [15:0]   data_reorder_66_imag;
  wire       [15:0]   data_reorder_67_real;
  wire       [15:0]   data_reorder_67_imag;
  wire       [15:0]   data_reorder_68_real;
  wire       [15:0]   data_reorder_68_imag;
  wire       [15:0]   data_reorder_69_real;
  wire       [15:0]   data_reorder_69_imag;
  wire       [15:0]   data_reorder_70_real;
  wire       [15:0]   data_reorder_70_imag;
  wire       [15:0]   data_reorder_71_real;
  wire       [15:0]   data_reorder_71_imag;
  wire       [15:0]   data_reorder_72_real;
  wire       [15:0]   data_reorder_72_imag;
  wire       [15:0]   data_reorder_73_real;
  wire       [15:0]   data_reorder_73_imag;
  wire       [15:0]   data_reorder_74_real;
  wire       [15:0]   data_reorder_74_imag;
  wire       [15:0]   data_reorder_75_real;
  wire       [15:0]   data_reorder_75_imag;
  wire       [15:0]   data_reorder_76_real;
  wire       [15:0]   data_reorder_76_imag;
  wire       [15:0]   data_reorder_77_real;
  wire       [15:0]   data_reorder_77_imag;
  wire       [15:0]   data_reorder_78_real;
  wire       [15:0]   data_reorder_78_imag;
  wire       [15:0]   data_reorder_79_real;
  wire       [15:0]   data_reorder_79_imag;
  wire       [15:0]   data_reorder_80_real;
  wire       [15:0]   data_reorder_80_imag;
  wire       [15:0]   data_reorder_81_real;
  wire       [15:0]   data_reorder_81_imag;
  wire       [15:0]   data_reorder_82_real;
  wire       [15:0]   data_reorder_82_imag;
  wire       [15:0]   data_reorder_83_real;
  wire       [15:0]   data_reorder_83_imag;
  wire       [15:0]   data_reorder_84_real;
  wire       [15:0]   data_reorder_84_imag;
  wire       [15:0]   data_reorder_85_real;
  wire       [15:0]   data_reorder_85_imag;
  wire       [15:0]   data_reorder_86_real;
  wire       [15:0]   data_reorder_86_imag;
  wire       [15:0]   data_reorder_87_real;
  wire       [15:0]   data_reorder_87_imag;
  wire       [15:0]   data_reorder_88_real;
  wire       [15:0]   data_reorder_88_imag;
  wire       [15:0]   data_reorder_89_real;
  wire       [15:0]   data_reorder_89_imag;
  wire       [15:0]   data_reorder_90_real;
  wire       [15:0]   data_reorder_90_imag;
  wire       [15:0]   data_reorder_91_real;
  wire       [15:0]   data_reorder_91_imag;
  wire       [15:0]   data_reorder_92_real;
  wire       [15:0]   data_reorder_92_imag;
  wire       [15:0]   data_reorder_93_real;
  wire       [15:0]   data_reorder_93_imag;
  wire       [15:0]   data_reorder_94_real;
  wire       [15:0]   data_reorder_94_imag;
  wire       [15:0]   data_reorder_95_real;
  wire       [15:0]   data_reorder_95_imag;
  wire       [15:0]   data_reorder_96_real;
  wire       [15:0]   data_reorder_96_imag;
  wire       [15:0]   data_reorder_97_real;
  wire       [15:0]   data_reorder_97_imag;
  wire       [15:0]   data_reorder_98_real;
  wire       [15:0]   data_reorder_98_imag;
  wire       [15:0]   data_reorder_99_real;
  wire       [15:0]   data_reorder_99_imag;
  wire       [15:0]   data_reorder_100_real;
  wire       [15:0]   data_reorder_100_imag;
  wire       [15:0]   data_reorder_101_real;
  wire       [15:0]   data_reorder_101_imag;
  wire       [15:0]   data_reorder_102_real;
  wire       [15:0]   data_reorder_102_imag;
  wire       [15:0]   data_reorder_103_real;
  wire       [15:0]   data_reorder_103_imag;
  wire       [15:0]   data_reorder_104_real;
  wire       [15:0]   data_reorder_104_imag;
  wire       [15:0]   data_reorder_105_real;
  wire       [15:0]   data_reorder_105_imag;
  wire       [15:0]   data_reorder_106_real;
  wire       [15:0]   data_reorder_106_imag;
  wire       [15:0]   data_reorder_107_real;
  wire       [15:0]   data_reorder_107_imag;
  wire       [15:0]   data_reorder_108_real;
  wire       [15:0]   data_reorder_108_imag;
  wire       [15:0]   data_reorder_109_real;
  wire       [15:0]   data_reorder_109_imag;
  wire       [15:0]   data_reorder_110_real;
  wire       [15:0]   data_reorder_110_imag;
  wire       [15:0]   data_reorder_111_real;
  wire       [15:0]   data_reorder_111_imag;
  wire       [15:0]   data_reorder_112_real;
  wire       [15:0]   data_reorder_112_imag;
  wire       [15:0]   data_reorder_113_real;
  wire       [15:0]   data_reorder_113_imag;
  wire       [15:0]   data_reorder_114_real;
  wire       [15:0]   data_reorder_114_imag;
  wire       [15:0]   data_reorder_115_real;
  wire       [15:0]   data_reorder_115_imag;
  wire       [15:0]   data_reorder_116_real;
  wire       [15:0]   data_reorder_116_imag;
  wire       [15:0]   data_reorder_117_real;
  wire       [15:0]   data_reorder_117_imag;
  wire       [15:0]   data_reorder_118_real;
  wire       [15:0]   data_reorder_118_imag;
  wire       [15:0]   data_reorder_119_real;
  wire       [15:0]   data_reorder_119_imag;
  wire       [15:0]   data_reorder_120_real;
  wire       [15:0]   data_reorder_120_imag;
  wire       [15:0]   data_reorder_121_real;
  wire       [15:0]   data_reorder_121_imag;
  wire       [15:0]   data_reorder_122_real;
  wire       [15:0]   data_reorder_122_imag;
  wire       [15:0]   data_reorder_123_real;
  wire       [15:0]   data_reorder_123_imag;
  wire       [15:0]   data_reorder_124_real;
  wire       [15:0]   data_reorder_124_imag;
  wire       [15:0]   data_reorder_125_real;
  wire       [15:0]   data_reorder_125_imag;
  wire       [15:0]   data_reorder_126_real;
  wire       [15:0]   data_reorder_126_imag;
  wire       [15:0]   data_reorder_127_real;
  wire       [15:0]   data_reorder_127_imag;
  reg        [15:0]   _zz_1;
  reg        [15:0]   _zz_2;
  reg        [15:0]   _zz_3;
  reg        [15:0]   _zz_4;
  reg        [15:0]   _zz_5;
  reg        [15:0]   _zz_6;
  reg        [15:0]   _zz_7;
  reg        [15:0]   _zz_8;
  reg        [15:0]   _zz_9;
  reg        [15:0]   _zz_10;
  reg        [15:0]   _zz_11;
  reg        [15:0]   _zz_12;
  reg        [15:0]   _zz_13;
  reg        [15:0]   _zz_14;
  reg        [15:0]   _zz_15;
  reg        [15:0]   _zz_16;
  reg        [15:0]   _zz_17;
  reg        [15:0]   _zz_18;
  reg        [15:0]   _zz_19;
  reg        [15:0]   _zz_20;
  reg        [15:0]   _zz_21;
  reg        [15:0]   _zz_22;
  reg        [15:0]   _zz_23;
  reg        [15:0]   _zz_24;
  reg        [15:0]   _zz_25;
  reg        [15:0]   _zz_26;
  reg        [15:0]   _zz_27;
  reg        [15:0]   _zz_28;
  reg        [15:0]   _zz_29;
  reg        [15:0]   _zz_30;
  reg        [15:0]   _zz_31;
  reg        [15:0]   _zz_32;
  reg        [15:0]   _zz_33;
  reg        [15:0]   _zz_34;
  reg        [15:0]   _zz_35;
  reg        [15:0]   _zz_36;
  reg        [15:0]   _zz_37;
  reg        [15:0]   _zz_38;
  reg        [15:0]   _zz_39;
  reg        [15:0]   _zz_40;
  reg        [15:0]   _zz_41;
  reg        [15:0]   _zz_42;
  reg        [15:0]   _zz_43;
  reg        [15:0]   _zz_44;
  reg        [15:0]   _zz_45;
  reg        [15:0]   _zz_46;
  reg        [15:0]   _zz_47;
  reg        [15:0]   _zz_48;
  reg        [15:0]   _zz_49;
  reg        [15:0]   _zz_50;
  reg        [15:0]   _zz_51;
  reg        [15:0]   _zz_52;
  reg        [15:0]   _zz_53;
  reg        [15:0]   _zz_54;
  reg        [15:0]   _zz_55;
  reg        [15:0]   _zz_56;
  reg        [15:0]   _zz_57;
  reg        [15:0]   _zz_58;
  reg        [15:0]   _zz_59;
  reg        [15:0]   _zz_60;
  reg        [15:0]   _zz_61;
  reg        [15:0]   _zz_62;
  reg        [15:0]   _zz_63;
  reg        [15:0]   _zz_64;
  reg        [15:0]   _zz_65;
  reg        [15:0]   _zz_66;
  reg        [15:0]   _zz_67;
  reg        [15:0]   _zz_68;
  reg        [15:0]   _zz_69;
  reg        [15:0]   _zz_70;
  reg        [15:0]   _zz_71;
  reg        [15:0]   _zz_72;
  reg        [15:0]   _zz_73;
  reg        [15:0]   _zz_74;
  reg        [15:0]   _zz_75;
  reg        [15:0]   _zz_76;
  reg        [15:0]   _zz_77;
  reg        [15:0]   _zz_78;
  reg        [15:0]   _zz_79;
  reg        [15:0]   _zz_80;
  reg        [15:0]   _zz_81;
  reg        [15:0]   _zz_82;
  reg        [15:0]   _zz_83;
  reg        [15:0]   _zz_84;
  reg        [15:0]   _zz_85;
  reg        [15:0]   _zz_86;
  reg        [15:0]   _zz_87;
  reg        [15:0]   _zz_88;
  reg        [15:0]   _zz_89;
  reg        [15:0]   _zz_90;
  reg        [15:0]   _zz_91;
  reg        [15:0]   _zz_92;
  reg        [15:0]   _zz_93;
  reg        [15:0]   _zz_94;
  reg        [15:0]   _zz_95;
  reg        [15:0]   _zz_96;
  reg        [15:0]   _zz_97;
  reg        [15:0]   _zz_98;
  reg        [15:0]   _zz_99;
  reg        [15:0]   _zz_100;
  reg        [15:0]   _zz_101;
  reg        [15:0]   _zz_102;
  reg        [15:0]   _zz_103;
  reg        [15:0]   _zz_104;
  reg        [15:0]   _zz_105;
  reg        [15:0]   _zz_106;
  reg        [15:0]   _zz_107;
  reg        [15:0]   _zz_108;
  reg        [15:0]   _zz_109;
  reg        [15:0]   _zz_110;
  reg        [15:0]   _zz_111;
  reg        [15:0]   _zz_112;
  reg        [15:0]   _zz_113;
  reg        [15:0]   _zz_114;
  reg        [15:0]   _zz_115;
  reg        [15:0]   _zz_116;
  reg        [15:0]   _zz_117;
  reg        [15:0]   _zz_118;
  reg        [15:0]   _zz_119;
  reg        [15:0]   _zz_120;
  reg        [15:0]   _zz_121;
  reg        [15:0]   _zz_122;
  reg        [15:0]   _zz_123;
  reg        [15:0]   _zz_124;
  reg        [15:0]   _zz_125;
  reg        [15:0]   _zz_126;
  reg        [15:0]   _zz_127;
  reg        [15:0]   _zz_128;
  reg        [15:0]   _zz_129;
  reg        [15:0]   _zz_130;
  reg        [15:0]   _zz_131;
  reg        [15:0]   _zz_132;
  reg        [15:0]   _zz_133;
  reg        [15:0]   _zz_134;
  reg        [15:0]   _zz_135;
  reg        [15:0]   _zz_136;
  reg        [15:0]   _zz_137;
  reg        [15:0]   _zz_138;
  reg        [15:0]   _zz_139;
  reg        [15:0]   _zz_140;
  reg        [15:0]   _zz_141;
  reg        [15:0]   _zz_142;
  reg        [15:0]   _zz_143;
  reg        [15:0]   _zz_144;
  reg        [15:0]   _zz_145;
  reg        [15:0]   _zz_146;
  reg        [15:0]   _zz_147;
  reg        [15:0]   _zz_148;
  reg        [15:0]   _zz_149;
  reg        [15:0]   _zz_150;
  reg        [15:0]   _zz_151;
  reg        [15:0]   _zz_152;
  reg        [15:0]   _zz_153;
  reg        [15:0]   _zz_154;
  reg        [15:0]   _zz_155;
  reg        [15:0]   _zz_156;
  reg        [15:0]   _zz_157;
  reg        [15:0]   _zz_158;
  reg        [15:0]   _zz_159;
  reg        [15:0]   _zz_160;
  reg        [15:0]   _zz_161;
  reg        [15:0]   _zz_162;
  reg        [15:0]   _zz_163;
  reg        [15:0]   _zz_164;
  reg        [15:0]   _zz_165;
  reg        [15:0]   _zz_166;
  reg        [15:0]   _zz_167;
  reg        [15:0]   _zz_168;
  reg        [15:0]   _zz_169;
  reg        [15:0]   _zz_170;
  reg        [15:0]   _zz_171;
  reg        [15:0]   _zz_172;
  reg        [15:0]   _zz_173;
  reg        [15:0]   _zz_174;
  reg        [15:0]   _zz_175;
  reg        [15:0]   _zz_176;
  reg        [15:0]   _zz_177;
  reg        [15:0]   _zz_178;
  reg        [15:0]   _zz_179;
  reg        [15:0]   _zz_180;
  reg        [15:0]   _zz_181;
  reg        [15:0]   _zz_182;
  reg        [15:0]   _zz_183;
  reg        [15:0]   _zz_184;
  reg        [15:0]   _zz_185;
  reg        [15:0]   _zz_186;
  reg        [15:0]   _zz_187;
  reg        [15:0]   _zz_188;
  reg        [15:0]   _zz_189;
  reg        [15:0]   _zz_190;
  reg        [15:0]   _zz_191;
  reg        [15:0]   _zz_192;
  reg        [15:0]   _zz_193;
  reg        [15:0]   _zz_194;
  reg        [15:0]   _zz_195;
  reg        [15:0]   _zz_196;
  reg        [15:0]   _zz_197;
  reg        [15:0]   _zz_198;
  reg        [15:0]   _zz_199;
  reg        [15:0]   _zz_200;
  reg        [15:0]   _zz_201;
  reg        [15:0]   _zz_202;
  reg        [15:0]   _zz_203;
  reg        [15:0]   _zz_204;
  reg        [15:0]   _zz_205;
  reg        [15:0]   _zz_206;
  reg        [15:0]   _zz_207;
  reg        [15:0]   _zz_208;
  reg        [15:0]   _zz_209;
  reg        [15:0]   _zz_210;
  reg        [15:0]   _zz_211;
  reg        [15:0]   _zz_212;
  reg        [15:0]   _zz_213;
  reg        [15:0]   _zz_214;
  reg        [15:0]   _zz_215;
  reg        [15:0]   _zz_216;
  reg        [15:0]   _zz_217;
  reg        [15:0]   _zz_218;
  reg        [15:0]   _zz_219;
  reg        [15:0]   _zz_220;
  reg        [15:0]   _zz_221;
  reg        [15:0]   _zz_222;
  reg        [15:0]   _zz_223;
  reg        [15:0]   _zz_224;
  reg        [15:0]   _zz_225;
  reg        [15:0]   _zz_226;
  reg        [15:0]   _zz_227;
  reg        [15:0]   _zz_228;
  reg        [15:0]   _zz_229;
  reg        [15:0]   _zz_230;
  reg        [15:0]   _zz_231;
  reg        [15:0]   _zz_232;
  reg        [15:0]   _zz_233;
  reg        [15:0]   _zz_234;
  reg        [15:0]   _zz_235;
  reg        [15:0]   _zz_236;
  reg        [15:0]   _zz_237;
  reg        [15:0]   _zz_238;
  reg        [15:0]   _zz_239;
  reg        [15:0]   _zz_240;
  reg        [15:0]   _zz_241;
  reg        [15:0]   _zz_242;
  reg        [15:0]   _zz_243;
  reg        [15:0]   _zz_244;
  reg        [15:0]   _zz_245;
  reg        [15:0]   _zz_246;
  reg        [15:0]   _zz_247;
  reg        [15:0]   _zz_248;
  reg        [15:0]   _zz_249;
  reg        [15:0]   _zz_250;
  reg        [15:0]   _zz_251;
  reg        [15:0]   _zz_252;
  reg        [15:0]   _zz_253;
  reg        [15:0]   _zz_254;
  reg        [15:0]   _zz_255;
  reg        [15:0]   _zz_256;
  reg        [15:0]   _zz_257;
  reg        [15:0]   _zz_258;
  reg        [15:0]   _zz_259;
  reg        [15:0]   _zz_260;
  reg        [15:0]   _zz_261;
  reg        [15:0]   _zz_262;
  reg        [15:0]   _zz_263;
  reg        [15:0]   _zz_264;
  reg        [15:0]   _zz_265;
  reg        [15:0]   _zz_266;
  reg        [15:0]   _zz_267;
  reg        [15:0]   _zz_268;
  reg        [15:0]   _zz_269;
  reg        [15:0]   _zz_270;
  reg        [15:0]   _zz_271;
  reg        [15:0]   _zz_272;
  reg        [15:0]   _zz_273;
  reg        [15:0]   _zz_274;
  reg        [15:0]   _zz_275;
  reg        [15:0]   _zz_276;
  reg        [15:0]   _zz_277;
  reg        [15:0]   _zz_278;
  reg        [15:0]   _zz_279;
  reg        [15:0]   _zz_280;
  reg        [15:0]   _zz_281;
  reg        [15:0]   _zz_282;
  reg        [15:0]   _zz_283;
  reg        [15:0]   _zz_284;
  reg        [15:0]   _zz_285;
  reg        [15:0]   _zz_286;
  reg        [15:0]   _zz_287;
  reg        [15:0]   _zz_288;
  reg        [15:0]   _zz_289;
  reg        [15:0]   _zz_290;
  reg        [15:0]   _zz_291;
  reg        [15:0]   _zz_292;
  reg        [15:0]   _zz_293;
  reg        [15:0]   _zz_294;
  reg        [15:0]   _zz_295;
  reg        [15:0]   _zz_296;
  reg        [15:0]   _zz_297;
  reg        [15:0]   _zz_298;
  reg        [15:0]   _zz_299;
  reg        [15:0]   _zz_300;
  reg        [15:0]   _zz_301;
  reg        [15:0]   _zz_302;
  reg        [15:0]   _zz_303;
  reg        [15:0]   _zz_304;
  reg        [15:0]   _zz_305;
  reg        [15:0]   _zz_306;
  reg        [15:0]   _zz_307;
  reg        [15:0]   _zz_308;
  reg        [15:0]   _zz_309;
  reg        [15:0]   _zz_310;
  reg        [15:0]   _zz_311;
  reg        [15:0]   _zz_312;
  reg        [15:0]   _zz_313;
  reg        [15:0]   _zz_314;
  reg        [15:0]   _zz_315;
  reg        [15:0]   _zz_316;
  reg        [15:0]   _zz_317;
  reg        [15:0]   _zz_318;
  reg        [15:0]   _zz_319;
  reg        [15:0]   _zz_320;
  reg        [15:0]   _zz_321;
  reg        [15:0]   _zz_322;
  reg        [15:0]   _zz_323;
  reg        [15:0]   _zz_324;
  reg        [15:0]   _zz_325;
  reg        [15:0]   _zz_326;
  reg        [15:0]   _zz_327;
  reg        [15:0]   _zz_328;
  reg        [15:0]   _zz_329;
  reg        [15:0]   _zz_330;
  reg        [15:0]   _zz_331;
  reg        [15:0]   _zz_332;
  reg        [15:0]   _zz_333;
  reg        [15:0]   _zz_334;
  reg        [15:0]   _zz_335;
  reg        [15:0]   _zz_336;
  reg        [15:0]   _zz_337;
  reg        [15:0]   _zz_338;
  reg        [15:0]   _zz_339;
  reg        [15:0]   _zz_340;
  reg        [15:0]   _zz_341;
  reg        [15:0]   _zz_342;
  reg        [15:0]   _zz_343;
  reg        [15:0]   _zz_344;
  reg        [15:0]   _zz_345;
  reg        [15:0]   _zz_346;
  reg        [15:0]   _zz_347;
  reg        [15:0]   _zz_348;
  reg        [15:0]   _zz_349;
  reg        [15:0]   _zz_350;
  reg        [15:0]   _zz_351;
  reg        [15:0]   _zz_352;
  reg        [15:0]   _zz_353;
  reg        [15:0]   _zz_354;
  reg        [15:0]   _zz_355;
  reg        [15:0]   _zz_356;
  reg        [15:0]   _zz_357;
  reg        [15:0]   _zz_358;
  reg        [15:0]   _zz_359;
  reg        [15:0]   _zz_360;
  reg        [15:0]   _zz_361;
  reg        [15:0]   _zz_362;
  reg        [15:0]   _zz_363;
  reg        [15:0]   _zz_364;
  reg        [15:0]   _zz_365;
  reg        [15:0]   _zz_366;
  reg        [15:0]   _zz_367;
  reg        [15:0]   _zz_368;
  reg        [15:0]   _zz_369;
  reg        [15:0]   _zz_370;
  reg        [15:0]   _zz_371;
  reg        [15:0]   _zz_372;
  reg        [15:0]   _zz_373;
  reg        [15:0]   _zz_374;
  reg        [15:0]   _zz_375;
  reg        [15:0]   _zz_376;
  reg        [15:0]   _zz_377;
  reg        [15:0]   _zz_378;
  reg        [15:0]   _zz_379;
  reg        [15:0]   _zz_380;
  reg        [15:0]   _zz_381;
  reg        [15:0]   _zz_382;
  reg        [15:0]   _zz_383;
  reg        [15:0]   _zz_384;
  reg        [15:0]   _zz_385;
  reg        [15:0]   _zz_386;
  reg        [15:0]   _zz_387;
  reg        [15:0]   _zz_388;
  reg        [15:0]   _zz_389;
  reg        [15:0]   _zz_390;
  reg        [15:0]   _zz_391;
  reg        [15:0]   _zz_392;
  reg        [15:0]   _zz_393;
  reg        [15:0]   _zz_394;
  reg        [15:0]   _zz_395;
  reg        [15:0]   _zz_396;
  reg        [15:0]   _zz_397;
  reg        [15:0]   _zz_398;
  reg        [15:0]   _zz_399;
  reg        [15:0]   _zz_400;
  reg        [15:0]   _zz_401;
  reg        [15:0]   _zz_402;
  reg        [15:0]   _zz_403;
  reg        [15:0]   _zz_404;
  reg        [15:0]   _zz_405;
  reg        [15:0]   _zz_406;
  reg        [15:0]   _zz_407;
  reg        [15:0]   _zz_408;
  reg        [15:0]   _zz_409;
  reg        [15:0]   _zz_410;
  reg        [15:0]   _zz_411;
  reg        [15:0]   _zz_412;
  reg        [15:0]   _zz_413;
  reg        [15:0]   _zz_414;
  reg        [15:0]   _zz_415;
  reg        [15:0]   _zz_416;
  reg        [15:0]   _zz_417;
  reg        [15:0]   _zz_418;
  reg        [15:0]   _zz_419;
  reg        [15:0]   _zz_420;
  reg        [15:0]   _zz_421;
  reg        [15:0]   _zz_422;
  reg        [15:0]   _zz_423;
  reg        [15:0]   _zz_424;
  reg        [15:0]   _zz_425;
  reg        [15:0]   _zz_426;
  reg        [15:0]   _zz_427;
  reg        [15:0]   _zz_428;
  reg        [15:0]   _zz_429;
  reg        [15:0]   _zz_430;
  reg        [15:0]   _zz_431;
  reg        [15:0]   _zz_432;
  reg        [15:0]   _zz_433;
  reg        [15:0]   _zz_434;
  reg        [15:0]   _zz_435;
  reg        [15:0]   _zz_436;
  reg        [15:0]   _zz_437;
  reg        [15:0]   _zz_438;
  reg        [15:0]   _zz_439;
  reg        [15:0]   _zz_440;
  reg        [15:0]   _zz_441;
  reg        [15:0]   _zz_442;
  reg        [15:0]   _zz_443;
  reg        [15:0]   _zz_444;
  reg        [15:0]   _zz_445;
  reg        [15:0]   _zz_446;
  reg        [15:0]   _zz_447;
  reg        [15:0]   _zz_448;
  reg        [15:0]   _zz_449;
  reg        [15:0]   _zz_450;
  reg        [15:0]   _zz_451;
  reg        [15:0]   _zz_452;
  reg        [15:0]   _zz_453;
  reg        [15:0]   _zz_454;
  reg        [15:0]   _zz_455;
  reg        [15:0]   _zz_456;
  reg        [15:0]   _zz_457;
  reg        [15:0]   _zz_458;
  reg        [15:0]   _zz_459;
  reg        [15:0]   _zz_460;
  reg        [15:0]   _zz_461;
  reg        [15:0]   _zz_462;
  reg        [15:0]   _zz_463;
  reg        [15:0]   _zz_464;
  reg        [15:0]   _zz_465;
  reg        [15:0]   _zz_466;
  reg        [15:0]   _zz_467;
  reg        [15:0]   _zz_468;
  reg        [15:0]   _zz_469;
  reg        [15:0]   _zz_470;
  reg        [15:0]   _zz_471;
  reg        [15:0]   _zz_472;
  reg        [15:0]   _zz_473;
  reg        [15:0]   _zz_474;
  reg        [15:0]   _zz_475;
  reg        [15:0]   _zz_476;
  reg        [15:0]   _zz_477;
  reg        [15:0]   _zz_478;
  reg        [15:0]   _zz_479;
  reg        [15:0]   _zz_480;
  reg        [15:0]   _zz_481;
  reg        [15:0]   _zz_482;
  reg        [15:0]   _zz_483;
  reg        [15:0]   _zz_484;
  reg        [15:0]   _zz_485;
  reg        [15:0]   _zz_486;
  reg        [15:0]   _zz_487;
  reg        [15:0]   _zz_488;
  reg        [15:0]   _zz_489;
  reg        [15:0]   _zz_490;
  reg        [15:0]   _zz_491;
  reg        [15:0]   _zz_492;
  reg        [15:0]   _zz_493;
  reg        [15:0]   _zz_494;
  reg        [15:0]   _zz_495;
  reg        [15:0]   _zz_496;
  reg        [15:0]   _zz_497;
  reg        [15:0]   _zz_498;
  reg        [15:0]   _zz_499;
  reg        [15:0]   _zz_500;
  reg        [15:0]   _zz_501;
  reg        [15:0]   _zz_502;
  reg        [15:0]   _zz_503;
  reg        [15:0]   _zz_504;
  reg        [15:0]   _zz_505;
  reg        [15:0]   _zz_506;
  reg        [15:0]   _zz_507;
  reg        [15:0]   _zz_508;
  reg        [15:0]   _zz_509;
  reg        [15:0]   _zz_510;
  reg        [15:0]   _zz_511;
  reg        [15:0]   _zz_512;
  reg        [15:0]   _zz_513;
  reg        [15:0]   _zz_514;
  reg        [15:0]   _zz_515;
  reg        [15:0]   _zz_516;
  reg        [15:0]   _zz_517;
  reg        [15:0]   _zz_518;
  reg        [15:0]   _zz_519;
  reg        [15:0]   _zz_520;
  reg        [15:0]   _zz_521;
  reg        [15:0]   _zz_522;
  reg        [15:0]   _zz_523;
  reg        [15:0]   _zz_524;
  reg        [15:0]   _zz_525;
  reg        [15:0]   _zz_526;
  reg        [15:0]   _zz_527;
  reg        [15:0]   _zz_528;
  reg        [15:0]   _zz_529;
  reg        [15:0]   _zz_530;
  reg        [15:0]   _zz_531;
  reg        [15:0]   _zz_532;
  reg        [15:0]   _zz_533;
  reg        [15:0]   _zz_534;
  reg        [15:0]   _zz_535;
  reg        [15:0]   _zz_536;
  reg        [15:0]   _zz_537;
  reg        [15:0]   _zz_538;
  reg        [15:0]   _zz_539;
  reg        [15:0]   _zz_540;
  reg        [15:0]   _zz_541;
  reg        [15:0]   _zz_542;
  reg        [15:0]   _zz_543;
  reg        [15:0]   _zz_544;
  reg        [15:0]   _zz_545;
  reg        [15:0]   _zz_546;
  reg        [15:0]   _zz_547;
  reg        [15:0]   _zz_548;
  reg        [15:0]   _zz_549;
  reg        [15:0]   _zz_550;
  reg        [15:0]   _zz_551;
  reg        [15:0]   _zz_552;
  reg        [15:0]   _zz_553;
  reg        [15:0]   _zz_554;
  reg        [15:0]   _zz_555;
  reg        [15:0]   _zz_556;
  reg        [15:0]   _zz_557;
  reg        [15:0]   _zz_558;
  reg        [15:0]   _zz_559;
  reg        [15:0]   _zz_560;
  reg        [15:0]   _zz_561;
  reg        [15:0]   _zz_562;
  reg        [15:0]   _zz_563;
  reg        [15:0]   _zz_564;
  reg        [15:0]   _zz_565;
  reg        [15:0]   _zz_566;
  reg        [15:0]   _zz_567;
  reg        [15:0]   _zz_568;
  reg        [15:0]   _zz_569;
  reg        [15:0]   _zz_570;
  reg        [15:0]   _zz_571;
  reg        [15:0]   _zz_572;
  reg        [15:0]   _zz_573;
  reg        [15:0]   _zz_574;
  reg        [15:0]   _zz_575;
  reg        [15:0]   _zz_576;
  reg        [15:0]   _zz_577;
  reg        [15:0]   _zz_578;
  reg        [15:0]   _zz_579;
  reg        [15:0]   _zz_580;
  reg        [15:0]   _zz_581;
  reg        [15:0]   _zz_582;
  reg        [15:0]   _zz_583;
  reg        [15:0]   _zz_584;
  reg        [15:0]   _zz_585;
  reg        [15:0]   _zz_586;
  reg        [15:0]   _zz_587;
  reg        [15:0]   _zz_588;
  reg        [15:0]   _zz_589;
  reg        [15:0]   _zz_590;
  reg        [15:0]   _zz_591;
  reg        [15:0]   _zz_592;
  reg        [15:0]   _zz_593;
  reg        [15:0]   _zz_594;
  reg        [15:0]   _zz_595;
  reg        [15:0]   _zz_596;
  reg        [15:0]   _zz_597;
  reg        [15:0]   _zz_598;
  reg        [15:0]   _zz_599;
  reg        [15:0]   _zz_600;
  reg        [15:0]   _zz_601;
  reg        [15:0]   _zz_602;
  reg        [15:0]   _zz_603;
  reg        [15:0]   _zz_604;
  reg        [15:0]   _zz_605;
  reg        [15:0]   _zz_606;
  reg        [15:0]   _zz_607;
  reg        [15:0]   _zz_608;
  reg        [15:0]   _zz_609;
  reg        [15:0]   _zz_610;
  reg        [15:0]   _zz_611;
  reg        [15:0]   _zz_612;
  reg        [15:0]   _zz_613;
  reg        [15:0]   _zz_614;
  reg        [15:0]   _zz_615;
  reg        [15:0]   _zz_616;
  reg        [15:0]   _zz_617;
  reg        [15:0]   _zz_618;
  reg        [15:0]   _zz_619;
  reg        [15:0]   _zz_620;
  reg        [15:0]   _zz_621;
  reg        [15:0]   _zz_622;
  reg        [15:0]   _zz_623;
  reg        [15:0]   _zz_624;
  reg        [15:0]   _zz_625;
  reg        [15:0]   _zz_626;
  reg        [15:0]   _zz_627;
  reg        [15:0]   _zz_628;
  reg        [15:0]   _zz_629;
  reg        [15:0]   _zz_630;
  reg        [15:0]   _zz_631;
  reg        [15:0]   _zz_632;
  reg        [15:0]   _zz_633;
  reg        [15:0]   _zz_634;
  reg        [15:0]   _zz_635;
  reg        [15:0]   _zz_636;
  reg        [15:0]   _zz_637;
  reg        [15:0]   _zz_638;
  reg        [15:0]   _zz_639;
  reg        [15:0]   _zz_640;
  reg        [15:0]   _zz_641;
  reg        [15:0]   _zz_642;
  reg        [15:0]   _zz_643;
  reg        [15:0]   _zz_644;
  reg        [15:0]   _zz_645;
  reg        [15:0]   _zz_646;
  reg        [15:0]   _zz_647;
  reg        [15:0]   _zz_648;
  reg        [15:0]   _zz_649;
  reg        [15:0]   _zz_650;
  reg        [15:0]   _zz_651;
  reg        [15:0]   _zz_652;
  reg        [15:0]   _zz_653;
  reg        [15:0]   _zz_654;
  reg        [15:0]   _zz_655;
  reg        [15:0]   _zz_656;
  reg        [15:0]   _zz_657;
  reg        [15:0]   _zz_658;
  reg        [15:0]   _zz_659;
  reg        [15:0]   _zz_660;
  reg        [15:0]   _zz_661;
  reg        [15:0]   _zz_662;
  reg        [15:0]   _zz_663;
  reg        [15:0]   _zz_664;
  reg        [15:0]   _zz_665;
  reg        [15:0]   _zz_666;
  reg        [15:0]   _zz_667;
  reg        [15:0]   _zz_668;
  reg        [15:0]   _zz_669;
  reg        [15:0]   _zz_670;
  reg        [15:0]   _zz_671;
  reg        [15:0]   _zz_672;
  reg        [15:0]   _zz_673;
  reg        [15:0]   _zz_674;
  reg        [15:0]   _zz_675;
  reg        [15:0]   _zz_676;
  reg        [15:0]   _zz_677;
  reg        [15:0]   _zz_678;
  reg        [15:0]   _zz_679;
  reg        [15:0]   _zz_680;
  reg        [15:0]   _zz_681;
  reg        [15:0]   _zz_682;
  reg        [15:0]   _zz_683;
  reg        [15:0]   _zz_684;
  reg        [15:0]   _zz_685;
  reg        [15:0]   _zz_686;
  reg        [15:0]   _zz_687;
  reg        [15:0]   _zz_688;
  reg        [15:0]   _zz_689;
  reg        [15:0]   _zz_690;
  reg        [15:0]   _zz_691;
  reg        [15:0]   _zz_692;
  reg        [15:0]   _zz_693;
  reg        [15:0]   _zz_694;
  reg        [15:0]   _zz_695;
  reg        [15:0]   _zz_696;
  reg        [15:0]   _zz_697;
  reg        [15:0]   _zz_698;
  reg        [15:0]   _zz_699;
  reg        [15:0]   _zz_700;
  reg        [15:0]   _zz_701;
  reg        [15:0]   _zz_702;
  reg        [15:0]   _zz_703;
  reg        [15:0]   _zz_704;
  reg        [15:0]   _zz_705;
  reg        [15:0]   _zz_706;
  reg        [15:0]   _zz_707;
  reg        [15:0]   _zz_708;
  reg        [15:0]   _zz_709;
  reg        [15:0]   _zz_710;
  reg        [15:0]   _zz_711;
  reg        [15:0]   _zz_712;
  reg        [15:0]   _zz_713;
  reg        [15:0]   _zz_714;
  reg        [15:0]   _zz_715;
  reg        [15:0]   _zz_716;
  reg        [15:0]   _zz_717;
  reg        [15:0]   _zz_718;
  reg        [15:0]   _zz_719;
  reg        [15:0]   _zz_720;
  reg        [15:0]   _zz_721;
  reg        [15:0]   _zz_722;
  reg        [15:0]   _zz_723;
  reg        [15:0]   _zz_724;
  reg        [15:0]   _zz_725;
  reg        [15:0]   _zz_726;
  reg        [15:0]   _zz_727;
  reg        [15:0]   _zz_728;
  reg        [15:0]   _zz_729;
  reg        [15:0]   _zz_730;
  reg        [15:0]   _zz_731;
  reg        [15:0]   _zz_732;
  reg        [15:0]   _zz_733;
  reg        [15:0]   _zz_734;
  reg        [15:0]   _zz_735;
  reg        [15:0]   _zz_736;
  reg        [15:0]   _zz_737;
  reg        [15:0]   _zz_738;
  reg        [15:0]   _zz_739;
  reg        [15:0]   _zz_740;
  reg        [15:0]   _zz_741;
  reg        [15:0]   _zz_742;
  reg        [15:0]   _zz_743;
  reg        [15:0]   _zz_744;
  reg        [15:0]   _zz_745;
  reg        [15:0]   _zz_746;
  reg        [15:0]   _zz_747;
  reg        [15:0]   _zz_748;
  reg        [15:0]   _zz_749;
  reg        [15:0]   _zz_750;
  reg        [15:0]   _zz_751;
  reg        [15:0]   _zz_752;
  reg        [15:0]   _zz_753;
  reg        [15:0]   _zz_754;
  reg        [15:0]   _zz_755;
  reg        [15:0]   _zz_756;
  reg        [15:0]   _zz_757;
  reg        [15:0]   _zz_758;
  reg        [15:0]   _zz_759;
  reg        [15:0]   _zz_760;
  reg        [15:0]   _zz_761;
  reg        [15:0]   _zz_762;
  reg        [15:0]   _zz_763;
  reg        [15:0]   _zz_764;
  reg        [15:0]   _zz_765;
  reg        [15:0]   _zz_766;
  reg        [15:0]   _zz_767;
  reg        [15:0]   _zz_768;
  reg        [15:0]   _zz_769;
  reg        [15:0]   _zz_770;
  reg        [15:0]   _zz_771;
  reg        [15:0]   _zz_772;
  reg        [15:0]   _zz_773;
  reg        [15:0]   _zz_774;
  reg        [15:0]   _zz_775;
  reg        [15:0]   _zz_776;
  reg        [15:0]   _zz_777;
  reg        [15:0]   _zz_778;
  reg        [15:0]   _zz_779;
  reg        [15:0]   _zz_780;
  reg        [15:0]   _zz_781;
  reg        [15:0]   _zz_782;
  reg        [15:0]   _zz_783;
  reg        [15:0]   _zz_784;
  reg        [15:0]   _zz_785;
  reg        [15:0]   _zz_786;
  reg        [15:0]   _zz_787;
  reg        [15:0]   _zz_788;
  reg        [15:0]   _zz_789;
  reg        [15:0]   _zz_790;
  reg        [15:0]   _zz_791;
  reg        [15:0]   _zz_792;
  reg        [15:0]   _zz_793;
  reg        [15:0]   _zz_794;
  reg        [15:0]   _zz_795;
  reg        [15:0]   _zz_796;
  reg        [15:0]   _zz_797;
  reg        [15:0]   _zz_798;
  reg        [15:0]   _zz_799;
  reg        [15:0]   _zz_800;
  reg        [15:0]   _zz_801;
  reg        [15:0]   _zz_802;
  reg        [15:0]   _zz_803;
  reg        [15:0]   _zz_804;
  reg        [15:0]   _zz_805;
  reg        [15:0]   _zz_806;
  reg        [15:0]   _zz_807;
  reg        [15:0]   _zz_808;
  reg        [15:0]   _zz_809;
  reg        [15:0]   _zz_810;
  reg        [15:0]   _zz_811;
  reg        [15:0]   _zz_812;
  reg        [15:0]   _zz_813;
  reg        [15:0]   _zz_814;
  reg        [15:0]   _zz_815;
  reg        [15:0]   _zz_816;
  reg        [15:0]   _zz_817;
  reg        [15:0]   _zz_818;
  reg        [15:0]   _zz_819;
  reg        [15:0]   _zz_820;
  reg        [15:0]   _zz_821;
  reg        [15:0]   _zz_822;
  reg        [15:0]   _zz_823;
  reg        [15:0]   _zz_824;
  reg        [15:0]   _zz_825;
  reg        [15:0]   _zz_826;
  reg        [15:0]   _zz_827;
  reg        [15:0]   _zz_828;
  reg        [15:0]   _zz_829;
  reg        [15:0]   _zz_830;
  reg        [15:0]   _zz_831;
  reg        [15:0]   _zz_832;
  reg        [15:0]   _zz_833;
  reg        [15:0]   _zz_834;
  reg        [15:0]   _zz_835;
  reg        [15:0]   _zz_836;
  reg        [15:0]   _zz_837;
  reg        [15:0]   _zz_838;
  reg        [15:0]   _zz_839;
  reg        [15:0]   _zz_840;
  reg        [15:0]   _zz_841;
  reg        [15:0]   _zz_842;
  reg        [15:0]   _zz_843;
  reg        [15:0]   _zz_844;
  reg        [15:0]   _zz_845;
  reg        [15:0]   _zz_846;
  reg        [15:0]   _zz_847;
  reg        [15:0]   _zz_848;
  reg        [15:0]   _zz_849;
  reg        [15:0]   _zz_850;
  reg        [15:0]   _zz_851;
  reg        [15:0]   _zz_852;
  reg        [15:0]   _zz_853;
  reg        [15:0]   _zz_854;
  reg        [15:0]   _zz_855;
  reg        [15:0]   _zz_856;
  reg        [15:0]   _zz_857;
  reg        [15:0]   _zz_858;
  reg        [15:0]   _zz_859;
  reg        [15:0]   _zz_860;
  reg        [15:0]   _zz_861;
  reg        [15:0]   _zz_862;
  reg        [15:0]   _zz_863;
  reg        [15:0]   _zz_864;
  reg        [15:0]   _zz_865;
  reg        [15:0]   _zz_866;
  reg        [15:0]   _zz_867;
  reg        [15:0]   _zz_868;
  reg        [15:0]   _zz_869;
  reg        [15:0]   _zz_870;
  reg        [15:0]   _zz_871;
  reg        [15:0]   _zz_872;
  reg        [15:0]   _zz_873;
  reg        [15:0]   _zz_874;
  reg        [15:0]   _zz_875;
  reg        [15:0]   _zz_876;
  reg        [15:0]   _zz_877;
  reg        [15:0]   _zz_878;
  reg        [15:0]   _zz_879;
  reg        [15:0]   _zz_880;
  reg        [15:0]   _zz_881;
  reg        [15:0]   _zz_882;
  reg        [15:0]   _zz_883;
  reg        [15:0]   _zz_884;
  reg        [15:0]   _zz_885;
  reg        [15:0]   _zz_886;
  reg        [15:0]   _zz_887;
  reg        [15:0]   _zz_888;
  reg        [15:0]   _zz_889;
  reg        [15:0]   _zz_890;
  reg        [15:0]   _zz_891;
  reg        [15:0]   _zz_892;
  reg        [15:0]   _zz_893;
  reg        [15:0]   _zz_894;
  reg        [15:0]   _zz_895;
  reg        [15:0]   _zz_896;
  reg        [15:0]   _zz_897;
  reg        [15:0]   _zz_898;
  reg        [15:0]   _zz_899;
  reg        [15:0]   _zz_900;
  reg        [15:0]   _zz_901;
  reg        [15:0]   _zz_902;
  reg        [15:0]   _zz_903;
  reg        [15:0]   _zz_904;
  reg        [15:0]   _zz_905;
  reg        [15:0]   _zz_906;
  reg        [15:0]   _zz_907;
  reg        [15:0]   _zz_908;
  reg        [15:0]   _zz_909;
  reg        [15:0]   _zz_910;
  reg        [15:0]   _zz_911;
  reg        [15:0]   _zz_912;
  reg        [15:0]   _zz_913;
  reg        [15:0]   _zz_914;
  reg        [15:0]   _zz_915;
  reg        [15:0]   _zz_916;
  reg        [15:0]   _zz_917;
  reg        [15:0]   _zz_918;
  reg        [15:0]   _zz_919;
  reg        [15:0]   _zz_920;
  reg        [15:0]   _zz_921;
  reg        [15:0]   _zz_922;
  reg        [15:0]   _zz_923;
  reg        [15:0]   _zz_924;
  reg        [15:0]   _zz_925;
  reg        [15:0]   _zz_926;
  reg        [15:0]   _zz_927;
  reg        [15:0]   _zz_928;
  reg        [15:0]   _zz_929;
  reg        [15:0]   _zz_930;
  reg        [15:0]   _zz_931;
  reg        [15:0]   _zz_932;
  reg        [15:0]   _zz_933;
  reg        [15:0]   _zz_934;
  reg        [15:0]   _zz_935;
  reg        [15:0]   _zz_936;
  reg        [15:0]   _zz_937;
  reg        [15:0]   _zz_938;
  reg        [15:0]   _zz_939;
  reg        [15:0]   _zz_940;
  reg        [15:0]   _zz_941;
  reg        [15:0]   _zz_942;
  reg        [15:0]   _zz_943;
  reg        [15:0]   _zz_944;
  reg        [15:0]   _zz_945;
  reg        [15:0]   _zz_946;
  reg        [15:0]   _zz_947;
  reg        [15:0]   _zz_948;
  reg        [15:0]   _zz_949;
  reg        [15:0]   _zz_950;
  reg        [15:0]   _zz_951;
  reg        [15:0]   _zz_952;
  reg        [15:0]   _zz_953;
  reg        [15:0]   _zz_954;
  reg        [15:0]   _zz_955;
  reg        [15:0]   _zz_956;
  reg        [15:0]   _zz_957;
  reg        [15:0]   _zz_958;
  reg        [15:0]   _zz_959;
  reg        [15:0]   _zz_960;
  reg        [15:0]   _zz_961;
  reg        [15:0]   _zz_962;
  reg        [15:0]   _zz_963;
  reg        [15:0]   _zz_964;
  reg        [15:0]   _zz_965;
  reg        [15:0]   _zz_966;
  reg        [15:0]   _zz_967;
  reg        [15:0]   _zz_968;
  reg        [15:0]   _zz_969;
  reg        [15:0]   _zz_970;
  reg        [15:0]   _zz_971;
  reg        [15:0]   _zz_972;
  reg        [15:0]   _zz_973;
  reg        [15:0]   _zz_974;
  reg        [15:0]   _zz_975;
  reg        [15:0]   _zz_976;
  reg        [15:0]   _zz_977;
  reg        [15:0]   _zz_978;
  reg        [15:0]   _zz_979;
  reg        [15:0]   _zz_980;
  reg        [15:0]   _zz_981;
  reg        [15:0]   _zz_982;
  reg        [15:0]   _zz_983;
  reg        [15:0]   _zz_984;
  reg        [15:0]   _zz_985;
  reg        [15:0]   _zz_986;
  reg        [15:0]   _zz_987;
  reg        [15:0]   _zz_988;
  reg        [15:0]   _zz_989;
  reg        [15:0]   _zz_990;
  reg        [15:0]   _zz_991;
  reg        [15:0]   _zz_992;
  reg        [15:0]   _zz_993;
  reg        [15:0]   _zz_994;
  reg        [15:0]   _zz_995;
  reg        [15:0]   _zz_996;
  reg        [15:0]   _zz_997;
  reg        [15:0]   _zz_998;
  reg        [15:0]   _zz_999;
  reg        [15:0]   _zz_1000;
  reg        [15:0]   _zz_1001;
  reg        [15:0]   _zz_1002;
  reg        [15:0]   _zz_1003;
  reg        [15:0]   _zz_1004;
  reg        [15:0]   _zz_1005;
  reg        [15:0]   _zz_1006;
  reg        [15:0]   _zz_1007;
  reg        [15:0]   _zz_1008;
  reg        [15:0]   _zz_1009;
  reg        [15:0]   _zz_1010;
  reg        [15:0]   _zz_1011;
  reg        [15:0]   _zz_1012;
  reg        [15:0]   _zz_1013;
  reg        [15:0]   _zz_1014;
  reg        [15:0]   _zz_1015;
  reg        [15:0]   _zz_1016;
  reg        [15:0]   _zz_1017;
  reg        [15:0]   _zz_1018;
  reg        [15:0]   _zz_1019;
  reg        [15:0]   _zz_1020;
  reg        [15:0]   _zz_1021;
  reg        [15:0]   _zz_1022;
  reg        [15:0]   _zz_1023;
  reg        [15:0]   _zz_1024;
  reg        [15:0]   _zz_1025;
  reg        [15:0]   _zz_1026;
  reg        [15:0]   _zz_1027;
  reg        [15:0]   _zz_1028;
  reg        [15:0]   _zz_1029;
  reg        [15:0]   _zz_1030;
  reg        [15:0]   _zz_1031;
  reg        [15:0]   _zz_1032;
  reg        [15:0]   _zz_1033;
  reg        [15:0]   _zz_1034;
  reg        [15:0]   _zz_1035;
  reg        [15:0]   _zz_1036;
  reg        [15:0]   _zz_1037;
  reg        [15:0]   _zz_1038;
  reg        [15:0]   _zz_1039;
  reg        [15:0]   _zz_1040;
  reg        [15:0]   _zz_1041;
  reg        [15:0]   _zz_1042;
  reg        [15:0]   _zz_1043;
  reg        [15:0]   _zz_1044;
  reg        [15:0]   _zz_1045;
  reg        [15:0]   _zz_1046;
  reg        [15:0]   _zz_1047;
  reg        [15:0]   _zz_1048;
  reg        [15:0]   _zz_1049;
  reg        [15:0]   _zz_1050;
  reg        [15:0]   _zz_1051;
  reg        [15:0]   _zz_1052;
  reg        [15:0]   _zz_1053;
  reg        [15:0]   _zz_1054;
  reg        [15:0]   _zz_1055;
  reg        [15:0]   _zz_1056;
  reg        [15:0]   _zz_1057;
  reg        [15:0]   _zz_1058;
  reg        [15:0]   _zz_1059;
  reg        [15:0]   _zz_1060;
  reg        [15:0]   _zz_1061;
  reg        [15:0]   _zz_1062;
  reg        [15:0]   _zz_1063;
  reg        [15:0]   _zz_1064;
  reg        [15:0]   _zz_1065;
  reg        [15:0]   _zz_1066;
  reg        [15:0]   _zz_1067;
  reg        [15:0]   _zz_1068;
  reg        [15:0]   _zz_1069;
  reg        [15:0]   _zz_1070;
  reg        [15:0]   _zz_1071;
  reg        [15:0]   _zz_1072;
  reg        [15:0]   _zz_1073;
  reg        [15:0]   _zz_1074;
  reg        [15:0]   _zz_1075;
  reg        [15:0]   _zz_1076;
  reg        [15:0]   _zz_1077;
  reg        [15:0]   _zz_1078;
  reg        [15:0]   _zz_1079;
  reg        [15:0]   _zz_1080;
  reg        [15:0]   _zz_1081;
  reg        [15:0]   _zz_1082;
  reg        [15:0]   _zz_1083;
  reg        [15:0]   _zz_1084;
  reg        [15:0]   _zz_1085;
  reg        [15:0]   _zz_1086;
  reg        [15:0]   _zz_1087;
  reg        [15:0]   _zz_1088;
  reg        [15:0]   _zz_1089;
  reg        [15:0]   _zz_1090;
  reg        [15:0]   _zz_1091;
  reg        [15:0]   _zz_1092;
  reg        [15:0]   _zz_1093;
  reg        [15:0]   _zz_1094;
  reg        [15:0]   _zz_1095;
  reg        [15:0]   _zz_1096;
  reg        [15:0]   _zz_1097;
  reg        [15:0]   _zz_1098;
  reg        [15:0]   _zz_1099;
  reg        [15:0]   _zz_1100;
  reg        [15:0]   _zz_1101;
  reg        [15:0]   _zz_1102;
  reg        [15:0]   _zz_1103;
  reg        [15:0]   _zz_1104;
  reg        [15:0]   _zz_1105;
  reg        [15:0]   _zz_1106;
  reg        [15:0]   _zz_1107;
  reg        [15:0]   _zz_1108;
  reg        [15:0]   _zz_1109;
  reg        [15:0]   _zz_1110;
  reg        [15:0]   _zz_1111;
  reg        [15:0]   _zz_1112;
  reg        [15:0]   _zz_1113;
  reg        [15:0]   _zz_1114;
  reg        [15:0]   _zz_1115;
  reg        [15:0]   _zz_1116;
  reg        [15:0]   _zz_1117;
  reg        [15:0]   _zz_1118;
  reg        [15:0]   _zz_1119;
  reg        [15:0]   _zz_1120;
  reg        [15:0]   _zz_1121;
  reg        [15:0]   _zz_1122;
  reg        [15:0]   _zz_1123;
  reg        [15:0]   _zz_1124;
  reg        [15:0]   _zz_1125;
  reg        [15:0]   _zz_1126;
  reg        [15:0]   _zz_1127;
  reg        [15:0]   _zz_1128;
  reg        [15:0]   _zz_1129;
  reg        [15:0]   _zz_1130;
  reg        [15:0]   _zz_1131;
  reg        [15:0]   _zz_1132;
  reg        [15:0]   _zz_1133;
  reg        [15:0]   _zz_1134;
  reg        [15:0]   _zz_1135;
  reg        [15:0]   _zz_1136;
  reg        [15:0]   _zz_1137;
  reg        [15:0]   _zz_1138;
  reg        [15:0]   _zz_1139;
  reg        [15:0]   _zz_1140;
  reg        [15:0]   _zz_1141;
  reg        [15:0]   _zz_1142;
  reg        [15:0]   _zz_1143;
  reg        [15:0]   _zz_1144;
  reg        [15:0]   _zz_1145;
  reg        [15:0]   _zz_1146;
  reg        [15:0]   _zz_1147;
  reg        [15:0]   _zz_1148;
  reg        [15:0]   _zz_1149;
  reg        [15:0]   _zz_1150;
  reg        [15:0]   _zz_1151;
  reg        [15:0]   _zz_1152;
  reg        [15:0]   _zz_1153;
  reg        [15:0]   _zz_1154;
  reg        [15:0]   _zz_1155;
  reg        [15:0]   _zz_1156;
  reg        [15:0]   _zz_1157;
  reg        [15:0]   _zz_1158;
  reg        [15:0]   _zz_1159;
  reg        [15:0]   _zz_1160;
  reg        [15:0]   _zz_1161;
  reg        [15:0]   _zz_1162;
  reg        [15:0]   _zz_1163;
  reg        [15:0]   _zz_1164;
  reg        [15:0]   _zz_1165;
  reg        [15:0]   _zz_1166;
  reg        [15:0]   _zz_1167;
  reg        [15:0]   _zz_1168;
  reg        [15:0]   _zz_1169;
  reg        [15:0]   _zz_1170;
  reg        [15:0]   _zz_1171;
  reg        [15:0]   _zz_1172;
  reg        [15:0]   _zz_1173;
  reg        [15:0]   _zz_1174;
  reg        [15:0]   _zz_1175;
  reg        [15:0]   _zz_1176;
  reg        [15:0]   _zz_1177;
  reg        [15:0]   _zz_1178;
  reg        [15:0]   _zz_1179;
  reg        [15:0]   _zz_1180;
  reg        [15:0]   _zz_1181;
  reg        [15:0]   _zz_1182;
  reg        [15:0]   _zz_1183;
  reg        [15:0]   _zz_1184;
  reg        [15:0]   _zz_1185;
  reg        [15:0]   _zz_1186;
  reg        [15:0]   _zz_1187;
  reg        [15:0]   _zz_1188;
  reg        [15:0]   _zz_1189;
  reg        [15:0]   _zz_1190;
  reg        [15:0]   _zz_1191;
  reg        [15:0]   _zz_1192;
  reg        [15:0]   _zz_1193;
  reg        [15:0]   _zz_1194;
  reg        [15:0]   _zz_1195;
  reg        [15:0]   _zz_1196;
  reg        [15:0]   _zz_1197;
  reg        [15:0]   _zz_1198;
  reg        [15:0]   _zz_1199;
  reg        [15:0]   _zz_1200;
  reg        [15:0]   _zz_1201;
  reg        [15:0]   _zz_1202;
  reg        [15:0]   _zz_1203;
  reg        [15:0]   _zz_1204;
  reg        [15:0]   _zz_1205;
  reg        [15:0]   _zz_1206;
  reg        [15:0]   _zz_1207;
  reg        [15:0]   _zz_1208;
  reg        [15:0]   _zz_1209;
  reg        [15:0]   _zz_1210;
  reg        [15:0]   _zz_1211;
  reg        [15:0]   _zz_1212;
  reg        [15:0]   _zz_1213;
  reg        [15:0]   _zz_1214;
  reg        [15:0]   _zz_1215;
  reg        [15:0]   _zz_1216;
  reg        [15:0]   _zz_1217;
  reg        [15:0]   _zz_1218;
  reg        [15:0]   _zz_1219;
  reg        [15:0]   _zz_1220;
  reg        [15:0]   _zz_1221;
  reg        [15:0]   _zz_1222;
  reg        [15:0]   _zz_1223;
  reg        [15:0]   _zz_1224;
  reg        [15:0]   _zz_1225;
  reg        [15:0]   _zz_1226;
  reg        [15:0]   _zz_1227;
  reg        [15:0]   _zz_1228;
  reg        [15:0]   _zz_1229;
  reg        [15:0]   _zz_1230;
  reg        [15:0]   _zz_1231;
  reg        [15:0]   _zz_1232;
  reg        [15:0]   _zz_1233;
  reg        [15:0]   _zz_1234;
  reg        [15:0]   _zz_1235;
  reg        [15:0]   _zz_1236;
  reg        [15:0]   _zz_1237;
  reg        [15:0]   _zz_1238;
  reg        [15:0]   _zz_1239;
  reg        [15:0]   _zz_1240;
  reg        [15:0]   _zz_1241;
  reg        [15:0]   _zz_1242;
  reg        [15:0]   _zz_1243;
  reg        [15:0]   _zz_1244;
  reg        [15:0]   _zz_1245;
  reg        [15:0]   _zz_1246;
  reg        [15:0]   _zz_1247;
  reg        [15:0]   _zz_1248;
  reg        [15:0]   _zz_1249;
  reg        [15:0]   _zz_1250;
  reg        [15:0]   _zz_1251;
  reg        [15:0]   _zz_1252;
  reg        [15:0]   _zz_1253;
  reg        [15:0]   _zz_1254;
  reg        [15:0]   _zz_1255;
  reg        [15:0]   _zz_1256;
  reg        [15:0]   _zz_1257;
  reg        [15:0]   _zz_1258;
  reg        [15:0]   _zz_1259;
  reg        [15:0]   _zz_1260;
  reg        [15:0]   _zz_1261;
  reg        [15:0]   _zz_1262;
  reg        [15:0]   _zz_1263;
  reg        [15:0]   _zz_1264;
  reg        [15:0]   _zz_1265;
  reg        [15:0]   _zz_1266;
  reg        [15:0]   _zz_1267;
  reg        [15:0]   _zz_1268;
  reg        [15:0]   _zz_1269;
  reg        [15:0]   _zz_1270;
  reg        [15:0]   _zz_1271;
  reg        [15:0]   _zz_1272;
  reg        [15:0]   _zz_1273;
  reg        [15:0]   _zz_1274;
  reg        [15:0]   _zz_1275;
  reg        [15:0]   _zz_1276;
  reg        [15:0]   _zz_1277;
  reg        [15:0]   _zz_1278;
  reg        [15:0]   _zz_1279;
  reg        [15:0]   _zz_1280;
  reg        [15:0]   _zz_1281;
  reg        [15:0]   _zz_1282;
  reg        [15:0]   _zz_1283;
  reg        [15:0]   _zz_1284;
  reg        [15:0]   _zz_1285;
  reg        [15:0]   _zz_1286;
  reg        [15:0]   _zz_1287;
  reg        [15:0]   _zz_1288;
  reg        [15:0]   _zz_1289;
  reg        [15:0]   _zz_1290;
  reg        [15:0]   _zz_1291;
  reg        [15:0]   _zz_1292;
  reg        [15:0]   _zz_1293;
  reg        [15:0]   _zz_1294;
  reg        [15:0]   _zz_1295;
  reg        [15:0]   _zz_1296;
  reg        [15:0]   _zz_1297;
  reg        [15:0]   _zz_1298;
  reg        [15:0]   _zz_1299;
  reg        [15:0]   _zz_1300;
  reg        [15:0]   _zz_1301;
  reg        [15:0]   _zz_1302;
  reg        [15:0]   _zz_1303;
  reg        [15:0]   _zz_1304;
  reg        [15:0]   _zz_1305;
  reg        [15:0]   _zz_1306;
  reg        [15:0]   _zz_1307;
  reg        [15:0]   _zz_1308;
  reg        [15:0]   _zz_1309;
  reg        [15:0]   _zz_1310;
  reg        [15:0]   _zz_1311;
  reg        [15:0]   _zz_1312;
  reg        [15:0]   _zz_1313;
  reg        [15:0]   _zz_1314;
  reg        [15:0]   _zz_1315;
  reg        [15:0]   _zz_1316;
  reg        [15:0]   _zz_1317;
  reg        [15:0]   _zz_1318;
  reg        [15:0]   _zz_1319;
  reg        [15:0]   _zz_1320;
  reg        [15:0]   _zz_1321;
  reg        [15:0]   _zz_1322;
  reg        [15:0]   _zz_1323;
  reg        [15:0]   _zz_1324;
  reg        [15:0]   _zz_1325;
  reg        [15:0]   _zz_1326;
  reg        [15:0]   _zz_1327;
  reg        [15:0]   _zz_1328;
  reg        [15:0]   _zz_1329;
  reg        [15:0]   _zz_1330;
  reg        [15:0]   _zz_1331;
  reg        [15:0]   _zz_1332;
  reg        [15:0]   _zz_1333;
  reg        [15:0]   _zz_1334;
  reg        [15:0]   _zz_1335;
  reg        [15:0]   _zz_1336;
  reg        [15:0]   _zz_1337;
  reg        [15:0]   _zz_1338;
  reg        [15:0]   _zz_1339;
  reg        [15:0]   _zz_1340;
  reg        [15:0]   _zz_1341;
  reg        [15:0]   _zz_1342;
  reg        [15:0]   _zz_1343;
  reg        [15:0]   _zz_1344;
  reg        [15:0]   _zz_1345;
  reg        [15:0]   _zz_1346;
  reg        [15:0]   _zz_1347;
  reg        [15:0]   _zz_1348;
  reg        [15:0]   _zz_1349;
  reg        [15:0]   _zz_1350;
  reg        [15:0]   _zz_1351;
  reg        [15:0]   _zz_1352;
  reg        [15:0]   _zz_1353;
  reg        [15:0]   _zz_1354;
  reg        [15:0]   _zz_1355;
  reg        [15:0]   _zz_1356;
  reg        [15:0]   _zz_1357;
  reg        [15:0]   _zz_1358;
  reg        [15:0]   _zz_1359;
  reg        [15:0]   _zz_1360;
  reg        [15:0]   _zz_1361;
  reg        [15:0]   _zz_1362;
  reg        [15:0]   _zz_1363;
  reg        [15:0]   _zz_1364;
  reg        [15:0]   _zz_1365;
  reg        [15:0]   _zz_1366;
  reg        [15:0]   _zz_1367;
  reg        [15:0]   _zz_1368;
  reg        [15:0]   _zz_1369;
  reg        [15:0]   _zz_1370;
  reg        [15:0]   _zz_1371;
  reg        [15:0]   _zz_1372;
  reg        [15:0]   _zz_1373;
  reg        [15:0]   _zz_1374;
  reg        [15:0]   _zz_1375;
  reg        [15:0]   _zz_1376;
  reg        [15:0]   _zz_1377;
  reg        [15:0]   _zz_1378;
  reg        [15:0]   _zz_1379;
  reg        [15:0]   _zz_1380;
  reg        [15:0]   _zz_1381;
  reg        [15:0]   _zz_1382;
  reg        [15:0]   _zz_1383;
  reg        [15:0]   _zz_1384;
  reg        [15:0]   _zz_1385;
  reg        [15:0]   _zz_1386;
  reg        [15:0]   _zz_1387;
  reg        [15:0]   _zz_1388;
  reg        [15:0]   _zz_1389;
  reg        [15:0]   _zz_1390;
  reg        [15:0]   _zz_1391;
  reg        [15:0]   _zz_1392;
  reg        [15:0]   _zz_1393;
  reg        [15:0]   _zz_1394;
  reg        [15:0]   _zz_1395;
  reg        [15:0]   _zz_1396;
  reg        [15:0]   _zz_1397;
  reg        [15:0]   _zz_1398;
  reg        [15:0]   _zz_1399;
  reg        [15:0]   _zz_1400;
  reg        [15:0]   _zz_1401;
  reg        [15:0]   _zz_1402;
  reg        [15:0]   _zz_1403;
  reg        [15:0]   _zz_1404;
  reg        [15:0]   _zz_1405;
  reg        [15:0]   _zz_1406;
  reg        [15:0]   _zz_1407;
  reg        [15:0]   _zz_1408;
  reg        [15:0]   _zz_1409;
  reg        [15:0]   _zz_1410;
  reg        [15:0]   _zz_1411;
  reg        [15:0]   _zz_1412;
  reg        [15:0]   _zz_1413;
  reg        [15:0]   _zz_1414;
  reg        [15:0]   _zz_1415;
  reg        [15:0]   _zz_1416;
  reg        [15:0]   _zz_1417;
  reg        [15:0]   _zz_1418;
  reg        [15:0]   _zz_1419;
  reg        [15:0]   _zz_1420;
  reg        [15:0]   _zz_1421;
  reg        [15:0]   _zz_1422;
  reg        [15:0]   _zz_1423;
  reg        [15:0]   _zz_1424;
  reg        [15:0]   _zz_1425;
  reg        [15:0]   _zz_1426;
  reg        [15:0]   _zz_1427;
  reg        [15:0]   _zz_1428;
  reg        [15:0]   _zz_1429;
  reg        [15:0]   _zz_1430;
  reg        [15:0]   _zz_1431;
  reg        [15:0]   _zz_1432;
  reg        [15:0]   _zz_1433;
  reg        [15:0]   _zz_1434;
  reg        [15:0]   _zz_1435;
  reg        [15:0]   _zz_1436;
  reg        [15:0]   _zz_1437;
  reg        [15:0]   _zz_1438;
  reg        [15:0]   _zz_1439;
  reg        [15:0]   _zz_1440;
  reg        [15:0]   _zz_1441;
  reg        [15:0]   _zz_1442;
  reg        [15:0]   _zz_1443;
  reg        [15:0]   _zz_1444;
  reg        [15:0]   _zz_1445;
  reg        [15:0]   _zz_1446;
  reg        [15:0]   _zz_1447;
  reg        [15:0]   _zz_1448;
  reg        [15:0]   _zz_1449;
  reg        [15:0]   _zz_1450;
  reg        [15:0]   _zz_1451;
  reg        [15:0]   _zz_1452;
  reg        [15:0]   _zz_1453;
  reg        [15:0]   _zz_1454;
  reg        [15:0]   _zz_1455;
  reg        [15:0]   _zz_1456;
  reg        [15:0]   _zz_1457;
  reg        [15:0]   _zz_1458;
  reg        [15:0]   _zz_1459;
  reg        [15:0]   _zz_1460;
  reg        [15:0]   _zz_1461;
  reg        [15:0]   _zz_1462;
  reg        [15:0]   _zz_1463;
  reg        [15:0]   _zz_1464;
  reg        [15:0]   _zz_1465;
  reg        [15:0]   _zz_1466;
  reg        [15:0]   _zz_1467;
  reg        [15:0]   _zz_1468;
  reg        [15:0]   _zz_1469;
  reg        [15:0]   _zz_1470;
  reg        [15:0]   _zz_1471;
  reg        [15:0]   _zz_1472;
  reg        [15:0]   _zz_1473;
  reg        [15:0]   _zz_1474;
  reg        [15:0]   _zz_1475;
  reg        [15:0]   _zz_1476;
  reg        [15:0]   _zz_1477;
  reg        [15:0]   _zz_1478;
  reg        [15:0]   _zz_1479;
  reg        [15:0]   _zz_1480;
  reg        [15:0]   _zz_1481;
  reg        [15:0]   _zz_1482;
  reg        [15:0]   _zz_1483;
  reg        [15:0]   _zz_1484;
  reg        [15:0]   _zz_1485;
  reg        [15:0]   _zz_1486;
  reg        [15:0]   _zz_1487;
  reg        [15:0]   _zz_1488;
  reg        [15:0]   _zz_1489;
  reg        [15:0]   _zz_1490;
  reg        [15:0]   _zz_1491;
  reg        [15:0]   _zz_1492;
  reg        [15:0]   _zz_1493;
  reg        [15:0]   _zz_1494;
  reg        [15:0]   _zz_1495;
  reg        [15:0]   _zz_1496;
  reg        [15:0]   _zz_1497;
  reg        [15:0]   _zz_1498;
  reg        [15:0]   _zz_1499;
  reg        [15:0]   _zz_1500;
  reg        [15:0]   _zz_1501;
  reg        [15:0]   _zz_1502;
  reg        [15:0]   _zz_1503;
  reg        [15:0]   _zz_1504;
  reg        [15:0]   _zz_1505;
  reg        [15:0]   _zz_1506;
  reg        [15:0]   _zz_1507;
  reg        [15:0]   _zz_1508;
  reg        [15:0]   _zz_1509;
  reg        [15:0]   _zz_1510;
  reg        [15:0]   _zz_1511;
  reg        [15:0]   _zz_1512;
  reg        [15:0]   _zz_1513;
  reg        [15:0]   _zz_1514;
  reg        [15:0]   _zz_1515;
  reg        [15:0]   _zz_1516;
  reg        [15:0]   _zz_1517;
  reg        [15:0]   _zz_1518;
  reg        [15:0]   _zz_1519;
  reg        [15:0]   _zz_1520;
  reg        [15:0]   _zz_1521;
  reg        [15:0]   _zz_1522;
  reg        [15:0]   _zz_1523;
  reg        [15:0]   _zz_1524;
  reg        [15:0]   _zz_1525;
  reg        [15:0]   _zz_1526;
  reg        [15:0]   _zz_1527;
  reg        [15:0]   _zz_1528;
  reg        [15:0]   _zz_1529;
  reg        [15:0]   _zz_1530;
  reg        [15:0]   _zz_1531;
  reg        [15:0]   _zz_1532;
  reg        [15:0]   _zz_1533;
  reg        [15:0]   _zz_1534;
  reg        [15:0]   _zz_1535;
  reg        [15:0]   _zz_1536;
  reg        [15:0]   _zz_1537;
  reg        [15:0]   _zz_1538;
  reg        [15:0]   _zz_1539;
  reg        [15:0]   _zz_1540;
  reg        [15:0]   _zz_1541;
  reg        [15:0]   _zz_1542;
  reg        [15:0]   _zz_1543;
  reg        [15:0]   _zz_1544;
  reg        [15:0]   _zz_1545;
  reg        [15:0]   _zz_1546;
  reg        [15:0]   _zz_1547;
  reg        [15:0]   _zz_1548;
  reg        [15:0]   _zz_1549;
  reg        [15:0]   _zz_1550;
  reg        [15:0]   _zz_1551;
  reg        [15:0]   _zz_1552;
  reg        [15:0]   _zz_1553;
  reg        [15:0]   _zz_1554;
  reg        [15:0]   _zz_1555;
  reg        [15:0]   _zz_1556;
  reg        [15:0]   _zz_1557;
  reg        [15:0]   _zz_1558;
  reg        [15:0]   _zz_1559;
  reg        [15:0]   _zz_1560;
  reg        [15:0]   _zz_1561;
  reg        [15:0]   _zz_1562;
  reg        [15:0]   _zz_1563;
  reg        [15:0]   _zz_1564;
  reg        [15:0]   _zz_1565;
  reg        [15:0]   _zz_1566;
  reg        [15:0]   _zz_1567;
  reg        [15:0]   _zz_1568;
  reg        [15:0]   _zz_1569;
  reg        [15:0]   _zz_1570;
  reg        [15:0]   _zz_1571;
  reg        [15:0]   _zz_1572;
  reg        [15:0]   _zz_1573;
  reg        [15:0]   _zz_1574;
  reg        [15:0]   _zz_1575;
  reg        [15:0]   _zz_1576;
  reg        [15:0]   _zz_1577;
  reg        [15:0]   _zz_1578;
  reg        [15:0]   _zz_1579;
  reg        [15:0]   _zz_1580;
  reg        [15:0]   _zz_1581;
  reg        [15:0]   _zz_1582;
  reg        [15:0]   _zz_1583;
  reg        [15:0]   _zz_1584;
  reg        [15:0]   _zz_1585;
  reg        [15:0]   _zz_1586;
  reg        [15:0]   _zz_1587;
  reg        [15:0]   _zz_1588;
  reg        [15:0]   _zz_1589;
  reg        [15:0]   _zz_1590;
  reg        [15:0]   _zz_1591;
  reg        [15:0]   _zz_1592;
  reg        [15:0]   _zz_1593;
  reg        [15:0]   _zz_1594;
  reg        [15:0]   _zz_1595;
  reg        [15:0]   _zz_1596;
  reg        [15:0]   _zz_1597;
  reg        [15:0]   _zz_1598;
  reg        [15:0]   _zz_1599;
  reg        [15:0]   _zz_1600;
  reg        [15:0]   _zz_1601;
  reg        [15:0]   _zz_1602;
  reg        [15:0]   _zz_1603;
  reg        [15:0]   _zz_1604;
  reg        [15:0]   _zz_1605;
  reg        [15:0]   _zz_1606;
  reg        [15:0]   _zz_1607;
  reg        [15:0]   _zz_1608;
  reg        [15:0]   _zz_1609;
  reg        [15:0]   _zz_1610;
  reg        [15:0]   _zz_1611;
  reg        [15:0]   _zz_1612;
  reg        [15:0]   _zz_1613;
  reg        [15:0]   _zz_1614;
  reg        [15:0]   _zz_1615;
  reg        [15:0]   _zz_1616;
  reg        [15:0]   _zz_1617;
  reg        [15:0]   _zz_1618;
  reg        [15:0]   _zz_1619;
  reg        [15:0]   _zz_1620;
  reg        [15:0]   _zz_1621;
  reg        [15:0]   _zz_1622;
  reg        [15:0]   _zz_1623;
  reg        [15:0]   _zz_1624;
  reg        [15:0]   _zz_1625;
  reg        [15:0]   _zz_1626;
  reg        [15:0]   _zz_1627;
  reg        [15:0]   _zz_1628;
  reg        [15:0]   _zz_1629;
  reg        [15:0]   _zz_1630;
  reg        [15:0]   _zz_1631;
  reg        [15:0]   _zz_1632;
  reg        [15:0]   _zz_1633;
  reg        [15:0]   _zz_1634;
  reg        [15:0]   _zz_1635;
  reg        [15:0]   _zz_1636;
  reg        [15:0]   _zz_1637;
  reg        [15:0]   _zz_1638;
  reg        [15:0]   _zz_1639;
  reg        [15:0]   _zz_1640;
  reg        [15:0]   _zz_1641;
  reg        [15:0]   _zz_1642;
  reg        [15:0]   _zz_1643;
  reg        [15:0]   _zz_1644;
  reg        [15:0]   _zz_1645;
  reg        [15:0]   _zz_1646;
  reg        [15:0]   _zz_1647;
  reg        [15:0]   _zz_1648;
  reg        [15:0]   _zz_1649;
  reg        [15:0]   _zz_1650;
  reg        [15:0]   _zz_1651;
  reg        [15:0]   _zz_1652;
  reg        [15:0]   _zz_1653;
  reg        [15:0]   _zz_1654;
  reg        [15:0]   _zz_1655;
  reg        [15:0]   _zz_1656;
  reg        [15:0]   _zz_1657;
  reg        [15:0]   _zz_1658;
  reg        [15:0]   _zz_1659;
  reg        [15:0]   _zz_1660;
  reg        [15:0]   _zz_1661;
  reg        [15:0]   _zz_1662;
  reg        [15:0]   _zz_1663;
  reg        [15:0]   _zz_1664;
  reg        [15:0]   _zz_1665;
  reg        [15:0]   _zz_1666;
  reg        [15:0]   _zz_1667;
  reg        [15:0]   _zz_1668;
  reg        [15:0]   _zz_1669;
  reg        [15:0]   _zz_1670;
  reg        [15:0]   _zz_1671;
  reg        [15:0]   _zz_1672;
  reg        [15:0]   _zz_1673;
  reg        [15:0]   _zz_1674;
  reg        [15:0]   _zz_1675;
  reg        [15:0]   _zz_1676;
  reg        [15:0]   _zz_1677;
  reg        [15:0]   _zz_1678;
  reg        [15:0]   _zz_1679;
  reg        [15:0]   _zz_1680;
  reg        [15:0]   _zz_1681;
  reg        [15:0]   _zz_1682;
  reg        [15:0]   _zz_1683;
  reg        [15:0]   _zz_1684;
  reg        [15:0]   _zz_1685;
  reg        [15:0]   _zz_1686;
  reg        [15:0]   _zz_1687;
  reg        [15:0]   _zz_1688;
  reg        [15:0]   _zz_1689;
  reg        [15:0]   _zz_1690;
  reg        [15:0]   _zz_1691;
  reg        [15:0]   _zz_1692;
  reg        [15:0]   _zz_1693;
  reg        [15:0]   _zz_1694;
  reg        [15:0]   _zz_1695;
  reg        [15:0]   _zz_1696;
  reg        [15:0]   _zz_1697;
  reg        [15:0]   _zz_1698;
  reg        [15:0]   _zz_1699;
  reg        [15:0]   _zz_1700;
  reg        [15:0]   _zz_1701;
  reg        [15:0]   _zz_1702;
  reg        [15:0]   _zz_1703;
  reg        [15:0]   _zz_1704;
  reg        [15:0]   _zz_1705;
  reg        [15:0]   _zz_1706;
  reg        [15:0]   _zz_1707;
  reg        [15:0]   _zz_1708;
  reg        [15:0]   _zz_1709;
  reg        [15:0]   _zz_1710;
  reg        [15:0]   _zz_1711;
  reg        [15:0]   _zz_1712;
  reg        [15:0]   _zz_1713;
  reg        [15:0]   _zz_1714;
  reg        [15:0]   _zz_1715;
  reg        [15:0]   _zz_1716;
  reg        [15:0]   _zz_1717;
  reg        [15:0]   _zz_1718;
  reg        [15:0]   _zz_1719;
  reg        [15:0]   _zz_1720;
  reg        [15:0]   _zz_1721;
  reg        [15:0]   _zz_1722;
  reg        [15:0]   _zz_1723;
  reg        [15:0]   _zz_1724;
  reg        [15:0]   _zz_1725;
  reg        [15:0]   _zz_1726;
  reg        [15:0]   _zz_1727;
  reg        [15:0]   _zz_1728;
  reg        [15:0]   _zz_1729;
  reg        [15:0]   _zz_1730;
  reg        [15:0]   _zz_1731;
  reg        [15:0]   _zz_1732;
  reg        [15:0]   _zz_1733;
  reg        [15:0]   _zz_1734;
  reg        [15:0]   _zz_1735;
  reg        [15:0]   _zz_1736;
  reg        [15:0]   _zz_1737;
  reg        [15:0]   _zz_1738;
  reg        [15:0]   _zz_1739;
  reg        [15:0]   _zz_1740;
  reg        [15:0]   _zz_1741;
  reg        [15:0]   _zz_1742;
  reg        [15:0]   _zz_1743;
  reg        [15:0]   _zz_1744;
  reg        [15:0]   _zz_1745;
  reg        [15:0]   _zz_1746;
  reg        [15:0]   _zz_1747;
  reg        [15:0]   _zz_1748;
  reg        [15:0]   _zz_1749;
  reg        [15:0]   _zz_1750;
  reg        [15:0]   _zz_1751;
  reg        [15:0]   _zz_1752;
  reg        [15:0]   _zz_1753;
  reg        [15:0]   _zz_1754;
  reg        [15:0]   _zz_1755;
  reg        [15:0]   _zz_1756;
  reg        [15:0]   _zz_1757;
  reg        [15:0]   _zz_1758;
  reg        [15:0]   _zz_1759;
  reg        [15:0]   _zz_1760;
  reg        [15:0]   _zz_1761;
  reg        [15:0]   _zz_1762;
  reg        [15:0]   _zz_1763;
  reg        [15:0]   _zz_1764;
  reg        [15:0]   _zz_1765;
  reg        [15:0]   _zz_1766;
  reg        [15:0]   _zz_1767;
  reg        [15:0]   _zz_1768;
  reg        [15:0]   _zz_1769;
  reg        [15:0]   _zz_1770;
  reg        [15:0]   _zz_1771;
  reg        [15:0]   _zz_1772;
  reg        [15:0]   _zz_1773;
  reg        [15:0]   _zz_1774;
  reg        [15:0]   _zz_1775;
  reg        [15:0]   _zz_1776;
  reg        [15:0]   _zz_1777;
  reg        [15:0]   _zz_1778;
  reg        [15:0]   _zz_1779;
  reg        [15:0]   _zz_1780;
  reg        [15:0]   _zz_1781;
  reg        [15:0]   _zz_1782;
  reg        [15:0]   _zz_1783;
  reg        [15:0]   _zz_1784;
  reg        [15:0]   _zz_1785;
  reg        [15:0]   _zz_1786;
  reg        [15:0]   _zz_1787;
  reg        [15:0]   _zz_1788;
  reg        [15:0]   _zz_1789;
  reg        [15:0]   _zz_1790;
  reg        [15:0]   _zz_1791;
  reg        [15:0]   _zz_1792;
  wire       [15:0]   _zz_1793;
  wire       [15:0]   _zz_1794;
  wire       [15:0]   _zz_1795;
  wire       [0:0]    _zz_1796;
  wire       [0:0]    _zz_1797;
  wire       [15:0]   _zz_1798;
  wire       [15:0]   _zz_1799;
  wire       [15:0]   _zz_1800;
  wire       [0:0]    _zz_1801;
  wire       [0:0]    _zz_1802;
  wire       [15:0]   _zz_1803;
  wire       [15:0]   _zz_1804;
  wire       [15:0]   _zz_1805;
  wire       [0:0]    _zz_1806;
  wire       [0:0]    _zz_1807;
  wire       [15:0]   _zz_1808;
  wire       [15:0]   _zz_1809;
  wire       [15:0]   _zz_1810;
  wire       [0:0]    _zz_1811;
  wire       [0:0]    _zz_1812;
  wire       [15:0]   _zz_1813;
  wire       [15:0]   _zz_1814;
  wire       [15:0]   _zz_1815;
  wire       [0:0]    _zz_1816;
  wire       [0:0]    _zz_1817;
  wire       [15:0]   _zz_1818;
  wire       [15:0]   _zz_1819;
  wire       [15:0]   _zz_1820;
  wire       [0:0]    _zz_1821;
  wire       [0:0]    _zz_1822;
  wire       [15:0]   _zz_1823;
  wire       [15:0]   _zz_1824;
  wire       [15:0]   _zz_1825;
  wire       [0:0]    _zz_1826;
  wire       [0:0]    _zz_1827;
  wire       [15:0]   _zz_1828;
  wire       [15:0]   _zz_1829;
  wire       [15:0]   _zz_1830;
  wire       [0:0]    _zz_1831;
  wire       [0:0]    _zz_1832;
  wire       [15:0]   _zz_1833;
  wire       [15:0]   _zz_1834;
  wire       [15:0]   _zz_1835;
  wire       [0:0]    _zz_1836;
  wire       [0:0]    _zz_1837;
  wire       [15:0]   _zz_1838;
  wire       [15:0]   _zz_1839;
  wire       [15:0]   _zz_1840;
  wire       [0:0]    _zz_1841;
  wire       [0:0]    _zz_1842;
  wire       [15:0]   _zz_1843;
  wire       [15:0]   _zz_1844;
  wire       [15:0]   _zz_1845;
  wire       [0:0]    _zz_1846;
  wire       [0:0]    _zz_1847;
  wire       [15:0]   _zz_1848;
  wire       [15:0]   _zz_1849;
  wire       [15:0]   _zz_1850;
  wire       [0:0]    _zz_1851;
  wire       [0:0]    _zz_1852;
  wire       [15:0]   _zz_1853;
  wire       [15:0]   _zz_1854;
  wire       [15:0]   _zz_1855;
  wire       [0:0]    _zz_1856;
  wire       [0:0]    _zz_1857;
  wire       [15:0]   _zz_1858;
  wire       [15:0]   _zz_1859;
  wire       [15:0]   _zz_1860;
  wire       [0:0]    _zz_1861;
  wire       [0:0]    _zz_1862;
  wire       [15:0]   _zz_1863;
  wire       [15:0]   _zz_1864;
  wire       [15:0]   _zz_1865;
  wire       [0:0]    _zz_1866;
  wire       [0:0]    _zz_1867;
  wire       [15:0]   _zz_1868;
  wire       [15:0]   _zz_1869;
  wire       [15:0]   _zz_1870;
  wire       [0:0]    _zz_1871;
  wire       [0:0]    _zz_1872;
  wire       [15:0]   _zz_1873;
  wire       [15:0]   _zz_1874;
  wire       [15:0]   _zz_1875;
  wire       [0:0]    _zz_1876;
  wire       [0:0]    _zz_1877;
  wire       [15:0]   _zz_1878;
  wire       [15:0]   _zz_1879;
  wire       [15:0]   _zz_1880;
  wire       [0:0]    _zz_1881;
  wire       [0:0]    _zz_1882;
  wire       [15:0]   _zz_1883;
  wire       [15:0]   _zz_1884;
  wire       [15:0]   _zz_1885;
  wire       [0:0]    _zz_1886;
  wire       [0:0]    _zz_1887;
  wire       [15:0]   _zz_1888;
  wire       [15:0]   _zz_1889;
  wire       [15:0]   _zz_1890;
  wire       [0:0]    _zz_1891;
  wire       [0:0]    _zz_1892;
  wire       [15:0]   _zz_1893;
  wire       [15:0]   _zz_1894;
  wire       [15:0]   _zz_1895;
  wire       [0:0]    _zz_1896;
  wire       [0:0]    _zz_1897;
  wire       [15:0]   _zz_1898;
  wire       [15:0]   _zz_1899;
  wire       [15:0]   _zz_1900;
  wire       [0:0]    _zz_1901;
  wire       [0:0]    _zz_1902;
  wire       [15:0]   _zz_1903;
  wire       [15:0]   _zz_1904;
  wire       [15:0]   _zz_1905;
  wire       [0:0]    _zz_1906;
  wire       [0:0]    _zz_1907;
  wire       [15:0]   _zz_1908;
  wire       [15:0]   _zz_1909;
  wire       [15:0]   _zz_1910;
  wire       [0:0]    _zz_1911;
  wire       [0:0]    _zz_1912;
  wire       [15:0]   _zz_1913;
  wire       [15:0]   _zz_1914;
  wire       [15:0]   _zz_1915;
  wire       [0:0]    _zz_1916;
  wire       [0:0]    _zz_1917;
  wire       [15:0]   _zz_1918;
  wire       [15:0]   _zz_1919;
  wire       [15:0]   _zz_1920;
  wire       [0:0]    _zz_1921;
  wire       [0:0]    _zz_1922;
  wire       [15:0]   _zz_1923;
  wire       [15:0]   _zz_1924;
  wire       [15:0]   _zz_1925;
  wire       [0:0]    _zz_1926;
  wire       [0:0]    _zz_1927;
  wire       [15:0]   _zz_1928;
  wire       [15:0]   _zz_1929;
  wire       [15:0]   _zz_1930;
  wire       [0:0]    _zz_1931;
  wire       [0:0]    _zz_1932;
  wire       [15:0]   _zz_1933;
  wire       [15:0]   _zz_1934;
  wire       [15:0]   _zz_1935;
  wire       [0:0]    _zz_1936;
  wire       [0:0]    _zz_1937;
  wire       [15:0]   _zz_1938;
  wire       [15:0]   _zz_1939;
  wire       [15:0]   _zz_1940;
  wire       [0:0]    _zz_1941;
  wire       [0:0]    _zz_1942;
  wire       [15:0]   _zz_1943;
  wire       [15:0]   _zz_1944;
  wire       [15:0]   _zz_1945;
  wire       [0:0]    _zz_1946;
  wire       [0:0]    _zz_1947;
  wire       [15:0]   _zz_1948;
  wire       [15:0]   _zz_1949;
  wire       [15:0]   _zz_1950;
  wire       [0:0]    _zz_1951;
  wire       [0:0]    _zz_1952;
  wire       [15:0]   _zz_1953;
  wire       [15:0]   _zz_1954;
  wire       [15:0]   _zz_1955;
  wire       [0:0]    _zz_1956;
  wire       [0:0]    _zz_1957;
  wire       [15:0]   _zz_1958;
  wire       [15:0]   _zz_1959;
  wire       [15:0]   _zz_1960;
  wire       [0:0]    _zz_1961;
  wire       [0:0]    _zz_1962;
  wire       [15:0]   _zz_1963;
  wire       [15:0]   _zz_1964;
  wire       [15:0]   _zz_1965;
  wire       [0:0]    _zz_1966;
  wire       [0:0]    _zz_1967;
  wire       [15:0]   _zz_1968;
  wire       [15:0]   _zz_1969;
  wire       [15:0]   _zz_1970;
  wire       [0:0]    _zz_1971;
  wire       [0:0]    _zz_1972;
  wire       [15:0]   _zz_1973;
  wire       [15:0]   _zz_1974;
  wire       [15:0]   _zz_1975;
  wire       [0:0]    _zz_1976;
  wire       [0:0]    _zz_1977;
  wire       [15:0]   _zz_1978;
  wire       [15:0]   _zz_1979;
  wire       [15:0]   _zz_1980;
  wire       [0:0]    _zz_1981;
  wire       [0:0]    _zz_1982;
  wire       [15:0]   _zz_1983;
  wire       [15:0]   _zz_1984;
  wire       [15:0]   _zz_1985;
  wire       [0:0]    _zz_1986;
  wire       [0:0]    _zz_1987;
  wire       [15:0]   _zz_1988;
  wire       [15:0]   _zz_1989;
  wire       [15:0]   _zz_1990;
  wire       [0:0]    _zz_1991;
  wire       [0:0]    _zz_1992;
  wire       [15:0]   _zz_1993;
  wire       [15:0]   _zz_1994;
  wire       [15:0]   _zz_1995;
  wire       [0:0]    _zz_1996;
  wire       [0:0]    _zz_1997;
  wire       [15:0]   _zz_1998;
  wire       [15:0]   _zz_1999;
  wire       [15:0]   _zz_2000;
  wire       [0:0]    _zz_2001;
  wire       [0:0]    _zz_2002;
  wire       [15:0]   _zz_2003;
  wire       [15:0]   _zz_2004;
  wire       [15:0]   _zz_2005;
  wire       [0:0]    _zz_2006;
  wire       [0:0]    _zz_2007;
  wire       [15:0]   _zz_2008;
  wire       [15:0]   _zz_2009;
  wire       [15:0]   _zz_2010;
  wire       [0:0]    _zz_2011;
  wire       [0:0]    _zz_2012;
  wire       [15:0]   _zz_2013;
  wire       [15:0]   _zz_2014;
  wire       [15:0]   _zz_2015;
  wire       [0:0]    _zz_2016;
  wire       [0:0]    _zz_2017;
  wire       [15:0]   _zz_2018;
  wire       [15:0]   _zz_2019;
  wire       [15:0]   _zz_2020;
  wire       [0:0]    _zz_2021;
  wire       [0:0]    _zz_2022;
  wire       [15:0]   _zz_2023;
  wire       [15:0]   _zz_2024;
  wire       [15:0]   _zz_2025;
  wire       [0:0]    _zz_2026;
  wire       [0:0]    _zz_2027;
  wire       [15:0]   _zz_2028;
  wire       [15:0]   _zz_2029;
  wire       [15:0]   _zz_2030;
  wire       [0:0]    _zz_2031;
  wire       [0:0]    _zz_2032;
  wire       [15:0]   _zz_2033;
  wire       [15:0]   _zz_2034;
  wire       [15:0]   _zz_2035;
  wire       [0:0]    _zz_2036;
  wire       [0:0]    _zz_2037;
  wire       [15:0]   _zz_2038;
  wire       [15:0]   _zz_2039;
  wire       [15:0]   _zz_2040;
  wire       [0:0]    _zz_2041;
  wire       [0:0]    _zz_2042;
  wire       [15:0]   _zz_2043;
  wire       [15:0]   _zz_2044;
  wire       [15:0]   _zz_2045;
  wire       [0:0]    _zz_2046;
  wire       [0:0]    _zz_2047;
  wire       [15:0]   _zz_2048;
  wire       [15:0]   _zz_2049;
  wire       [15:0]   _zz_2050;
  wire       [0:0]    _zz_2051;
  wire       [0:0]    _zz_2052;
  wire       [15:0]   _zz_2053;
  wire       [15:0]   _zz_2054;
  wire       [15:0]   _zz_2055;
  wire       [0:0]    _zz_2056;
  wire       [0:0]    _zz_2057;
  wire       [15:0]   _zz_2058;
  wire       [15:0]   _zz_2059;
  wire       [15:0]   _zz_2060;
  wire       [0:0]    _zz_2061;
  wire       [0:0]    _zz_2062;
  wire       [15:0]   _zz_2063;
  wire       [15:0]   _zz_2064;
  wire       [15:0]   _zz_2065;
  wire       [0:0]    _zz_2066;
  wire       [0:0]    _zz_2067;
  wire       [15:0]   _zz_2068;
  wire       [15:0]   _zz_2069;
  wire       [15:0]   _zz_2070;
  wire       [0:0]    _zz_2071;
  wire       [0:0]    _zz_2072;
  wire       [15:0]   _zz_2073;
  wire       [15:0]   _zz_2074;
  wire       [15:0]   _zz_2075;
  wire       [0:0]    _zz_2076;
  wire       [0:0]    _zz_2077;
  wire       [15:0]   _zz_2078;
  wire       [15:0]   _zz_2079;
  wire       [15:0]   _zz_2080;
  wire       [0:0]    _zz_2081;
  wire       [0:0]    _zz_2082;
  wire       [15:0]   _zz_2083;
  wire       [15:0]   _zz_2084;
  wire       [15:0]   _zz_2085;
  wire       [0:0]    _zz_2086;
  wire       [0:0]    _zz_2087;
  wire       [15:0]   _zz_2088;
  wire       [15:0]   _zz_2089;
  wire       [15:0]   _zz_2090;
  wire       [0:0]    _zz_2091;
  wire       [0:0]    _zz_2092;
  wire       [15:0]   _zz_2093;
  wire       [15:0]   _zz_2094;
  wire       [15:0]   _zz_2095;
  wire       [0:0]    _zz_2096;
  wire       [0:0]    _zz_2097;
  wire       [15:0]   _zz_2098;
  wire       [15:0]   _zz_2099;
  wire       [15:0]   _zz_2100;
  wire       [0:0]    _zz_2101;
  wire       [0:0]    _zz_2102;
  wire       [15:0]   _zz_2103;
  wire       [15:0]   _zz_2104;
  wire       [15:0]   _zz_2105;
  wire       [0:0]    _zz_2106;
  wire       [0:0]    _zz_2107;
  wire       [15:0]   _zz_2108;
  wire       [15:0]   _zz_2109;
  wire       [15:0]   _zz_2110;
  wire       [0:0]    _zz_2111;
  wire       [0:0]    _zz_2112;
  wire       [15:0]   _zz_2113;
  wire       [15:0]   _zz_2114;
  wire       [15:0]   _zz_2115;
  wire       [0:0]    _zz_2116;
  wire       [0:0]    _zz_2117;
  wire       [15:0]   _zz_2118;
  wire       [15:0]   _zz_2119;
  wire       [15:0]   _zz_2120;
  wire       [0:0]    _zz_2121;
  wire       [0:0]    _zz_2122;
  wire       [15:0]   _zz_2123;
  wire       [15:0]   _zz_2124;
  wire       [15:0]   _zz_2125;
  wire       [0:0]    _zz_2126;
  wire       [0:0]    _zz_2127;
  wire       [15:0]   _zz_2128;
  wire       [15:0]   _zz_2129;
  wire       [15:0]   _zz_2130;
  wire       [0:0]    _zz_2131;
  wire       [0:0]    _zz_2132;
  wire       [15:0]   _zz_2133;
  wire       [15:0]   _zz_2134;
  wire       [15:0]   _zz_2135;
  wire       [0:0]    _zz_2136;
  wire       [0:0]    _zz_2137;
  wire       [15:0]   _zz_2138;
  wire       [15:0]   _zz_2139;
  wire       [15:0]   _zz_2140;
  wire       [0:0]    _zz_2141;
  wire       [0:0]    _zz_2142;
  wire       [15:0]   _zz_2143;
  wire       [15:0]   _zz_2144;
  wire       [15:0]   _zz_2145;
  wire       [0:0]    _zz_2146;
  wire       [0:0]    _zz_2147;
  wire       [15:0]   _zz_2148;
  wire       [15:0]   _zz_2149;
  wire       [15:0]   _zz_2150;
  wire       [0:0]    _zz_2151;
  wire       [0:0]    _zz_2152;
  wire       [15:0]   _zz_2153;
  wire       [15:0]   _zz_2154;
  wire       [15:0]   _zz_2155;
  wire       [0:0]    _zz_2156;
  wire       [0:0]    _zz_2157;
  wire       [15:0]   _zz_2158;
  wire       [15:0]   _zz_2159;
  wire       [15:0]   _zz_2160;
  wire       [0:0]    _zz_2161;
  wire       [0:0]    _zz_2162;
  wire       [15:0]   _zz_2163;
  wire       [15:0]   _zz_2164;
  wire       [15:0]   _zz_2165;
  wire       [0:0]    _zz_2166;
  wire       [0:0]    _zz_2167;
  wire       [15:0]   _zz_2168;
  wire       [15:0]   _zz_2169;
  wire       [15:0]   _zz_2170;
  wire       [0:0]    _zz_2171;
  wire       [0:0]    _zz_2172;
  wire       [15:0]   _zz_2173;
  wire       [15:0]   _zz_2174;
  wire       [15:0]   _zz_2175;
  wire       [0:0]    _zz_2176;
  wire       [0:0]    _zz_2177;
  wire       [15:0]   _zz_2178;
  wire       [15:0]   _zz_2179;
  wire       [15:0]   _zz_2180;
  wire       [0:0]    _zz_2181;
  wire       [0:0]    _zz_2182;
  wire       [15:0]   _zz_2183;
  wire       [15:0]   _zz_2184;
  wire       [15:0]   _zz_2185;
  wire       [0:0]    _zz_2186;
  wire       [0:0]    _zz_2187;
  wire       [15:0]   _zz_2188;
  wire       [15:0]   _zz_2189;
  wire       [15:0]   _zz_2190;
  wire       [0:0]    _zz_2191;
  wire       [0:0]    _zz_2192;
  wire       [15:0]   _zz_2193;
  wire       [15:0]   _zz_2194;
  wire       [15:0]   _zz_2195;
  wire       [0:0]    _zz_2196;
  wire       [0:0]    _zz_2197;
  wire       [15:0]   _zz_2198;
  wire       [15:0]   _zz_2199;
  wire       [15:0]   _zz_2200;
  wire       [0:0]    _zz_2201;
  wire       [0:0]    _zz_2202;
  wire       [15:0]   _zz_2203;
  wire       [15:0]   _zz_2204;
  wire       [15:0]   _zz_2205;
  wire       [0:0]    _zz_2206;
  wire       [0:0]    _zz_2207;
  wire       [15:0]   _zz_2208;
  wire       [15:0]   _zz_2209;
  wire       [15:0]   _zz_2210;
  wire       [0:0]    _zz_2211;
  wire       [0:0]    _zz_2212;
  wire       [15:0]   _zz_2213;
  wire       [15:0]   _zz_2214;
  wire       [15:0]   _zz_2215;
  wire       [0:0]    _zz_2216;
  wire       [0:0]    _zz_2217;
  wire       [15:0]   _zz_2218;
  wire       [15:0]   _zz_2219;
  wire       [15:0]   _zz_2220;
  wire       [0:0]    _zz_2221;
  wire       [0:0]    _zz_2222;
  wire       [15:0]   _zz_2223;
  wire       [15:0]   _zz_2224;
  wire       [15:0]   _zz_2225;
  wire       [0:0]    _zz_2226;
  wire       [0:0]    _zz_2227;
  wire       [15:0]   _zz_2228;
  wire       [15:0]   _zz_2229;
  wire       [15:0]   _zz_2230;
  wire       [0:0]    _zz_2231;
  wire       [0:0]    _zz_2232;
  wire       [15:0]   _zz_2233;
  wire       [15:0]   _zz_2234;
  wire       [15:0]   _zz_2235;
  wire       [0:0]    _zz_2236;
  wire       [0:0]    _zz_2237;
  wire       [15:0]   _zz_2238;
  wire       [15:0]   _zz_2239;
  wire       [15:0]   _zz_2240;
  wire       [0:0]    _zz_2241;
  wire       [0:0]    _zz_2242;
  wire       [15:0]   _zz_2243;
  wire       [15:0]   _zz_2244;
  wire       [15:0]   _zz_2245;
  wire       [0:0]    _zz_2246;
  wire       [0:0]    _zz_2247;
  wire       [15:0]   _zz_2248;
  wire       [15:0]   _zz_2249;
  wire       [15:0]   _zz_2250;
  wire       [0:0]    _zz_2251;
  wire       [0:0]    _zz_2252;
  wire       [15:0]   _zz_2253;
  wire       [15:0]   _zz_2254;
  wire       [15:0]   _zz_2255;
  wire       [0:0]    _zz_2256;
  wire       [0:0]    _zz_2257;
  wire       [15:0]   _zz_2258;
  wire       [15:0]   _zz_2259;
  wire       [15:0]   _zz_2260;
  wire       [0:0]    _zz_2261;
  wire       [0:0]    _zz_2262;
  wire       [15:0]   _zz_2263;
  wire       [15:0]   _zz_2264;
  wire       [15:0]   _zz_2265;
  wire       [0:0]    _zz_2266;
  wire       [0:0]    _zz_2267;
  wire       [15:0]   _zz_2268;
  wire       [15:0]   _zz_2269;
  wire       [15:0]   _zz_2270;
  wire       [0:0]    _zz_2271;
  wire       [0:0]    _zz_2272;
  wire       [15:0]   _zz_2273;
  wire       [15:0]   _zz_2274;
  wire       [15:0]   _zz_2275;
  wire       [0:0]    _zz_2276;
  wire       [0:0]    _zz_2277;
  wire       [15:0]   _zz_2278;
  wire       [15:0]   _zz_2279;
  wire       [15:0]   _zz_2280;
  wire       [0:0]    _zz_2281;
  wire       [0:0]    _zz_2282;
  wire       [15:0]   _zz_2283;
  wire       [15:0]   _zz_2284;
  wire       [15:0]   _zz_2285;
  wire       [0:0]    _zz_2286;
  wire       [0:0]    _zz_2287;
  wire       [15:0]   _zz_2288;
  wire       [15:0]   _zz_2289;
  wire       [15:0]   _zz_2290;
  wire       [0:0]    _zz_2291;
  wire       [0:0]    _zz_2292;
  wire       [15:0]   _zz_2293;
  wire       [15:0]   _zz_2294;
  wire       [15:0]   _zz_2295;
  wire       [0:0]    _zz_2296;
  wire       [0:0]    _zz_2297;
  wire       [15:0]   _zz_2298;
  wire       [15:0]   _zz_2299;
  wire       [15:0]   _zz_2300;
  wire       [0:0]    _zz_2301;
  wire       [0:0]    _zz_2302;
  wire       [15:0]   _zz_2303;
  wire       [15:0]   _zz_2304;
  wire       [15:0]   _zz_2305;
  wire       [0:0]    _zz_2306;
  wire       [0:0]    _zz_2307;
  wire       [15:0]   _zz_2308;
  wire       [15:0]   _zz_2309;
  wire       [15:0]   _zz_2310;
  wire       [0:0]    _zz_2311;
  wire       [0:0]    _zz_2312;
  wire       [15:0]   _zz_2313;
  wire       [15:0]   _zz_2314;
  wire       [15:0]   _zz_2315;
  wire       [0:0]    _zz_2316;
  wire       [0:0]    _zz_2317;
  wire       [15:0]   _zz_2318;
  wire       [15:0]   _zz_2319;
  wire       [15:0]   _zz_2320;
  wire       [0:0]    _zz_2321;
  wire       [0:0]    _zz_2322;
  wire       [15:0]   _zz_2323;
  wire       [15:0]   _zz_2324;
  wire       [15:0]   _zz_2325;
  wire       [0:0]    _zz_2326;
  wire       [0:0]    _zz_2327;
  wire       [15:0]   _zz_2328;
  wire       [15:0]   _zz_2329;
  wire       [15:0]   _zz_2330;
  wire       [0:0]    _zz_2331;
  wire       [0:0]    _zz_2332;
  wire       [15:0]   _zz_2333;
  wire       [15:0]   _zz_2334;
  wire       [15:0]   _zz_2335;
  wire       [0:0]    _zz_2336;
  wire       [0:0]    _zz_2337;
  wire       [15:0]   _zz_2338;
  wire       [15:0]   _zz_2339;
  wire       [15:0]   _zz_2340;
  wire       [0:0]    _zz_2341;
  wire       [0:0]    _zz_2342;
  wire       [15:0]   _zz_2343;
  wire       [15:0]   _zz_2344;
  wire       [15:0]   _zz_2345;
  wire       [0:0]    _zz_2346;
  wire       [0:0]    _zz_2347;
  wire       [15:0]   _zz_2348;
  wire       [15:0]   _zz_2349;
  wire       [15:0]   _zz_2350;
  wire       [0:0]    _zz_2351;
  wire       [0:0]    _zz_2352;
  wire       [15:0]   _zz_2353;
  wire       [15:0]   _zz_2354;
  wire       [15:0]   _zz_2355;
  wire       [0:0]    _zz_2356;
  wire       [0:0]    _zz_2357;
  wire       [15:0]   _zz_2358;
  wire       [15:0]   _zz_2359;
  wire       [15:0]   _zz_2360;
  wire       [0:0]    _zz_2361;
  wire       [0:0]    _zz_2362;
  wire       [15:0]   _zz_2363;
  wire       [15:0]   _zz_2364;
  wire       [15:0]   _zz_2365;
  wire       [0:0]    _zz_2366;
  wire       [0:0]    _zz_2367;
  wire       [15:0]   _zz_2368;
  wire       [15:0]   _zz_2369;
  wire       [15:0]   _zz_2370;
  wire       [0:0]    _zz_2371;
  wire       [0:0]    _zz_2372;
  wire       [15:0]   _zz_2373;
  wire       [15:0]   _zz_2374;
  wire       [15:0]   _zz_2375;
  wire       [0:0]    _zz_2376;
  wire       [0:0]    _zz_2377;
  wire       [15:0]   _zz_2378;
  wire       [15:0]   _zz_2379;
  wire       [15:0]   _zz_2380;
  wire       [0:0]    _zz_2381;
  wire       [0:0]    _zz_2382;
  wire       [15:0]   _zz_2383;
  wire       [15:0]   _zz_2384;
  wire       [15:0]   _zz_2385;
  wire       [0:0]    _zz_2386;
  wire       [0:0]    _zz_2387;
  wire       [15:0]   _zz_2388;
  wire       [15:0]   _zz_2389;
  wire       [15:0]   _zz_2390;
  wire       [0:0]    _zz_2391;
  wire       [0:0]    _zz_2392;
  wire       [15:0]   _zz_2393;
  wire       [15:0]   _zz_2394;
  wire       [15:0]   _zz_2395;
  wire       [0:0]    _zz_2396;
  wire       [0:0]    _zz_2397;
  wire       [15:0]   _zz_2398;
  wire       [15:0]   _zz_2399;
  wire       [15:0]   _zz_2400;
  wire       [0:0]    _zz_2401;
  wire       [0:0]    _zz_2402;
  wire       [15:0]   _zz_2403;
  wire       [15:0]   _zz_2404;
  wire       [15:0]   _zz_2405;
  wire       [0:0]    _zz_2406;
  wire       [0:0]    _zz_2407;
  wire       [15:0]   _zz_2408;
  wire       [15:0]   _zz_2409;
  wire       [15:0]   _zz_2410;
  wire       [0:0]    _zz_2411;
  wire       [0:0]    _zz_2412;
  wire       [15:0]   _zz_2413;
  wire       [15:0]   _zz_2414;
  wire       [15:0]   _zz_2415;
  wire       [0:0]    _zz_2416;
  wire       [0:0]    _zz_2417;
  wire       [15:0]   _zz_2418;
  wire       [15:0]   _zz_2419;
  wire       [15:0]   _zz_2420;
  wire       [0:0]    _zz_2421;
  wire       [0:0]    _zz_2422;
  wire       [15:0]   _zz_2423;
  wire       [15:0]   _zz_2424;
  wire       [15:0]   _zz_2425;
  wire       [0:0]    _zz_2426;
  wire       [0:0]    _zz_2427;
  wire       [15:0]   _zz_2428;
  wire       [15:0]   _zz_2429;
  wire       [15:0]   _zz_2430;
  wire       [0:0]    _zz_2431;
  wire       [0:0]    _zz_2432;
  wire       [15:0]   _zz_2433;
  wire       [15:0]   _zz_2434;
  wire       [15:0]   _zz_2435;
  wire       [0:0]    _zz_2436;
  wire       [0:0]    _zz_2437;
  wire       [15:0]   _zz_2438;
  wire       [15:0]   _zz_2439;
  wire       [15:0]   _zz_2440;
  wire       [0:0]    _zz_2441;
  wire       [0:0]    _zz_2442;
  wire       [15:0]   _zz_2443;
  wire       [15:0]   _zz_2444;
  wire       [15:0]   _zz_2445;
  wire       [0:0]    _zz_2446;
  wire       [0:0]    _zz_2447;
  wire       [15:0]   _zz_2448;
  wire       [15:0]   _zz_2449;
  wire       [15:0]   _zz_2450;
  wire       [0:0]    _zz_2451;
  wire       [0:0]    _zz_2452;
  wire       [15:0]   _zz_2453;
  wire       [15:0]   _zz_2454;
  wire       [15:0]   _zz_2455;
  wire       [0:0]    _zz_2456;
  wire       [0:0]    _zz_2457;
  wire       [15:0]   _zz_2458;
  wire       [15:0]   _zz_2459;
  wire       [15:0]   _zz_2460;
  wire       [0:0]    _zz_2461;
  wire       [0:0]    _zz_2462;
  wire       [15:0]   _zz_2463;
  wire       [15:0]   _zz_2464;
  wire       [15:0]   _zz_2465;
  wire       [0:0]    _zz_2466;
  wire       [0:0]    _zz_2467;
  wire       [15:0]   _zz_2468;
  wire       [15:0]   _zz_2469;
  wire       [15:0]   _zz_2470;
  wire       [0:0]    _zz_2471;
  wire       [0:0]    _zz_2472;
  wire       [15:0]   _zz_2473;
  wire       [15:0]   _zz_2474;
  wire       [15:0]   _zz_2475;
  wire       [0:0]    _zz_2476;
  wire       [0:0]    _zz_2477;
  wire       [15:0]   _zz_2478;
  wire       [15:0]   _zz_2479;
  wire       [15:0]   _zz_2480;
  wire       [0:0]    _zz_2481;
  wire       [0:0]    _zz_2482;
  wire       [15:0]   _zz_2483;
  wire       [15:0]   _zz_2484;
  wire       [15:0]   _zz_2485;
  wire       [0:0]    _zz_2486;
  wire       [0:0]    _zz_2487;
  wire       [15:0]   _zz_2488;
  wire       [15:0]   _zz_2489;
  wire       [15:0]   _zz_2490;
  wire       [0:0]    _zz_2491;
  wire       [0:0]    _zz_2492;
  wire       [15:0]   _zz_2493;
  wire       [15:0]   _zz_2494;
  wire       [15:0]   _zz_2495;
  wire       [0:0]    _zz_2496;
  wire       [0:0]    _zz_2497;
  wire       [15:0]   _zz_2498;
  wire       [15:0]   _zz_2499;
  wire       [15:0]   _zz_2500;
  wire       [0:0]    _zz_2501;
  wire       [0:0]    _zz_2502;
  wire       [15:0]   _zz_2503;
  wire       [15:0]   _zz_2504;
  wire       [15:0]   _zz_2505;
  wire       [0:0]    _zz_2506;
  wire       [0:0]    _zz_2507;
  wire       [15:0]   _zz_2508;
  wire       [15:0]   _zz_2509;
  wire       [15:0]   _zz_2510;
  wire       [0:0]    _zz_2511;
  wire       [0:0]    _zz_2512;
  wire       [15:0]   _zz_2513;
  wire       [15:0]   _zz_2514;
  wire       [15:0]   _zz_2515;
  wire       [0:0]    _zz_2516;
  wire       [0:0]    _zz_2517;
  wire       [15:0]   _zz_2518;
  wire       [15:0]   _zz_2519;
  wire       [15:0]   _zz_2520;
  wire       [0:0]    _zz_2521;
  wire       [0:0]    _zz_2522;
  wire       [15:0]   _zz_2523;
  wire       [15:0]   _zz_2524;
  wire       [15:0]   _zz_2525;
  wire       [0:0]    _zz_2526;
  wire       [0:0]    _zz_2527;
  wire       [15:0]   _zz_2528;
  wire       [15:0]   _zz_2529;
  wire       [15:0]   _zz_2530;
  wire       [0:0]    _zz_2531;
  wire       [0:0]    _zz_2532;
  wire       [15:0]   _zz_2533;
  wire       [15:0]   _zz_2534;
  wire       [15:0]   _zz_2535;
  wire       [0:0]    _zz_2536;
  wire       [0:0]    _zz_2537;
  wire       [15:0]   _zz_2538;
  wire       [15:0]   _zz_2539;
  wire       [15:0]   _zz_2540;
  wire       [0:0]    _zz_2541;
  wire       [0:0]    _zz_2542;
  wire       [15:0]   _zz_2543;
  wire       [15:0]   _zz_2544;
  wire       [15:0]   _zz_2545;
  wire       [0:0]    _zz_2546;
  wire       [0:0]    _zz_2547;
  wire       [15:0]   _zz_2548;
  wire       [15:0]   _zz_2549;
  wire       [15:0]   _zz_2550;
  wire       [0:0]    _zz_2551;
  wire       [0:0]    _zz_2552;
  wire       [15:0]   _zz_2553;
  wire       [15:0]   _zz_2554;
  wire       [15:0]   _zz_2555;
  wire       [0:0]    _zz_2556;
  wire       [0:0]    _zz_2557;
  wire       [15:0]   _zz_2558;
  wire       [15:0]   _zz_2559;
  wire       [15:0]   _zz_2560;
  wire       [0:0]    _zz_2561;
  wire       [0:0]    _zz_2562;
  wire       [15:0]   _zz_2563;
  wire       [15:0]   _zz_2564;
  wire       [15:0]   _zz_2565;
  wire       [0:0]    _zz_2566;
  wire       [0:0]    _zz_2567;
  wire       [15:0]   _zz_2568;
  wire       [15:0]   _zz_2569;
  wire       [15:0]   _zz_2570;
  wire       [0:0]    _zz_2571;
  wire       [0:0]    _zz_2572;
  wire       [15:0]   _zz_2573;
  wire       [15:0]   _zz_2574;
  wire       [15:0]   _zz_2575;
  wire       [0:0]    _zz_2576;
  wire       [0:0]    _zz_2577;
  wire       [15:0]   _zz_2578;
  wire       [15:0]   _zz_2579;
  wire       [15:0]   _zz_2580;
  wire       [0:0]    _zz_2581;
  wire       [0:0]    _zz_2582;
  wire       [15:0]   _zz_2583;
  wire       [15:0]   _zz_2584;
  wire       [15:0]   _zz_2585;
  wire       [0:0]    _zz_2586;
  wire       [0:0]    _zz_2587;
  wire       [15:0]   _zz_2588;
  wire       [15:0]   _zz_2589;
  wire       [15:0]   _zz_2590;
  wire       [0:0]    _zz_2591;
  wire       [0:0]    _zz_2592;
  wire       [15:0]   _zz_2593;
  wire       [15:0]   _zz_2594;
  wire       [15:0]   _zz_2595;
  wire       [0:0]    _zz_2596;
  wire       [0:0]    _zz_2597;
  wire       [15:0]   _zz_2598;
  wire       [15:0]   _zz_2599;
  wire       [15:0]   _zz_2600;
  wire       [0:0]    _zz_2601;
  wire       [0:0]    _zz_2602;
  wire       [15:0]   _zz_2603;
  wire       [15:0]   _zz_2604;
  wire       [15:0]   _zz_2605;
  wire       [0:0]    _zz_2606;
  wire       [0:0]    _zz_2607;
  wire       [15:0]   _zz_2608;
  wire       [15:0]   _zz_2609;
  wire       [15:0]   _zz_2610;
  wire       [0:0]    _zz_2611;
  wire       [0:0]    _zz_2612;
  wire       [15:0]   _zz_2613;
  wire       [15:0]   _zz_2614;
  wire       [15:0]   _zz_2615;
  wire       [0:0]    _zz_2616;
  wire       [0:0]    _zz_2617;
  wire       [15:0]   _zz_2618;
  wire       [15:0]   _zz_2619;
  wire       [15:0]   _zz_2620;
  wire       [0:0]    _zz_2621;
  wire       [0:0]    _zz_2622;
  wire       [15:0]   _zz_2623;
  wire       [15:0]   _zz_2624;
  wire       [15:0]   _zz_2625;
  wire       [0:0]    _zz_2626;
  wire       [0:0]    _zz_2627;
  wire       [15:0]   _zz_2628;
  wire       [15:0]   _zz_2629;
  wire       [15:0]   _zz_2630;
  wire       [0:0]    _zz_2631;
  wire       [0:0]    _zz_2632;
  wire       [15:0]   _zz_2633;
  wire       [15:0]   _zz_2634;
  wire       [15:0]   _zz_2635;
  wire       [0:0]    _zz_2636;
  wire       [0:0]    _zz_2637;
  wire       [15:0]   _zz_2638;
  wire       [15:0]   _zz_2639;
  wire       [15:0]   _zz_2640;
  wire       [0:0]    _zz_2641;
  wire       [0:0]    _zz_2642;
  wire       [15:0]   _zz_2643;
  wire       [15:0]   _zz_2644;
  wire       [15:0]   _zz_2645;
  wire       [0:0]    _zz_2646;
  wire       [0:0]    _zz_2647;
  wire       [15:0]   _zz_2648;
  wire       [15:0]   _zz_2649;
  wire       [15:0]   _zz_2650;
  wire       [0:0]    _zz_2651;
  wire       [0:0]    _zz_2652;
  wire       [15:0]   _zz_2653;
  wire       [15:0]   _zz_2654;
  wire       [15:0]   _zz_2655;
  wire       [0:0]    _zz_2656;
  wire       [0:0]    _zz_2657;
  wire       [15:0]   _zz_2658;
  wire       [15:0]   _zz_2659;
  wire       [15:0]   _zz_2660;
  wire       [0:0]    _zz_2661;
  wire       [0:0]    _zz_2662;
  wire       [15:0]   _zz_2663;
  wire       [15:0]   _zz_2664;
  wire       [15:0]   _zz_2665;
  wire       [0:0]    _zz_2666;
  wire       [0:0]    _zz_2667;
  wire       [15:0]   _zz_2668;
  wire       [15:0]   _zz_2669;
  wire       [15:0]   _zz_2670;
  wire       [0:0]    _zz_2671;
  wire       [0:0]    _zz_2672;
  wire       [15:0]   _zz_2673;
  wire       [15:0]   _zz_2674;
  wire       [15:0]   _zz_2675;
  wire       [0:0]    _zz_2676;
  wire       [0:0]    _zz_2677;
  wire       [15:0]   _zz_2678;
  wire       [15:0]   _zz_2679;
  wire       [15:0]   _zz_2680;
  wire       [0:0]    _zz_2681;
  wire       [0:0]    _zz_2682;
  wire       [15:0]   _zz_2683;
  wire       [15:0]   _zz_2684;
  wire       [15:0]   _zz_2685;
  wire       [0:0]    _zz_2686;
  wire       [0:0]    _zz_2687;
  wire       [15:0]   _zz_2688;
  wire       [15:0]   _zz_2689;
  wire       [15:0]   _zz_2690;
  wire       [0:0]    _zz_2691;
  wire       [0:0]    _zz_2692;
  wire       [15:0]   _zz_2693;
  wire       [15:0]   _zz_2694;
  wire       [15:0]   _zz_2695;
  wire       [0:0]    _zz_2696;
  wire       [0:0]    _zz_2697;
  wire       [15:0]   _zz_2698;
  wire       [15:0]   _zz_2699;
  wire       [15:0]   _zz_2700;
  wire       [0:0]    _zz_2701;
  wire       [0:0]    _zz_2702;
  wire       [15:0]   _zz_2703;
  wire       [15:0]   _zz_2704;
  wire       [15:0]   _zz_2705;
  wire       [0:0]    _zz_2706;
  wire       [0:0]    _zz_2707;
  wire       [15:0]   _zz_2708;
  wire       [15:0]   _zz_2709;
  wire       [15:0]   _zz_2710;
  wire       [0:0]    _zz_2711;
  wire       [0:0]    _zz_2712;
  wire       [15:0]   _zz_2713;
  wire       [15:0]   _zz_2714;
  wire       [15:0]   _zz_2715;
  wire       [0:0]    _zz_2716;
  wire       [0:0]    _zz_2717;
  wire       [15:0]   _zz_2718;
  wire       [15:0]   _zz_2719;
  wire       [15:0]   _zz_2720;
  wire       [0:0]    _zz_2721;
  wire       [0:0]    _zz_2722;
  wire       [15:0]   _zz_2723;
  wire       [15:0]   _zz_2724;
  wire       [15:0]   _zz_2725;
  wire       [0:0]    _zz_2726;
  wire       [0:0]    _zz_2727;
  wire       [15:0]   _zz_2728;
  wire       [15:0]   _zz_2729;
  wire       [15:0]   _zz_2730;
  wire       [0:0]    _zz_2731;
  wire       [0:0]    _zz_2732;
  wire       [15:0]   _zz_2733;
  wire       [15:0]   _zz_2734;
  wire       [15:0]   _zz_2735;
  wire       [0:0]    _zz_2736;
  wire       [0:0]    _zz_2737;
  wire       [15:0]   _zz_2738;
  wire       [15:0]   _zz_2739;
  wire       [15:0]   _zz_2740;
  wire       [0:0]    _zz_2741;
  wire       [0:0]    _zz_2742;
  wire       [15:0]   _zz_2743;
  wire       [15:0]   _zz_2744;
  wire       [15:0]   _zz_2745;
  wire       [0:0]    _zz_2746;
  wire       [0:0]    _zz_2747;
  wire       [15:0]   _zz_2748;
  wire       [15:0]   _zz_2749;
  wire       [15:0]   _zz_2750;
  wire       [0:0]    _zz_2751;
  wire       [0:0]    _zz_2752;
  wire       [15:0]   _zz_2753;
  wire       [15:0]   _zz_2754;
  wire       [15:0]   _zz_2755;
  wire       [0:0]    _zz_2756;
  wire       [0:0]    _zz_2757;
  wire       [15:0]   _zz_2758;
  wire       [15:0]   _zz_2759;
  wire       [15:0]   _zz_2760;
  wire       [0:0]    _zz_2761;
  wire       [0:0]    _zz_2762;
  wire       [15:0]   _zz_2763;
  wire       [15:0]   _zz_2764;
  wire       [15:0]   _zz_2765;
  wire       [0:0]    _zz_2766;
  wire       [0:0]    _zz_2767;
  wire       [15:0]   _zz_2768;
  wire       [15:0]   _zz_2769;
  wire       [15:0]   _zz_2770;
  wire       [0:0]    _zz_2771;
  wire       [0:0]    _zz_2772;
  wire       [15:0]   _zz_2773;
  wire       [15:0]   _zz_2774;
  wire       [15:0]   _zz_2775;
  wire       [0:0]    _zz_2776;
  wire       [0:0]    _zz_2777;
  wire       [15:0]   _zz_2778;
  wire       [15:0]   _zz_2779;
  wire       [15:0]   _zz_2780;
  wire       [0:0]    _zz_2781;
  wire       [0:0]    _zz_2782;
  wire       [15:0]   _zz_2783;
  wire       [15:0]   _zz_2784;
  wire       [15:0]   _zz_2785;
  wire       [0:0]    _zz_2786;
  wire       [0:0]    _zz_2787;
  wire       [15:0]   _zz_2788;
  wire       [15:0]   _zz_2789;
  wire       [15:0]   _zz_2790;
  wire       [0:0]    _zz_2791;
  wire       [0:0]    _zz_2792;
  wire       [15:0]   _zz_2793;
  wire       [15:0]   _zz_2794;
  wire       [15:0]   _zz_2795;
  wire       [0:0]    _zz_2796;
  wire       [0:0]    _zz_2797;
  wire       [15:0]   _zz_2798;
  wire       [15:0]   _zz_2799;
  wire       [15:0]   _zz_2800;
  wire       [0:0]    _zz_2801;
  wire       [0:0]    _zz_2802;
  wire       [15:0]   _zz_2803;
  wire       [15:0]   _zz_2804;
  wire       [15:0]   _zz_2805;
  wire       [0:0]    _zz_2806;
  wire       [0:0]    _zz_2807;
  wire       [15:0]   _zz_2808;
  wire       [15:0]   _zz_2809;
  wire       [15:0]   _zz_2810;
  wire       [0:0]    _zz_2811;
  wire       [0:0]    _zz_2812;
  wire       [15:0]   _zz_2813;
  wire       [15:0]   _zz_2814;
  wire       [15:0]   _zz_2815;
  wire       [0:0]    _zz_2816;
  wire       [0:0]    _zz_2817;
  wire       [15:0]   _zz_2818;
  wire       [15:0]   _zz_2819;
  wire       [15:0]   _zz_2820;
  wire       [0:0]    _zz_2821;
  wire       [0:0]    _zz_2822;
  wire       [15:0]   _zz_2823;
  wire       [15:0]   _zz_2824;
  wire       [15:0]   _zz_2825;
  wire       [0:0]    _zz_2826;
  wire       [0:0]    _zz_2827;
  wire       [15:0]   _zz_2828;
  wire       [15:0]   _zz_2829;
  wire       [15:0]   _zz_2830;
  wire       [0:0]    _zz_2831;
  wire       [0:0]    _zz_2832;
  wire       [15:0]   _zz_2833;
  wire       [15:0]   _zz_2834;
  wire       [15:0]   _zz_2835;
  wire       [0:0]    _zz_2836;
  wire       [0:0]    _zz_2837;
  wire       [15:0]   _zz_2838;
  wire       [15:0]   _zz_2839;
  wire       [15:0]   _zz_2840;
  wire       [0:0]    _zz_2841;
  wire       [0:0]    _zz_2842;
  wire       [15:0]   _zz_2843;
  wire       [15:0]   _zz_2844;
  wire       [15:0]   _zz_2845;
  wire       [0:0]    _zz_2846;
  wire       [0:0]    _zz_2847;
  wire       [15:0]   _zz_2848;
  wire       [15:0]   _zz_2849;
  wire       [15:0]   _zz_2850;
  wire       [0:0]    _zz_2851;
  wire       [0:0]    _zz_2852;
  wire       [15:0]   _zz_2853;
  wire       [15:0]   _zz_2854;
  wire       [15:0]   _zz_2855;
  wire       [0:0]    _zz_2856;
  wire       [0:0]    _zz_2857;
  wire       [15:0]   _zz_2858;
  wire       [15:0]   _zz_2859;
  wire       [15:0]   _zz_2860;
  wire       [0:0]    _zz_2861;
  wire       [0:0]    _zz_2862;
  wire       [15:0]   _zz_2863;
  wire       [15:0]   _zz_2864;
  wire       [15:0]   _zz_2865;
  wire       [0:0]    _zz_2866;
  wire       [0:0]    _zz_2867;
  wire       [15:0]   _zz_2868;
  wire       [15:0]   _zz_2869;
  wire       [15:0]   _zz_2870;
  wire       [0:0]    _zz_2871;
  wire       [0:0]    _zz_2872;
  wire       [15:0]   _zz_2873;
  wire       [15:0]   _zz_2874;
  wire       [15:0]   _zz_2875;
  wire       [0:0]    _zz_2876;
  wire       [0:0]    _zz_2877;
  wire       [15:0]   _zz_2878;
  wire       [15:0]   _zz_2879;
  wire       [15:0]   _zz_2880;
  wire       [0:0]    _zz_2881;
  wire       [0:0]    _zz_2882;
  wire       [15:0]   _zz_2883;
  wire       [15:0]   _zz_2884;
  wire       [15:0]   _zz_2885;
  wire       [0:0]    _zz_2886;
  wire       [0:0]    _zz_2887;
  wire       [15:0]   _zz_2888;
  wire       [15:0]   _zz_2889;
  wire       [15:0]   _zz_2890;
  wire       [0:0]    _zz_2891;
  wire       [0:0]    _zz_2892;
  wire       [15:0]   _zz_2893;
  wire       [15:0]   _zz_2894;
  wire       [15:0]   _zz_2895;
  wire       [0:0]    _zz_2896;
  wire       [0:0]    _zz_2897;
  wire       [15:0]   _zz_2898;
  wire       [15:0]   _zz_2899;
  wire       [15:0]   _zz_2900;
  wire       [0:0]    _zz_2901;
  wire       [0:0]    _zz_2902;
  wire       [15:0]   _zz_2903;
  wire       [15:0]   _zz_2904;
  wire       [15:0]   _zz_2905;
  wire       [0:0]    _zz_2906;
  wire       [0:0]    _zz_2907;
  wire       [15:0]   _zz_2908;
  wire       [15:0]   _zz_2909;
  wire       [15:0]   _zz_2910;
  wire       [0:0]    _zz_2911;
  wire       [0:0]    _zz_2912;
  wire       [15:0]   _zz_2913;
  wire       [15:0]   _zz_2914;
  wire       [15:0]   _zz_2915;
  wire       [0:0]    _zz_2916;
  wire       [0:0]    _zz_2917;
  wire       [15:0]   _zz_2918;
  wire       [15:0]   _zz_2919;
  wire       [15:0]   _zz_2920;
  wire       [0:0]    _zz_2921;
  wire       [0:0]    _zz_2922;
  wire       [15:0]   _zz_2923;
  wire       [15:0]   _zz_2924;
  wire       [15:0]   _zz_2925;
  wire       [0:0]    _zz_2926;
  wire       [0:0]    _zz_2927;
  wire       [15:0]   _zz_2928;
  wire       [15:0]   _zz_2929;
  wire       [15:0]   _zz_2930;
  wire       [0:0]    _zz_2931;
  wire       [0:0]    _zz_2932;
  wire       [15:0]   _zz_2933;
  wire       [15:0]   _zz_2934;
  wire       [15:0]   _zz_2935;
  wire       [0:0]    _zz_2936;
  wire       [0:0]    _zz_2937;
  wire       [15:0]   _zz_2938;
  wire       [15:0]   _zz_2939;
  wire       [15:0]   _zz_2940;
  wire       [0:0]    _zz_2941;
  wire       [0:0]    _zz_2942;
  wire       [15:0]   _zz_2943;
  wire       [15:0]   _zz_2944;
  wire       [15:0]   _zz_2945;
  wire       [0:0]    _zz_2946;
  wire       [0:0]    _zz_2947;
  wire       [15:0]   _zz_2948;
  wire       [15:0]   _zz_2949;
  wire       [15:0]   _zz_2950;
  wire       [0:0]    _zz_2951;
  wire       [0:0]    _zz_2952;
  wire       [15:0]   _zz_2953;
  wire       [15:0]   _zz_2954;
  wire       [15:0]   _zz_2955;
  wire       [0:0]    _zz_2956;
  wire       [0:0]    _zz_2957;
  wire       [15:0]   _zz_2958;
  wire       [15:0]   _zz_2959;
  wire       [15:0]   _zz_2960;
  wire       [0:0]    _zz_2961;
  wire       [0:0]    _zz_2962;
  wire       [15:0]   _zz_2963;
  wire       [15:0]   _zz_2964;
  wire       [15:0]   _zz_2965;
  wire       [0:0]    _zz_2966;
  wire       [0:0]    _zz_2967;
  wire       [15:0]   _zz_2968;
  wire       [15:0]   _zz_2969;
  wire       [15:0]   _zz_2970;
  wire       [0:0]    _zz_2971;
  wire       [0:0]    _zz_2972;
  wire       [15:0]   _zz_2973;
  wire       [15:0]   _zz_2974;
  wire       [15:0]   _zz_2975;
  wire       [0:0]    _zz_2976;
  wire       [0:0]    _zz_2977;
  wire       [15:0]   _zz_2978;
  wire       [15:0]   _zz_2979;
  wire       [15:0]   _zz_2980;
  wire       [0:0]    _zz_2981;
  wire       [0:0]    _zz_2982;
  wire       [15:0]   _zz_2983;
  wire       [15:0]   _zz_2984;
  wire       [15:0]   _zz_2985;
  wire       [0:0]    _zz_2986;
  wire       [0:0]    _zz_2987;
  wire       [15:0]   _zz_2988;
  wire       [15:0]   _zz_2989;
  wire       [15:0]   _zz_2990;
  wire       [0:0]    _zz_2991;
  wire       [0:0]    _zz_2992;
  wire       [15:0]   _zz_2993;
  wire       [15:0]   _zz_2994;
  wire       [15:0]   _zz_2995;
  wire       [0:0]    _zz_2996;
  wire       [0:0]    _zz_2997;
  wire       [15:0]   _zz_2998;
  wire       [15:0]   _zz_2999;
  wire       [15:0]   _zz_3000;
  wire       [0:0]    _zz_3001;
  wire       [0:0]    _zz_3002;
  wire       [15:0]   _zz_3003;
  wire       [15:0]   _zz_3004;
  wire       [15:0]   _zz_3005;
  wire       [0:0]    _zz_3006;
  wire       [0:0]    _zz_3007;
  wire       [15:0]   _zz_3008;
  wire       [15:0]   _zz_3009;
  wire       [15:0]   _zz_3010;
  wire       [0:0]    _zz_3011;
  wire       [0:0]    _zz_3012;
  wire       [15:0]   _zz_3013;
  wire       [15:0]   _zz_3014;
  wire       [15:0]   _zz_3015;
  wire       [0:0]    _zz_3016;
  wire       [0:0]    _zz_3017;
  wire       [15:0]   _zz_3018;
  wire       [15:0]   _zz_3019;
  wire       [15:0]   _zz_3020;
  wire       [0:0]    _zz_3021;
  wire       [0:0]    _zz_3022;
  wire       [15:0]   _zz_3023;
  wire       [15:0]   _zz_3024;
  wire       [15:0]   _zz_3025;
  wire       [0:0]    _zz_3026;
  wire       [0:0]    _zz_3027;
  wire       [15:0]   _zz_3028;
  wire       [15:0]   _zz_3029;
  wire       [15:0]   _zz_3030;
  wire       [0:0]    _zz_3031;
  wire       [0:0]    _zz_3032;
  wire       [15:0]   _zz_3033;
  wire       [15:0]   _zz_3034;
  wire       [15:0]   _zz_3035;
  wire       [0:0]    _zz_3036;
  wire       [0:0]    _zz_3037;
  wire       [15:0]   _zz_3038;
  wire       [15:0]   _zz_3039;
  wire       [15:0]   _zz_3040;
  wire       [0:0]    _zz_3041;
  wire       [0:0]    _zz_3042;
  wire       [15:0]   _zz_3043;
  wire       [15:0]   _zz_3044;
  wire       [15:0]   _zz_3045;
  wire       [0:0]    _zz_3046;
  wire       [0:0]    _zz_3047;
  wire       [15:0]   _zz_3048;
  wire       [15:0]   _zz_3049;
  wire       [15:0]   _zz_3050;
  wire       [0:0]    _zz_3051;
  wire       [0:0]    _zz_3052;
  wire       [15:0]   _zz_3053;
  wire       [15:0]   _zz_3054;
  wire       [15:0]   _zz_3055;
  wire       [0:0]    _zz_3056;
  wire       [0:0]    _zz_3057;
  wire       [15:0]   _zz_3058;
  wire       [15:0]   _zz_3059;
  wire       [15:0]   _zz_3060;
  wire       [0:0]    _zz_3061;
  wire       [0:0]    _zz_3062;
  wire       [15:0]   _zz_3063;
  wire       [15:0]   _zz_3064;
  wire       [15:0]   _zz_3065;
  wire       [0:0]    _zz_3066;
  wire       [0:0]    _zz_3067;
  wire       [15:0]   _zz_3068;
  wire       [15:0]   _zz_3069;
  wire       [15:0]   _zz_3070;
  wire       [0:0]    _zz_3071;
  wire       [0:0]    _zz_3072;
  wire       [15:0]   _zz_3073;
  wire       [15:0]   _zz_3074;
  wire       [15:0]   _zz_3075;
  wire       [0:0]    _zz_3076;
  wire       [0:0]    _zz_3077;
  wire       [15:0]   _zz_3078;
  wire       [15:0]   _zz_3079;
  wire       [15:0]   _zz_3080;
  wire       [0:0]    _zz_3081;
  wire       [0:0]    _zz_3082;
  wire       [15:0]   _zz_3083;
  wire       [15:0]   _zz_3084;
  wire       [15:0]   _zz_3085;
  wire       [0:0]    _zz_3086;
  wire       [0:0]    _zz_3087;
  wire       [15:0]   _zz_3088;
  wire       [15:0]   _zz_3089;
  wire       [15:0]   _zz_3090;
  wire       [0:0]    _zz_3091;
  wire       [0:0]    _zz_3092;
  wire       [15:0]   _zz_3093;
  wire       [15:0]   _zz_3094;
  wire       [15:0]   _zz_3095;
  wire       [0:0]    _zz_3096;
  wire       [0:0]    _zz_3097;
  wire       [15:0]   _zz_3098;
  wire       [15:0]   _zz_3099;
  wire       [15:0]   _zz_3100;
  wire       [0:0]    _zz_3101;
  wire       [0:0]    _zz_3102;
  wire       [15:0]   _zz_3103;
  wire       [15:0]   _zz_3104;
  wire       [15:0]   _zz_3105;
  wire       [0:0]    _zz_3106;
  wire       [0:0]    _zz_3107;
  wire       [15:0]   _zz_3108;
  wire       [15:0]   _zz_3109;
  wire       [15:0]   _zz_3110;
  wire       [0:0]    _zz_3111;
  wire       [0:0]    _zz_3112;
  wire       [15:0]   _zz_3113;
  wire       [15:0]   _zz_3114;
  wire       [15:0]   _zz_3115;
  wire       [0:0]    _zz_3116;
  wire       [0:0]    _zz_3117;
  wire       [15:0]   _zz_3118;
  wire       [15:0]   _zz_3119;
  wire       [15:0]   _zz_3120;
  wire       [0:0]    _zz_3121;
  wire       [0:0]    _zz_3122;
  wire       [15:0]   _zz_3123;
  wire       [15:0]   _zz_3124;
  wire       [15:0]   _zz_3125;
  wire       [0:0]    _zz_3126;
  wire       [0:0]    _zz_3127;
  wire       [15:0]   _zz_3128;
  wire       [15:0]   _zz_3129;
  wire       [15:0]   _zz_3130;
  wire       [0:0]    _zz_3131;
  wire       [0:0]    _zz_3132;
  wire       [15:0]   _zz_3133;
  wire       [15:0]   _zz_3134;
  wire       [15:0]   _zz_3135;
  wire       [0:0]    _zz_3136;
  wire       [0:0]    _zz_3137;
  wire       [15:0]   _zz_3138;
  wire       [15:0]   _zz_3139;
  wire       [15:0]   _zz_3140;
  wire       [0:0]    _zz_3141;
  wire       [0:0]    _zz_3142;
  wire       [15:0]   _zz_3143;
  wire       [15:0]   _zz_3144;
  wire       [15:0]   _zz_3145;
  wire       [0:0]    _zz_3146;
  wire       [0:0]    _zz_3147;
  wire       [15:0]   _zz_3148;
  wire       [15:0]   _zz_3149;
  wire       [15:0]   _zz_3150;
  wire       [0:0]    _zz_3151;
  wire       [0:0]    _zz_3152;
  wire       [15:0]   _zz_3153;
  wire       [15:0]   _zz_3154;
  wire       [15:0]   _zz_3155;
  wire       [0:0]    _zz_3156;
  wire       [0:0]    _zz_3157;
  wire       [15:0]   _zz_3158;
  wire       [15:0]   _zz_3159;
  wire       [15:0]   _zz_3160;
  wire       [0:0]    _zz_3161;
  wire       [0:0]    _zz_3162;
  wire       [15:0]   _zz_3163;
  wire       [15:0]   _zz_3164;
  wire       [15:0]   _zz_3165;
  wire       [0:0]    _zz_3166;
  wire       [0:0]    _zz_3167;
  wire       [15:0]   _zz_3168;
  wire       [15:0]   _zz_3169;
  wire       [15:0]   _zz_3170;
  wire       [0:0]    _zz_3171;
  wire       [0:0]    _zz_3172;
  wire       [15:0]   _zz_3173;
  wire       [15:0]   _zz_3174;
  wire       [15:0]   _zz_3175;
  wire       [0:0]    _zz_3176;
  wire       [0:0]    _zz_3177;
  wire       [15:0]   _zz_3178;
  wire       [15:0]   _zz_3179;
  wire       [15:0]   _zz_3180;
  wire       [0:0]    _zz_3181;
  wire       [0:0]    _zz_3182;
  wire       [15:0]   _zz_3183;
  wire       [15:0]   _zz_3184;
  wire       [15:0]   _zz_3185;
  wire       [0:0]    _zz_3186;
  wire       [0:0]    _zz_3187;
  wire       [15:0]   _zz_3188;
  wire       [15:0]   _zz_3189;
  wire       [15:0]   _zz_3190;
  wire       [0:0]    _zz_3191;
  wire       [0:0]    _zz_3192;
  wire       [15:0]   _zz_3193;
  wire       [15:0]   _zz_3194;
  wire       [15:0]   _zz_3195;
  wire       [0:0]    _zz_3196;
  wire       [0:0]    _zz_3197;
  wire       [15:0]   _zz_3198;
  wire       [15:0]   _zz_3199;
  wire       [15:0]   _zz_3200;
  wire       [0:0]    _zz_3201;
  wire       [0:0]    _zz_3202;
  wire       [15:0]   _zz_3203;
  wire       [15:0]   _zz_3204;
  wire       [15:0]   _zz_3205;
  wire       [0:0]    _zz_3206;
  wire       [0:0]    _zz_3207;
  wire       [15:0]   _zz_3208;
  wire       [15:0]   _zz_3209;
  wire       [15:0]   _zz_3210;
  wire       [0:0]    _zz_3211;
  wire       [0:0]    _zz_3212;
  wire       [15:0]   _zz_3213;
  wire       [15:0]   _zz_3214;
  wire       [15:0]   _zz_3215;
  wire       [0:0]    _zz_3216;
  wire       [0:0]    _zz_3217;
  wire       [15:0]   _zz_3218;
  wire       [15:0]   _zz_3219;
  wire       [15:0]   _zz_3220;
  wire       [0:0]    _zz_3221;
  wire       [0:0]    _zz_3222;
  wire       [15:0]   _zz_3223;
  wire       [15:0]   _zz_3224;
  wire       [15:0]   _zz_3225;
  wire       [0:0]    _zz_3226;
  wire       [0:0]    _zz_3227;
  wire       [15:0]   _zz_3228;
  wire       [15:0]   _zz_3229;
  wire       [15:0]   _zz_3230;
  wire       [0:0]    _zz_3231;
  wire       [0:0]    _zz_3232;
  wire       [15:0]   _zz_3233;
  wire       [15:0]   _zz_3234;
  wire       [15:0]   _zz_3235;
  wire       [0:0]    _zz_3236;
  wire       [0:0]    _zz_3237;
  wire       [15:0]   _zz_3238;
  wire       [15:0]   _zz_3239;
  wire       [15:0]   _zz_3240;
  wire       [0:0]    _zz_3241;
  wire       [0:0]    _zz_3242;
  wire       [15:0]   _zz_3243;
  wire       [15:0]   _zz_3244;
  wire       [15:0]   _zz_3245;
  wire       [0:0]    _zz_3246;
  wire       [0:0]    _zz_3247;
  wire       [15:0]   _zz_3248;
  wire       [15:0]   _zz_3249;
  wire       [15:0]   _zz_3250;
  wire       [0:0]    _zz_3251;
  wire       [0:0]    _zz_3252;
  wire       [15:0]   _zz_3253;
  wire       [15:0]   _zz_3254;
  wire       [15:0]   _zz_3255;
  wire       [0:0]    _zz_3256;
  wire       [0:0]    _zz_3257;
  wire       [15:0]   _zz_3258;
  wire       [15:0]   _zz_3259;
  wire       [15:0]   _zz_3260;
  wire       [0:0]    _zz_3261;
  wire       [0:0]    _zz_3262;
  wire       [15:0]   _zz_3263;
  wire       [15:0]   _zz_3264;
  wire       [15:0]   _zz_3265;
  wire       [0:0]    _zz_3266;
  wire       [0:0]    _zz_3267;
  wire       [15:0]   _zz_3268;
  wire       [15:0]   _zz_3269;
  wire       [15:0]   _zz_3270;
  wire       [0:0]    _zz_3271;
  wire       [0:0]    _zz_3272;
  wire       [15:0]   _zz_3273;
  wire       [15:0]   _zz_3274;
  wire       [15:0]   _zz_3275;
  wire       [0:0]    _zz_3276;
  wire       [0:0]    _zz_3277;
  wire       [15:0]   _zz_3278;
  wire       [15:0]   _zz_3279;
  wire       [15:0]   _zz_3280;
  wire       [0:0]    _zz_3281;
  wire       [0:0]    _zz_3282;
  wire       [15:0]   _zz_3283;
  wire       [15:0]   _zz_3284;
  wire       [15:0]   _zz_3285;
  wire       [0:0]    _zz_3286;
  wire       [0:0]    _zz_3287;
  wire       [15:0]   _zz_3288;
  wire       [15:0]   _zz_3289;
  wire       [15:0]   _zz_3290;
  wire       [0:0]    _zz_3291;
  wire       [0:0]    _zz_3292;
  wire       [15:0]   _zz_3293;
  wire       [15:0]   _zz_3294;
  wire       [15:0]   _zz_3295;
  wire       [0:0]    _zz_3296;
  wire       [0:0]    _zz_3297;
  wire       [15:0]   _zz_3298;
  wire       [15:0]   _zz_3299;
  wire       [15:0]   _zz_3300;
  wire       [0:0]    _zz_3301;
  wire       [0:0]    _zz_3302;
  wire       [15:0]   _zz_3303;
  wire       [15:0]   _zz_3304;
  wire       [15:0]   _zz_3305;
  wire       [0:0]    _zz_3306;
  wire       [0:0]    _zz_3307;
  wire       [15:0]   _zz_3308;
  wire       [15:0]   _zz_3309;
  wire       [15:0]   _zz_3310;
  wire       [0:0]    _zz_3311;
  wire       [0:0]    _zz_3312;
  wire       [15:0]   _zz_3313;
  wire       [15:0]   _zz_3314;
  wire       [15:0]   _zz_3315;
  wire       [0:0]    _zz_3316;
  wire       [0:0]    _zz_3317;
  wire       [15:0]   _zz_3318;
  wire       [15:0]   _zz_3319;
  wire       [15:0]   _zz_3320;
  wire       [0:0]    _zz_3321;
  wire       [0:0]    _zz_3322;
  wire       [15:0]   _zz_3323;
  wire       [15:0]   _zz_3324;
  wire       [15:0]   _zz_3325;
  wire       [0:0]    _zz_3326;
  wire       [0:0]    _zz_3327;
  wire       [15:0]   _zz_3328;
  wire       [15:0]   _zz_3329;
  wire       [15:0]   _zz_3330;
  wire       [0:0]    _zz_3331;
  wire       [0:0]    _zz_3332;
  wire       [15:0]   _zz_3333;
  wire       [15:0]   _zz_3334;
  wire       [15:0]   _zz_3335;
  wire       [0:0]    _zz_3336;
  wire       [0:0]    _zz_3337;
  wire       [15:0]   _zz_3338;
  wire       [15:0]   _zz_3339;
  wire       [15:0]   _zz_3340;
  wire       [0:0]    _zz_3341;
  wire       [0:0]    _zz_3342;
  wire       [15:0]   _zz_3343;
  wire       [15:0]   _zz_3344;
  wire       [15:0]   _zz_3345;
  wire       [0:0]    _zz_3346;
  wire       [0:0]    _zz_3347;
  wire       [15:0]   _zz_3348;
  wire       [15:0]   _zz_3349;
  wire       [15:0]   _zz_3350;
  wire       [0:0]    _zz_3351;
  wire       [0:0]    _zz_3352;
  wire       [15:0]   _zz_3353;
  wire       [15:0]   _zz_3354;
  wire       [15:0]   _zz_3355;
  wire       [0:0]    _zz_3356;
  wire       [0:0]    _zz_3357;
  wire       [15:0]   _zz_3358;
  wire       [15:0]   _zz_3359;
  wire       [15:0]   _zz_3360;
  wire       [0:0]    _zz_3361;
  wire       [0:0]    _zz_3362;
  wire       [15:0]   _zz_3363;
  wire       [15:0]   _zz_3364;
  wire       [15:0]   _zz_3365;
  wire       [0:0]    _zz_3366;
  wire       [0:0]    _zz_3367;
  wire       [15:0]   _zz_3368;
  wire       [15:0]   _zz_3369;
  wire       [15:0]   _zz_3370;
  wire       [0:0]    _zz_3371;
  wire       [0:0]    _zz_3372;
  wire       [15:0]   _zz_3373;
  wire       [15:0]   _zz_3374;
  wire       [15:0]   _zz_3375;
  wire       [0:0]    _zz_3376;
  wire       [0:0]    _zz_3377;
  wire       [15:0]   _zz_3378;
  wire       [15:0]   _zz_3379;
  wire       [15:0]   _zz_3380;
  wire       [0:0]    _zz_3381;
  wire       [0:0]    _zz_3382;
  wire       [15:0]   _zz_3383;
  wire       [15:0]   _zz_3384;
  wire       [15:0]   _zz_3385;
  wire       [0:0]    _zz_3386;
  wire       [0:0]    _zz_3387;
  wire       [15:0]   _zz_3388;
  wire       [15:0]   _zz_3389;
  wire       [15:0]   _zz_3390;
  wire       [0:0]    _zz_3391;
  wire       [0:0]    _zz_3392;
  wire       [15:0]   _zz_3393;
  wire       [15:0]   _zz_3394;
  wire       [15:0]   _zz_3395;
  wire       [0:0]    _zz_3396;
  wire       [0:0]    _zz_3397;
  wire       [15:0]   _zz_3398;
  wire       [15:0]   _zz_3399;
  wire       [15:0]   _zz_3400;
  wire       [0:0]    _zz_3401;
  wire       [0:0]    _zz_3402;
  wire       [15:0]   _zz_3403;
  wire       [15:0]   _zz_3404;
  wire       [15:0]   _zz_3405;
  wire       [0:0]    _zz_3406;
  wire       [0:0]    _zz_3407;
  wire       [15:0]   _zz_3408;
  wire       [15:0]   _zz_3409;
  wire       [15:0]   _zz_3410;
  wire       [0:0]    _zz_3411;
  wire       [0:0]    _zz_3412;
  wire       [15:0]   _zz_3413;
  wire       [15:0]   _zz_3414;
  wire       [15:0]   _zz_3415;
  wire       [0:0]    _zz_3416;
  wire       [0:0]    _zz_3417;
  wire       [15:0]   _zz_3418;
  wire       [15:0]   _zz_3419;
  wire       [15:0]   _zz_3420;
  wire       [0:0]    _zz_3421;
  wire       [0:0]    _zz_3422;
  wire       [15:0]   _zz_3423;
  wire       [15:0]   _zz_3424;
  wire       [15:0]   _zz_3425;
  wire       [0:0]    _zz_3426;
  wire       [0:0]    _zz_3427;
  wire       [15:0]   _zz_3428;
  wire       [15:0]   _zz_3429;
  wire       [15:0]   _zz_3430;
  wire       [0:0]    _zz_3431;
  wire       [0:0]    _zz_3432;
  wire       [15:0]   _zz_3433;
  wire       [15:0]   _zz_3434;
  wire       [15:0]   _zz_3435;
  wire       [0:0]    _zz_3436;
  wire       [0:0]    _zz_3437;
  wire       [15:0]   _zz_3438;
  wire       [15:0]   _zz_3439;
  wire       [15:0]   _zz_3440;
  wire       [0:0]    _zz_3441;
  wire       [0:0]    _zz_3442;
  wire       [15:0]   _zz_3443;
  wire       [15:0]   _zz_3444;
  wire       [15:0]   _zz_3445;
  wire       [0:0]    _zz_3446;
  wire       [0:0]    _zz_3447;
  wire       [15:0]   _zz_3448;
  wire       [15:0]   _zz_3449;
  wire       [15:0]   _zz_3450;
  wire       [0:0]    _zz_3451;
  wire       [0:0]    _zz_3452;
  wire       [15:0]   _zz_3453;
  wire       [15:0]   _zz_3454;
  wire       [15:0]   _zz_3455;
  wire       [0:0]    _zz_3456;
  wire       [0:0]    _zz_3457;
  wire       [15:0]   _zz_3458;
  wire       [15:0]   _zz_3459;
  wire       [15:0]   _zz_3460;
  wire       [0:0]    _zz_3461;
  wire       [0:0]    _zz_3462;
  wire       [15:0]   _zz_3463;
  wire       [15:0]   _zz_3464;
  wire       [15:0]   _zz_3465;
  wire       [0:0]    _zz_3466;
  wire       [0:0]    _zz_3467;
  wire       [15:0]   _zz_3468;
  wire       [15:0]   _zz_3469;
  wire       [15:0]   _zz_3470;
  wire       [0:0]    _zz_3471;
  wire       [0:0]    _zz_3472;
  wire       [15:0]   _zz_3473;
  wire       [15:0]   _zz_3474;
  wire       [15:0]   _zz_3475;
  wire       [0:0]    _zz_3476;
  wire       [0:0]    _zz_3477;
  wire       [15:0]   _zz_3478;
  wire       [15:0]   _zz_3479;
  wire       [15:0]   _zz_3480;
  wire       [0:0]    _zz_3481;
  wire       [0:0]    _zz_3482;
  wire       [15:0]   _zz_3483;
  wire       [15:0]   _zz_3484;
  wire       [15:0]   _zz_3485;
  wire       [0:0]    _zz_3486;
  wire       [0:0]    _zz_3487;
  wire       [15:0]   _zz_3488;
  wire       [15:0]   _zz_3489;
  wire       [15:0]   _zz_3490;
  wire       [0:0]    _zz_3491;
  wire       [0:0]    _zz_3492;
  wire       [15:0]   _zz_3493;
  wire       [15:0]   _zz_3494;
  wire       [15:0]   _zz_3495;
  wire       [0:0]    _zz_3496;
  wire       [0:0]    _zz_3497;
  wire       [15:0]   _zz_3498;
  wire       [15:0]   _zz_3499;
  wire       [15:0]   _zz_3500;
  wire       [0:0]    _zz_3501;
  wire       [0:0]    _zz_3502;
  wire       [15:0]   _zz_3503;
  wire       [15:0]   _zz_3504;
  wire       [15:0]   _zz_3505;
  wire       [0:0]    _zz_3506;
  wire       [0:0]    _zz_3507;
  wire       [15:0]   _zz_3508;
  wire       [15:0]   _zz_3509;
  wire       [15:0]   _zz_3510;
  wire       [0:0]    _zz_3511;
  wire       [0:0]    _zz_3512;
  wire       [15:0]   _zz_3513;
  wire       [15:0]   _zz_3514;
  wire       [15:0]   _zz_3515;
  wire       [0:0]    _zz_3516;
  wire       [0:0]    _zz_3517;
  wire       [15:0]   _zz_3518;
  wire       [15:0]   _zz_3519;
  wire       [15:0]   _zz_3520;
  wire       [0:0]    _zz_3521;
  wire       [0:0]    _zz_3522;
  wire       [15:0]   _zz_3523;
  wire       [15:0]   _zz_3524;
  wire       [15:0]   _zz_3525;
  wire       [0:0]    _zz_3526;
  wire       [0:0]    _zz_3527;
  wire       [15:0]   _zz_3528;
  wire       [15:0]   _zz_3529;
  wire       [15:0]   _zz_3530;
  wire       [0:0]    _zz_3531;
  wire       [0:0]    _zz_3532;
  wire       [15:0]   _zz_3533;
  wire       [15:0]   _zz_3534;
  wire       [15:0]   _zz_3535;
  wire       [0:0]    _zz_3536;
  wire       [0:0]    _zz_3537;
  wire       [15:0]   _zz_3538;
  wire       [15:0]   _zz_3539;
  wire       [15:0]   _zz_3540;
  wire       [0:0]    _zz_3541;
  wire       [0:0]    _zz_3542;
  wire       [15:0]   _zz_3543;
  wire       [15:0]   _zz_3544;
  wire       [15:0]   _zz_3545;
  wire       [0:0]    _zz_3546;
  wire       [0:0]    _zz_3547;
  wire       [15:0]   _zz_3548;
  wire       [15:0]   _zz_3549;
  wire       [15:0]   _zz_3550;
  wire       [0:0]    _zz_3551;
  wire       [0:0]    _zz_3552;
  wire       [15:0]   _zz_3553;
  wire       [15:0]   _zz_3554;
  wire       [15:0]   _zz_3555;
  wire       [0:0]    _zz_3556;
  wire       [0:0]    _zz_3557;
  wire       [15:0]   _zz_3558;
  wire       [15:0]   _zz_3559;
  wire       [15:0]   _zz_3560;
  wire       [0:0]    _zz_3561;
  wire       [0:0]    _zz_3562;
  wire       [15:0]   _zz_3563;
  wire       [15:0]   _zz_3564;
  wire       [15:0]   _zz_3565;
  wire       [0:0]    _zz_3566;
  wire       [0:0]    _zz_3567;
  wire       [15:0]   _zz_3568;
  wire       [15:0]   _zz_3569;
  wire       [15:0]   _zz_3570;
  wire       [0:0]    _zz_3571;
  wire       [0:0]    _zz_3572;
  wire       [15:0]   _zz_3573;
  wire       [15:0]   _zz_3574;
  wire       [15:0]   _zz_3575;
  wire       [0:0]    _zz_3576;
  wire       [0:0]    _zz_3577;
  wire       [15:0]   _zz_3578;
  wire       [15:0]   _zz_3579;
  wire       [15:0]   _zz_3580;
  wire       [0:0]    _zz_3581;
  wire       [0:0]    _zz_3582;
  wire       [15:0]   _zz_3583;
  wire       [15:0]   _zz_3584;
  wire       [15:0]   _zz_3585;
  wire       [0:0]    _zz_3586;
  wire       [0:0]    _zz_3587;
  wire       [15:0]   _zz_3588;
  wire       [15:0]   _zz_3589;
  wire       [15:0]   _zz_3590;
  wire       [0:0]    _zz_3591;
  wire       [0:0]    _zz_3592;
  wire       [15:0]   _zz_3593;
  wire       [15:0]   _zz_3594;
  wire       [15:0]   _zz_3595;
  wire       [0:0]    _zz_3596;
  wire       [0:0]    _zz_3597;
  wire       [15:0]   _zz_3598;
  wire       [15:0]   _zz_3599;
  wire       [15:0]   _zz_3600;
  wire       [0:0]    _zz_3601;
  wire       [0:0]    _zz_3602;
  wire       [15:0]   _zz_3603;
  wire       [15:0]   _zz_3604;
  wire       [15:0]   _zz_3605;
  wire       [0:0]    _zz_3606;
  wire       [0:0]    _zz_3607;
  wire       [15:0]   _zz_3608;
  wire       [15:0]   _zz_3609;
  wire       [15:0]   _zz_3610;
  wire       [0:0]    _zz_3611;
  wire       [0:0]    _zz_3612;
  wire       [15:0]   _zz_3613;
  wire       [15:0]   _zz_3614;
  wire       [15:0]   _zz_3615;
  wire       [0:0]    _zz_3616;
  wire       [0:0]    _zz_3617;
  wire       [15:0]   _zz_3618;
  wire       [15:0]   _zz_3619;
  wire       [15:0]   _zz_3620;
  wire       [0:0]    _zz_3621;
  wire       [0:0]    _zz_3622;
  wire       [15:0]   _zz_3623;
  wire       [15:0]   _zz_3624;
  wire       [15:0]   _zz_3625;
  wire       [0:0]    _zz_3626;
  wire       [0:0]    _zz_3627;
  wire       [15:0]   _zz_3628;
  wire       [15:0]   _zz_3629;
  wire       [15:0]   _zz_3630;
  wire       [0:0]    _zz_3631;
  wire       [0:0]    _zz_3632;
  wire       [15:0]   _zz_3633;
  wire       [15:0]   _zz_3634;
  wire       [15:0]   _zz_3635;
  wire       [0:0]    _zz_3636;
  wire       [0:0]    _zz_3637;
  wire       [15:0]   _zz_3638;
  wire       [15:0]   _zz_3639;
  wire       [15:0]   _zz_3640;
  wire       [0:0]    _zz_3641;
  wire       [0:0]    _zz_3642;
  wire       [15:0]   _zz_3643;
  wire       [15:0]   _zz_3644;
  wire       [15:0]   _zz_3645;
  wire       [0:0]    _zz_3646;
  wire       [0:0]    _zz_3647;
  wire       [15:0]   _zz_3648;
  wire       [15:0]   _zz_3649;
  wire       [15:0]   _zz_3650;
  wire       [0:0]    _zz_3651;
  wire       [0:0]    _zz_3652;
  wire       [15:0]   _zz_3653;
  wire       [15:0]   _zz_3654;
  wire       [15:0]   _zz_3655;
  wire       [0:0]    _zz_3656;
  wire       [0:0]    _zz_3657;
  wire       [15:0]   _zz_3658;
  wire       [15:0]   _zz_3659;
  wire       [15:0]   _zz_3660;
  wire       [0:0]    _zz_3661;
  wire       [0:0]    _zz_3662;
  wire       [15:0]   _zz_3663;
  wire       [15:0]   _zz_3664;
  wire       [15:0]   _zz_3665;
  wire       [0:0]    _zz_3666;
  wire       [0:0]    _zz_3667;
  wire       [15:0]   _zz_3668;
  wire       [15:0]   _zz_3669;
  wire       [15:0]   _zz_3670;
  wire       [0:0]    _zz_3671;
  wire       [0:0]    _zz_3672;
  wire       [15:0]   _zz_3673;
  wire       [15:0]   _zz_3674;
  wire       [15:0]   _zz_3675;
  wire       [0:0]    _zz_3676;
  wire       [0:0]    _zz_3677;
  wire       [15:0]   _zz_3678;
  wire       [15:0]   _zz_3679;
  wire       [15:0]   _zz_3680;
  wire       [0:0]    _zz_3681;
  wire       [0:0]    _zz_3682;
  wire       [15:0]   _zz_3683;
  wire       [15:0]   _zz_3684;
  wire       [15:0]   _zz_3685;
  wire       [0:0]    _zz_3686;
  wire       [0:0]    _zz_3687;
  wire       [15:0]   _zz_3688;
  wire       [15:0]   _zz_3689;
  wire       [15:0]   _zz_3690;
  wire       [0:0]    _zz_3691;
  wire       [0:0]    _zz_3692;
  wire       [15:0]   _zz_3693;
  wire       [15:0]   _zz_3694;
  wire       [15:0]   _zz_3695;
  wire       [0:0]    _zz_3696;
  wire       [0:0]    _zz_3697;
  wire       [15:0]   _zz_3698;
  wire       [15:0]   _zz_3699;
  wire       [15:0]   _zz_3700;
  wire       [0:0]    _zz_3701;
  wire       [0:0]    _zz_3702;
  wire       [15:0]   _zz_3703;
  wire       [15:0]   _zz_3704;
  wire       [15:0]   _zz_3705;
  wire       [0:0]    _zz_3706;
  wire       [0:0]    _zz_3707;
  wire       [15:0]   _zz_3708;
  wire       [15:0]   _zz_3709;
  wire       [15:0]   _zz_3710;
  wire       [0:0]    _zz_3711;
  wire       [0:0]    _zz_3712;
  wire       [15:0]   _zz_3713;
  wire       [15:0]   _zz_3714;
  wire       [15:0]   _zz_3715;
  wire       [0:0]    _zz_3716;
  wire       [0:0]    _zz_3717;
  wire       [15:0]   _zz_3718;
  wire       [15:0]   _zz_3719;
  wire       [15:0]   _zz_3720;
  wire       [0:0]    _zz_3721;
  wire       [0:0]    _zz_3722;
  wire       [15:0]   _zz_3723;
  wire       [15:0]   _zz_3724;
  wire       [15:0]   _zz_3725;
  wire       [0:0]    _zz_3726;
  wire       [0:0]    _zz_3727;
  wire       [15:0]   _zz_3728;
  wire       [15:0]   _zz_3729;
  wire       [15:0]   _zz_3730;
  wire       [0:0]    _zz_3731;
  wire       [0:0]    _zz_3732;
  wire       [15:0]   _zz_3733;
  wire       [15:0]   _zz_3734;
  wire       [15:0]   _zz_3735;
  wire       [0:0]    _zz_3736;
  wire       [0:0]    _zz_3737;
  wire       [15:0]   _zz_3738;
  wire       [15:0]   _zz_3739;
  wire       [15:0]   _zz_3740;
  wire       [0:0]    _zz_3741;
  wire       [0:0]    _zz_3742;
  wire       [15:0]   _zz_3743;
  wire       [15:0]   _zz_3744;
  wire       [15:0]   _zz_3745;
  wire       [0:0]    _zz_3746;
  wire       [0:0]    _zz_3747;
  wire       [15:0]   _zz_3748;
  wire       [15:0]   _zz_3749;
  wire       [15:0]   _zz_3750;
  wire       [0:0]    _zz_3751;
  wire       [0:0]    _zz_3752;
  wire       [15:0]   _zz_3753;
  wire       [15:0]   _zz_3754;
  wire       [15:0]   _zz_3755;
  wire       [0:0]    _zz_3756;
  wire       [0:0]    _zz_3757;
  wire       [15:0]   _zz_3758;
  wire       [15:0]   _zz_3759;
  wire       [15:0]   _zz_3760;
  wire       [0:0]    _zz_3761;
  wire       [0:0]    _zz_3762;
  wire       [15:0]   _zz_3763;
  wire       [15:0]   _zz_3764;
  wire       [15:0]   _zz_3765;
  wire       [0:0]    _zz_3766;
  wire       [0:0]    _zz_3767;
  wire       [15:0]   _zz_3768;
  wire       [15:0]   _zz_3769;
  wire       [15:0]   _zz_3770;
  wire       [0:0]    _zz_3771;
  wire       [0:0]    _zz_3772;
  wire       [15:0]   _zz_3773;
  wire       [15:0]   _zz_3774;
  wire       [15:0]   _zz_3775;
  wire       [0:0]    _zz_3776;
  wire       [0:0]    _zz_3777;
  wire       [15:0]   _zz_3778;
  wire       [15:0]   _zz_3779;
  wire       [15:0]   _zz_3780;
  wire       [0:0]    _zz_3781;
  wire       [0:0]    _zz_3782;
  wire       [15:0]   _zz_3783;
  wire       [15:0]   _zz_3784;
  wire       [15:0]   _zz_3785;
  wire       [0:0]    _zz_3786;
  wire       [0:0]    _zz_3787;
  wire       [15:0]   _zz_3788;
  wire       [15:0]   _zz_3789;
  wire       [15:0]   _zz_3790;
  wire       [0:0]    _zz_3791;
  wire       [0:0]    _zz_3792;
  wire       [15:0]   _zz_3793;
  wire       [15:0]   _zz_3794;
  wire       [15:0]   _zz_3795;
  wire       [0:0]    _zz_3796;
  wire       [0:0]    _zz_3797;
  wire       [15:0]   _zz_3798;
  wire       [15:0]   _zz_3799;
  wire       [15:0]   _zz_3800;
  wire       [0:0]    _zz_3801;
  wire       [0:0]    _zz_3802;
  wire       [15:0]   _zz_3803;
  wire       [15:0]   _zz_3804;
  wire       [15:0]   _zz_3805;
  wire       [0:0]    _zz_3806;
  wire       [0:0]    _zz_3807;
  wire       [15:0]   _zz_3808;
  wire       [15:0]   _zz_3809;
  wire       [15:0]   _zz_3810;
  wire       [0:0]    _zz_3811;
  wire       [0:0]    _zz_3812;
  wire       [15:0]   _zz_3813;
  wire       [15:0]   _zz_3814;
  wire       [15:0]   _zz_3815;
  wire       [0:0]    _zz_3816;
  wire       [0:0]    _zz_3817;
  wire       [15:0]   _zz_3818;
  wire       [15:0]   _zz_3819;
  wire       [15:0]   _zz_3820;
  wire       [0:0]    _zz_3821;
  wire       [0:0]    _zz_3822;
  wire       [15:0]   _zz_3823;
  wire       [15:0]   _zz_3824;
  wire       [15:0]   _zz_3825;
  wire       [0:0]    _zz_3826;
  wire       [0:0]    _zz_3827;
  wire       [15:0]   _zz_3828;
  wire       [15:0]   _zz_3829;
  wire       [15:0]   _zz_3830;
  wire       [0:0]    _zz_3831;
  wire       [0:0]    _zz_3832;
  wire       [15:0]   _zz_3833;
  wire       [15:0]   _zz_3834;
  wire       [15:0]   _zz_3835;
  wire       [0:0]    _zz_3836;
  wire       [0:0]    _zz_3837;
  wire       [15:0]   _zz_3838;
  wire       [15:0]   _zz_3839;
  wire       [15:0]   _zz_3840;
  wire       [0:0]    _zz_3841;
  wire       [0:0]    _zz_3842;
  wire       [15:0]   _zz_3843;
  wire       [15:0]   _zz_3844;
  wire       [15:0]   _zz_3845;
  wire       [0:0]    _zz_3846;
  wire       [0:0]    _zz_3847;
  wire       [15:0]   _zz_3848;
  wire       [15:0]   _zz_3849;
  wire       [15:0]   _zz_3850;
  wire       [0:0]    _zz_3851;
  wire       [0:0]    _zz_3852;
  wire       [15:0]   _zz_3853;
  wire       [15:0]   _zz_3854;
  wire       [15:0]   _zz_3855;
  wire       [0:0]    _zz_3856;
  wire       [0:0]    _zz_3857;
  wire       [15:0]   _zz_3858;
  wire       [15:0]   _zz_3859;
  wire       [15:0]   _zz_3860;
  wire       [0:0]    _zz_3861;
  wire       [0:0]    _zz_3862;
  wire       [15:0]   _zz_3863;
  wire       [15:0]   _zz_3864;
  wire       [15:0]   _zz_3865;
  wire       [0:0]    _zz_3866;
  wire       [0:0]    _zz_3867;
  wire       [15:0]   _zz_3868;
  wire       [15:0]   _zz_3869;
  wire       [15:0]   _zz_3870;
  wire       [0:0]    _zz_3871;
  wire       [0:0]    _zz_3872;
  wire       [15:0]   _zz_3873;
  wire       [15:0]   _zz_3874;
  wire       [15:0]   _zz_3875;
  wire       [0:0]    _zz_3876;
  wire       [0:0]    _zz_3877;
  wire       [15:0]   _zz_3878;
  wire       [15:0]   _zz_3879;
  wire       [15:0]   _zz_3880;
  wire       [0:0]    _zz_3881;
  wire       [0:0]    _zz_3882;
  wire       [15:0]   _zz_3883;
  wire       [15:0]   _zz_3884;
  wire       [15:0]   _zz_3885;
  wire       [0:0]    _zz_3886;
  wire       [0:0]    _zz_3887;
  wire       [15:0]   _zz_3888;
  wire       [15:0]   _zz_3889;
  wire       [15:0]   _zz_3890;
  wire       [0:0]    _zz_3891;
  wire       [0:0]    _zz_3892;
  wire       [15:0]   _zz_3893;
  wire       [15:0]   _zz_3894;
  wire       [15:0]   _zz_3895;
  wire       [0:0]    _zz_3896;
  wire       [0:0]    _zz_3897;
  wire       [15:0]   _zz_3898;
  wire       [15:0]   _zz_3899;
  wire       [15:0]   _zz_3900;
  wire       [0:0]    _zz_3901;
  wire       [0:0]    _zz_3902;
  wire       [15:0]   _zz_3903;
  wire       [15:0]   _zz_3904;
  wire       [15:0]   _zz_3905;
  wire       [0:0]    _zz_3906;
  wire       [0:0]    _zz_3907;
  wire       [15:0]   _zz_3908;
  wire       [15:0]   _zz_3909;
  wire       [15:0]   _zz_3910;
  wire       [0:0]    _zz_3911;
  wire       [0:0]    _zz_3912;
  wire       [15:0]   _zz_3913;
  wire       [15:0]   _zz_3914;
  wire       [15:0]   _zz_3915;
  wire       [0:0]    _zz_3916;
  wire       [0:0]    _zz_3917;
  wire       [15:0]   _zz_3918;
  wire       [15:0]   _zz_3919;
  wire       [15:0]   _zz_3920;
  wire       [0:0]    _zz_3921;
  wire       [0:0]    _zz_3922;
  wire       [15:0]   _zz_3923;
  wire       [15:0]   _zz_3924;
  wire       [15:0]   _zz_3925;
  wire       [0:0]    _zz_3926;
  wire       [0:0]    _zz_3927;
  wire       [15:0]   _zz_3928;
  wire       [15:0]   _zz_3929;
  wire       [15:0]   _zz_3930;
  wire       [0:0]    _zz_3931;
  wire       [0:0]    _zz_3932;
  wire       [15:0]   _zz_3933;
  wire       [15:0]   _zz_3934;
  wire       [15:0]   _zz_3935;
  wire       [0:0]    _zz_3936;
  wire       [0:0]    _zz_3937;
  wire       [15:0]   _zz_3938;
  wire       [15:0]   _zz_3939;
  wire       [15:0]   _zz_3940;
  wire       [0:0]    _zz_3941;
  wire       [0:0]    _zz_3942;
  wire       [15:0]   _zz_3943;
  wire       [15:0]   _zz_3944;
  wire       [15:0]   _zz_3945;
  wire       [0:0]    _zz_3946;
  wire       [0:0]    _zz_3947;
  wire       [15:0]   _zz_3948;
  wire       [15:0]   _zz_3949;
  wire       [15:0]   _zz_3950;
  wire       [0:0]    _zz_3951;
  wire       [0:0]    _zz_3952;
  wire       [15:0]   _zz_3953;
  wire       [15:0]   _zz_3954;
  wire       [15:0]   _zz_3955;
  wire       [0:0]    _zz_3956;
  wire       [0:0]    _zz_3957;
  wire       [15:0]   _zz_3958;
  wire       [15:0]   _zz_3959;
  wire       [15:0]   _zz_3960;
  wire       [0:0]    _zz_3961;
  wire       [0:0]    _zz_3962;
  wire       [15:0]   _zz_3963;
  wire       [15:0]   _zz_3964;
  wire       [15:0]   _zz_3965;
  wire       [0:0]    _zz_3966;
  wire       [0:0]    _zz_3967;
  wire       [15:0]   _zz_3968;
  wire       [15:0]   _zz_3969;
  wire       [15:0]   _zz_3970;
  wire       [0:0]    _zz_3971;
  wire       [0:0]    _zz_3972;
  wire       [15:0]   _zz_3973;
  wire       [15:0]   _zz_3974;
  wire       [15:0]   _zz_3975;
  wire       [0:0]    _zz_3976;
  wire       [0:0]    _zz_3977;
  wire       [15:0]   _zz_3978;
  wire       [15:0]   _zz_3979;
  wire       [15:0]   _zz_3980;
  wire       [0:0]    _zz_3981;
  wire       [0:0]    _zz_3982;
  wire       [15:0]   _zz_3983;
  wire       [15:0]   _zz_3984;
  wire       [15:0]   _zz_3985;
  wire       [0:0]    _zz_3986;
  wire       [0:0]    _zz_3987;
  wire       [15:0]   _zz_3988;
  wire       [15:0]   _zz_3989;
  wire       [15:0]   _zz_3990;
  wire       [0:0]    _zz_3991;
  wire       [0:0]    _zz_3992;
  wire       [15:0]   _zz_3993;
  wire       [15:0]   _zz_3994;
  wire       [15:0]   _zz_3995;
  wire       [0:0]    _zz_3996;
  wire       [0:0]    _zz_3997;
  wire       [15:0]   _zz_3998;
  wire       [15:0]   _zz_3999;
  wire       [15:0]   _zz_4000;
  wire       [0:0]    _zz_4001;
  wire       [0:0]    _zz_4002;
  wire       [15:0]   _zz_4003;
  wire       [15:0]   _zz_4004;
  wire       [15:0]   _zz_4005;
  wire       [0:0]    _zz_4006;
  wire       [0:0]    _zz_4007;
  wire       [15:0]   _zz_4008;
  wire       [15:0]   _zz_4009;
  wire       [15:0]   _zz_4010;
  wire       [0:0]    _zz_4011;
  wire       [0:0]    _zz_4012;
  wire       [15:0]   _zz_4013;
  wire       [15:0]   _zz_4014;
  wire       [15:0]   _zz_4015;
  wire       [0:0]    _zz_4016;
  wire       [0:0]    _zz_4017;
  wire       [15:0]   _zz_4018;
  wire       [15:0]   _zz_4019;
  wire       [15:0]   _zz_4020;
  wire       [0:0]    _zz_4021;
  wire       [0:0]    _zz_4022;
  wire       [15:0]   _zz_4023;
  wire       [15:0]   _zz_4024;
  wire       [15:0]   _zz_4025;
  wire       [0:0]    _zz_4026;
  wire       [0:0]    _zz_4027;
  wire       [15:0]   _zz_4028;
  wire       [15:0]   _zz_4029;
  wire       [15:0]   _zz_4030;
  wire       [0:0]    _zz_4031;
  wire       [0:0]    _zz_4032;
  reg                 io_data_in_valid_regNext;
  reg                 _zz_4033;
  reg        [3:0]    _zz_4034;
  reg        [3:0]    _zz_4035;
  wire                _zz_4036;
  wire                _zz_4037;
  reg                 _zz_4038;

  assign _zz_5383 = ($signed(twiddle_factor_table_0_real) + $signed(twiddle_factor_table_0_imag));
  assign _zz_5384 = fixTo_dout;
  assign _zz_5385 = ($signed(_zz_4) - $signed(_zz_3));
  assign _zz_5386 = ($signed(_zz_3) + $signed(_zz_4));
  assign _zz_5387 = _zz_5388[15 : 0];
  assign _zz_5388 = fixTo_2_dout;
  assign _zz_5389 = _zz_5390[15 : 0];
  assign _zz_5390 = fixTo_1_dout;
  assign _zz_5391 = _zz_5392;
  assign _zz_5392 = ($signed(_zz_5393) >>> _zz_1796);
  assign _zz_5393 = _zz_5394;
  assign _zz_5394 = ($signed(_zz_1) - $signed(_zz_1793));
  assign _zz_5395 = _zz_5396;
  assign _zz_5396 = ($signed(_zz_5397) >>> _zz_1796);
  assign _zz_5397 = _zz_5398;
  assign _zz_5398 = ($signed(_zz_2) - $signed(_zz_1794));
  assign _zz_5399 = _zz_5400;
  assign _zz_5400 = ($signed(_zz_5401) >>> _zz_1797);
  assign _zz_5401 = _zz_5402;
  assign _zz_5402 = ($signed(_zz_1) + $signed(_zz_1793));
  assign _zz_5403 = _zz_5404;
  assign _zz_5404 = ($signed(_zz_5405) >>> _zz_1797);
  assign _zz_5405 = _zz_5406;
  assign _zz_5406 = ($signed(_zz_2) + $signed(_zz_1794));
  assign _zz_5407 = ($signed(twiddle_factor_table_0_real) + $signed(twiddle_factor_table_0_imag));
  assign _zz_5408 = fixTo_3_dout;
  assign _zz_5409 = ($signed(_zz_8) - $signed(_zz_7));
  assign _zz_5410 = ($signed(_zz_7) + $signed(_zz_8));
  assign _zz_5411 = _zz_5412[15 : 0];
  assign _zz_5412 = fixTo_5_dout;
  assign _zz_5413 = _zz_5414[15 : 0];
  assign _zz_5414 = fixTo_4_dout;
  assign _zz_5415 = _zz_5416;
  assign _zz_5416 = ($signed(_zz_5417) >>> _zz_1801);
  assign _zz_5417 = _zz_5418;
  assign _zz_5418 = ($signed(_zz_5) - $signed(_zz_1798));
  assign _zz_5419 = _zz_5420;
  assign _zz_5420 = ($signed(_zz_5421) >>> _zz_1801);
  assign _zz_5421 = _zz_5422;
  assign _zz_5422 = ($signed(_zz_6) - $signed(_zz_1799));
  assign _zz_5423 = _zz_5424;
  assign _zz_5424 = ($signed(_zz_5425) >>> _zz_1802);
  assign _zz_5425 = _zz_5426;
  assign _zz_5426 = ($signed(_zz_5) + $signed(_zz_1798));
  assign _zz_5427 = _zz_5428;
  assign _zz_5428 = ($signed(_zz_5429) >>> _zz_1802);
  assign _zz_5429 = _zz_5430;
  assign _zz_5430 = ($signed(_zz_6) + $signed(_zz_1799));
  assign _zz_5431 = ($signed(twiddle_factor_table_0_real) + $signed(twiddle_factor_table_0_imag));
  assign _zz_5432 = fixTo_6_dout;
  assign _zz_5433 = ($signed(_zz_12) - $signed(_zz_11));
  assign _zz_5434 = ($signed(_zz_11) + $signed(_zz_12));
  assign _zz_5435 = _zz_5436[15 : 0];
  assign _zz_5436 = fixTo_8_dout;
  assign _zz_5437 = _zz_5438[15 : 0];
  assign _zz_5438 = fixTo_7_dout;
  assign _zz_5439 = _zz_5440;
  assign _zz_5440 = ($signed(_zz_5441) >>> _zz_1806);
  assign _zz_5441 = _zz_5442;
  assign _zz_5442 = ($signed(_zz_9) - $signed(_zz_1803));
  assign _zz_5443 = _zz_5444;
  assign _zz_5444 = ($signed(_zz_5445) >>> _zz_1806);
  assign _zz_5445 = _zz_5446;
  assign _zz_5446 = ($signed(_zz_10) - $signed(_zz_1804));
  assign _zz_5447 = _zz_5448;
  assign _zz_5448 = ($signed(_zz_5449) >>> _zz_1807);
  assign _zz_5449 = _zz_5450;
  assign _zz_5450 = ($signed(_zz_9) + $signed(_zz_1803));
  assign _zz_5451 = _zz_5452;
  assign _zz_5452 = ($signed(_zz_5453) >>> _zz_1807);
  assign _zz_5453 = _zz_5454;
  assign _zz_5454 = ($signed(_zz_10) + $signed(_zz_1804));
  assign _zz_5455 = ($signed(twiddle_factor_table_0_real) + $signed(twiddle_factor_table_0_imag));
  assign _zz_5456 = fixTo_9_dout;
  assign _zz_5457 = ($signed(_zz_16) - $signed(_zz_15));
  assign _zz_5458 = ($signed(_zz_15) + $signed(_zz_16));
  assign _zz_5459 = _zz_5460[15 : 0];
  assign _zz_5460 = fixTo_11_dout;
  assign _zz_5461 = _zz_5462[15 : 0];
  assign _zz_5462 = fixTo_10_dout;
  assign _zz_5463 = _zz_5464;
  assign _zz_5464 = ($signed(_zz_5465) >>> _zz_1811);
  assign _zz_5465 = _zz_5466;
  assign _zz_5466 = ($signed(_zz_13) - $signed(_zz_1808));
  assign _zz_5467 = _zz_5468;
  assign _zz_5468 = ($signed(_zz_5469) >>> _zz_1811);
  assign _zz_5469 = _zz_5470;
  assign _zz_5470 = ($signed(_zz_14) - $signed(_zz_1809));
  assign _zz_5471 = _zz_5472;
  assign _zz_5472 = ($signed(_zz_5473) >>> _zz_1812);
  assign _zz_5473 = _zz_5474;
  assign _zz_5474 = ($signed(_zz_13) + $signed(_zz_1808));
  assign _zz_5475 = _zz_5476;
  assign _zz_5476 = ($signed(_zz_5477) >>> _zz_1812);
  assign _zz_5477 = _zz_5478;
  assign _zz_5478 = ($signed(_zz_14) + $signed(_zz_1809));
  assign _zz_5479 = ($signed(twiddle_factor_table_0_real) + $signed(twiddle_factor_table_0_imag));
  assign _zz_5480 = fixTo_12_dout;
  assign _zz_5481 = ($signed(_zz_20) - $signed(_zz_19));
  assign _zz_5482 = ($signed(_zz_19) + $signed(_zz_20));
  assign _zz_5483 = _zz_5484[15 : 0];
  assign _zz_5484 = fixTo_14_dout;
  assign _zz_5485 = _zz_5486[15 : 0];
  assign _zz_5486 = fixTo_13_dout;
  assign _zz_5487 = _zz_5488;
  assign _zz_5488 = ($signed(_zz_5489) >>> _zz_1816);
  assign _zz_5489 = _zz_5490;
  assign _zz_5490 = ($signed(_zz_17) - $signed(_zz_1813));
  assign _zz_5491 = _zz_5492;
  assign _zz_5492 = ($signed(_zz_5493) >>> _zz_1816);
  assign _zz_5493 = _zz_5494;
  assign _zz_5494 = ($signed(_zz_18) - $signed(_zz_1814));
  assign _zz_5495 = _zz_5496;
  assign _zz_5496 = ($signed(_zz_5497) >>> _zz_1817);
  assign _zz_5497 = _zz_5498;
  assign _zz_5498 = ($signed(_zz_17) + $signed(_zz_1813));
  assign _zz_5499 = _zz_5500;
  assign _zz_5500 = ($signed(_zz_5501) >>> _zz_1817);
  assign _zz_5501 = _zz_5502;
  assign _zz_5502 = ($signed(_zz_18) + $signed(_zz_1814));
  assign _zz_5503 = ($signed(twiddle_factor_table_0_real) + $signed(twiddle_factor_table_0_imag));
  assign _zz_5504 = fixTo_15_dout;
  assign _zz_5505 = ($signed(_zz_24) - $signed(_zz_23));
  assign _zz_5506 = ($signed(_zz_23) + $signed(_zz_24));
  assign _zz_5507 = _zz_5508[15 : 0];
  assign _zz_5508 = fixTo_17_dout;
  assign _zz_5509 = _zz_5510[15 : 0];
  assign _zz_5510 = fixTo_16_dout;
  assign _zz_5511 = _zz_5512;
  assign _zz_5512 = ($signed(_zz_5513) >>> _zz_1821);
  assign _zz_5513 = _zz_5514;
  assign _zz_5514 = ($signed(_zz_21) - $signed(_zz_1818));
  assign _zz_5515 = _zz_5516;
  assign _zz_5516 = ($signed(_zz_5517) >>> _zz_1821);
  assign _zz_5517 = _zz_5518;
  assign _zz_5518 = ($signed(_zz_22) - $signed(_zz_1819));
  assign _zz_5519 = _zz_5520;
  assign _zz_5520 = ($signed(_zz_5521) >>> _zz_1822);
  assign _zz_5521 = _zz_5522;
  assign _zz_5522 = ($signed(_zz_21) + $signed(_zz_1818));
  assign _zz_5523 = _zz_5524;
  assign _zz_5524 = ($signed(_zz_5525) >>> _zz_1822);
  assign _zz_5525 = _zz_5526;
  assign _zz_5526 = ($signed(_zz_22) + $signed(_zz_1819));
  assign _zz_5527 = ($signed(twiddle_factor_table_0_real) + $signed(twiddle_factor_table_0_imag));
  assign _zz_5528 = fixTo_18_dout;
  assign _zz_5529 = ($signed(_zz_28) - $signed(_zz_27));
  assign _zz_5530 = ($signed(_zz_27) + $signed(_zz_28));
  assign _zz_5531 = _zz_5532[15 : 0];
  assign _zz_5532 = fixTo_20_dout;
  assign _zz_5533 = _zz_5534[15 : 0];
  assign _zz_5534 = fixTo_19_dout;
  assign _zz_5535 = _zz_5536;
  assign _zz_5536 = ($signed(_zz_5537) >>> _zz_1826);
  assign _zz_5537 = _zz_5538;
  assign _zz_5538 = ($signed(_zz_25) - $signed(_zz_1823));
  assign _zz_5539 = _zz_5540;
  assign _zz_5540 = ($signed(_zz_5541) >>> _zz_1826);
  assign _zz_5541 = _zz_5542;
  assign _zz_5542 = ($signed(_zz_26) - $signed(_zz_1824));
  assign _zz_5543 = _zz_5544;
  assign _zz_5544 = ($signed(_zz_5545) >>> _zz_1827);
  assign _zz_5545 = _zz_5546;
  assign _zz_5546 = ($signed(_zz_25) + $signed(_zz_1823));
  assign _zz_5547 = _zz_5548;
  assign _zz_5548 = ($signed(_zz_5549) >>> _zz_1827);
  assign _zz_5549 = _zz_5550;
  assign _zz_5550 = ($signed(_zz_26) + $signed(_zz_1824));
  assign _zz_5551 = ($signed(twiddle_factor_table_0_real) + $signed(twiddle_factor_table_0_imag));
  assign _zz_5552 = fixTo_21_dout;
  assign _zz_5553 = ($signed(_zz_32) - $signed(_zz_31));
  assign _zz_5554 = ($signed(_zz_31) + $signed(_zz_32));
  assign _zz_5555 = _zz_5556[15 : 0];
  assign _zz_5556 = fixTo_23_dout;
  assign _zz_5557 = _zz_5558[15 : 0];
  assign _zz_5558 = fixTo_22_dout;
  assign _zz_5559 = _zz_5560;
  assign _zz_5560 = ($signed(_zz_5561) >>> _zz_1831);
  assign _zz_5561 = _zz_5562;
  assign _zz_5562 = ($signed(_zz_29) - $signed(_zz_1828));
  assign _zz_5563 = _zz_5564;
  assign _zz_5564 = ($signed(_zz_5565) >>> _zz_1831);
  assign _zz_5565 = _zz_5566;
  assign _zz_5566 = ($signed(_zz_30) - $signed(_zz_1829));
  assign _zz_5567 = _zz_5568;
  assign _zz_5568 = ($signed(_zz_5569) >>> _zz_1832);
  assign _zz_5569 = _zz_5570;
  assign _zz_5570 = ($signed(_zz_29) + $signed(_zz_1828));
  assign _zz_5571 = _zz_5572;
  assign _zz_5572 = ($signed(_zz_5573) >>> _zz_1832);
  assign _zz_5573 = _zz_5574;
  assign _zz_5574 = ($signed(_zz_30) + $signed(_zz_1829));
  assign _zz_5575 = ($signed(twiddle_factor_table_0_real) + $signed(twiddle_factor_table_0_imag));
  assign _zz_5576 = fixTo_24_dout;
  assign _zz_5577 = ($signed(_zz_36) - $signed(_zz_35));
  assign _zz_5578 = ($signed(_zz_35) + $signed(_zz_36));
  assign _zz_5579 = _zz_5580[15 : 0];
  assign _zz_5580 = fixTo_26_dout;
  assign _zz_5581 = _zz_5582[15 : 0];
  assign _zz_5582 = fixTo_25_dout;
  assign _zz_5583 = _zz_5584;
  assign _zz_5584 = ($signed(_zz_5585) >>> _zz_1836);
  assign _zz_5585 = _zz_5586;
  assign _zz_5586 = ($signed(_zz_33) - $signed(_zz_1833));
  assign _zz_5587 = _zz_5588;
  assign _zz_5588 = ($signed(_zz_5589) >>> _zz_1836);
  assign _zz_5589 = _zz_5590;
  assign _zz_5590 = ($signed(_zz_34) - $signed(_zz_1834));
  assign _zz_5591 = _zz_5592;
  assign _zz_5592 = ($signed(_zz_5593) >>> _zz_1837);
  assign _zz_5593 = _zz_5594;
  assign _zz_5594 = ($signed(_zz_33) + $signed(_zz_1833));
  assign _zz_5595 = _zz_5596;
  assign _zz_5596 = ($signed(_zz_5597) >>> _zz_1837);
  assign _zz_5597 = _zz_5598;
  assign _zz_5598 = ($signed(_zz_34) + $signed(_zz_1834));
  assign _zz_5599 = ($signed(twiddle_factor_table_0_real) + $signed(twiddle_factor_table_0_imag));
  assign _zz_5600 = fixTo_27_dout;
  assign _zz_5601 = ($signed(_zz_40) - $signed(_zz_39));
  assign _zz_5602 = ($signed(_zz_39) + $signed(_zz_40));
  assign _zz_5603 = _zz_5604[15 : 0];
  assign _zz_5604 = fixTo_29_dout;
  assign _zz_5605 = _zz_5606[15 : 0];
  assign _zz_5606 = fixTo_28_dout;
  assign _zz_5607 = _zz_5608;
  assign _zz_5608 = ($signed(_zz_5609) >>> _zz_1841);
  assign _zz_5609 = _zz_5610;
  assign _zz_5610 = ($signed(_zz_37) - $signed(_zz_1838));
  assign _zz_5611 = _zz_5612;
  assign _zz_5612 = ($signed(_zz_5613) >>> _zz_1841);
  assign _zz_5613 = _zz_5614;
  assign _zz_5614 = ($signed(_zz_38) - $signed(_zz_1839));
  assign _zz_5615 = _zz_5616;
  assign _zz_5616 = ($signed(_zz_5617) >>> _zz_1842);
  assign _zz_5617 = _zz_5618;
  assign _zz_5618 = ($signed(_zz_37) + $signed(_zz_1838));
  assign _zz_5619 = _zz_5620;
  assign _zz_5620 = ($signed(_zz_5621) >>> _zz_1842);
  assign _zz_5621 = _zz_5622;
  assign _zz_5622 = ($signed(_zz_38) + $signed(_zz_1839));
  assign _zz_5623 = ($signed(twiddle_factor_table_0_real) + $signed(twiddle_factor_table_0_imag));
  assign _zz_5624 = fixTo_30_dout;
  assign _zz_5625 = ($signed(_zz_44) - $signed(_zz_43));
  assign _zz_5626 = ($signed(_zz_43) + $signed(_zz_44));
  assign _zz_5627 = _zz_5628[15 : 0];
  assign _zz_5628 = fixTo_32_dout;
  assign _zz_5629 = _zz_5630[15 : 0];
  assign _zz_5630 = fixTo_31_dout;
  assign _zz_5631 = _zz_5632;
  assign _zz_5632 = ($signed(_zz_5633) >>> _zz_1846);
  assign _zz_5633 = _zz_5634;
  assign _zz_5634 = ($signed(_zz_41) - $signed(_zz_1843));
  assign _zz_5635 = _zz_5636;
  assign _zz_5636 = ($signed(_zz_5637) >>> _zz_1846);
  assign _zz_5637 = _zz_5638;
  assign _zz_5638 = ($signed(_zz_42) - $signed(_zz_1844));
  assign _zz_5639 = _zz_5640;
  assign _zz_5640 = ($signed(_zz_5641) >>> _zz_1847);
  assign _zz_5641 = _zz_5642;
  assign _zz_5642 = ($signed(_zz_41) + $signed(_zz_1843));
  assign _zz_5643 = _zz_5644;
  assign _zz_5644 = ($signed(_zz_5645) >>> _zz_1847);
  assign _zz_5645 = _zz_5646;
  assign _zz_5646 = ($signed(_zz_42) + $signed(_zz_1844));
  assign _zz_5647 = ($signed(twiddle_factor_table_0_real) + $signed(twiddle_factor_table_0_imag));
  assign _zz_5648 = fixTo_33_dout;
  assign _zz_5649 = ($signed(_zz_48) - $signed(_zz_47));
  assign _zz_5650 = ($signed(_zz_47) + $signed(_zz_48));
  assign _zz_5651 = _zz_5652[15 : 0];
  assign _zz_5652 = fixTo_35_dout;
  assign _zz_5653 = _zz_5654[15 : 0];
  assign _zz_5654 = fixTo_34_dout;
  assign _zz_5655 = _zz_5656;
  assign _zz_5656 = ($signed(_zz_5657) >>> _zz_1851);
  assign _zz_5657 = _zz_5658;
  assign _zz_5658 = ($signed(_zz_45) - $signed(_zz_1848));
  assign _zz_5659 = _zz_5660;
  assign _zz_5660 = ($signed(_zz_5661) >>> _zz_1851);
  assign _zz_5661 = _zz_5662;
  assign _zz_5662 = ($signed(_zz_46) - $signed(_zz_1849));
  assign _zz_5663 = _zz_5664;
  assign _zz_5664 = ($signed(_zz_5665) >>> _zz_1852);
  assign _zz_5665 = _zz_5666;
  assign _zz_5666 = ($signed(_zz_45) + $signed(_zz_1848));
  assign _zz_5667 = _zz_5668;
  assign _zz_5668 = ($signed(_zz_5669) >>> _zz_1852);
  assign _zz_5669 = _zz_5670;
  assign _zz_5670 = ($signed(_zz_46) + $signed(_zz_1849));
  assign _zz_5671 = ($signed(twiddle_factor_table_0_real) + $signed(twiddle_factor_table_0_imag));
  assign _zz_5672 = fixTo_36_dout;
  assign _zz_5673 = ($signed(_zz_52) - $signed(_zz_51));
  assign _zz_5674 = ($signed(_zz_51) + $signed(_zz_52));
  assign _zz_5675 = _zz_5676[15 : 0];
  assign _zz_5676 = fixTo_38_dout;
  assign _zz_5677 = _zz_5678[15 : 0];
  assign _zz_5678 = fixTo_37_dout;
  assign _zz_5679 = _zz_5680;
  assign _zz_5680 = ($signed(_zz_5681) >>> _zz_1856);
  assign _zz_5681 = _zz_5682;
  assign _zz_5682 = ($signed(_zz_49) - $signed(_zz_1853));
  assign _zz_5683 = _zz_5684;
  assign _zz_5684 = ($signed(_zz_5685) >>> _zz_1856);
  assign _zz_5685 = _zz_5686;
  assign _zz_5686 = ($signed(_zz_50) - $signed(_zz_1854));
  assign _zz_5687 = _zz_5688;
  assign _zz_5688 = ($signed(_zz_5689) >>> _zz_1857);
  assign _zz_5689 = _zz_5690;
  assign _zz_5690 = ($signed(_zz_49) + $signed(_zz_1853));
  assign _zz_5691 = _zz_5692;
  assign _zz_5692 = ($signed(_zz_5693) >>> _zz_1857);
  assign _zz_5693 = _zz_5694;
  assign _zz_5694 = ($signed(_zz_50) + $signed(_zz_1854));
  assign _zz_5695 = ($signed(twiddle_factor_table_0_real) + $signed(twiddle_factor_table_0_imag));
  assign _zz_5696 = fixTo_39_dout;
  assign _zz_5697 = ($signed(_zz_56) - $signed(_zz_55));
  assign _zz_5698 = ($signed(_zz_55) + $signed(_zz_56));
  assign _zz_5699 = _zz_5700[15 : 0];
  assign _zz_5700 = fixTo_41_dout;
  assign _zz_5701 = _zz_5702[15 : 0];
  assign _zz_5702 = fixTo_40_dout;
  assign _zz_5703 = _zz_5704;
  assign _zz_5704 = ($signed(_zz_5705) >>> _zz_1861);
  assign _zz_5705 = _zz_5706;
  assign _zz_5706 = ($signed(_zz_53) - $signed(_zz_1858));
  assign _zz_5707 = _zz_5708;
  assign _zz_5708 = ($signed(_zz_5709) >>> _zz_1861);
  assign _zz_5709 = _zz_5710;
  assign _zz_5710 = ($signed(_zz_54) - $signed(_zz_1859));
  assign _zz_5711 = _zz_5712;
  assign _zz_5712 = ($signed(_zz_5713) >>> _zz_1862);
  assign _zz_5713 = _zz_5714;
  assign _zz_5714 = ($signed(_zz_53) + $signed(_zz_1858));
  assign _zz_5715 = _zz_5716;
  assign _zz_5716 = ($signed(_zz_5717) >>> _zz_1862);
  assign _zz_5717 = _zz_5718;
  assign _zz_5718 = ($signed(_zz_54) + $signed(_zz_1859));
  assign _zz_5719 = ($signed(twiddle_factor_table_0_real) + $signed(twiddle_factor_table_0_imag));
  assign _zz_5720 = fixTo_42_dout;
  assign _zz_5721 = ($signed(_zz_60) - $signed(_zz_59));
  assign _zz_5722 = ($signed(_zz_59) + $signed(_zz_60));
  assign _zz_5723 = _zz_5724[15 : 0];
  assign _zz_5724 = fixTo_44_dout;
  assign _zz_5725 = _zz_5726[15 : 0];
  assign _zz_5726 = fixTo_43_dout;
  assign _zz_5727 = _zz_5728;
  assign _zz_5728 = ($signed(_zz_5729) >>> _zz_1866);
  assign _zz_5729 = _zz_5730;
  assign _zz_5730 = ($signed(_zz_57) - $signed(_zz_1863));
  assign _zz_5731 = _zz_5732;
  assign _zz_5732 = ($signed(_zz_5733) >>> _zz_1866);
  assign _zz_5733 = _zz_5734;
  assign _zz_5734 = ($signed(_zz_58) - $signed(_zz_1864));
  assign _zz_5735 = _zz_5736;
  assign _zz_5736 = ($signed(_zz_5737) >>> _zz_1867);
  assign _zz_5737 = _zz_5738;
  assign _zz_5738 = ($signed(_zz_57) + $signed(_zz_1863));
  assign _zz_5739 = _zz_5740;
  assign _zz_5740 = ($signed(_zz_5741) >>> _zz_1867);
  assign _zz_5741 = _zz_5742;
  assign _zz_5742 = ($signed(_zz_58) + $signed(_zz_1864));
  assign _zz_5743 = ($signed(twiddle_factor_table_0_real) + $signed(twiddle_factor_table_0_imag));
  assign _zz_5744 = fixTo_45_dout;
  assign _zz_5745 = ($signed(_zz_64) - $signed(_zz_63));
  assign _zz_5746 = ($signed(_zz_63) + $signed(_zz_64));
  assign _zz_5747 = _zz_5748[15 : 0];
  assign _zz_5748 = fixTo_47_dout;
  assign _zz_5749 = _zz_5750[15 : 0];
  assign _zz_5750 = fixTo_46_dout;
  assign _zz_5751 = _zz_5752;
  assign _zz_5752 = ($signed(_zz_5753) >>> _zz_1871);
  assign _zz_5753 = _zz_5754;
  assign _zz_5754 = ($signed(_zz_61) - $signed(_zz_1868));
  assign _zz_5755 = _zz_5756;
  assign _zz_5756 = ($signed(_zz_5757) >>> _zz_1871);
  assign _zz_5757 = _zz_5758;
  assign _zz_5758 = ($signed(_zz_62) - $signed(_zz_1869));
  assign _zz_5759 = _zz_5760;
  assign _zz_5760 = ($signed(_zz_5761) >>> _zz_1872);
  assign _zz_5761 = _zz_5762;
  assign _zz_5762 = ($signed(_zz_61) + $signed(_zz_1868));
  assign _zz_5763 = _zz_5764;
  assign _zz_5764 = ($signed(_zz_5765) >>> _zz_1872);
  assign _zz_5765 = _zz_5766;
  assign _zz_5766 = ($signed(_zz_62) + $signed(_zz_1869));
  assign _zz_5767 = ($signed(twiddle_factor_table_0_real) + $signed(twiddle_factor_table_0_imag));
  assign _zz_5768 = fixTo_48_dout;
  assign _zz_5769 = ($signed(_zz_68) - $signed(_zz_67));
  assign _zz_5770 = ($signed(_zz_67) + $signed(_zz_68));
  assign _zz_5771 = _zz_5772[15 : 0];
  assign _zz_5772 = fixTo_50_dout;
  assign _zz_5773 = _zz_5774[15 : 0];
  assign _zz_5774 = fixTo_49_dout;
  assign _zz_5775 = _zz_5776;
  assign _zz_5776 = ($signed(_zz_5777) >>> _zz_1876);
  assign _zz_5777 = _zz_5778;
  assign _zz_5778 = ($signed(_zz_65) - $signed(_zz_1873));
  assign _zz_5779 = _zz_5780;
  assign _zz_5780 = ($signed(_zz_5781) >>> _zz_1876);
  assign _zz_5781 = _zz_5782;
  assign _zz_5782 = ($signed(_zz_66) - $signed(_zz_1874));
  assign _zz_5783 = _zz_5784;
  assign _zz_5784 = ($signed(_zz_5785) >>> _zz_1877);
  assign _zz_5785 = _zz_5786;
  assign _zz_5786 = ($signed(_zz_65) + $signed(_zz_1873));
  assign _zz_5787 = _zz_5788;
  assign _zz_5788 = ($signed(_zz_5789) >>> _zz_1877);
  assign _zz_5789 = _zz_5790;
  assign _zz_5790 = ($signed(_zz_66) + $signed(_zz_1874));
  assign _zz_5791 = ($signed(twiddle_factor_table_0_real) + $signed(twiddle_factor_table_0_imag));
  assign _zz_5792 = fixTo_51_dout;
  assign _zz_5793 = ($signed(_zz_72) - $signed(_zz_71));
  assign _zz_5794 = ($signed(_zz_71) + $signed(_zz_72));
  assign _zz_5795 = _zz_5796[15 : 0];
  assign _zz_5796 = fixTo_53_dout;
  assign _zz_5797 = _zz_5798[15 : 0];
  assign _zz_5798 = fixTo_52_dout;
  assign _zz_5799 = _zz_5800;
  assign _zz_5800 = ($signed(_zz_5801) >>> _zz_1881);
  assign _zz_5801 = _zz_5802;
  assign _zz_5802 = ($signed(_zz_69) - $signed(_zz_1878));
  assign _zz_5803 = _zz_5804;
  assign _zz_5804 = ($signed(_zz_5805) >>> _zz_1881);
  assign _zz_5805 = _zz_5806;
  assign _zz_5806 = ($signed(_zz_70) - $signed(_zz_1879));
  assign _zz_5807 = _zz_5808;
  assign _zz_5808 = ($signed(_zz_5809) >>> _zz_1882);
  assign _zz_5809 = _zz_5810;
  assign _zz_5810 = ($signed(_zz_69) + $signed(_zz_1878));
  assign _zz_5811 = _zz_5812;
  assign _zz_5812 = ($signed(_zz_5813) >>> _zz_1882);
  assign _zz_5813 = _zz_5814;
  assign _zz_5814 = ($signed(_zz_70) + $signed(_zz_1879));
  assign _zz_5815 = ($signed(twiddle_factor_table_0_real) + $signed(twiddle_factor_table_0_imag));
  assign _zz_5816 = fixTo_54_dout;
  assign _zz_5817 = ($signed(_zz_76) - $signed(_zz_75));
  assign _zz_5818 = ($signed(_zz_75) + $signed(_zz_76));
  assign _zz_5819 = _zz_5820[15 : 0];
  assign _zz_5820 = fixTo_56_dout;
  assign _zz_5821 = _zz_5822[15 : 0];
  assign _zz_5822 = fixTo_55_dout;
  assign _zz_5823 = _zz_5824;
  assign _zz_5824 = ($signed(_zz_5825) >>> _zz_1886);
  assign _zz_5825 = _zz_5826;
  assign _zz_5826 = ($signed(_zz_73) - $signed(_zz_1883));
  assign _zz_5827 = _zz_5828;
  assign _zz_5828 = ($signed(_zz_5829) >>> _zz_1886);
  assign _zz_5829 = _zz_5830;
  assign _zz_5830 = ($signed(_zz_74) - $signed(_zz_1884));
  assign _zz_5831 = _zz_5832;
  assign _zz_5832 = ($signed(_zz_5833) >>> _zz_1887);
  assign _zz_5833 = _zz_5834;
  assign _zz_5834 = ($signed(_zz_73) + $signed(_zz_1883));
  assign _zz_5835 = _zz_5836;
  assign _zz_5836 = ($signed(_zz_5837) >>> _zz_1887);
  assign _zz_5837 = _zz_5838;
  assign _zz_5838 = ($signed(_zz_74) + $signed(_zz_1884));
  assign _zz_5839 = ($signed(twiddle_factor_table_0_real) + $signed(twiddle_factor_table_0_imag));
  assign _zz_5840 = fixTo_57_dout;
  assign _zz_5841 = ($signed(_zz_80) - $signed(_zz_79));
  assign _zz_5842 = ($signed(_zz_79) + $signed(_zz_80));
  assign _zz_5843 = _zz_5844[15 : 0];
  assign _zz_5844 = fixTo_59_dout;
  assign _zz_5845 = _zz_5846[15 : 0];
  assign _zz_5846 = fixTo_58_dout;
  assign _zz_5847 = _zz_5848;
  assign _zz_5848 = ($signed(_zz_5849) >>> _zz_1891);
  assign _zz_5849 = _zz_5850;
  assign _zz_5850 = ($signed(_zz_77) - $signed(_zz_1888));
  assign _zz_5851 = _zz_5852;
  assign _zz_5852 = ($signed(_zz_5853) >>> _zz_1891);
  assign _zz_5853 = _zz_5854;
  assign _zz_5854 = ($signed(_zz_78) - $signed(_zz_1889));
  assign _zz_5855 = _zz_5856;
  assign _zz_5856 = ($signed(_zz_5857) >>> _zz_1892);
  assign _zz_5857 = _zz_5858;
  assign _zz_5858 = ($signed(_zz_77) + $signed(_zz_1888));
  assign _zz_5859 = _zz_5860;
  assign _zz_5860 = ($signed(_zz_5861) >>> _zz_1892);
  assign _zz_5861 = _zz_5862;
  assign _zz_5862 = ($signed(_zz_78) + $signed(_zz_1889));
  assign _zz_5863 = ($signed(twiddle_factor_table_0_real) + $signed(twiddle_factor_table_0_imag));
  assign _zz_5864 = fixTo_60_dout;
  assign _zz_5865 = ($signed(_zz_84) - $signed(_zz_83));
  assign _zz_5866 = ($signed(_zz_83) + $signed(_zz_84));
  assign _zz_5867 = _zz_5868[15 : 0];
  assign _zz_5868 = fixTo_62_dout;
  assign _zz_5869 = _zz_5870[15 : 0];
  assign _zz_5870 = fixTo_61_dout;
  assign _zz_5871 = _zz_5872;
  assign _zz_5872 = ($signed(_zz_5873) >>> _zz_1896);
  assign _zz_5873 = _zz_5874;
  assign _zz_5874 = ($signed(_zz_81) - $signed(_zz_1893));
  assign _zz_5875 = _zz_5876;
  assign _zz_5876 = ($signed(_zz_5877) >>> _zz_1896);
  assign _zz_5877 = _zz_5878;
  assign _zz_5878 = ($signed(_zz_82) - $signed(_zz_1894));
  assign _zz_5879 = _zz_5880;
  assign _zz_5880 = ($signed(_zz_5881) >>> _zz_1897);
  assign _zz_5881 = _zz_5882;
  assign _zz_5882 = ($signed(_zz_81) + $signed(_zz_1893));
  assign _zz_5883 = _zz_5884;
  assign _zz_5884 = ($signed(_zz_5885) >>> _zz_1897);
  assign _zz_5885 = _zz_5886;
  assign _zz_5886 = ($signed(_zz_82) + $signed(_zz_1894));
  assign _zz_5887 = ($signed(twiddle_factor_table_0_real) + $signed(twiddle_factor_table_0_imag));
  assign _zz_5888 = fixTo_63_dout;
  assign _zz_5889 = ($signed(_zz_88) - $signed(_zz_87));
  assign _zz_5890 = ($signed(_zz_87) + $signed(_zz_88));
  assign _zz_5891 = _zz_5892[15 : 0];
  assign _zz_5892 = fixTo_65_dout;
  assign _zz_5893 = _zz_5894[15 : 0];
  assign _zz_5894 = fixTo_64_dout;
  assign _zz_5895 = _zz_5896;
  assign _zz_5896 = ($signed(_zz_5897) >>> _zz_1901);
  assign _zz_5897 = _zz_5898;
  assign _zz_5898 = ($signed(_zz_85) - $signed(_zz_1898));
  assign _zz_5899 = _zz_5900;
  assign _zz_5900 = ($signed(_zz_5901) >>> _zz_1901);
  assign _zz_5901 = _zz_5902;
  assign _zz_5902 = ($signed(_zz_86) - $signed(_zz_1899));
  assign _zz_5903 = _zz_5904;
  assign _zz_5904 = ($signed(_zz_5905) >>> _zz_1902);
  assign _zz_5905 = _zz_5906;
  assign _zz_5906 = ($signed(_zz_85) + $signed(_zz_1898));
  assign _zz_5907 = _zz_5908;
  assign _zz_5908 = ($signed(_zz_5909) >>> _zz_1902);
  assign _zz_5909 = _zz_5910;
  assign _zz_5910 = ($signed(_zz_86) + $signed(_zz_1899));
  assign _zz_5911 = ($signed(twiddle_factor_table_0_real) + $signed(twiddle_factor_table_0_imag));
  assign _zz_5912 = fixTo_66_dout;
  assign _zz_5913 = ($signed(_zz_92) - $signed(_zz_91));
  assign _zz_5914 = ($signed(_zz_91) + $signed(_zz_92));
  assign _zz_5915 = _zz_5916[15 : 0];
  assign _zz_5916 = fixTo_68_dout;
  assign _zz_5917 = _zz_5918[15 : 0];
  assign _zz_5918 = fixTo_67_dout;
  assign _zz_5919 = _zz_5920;
  assign _zz_5920 = ($signed(_zz_5921) >>> _zz_1906);
  assign _zz_5921 = _zz_5922;
  assign _zz_5922 = ($signed(_zz_89) - $signed(_zz_1903));
  assign _zz_5923 = _zz_5924;
  assign _zz_5924 = ($signed(_zz_5925) >>> _zz_1906);
  assign _zz_5925 = _zz_5926;
  assign _zz_5926 = ($signed(_zz_90) - $signed(_zz_1904));
  assign _zz_5927 = _zz_5928;
  assign _zz_5928 = ($signed(_zz_5929) >>> _zz_1907);
  assign _zz_5929 = _zz_5930;
  assign _zz_5930 = ($signed(_zz_89) + $signed(_zz_1903));
  assign _zz_5931 = _zz_5932;
  assign _zz_5932 = ($signed(_zz_5933) >>> _zz_1907);
  assign _zz_5933 = _zz_5934;
  assign _zz_5934 = ($signed(_zz_90) + $signed(_zz_1904));
  assign _zz_5935 = ($signed(twiddle_factor_table_0_real) + $signed(twiddle_factor_table_0_imag));
  assign _zz_5936 = fixTo_69_dout;
  assign _zz_5937 = ($signed(_zz_96) - $signed(_zz_95));
  assign _zz_5938 = ($signed(_zz_95) + $signed(_zz_96));
  assign _zz_5939 = _zz_5940[15 : 0];
  assign _zz_5940 = fixTo_71_dout;
  assign _zz_5941 = _zz_5942[15 : 0];
  assign _zz_5942 = fixTo_70_dout;
  assign _zz_5943 = _zz_5944;
  assign _zz_5944 = ($signed(_zz_5945) >>> _zz_1911);
  assign _zz_5945 = _zz_5946;
  assign _zz_5946 = ($signed(_zz_93) - $signed(_zz_1908));
  assign _zz_5947 = _zz_5948;
  assign _zz_5948 = ($signed(_zz_5949) >>> _zz_1911);
  assign _zz_5949 = _zz_5950;
  assign _zz_5950 = ($signed(_zz_94) - $signed(_zz_1909));
  assign _zz_5951 = _zz_5952;
  assign _zz_5952 = ($signed(_zz_5953) >>> _zz_1912);
  assign _zz_5953 = _zz_5954;
  assign _zz_5954 = ($signed(_zz_93) + $signed(_zz_1908));
  assign _zz_5955 = _zz_5956;
  assign _zz_5956 = ($signed(_zz_5957) >>> _zz_1912);
  assign _zz_5957 = _zz_5958;
  assign _zz_5958 = ($signed(_zz_94) + $signed(_zz_1909));
  assign _zz_5959 = ($signed(twiddle_factor_table_0_real) + $signed(twiddle_factor_table_0_imag));
  assign _zz_5960 = fixTo_72_dout;
  assign _zz_5961 = ($signed(_zz_100) - $signed(_zz_99));
  assign _zz_5962 = ($signed(_zz_99) + $signed(_zz_100));
  assign _zz_5963 = _zz_5964[15 : 0];
  assign _zz_5964 = fixTo_74_dout;
  assign _zz_5965 = _zz_5966[15 : 0];
  assign _zz_5966 = fixTo_73_dout;
  assign _zz_5967 = _zz_5968;
  assign _zz_5968 = ($signed(_zz_5969) >>> _zz_1916);
  assign _zz_5969 = _zz_5970;
  assign _zz_5970 = ($signed(_zz_97) - $signed(_zz_1913));
  assign _zz_5971 = _zz_5972;
  assign _zz_5972 = ($signed(_zz_5973) >>> _zz_1916);
  assign _zz_5973 = _zz_5974;
  assign _zz_5974 = ($signed(_zz_98) - $signed(_zz_1914));
  assign _zz_5975 = _zz_5976;
  assign _zz_5976 = ($signed(_zz_5977) >>> _zz_1917);
  assign _zz_5977 = _zz_5978;
  assign _zz_5978 = ($signed(_zz_97) + $signed(_zz_1913));
  assign _zz_5979 = _zz_5980;
  assign _zz_5980 = ($signed(_zz_5981) >>> _zz_1917);
  assign _zz_5981 = _zz_5982;
  assign _zz_5982 = ($signed(_zz_98) + $signed(_zz_1914));
  assign _zz_5983 = ($signed(twiddle_factor_table_0_real) + $signed(twiddle_factor_table_0_imag));
  assign _zz_5984 = fixTo_75_dout;
  assign _zz_5985 = ($signed(_zz_104) - $signed(_zz_103));
  assign _zz_5986 = ($signed(_zz_103) + $signed(_zz_104));
  assign _zz_5987 = _zz_5988[15 : 0];
  assign _zz_5988 = fixTo_77_dout;
  assign _zz_5989 = _zz_5990[15 : 0];
  assign _zz_5990 = fixTo_76_dout;
  assign _zz_5991 = _zz_5992;
  assign _zz_5992 = ($signed(_zz_5993) >>> _zz_1921);
  assign _zz_5993 = _zz_5994;
  assign _zz_5994 = ($signed(_zz_101) - $signed(_zz_1918));
  assign _zz_5995 = _zz_5996;
  assign _zz_5996 = ($signed(_zz_5997) >>> _zz_1921);
  assign _zz_5997 = _zz_5998;
  assign _zz_5998 = ($signed(_zz_102) - $signed(_zz_1919));
  assign _zz_5999 = _zz_6000;
  assign _zz_6000 = ($signed(_zz_6001) >>> _zz_1922);
  assign _zz_6001 = _zz_6002;
  assign _zz_6002 = ($signed(_zz_101) + $signed(_zz_1918));
  assign _zz_6003 = _zz_6004;
  assign _zz_6004 = ($signed(_zz_6005) >>> _zz_1922);
  assign _zz_6005 = _zz_6006;
  assign _zz_6006 = ($signed(_zz_102) + $signed(_zz_1919));
  assign _zz_6007 = ($signed(twiddle_factor_table_0_real) + $signed(twiddle_factor_table_0_imag));
  assign _zz_6008 = fixTo_78_dout;
  assign _zz_6009 = ($signed(_zz_108) - $signed(_zz_107));
  assign _zz_6010 = ($signed(_zz_107) + $signed(_zz_108));
  assign _zz_6011 = _zz_6012[15 : 0];
  assign _zz_6012 = fixTo_80_dout;
  assign _zz_6013 = _zz_6014[15 : 0];
  assign _zz_6014 = fixTo_79_dout;
  assign _zz_6015 = _zz_6016;
  assign _zz_6016 = ($signed(_zz_6017) >>> _zz_1926);
  assign _zz_6017 = _zz_6018;
  assign _zz_6018 = ($signed(_zz_105) - $signed(_zz_1923));
  assign _zz_6019 = _zz_6020;
  assign _zz_6020 = ($signed(_zz_6021) >>> _zz_1926);
  assign _zz_6021 = _zz_6022;
  assign _zz_6022 = ($signed(_zz_106) - $signed(_zz_1924));
  assign _zz_6023 = _zz_6024;
  assign _zz_6024 = ($signed(_zz_6025) >>> _zz_1927);
  assign _zz_6025 = _zz_6026;
  assign _zz_6026 = ($signed(_zz_105) + $signed(_zz_1923));
  assign _zz_6027 = _zz_6028;
  assign _zz_6028 = ($signed(_zz_6029) >>> _zz_1927);
  assign _zz_6029 = _zz_6030;
  assign _zz_6030 = ($signed(_zz_106) + $signed(_zz_1924));
  assign _zz_6031 = ($signed(twiddle_factor_table_0_real) + $signed(twiddle_factor_table_0_imag));
  assign _zz_6032 = fixTo_81_dout;
  assign _zz_6033 = ($signed(_zz_112) - $signed(_zz_111));
  assign _zz_6034 = ($signed(_zz_111) + $signed(_zz_112));
  assign _zz_6035 = _zz_6036[15 : 0];
  assign _zz_6036 = fixTo_83_dout;
  assign _zz_6037 = _zz_6038[15 : 0];
  assign _zz_6038 = fixTo_82_dout;
  assign _zz_6039 = _zz_6040;
  assign _zz_6040 = ($signed(_zz_6041) >>> _zz_1931);
  assign _zz_6041 = _zz_6042;
  assign _zz_6042 = ($signed(_zz_109) - $signed(_zz_1928));
  assign _zz_6043 = _zz_6044;
  assign _zz_6044 = ($signed(_zz_6045) >>> _zz_1931);
  assign _zz_6045 = _zz_6046;
  assign _zz_6046 = ($signed(_zz_110) - $signed(_zz_1929));
  assign _zz_6047 = _zz_6048;
  assign _zz_6048 = ($signed(_zz_6049) >>> _zz_1932);
  assign _zz_6049 = _zz_6050;
  assign _zz_6050 = ($signed(_zz_109) + $signed(_zz_1928));
  assign _zz_6051 = _zz_6052;
  assign _zz_6052 = ($signed(_zz_6053) >>> _zz_1932);
  assign _zz_6053 = _zz_6054;
  assign _zz_6054 = ($signed(_zz_110) + $signed(_zz_1929));
  assign _zz_6055 = ($signed(twiddle_factor_table_0_real) + $signed(twiddle_factor_table_0_imag));
  assign _zz_6056 = fixTo_84_dout;
  assign _zz_6057 = ($signed(_zz_116) - $signed(_zz_115));
  assign _zz_6058 = ($signed(_zz_115) + $signed(_zz_116));
  assign _zz_6059 = _zz_6060[15 : 0];
  assign _zz_6060 = fixTo_86_dout;
  assign _zz_6061 = _zz_6062[15 : 0];
  assign _zz_6062 = fixTo_85_dout;
  assign _zz_6063 = _zz_6064;
  assign _zz_6064 = ($signed(_zz_6065) >>> _zz_1936);
  assign _zz_6065 = _zz_6066;
  assign _zz_6066 = ($signed(_zz_113) - $signed(_zz_1933));
  assign _zz_6067 = _zz_6068;
  assign _zz_6068 = ($signed(_zz_6069) >>> _zz_1936);
  assign _zz_6069 = _zz_6070;
  assign _zz_6070 = ($signed(_zz_114) - $signed(_zz_1934));
  assign _zz_6071 = _zz_6072;
  assign _zz_6072 = ($signed(_zz_6073) >>> _zz_1937);
  assign _zz_6073 = _zz_6074;
  assign _zz_6074 = ($signed(_zz_113) + $signed(_zz_1933));
  assign _zz_6075 = _zz_6076;
  assign _zz_6076 = ($signed(_zz_6077) >>> _zz_1937);
  assign _zz_6077 = _zz_6078;
  assign _zz_6078 = ($signed(_zz_114) + $signed(_zz_1934));
  assign _zz_6079 = ($signed(twiddle_factor_table_0_real) + $signed(twiddle_factor_table_0_imag));
  assign _zz_6080 = fixTo_87_dout;
  assign _zz_6081 = ($signed(_zz_120) - $signed(_zz_119));
  assign _zz_6082 = ($signed(_zz_119) + $signed(_zz_120));
  assign _zz_6083 = _zz_6084[15 : 0];
  assign _zz_6084 = fixTo_89_dout;
  assign _zz_6085 = _zz_6086[15 : 0];
  assign _zz_6086 = fixTo_88_dout;
  assign _zz_6087 = _zz_6088;
  assign _zz_6088 = ($signed(_zz_6089) >>> _zz_1941);
  assign _zz_6089 = _zz_6090;
  assign _zz_6090 = ($signed(_zz_117) - $signed(_zz_1938));
  assign _zz_6091 = _zz_6092;
  assign _zz_6092 = ($signed(_zz_6093) >>> _zz_1941);
  assign _zz_6093 = _zz_6094;
  assign _zz_6094 = ($signed(_zz_118) - $signed(_zz_1939));
  assign _zz_6095 = _zz_6096;
  assign _zz_6096 = ($signed(_zz_6097) >>> _zz_1942);
  assign _zz_6097 = _zz_6098;
  assign _zz_6098 = ($signed(_zz_117) + $signed(_zz_1938));
  assign _zz_6099 = _zz_6100;
  assign _zz_6100 = ($signed(_zz_6101) >>> _zz_1942);
  assign _zz_6101 = _zz_6102;
  assign _zz_6102 = ($signed(_zz_118) + $signed(_zz_1939));
  assign _zz_6103 = ($signed(twiddle_factor_table_0_real) + $signed(twiddle_factor_table_0_imag));
  assign _zz_6104 = fixTo_90_dout;
  assign _zz_6105 = ($signed(_zz_124) - $signed(_zz_123));
  assign _zz_6106 = ($signed(_zz_123) + $signed(_zz_124));
  assign _zz_6107 = _zz_6108[15 : 0];
  assign _zz_6108 = fixTo_92_dout;
  assign _zz_6109 = _zz_6110[15 : 0];
  assign _zz_6110 = fixTo_91_dout;
  assign _zz_6111 = _zz_6112;
  assign _zz_6112 = ($signed(_zz_6113) >>> _zz_1946);
  assign _zz_6113 = _zz_6114;
  assign _zz_6114 = ($signed(_zz_121) - $signed(_zz_1943));
  assign _zz_6115 = _zz_6116;
  assign _zz_6116 = ($signed(_zz_6117) >>> _zz_1946);
  assign _zz_6117 = _zz_6118;
  assign _zz_6118 = ($signed(_zz_122) - $signed(_zz_1944));
  assign _zz_6119 = _zz_6120;
  assign _zz_6120 = ($signed(_zz_6121) >>> _zz_1947);
  assign _zz_6121 = _zz_6122;
  assign _zz_6122 = ($signed(_zz_121) + $signed(_zz_1943));
  assign _zz_6123 = _zz_6124;
  assign _zz_6124 = ($signed(_zz_6125) >>> _zz_1947);
  assign _zz_6125 = _zz_6126;
  assign _zz_6126 = ($signed(_zz_122) + $signed(_zz_1944));
  assign _zz_6127 = ($signed(twiddle_factor_table_0_real) + $signed(twiddle_factor_table_0_imag));
  assign _zz_6128 = fixTo_93_dout;
  assign _zz_6129 = ($signed(_zz_128) - $signed(_zz_127));
  assign _zz_6130 = ($signed(_zz_127) + $signed(_zz_128));
  assign _zz_6131 = _zz_6132[15 : 0];
  assign _zz_6132 = fixTo_95_dout;
  assign _zz_6133 = _zz_6134[15 : 0];
  assign _zz_6134 = fixTo_94_dout;
  assign _zz_6135 = _zz_6136;
  assign _zz_6136 = ($signed(_zz_6137) >>> _zz_1951);
  assign _zz_6137 = _zz_6138;
  assign _zz_6138 = ($signed(_zz_125) - $signed(_zz_1948));
  assign _zz_6139 = _zz_6140;
  assign _zz_6140 = ($signed(_zz_6141) >>> _zz_1951);
  assign _zz_6141 = _zz_6142;
  assign _zz_6142 = ($signed(_zz_126) - $signed(_zz_1949));
  assign _zz_6143 = _zz_6144;
  assign _zz_6144 = ($signed(_zz_6145) >>> _zz_1952);
  assign _zz_6145 = _zz_6146;
  assign _zz_6146 = ($signed(_zz_125) + $signed(_zz_1948));
  assign _zz_6147 = _zz_6148;
  assign _zz_6148 = ($signed(_zz_6149) >>> _zz_1952);
  assign _zz_6149 = _zz_6150;
  assign _zz_6150 = ($signed(_zz_126) + $signed(_zz_1949));
  assign _zz_6151 = ($signed(twiddle_factor_table_0_real) + $signed(twiddle_factor_table_0_imag));
  assign _zz_6152 = fixTo_96_dout;
  assign _zz_6153 = ($signed(_zz_132) - $signed(_zz_131));
  assign _zz_6154 = ($signed(_zz_131) + $signed(_zz_132));
  assign _zz_6155 = _zz_6156[15 : 0];
  assign _zz_6156 = fixTo_98_dout;
  assign _zz_6157 = _zz_6158[15 : 0];
  assign _zz_6158 = fixTo_97_dout;
  assign _zz_6159 = _zz_6160;
  assign _zz_6160 = ($signed(_zz_6161) >>> _zz_1956);
  assign _zz_6161 = _zz_6162;
  assign _zz_6162 = ($signed(_zz_129) - $signed(_zz_1953));
  assign _zz_6163 = _zz_6164;
  assign _zz_6164 = ($signed(_zz_6165) >>> _zz_1956);
  assign _zz_6165 = _zz_6166;
  assign _zz_6166 = ($signed(_zz_130) - $signed(_zz_1954));
  assign _zz_6167 = _zz_6168;
  assign _zz_6168 = ($signed(_zz_6169) >>> _zz_1957);
  assign _zz_6169 = _zz_6170;
  assign _zz_6170 = ($signed(_zz_129) + $signed(_zz_1953));
  assign _zz_6171 = _zz_6172;
  assign _zz_6172 = ($signed(_zz_6173) >>> _zz_1957);
  assign _zz_6173 = _zz_6174;
  assign _zz_6174 = ($signed(_zz_130) + $signed(_zz_1954));
  assign _zz_6175 = ($signed(twiddle_factor_table_0_real) + $signed(twiddle_factor_table_0_imag));
  assign _zz_6176 = fixTo_99_dout;
  assign _zz_6177 = ($signed(_zz_136) - $signed(_zz_135));
  assign _zz_6178 = ($signed(_zz_135) + $signed(_zz_136));
  assign _zz_6179 = _zz_6180[15 : 0];
  assign _zz_6180 = fixTo_101_dout;
  assign _zz_6181 = _zz_6182[15 : 0];
  assign _zz_6182 = fixTo_100_dout;
  assign _zz_6183 = _zz_6184;
  assign _zz_6184 = ($signed(_zz_6185) >>> _zz_1961);
  assign _zz_6185 = _zz_6186;
  assign _zz_6186 = ($signed(_zz_133) - $signed(_zz_1958));
  assign _zz_6187 = _zz_6188;
  assign _zz_6188 = ($signed(_zz_6189) >>> _zz_1961);
  assign _zz_6189 = _zz_6190;
  assign _zz_6190 = ($signed(_zz_134) - $signed(_zz_1959));
  assign _zz_6191 = _zz_6192;
  assign _zz_6192 = ($signed(_zz_6193) >>> _zz_1962);
  assign _zz_6193 = _zz_6194;
  assign _zz_6194 = ($signed(_zz_133) + $signed(_zz_1958));
  assign _zz_6195 = _zz_6196;
  assign _zz_6196 = ($signed(_zz_6197) >>> _zz_1962);
  assign _zz_6197 = _zz_6198;
  assign _zz_6198 = ($signed(_zz_134) + $signed(_zz_1959));
  assign _zz_6199 = ($signed(twiddle_factor_table_0_real) + $signed(twiddle_factor_table_0_imag));
  assign _zz_6200 = fixTo_102_dout;
  assign _zz_6201 = ($signed(_zz_140) - $signed(_zz_139));
  assign _zz_6202 = ($signed(_zz_139) + $signed(_zz_140));
  assign _zz_6203 = _zz_6204[15 : 0];
  assign _zz_6204 = fixTo_104_dout;
  assign _zz_6205 = _zz_6206[15 : 0];
  assign _zz_6206 = fixTo_103_dout;
  assign _zz_6207 = _zz_6208;
  assign _zz_6208 = ($signed(_zz_6209) >>> _zz_1966);
  assign _zz_6209 = _zz_6210;
  assign _zz_6210 = ($signed(_zz_137) - $signed(_zz_1963));
  assign _zz_6211 = _zz_6212;
  assign _zz_6212 = ($signed(_zz_6213) >>> _zz_1966);
  assign _zz_6213 = _zz_6214;
  assign _zz_6214 = ($signed(_zz_138) - $signed(_zz_1964));
  assign _zz_6215 = _zz_6216;
  assign _zz_6216 = ($signed(_zz_6217) >>> _zz_1967);
  assign _zz_6217 = _zz_6218;
  assign _zz_6218 = ($signed(_zz_137) + $signed(_zz_1963));
  assign _zz_6219 = _zz_6220;
  assign _zz_6220 = ($signed(_zz_6221) >>> _zz_1967);
  assign _zz_6221 = _zz_6222;
  assign _zz_6222 = ($signed(_zz_138) + $signed(_zz_1964));
  assign _zz_6223 = ($signed(twiddle_factor_table_0_real) + $signed(twiddle_factor_table_0_imag));
  assign _zz_6224 = fixTo_105_dout;
  assign _zz_6225 = ($signed(_zz_144) - $signed(_zz_143));
  assign _zz_6226 = ($signed(_zz_143) + $signed(_zz_144));
  assign _zz_6227 = _zz_6228[15 : 0];
  assign _zz_6228 = fixTo_107_dout;
  assign _zz_6229 = _zz_6230[15 : 0];
  assign _zz_6230 = fixTo_106_dout;
  assign _zz_6231 = _zz_6232;
  assign _zz_6232 = ($signed(_zz_6233) >>> _zz_1971);
  assign _zz_6233 = _zz_6234;
  assign _zz_6234 = ($signed(_zz_141) - $signed(_zz_1968));
  assign _zz_6235 = _zz_6236;
  assign _zz_6236 = ($signed(_zz_6237) >>> _zz_1971);
  assign _zz_6237 = _zz_6238;
  assign _zz_6238 = ($signed(_zz_142) - $signed(_zz_1969));
  assign _zz_6239 = _zz_6240;
  assign _zz_6240 = ($signed(_zz_6241) >>> _zz_1972);
  assign _zz_6241 = _zz_6242;
  assign _zz_6242 = ($signed(_zz_141) + $signed(_zz_1968));
  assign _zz_6243 = _zz_6244;
  assign _zz_6244 = ($signed(_zz_6245) >>> _zz_1972);
  assign _zz_6245 = _zz_6246;
  assign _zz_6246 = ($signed(_zz_142) + $signed(_zz_1969));
  assign _zz_6247 = ($signed(twiddle_factor_table_0_real) + $signed(twiddle_factor_table_0_imag));
  assign _zz_6248 = fixTo_108_dout;
  assign _zz_6249 = ($signed(_zz_148) - $signed(_zz_147));
  assign _zz_6250 = ($signed(_zz_147) + $signed(_zz_148));
  assign _zz_6251 = _zz_6252[15 : 0];
  assign _zz_6252 = fixTo_110_dout;
  assign _zz_6253 = _zz_6254[15 : 0];
  assign _zz_6254 = fixTo_109_dout;
  assign _zz_6255 = _zz_6256;
  assign _zz_6256 = ($signed(_zz_6257) >>> _zz_1976);
  assign _zz_6257 = _zz_6258;
  assign _zz_6258 = ($signed(_zz_145) - $signed(_zz_1973));
  assign _zz_6259 = _zz_6260;
  assign _zz_6260 = ($signed(_zz_6261) >>> _zz_1976);
  assign _zz_6261 = _zz_6262;
  assign _zz_6262 = ($signed(_zz_146) - $signed(_zz_1974));
  assign _zz_6263 = _zz_6264;
  assign _zz_6264 = ($signed(_zz_6265) >>> _zz_1977);
  assign _zz_6265 = _zz_6266;
  assign _zz_6266 = ($signed(_zz_145) + $signed(_zz_1973));
  assign _zz_6267 = _zz_6268;
  assign _zz_6268 = ($signed(_zz_6269) >>> _zz_1977);
  assign _zz_6269 = _zz_6270;
  assign _zz_6270 = ($signed(_zz_146) + $signed(_zz_1974));
  assign _zz_6271 = ($signed(twiddle_factor_table_0_real) + $signed(twiddle_factor_table_0_imag));
  assign _zz_6272 = fixTo_111_dout;
  assign _zz_6273 = ($signed(_zz_152) - $signed(_zz_151));
  assign _zz_6274 = ($signed(_zz_151) + $signed(_zz_152));
  assign _zz_6275 = _zz_6276[15 : 0];
  assign _zz_6276 = fixTo_113_dout;
  assign _zz_6277 = _zz_6278[15 : 0];
  assign _zz_6278 = fixTo_112_dout;
  assign _zz_6279 = _zz_6280;
  assign _zz_6280 = ($signed(_zz_6281) >>> _zz_1981);
  assign _zz_6281 = _zz_6282;
  assign _zz_6282 = ($signed(_zz_149) - $signed(_zz_1978));
  assign _zz_6283 = _zz_6284;
  assign _zz_6284 = ($signed(_zz_6285) >>> _zz_1981);
  assign _zz_6285 = _zz_6286;
  assign _zz_6286 = ($signed(_zz_150) - $signed(_zz_1979));
  assign _zz_6287 = _zz_6288;
  assign _zz_6288 = ($signed(_zz_6289) >>> _zz_1982);
  assign _zz_6289 = _zz_6290;
  assign _zz_6290 = ($signed(_zz_149) + $signed(_zz_1978));
  assign _zz_6291 = _zz_6292;
  assign _zz_6292 = ($signed(_zz_6293) >>> _zz_1982);
  assign _zz_6293 = _zz_6294;
  assign _zz_6294 = ($signed(_zz_150) + $signed(_zz_1979));
  assign _zz_6295 = ($signed(twiddle_factor_table_0_real) + $signed(twiddle_factor_table_0_imag));
  assign _zz_6296 = fixTo_114_dout;
  assign _zz_6297 = ($signed(_zz_156) - $signed(_zz_155));
  assign _zz_6298 = ($signed(_zz_155) + $signed(_zz_156));
  assign _zz_6299 = _zz_6300[15 : 0];
  assign _zz_6300 = fixTo_116_dout;
  assign _zz_6301 = _zz_6302[15 : 0];
  assign _zz_6302 = fixTo_115_dout;
  assign _zz_6303 = _zz_6304;
  assign _zz_6304 = ($signed(_zz_6305) >>> _zz_1986);
  assign _zz_6305 = _zz_6306;
  assign _zz_6306 = ($signed(_zz_153) - $signed(_zz_1983));
  assign _zz_6307 = _zz_6308;
  assign _zz_6308 = ($signed(_zz_6309) >>> _zz_1986);
  assign _zz_6309 = _zz_6310;
  assign _zz_6310 = ($signed(_zz_154) - $signed(_zz_1984));
  assign _zz_6311 = _zz_6312;
  assign _zz_6312 = ($signed(_zz_6313) >>> _zz_1987);
  assign _zz_6313 = _zz_6314;
  assign _zz_6314 = ($signed(_zz_153) + $signed(_zz_1983));
  assign _zz_6315 = _zz_6316;
  assign _zz_6316 = ($signed(_zz_6317) >>> _zz_1987);
  assign _zz_6317 = _zz_6318;
  assign _zz_6318 = ($signed(_zz_154) + $signed(_zz_1984));
  assign _zz_6319 = ($signed(twiddle_factor_table_0_real) + $signed(twiddle_factor_table_0_imag));
  assign _zz_6320 = fixTo_117_dout;
  assign _zz_6321 = ($signed(_zz_160) - $signed(_zz_159));
  assign _zz_6322 = ($signed(_zz_159) + $signed(_zz_160));
  assign _zz_6323 = _zz_6324[15 : 0];
  assign _zz_6324 = fixTo_119_dout;
  assign _zz_6325 = _zz_6326[15 : 0];
  assign _zz_6326 = fixTo_118_dout;
  assign _zz_6327 = _zz_6328;
  assign _zz_6328 = ($signed(_zz_6329) >>> _zz_1991);
  assign _zz_6329 = _zz_6330;
  assign _zz_6330 = ($signed(_zz_157) - $signed(_zz_1988));
  assign _zz_6331 = _zz_6332;
  assign _zz_6332 = ($signed(_zz_6333) >>> _zz_1991);
  assign _zz_6333 = _zz_6334;
  assign _zz_6334 = ($signed(_zz_158) - $signed(_zz_1989));
  assign _zz_6335 = _zz_6336;
  assign _zz_6336 = ($signed(_zz_6337) >>> _zz_1992);
  assign _zz_6337 = _zz_6338;
  assign _zz_6338 = ($signed(_zz_157) + $signed(_zz_1988));
  assign _zz_6339 = _zz_6340;
  assign _zz_6340 = ($signed(_zz_6341) >>> _zz_1992);
  assign _zz_6341 = _zz_6342;
  assign _zz_6342 = ($signed(_zz_158) + $signed(_zz_1989));
  assign _zz_6343 = ($signed(twiddle_factor_table_0_real) + $signed(twiddle_factor_table_0_imag));
  assign _zz_6344 = fixTo_120_dout;
  assign _zz_6345 = ($signed(_zz_164) - $signed(_zz_163));
  assign _zz_6346 = ($signed(_zz_163) + $signed(_zz_164));
  assign _zz_6347 = _zz_6348[15 : 0];
  assign _zz_6348 = fixTo_122_dout;
  assign _zz_6349 = _zz_6350[15 : 0];
  assign _zz_6350 = fixTo_121_dout;
  assign _zz_6351 = _zz_6352;
  assign _zz_6352 = ($signed(_zz_6353) >>> _zz_1996);
  assign _zz_6353 = _zz_6354;
  assign _zz_6354 = ($signed(_zz_161) - $signed(_zz_1993));
  assign _zz_6355 = _zz_6356;
  assign _zz_6356 = ($signed(_zz_6357) >>> _zz_1996);
  assign _zz_6357 = _zz_6358;
  assign _zz_6358 = ($signed(_zz_162) - $signed(_zz_1994));
  assign _zz_6359 = _zz_6360;
  assign _zz_6360 = ($signed(_zz_6361) >>> _zz_1997);
  assign _zz_6361 = _zz_6362;
  assign _zz_6362 = ($signed(_zz_161) + $signed(_zz_1993));
  assign _zz_6363 = _zz_6364;
  assign _zz_6364 = ($signed(_zz_6365) >>> _zz_1997);
  assign _zz_6365 = _zz_6366;
  assign _zz_6366 = ($signed(_zz_162) + $signed(_zz_1994));
  assign _zz_6367 = ($signed(twiddle_factor_table_0_real) + $signed(twiddle_factor_table_0_imag));
  assign _zz_6368 = fixTo_123_dout;
  assign _zz_6369 = ($signed(_zz_168) - $signed(_zz_167));
  assign _zz_6370 = ($signed(_zz_167) + $signed(_zz_168));
  assign _zz_6371 = _zz_6372[15 : 0];
  assign _zz_6372 = fixTo_125_dout;
  assign _zz_6373 = _zz_6374[15 : 0];
  assign _zz_6374 = fixTo_124_dout;
  assign _zz_6375 = _zz_6376;
  assign _zz_6376 = ($signed(_zz_6377) >>> _zz_2001);
  assign _zz_6377 = _zz_6378;
  assign _zz_6378 = ($signed(_zz_165) - $signed(_zz_1998));
  assign _zz_6379 = _zz_6380;
  assign _zz_6380 = ($signed(_zz_6381) >>> _zz_2001);
  assign _zz_6381 = _zz_6382;
  assign _zz_6382 = ($signed(_zz_166) - $signed(_zz_1999));
  assign _zz_6383 = _zz_6384;
  assign _zz_6384 = ($signed(_zz_6385) >>> _zz_2002);
  assign _zz_6385 = _zz_6386;
  assign _zz_6386 = ($signed(_zz_165) + $signed(_zz_1998));
  assign _zz_6387 = _zz_6388;
  assign _zz_6388 = ($signed(_zz_6389) >>> _zz_2002);
  assign _zz_6389 = _zz_6390;
  assign _zz_6390 = ($signed(_zz_166) + $signed(_zz_1999));
  assign _zz_6391 = ($signed(twiddle_factor_table_0_real) + $signed(twiddle_factor_table_0_imag));
  assign _zz_6392 = fixTo_126_dout;
  assign _zz_6393 = ($signed(_zz_172) - $signed(_zz_171));
  assign _zz_6394 = ($signed(_zz_171) + $signed(_zz_172));
  assign _zz_6395 = _zz_6396[15 : 0];
  assign _zz_6396 = fixTo_128_dout;
  assign _zz_6397 = _zz_6398[15 : 0];
  assign _zz_6398 = fixTo_127_dout;
  assign _zz_6399 = _zz_6400;
  assign _zz_6400 = ($signed(_zz_6401) >>> _zz_2006);
  assign _zz_6401 = _zz_6402;
  assign _zz_6402 = ($signed(_zz_169) - $signed(_zz_2003));
  assign _zz_6403 = _zz_6404;
  assign _zz_6404 = ($signed(_zz_6405) >>> _zz_2006);
  assign _zz_6405 = _zz_6406;
  assign _zz_6406 = ($signed(_zz_170) - $signed(_zz_2004));
  assign _zz_6407 = _zz_6408;
  assign _zz_6408 = ($signed(_zz_6409) >>> _zz_2007);
  assign _zz_6409 = _zz_6410;
  assign _zz_6410 = ($signed(_zz_169) + $signed(_zz_2003));
  assign _zz_6411 = _zz_6412;
  assign _zz_6412 = ($signed(_zz_6413) >>> _zz_2007);
  assign _zz_6413 = _zz_6414;
  assign _zz_6414 = ($signed(_zz_170) + $signed(_zz_2004));
  assign _zz_6415 = ($signed(twiddle_factor_table_0_real) + $signed(twiddle_factor_table_0_imag));
  assign _zz_6416 = fixTo_129_dout;
  assign _zz_6417 = ($signed(_zz_176) - $signed(_zz_175));
  assign _zz_6418 = ($signed(_zz_175) + $signed(_zz_176));
  assign _zz_6419 = _zz_6420[15 : 0];
  assign _zz_6420 = fixTo_131_dout;
  assign _zz_6421 = _zz_6422[15 : 0];
  assign _zz_6422 = fixTo_130_dout;
  assign _zz_6423 = _zz_6424;
  assign _zz_6424 = ($signed(_zz_6425) >>> _zz_2011);
  assign _zz_6425 = _zz_6426;
  assign _zz_6426 = ($signed(_zz_173) - $signed(_zz_2008));
  assign _zz_6427 = _zz_6428;
  assign _zz_6428 = ($signed(_zz_6429) >>> _zz_2011);
  assign _zz_6429 = _zz_6430;
  assign _zz_6430 = ($signed(_zz_174) - $signed(_zz_2009));
  assign _zz_6431 = _zz_6432;
  assign _zz_6432 = ($signed(_zz_6433) >>> _zz_2012);
  assign _zz_6433 = _zz_6434;
  assign _zz_6434 = ($signed(_zz_173) + $signed(_zz_2008));
  assign _zz_6435 = _zz_6436;
  assign _zz_6436 = ($signed(_zz_6437) >>> _zz_2012);
  assign _zz_6437 = _zz_6438;
  assign _zz_6438 = ($signed(_zz_174) + $signed(_zz_2009));
  assign _zz_6439 = ($signed(twiddle_factor_table_0_real) + $signed(twiddle_factor_table_0_imag));
  assign _zz_6440 = fixTo_132_dout;
  assign _zz_6441 = ($signed(_zz_180) - $signed(_zz_179));
  assign _zz_6442 = ($signed(_zz_179) + $signed(_zz_180));
  assign _zz_6443 = _zz_6444[15 : 0];
  assign _zz_6444 = fixTo_134_dout;
  assign _zz_6445 = _zz_6446[15 : 0];
  assign _zz_6446 = fixTo_133_dout;
  assign _zz_6447 = _zz_6448;
  assign _zz_6448 = ($signed(_zz_6449) >>> _zz_2016);
  assign _zz_6449 = _zz_6450;
  assign _zz_6450 = ($signed(_zz_177) - $signed(_zz_2013));
  assign _zz_6451 = _zz_6452;
  assign _zz_6452 = ($signed(_zz_6453) >>> _zz_2016);
  assign _zz_6453 = _zz_6454;
  assign _zz_6454 = ($signed(_zz_178) - $signed(_zz_2014));
  assign _zz_6455 = _zz_6456;
  assign _zz_6456 = ($signed(_zz_6457) >>> _zz_2017);
  assign _zz_6457 = _zz_6458;
  assign _zz_6458 = ($signed(_zz_177) + $signed(_zz_2013));
  assign _zz_6459 = _zz_6460;
  assign _zz_6460 = ($signed(_zz_6461) >>> _zz_2017);
  assign _zz_6461 = _zz_6462;
  assign _zz_6462 = ($signed(_zz_178) + $signed(_zz_2014));
  assign _zz_6463 = ($signed(twiddle_factor_table_0_real) + $signed(twiddle_factor_table_0_imag));
  assign _zz_6464 = fixTo_135_dout;
  assign _zz_6465 = ($signed(_zz_184) - $signed(_zz_183));
  assign _zz_6466 = ($signed(_zz_183) + $signed(_zz_184));
  assign _zz_6467 = _zz_6468[15 : 0];
  assign _zz_6468 = fixTo_137_dout;
  assign _zz_6469 = _zz_6470[15 : 0];
  assign _zz_6470 = fixTo_136_dout;
  assign _zz_6471 = _zz_6472;
  assign _zz_6472 = ($signed(_zz_6473) >>> _zz_2021);
  assign _zz_6473 = _zz_6474;
  assign _zz_6474 = ($signed(_zz_181) - $signed(_zz_2018));
  assign _zz_6475 = _zz_6476;
  assign _zz_6476 = ($signed(_zz_6477) >>> _zz_2021);
  assign _zz_6477 = _zz_6478;
  assign _zz_6478 = ($signed(_zz_182) - $signed(_zz_2019));
  assign _zz_6479 = _zz_6480;
  assign _zz_6480 = ($signed(_zz_6481) >>> _zz_2022);
  assign _zz_6481 = _zz_6482;
  assign _zz_6482 = ($signed(_zz_181) + $signed(_zz_2018));
  assign _zz_6483 = _zz_6484;
  assign _zz_6484 = ($signed(_zz_6485) >>> _zz_2022);
  assign _zz_6485 = _zz_6486;
  assign _zz_6486 = ($signed(_zz_182) + $signed(_zz_2019));
  assign _zz_6487 = ($signed(twiddle_factor_table_0_real) + $signed(twiddle_factor_table_0_imag));
  assign _zz_6488 = fixTo_138_dout;
  assign _zz_6489 = ($signed(_zz_188) - $signed(_zz_187));
  assign _zz_6490 = ($signed(_zz_187) + $signed(_zz_188));
  assign _zz_6491 = _zz_6492[15 : 0];
  assign _zz_6492 = fixTo_140_dout;
  assign _zz_6493 = _zz_6494[15 : 0];
  assign _zz_6494 = fixTo_139_dout;
  assign _zz_6495 = _zz_6496;
  assign _zz_6496 = ($signed(_zz_6497) >>> _zz_2026);
  assign _zz_6497 = _zz_6498;
  assign _zz_6498 = ($signed(_zz_185) - $signed(_zz_2023));
  assign _zz_6499 = _zz_6500;
  assign _zz_6500 = ($signed(_zz_6501) >>> _zz_2026);
  assign _zz_6501 = _zz_6502;
  assign _zz_6502 = ($signed(_zz_186) - $signed(_zz_2024));
  assign _zz_6503 = _zz_6504;
  assign _zz_6504 = ($signed(_zz_6505) >>> _zz_2027);
  assign _zz_6505 = _zz_6506;
  assign _zz_6506 = ($signed(_zz_185) + $signed(_zz_2023));
  assign _zz_6507 = _zz_6508;
  assign _zz_6508 = ($signed(_zz_6509) >>> _zz_2027);
  assign _zz_6509 = _zz_6510;
  assign _zz_6510 = ($signed(_zz_186) + $signed(_zz_2024));
  assign _zz_6511 = ($signed(twiddle_factor_table_0_real) + $signed(twiddle_factor_table_0_imag));
  assign _zz_6512 = fixTo_141_dout;
  assign _zz_6513 = ($signed(_zz_192) - $signed(_zz_191));
  assign _zz_6514 = ($signed(_zz_191) + $signed(_zz_192));
  assign _zz_6515 = _zz_6516[15 : 0];
  assign _zz_6516 = fixTo_143_dout;
  assign _zz_6517 = _zz_6518[15 : 0];
  assign _zz_6518 = fixTo_142_dout;
  assign _zz_6519 = _zz_6520;
  assign _zz_6520 = ($signed(_zz_6521) >>> _zz_2031);
  assign _zz_6521 = _zz_6522;
  assign _zz_6522 = ($signed(_zz_189) - $signed(_zz_2028));
  assign _zz_6523 = _zz_6524;
  assign _zz_6524 = ($signed(_zz_6525) >>> _zz_2031);
  assign _zz_6525 = _zz_6526;
  assign _zz_6526 = ($signed(_zz_190) - $signed(_zz_2029));
  assign _zz_6527 = _zz_6528;
  assign _zz_6528 = ($signed(_zz_6529) >>> _zz_2032);
  assign _zz_6529 = _zz_6530;
  assign _zz_6530 = ($signed(_zz_189) + $signed(_zz_2028));
  assign _zz_6531 = _zz_6532;
  assign _zz_6532 = ($signed(_zz_6533) >>> _zz_2032);
  assign _zz_6533 = _zz_6534;
  assign _zz_6534 = ($signed(_zz_190) + $signed(_zz_2029));
  assign _zz_6535 = ($signed(twiddle_factor_table_0_real) + $signed(twiddle_factor_table_0_imag));
  assign _zz_6536 = fixTo_144_dout;
  assign _zz_6537 = ($signed(_zz_196) - $signed(_zz_195));
  assign _zz_6538 = ($signed(_zz_195) + $signed(_zz_196));
  assign _zz_6539 = _zz_6540[15 : 0];
  assign _zz_6540 = fixTo_146_dout;
  assign _zz_6541 = _zz_6542[15 : 0];
  assign _zz_6542 = fixTo_145_dout;
  assign _zz_6543 = _zz_6544;
  assign _zz_6544 = ($signed(_zz_6545) >>> _zz_2036);
  assign _zz_6545 = _zz_6546;
  assign _zz_6546 = ($signed(_zz_193) - $signed(_zz_2033));
  assign _zz_6547 = _zz_6548;
  assign _zz_6548 = ($signed(_zz_6549) >>> _zz_2036);
  assign _zz_6549 = _zz_6550;
  assign _zz_6550 = ($signed(_zz_194) - $signed(_zz_2034));
  assign _zz_6551 = _zz_6552;
  assign _zz_6552 = ($signed(_zz_6553) >>> _zz_2037);
  assign _zz_6553 = _zz_6554;
  assign _zz_6554 = ($signed(_zz_193) + $signed(_zz_2033));
  assign _zz_6555 = _zz_6556;
  assign _zz_6556 = ($signed(_zz_6557) >>> _zz_2037);
  assign _zz_6557 = _zz_6558;
  assign _zz_6558 = ($signed(_zz_194) + $signed(_zz_2034));
  assign _zz_6559 = ($signed(twiddle_factor_table_0_real) + $signed(twiddle_factor_table_0_imag));
  assign _zz_6560 = fixTo_147_dout;
  assign _zz_6561 = ($signed(_zz_200) - $signed(_zz_199));
  assign _zz_6562 = ($signed(_zz_199) + $signed(_zz_200));
  assign _zz_6563 = _zz_6564[15 : 0];
  assign _zz_6564 = fixTo_149_dout;
  assign _zz_6565 = _zz_6566[15 : 0];
  assign _zz_6566 = fixTo_148_dout;
  assign _zz_6567 = _zz_6568;
  assign _zz_6568 = ($signed(_zz_6569) >>> _zz_2041);
  assign _zz_6569 = _zz_6570;
  assign _zz_6570 = ($signed(_zz_197) - $signed(_zz_2038));
  assign _zz_6571 = _zz_6572;
  assign _zz_6572 = ($signed(_zz_6573) >>> _zz_2041);
  assign _zz_6573 = _zz_6574;
  assign _zz_6574 = ($signed(_zz_198) - $signed(_zz_2039));
  assign _zz_6575 = _zz_6576;
  assign _zz_6576 = ($signed(_zz_6577) >>> _zz_2042);
  assign _zz_6577 = _zz_6578;
  assign _zz_6578 = ($signed(_zz_197) + $signed(_zz_2038));
  assign _zz_6579 = _zz_6580;
  assign _zz_6580 = ($signed(_zz_6581) >>> _zz_2042);
  assign _zz_6581 = _zz_6582;
  assign _zz_6582 = ($signed(_zz_198) + $signed(_zz_2039));
  assign _zz_6583 = ($signed(twiddle_factor_table_0_real) + $signed(twiddle_factor_table_0_imag));
  assign _zz_6584 = fixTo_150_dout;
  assign _zz_6585 = ($signed(_zz_204) - $signed(_zz_203));
  assign _zz_6586 = ($signed(_zz_203) + $signed(_zz_204));
  assign _zz_6587 = _zz_6588[15 : 0];
  assign _zz_6588 = fixTo_152_dout;
  assign _zz_6589 = _zz_6590[15 : 0];
  assign _zz_6590 = fixTo_151_dout;
  assign _zz_6591 = _zz_6592;
  assign _zz_6592 = ($signed(_zz_6593) >>> _zz_2046);
  assign _zz_6593 = _zz_6594;
  assign _zz_6594 = ($signed(_zz_201) - $signed(_zz_2043));
  assign _zz_6595 = _zz_6596;
  assign _zz_6596 = ($signed(_zz_6597) >>> _zz_2046);
  assign _zz_6597 = _zz_6598;
  assign _zz_6598 = ($signed(_zz_202) - $signed(_zz_2044));
  assign _zz_6599 = _zz_6600;
  assign _zz_6600 = ($signed(_zz_6601) >>> _zz_2047);
  assign _zz_6601 = _zz_6602;
  assign _zz_6602 = ($signed(_zz_201) + $signed(_zz_2043));
  assign _zz_6603 = _zz_6604;
  assign _zz_6604 = ($signed(_zz_6605) >>> _zz_2047);
  assign _zz_6605 = _zz_6606;
  assign _zz_6606 = ($signed(_zz_202) + $signed(_zz_2044));
  assign _zz_6607 = ($signed(twiddle_factor_table_0_real) + $signed(twiddle_factor_table_0_imag));
  assign _zz_6608 = fixTo_153_dout;
  assign _zz_6609 = ($signed(_zz_208) - $signed(_zz_207));
  assign _zz_6610 = ($signed(_zz_207) + $signed(_zz_208));
  assign _zz_6611 = _zz_6612[15 : 0];
  assign _zz_6612 = fixTo_155_dout;
  assign _zz_6613 = _zz_6614[15 : 0];
  assign _zz_6614 = fixTo_154_dout;
  assign _zz_6615 = _zz_6616;
  assign _zz_6616 = ($signed(_zz_6617) >>> _zz_2051);
  assign _zz_6617 = _zz_6618;
  assign _zz_6618 = ($signed(_zz_205) - $signed(_zz_2048));
  assign _zz_6619 = _zz_6620;
  assign _zz_6620 = ($signed(_zz_6621) >>> _zz_2051);
  assign _zz_6621 = _zz_6622;
  assign _zz_6622 = ($signed(_zz_206) - $signed(_zz_2049));
  assign _zz_6623 = _zz_6624;
  assign _zz_6624 = ($signed(_zz_6625) >>> _zz_2052);
  assign _zz_6625 = _zz_6626;
  assign _zz_6626 = ($signed(_zz_205) + $signed(_zz_2048));
  assign _zz_6627 = _zz_6628;
  assign _zz_6628 = ($signed(_zz_6629) >>> _zz_2052);
  assign _zz_6629 = _zz_6630;
  assign _zz_6630 = ($signed(_zz_206) + $signed(_zz_2049));
  assign _zz_6631 = ($signed(twiddle_factor_table_0_real) + $signed(twiddle_factor_table_0_imag));
  assign _zz_6632 = fixTo_156_dout;
  assign _zz_6633 = ($signed(_zz_212) - $signed(_zz_211));
  assign _zz_6634 = ($signed(_zz_211) + $signed(_zz_212));
  assign _zz_6635 = _zz_6636[15 : 0];
  assign _zz_6636 = fixTo_158_dout;
  assign _zz_6637 = _zz_6638[15 : 0];
  assign _zz_6638 = fixTo_157_dout;
  assign _zz_6639 = _zz_6640;
  assign _zz_6640 = ($signed(_zz_6641) >>> _zz_2056);
  assign _zz_6641 = _zz_6642;
  assign _zz_6642 = ($signed(_zz_209) - $signed(_zz_2053));
  assign _zz_6643 = _zz_6644;
  assign _zz_6644 = ($signed(_zz_6645) >>> _zz_2056);
  assign _zz_6645 = _zz_6646;
  assign _zz_6646 = ($signed(_zz_210) - $signed(_zz_2054));
  assign _zz_6647 = _zz_6648;
  assign _zz_6648 = ($signed(_zz_6649) >>> _zz_2057);
  assign _zz_6649 = _zz_6650;
  assign _zz_6650 = ($signed(_zz_209) + $signed(_zz_2053));
  assign _zz_6651 = _zz_6652;
  assign _zz_6652 = ($signed(_zz_6653) >>> _zz_2057);
  assign _zz_6653 = _zz_6654;
  assign _zz_6654 = ($signed(_zz_210) + $signed(_zz_2054));
  assign _zz_6655 = ($signed(twiddle_factor_table_0_real) + $signed(twiddle_factor_table_0_imag));
  assign _zz_6656 = fixTo_159_dout;
  assign _zz_6657 = ($signed(_zz_216) - $signed(_zz_215));
  assign _zz_6658 = ($signed(_zz_215) + $signed(_zz_216));
  assign _zz_6659 = _zz_6660[15 : 0];
  assign _zz_6660 = fixTo_161_dout;
  assign _zz_6661 = _zz_6662[15 : 0];
  assign _zz_6662 = fixTo_160_dout;
  assign _zz_6663 = _zz_6664;
  assign _zz_6664 = ($signed(_zz_6665) >>> _zz_2061);
  assign _zz_6665 = _zz_6666;
  assign _zz_6666 = ($signed(_zz_213) - $signed(_zz_2058));
  assign _zz_6667 = _zz_6668;
  assign _zz_6668 = ($signed(_zz_6669) >>> _zz_2061);
  assign _zz_6669 = _zz_6670;
  assign _zz_6670 = ($signed(_zz_214) - $signed(_zz_2059));
  assign _zz_6671 = _zz_6672;
  assign _zz_6672 = ($signed(_zz_6673) >>> _zz_2062);
  assign _zz_6673 = _zz_6674;
  assign _zz_6674 = ($signed(_zz_213) + $signed(_zz_2058));
  assign _zz_6675 = _zz_6676;
  assign _zz_6676 = ($signed(_zz_6677) >>> _zz_2062);
  assign _zz_6677 = _zz_6678;
  assign _zz_6678 = ($signed(_zz_214) + $signed(_zz_2059));
  assign _zz_6679 = ($signed(twiddle_factor_table_0_real) + $signed(twiddle_factor_table_0_imag));
  assign _zz_6680 = fixTo_162_dout;
  assign _zz_6681 = ($signed(_zz_220) - $signed(_zz_219));
  assign _zz_6682 = ($signed(_zz_219) + $signed(_zz_220));
  assign _zz_6683 = _zz_6684[15 : 0];
  assign _zz_6684 = fixTo_164_dout;
  assign _zz_6685 = _zz_6686[15 : 0];
  assign _zz_6686 = fixTo_163_dout;
  assign _zz_6687 = _zz_6688;
  assign _zz_6688 = ($signed(_zz_6689) >>> _zz_2066);
  assign _zz_6689 = _zz_6690;
  assign _zz_6690 = ($signed(_zz_217) - $signed(_zz_2063));
  assign _zz_6691 = _zz_6692;
  assign _zz_6692 = ($signed(_zz_6693) >>> _zz_2066);
  assign _zz_6693 = _zz_6694;
  assign _zz_6694 = ($signed(_zz_218) - $signed(_zz_2064));
  assign _zz_6695 = _zz_6696;
  assign _zz_6696 = ($signed(_zz_6697) >>> _zz_2067);
  assign _zz_6697 = _zz_6698;
  assign _zz_6698 = ($signed(_zz_217) + $signed(_zz_2063));
  assign _zz_6699 = _zz_6700;
  assign _zz_6700 = ($signed(_zz_6701) >>> _zz_2067);
  assign _zz_6701 = _zz_6702;
  assign _zz_6702 = ($signed(_zz_218) + $signed(_zz_2064));
  assign _zz_6703 = ($signed(twiddle_factor_table_0_real) + $signed(twiddle_factor_table_0_imag));
  assign _zz_6704 = fixTo_165_dout;
  assign _zz_6705 = ($signed(_zz_224) - $signed(_zz_223));
  assign _zz_6706 = ($signed(_zz_223) + $signed(_zz_224));
  assign _zz_6707 = _zz_6708[15 : 0];
  assign _zz_6708 = fixTo_167_dout;
  assign _zz_6709 = _zz_6710[15 : 0];
  assign _zz_6710 = fixTo_166_dout;
  assign _zz_6711 = _zz_6712;
  assign _zz_6712 = ($signed(_zz_6713) >>> _zz_2071);
  assign _zz_6713 = _zz_6714;
  assign _zz_6714 = ($signed(_zz_221) - $signed(_zz_2068));
  assign _zz_6715 = _zz_6716;
  assign _zz_6716 = ($signed(_zz_6717) >>> _zz_2071);
  assign _zz_6717 = _zz_6718;
  assign _zz_6718 = ($signed(_zz_222) - $signed(_zz_2069));
  assign _zz_6719 = _zz_6720;
  assign _zz_6720 = ($signed(_zz_6721) >>> _zz_2072);
  assign _zz_6721 = _zz_6722;
  assign _zz_6722 = ($signed(_zz_221) + $signed(_zz_2068));
  assign _zz_6723 = _zz_6724;
  assign _zz_6724 = ($signed(_zz_6725) >>> _zz_2072);
  assign _zz_6725 = _zz_6726;
  assign _zz_6726 = ($signed(_zz_222) + $signed(_zz_2069));
  assign _zz_6727 = ($signed(twiddle_factor_table_0_real) + $signed(twiddle_factor_table_0_imag));
  assign _zz_6728 = fixTo_168_dout;
  assign _zz_6729 = ($signed(_zz_228) - $signed(_zz_227));
  assign _zz_6730 = ($signed(_zz_227) + $signed(_zz_228));
  assign _zz_6731 = _zz_6732[15 : 0];
  assign _zz_6732 = fixTo_170_dout;
  assign _zz_6733 = _zz_6734[15 : 0];
  assign _zz_6734 = fixTo_169_dout;
  assign _zz_6735 = _zz_6736;
  assign _zz_6736 = ($signed(_zz_6737) >>> _zz_2076);
  assign _zz_6737 = _zz_6738;
  assign _zz_6738 = ($signed(_zz_225) - $signed(_zz_2073));
  assign _zz_6739 = _zz_6740;
  assign _zz_6740 = ($signed(_zz_6741) >>> _zz_2076);
  assign _zz_6741 = _zz_6742;
  assign _zz_6742 = ($signed(_zz_226) - $signed(_zz_2074));
  assign _zz_6743 = _zz_6744;
  assign _zz_6744 = ($signed(_zz_6745) >>> _zz_2077);
  assign _zz_6745 = _zz_6746;
  assign _zz_6746 = ($signed(_zz_225) + $signed(_zz_2073));
  assign _zz_6747 = _zz_6748;
  assign _zz_6748 = ($signed(_zz_6749) >>> _zz_2077);
  assign _zz_6749 = _zz_6750;
  assign _zz_6750 = ($signed(_zz_226) + $signed(_zz_2074));
  assign _zz_6751 = ($signed(twiddle_factor_table_0_real) + $signed(twiddle_factor_table_0_imag));
  assign _zz_6752 = fixTo_171_dout;
  assign _zz_6753 = ($signed(_zz_232) - $signed(_zz_231));
  assign _zz_6754 = ($signed(_zz_231) + $signed(_zz_232));
  assign _zz_6755 = _zz_6756[15 : 0];
  assign _zz_6756 = fixTo_173_dout;
  assign _zz_6757 = _zz_6758[15 : 0];
  assign _zz_6758 = fixTo_172_dout;
  assign _zz_6759 = _zz_6760;
  assign _zz_6760 = ($signed(_zz_6761) >>> _zz_2081);
  assign _zz_6761 = _zz_6762;
  assign _zz_6762 = ($signed(_zz_229) - $signed(_zz_2078));
  assign _zz_6763 = _zz_6764;
  assign _zz_6764 = ($signed(_zz_6765) >>> _zz_2081);
  assign _zz_6765 = _zz_6766;
  assign _zz_6766 = ($signed(_zz_230) - $signed(_zz_2079));
  assign _zz_6767 = _zz_6768;
  assign _zz_6768 = ($signed(_zz_6769) >>> _zz_2082);
  assign _zz_6769 = _zz_6770;
  assign _zz_6770 = ($signed(_zz_229) + $signed(_zz_2078));
  assign _zz_6771 = _zz_6772;
  assign _zz_6772 = ($signed(_zz_6773) >>> _zz_2082);
  assign _zz_6773 = _zz_6774;
  assign _zz_6774 = ($signed(_zz_230) + $signed(_zz_2079));
  assign _zz_6775 = ($signed(twiddle_factor_table_0_real) + $signed(twiddle_factor_table_0_imag));
  assign _zz_6776 = fixTo_174_dout;
  assign _zz_6777 = ($signed(_zz_236) - $signed(_zz_235));
  assign _zz_6778 = ($signed(_zz_235) + $signed(_zz_236));
  assign _zz_6779 = _zz_6780[15 : 0];
  assign _zz_6780 = fixTo_176_dout;
  assign _zz_6781 = _zz_6782[15 : 0];
  assign _zz_6782 = fixTo_175_dout;
  assign _zz_6783 = _zz_6784;
  assign _zz_6784 = ($signed(_zz_6785) >>> _zz_2086);
  assign _zz_6785 = _zz_6786;
  assign _zz_6786 = ($signed(_zz_233) - $signed(_zz_2083));
  assign _zz_6787 = _zz_6788;
  assign _zz_6788 = ($signed(_zz_6789) >>> _zz_2086);
  assign _zz_6789 = _zz_6790;
  assign _zz_6790 = ($signed(_zz_234) - $signed(_zz_2084));
  assign _zz_6791 = _zz_6792;
  assign _zz_6792 = ($signed(_zz_6793) >>> _zz_2087);
  assign _zz_6793 = _zz_6794;
  assign _zz_6794 = ($signed(_zz_233) + $signed(_zz_2083));
  assign _zz_6795 = _zz_6796;
  assign _zz_6796 = ($signed(_zz_6797) >>> _zz_2087);
  assign _zz_6797 = _zz_6798;
  assign _zz_6798 = ($signed(_zz_234) + $signed(_zz_2084));
  assign _zz_6799 = ($signed(twiddle_factor_table_0_real) + $signed(twiddle_factor_table_0_imag));
  assign _zz_6800 = fixTo_177_dout;
  assign _zz_6801 = ($signed(_zz_240) - $signed(_zz_239));
  assign _zz_6802 = ($signed(_zz_239) + $signed(_zz_240));
  assign _zz_6803 = _zz_6804[15 : 0];
  assign _zz_6804 = fixTo_179_dout;
  assign _zz_6805 = _zz_6806[15 : 0];
  assign _zz_6806 = fixTo_178_dout;
  assign _zz_6807 = _zz_6808;
  assign _zz_6808 = ($signed(_zz_6809) >>> _zz_2091);
  assign _zz_6809 = _zz_6810;
  assign _zz_6810 = ($signed(_zz_237) - $signed(_zz_2088));
  assign _zz_6811 = _zz_6812;
  assign _zz_6812 = ($signed(_zz_6813) >>> _zz_2091);
  assign _zz_6813 = _zz_6814;
  assign _zz_6814 = ($signed(_zz_238) - $signed(_zz_2089));
  assign _zz_6815 = _zz_6816;
  assign _zz_6816 = ($signed(_zz_6817) >>> _zz_2092);
  assign _zz_6817 = _zz_6818;
  assign _zz_6818 = ($signed(_zz_237) + $signed(_zz_2088));
  assign _zz_6819 = _zz_6820;
  assign _zz_6820 = ($signed(_zz_6821) >>> _zz_2092);
  assign _zz_6821 = _zz_6822;
  assign _zz_6822 = ($signed(_zz_238) + $signed(_zz_2089));
  assign _zz_6823 = ($signed(twiddle_factor_table_0_real) + $signed(twiddle_factor_table_0_imag));
  assign _zz_6824 = fixTo_180_dout;
  assign _zz_6825 = ($signed(_zz_244) - $signed(_zz_243));
  assign _zz_6826 = ($signed(_zz_243) + $signed(_zz_244));
  assign _zz_6827 = _zz_6828[15 : 0];
  assign _zz_6828 = fixTo_182_dout;
  assign _zz_6829 = _zz_6830[15 : 0];
  assign _zz_6830 = fixTo_181_dout;
  assign _zz_6831 = _zz_6832;
  assign _zz_6832 = ($signed(_zz_6833) >>> _zz_2096);
  assign _zz_6833 = _zz_6834;
  assign _zz_6834 = ($signed(_zz_241) - $signed(_zz_2093));
  assign _zz_6835 = _zz_6836;
  assign _zz_6836 = ($signed(_zz_6837) >>> _zz_2096);
  assign _zz_6837 = _zz_6838;
  assign _zz_6838 = ($signed(_zz_242) - $signed(_zz_2094));
  assign _zz_6839 = _zz_6840;
  assign _zz_6840 = ($signed(_zz_6841) >>> _zz_2097);
  assign _zz_6841 = _zz_6842;
  assign _zz_6842 = ($signed(_zz_241) + $signed(_zz_2093));
  assign _zz_6843 = _zz_6844;
  assign _zz_6844 = ($signed(_zz_6845) >>> _zz_2097);
  assign _zz_6845 = _zz_6846;
  assign _zz_6846 = ($signed(_zz_242) + $signed(_zz_2094));
  assign _zz_6847 = ($signed(twiddle_factor_table_0_real) + $signed(twiddle_factor_table_0_imag));
  assign _zz_6848 = fixTo_183_dout;
  assign _zz_6849 = ($signed(_zz_248) - $signed(_zz_247));
  assign _zz_6850 = ($signed(_zz_247) + $signed(_zz_248));
  assign _zz_6851 = _zz_6852[15 : 0];
  assign _zz_6852 = fixTo_185_dout;
  assign _zz_6853 = _zz_6854[15 : 0];
  assign _zz_6854 = fixTo_184_dout;
  assign _zz_6855 = _zz_6856;
  assign _zz_6856 = ($signed(_zz_6857) >>> _zz_2101);
  assign _zz_6857 = _zz_6858;
  assign _zz_6858 = ($signed(_zz_245) - $signed(_zz_2098));
  assign _zz_6859 = _zz_6860;
  assign _zz_6860 = ($signed(_zz_6861) >>> _zz_2101);
  assign _zz_6861 = _zz_6862;
  assign _zz_6862 = ($signed(_zz_246) - $signed(_zz_2099));
  assign _zz_6863 = _zz_6864;
  assign _zz_6864 = ($signed(_zz_6865) >>> _zz_2102);
  assign _zz_6865 = _zz_6866;
  assign _zz_6866 = ($signed(_zz_245) + $signed(_zz_2098));
  assign _zz_6867 = _zz_6868;
  assign _zz_6868 = ($signed(_zz_6869) >>> _zz_2102);
  assign _zz_6869 = _zz_6870;
  assign _zz_6870 = ($signed(_zz_246) + $signed(_zz_2099));
  assign _zz_6871 = ($signed(twiddle_factor_table_0_real) + $signed(twiddle_factor_table_0_imag));
  assign _zz_6872 = fixTo_186_dout;
  assign _zz_6873 = ($signed(_zz_252) - $signed(_zz_251));
  assign _zz_6874 = ($signed(_zz_251) + $signed(_zz_252));
  assign _zz_6875 = _zz_6876[15 : 0];
  assign _zz_6876 = fixTo_188_dout;
  assign _zz_6877 = _zz_6878[15 : 0];
  assign _zz_6878 = fixTo_187_dout;
  assign _zz_6879 = _zz_6880;
  assign _zz_6880 = ($signed(_zz_6881) >>> _zz_2106);
  assign _zz_6881 = _zz_6882;
  assign _zz_6882 = ($signed(_zz_249) - $signed(_zz_2103));
  assign _zz_6883 = _zz_6884;
  assign _zz_6884 = ($signed(_zz_6885) >>> _zz_2106);
  assign _zz_6885 = _zz_6886;
  assign _zz_6886 = ($signed(_zz_250) - $signed(_zz_2104));
  assign _zz_6887 = _zz_6888;
  assign _zz_6888 = ($signed(_zz_6889) >>> _zz_2107);
  assign _zz_6889 = _zz_6890;
  assign _zz_6890 = ($signed(_zz_249) + $signed(_zz_2103));
  assign _zz_6891 = _zz_6892;
  assign _zz_6892 = ($signed(_zz_6893) >>> _zz_2107);
  assign _zz_6893 = _zz_6894;
  assign _zz_6894 = ($signed(_zz_250) + $signed(_zz_2104));
  assign _zz_6895 = ($signed(twiddle_factor_table_0_real) + $signed(twiddle_factor_table_0_imag));
  assign _zz_6896 = fixTo_189_dout;
  assign _zz_6897 = ($signed(_zz_256) - $signed(_zz_255));
  assign _zz_6898 = ($signed(_zz_255) + $signed(_zz_256));
  assign _zz_6899 = _zz_6900[15 : 0];
  assign _zz_6900 = fixTo_191_dout;
  assign _zz_6901 = _zz_6902[15 : 0];
  assign _zz_6902 = fixTo_190_dout;
  assign _zz_6903 = _zz_6904;
  assign _zz_6904 = ($signed(_zz_6905) >>> _zz_2111);
  assign _zz_6905 = _zz_6906;
  assign _zz_6906 = ($signed(_zz_253) - $signed(_zz_2108));
  assign _zz_6907 = _zz_6908;
  assign _zz_6908 = ($signed(_zz_6909) >>> _zz_2111);
  assign _zz_6909 = _zz_6910;
  assign _zz_6910 = ($signed(_zz_254) - $signed(_zz_2109));
  assign _zz_6911 = _zz_6912;
  assign _zz_6912 = ($signed(_zz_6913) >>> _zz_2112);
  assign _zz_6913 = _zz_6914;
  assign _zz_6914 = ($signed(_zz_253) + $signed(_zz_2108));
  assign _zz_6915 = _zz_6916;
  assign _zz_6916 = ($signed(_zz_6917) >>> _zz_2112);
  assign _zz_6917 = _zz_6918;
  assign _zz_6918 = ($signed(_zz_254) + $signed(_zz_2109));
  assign _zz_6919 = ($signed(twiddle_factor_table_1_real) + $signed(twiddle_factor_table_1_imag));
  assign _zz_6920 = fixTo_192_dout;
  assign _zz_6921 = ($signed(_zz_262) - $signed(_zz_261));
  assign _zz_6922 = ($signed(_zz_261) + $signed(_zz_262));
  assign _zz_6923 = _zz_6924[15 : 0];
  assign _zz_6924 = fixTo_194_dout;
  assign _zz_6925 = _zz_6926[15 : 0];
  assign _zz_6926 = fixTo_193_dout;
  assign _zz_6927 = _zz_6928;
  assign _zz_6928 = ($signed(_zz_6929) >>> _zz_2116);
  assign _zz_6929 = _zz_6930;
  assign _zz_6930 = ($signed(_zz_257) - $signed(_zz_2113));
  assign _zz_6931 = _zz_6932;
  assign _zz_6932 = ($signed(_zz_6933) >>> _zz_2116);
  assign _zz_6933 = _zz_6934;
  assign _zz_6934 = ($signed(_zz_258) - $signed(_zz_2114));
  assign _zz_6935 = _zz_6936;
  assign _zz_6936 = ($signed(_zz_6937) >>> _zz_2117);
  assign _zz_6937 = _zz_6938;
  assign _zz_6938 = ($signed(_zz_257) + $signed(_zz_2113));
  assign _zz_6939 = _zz_6940;
  assign _zz_6940 = ($signed(_zz_6941) >>> _zz_2117);
  assign _zz_6941 = _zz_6942;
  assign _zz_6942 = ($signed(_zz_258) + $signed(_zz_2114));
  assign _zz_6943 = ($signed(twiddle_factor_table_2_real) + $signed(twiddle_factor_table_2_imag));
  assign _zz_6944 = fixTo_195_dout;
  assign _zz_6945 = ($signed(_zz_264) - $signed(_zz_263));
  assign _zz_6946 = ($signed(_zz_263) + $signed(_zz_264));
  assign _zz_6947 = _zz_6948[15 : 0];
  assign _zz_6948 = fixTo_197_dout;
  assign _zz_6949 = _zz_6950[15 : 0];
  assign _zz_6950 = fixTo_196_dout;
  assign _zz_6951 = _zz_6952;
  assign _zz_6952 = ($signed(_zz_6953) >>> _zz_2121);
  assign _zz_6953 = _zz_6954;
  assign _zz_6954 = ($signed(_zz_259) - $signed(_zz_2118));
  assign _zz_6955 = _zz_6956;
  assign _zz_6956 = ($signed(_zz_6957) >>> _zz_2121);
  assign _zz_6957 = _zz_6958;
  assign _zz_6958 = ($signed(_zz_260) - $signed(_zz_2119));
  assign _zz_6959 = _zz_6960;
  assign _zz_6960 = ($signed(_zz_6961) >>> _zz_2122);
  assign _zz_6961 = _zz_6962;
  assign _zz_6962 = ($signed(_zz_259) + $signed(_zz_2118));
  assign _zz_6963 = _zz_6964;
  assign _zz_6964 = ($signed(_zz_6965) >>> _zz_2122);
  assign _zz_6965 = _zz_6966;
  assign _zz_6966 = ($signed(_zz_260) + $signed(_zz_2119));
  assign _zz_6967 = ($signed(twiddle_factor_table_1_real) + $signed(twiddle_factor_table_1_imag));
  assign _zz_6968 = fixTo_198_dout;
  assign _zz_6969 = ($signed(_zz_270) - $signed(_zz_269));
  assign _zz_6970 = ($signed(_zz_269) + $signed(_zz_270));
  assign _zz_6971 = _zz_6972[15 : 0];
  assign _zz_6972 = fixTo_200_dout;
  assign _zz_6973 = _zz_6974[15 : 0];
  assign _zz_6974 = fixTo_199_dout;
  assign _zz_6975 = _zz_6976;
  assign _zz_6976 = ($signed(_zz_6977) >>> _zz_2126);
  assign _zz_6977 = _zz_6978;
  assign _zz_6978 = ($signed(_zz_265) - $signed(_zz_2123));
  assign _zz_6979 = _zz_6980;
  assign _zz_6980 = ($signed(_zz_6981) >>> _zz_2126);
  assign _zz_6981 = _zz_6982;
  assign _zz_6982 = ($signed(_zz_266) - $signed(_zz_2124));
  assign _zz_6983 = _zz_6984;
  assign _zz_6984 = ($signed(_zz_6985) >>> _zz_2127);
  assign _zz_6985 = _zz_6986;
  assign _zz_6986 = ($signed(_zz_265) + $signed(_zz_2123));
  assign _zz_6987 = _zz_6988;
  assign _zz_6988 = ($signed(_zz_6989) >>> _zz_2127);
  assign _zz_6989 = _zz_6990;
  assign _zz_6990 = ($signed(_zz_266) + $signed(_zz_2124));
  assign _zz_6991 = ($signed(twiddle_factor_table_2_real) + $signed(twiddle_factor_table_2_imag));
  assign _zz_6992 = fixTo_201_dout;
  assign _zz_6993 = ($signed(_zz_272) - $signed(_zz_271));
  assign _zz_6994 = ($signed(_zz_271) + $signed(_zz_272));
  assign _zz_6995 = _zz_6996[15 : 0];
  assign _zz_6996 = fixTo_203_dout;
  assign _zz_6997 = _zz_6998[15 : 0];
  assign _zz_6998 = fixTo_202_dout;
  assign _zz_6999 = _zz_7000;
  assign _zz_7000 = ($signed(_zz_7001) >>> _zz_2131);
  assign _zz_7001 = _zz_7002;
  assign _zz_7002 = ($signed(_zz_267) - $signed(_zz_2128));
  assign _zz_7003 = _zz_7004;
  assign _zz_7004 = ($signed(_zz_7005) >>> _zz_2131);
  assign _zz_7005 = _zz_7006;
  assign _zz_7006 = ($signed(_zz_268) - $signed(_zz_2129));
  assign _zz_7007 = _zz_7008;
  assign _zz_7008 = ($signed(_zz_7009) >>> _zz_2132);
  assign _zz_7009 = _zz_7010;
  assign _zz_7010 = ($signed(_zz_267) + $signed(_zz_2128));
  assign _zz_7011 = _zz_7012;
  assign _zz_7012 = ($signed(_zz_7013) >>> _zz_2132);
  assign _zz_7013 = _zz_7014;
  assign _zz_7014 = ($signed(_zz_268) + $signed(_zz_2129));
  assign _zz_7015 = ($signed(twiddle_factor_table_1_real) + $signed(twiddle_factor_table_1_imag));
  assign _zz_7016 = fixTo_204_dout;
  assign _zz_7017 = ($signed(_zz_278) - $signed(_zz_277));
  assign _zz_7018 = ($signed(_zz_277) + $signed(_zz_278));
  assign _zz_7019 = _zz_7020[15 : 0];
  assign _zz_7020 = fixTo_206_dout;
  assign _zz_7021 = _zz_7022[15 : 0];
  assign _zz_7022 = fixTo_205_dout;
  assign _zz_7023 = _zz_7024;
  assign _zz_7024 = ($signed(_zz_7025) >>> _zz_2136);
  assign _zz_7025 = _zz_7026;
  assign _zz_7026 = ($signed(_zz_273) - $signed(_zz_2133));
  assign _zz_7027 = _zz_7028;
  assign _zz_7028 = ($signed(_zz_7029) >>> _zz_2136);
  assign _zz_7029 = _zz_7030;
  assign _zz_7030 = ($signed(_zz_274) - $signed(_zz_2134));
  assign _zz_7031 = _zz_7032;
  assign _zz_7032 = ($signed(_zz_7033) >>> _zz_2137);
  assign _zz_7033 = _zz_7034;
  assign _zz_7034 = ($signed(_zz_273) + $signed(_zz_2133));
  assign _zz_7035 = _zz_7036;
  assign _zz_7036 = ($signed(_zz_7037) >>> _zz_2137);
  assign _zz_7037 = _zz_7038;
  assign _zz_7038 = ($signed(_zz_274) + $signed(_zz_2134));
  assign _zz_7039 = ($signed(twiddle_factor_table_2_real) + $signed(twiddle_factor_table_2_imag));
  assign _zz_7040 = fixTo_207_dout;
  assign _zz_7041 = ($signed(_zz_280) - $signed(_zz_279));
  assign _zz_7042 = ($signed(_zz_279) + $signed(_zz_280));
  assign _zz_7043 = _zz_7044[15 : 0];
  assign _zz_7044 = fixTo_209_dout;
  assign _zz_7045 = _zz_7046[15 : 0];
  assign _zz_7046 = fixTo_208_dout;
  assign _zz_7047 = _zz_7048;
  assign _zz_7048 = ($signed(_zz_7049) >>> _zz_2141);
  assign _zz_7049 = _zz_7050;
  assign _zz_7050 = ($signed(_zz_275) - $signed(_zz_2138));
  assign _zz_7051 = _zz_7052;
  assign _zz_7052 = ($signed(_zz_7053) >>> _zz_2141);
  assign _zz_7053 = _zz_7054;
  assign _zz_7054 = ($signed(_zz_276) - $signed(_zz_2139));
  assign _zz_7055 = _zz_7056;
  assign _zz_7056 = ($signed(_zz_7057) >>> _zz_2142);
  assign _zz_7057 = _zz_7058;
  assign _zz_7058 = ($signed(_zz_275) + $signed(_zz_2138));
  assign _zz_7059 = _zz_7060;
  assign _zz_7060 = ($signed(_zz_7061) >>> _zz_2142);
  assign _zz_7061 = _zz_7062;
  assign _zz_7062 = ($signed(_zz_276) + $signed(_zz_2139));
  assign _zz_7063 = ($signed(twiddle_factor_table_1_real) + $signed(twiddle_factor_table_1_imag));
  assign _zz_7064 = fixTo_210_dout;
  assign _zz_7065 = ($signed(_zz_286) - $signed(_zz_285));
  assign _zz_7066 = ($signed(_zz_285) + $signed(_zz_286));
  assign _zz_7067 = _zz_7068[15 : 0];
  assign _zz_7068 = fixTo_212_dout;
  assign _zz_7069 = _zz_7070[15 : 0];
  assign _zz_7070 = fixTo_211_dout;
  assign _zz_7071 = _zz_7072;
  assign _zz_7072 = ($signed(_zz_7073) >>> _zz_2146);
  assign _zz_7073 = _zz_7074;
  assign _zz_7074 = ($signed(_zz_281) - $signed(_zz_2143));
  assign _zz_7075 = _zz_7076;
  assign _zz_7076 = ($signed(_zz_7077) >>> _zz_2146);
  assign _zz_7077 = _zz_7078;
  assign _zz_7078 = ($signed(_zz_282) - $signed(_zz_2144));
  assign _zz_7079 = _zz_7080;
  assign _zz_7080 = ($signed(_zz_7081) >>> _zz_2147);
  assign _zz_7081 = _zz_7082;
  assign _zz_7082 = ($signed(_zz_281) + $signed(_zz_2143));
  assign _zz_7083 = _zz_7084;
  assign _zz_7084 = ($signed(_zz_7085) >>> _zz_2147);
  assign _zz_7085 = _zz_7086;
  assign _zz_7086 = ($signed(_zz_282) + $signed(_zz_2144));
  assign _zz_7087 = ($signed(twiddle_factor_table_2_real) + $signed(twiddle_factor_table_2_imag));
  assign _zz_7088 = fixTo_213_dout;
  assign _zz_7089 = ($signed(_zz_288) - $signed(_zz_287));
  assign _zz_7090 = ($signed(_zz_287) + $signed(_zz_288));
  assign _zz_7091 = _zz_7092[15 : 0];
  assign _zz_7092 = fixTo_215_dout;
  assign _zz_7093 = _zz_7094[15 : 0];
  assign _zz_7094 = fixTo_214_dout;
  assign _zz_7095 = _zz_7096;
  assign _zz_7096 = ($signed(_zz_7097) >>> _zz_2151);
  assign _zz_7097 = _zz_7098;
  assign _zz_7098 = ($signed(_zz_283) - $signed(_zz_2148));
  assign _zz_7099 = _zz_7100;
  assign _zz_7100 = ($signed(_zz_7101) >>> _zz_2151);
  assign _zz_7101 = _zz_7102;
  assign _zz_7102 = ($signed(_zz_284) - $signed(_zz_2149));
  assign _zz_7103 = _zz_7104;
  assign _zz_7104 = ($signed(_zz_7105) >>> _zz_2152);
  assign _zz_7105 = _zz_7106;
  assign _zz_7106 = ($signed(_zz_283) + $signed(_zz_2148));
  assign _zz_7107 = _zz_7108;
  assign _zz_7108 = ($signed(_zz_7109) >>> _zz_2152);
  assign _zz_7109 = _zz_7110;
  assign _zz_7110 = ($signed(_zz_284) + $signed(_zz_2149));
  assign _zz_7111 = ($signed(twiddle_factor_table_1_real) + $signed(twiddle_factor_table_1_imag));
  assign _zz_7112 = fixTo_216_dout;
  assign _zz_7113 = ($signed(_zz_294) - $signed(_zz_293));
  assign _zz_7114 = ($signed(_zz_293) + $signed(_zz_294));
  assign _zz_7115 = _zz_7116[15 : 0];
  assign _zz_7116 = fixTo_218_dout;
  assign _zz_7117 = _zz_7118[15 : 0];
  assign _zz_7118 = fixTo_217_dout;
  assign _zz_7119 = _zz_7120;
  assign _zz_7120 = ($signed(_zz_7121) >>> _zz_2156);
  assign _zz_7121 = _zz_7122;
  assign _zz_7122 = ($signed(_zz_289) - $signed(_zz_2153));
  assign _zz_7123 = _zz_7124;
  assign _zz_7124 = ($signed(_zz_7125) >>> _zz_2156);
  assign _zz_7125 = _zz_7126;
  assign _zz_7126 = ($signed(_zz_290) - $signed(_zz_2154));
  assign _zz_7127 = _zz_7128;
  assign _zz_7128 = ($signed(_zz_7129) >>> _zz_2157);
  assign _zz_7129 = _zz_7130;
  assign _zz_7130 = ($signed(_zz_289) + $signed(_zz_2153));
  assign _zz_7131 = _zz_7132;
  assign _zz_7132 = ($signed(_zz_7133) >>> _zz_2157);
  assign _zz_7133 = _zz_7134;
  assign _zz_7134 = ($signed(_zz_290) + $signed(_zz_2154));
  assign _zz_7135 = ($signed(twiddle_factor_table_2_real) + $signed(twiddle_factor_table_2_imag));
  assign _zz_7136 = fixTo_219_dout;
  assign _zz_7137 = ($signed(_zz_296) - $signed(_zz_295));
  assign _zz_7138 = ($signed(_zz_295) + $signed(_zz_296));
  assign _zz_7139 = _zz_7140[15 : 0];
  assign _zz_7140 = fixTo_221_dout;
  assign _zz_7141 = _zz_7142[15 : 0];
  assign _zz_7142 = fixTo_220_dout;
  assign _zz_7143 = _zz_7144;
  assign _zz_7144 = ($signed(_zz_7145) >>> _zz_2161);
  assign _zz_7145 = _zz_7146;
  assign _zz_7146 = ($signed(_zz_291) - $signed(_zz_2158));
  assign _zz_7147 = _zz_7148;
  assign _zz_7148 = ($signed(_zz_7149) >>> _zz_2161);
  assign _zz_7149 = _zz_7150;
  assign _zz_7150 = ($signed(_zz_292) - $signed(_zz_2159));
  assign _zz_7151 = _zz_7152;
  assign _zz_7152 = ($signed(_zz_7153) >>> _zz_2162);
  assign _zz_7153 = _zz_7154;
  assign _zz_7154 = ($signed(_zz_291) + $signed(_zz_2158));
  assign _zz_7155 = _zz_7156;
  assign _zz_7156 = ($signed(_zz_7157) >>> _zz_2162);
  assign _zz_7157 = _zz_7158;
  assign _zz_7158 = ($signed(_zz_292) + $signed(_zz_2159));
  assign _zz_7159 = ($signed(twiddle_factor_table_1_real) + $signed(twiddle_factor_table_1_imag));
  assign _zz_7160 = fixTo_222_dout;
  assign _zz_7161 = ($signed(_zz_302) - $signed(_zz_301));
  assign _zz_7162 = ($signed(_zz_301) + $signed(_zz_302));
  assign _zz_7163 = _zz_7164[15 : 0];
  assign _zz_7164 = fixTo_224_dout;
  assign _zz_7165 = _zz_7166[15 : 0];
  assign _zz_7166 = fixTo_223_dout;
  assign _zz_7167 = _zz_7168;
  assign _zz_7168 = ($signed(_zz_7169) >>> _zz_2166);
  assign _zz_7169 = _zz_7170;
  assign _zz_7170 = ($signed(_zz_297) - $signed(_zz_2163));
  assign _zz_7171 = _zz_7172;
  assign _zz_7172 = ($signed(_zz_7173) >>> _zz_2166);
  assign _zz_7173 = _zz_7174;
  assign _zz_7174 = ($signed(_zz_298) - $signed(_zz_2164));
  assign _zz_7175 = _zz_7176;
  assign _zz_7176 = ($signed(_zz_7177) >>> _zz_2167);
  assign _zz_7177 = _zz_7178;
  assign _zz_7178 = ($signed(_zz_297) + $signed(_zz_2163));
  assign _zz_7179 = _zz_7180;
  assign _zz_7180 = ($signed(_zz_7181) >>> _zz_2167);
  assign _zz_7181 = _zz_7182;
  assign _zz_7182 = ($signed(_zz_298) + $signed(_zz_2164));
  assign _zz_7183 = ($signed(twiddle_factor_table_2_real) + $signed(twiddle_factor_table_2_imag));
  assign _zz_7184 = fixTo_225_dout;
  assign _zz_7185 = ($signed(_zz_304) - $signed(_zz_303));
  assign _zz_7186 = ($signed(_zz_303) + $signed(_zz_304));
  assign _zz_7187 = _zz_7188[15 : 0];
  assign _zz_7188 = fixTo_227_dout;
  assign _zz_7189 = _zz_7190[15 : 0];
  assign _zz_7190 = fixTo_226_dout;
  assign _zz_7191 = _zz_7192;
  assign _zz_7192 = ($signed(_zz_7193) >>> _zz_2171);
  assign _zz_7193 = _zz_7194;
  assign _zz_7194 = ($signed(_zz_299) - $signed(_zz_2168));
  assign _zz_7195 = _zz_7196;
  assign _zz_7196 = ($signed(_zz_7197) >>> _zz_2171);
  assign _zz_7197 = _zz_7198;
  assign _zz_7198 = ($signed(_zz_300) - $signed(_zz_2169));
  assign _zz_7199 = _zz_7200;
  assign _zz_7200 = ($signed(_zz_7201) >>> _zz_2172);
  assign _zz_7201 = _zz_7202;
  assign _zz_7202 = ($signed(_zz_299) + $signed(_zz_2168));
  assign _zz_7203 = _zz_7204;
  assign _zz_7204 = ($signed(_zz_7205) >>> _zz_2172);
  assign _zz_7205 = _zz_7206;
  assign _zz_7206 = ($signed(_zz_300) + $signed(_zz_2169));
  assign _zz_7207 = ($signed(twiddle_factor_table_1_real) + $signed(twiddle_factor_table_1_imag));
  assign _zz_7208 = fixTo_228_dout;
  assign _zz_7209 = ($signed(_zz_310) - $signed(_zz_309));
  assign _zz_7210 = ($signed(_zz_309) + $signed(_zz_310));
  assign _zz_7211 = _zz_7212[15 : 0];
  assign _zz_7212 = fixTo_230_dout;
  assign _zz_7213 = _zz_7214[15 : 0];
  assign _zz_7214 = fixTo_229_dout;
  assign _zz_7215 = _zz_7216;
  assign _zz_7216 = ($signed(_zz_7217) >>> _zz_2176);
  assign _zz_7217 = _zz_7218;
  assign _zz_7218 = ($signed(_zz_305) - $signed(_zz_2173));
  assign _zz_7219 = _zz_7220;
  assign _zz_7220 = ($signed(_zz_7221) >>> _zz_2176);
  assign _zz_7221 = _zz_7222;
  assign _zz_7222 = ($signed(_zz_306) - $signed(_zz_2174));
  assign _zz_7223 = _zz_7224;
  assign _zz_7224 = ($signed(_zz_7225) >>> _zz_2177);
  assign _zz_7225 = _zz_7226;
  assign _zz_7226 = ($signed(_zz_305) + $signed(_zz_2173));
  assign _zz_7227 = _zz_7228;
  assign _zz_7228 = ($signed(_zz_7229) >>> _zz_2177);
  assign _zz_7229 = _zz_7230;
  assign _zz_7230 = ($signed(_zz_306) + $signed(_zz_2174));
  assign _zz_7231 = ($signed(twiddle_factor_table_2_real) + $signed(twiddle_factor_table_2_imag));
  assign _zz_7232 = fixTo_231_dout;
  assign _zz_7233 = ($signed(_zz_312) - $signed(_zz_311));
  assign _zz_7234 = ($signed(_zz_311) + $signed(_zz_312));
  assign _zz_7235 = _zz_7236[15 : 0];
  assign _zz_7236 = fixTo_233_dout;
  assign _zz_7237 = _zz_7238[15 : 0];
  assign _zz_7238 = fixTo_232_dout;
  assign _zz_7239 = _zz_7240;
  assign _zz_7240 = ($signed(_zz_7241) >>> _zz_2181);
  assign _zz_7241 = _zz_7242;
  assign _zz_7242 = ($signed(_zz_307) - $signed(_zz_2178));
  assign _zz_7243 = _zz_7244;
  assign _zz_7244 = ($signed(_zz_7245) >>> _zz_2181);
  assign _zz_7245 = _zz_7246;
  assign _zz_7246 = ($signed(_zz_308) - $signed(_zz_2179));
  assign _zz_7247 = _zz_7248;
  assign _zz_7248 = ($signed(_zz_7249) >>> _zz_2182);
  assign _zz_7249 = _zz_7250;
  assign _zz_7250 = ($signed(_zz_307) + $signed(_zz_2178));
  assign _zz_7251 = _zz_7252;
  assign _zz_7252 = ($signed(_zz_7253) >>> _zz_2182);
  assign _zz_7253 = _zz_7254;
  assign _zz_7254 = ($signed(_zz_308) + $signed(_zz_2179));
  assign _zz_7255 = ($signed(twiddle_factor_table_1_real) + $signed(twiddle_factor_table_1_imag));
  assign _zz_7256 = fixTo_234_dout;
  assign _zz_7257 = ($signed(_zz_318) - $signed(_zz_317));
  assign _zz_7258 = ($signed(_zz_317) + $signed(_zz_318));
  assign _zz_7259 = _zz_7260[15 : 0];
  assign _zz_7260 = fixTo_236_dout;
  assign _zz_7261 = _zz_7262[15 : 0];
  assign _zz_7262 = fixTo_235_dout;
  assign _zz_7263 = _zz_7264;
  assign _zz_7264 = ($signed(_zz_7265) >>> _zz_2186);
  assign _zz_7265 = _zz_7266;
  assign _zz_7266 = ($signed(_zz_313) - $signed(_zz_2183));
  assign _zz_7267 = _zz_7268;
  assign _zz_7268 = ($signed(_zz_7269) >>> _zz_2186);
  assign _zz_7269 = _zz_7270;
  assign _zz_7270 = ($signed(_zz_314) - $signed(_zz_2184));
  assign _zz_7271 = _zz_7272;
  assign _zz_7272 = ($signed(_zz_7273) >>> _zz_2187);
  assign _zz_7273 = _zz_7274;
  assign _zz_7274 = ($signed(_zz_313) + $signed(_zz_2183));
  assign _zz_7275 = _zz_7276;
  assign _zz_7276 = ($signed(_zz_7277) >>> _zz_2187);
  assign _zz_7277 = _zz_7278;
  assign _zz_7278 = ($signed(_zz_314) + $signed(_zz_2184));
  assign _zz_7279 = ($signed(twiddle_factor_table_2_real) + $signed(twiddle_factor_table_2_imag));
  assign _zz_7280 = fixTo_237_dout;
  assign _zz_7281 = ($signed(_zz_320) - $signed(_zz_319));
  assign _zz_7282 = ($signed(_zz_319) + $signed(_zz_320));
  assign _zz_7283 = _zz_7284[15 : 0];
  assign _zz_7284 = fixTo_239_dout;
  assign _zz_7285 = _zz_7286[15 : 0];
  assign _zz_7286 = fixTo_238_dout;
  assign _zz_7287 = _zz_7288;
  assign _zz_7288 = ($signed(_zz_7289) >>> _zz_2191);
  assign _zz_7289 = _zz_7290;
  assign _zz_7290 = ($signed(_zz_315) - $signed(_zz_2188));
  assign _zz_7291 = _zz_7292;
  assign _zz_7292 = ($signed(_zz_7293) >>> _zz_2191);
  assign _zz_7293 = _zz_7294;
  assign _zz_7294 = ($signed(_zz_316) - $signed(_zz_2189));
  assign _zz_7295 = _zz_7296;
  assign _zz_7296 = ($signed(_zz_7297) >>> _zz_2192);
  assign _zz_7297 = _zz_7298;
  assign _zz_7298 = ($signed(_zz_315) + $signed(_zz_2188));
  assign _zz_7299 = _zz_7300;
  assign _zz_7300 = ($signed(_zz_7301) >>> _zz_2192);
  assign _zz_7301 = _zz_7302;
  assign _zz_7302 = ($signed(_zz_316) + $signed(_zz_2189));
  assign _zz_7303 = ($signed(twiddle_factor_table_1_real) + $signed(twiddle_factor_table_1_imag));
  assign _zz_7304 = fixTo_240_dout;
  assign _zz_7305 = ($signed(_zz_326) - $signed(_zz_325));
  assign _zz_7306 = ($signed(_zz_325) + $signed(_zz_326));
  assign _zz_7307 = _zz_7308[15 : 0];
  assign _zz_7308 = fixTo_242_dout;
  assign _zz_7309 = _zz_7310[15 : 0];
  assign _zz_7310 = fixTo_241_dout;
  assign _zz_7311 = _zz_7312;
  assign _zz_7312 = ($signed(_zz_7313) >>> _zz_2196);
  assign _zz_7313 = _zz_7314;
  assign _zz_7314 = ($signed(_zz_321) - $signed(_zz_2193));
  assign _zz_7315 = _zz_7316;
  assign _zz_7316 = ($signed(_zz_7317) >>> _zz_2196);
  assign _zz_7317 = _zz_7318;
  assign _zz_7318 = ($signed(_zz_322) - $signed(_zz_2194));
  assign _zz_7319 = _zz_7320;
  assign _zz_7320 = ($signed(_zz_7321) >>> _zz_2197);
  assign _zz_7321 = _zz_7322;
  assign _zz_7322 = ($signed(_zz_321) + $signed(_zz_2193));
  assign _zz_7323 = _zz_7324;
  assign _zz_7324 = ($signed(_zz_7325) >>> _zz_2197);
  assign _zz_7325 = _zz_7326;
  assign _zz_7326 = ($signed(_zz_322) + $signed(_zz_2194));
  assign _zz_7327 = ($signed(twiddle_factor_table_2_real) + $signed(twiddle_factor_table_2_imag));
  assign _zz_7328 = fixTo_243_dout;
  assign _zz_7329 = ($signed(_zz_328) - $signed(_zz_327));
  assign _zz_7330 = ($signed(_zz_327) + $signed(_zz_328));
  assign _zz_7331 = _zz_7332[15 : 0];
  assign _zz_7332 = fixTo_245_dout;
  assign _zz_7333 = _zz_7334[15 : 0];
  assign _zz_7334 = fixTo_244_dout;
  assign _zz_7335 = _zz_7336;
  assign _zz_7336 = ($signed(_zz_7337) >>> _zz_2201);
  assign _zz_7337 = _zz_7338;
  assign _zz_7338 = ($signed(_zz_323) - $signed(_zz_2198));
  assign _zz_7339 = _zz_7340;
  assign _zz_7340 = ($signed(_zz_7341) >>> _zz_2201);
  assign _zz_7341 = _zz_7342;
  assign _zz_7342 = ($signed(_zz_324) - $signed(_zz_2199));
  assign _zz_7343 = _zz_7344;
  assign _zz_7344 = ($signed(_zz_7345) >>> _zz_2202);
  assign _zz_7345 = _zz_7346;
  assign _zz_7346 = ($signed(_zz_323) + $signed(_zz_2198));
  assign _zz_7347 = _zz_7348;
  assign _zz_7348 = ($signed(_zz_7349) >>> _zz_2202);
  assign _zz_7349 = _zz_7350;
  assign _zz_7350 = ($signed(_zz_324) + $signed(_zz_2199));
  assign _zz_7351 = ($signed(twiddle_factor_table_1_real) + $signed(twiddle_factor_table_1_imag));
  assign _zz_7352 = fixTo_246_dout;
  assign _zz_7353 = ($signed(_zz_334) - $signed(_zz_333));
  assign _zz_7354 = ($signed(_zz_333) + $signed(_zz_334));
  assign _zz_7355 = _zz_7356[15 : 0];
  assign _zz_7356 = fixTo_248_dout;
  assign _zz_7357 = _zz_7358[15 : 0];
  assign _zz_7358 = fixTo_247_dout;
  assign _zz_7359 = _zz_7360;
  assign _zz_7360 = ($signed(_zz_7361) >>> _zz_2206);
  assign _zz_7361 = _zz_7362;
  assign _zz_7362 = ($signed(_zz_329) - $signed(_zz_2203));
  assign _zz_7363 = _zz_7364;
  assign _zz_7364 = ($signed(_zz_7365) >>> _zz_2206);
  assign _zz_7365 = _zz_7366;
  assign _zz_7366 = ($signed(_zz_330) - $signed(_zz_2204));
  assign _zz_7367 = _zz_7368;
  assign _zz_7368 = ($signed(_zz_7369) >>> _zz_2207);
  assign _zz_7369 = _zz_7370;
  assign _zz_7370 = ($signed(_zz_329) + $signed(_zz_2203));
  assign _zz_7371 = _zz_7372;
  assign _zz_7372 = ($signed(_zz_7373) >>> _zz_2207);
  assign _zz_7373 = _zz_7374;
  assign _zz_7374 = ($signed(_zz_330) + $signed(_zz_2204));
  assign _zz_7375 = ($signed(twiddle_factor_table_2_real) + $signed(twiddle_factor_table_2_imag));
  assign _zz_7376 = fixTo_249_dout;
  assign _zz_7377 = ($signed(_zz_336) - $signed(_zz_335));
  assign _zz_7378 = ($signed(_zz_335) + $signed(_zz_336));
  assign _zz_7379 = _zz_7380[15 : 0];
  assign _zz_7380 = fixTo_251_dout;
  assign _zz_7381 = _zz_7382[15 : 0];
  assign _zz_7382 = fixTo_250_dout;
  assign _zz_7383 = _zz_7384;
  assign _zz_7384 = ($signed(_zz_7385) >>> _zz_2211);
  assign _zz_7385 = _zz_7386;
  assign _zz_7386 = ($signed(_zz_331) - $signed(_zz_2208));
  assign _zz_7387 = _zz_7388;
  assign _zz_7388 = ($signed(_zz_7389) >>> _zz_2211);
  assign _zz_7389 = _zz_7390;
  assign _zz_7390 = ($signed(_zz_332) - $signed(_zz_2209));
  assign _zz_7391 = _zz_7392;
  assign _zz_7392 = ($signed(_zz_7393) >>> _zz_2212);
  assign _zz_7393 = _zz_7394;
  assign _zz_7394 = ($signed(_zz_331) + $signed(_zz_2208));
  assign _zz_7395 = _zz_7396;
  assign _zz_7396 = ($signed(_zz_7397) >>> _zz_2212);
  assign _zz_7397 = _zz_7398;
  assign _zz_7398 = ($signed(_zz_332) + $signed(_zz_2209));
  assign _zz_7399 = ($signed(twiddle_factor_table_1_real) + $signed(twiddle_factor_table_1_imag));
  assign _zz_7400 = fixTo_252_dout;
  assign _zz_7401 = ($signed(_zz_342) - $signed(_zz_341));
  assign _zz_7402 = ($signed(_zz_341) + $signed(_zz_342));
  assign _zz_7403 = _zz_7404[15 : 0];
  assign _zz_7404 = fixTo_254_dout;
  assign _zz_7405 = _zz_7406[15 : 0];
  assign _zz_7406 = fixTo_253_dout;
  assign _zz_7407 = _zz_7408;
  assign _zz_7408 = ($signed(_zz_7409) >>> _zz_2216);
  assign _zz_7409 = _zz_7410;
  assign _zz_7410 = ($signed(_zz_337) - $signed(_zz_2213));
  assign _zz_7411 = _zz_7412;
  assign _zz_7412 = ($signed(_zz_7413) >>> _zz_2216);
  assign _zz_7413 = _zz_7414;
  assign _zz_7414 = ($signed(_zz_338) - $signed(_zz_2214));
  assign _zz_7415 = _zz_7416;
  assign _zz_7416 = ($signed(_zz_7417) >>> _zz_2217);
  assign _zz_7417 = _zz_7418;
  assign _zz_7418 = ($signed(_zz_337) + $signed(_zz_2213));
  assign _zz_7419 = _zz_7420;
  assign _zz_7420 = ($signed(_zz_7421) >>> _zz_2217);
  assign _zz_7421 = _zz_7422;
  assign _zz_7422 = ($signed(_zz_338) + $signed(_zz_2214));
  assign _zz_7423 = ($signed(twiddle_factor_table_2_real) + $signed(twiddle_factor_table_2_imag));
  assign _zz_7424 = fixTo_255_dout;
  assign _zz_7425 = ($signed(_zz_344) - $signed(_zz_343));
  assign _zz_7426 = ($signed(_zz_343) + $signed(_zz_344));
  assign _zz_7427 = _zz_7428[15 : 0];
  assign _zz_7428 = fixTo_257_dout;
  assign _zz_7429 = _zz_7430[15 : 0];
  assign _zz_7430 = fixTo_256_dout;
  assign _zz_7431 = _zz_7432;
  assign _zz_7432 = ($signed(_zz_7433) >>> _zz_2221);
  assign _zz_7433 = _zz_7434;
  assign _zz_7434 = ($signed(_zz_339) - $signed(_zz_2218));
  assign _zz_7435 = _zz_7436;
  assign _zz_7436 = ($signed(_zz_7437) >>> _zz_2221);
  assign _zz_7437 = _zz_7438;
  assign _zz_7438 = ($signed(_zz_340) - $signed(_zz_2219));
  assign _zz_7439 = _zz_7440;
  assign _zz_7440 = ($signed(_zz_7441) >>> _zz_2222);
  assign _zz_7441 = _zz_7442;
  assign _zz_7442 = ($signed(_zz_339) + $signed(_zz_2218));
  assign _zz_7443 = _zz_7444;
  assign _zz_7444 = ($signed(_zz_7445) >>> _zz_2222);
  assign _zz_7445 = _zz_7446;
  assign _zz_7446 = ($signed(_zz_340) + $signed(_zz_2219));
  assign _zz_7447 = ($signed(twiddle_factor_table_1_real) + $signed(twiddle_factor_table_1_imag));
  assign _zz_7448 = fixTo_258_dout;
  assign _zz_7449 = ($signed(_zz_350) - $signed(_zz_349));
  assign _zz_7450 = ($signed(_zz_349) + $signed(_zz_350));
  assign _zz_7451 = _zz_7452[15 : 0];
  assign _zz_7452 = fixTo_260_dout;
  assign _zz_7453 = _zz_7454[15 : 0];
  assign _zz_7454 = fixTo_259_dout;
  assign _zz_7455 = _zz_7456;
  assign _zz_7456 = ($signed(_zz_7457) >>> _zz_2226);
  assign _zz_7457 = _zz_7458;
  assign _zz_7458 = ($signed(_zz_345) - $signed(_zz_2223));
  assign _zz_7459 = _zz_7460;
  assign _zz_7460 = ($signed(_zz_7461) >>> _zz_2226);
  assign _zz_7461 = _zz_7462;
  assign _zz_7462 = ($signed(_zz_346) - $signed(_zz_2224));
  assign _zz_7463 = _zz_7464;
  assign _zz_7464 = ($signed(_zz_7465) >>> _zz_2227);
  assign _zz_7465 = _zz_7466;
  assign _zz_7466 = ($signed(_zz_345) + $signed(_zz_2223));
  assign _zz_7467 = _zz_7468;
  assign _zz_7468 = ($signed(_zz_7469) >>> _zz_2227);
  assign _zz_7469 = _zz_7470;
  assign _zz_7470 = ($signed(_zz_346) + $signed(_zz_2224));
  assign _zz_7471 = ($signed(twiddle_factor_table_2_real) + $signed(twiddle_factor_table_2_imag));
  assign _zz_7472 = fixTo_261_dout;
  assign _zz_7473 = ($signed(_zz_352) - $signed(_zz_351));
  assign _zz_7474 = ($signed(_zz_351) + $signed(_zz_352));
  assign _zz_7475 = _zz_7476[15 : 0];
  assign _zz_7476 = fixTo_263_dout;
  assign _zz_7477 = _zz_7478[15 : 0];
  assign _zz_7478 = fixTo_262_dout;
  assign _zz_7479 = _zz_7480;
  assign _zz_7480 = ($signed(_zz_7481) >>> _zz_2231);
  assign _zz_7481 = _zz_7482;
  assign _zz_7482 = ($signed(_zz_347) - $signed(_zz_2228));
  assign _zz_7483 = _zz_7484;
  assign _zz_7484 = ($signed(_zz_7485) >>> _zz_2231);
  assign _zz_7485 = _zz_7486;
  assign _zz_7486 = ($signed(_zz_348) - $signed(_zz_2229));
  assign _zz_7487 = _zz_7488;
  assign _zz_7488 = ($signed(_zz_7489) >>> _zz_2232);
  assign _zz_7489 = _zz_7490;
  assign _zz_7490 = ($signed(_zz_347) + $signed(_zz_2228));
  assign _zz_7491 = _zz_7492;
  assign _zz_7492 = ($signed(_zz_7493) >>> _zz_2232);
  assign _zz_7493 = _zz_7494;
  assign _zz_7494 = ($signed(_zz_348) + $signed(_zz_2229));
  assign _zz_7495 = ($signed(twiddle_factor_table_1_real) + $signed(twiddle_factor_table_1_imag));
  assign _zz_7496 = fixTo_264_dout;
  assign _zz_7497 = ($signed(_zz_358) - $signed(_zz_357));
  assign _zz_7498 = ($signed(_zz_357) + $signed(_zz_358));
  assign _zz_7499 = _zz_7500[15 : 0];
  assign _zz_7500 = fixTo_266_dout;
  assign _zz_7501 = _zz_7502[15 : 0];
  assign _zz_7502 = fixTo_265_dout;
  assign _zz_7503 = _zz_7504;
  assign _zz_7504 = ($signed(_zz_7505) >>> _zz_2236);
  assign _zz_7505 = _zz_7506;
  assign _zz_7506 = ($signed(_zz_353) - $signed(_zz_2233));
  assign _zz_7507 = _zz_7508;
  assign _zz_7508 = ($signed(_zz_7509) >>> _zz_2236);
  assign _zz_7509 = _zz_7510;
  assign _zz_7510 = ($signed(_zz_354) - $signed(_zz_2234));
  assign _zz_7511 = _zz_7512;
  assign _zz_7512 = ($signed(_zz_7513) >>> _zz_2237);
  assign _zz_7513 = _zz_7514;
  assign _zz_7514 = ($signed(_zz_353) + $signed(_zz_2233));
  assign _zz_7515 = _zz_7516;
  assign _zz_7516 = ($signed(_zz_7517) >>> _zz_2237);
  assign _zz_7517 = _zz_7518;
  assign _zz_7518 = ($signed(_zz_354) + $signed(_zz_2234));
  assign _zz_7519 = ($signed(twiddle_factor_table_2_real) + $signed(twiddle_factor_table_2_imag));
  assign _zz_7520 = fixTo_267_dout;
  assign _zz_7521 = ($signed(_zz_360) - $signed(_zz_359));
  assign _zz_7522 = ($signed(_zz_359) + $signed(_zz_360));
  assign _zz_7523 = _zz_7524[15 : 0];
  assign _zz_7524 = fixTo_269_dout;
  assign _zz_7525 = _zz_7526[15 : 0];
  assign _zz_7526 = fixTo_268_dout;
  assign _zz_7527 = _zz_7528;
  assign _zz_7528 = ($signed(_zz_7529) >>> _zz_2241);
  assign _zz_7529 = _zz_7530;
  assign _zz_7530 = ($signed(_zz_355) - $signed(_zz_2238));
  assign _zz_7531 = _zz_7532;
  assign _zz_7532 = ($signed(_zz_7533) >>> _zz_2241);
  assign _zz_7533 = _zz_7534;
  assign _zz_7534 = ($signed(_zz_356) - $signed(_zz_2239));
  assign _zz_7535 = _zz_7536;
  assign _zz_7536 = ($signed(_zz_7537) >>> _zz_2242);
  assign _zz_7537 = _zz_7538;
  assign _zz_7538 = ($signed(_zz_355) + $signed(_zz_2238));
  assign _zz_7539 = _zz_7540;
  assign _zz_7540 = ($signed(_zz_7541) >>> _zz_2242);
  assign _zz_7541 = _zz_7542;
  assign _zz_7542 = ($signed(_zz_356) + $signed(_zz_2239));
  assign _zz_7543 = ($signed(twiddle_factor_table_1_real) + $signed(twiddle_factor_table_1_imag));
  assign _zz_7544 = fixTo_270_dout;
  assign _zz_7545 = ($signed(_zz_366) - $signed(_zz_365));
  assign _zz_7546 = ($signed(_zz_365) + $signed(_zz_366));
  assign _zz_7547 = _zz_7548[15 : 0];
  assign _zz_7548 = fixTo_272_dout;
  assign _zz_7549 = _zz_7550[15 : 0];
  assign _zz_7550 = fixTo_271_dout;
  assign _zz_7551 = _zz_7552;
  assign _zz_7552 = ($signed(_zz_7553) >>> _zz_2246);
  assign _zz_7553 = _zz_7554;
  assign _zz_7554 = ($signed(_zz_361) - $signed(_zz_2243));
  assign _zz_7555 = _zz_7556;
  assign _zz_7556 = ($signed(_zz_7557) >>> _zz_2246);
  assign _zz_7557 = _zz_7558;
  assign _zz_7558 = ($signed(_zz_362) - $signed(_zz_2244));
  assign _zz_7559 = _zz_7560;
  assign _zz_7560 = ($signed(_zz_7561) >>> _zz_2247);
  assign _zz_7561 = _zz_7562;
  assign _zz_7562 = ($signed(_zz_361) + $signed(_zz_2243));
  assign _zz_7563 = _zz_7564;
  assign _zz_7564 = ($signed(_zz_7565) >>> _zz_2247);
  assign _zz_7565 = _zz_7566;
  assign _zz_7566 = ($signed(_zz_362) + $signed(_zz_2244));
  assign _zz_7567 = ($signed(twiddle_factor_table_2_real) + $signed(twiddle_factor_table_2_imag));
  assign _zz_7568 = fixTo_273_dout;
  assign _zz_7569 = ($signed(_zz_368) - $signed(_zz_367));
  assign _zz_7570 = ($signed(_zz_367) + $signed(_zz_368));
  assign _zz_7571 = _zz_7572[15 : 0];
  assign _zz_7572 = fixTo_275_dout;
  assign _zz_7573 = _zz_7574[15 : 0];
  assign _zz_7574 = fixTo_274_dout;
  assign _zz_7575 = _zz_7576;
  assign _zz_7576 = ($signed(_zz_7577) >>> _zz_2251);
  assign _zz_7577 = _zz_7578;
  assign _zz_7578 = ($signed(_zz_363) - $signed(_zz_2248));
  assign _zz_7579 = _zz_7580;
  assign _zz_7580 = ($signed(_zz_7581) >>> _zz_2251);
  assign _zz_7581 = _zz_7582;
  assign _zz_7582 = ($signed(_zz_364) - $signed(_zz_2249));
  assign _zz_7583 = _zz_7584;
  assign _zz_7584 = ($signed(_zz_7585) >>> _zz_2252);
  assign _zz_7585 = _zz_7586;
  assign _zz_7586 = ($signed(_zz_363) + $signed(_zz_2248));
  assign _zz_7587 = _zz_7588;
  assign _zz_7588 = ($signed(_zz_7589) >>> _zz_2252);
  assign _zz_7589 = _zz_7590;
  assign _zz_7590 = ($signed(_zz_364) + $signed(_zz_2249));
  assign _zz_7591 = ($signed(twiddle_factor_table_1_real) + $signed(twiddle_factor_table_1_imag));
  assign _zz_7592 = fixTo_276_dout;
  assign _zz_7593 = ($signed(_zz_374) - $signed(_zz_373));
  assign _zz_7594 = ($signed(_zz_373) + $signed(_zz_374));
  assign _zz_7595 = _zz_7596[15 : 0];
  assign _zz_7596 = fixTo_278_dout;
  assign _zz_7597 = _zz_7598[15 : 0];
  assign _zz_7598 = fixTo_277_dout;
  assign _zz_7599 = _zz_7600;
  assign _zz_7600 = ($signed(_zz_7601) >>> _zz_2256);
  assign _zz_7601 = _zz_7602;
  assign _zz_7602 = ($signed(_zz_369) - $signed(_zz_2253));
  assign _zz_7603 = _zz_7604;
  assign _zz_7604 = ($signed(_zz_7605) >>> _zz_2256);
  assign _zz_7605 = _zz_7606;
  assign _zz_7606 = ($signed(_zz_370) - $signed(_zz_2254));
  assign _zz_7607 = _zz_7608;
  assign _zz_7608 = ($signed(_zz_7609) >>> _zz_2257);
  assign _zz_7609 = _zz_7610;
  assign _zz_7610 = ($signed(_zz_369) + $signed(_zz_2253));
  assign _zz_7611 = _zz_7612;
  assign _zz_7612 = ($signed(_zz_7613) >>> _zz_2257);
  assign _zz_7613 = _zz_7614;
  assign _zz_7614 = ($signed(_zz_370) + $signed(_zz_2254));
  assign _zz_7615 = ($signed(twiddle_factor_table_2_real) + $signed(twiddle_factor_table_2_imag));
  assign _zz_7616 = fixTo_279_dout;
  assign _zz_7617 = ($signed(_zz_376) - $signed(_zz_375));
  assign _zz_7618 = ($signed(_zz_375) + $signed(_zz_376));
  assign _zz_7619 = _zz_7620[15 : 0];
  assign _zz_7620 = fixTo_281_dout;
  assign _zz_7621 = _zz_7622[15 : 0];
  assign _zz_7622 = fixTo_280_dout;
  assign _zz_7623 = _zz_7624;
  assign _zz_7624 = ($signed(_zz_7625) >>> _zz_2261);
  assign _zz_7625 = _zz_7626;
  assign _zz_7626 = ($signed(_zz_371) - $signed(_zz_2258));
  assign _zz_7627 = _zz_7628;
  assign _zz_7628 = ($signed(_zz_7629) >>> _zz_2261);
  assign _zz_7629 = _zz_7630;
  assign _zz_7630 = ($signed(_zz_372) - $signed(_zz_2259));
  assign _zz_7631 = _zz_7632;
  assign _zz_7632 = ($signed(_zz_7633) >>> _zz_2262);
  assign _zz_7633 = _zz_7634;
  assign _zz_7634 = ($signed(_zz_371) + $signed(_zz_2258));
  assign _zz_7635 = _zz_7636;
  assign _zz_7636 = ($signed(_zz_7637) >>> _zz_2262);
  assign _zz_7637 = _zz_7638;
  assign _zz_7638 = ($signed(_zz_372) + $signed(_zz_2259));
  assign _zz_7639 = ($signed(twiddle_factor_table_1_real) + $signed(twiddle_factor_table_1_imag));
  assign _zz_7640 = fixTo_282_dout;
  assign _zz_7641 = ($signed(_zz_382) - $signed(_zz_381));
  assign _zz_7642 = ($signed(_zz_381) + $signed(_zz_382));
  assign _zz_7643 = _zz_7644[15 : 0];
  assign _zz_7644 = fixTo_284_dout;
  assign _zz_7645 = _zz_7646[15 : 0];
  assign _zz_7646 = fixTo_283_dout;
  assign _zz_7647 = _zz_7648;
  assign _zz_7648 = ($signed(_zz_7649) >>> _zz_2266);
  assign _zz_7649 = _zz_7650;
  assign _zz_7650 = ($signed(_zz_377) - $signed(_zz_2263));
  assign _zz_7651 = _zz_7652;
  assign _zz_7652 = ($signed(_zz_7653) >>> _zz_2266);
  assign _zz_7653 = _zz_7654;
  assign _zz_7654 = ($signed(_zz_378) - $signed(_zz_2264));
  assign _zz_7655 = _zz_7656;
  assign _zz_7656 = ($signed(_zz_7657) >>> _zz_2267);
  assign _zz_7657 = _zz_7658;
  assign _zz_7658 = ($signed(_zz_377) + $signed(_zz_2263));
  assign _zz_7659 = _zz_7660;
  assign _zz_7660 = ($signed(_zz_7661) >>> _zz_2267);
  assign _zz_7661 = _zz_7662;
  assign _zz_7662 = ($signed(_zz_378) + $signed(_zz_2264));
  assign _zz_7663 = ($signed(twiddle_factor_table_2_real) + $signed(twiddle_factor_table_2_imag));
  assign _zz_7664 = fixTo_285_dout;
  assign _zz_7665 = ($signed(_zz_384) - $signed(_zz_383));
  assign _zz_7666 = ($signed(_zz_383) + $signed(_zz_384));
  assign _zz_7667 = _zz_7668[15 : 0];
  assign _zz_7668 = fixTo_287_dout;
  assign _zz_7669 = _zz_7670[15 : 0];
  assign _zz_7670 = fixTo_286_dout;
  assign _zz_7671 = _zz_7672;
  assign _zz_7672 = ($signed(_zz_7673) >>> _zz_2271);
  assign _zz_7673 = _zz_7674;
  assign _zz_7674 = ($signed(_zz_379) - $signed(_zz_2268));
  assign _zz_7675 = _zz_7676;
  assign _zz_7676 = ($signed(_zz_7677) >>> _zz_2271);
  assign _zz_7677 = _zz_7678;
  assign _zz_7678 = ($signed(_zz_380) - $signed(_zz_2269));
  assign _zz_7679 = _zz_7680;
  assign _zz_7680 = ($signed(_zz_7681) >>> _zz_2272);
  assign _zz_7681 = _zz_7682;
  assign _zz_7682 = ($signed(_zz_379) + $signed(_zz_2268));
  assign _zz_7683 = _zz_7684;
  assign _zz_7684 = ($signed(_zz_7685) >>> _zz_2272);
  assign _zz_7685 = _zz_7686;
  assign _zz_7686 = ($signed(_zz_380) + $signed(_zz_2269));
  assign _zz_7687 = ($signed(twiddle_factor_table_1_real) + $signed(twiddle_factor_table_1_imag));
  assign _zz_7688 = fixTo_288_dout;
  assign _zz_7689 = ($signed(_zz_390) - $signed(_zz_389));
  assign _zz_7690 = ($signed(_zz_389) + $signed(_zz_390));
  assign _zz_7691 = _zz_7692[15 : 0];
  assign _zz_7692 = fixTo_290_dout;
  assign _zz_7693 = _zz_7694[15 : 0];
  assign _zz_7694 = fixTo_289_dout;
  assign _zz_7695 = _zz_7696;
  assign _zz_7696 = ($signed(_zz_7697) >>> _zz_2276);
  assign _zz_7697 = _zz_7698;
  assign _zz_7698 = ($signed(_zz_385) - $signed(_zz_2273));
  assign _zz_7699 = _zz_7700;
  assign _zz_7700 = ($signed(_zz_7701) >>> _zz_2276);
  assign _zz_7701 = _zz_7702;
  assign _zz_7702 = ($signed(_zz_386) - $signed(_zz_2274));
  assign _zz_7703 = _zz_7704;
  assign _zz_7704 = ($signed(_zz_7705) >>> _zz_2277);
  assign _zz_7705 = _zz_7706;
  assign _zz_7706 = ($signed(_zz_385) + $signed(_zz_2273));
  assign _zz_7707 = _zz_7708;
  assign _zz_7708 = ($signed(_zz_7709) >>> _zz_2277);
  assign _zz_7709 = _zz_7710;
  assign _zz_7710 = ($signed(_zz_386) + $signed(_zz_2274));
  assign _zz_7711 = ($signed(twiddle_factor_table_2_real) + $signed(twiddle_factor_table_2_imag));
  assign _zz_7712 = fixTo_291_dout;
  assign _zz_7713 = ($signed(_zz_392) - $signed(_zz_391));
  assign _zz_7714 = ($signed(_zz_391) + $signed(_zz_392));
  assign _zz_7715 = _zz_7716[15 : 0];
  assign _zz_7716 = fixTo_293_dout;
  assign _zz_7717 = _zz_7718[15 : 0];
  assign _zz_7718 = fixTo_292_dout;
  assign _zz_7719 = _zz_7720;
  assign _zz_7720 = ($signed(_zz_7721) >>> _zz_2281);
  assign _zz_7721 = _zz_7722;
  assign _zz_7722 = ($signed(_zz_387) - $signed(_zz_2278));
  assign _zz_7723 = _zz_7724;
  assign _zz_7724 = ($signed(_zz_7725) >>> _zz_2281);
  assign _zz_7725 = _zz_7726;
  assign _zz_7726 = ($signed(_zz_388) - $signed(_zz_2279));
  assign _zz_7727 = _zz_7728;
  assign _zz_7728 = ($signed(_zz_7729) >>> _zz_2282);
  assign _zz_7729 = _zz_7730;
  assign _zz_7730 = ($signed(_zz_387) + $signed(_zz_2278));
  assign _zz_7731 = _zz_7732;
  assign _zz_7732 = ($signed(_zz_7733) >>> _zz_2282);
  assign _zz_7733 = _zz_7734;
  assign _zz_7734 = ($signed(_zz_388) + $signed(_zz_2279));
  assign _zz_7735 = ($signed(twiddle_factor_table_1_real) + $signed(twiddle_factor_table_1_imag));
  assign _zz_7736 = fixTo_294_dout;
  assign _zz_7737 = ($signed(_zz_398) - $signed(_zz_397));
  assign _zz_7738 = ($signed(_zz_397) + $signed(_zz_398));
  assign _zz_7739 = _zz_7740[15 : 0];
  assign _zz_7740 = fixTo_296_dout;
  assign _zz_7741 = _zz_7742[15 : 0];
  assign _zz_7742 = fixTo_295_dout;
  assign _zz_7743 = _zz_7744;
  assign _zz_7744 = ($signed(_zz_7745) >>> _zz_2286);
  assign _zz_7745 = _zz_7746;
  assign _zz_7746 = ($signed(_zz_393) - $signed(_zz_2283));
  assign _zz_7747 = _zz_7748;
  assign _zz_7748 = ($signed(_zz_7749) >>> _zz_2286);
  assign _zz_7749 = _zz_7750;
  assign _zz_7750 = ($signed(_zz_394) - $signed(_zz_2284));
  assign _zz_7751 = _zz_7752;
  assign _zz_7752 = ($signed(_zz_7753) >>> _zz_2287);
  assign _zz_7753 = _zz_7754;
  assign _zz_7754 = ($signed(_zz_393) + $signed(_zz_2283));
  assign _zz_7755 = _zz_7756;
  assign _zz_7756 = ($signed(_zz_7757) >>> _zz_2287);
  assign _zz_7757 = _zz_7758;
  assign _zz_7758 = ($signed(_zz_394) + $signed(_zz_2284));
  assign _zz_7759 = ($signed(twiddle_factor_table_2_real) + $signed(twiddle_factor_table_2_imag));
  assign _zz_7760 = fixTo_297_dout;
  assign _zz_7761 = ($signed(_zz_400) - $signed(_zz_399));
  assign _zz_7762 = ($signed(_zz_399) + $signed(_zz_400));
  assign _zz_7763 = _zz_7764[15 : 0];
  assign _zz_7764 = fixTo_299_dout;
  assign _zz_7765 = _zz_7766[15 : 0];
  assign _zz_7766 = fixTo_298_dout;
  assign _zz_7767 = _zz_7768;
  assign _zz_7768 = ($signed(_zz_7769) >>> _zz_2291);
  assign _zz_7769 = _zz_7770;
  assign _zz_7770 = ($signed(_zz_395) - $signed(_zz_2288));
  assign _zz_7771 = _zz_7772;
  assign _zz_7772 = ($signed(_zz_7773) >>> _zz_2291);
  assign _zz_7773 = _zz_7774;
  assign _zz_7774 = ($signed(_zz_396) - $signed(_zz_2289));
  assign _zz_7775 = _zz_7776;
  assign _zz_7776 = ($signed(_zz_7777) >>> _zz_2292);
  assign _zz_7777 = _zz_7778;
  assign _zz_7778 = ($signed(_zz_395) + $signed(_zz_2288));
  assign _zz_7779 = _zz_7780;
  assign _zz_7780 = ($signed(_zz_7781) >>> _zz_2292);
  assign _zz_7781 = _zz_7782;
  assign _zz_7782 = ($signed(_zz_396) + $signed(_zz_2289));
  assign _zz_7783 = ($signed(twiddle_factor_table_1_real) + $signed(twiddle_factor_table_1_imag));
  assign _zz_7784 = fixTo_300_dout;
  assign _zz_7785 = ($signed(_zz_406) - $signed(_zz_405));
  assign _zz_7786 = ($signed(_zz_405) + $signed(_zz_406));
  assign _zz_7787 = _zz_7788[15 : 0];
  assign _zz_7788 = fixTo_302_dout;
  assign _zz_7789 = _zz_7790[15 : 0];
  assign _zz_7790 = fixTo_301_dout;
  assign _zz_7791 = _zz_7792;
  assign _zz_7792 = ($signed(_zz_7793) >>> _zz_2296);
  assign _zz_7793 = _zz_7794;
  assign _zz_7794 = ($signed(_zz_401) - $signed(_zz_2293));
  assign _zz_7795 = _zz_7796;
  assign _zz_7796 = ($signed(_zz_7797) >>> _zz_2296);
  assign _zz_7797 = _zz_7798;
  assign _zz_7798 = ($signed(_zz_402) - $signed(_zz_2294));
  assign _zz_7799 = _zz_7800;
  assign _zz_7800 = ($signed(_zz_7801) >>> _zz_2297);
  assign _zz_7801 = _zz_7802;
  assign _zz_7802 = ($signed(_zz_401) + $signed(_zz_2293));
  assign _zz_7803 = _zz_7804;
  assign _zz_7804 = ($signed(_zz_7805) >>> _zz_2297);
  assign _zz_7805 = _zz_7806;
  assign _zz_7806 = ($signed(_zz_402) + $signed(_zz_2294));
  assign _zz_7807 = ($signed(twiddle_factor_table_2_real) + $signed(twiddle_factor_table_2_imag));
  assign _zz_7808 = fixTo_303_dout;
  assign _zz_7809 = ($signed(_zz_408) - $signed(_zz_407));
  assign _zz_7810 = ($signed(_zz_407) + $signed(_zz_408));
  assign _zz_7811 = _zz_7812[15 : 0];
  assign _zz_7812 = fixTo_305_dout;
  assign _zz_7813 = _zz_7814[15 : 0];
  assign _zz_7814 = fixTo_304_dout;
  assign _zz_7815 = _zz_7816;
  assign _zz_7816 = ($signed(_zz_7817) >>> _zz_2301);
  assign _zz_7817 = _zz_7818;
  assign _zz_7818 = ($signed(_zz_403) - $signed(_zz_2298));
  assign _zz_7819 = _zz_7820;
  assign _zz_7820 = ($signed(_zz_7821) >>> _zz_2301);
  assign _zz_7821 = _zz_7822;
  assign _zz_7822 = ($signed(_zz_404) - $signed(_zz_2299));
  assign _zz_7823 = _zz_7824;
  assign _zz_7824 = ($signed(_zz_7825) >>> _zz_2302);
  assign _zz_7825 = _zz_7826;
  assign _zz_7826 = ($signed(_zz_403) + $signed(_zz_2298));
  assign _zz_7827 = _zz_7828;
  assign _zz_7828 = ($signed(_zz_7829) >>> _zz_2302);
  assign _zz_7829 = _zz_7830;
  assign _zz_7830 = ($signed(_zz_404) + $signed(_zz_2299));
  assign _zz_7831 = ($signed(twiddle_factor_table_1_real) + $signed(twiddle_factor_table_1_imag));
  assign _zz_7832 = fixTo_306_dout;
  assign _zz_7833 = ($signed(_zz_414) - $signed(_zz_413));
  assign _zz_7834 = ($signed(_zz_413) + $signed(_zz_414));
  assign _zz_7835 = _zz_7836[15 : 0];
  assign _zz_7836 = fixTo_308_dout;
  assign _zz_7837 = _zz_7838[15 : 0];
  assign _zz_7838 = fixTo_307_dout;
  assign _zz_7839 = _zz_7840;
  assign _zz_7840 = ($signed(_zz_7841) >>> _zz_2306);
  assign _zz_7841 = _zz_7842;
  assign _zz_7842 = ($signed(_zz_409) - $signed(_zz_2303));
  assign _zz_7843 = _zz_7844;
  assign _zz_7844 = ($signed(_zz_7845) >>> _zz_2306);
  assign _zz_7845 = _zz_7846;
  assign _zz_7846 = ($signed(_zz_410) - $signed(_zz_2304));
  assign _zz_7847 = _zz_7848;
  assign _zz_7848 = ($signed(_zz_7849) >>> _zz_2307);
  assign _zz_7849 = _zz_7850;
  assign _zz_7850 = ($signed(_zz_409) + $signed(_zz_2303));
  assign _zz_7851 = _zz_7852;
  assign _zz_7852 = ($signed(_zz_7853) >>> _zz_2307);
  assign _zz_7853 = _zz_7854;
  assign _zz_7854 = ($signed(_zz_410) + $signed(_zz_2304));
  assign _zz_7855 = ($signed(twiddle_factor_table_2_real) + $signed(twiddle_factor_table_2_imag));
  assign _zz_7856 = fixTo_309_dout;
  assign _zz_7857 = ($signed(_zz_416) - $signed(_zz_415));
  assign _zz_7858 = ($signed(_zz_415) + $signed(_zz_416));
  assign _zz_7859 = _zz_7860[15 : 0];
  assign _zz_7860 = fixTo_311_dout;
  assign _zz_7861 = _zz_7862[15 : 0];
  assign _zz_7862 = fixTo_310_dout;
  assign _zz_7863 = _zz_7864;
  assign _zz_7864 = ($signed(_zz_7865) >>> _zz_2311);
  assign _zz_7865 = _zz_7866;
  assign _zz_7866 = ($signed(_zz_411) - $signed(_zz_2308));
  assign _zz_7867 = _zz_7868;
  assign _zz_7868 = ($signed(_zz_7869) >>> _zz_2311);
  assign _zz_7869 = _zz_7870;
  assign _zz_7870 = ($signed(_zz_412) - $signed(_zz_2309));
  assign _zz_7871 = _zz_7872;
  assign _zz_7872 = ($signed(_zz_7873) >>> _zz_2312);
  assign _zz_7873 = _zz_7874;
  assign _zz_7874 = ($signed(_zz_411) + $signed(_zz_2308));
  assign _zz_7875 = _zz_7876;
  assign _zz_7876 = ($signed(_zz_7877) >>> _zz_2312);
  assign _zz_7877 = _zz_7878;
  assign _zz_7878 = ($signed(_zz_412) + $signed(_zz_2309));
  assign _zz_7879 = ($signed(twiddle_factor_table_1_real) + $signed(twiddle_factor_table_1_imag));
  assign _zz_7880 = fixTo_312_dout;
  assign _zz_7881 = ($signed(_zz_422) - $signed(_zz_421));
  assign _zz_7882 = ($signed(_zz_421) + $signed(_zz_422));
  assign _zz_7883 = _zz_7884[15 : 0];
  assign _zz_7884 = fixTo_314_dout;
  assign _zz_7885 = _zz_7886[15 : 0];
  assign _zz_7886 = fixTo_313_dout;
  assign _zz_7887 = _zz_7888;
  assign _zz_7888 = ($signed(_zz_7889) >>> _zz_2316);
  assign _zz_7889 = _zz_7890;
  assign _zz_7890 = ($signed(_zz_417) - $signed(_zz_2313));
  assign _zz_7891 = _zz_7892;
  assign _zz_7892 = ($signed(_zz_7893) >>> _zz_2316);
  assign _zz_7893 = _zz_7894;
  assign _zz_7894 = ($signed(_zz_418) - $signed(_zz_2314));
  assign _zz_7895 = _zz_7896;
  assign _zz_7896 = ($signed(_zz_7897) >>> _zz_2317);
  assign _zz_7897 = _zz_7898;
  assign _zz_7898 = ($signed(_zz_417) + $signed(_zz_2313));
  assign _zz_7899 = _zz_7900;
  assign _zz_7900 = ($signed(_zz_7901) >>> _zz_2317);
  assign _zz_7901 = _zz_7902;
  assign _zz_7902 = ($signed(_zz_418) + $signed(_zz_2314));
  assign _zz_7903 = ($signed(twiddle_factor_table_2_real) + $signed(twiddle_factor_table_2_imag));
  assign _zz_7904 = fixTo_315_dout;
  assign _zz_7905 = ($signed(_zz_424) - $signed(_zz_423));
  assign _zz_7906 = ($signed(_zz_423) + $signed(_zz_424));
  assign _zz_7907 = _zz_7908[15 : 0];
  assign _zz_7908 = fixTo_317_dout;
  assign _zz_7909 = _zz_7910[15 : 0];
  assign _zz_7910 = fixTo_316_dout;
  assign _zz_7911 = _zz_7912;
  assign _zz_7912 = ($signed(_zz_7913) >>> _zz_2321);
  assign _zz_7913 = _zz_7914;
  assign _zz_7914 = ($signed(_zz_419) - $signed(_zz_2318));
  assign _zz_7915 = _zz_7916;
  assign _zz_7916 = ($signed(_zz_7917) >>> _zz_2321);
  assign _zz_7917 = _zz_7918;
  assign _zz_7918 = ($signed(_zz_420) - $signed(_zz_2319));
  assign _zz_7919 = _zz_7920;
  assign _zz_7920 = ($signed(_zz_7921) >>> _zz_2322);
  assign _zz_7921 = _zz_7922;
  assign _zz_7922 = ($signed(_zz_419) + $signed(_zz_2318));
  assign _zz_7923 = _zz_7924;
  assign _zz_7924 = ($signed(_zz_7925) >>> _zz_2322);
  assign _zz_7925 = _zz_7926;
  assign _zz_7926 = ($signed(_zz_420) + $signed(_zz_2319));
  assign _zz_7927 = ($signed(twiddle_factor_table_1_real) + $signed(twiddle_factor_table_1_imag));
  assign _zz_7928 = fixTo_318_dout;
  assign _zz_7929 = ($signed(_zz_430) - $signed(_zz_429));
  assign _zz_7930 = ($signed(_zz_429) + $signed(_zz_430));
  assign _zz_7931 = _zz_7932[15 : 0];
  assign _zz_7932 = fixTo_320_dout;
  assign _zz_7933 = _zz_7934[15 : 0];
  assign _zz_7934 = fixTo_319_dout;
  assign _zz_7935 = _zz_7936;
  assign _zz_7936 = ($signed(_zz_7937) >>> _zz_2326);
  assign _zz_7937 = _zz_7938;
  assign _zz_7938 = ($signed(_zz_425) - $signed(_zz_2323));
  assign _zz_7939 = _zz_7940;
  assign _zz_7940 = ($signed(_zz_7941) >>> _zz_2326);
  assign _zz_7941 = _zz_7942;
  assign _zz_7942 = ($signed(_zz_426) - $signed(_zz_2324));
  assign _zz_7943 = _zz_7944;
  assign _zz_7944 = ($signed(_zz_7945) >>> _zz_2327);
  assign _zz_7945 = _zz_7946;
  assign _zz_7946 = ($signed(_zz_425) + $signed(_zz_2323));
  assign _zz_7947 = _zz_7948;
  assign _zz_7948 = ($signed(_zz_7949) >>> _zz_2327);
  assign _zz_7949 = _zz_7950;
  assign _zz_7950 = ($signed(_zz_426) + $signed(_zz_2324));
  assign _zz_7951 = ($signed(twiddle_factor_table_2_real) + $signed(twiddle_factor_table_2_imag));
  assign _zz_7952 = fixTo_321_dout;
  assign _zz_7953 = ($signed(_zz_432) - $signed(_zz_431));
  assign _zz_7954 = ($signed(_zz_431) + $signed(_zz_432));
  assign _zz_7955 = _zz_7956[15 : 0];
  assign _zz_7956 = fixTo_323_dout;
  assign _zz_7957 = _zz_7958[15 : 0];
  assign _zz_7958 = fixTo_322_dout;
  assign _zz_7959 = _zz_7960;
  assign _zz_7960 = ($signed(_zz_7961) >>> _zz_2331);
  assign _zz_7961 = _zz_7962;
  assign _zz_7962 = ($signed(_zz_427) - $signed(_zz_2328));
  assign _zz_7963 = _zz_7964;
  assign _zz_7964 = ($signed(_zz_7965) >>> _zz_2331);
  assign _zz_7965 = _zz_7966;
  assign _zz_7966 = ($signed(_zz_428) - $signed(_zz_2329));
  assign _zz_7967 = _zz_7968;
  assign _zz_7968 = ($signed(_zz_7969) >>> _zz_2332);
  assign _zz_7969 = _zz_7970;
  assign _zz_7970 = ($signed(_zz_427) + $signed(_zz_2328));
  assign _zz_7971 = _zz_7972;
  assign _zz_7972 = ($signed(_zz_7973) >>> _zz_2332);
  assign _zz_7973 = _zz_7974;
  assign _zz_7974 = ($signed(_zz_428) + $signed(_zz_2329));
  assign _zz_7975 = ($signed(twiddle_factor_table_1_real) + $signed(twiddle_factor_table_1_imag));
  assign _zz_7976 = fixTo_324_dout;
  assign _zz_7977 = ($signed(_zz_438) - $signed(_zz_437));
  assign _zz_7978 = ($signed(_zz_437) + $signed(_zz_438));
  assign _zz_7979 = _zz_7980[15 : 0];
  assign _zz_7980 = fixTo_326_dout;
  assign _zz_7981 = _zz_7982[15 : 0];
  assign _zz_7982 = fixTo_325_dout;
  assign _zz_7983 = _zz_7984;
  assign _zz_7984 = ($signed(_zz_7985) >>> _zz_2336);
  assign _zz_7985 = _zz_7986;
  assign _zz_7986 = ($signed(_zz_433) - $signed(_zz_2333));
  assign _zz_7987 = _zz_7988;
  assign _zz_7988 = ($signed(_zz_7989) >>> _zz_2336);
  assign _zz_7989 = _zz_7990;
  assign _zz_7990 = ($signed(_zz_434) - $signed(_zz_2334));
  assign _zz_7991 = _zz_7992;
  assign _zz_7992 = ($signed(_zz_7993) >>> _zz_2337);
  assign _zz_7993 = _zz_7994;
  assign _zz_7994 = ($signed(_zz_433) + $signed(_zz_2333));
  assign _zz_7995 = _zz_7996;
  assign _zz_7996 = ($signed(_zz_7997) >>> _zz_2337);
  assign _zz_7997 = _zz_7998;
  assign _zz_7998 = ($signed(_zz_434) + $signed(_zz_2334));
  assign _zz_7999 = ($signed(twiddle_factor_table_2_real) + $signed(twiddle_factor_table_2_imag));
  assign _zz_8000 = fixTo_327_dout;
  assign _zz_8001 = ($signed(_zz_440) - $signed(_zz_439));
  assign _zz_8002 = ($signed(_zz_439) + $signed(_zz_440));
  assign _zz_8003 = _zz_8004[15 : 0];
  assign _zz_8004 = fixTo_329_dout;
  assign _zz_8005 = _zz_8006[15 : 0];
  assign _zz_8006 = fixTo_328_dout;
  assign _zz_8007 = _zz_8008;
  assign _zz_8008 = ($signed(_zz_8009) >>> _zz_2341);
  assign _zz_8009 = _zz_8010;
  assign _zz_8010 = ($signed(_zz_435) - $signed(_zz_2338));
  assign _zz_8011 = _zz_8012;
  assign _zz_8012 = ($signed(_zz_8013) >>> _zz_2341);
  assign _zz_8013 = _zz_8014;
  assign _zz_8014 = ($signed(_zz_436) - $signed(_zz_2339));
  assign _zz_8015 = _zz_8016;
  assign _zz_8016 = ($signed(_zz_8017) >>> _zz_2342);
  assign _zz_8017 = _zz_8018;
  assign _zz_8018 = ($signed(_zz_435) + $signed(_zz_2338));
  assign _zz_8019 = _zz_8020;
  assign _zz_8020 = ($signed(_zz_8021) >>> _zz_2342);
  assign _zz_8021 = _zz_8022;
  assign _zz_8022 = ($signed(_zz_436) + $signed(_zz_2339));
  assign _zz_8023 = ($signed(twiddle_factor_table_1_real) + $signed(twiddle_factor_table_1_imag));
  assign _zz_8024 = fixTo_330_dout;
  assign _zz_8025 = ($signed(_zz_446) - $signed(_zz_445));
  assign _zz_8026 = ($signed(_zz_445) + $signed(_zz_446));
  assign _zz_8027 = _zz_8028[15 : 0];
  assign _zz_8028 = fixTo_332_dout;
  assign _zz_8029 = _zz_8030[15 : 0];
  assign _zz_8030 = fixTo_331_dout;
  assign _zz_8031 = _zz_8032;
  assign _zz_8032 = ($signed(_zz_8033) >>> _zz_2346);
  assign _zz_8033 = _zz_8034;
  assign _zz_8034 = ($signed(_zz_441) - $signed(_zz_2343));
  assign _zz_8035 = _zz_8036;
  assign _zz_8036 = ($signed(_zz_8037) >>> _zz_2346);
  assign _zz_8037 = _zz_8038;
  assign _zz_8038 = ($signed(_zz_442) - $signed(_zz_2344));
  assign _zz_8039 = _zz_8040;
  assign _zz_8040 = ($signed(_zz_8041) >>> _zz_2347);
  assign _zz_8041 = _zz_8042;
  assign _zz_8042 = ($signed(_zz_441) + $signed(_zz_2343));
  assign _zz_8043 = _zz_8044;
  assign _zz_8044 = ($signed(_zz_8045) >>> _zz_2347);
  assign _zz_8045 = _zz_8046;
  assign _zz_8046 = ($signed(_zz_442) + $signed(_zz_2344));
  assign _zz_8047 = ($signed(twiddle_factor_table_2_real) + $signed(twiddle_factor_table_2_imag));
  assign _zz_8048 = fixTo_333_dout;
  assign _zz_8049 = ($signed(_zz_448) - $signed(_zz_447));
  assign _zz_8050 = ($signed(_zz_447) + $signed(_zz_448));
  assign _zz_8051 = _zz_8052[15 : 0];
  assign _zz_8052 = fixTo_335_dout;
  assign _zz_8053 = _zz_8054[15 : 0];
  assign _zz_8054 = fixTo_334_dout;
  assign _zz_8055 = _zz_8056;
  assign _zz_8056 = ($signed(_zz_8057) >>> _zz_2351);
  assign _zz_8057 = _zz_8058;
  assign _zz_8058 = ($signed(_zz_443) - $signed(_zz_2348));
  assign _zz_8059 = _zz_8060;
  assign _zz_8060 = ($signed(_zz_8061) >>> _zz_2351);
  assign _zz_8061 = _zz_8062;
  assign _zz_8062 = ($signed(_zz_444) - $signed(_zz_2349));
  assign _zz_8063 = _zz_8064;
  assign _zz_8064 = ($signed(_zz_8065) >>> _zz_2352);
  assign _zz_8065 = _zz_8066;
  assign _zz_8066 = ($signed(_zz_443) + $signed(_zz_2348));
  assign _zz_8067 = _zz_8068;
  assign _zz_8068 = ($signed(_zz_8069) >>> _zz_2352);
  assign _zz_8069 = _zz_8070;
  assign _zz_8070 = ($signed(_zz_444) + $signed(_zz_2349));
  assign _zz_8071 = ($signed(twiddle_factor_table_1_real) + $signed(twiddle_factor_table_1_imag));
  assign _zz_8072 = fixTo_336_dout;
  assign _zz_8073 = ($signed(_zz_454) - $signed(_zz_453));
  assign _zz_8074 = ($signed(_zz_453) + $signed(_zz_454));
  assign _zz_8075 = _zz_8076[15 : 0];
  assign _zz_8076 = fixTo_338_dout;
  assign _zz_8077 = _zz_8078[15 : 0];
  assign _zz_8078 = fixTo_337_dout;
  assign _zz_8079 = _zz_8080;
  assign _zz_8080 = ($signed(_zz_8081) >>> _zz_2356);
  assign _zz_8081 = _zz_8082;
  assign _zz_8082 = ($signed(_zz_449) - $signed(_zz_2353));
  assign _zz_8083 = _zz_8084;
  assign _zz_8084 = ($signed(_zz_8085) >>> _zz_2356);
  assign _zz_8085 = _zz_8086;
  assign _zz_8086 = ($signed(_zz_450) - $signed(_zz_2354));
  assign _zz_8087 = _zz_8088;
  assign _zz_8088 = ($signed(_zz_8089) >>> _zz_2357);
  assign _zz_8089 = _zz_8090;
  assign _zz_8090 = ($signed(_zz_449) + $signed(_zz_2353));
  assign _zz_8091 = _zz_8092;
  assign _zz_8092 = ($signed(_zz_8093) >>> _zz_2357);
  assign _zz_8093 = _zz_8094;
  assign _zz_8094 = ($signed(_zz_450) + $signed(_zz_2354));
  assign _zz_8095 = ($signed(twiddle_factor_table_2_real) + $signed(twiddle_factor_table_2_imag));
  assign _zz_8096 = fixTo_339_dout;
  assign _zz_8097 = ($signed(_zz_456) - $signed(_zz_455));
  assign _zz_8098 = ($signed(_zz_455) + $signed(_zz_456));
  assign _zz_8099 = _zz_8100[15 : 0];
  assign _zz_8100 = fixTo_341_dout;
  assign _zz_8101 = _zz_8102[15 : 0];
  assign _zz_8102 = fixTo_340_dout;
  assign _zz_8103 = _zz_8104;
  assign _zz_8104 = ($signed(_zz_8105) >>> _zz_2361);
  assign _zz_8105 = _zz_8106;
  assign _zz_8106 = ($signed(_zz_451) - $signed(_zz_2358));
  assign _zz_8107 = _zz_8108;
  assign _zz_8108 = ($signed(_zz_8109) >>> _zz_2361);
  assign _zz_8109 = _zz_8110;
  assign _zz_8110 = ($signed(_zz_452) - $signed(_zz_2359));
  assign _zz_8111 = _zz_8112;
  assign _zz_8112 = ($signed(_zz_8113) >>> _zz_2362);
  assign _zz_8113 = _zz_8114;
  assign _zz_8114 = ($signed(_zz_451) + $signed(_zz_2358));
  assign _zz_8115 = _zz_8116;
  assign _zz_8116 = ($signed(_zz_8117) >>> _zz_2362);
  assign _zz_8117 = _zz_8118;
  assign _zz_8118 = ($signed(_zz_452) + $signed(_zz_2359));
  assign _zz_8119 = ($signed(twiddle_factor_table_1_real) + $signed(twiddle_factor_table_1_imag));
  assign _zz_8120 = fixTo_342_dout;
  assign _zz_8121 = ($signed(_zz_462) - $signed(_zz_461));
  assign _zz_8122 = ($signed(_zz_461) + $signed(_zz_462));
  assign _zz_8123 = _zz_8124[15 : 0];
  assign _zz_8124 = fixTo_344_dout;
  assign _zz_8125 = _zz_8126[15 : 0];
  assign _zz_8126 = fixTo_343_dout;
  assign _zz_8127 = _zz_8128;
  assign _zz_8128 = ($signed(_zz_8129) >>> _zz_2366);
  assign _zz_8129 = _zz_8130;
  assign _zz_8130 = ($signed(_zz_457) - $signed(_zz_2363));
  assign _zz_8131 = _zz_8132;
  assign _zz_8132 = ($signed(_zz_8133) >>> _zz_2366);
  assign _zz_8133 = _zz_8134;
  assign _zz_8134 = ($signed(_zz_458) - $signed(_zz_2364));
  assign _zz_8135 = _zz_8136;
  assign _zz_8136 = ($signed(_zz_8137) >>> _zz_2367);
  assign _zz_8137 = _zz_8138;
  assign _zz_8138 = ($signed(_zz_457) + $signed(_zz_2363));
  assign _zz_8139 = _zz_8140;
  assign _zz_8140 = ($signed(_zz_8141) >>> _zz_2367);
  assign _zz_8141 = _zz_8142;
  assign _zz_8142 = ($signed(_zz_458) + $signed(_zz_2364));
  assign _zz_8143 = ($signed(twiddle_factor_table_2_real) + $signed(twiddle_factor_table_2_imag));
  assign _zz_8144 = fixTo_345_dout;
  assign _zz_8145 = ($signed(_zz_464) - $signed(_zz_463));
  assign _zz_8146 = ($signed(_zz_463) + $signed(_zz_464));
  assign _zz_8147 = _zz_8148[15 : 0];
  assign _zz_8148 = fixTo_347_dout;
  assign _zz_8149 = _zz_8150[15 : 0];
  assign _zz_8150 = fixTo_346_dout;
  assign _zz_8151 = _zz_8152;
  assign _zz_8152 = ($signed(_zz_8153) >>> _zz_2371);
  assign _zz_8153 = _zz_8154;
  assign _zz_8154 = ($signed(_zz_459) - $signed(_zz_2368));
  assign _zz_8155 = _zz_8156;
  assign _zz_8156 = ($signed(_zz_8157) >>> _zz_2371);
  assign _zz_8157 = _zz_8158;
  assign _zz_8158 = ($signed(_zz_460) - $signed(_zz_2369));
  assign _zz_8159 = _zz_8160;
  assign _zz_8160 = ($signed(_zz_8161) >>> _zz_2372);
  assign _zz_8161 = _zz_8162;
  assign _zz_8162 = ($signed(_zz_459) + $signed(_zz_2368));
  assign _zz_8163 = _zz_8164;
  assign _zz_8164 = ($signed(_zz_8165) >>> _zz_2372);
  assign _zz_8165 = _zz_8166;
  assign _zz_8166 = ($signed(_zz_460) + $signed(_zz_2369));
  assign _zz_8167 = ($signed(twiddle_factor_table_1_real) + $signed(twiddle_factor_table_1_imag));
  assign _zz_8168 = fixTo_348_dout;
  assign _zz_8169 = ($signed(_zz_470) - $signed(_zz_469));
  assign _zz_8170 = ($signed(_zz_469) + $signed(_zz_470));
  assign _zz_8171 = _zz_8172[15 : 0];
  assign _zz_8172 = fixTo_350_dout;
  assign _zz_8173 = _zz_8174[15 : 0];
  assign _zz_8174 = fixTo_349_dout;
  assign _zz_8175 = _zz_8176;
  assign _zz_8176 = ($signed(_zz_8177) >>> _zz_2376);
  assign _zz_8177 = _zz_8178;
  assign _zz_8178 = ($signed(_zz_465) - $signed(_zz_2373));
  assign _zz_8179 = _zz_8180;
  assign _zz_8180 = ($signed(_zz_8181) >>> _zz_2376);
  assign _zz_8181 = _zz_8182;
  assign _zz_8182 = ($signed(_zz_466) - $signed(_zz_2374));
  assign _zz_8183 = _zz_8184;
  assign _zz_8184 = ($signed(_zz_8185) >>> _zz_2377);
  assign _zz_8185 = _zz_8186;
  assign _zz_8186 = ($signed(_zz_465) + $signed(_zz_2373));
  assign _zz_8187 = _zz_8188;
  assign _zz_8188 = ($signed(_zz_8189) >>> _zz_2377);
  assign _zz_8189 = _zz_8190;
  assign _zz_8190 = ($signed(_zz_466) + $signed(_zz_2374));
  assign _zz_8191 = ($signed(twiddle_factor_table_2_real) + $signed(twiddle_factor_table_2_imag));
  assign _zz_8192 = fixTo_351_dout;
  assign _zz_8193 = ($signed(_zz_472) - $signed(_zz_471));
  assign _zz_8194 = ($signed(_zz_471) + $signed(_zz_472));
  assign _zz_8195 = _zz_8196[15 : 0];
  assign _zz_8196 = fixTo_353_dout;
  assign _zz_8197 = _zz_8198[15 : 0];
  assign _zz_8198 = fixTo_352_dout;
  assign _zz_8199 = _zz_8200;
  assign _zz_8200 = ($signed(_zz_8201) >>> _zz_2381);
  assign _zz_8201 = _zz_8202;
  assign _zz_8202 = ($signed(_zz_467) - $signed(_zz_2378));
  assign _zz_8203 = _zz_8204;
  assign _zz_8204 = ($signed(_zz_8205) >>> _zz_2381);
  assign _zz_8205 = _zz_8206;
  assign _zz_8206 = ($signed(_zz_468) - $signed(_zz_2379));
  assign _zz_8207 = _zz_8208;
  assign _zz_8208 = ($signed(_zz_8209) >>> _zz_2382);
  assign _zz_8209 = _zz_8210;
  assign _zz_8210 = ($signed(_zz_467) + $signed(_zz_2378));
  assign _zz_8211 = _zz_8212;
  assign _zz_8212 = ($signed(_zz_8213) >>> _zz_2382);
  assign _zz_8213 = _zz_8214;
  assign _zz_8214 = ($signed(_zz_468) + $signed(_zz_2379));
  assign _zz_8215 = ($signed(twiddle_factor_table_1_real) + $signed(twiddle_factor_table_1_imag));
  assign _zz_8216 = fixTo_354_dout;
  assign _zz_8217 = ($signed(_zz_478) - $signed(_zz_477));
  assign _zz_8218 = ($signed(_zz_477) + $signed(_zz_478));
  assign _zz_8219 = _zz_8220[15 : 0];
  assign _zz_8220 = fixTo_356_dout;
  assign _zz_8221 = _zz_8222[15 : 0];
  assign _zz_8222 = fixTo_355_dout;
  assign _zz_8223 = _zz_8224;
  assign _zz_8224 = ($signed(_zz_8225) >>> _zz_2386);
  assign _zz_8225 = _zz_8226;
  assign _zz_8226 = ($signed(_zz_473) - $signed(_zz_2383));
  assign _zz_8227 = _zz_8228;
  assign _zz_8228 = ($signed(_zz_8229) >>> _zz_2386);
  assign _zz_8229 = _zz_8230;
  assign _zz_8230 = ($signed(_zz_474) - $signed(_zz_2384));
  assign _zz_8231 = _zz_8232;
  assign _zz_8232 = ($signed(_zz_8233) >>> _zz_2387);
  assign _zz_8233 = _zz_8234;
  assign _zz_8234 = ($signed(_zz_473) + $signed(_zz_2383));
  assign _zz_8235 = _zz_8236;
  assign _zz_8236 = ($signed(_zz_8237) >>> _zz_2387);
  assign _zz_8237 = _zz_8238;
  assign _zz_8238 = ($signed(_zz_474) + $signed(_zz_2384));
  assign _zz_8239 = ($signed(twiddle_factor_table_2_real) + $signed(twiddle_factor_table_2_imag));
  assign _zz_8240 = fixTo_357_dout;
  assign _zz_8241 = ($signed(_zz_480) - $signed(_zz_479));
  assign _zz_8242 = ($signed(_zz_479) + $signed(_zz_480));
  assign _zz_8243 = _zz_8244[15 : 0];
  assign _zz_8244 = fixTo_359_dout;
  assign _zz_8245 = _zz_8246[15 : 0];
  assign _zz_8246 = fixTo_358_dout;
  assign _zz_8247 = _zz_8248;
  assign _zz_8248 = ($signed(_zz_8249) >>> _zz_2391);
  assign _zz_8249 = _zz_8250;
  assign _zz_8250 = ($signed(_zz_475) - $signed(_zz_2388));
  assign _zz_8251 = _zz_8252;
  assign _zz_8252 = ($signed(_zz_8253) >>> _zz_2391);
  assign _zz_8253 = _zz_8254;
  assign _zz_8254 = ($signed(_zz_476) - $signed(_zz_2389));
  assign _zz_8255 = _zz_8256;
  assign _zz_8256 = ($signed(_zz_8257) >>> _zz_2392);
  assign _zz_8257 = _zz_8258;
  assign _zz_8258 = ($signed(_zz_475) + $signed(_zz_2388));
  assign _zz_8259 = _zz_8260;
  assign _zz_8260 = ($signed(_zz_8261) >>> _zz_2392);
  assign _zz_8261 = _zz_8262;
  assign _zz_8262 = ($signed(_zz_476) + $signed(_zz_2389));
  assign _zz_8263 = ($signed(twiddle_factor_table_1_real) + $signed(twiddle_factor_table_1_imag));
  assign _zz_8264 = fixTo_360_dout;
  assign _zz_8265 = ($signed(_zz_486) - $signed(_zz_485));
  assign _zz_8266 = ($signed(_zz_485) + $signed(_zz_486));
  assign _zz_8267 = _zz_8268[15 : 0];
  assign _zz_8268 = fixTo_362_dout;
  assign _zz_8269 = _zz_8270[15 : 0];
  assign _zz_8270 = fixTo_361_dout;
  assign _zz_8271 = _zz_8272;
  assign _zz_8272 = ($signed(_zz_8273) >>> _zz_2396);
  assign _zz_8273 = _zz_8274;
  assign _zz_8274 = ($signed(_zz_481) - $signed(_zz_2393));
  assign _zz_8275 = _zz_8276;
  assign _zz_8276 = ($signed(_zz_8277) >>> _zz_2396);
  assign _zz_8277 = _zz_8278;
  assign _zz_8278 = ($signed(_zz_482) - $signed(_zz_2394));
  assign _zz_8279 = _zz_8280;
  assign _zz_8280 = ($signed(_zz_8281) >>> _zz_2397);
  assign _zz_8281 = _zz_8282;
  assign _zz_8282 = ($signed(_zz_481) + $signed(_zz_2393));
  assign _zz_8283 = _zz_8284;
  assign _zz_8284 = ($signed(_zz_8285) >>> _zz_2397);
  assign _zz_8285 = _zz_8286;
  assign _zz_8286 = ($signed(_zz_482) + $signed(_zz_2394));
  assign _zz_8287 = ($signed(twiddle_factor_table_2_real) + $signed(twiddle_factor_table_2_imag));
  assign _zz_8288 = fixTo_363_dout;
  assign _zz_8289 = ($signed(_zz_488) - $signed(_zz_487));
  assign _zz_8290 = ($signed(_zz_487) + $signed(_zz_488));
  assign _zz_8291 = _zz_8292[15 : 0];
  assign _zz_8292 = fixTo_365_dout;
  assign _zz_8293 = _zz_8294[15 : 0];
  assign _zz_8294 = fixTo_364_dout;
  assign _zz_8295 = _zz_8296;
  assign _zz_8296 = ($signed(_zz_8297) >>> _zz_2401);
  assign _zz_8297 = _zz_8298;
  assign _zz_8298 = ($signed(_zz_483) - $signed(_zz_2398));
  assign _zz_8299 = _zz_8300;
  assign _zz_8300 = ($signed(_zz_8301) >>> _zz_2401);
  assign _zz_8301 = _zz_8302;
  assign _zz_8302 = ($signed(_zz_484) - $signed(_zz_2399));
  assign _zz_8303 = _zz_8304;
  assign _zz_8304 = ($signed(_zz_8305) >>> _zz_2402);
  assign _zz_8305 = _zz_8306;
  assign _zz_8306 = ($signed(_zz_483) + $signed(_zz_2398));
  assign _zz_8307 = _zz_8308;
  assign _zz_8308 = ($signed(_zz_8309) >>> _zz_2402);
  assign _zz_8309 = _zz_8310;
  assign _zz_8310 = ($signed(_zz_484) + $signed(_zz_2399));
  assign _zz_8311 = ($signed(twiddle_factor_table_1_real) + $signed(twiddle_factor_table_1_imag));
  assign _zz_8312 = fixTo_366_dout;
  assign _zz_8313 = ($signed(_zz_494) - $signed(_zz_493));
  assign _zz_8314 = ($signed(_zz_493) + $signed(_zz_494));
  assign _zz_8315 = _zz_8316[15 : 0];
  assign _zz_8316 = fixTo_368_dout;
  assign _zz_8317 = _zz_8318[15 : 0];
  assign _zz_8318 = fixTo_367_dout;
  assign _zz_8319 = _zz_8320;
  assign _zz_8320 = ($signed(_zz_8321) >>> _zz_2406);
  assign _zz_8321 = _zz_8322;
  assign _zz_8322 = ($signed(_zz_489) - $signed(_zz_2403));
  assign _zz_8323 = _zz_8324;
  assign _zz_8324 = ($signed(_zz_8325) >>> _zz_2406);
  assign _zz_8325 = _zz_8326;
  assign _zz_8326 = ($signed(_zz_490) - $signed(_zz_2404));
  assign _zz_8327 = _zz_8328;
  assign _zz_8328 = ($signed(_zz_8329) >>> _zz_2407);
  assign _zz_8329 = _zz_8330;
  assign _zz_8330 = ($signed(_zz_489) + $signed(_zz_2403));
  assign _zz_8331 = _zz_8332;
  assign _zz_8332 = ($signed(_zz_8333) >>> _zz_2407);
  assign _zz_8333 = _zz_8334;
  assign _zz_8334 = ($signed(_zz_490) + $signed(_zz_2404));
  assign _zz_8335 = ($signed(twiddle_factor_table_2_real) + $signed(twiddle_factor_table_2_imag));
  assign _zz_8336 = fixTo_369_dout;
  assign _zz_8337 = ($signed(_zz_496) - $signed(_zz_495));
  assign _zz_8338 = ($signed(_zz_495) + $signed(_zz_496));
  assign _zz_8339 = _zz_8340[15 : 0];
  assign _zz_8340 = fixTo_371_dout;
  assign _zz_8341 = _zz_8342[15 : 0];
  assign _zz_8342 = fixTo_370_dout;
  assign _zz_8343 = _zz_8344;
  assign _zz_8344 = ($signed(_zz_8345) >>> _zz_2411);
  assign _zz_8345 = _zz_8346;
  assign _zz_8346 = ($signed(_zz_491) - $signed(_zz_2408));
  assign _zz_8347 = _zz_8348;
  assign _zz_8348 = ($signed(_zz_8349) >>> _zz_2411);
  assign _zz_8349 = _zz_8350;
  assign _zz_8350 = ($signed(_zz_492) - $signed(_zz_2409));
  assign _zz_8351 = _zz_8352;
  assign _zz_8352 = ($signed(_zz_8353) >>> _zz_2412);
  assign _zz_8353 = _zz_8354;
  assign _zz_8354 = ($signed(_zz_491) + $signed(_zz_2408));
  assign _zz_8355 = _zz_8356;
  assign _zz_8356 = ($signed(_zz_8357) >>> _zz_2412);
  assign _zz_8357 = _zz_8358;
  assign _zz_8358 = ($signed(_zz_492) + $signed(_zz_2409));
  assign _zz_8359 = ($signed(twiddle_factor_table_1_real) + $signed(twiddle_factor_table_1_imag));
  assign _zz_8360 = fixTo_372_dout;
  assign _zz_8361 = ($signed(_zz_502) - $signed(_zz_501));
  assign _zz_8362 = ($signed(_zz_501) + $signed(_zz_502));
  assign _zz_8363 = _zz_8364[15 : 0];
  assign _zz_8364 = fixTo_374_dout;
  assign _zz_8365 = _zz_8366[15 : 0];
  assign _zz_8366 = fixTo_373_dout;
  assign _zz_8367 = _zz_8368;
  assign _zz_8368 = ($signed(_zz_8369) >>> _zz_2416);
  assign _zz_8369 = _zz_8370;
  assign _zz_8370 = ($signed(_zz_497) - $signed(_zz_2413));
  assign _zz_8371 = _zz_8372;
  assign _zz_8372 = ($signed(_zz_8373) >>> _zz_2416);
  assign _zz_8373 = _zz_8374;
  assign _zz_8374 = ($signed(_zz_498) - $signed(_zz_2414));
  assign _zz_8375 = _zz_8376;
  assign _zz_8376 = ($signed(_zz_8377) >>> _zz_2417);
  assign _zz_8377 = _zz_8378;
  assign _zz_8378 = ($signed(_zz_497) + $signed(_zz_2413));
  assign _zz_8379 = _zz_8380;
  assign _zz_8380 = ($signed(_zz_8381) >>> _zz_2417);
  assign _zz_8381 = _zz_8382;
  assign _zz_8382 = ($signed(_zz_498) + $signed(_zz_2414));
  assign _zz_8383 = ($signed(twiddle_factor_table_2_real) + $signed(twiddle_factor_table_2_imag));
  assign _zz_8384 = fixTo_375_dout;
  assign _zz_8385 = ($signed(_zz_504) - $signed(_zz_503));
  assign _zz_8386 = ($signed(_zz_503) + $signed(_zz_504));
  assign _zz_8387 = _zz_8388[15 : 0];
  assign _zz_8388 = fixTo_377_dout;
  assign _zz_8389 = _zz_8390[15 : 0];
  assign _zz_8390 = fixTo_376_dout;
  assign _zz_8391 = _zz_8392;
  assign _zz_8392 = ($signed(_zz_8393) >>> _zz_2421);
  assign _zz_8393 = _zz_8394;
  assign _zz_8394 = ($signed(_zz_499) - $signed(_zz_2418));
  assign _zz_8395 = _zz_8396;
  assign _zz_8396 = ($signed(_zz_8397) >>> _zz_2421);
  assign _zz_8397 = _zz_8398;
  assign _zz_8398 = ($signed(_zz_500) - $signed(_zz_2419));
  assign _zz_8399 = _zz_8400;
  assign _zz_8400 = ($signed(_zz_8401) >>> _zz_2422);
  assign _zz_8401 = _zz_8402;
  assign _zz_8402 = ($signed(_zz_499) + $signed(_zz_2418));
  assign _zz_8403 = _zz_8404;
  assign _zz_8404 = ($signed(_zz_8405) >>> _zz_2422);
  assign _zz_8405 = _zz_8406;
  assign _zz_8406 = ($signed(_zz_500) + $signed(_zz_2419));
  assign _zz_8407 = ($signed(twiddle_factor_table_1_real) + $signed(twiddle_factor_table_1_imag));
  assign _zz_8408 = fixTo_378_dout;
  assign _zz_8409 = ($signed(_zz_510) - $signed(_zz_509));
  assign _zz_8410 = ($signed(_zz_509) + $signed(_zz_510));
  assign _zz_8411 = _zz_8412[15 : 0];
  assign _zz_8412 = fixTo_380_dout;
  assign _zz_8413 = _zz_8414[15 : 0];
  assign _zz_8414 = fixTo_379_dout;
  assign _zz_8415 = _zz_8416;
  assign _zz_8416 = ($signed(_zz_8417) >>> _zz_2426);
  assign _zz_8417 = _zz_8418;
  assign _zz_8418 = ($signed(_zz_505) - $signed(_zz_2423));
  assign _zz_8419 = _zz_8420;
  assign _zz_8420 = ($signed(_zz_8421) >>> _zz_2426);
  assign _zz_8421 = _zz_8422;
  assign _zz_8422 = ($signed(_zz_506) - $signed(_zz_2424));
  assign _zz_8423 = _zz_8424;
  assign _zz_8424 = ($signed(_zz_8425) >>> _zz_2427);
  assign _zz_8425 = _zz_8426;
  assign _zz_8426 = ($signed(_zz_505) + $signed(_zz_2423));
  assign _zz_8427 = _zz_8428;
  assign _zz_8428 = ($signed(_zz_8429) >>> _zz_2427);
  assign _zz_8429 = _zz_8430;
  assign _zz_8430 = ($signed(_zz_506) + $signed(_zz_2424));
  assign _zz_8431 = ($signed(twiddle_factor_table_2_real) + $signed(twiddle_factor_table_2_imag));
  assign _zz_8432 = fixTo_381_dout;
  assign _zz_8433 = ($signed(_zz_512) - $signed(_zz_511));
  assign _zz_8434 = ($signed(_zz_511) + $signed(_zz_512));
  assign _zz_8435 = _zz_8436[15 : 0];
  assign _zz_8436 = fixTo_383_dout;
  assign _zz_8437 = _zz_8438[15 : 0];
  assign _zz_8438 = fixTo_382_dout;
  assign _zz_8439 = _zz_8440;
  assign _zz_8440 = ($signed(_zz_8441) >>> _zz_2431);
  assign _zz_8441 = _zz_8442;
  assign _zz_8442 = ($signed(_zz_507) - $signed(_zz_2428));
  assign _zz_8443 = _zz_8444;
  assign _zz_8444 = ($signed(_zz_8445) >>> _zz_2431);
  assign _zz_8445 = _zz_8446;
  assign _zz_8446 = ($signed(_zz_508) - $signed(_zz_2429));
  assign _zz_8447 = _zz_8448;
  assign _zz_8448 = ($signed(_zz_8449) >>> _zz_2432);
  assign _zz_8449 = _zz_8450;
  assign _zz_8450 = ($signed(_zz_507) + $signed(_zz_2428));
  assign _zz_8451 = _zz_8452;
  assign _zz_8452 = ($signed(_zz_8453) >>> _zz_2432);
  assign _zz_8453 = _zz_8454;
  assign _zz_8454 = ($signed(_zz_508) + $signed(_zz_2429));
  assign _zz_8455 = ($signed(twiddle_factor_table_3_real) + $signed(twiddle_factor_table_3_imag));
  assign _zz_8456 = fixTo_384_dout;
  assign _zz_8457 = ($signed(_zz_522) - $signed(_zz_521));
  assign _zz_8458 = ($signed(_zz_521) + $signed(_zz_522));
  assign _zz_8459 = _zz_8460[15 : 0];
  assign _zz_8460 = fixTo_386_dout;
  assign _zz_8461 = _zz_8462[15 : 0];
  assign _zz_8462 = fixTo_385_dout;
  assign _zz_8463 = _zz_8464;
  assign _zz_8464 = ($signed(_zz_8465) >>> _zz_2436);
  assign _zz_8465 = _zz_8466;
  assign _zz_8466 = ($signed(_zz_513) - $signed(_zz_2433));
  assign _zz_8467 = _zz_8468;
  assign _zz_8468 = ($signed(_zz_8469) >>> _zz_2436);
  assign _zz_8469 = _zz_8470;
  assign _zz_8470 = ($signed(_zz_514) - $signed(_zz_2434));
  assign _zz_8471 = _zz_8472;
  assign _zz_8472 = ($signed(_zz_8473) >>> _zz_2437);
  assign _zz_8473 = _zz_8474;
  assign _zz_8474 = ($signed(_zz_513) + $signed(_zz_2433));
  assign _zz_8475 = _zz_8476;
  assign _zz_8476 = ($signed(_zz_8477) >>> _zz_2437);
  assign _zz_8477 = _zz_8478;
  assign _zz_8478 = ($signed(_zz_514) + $signed(_zz_2434));
  assign _zz_8479 = ($signed(twiddle_factor_table_4_real) + $signed(twiddle_factor_table_4_imag));
  assign _zz_8480 = fixTo_387_dout;
  assign _zz_8481 = ($signed(_zz_524) - $signed(_zz_523));
  assign _zz_8482 = ($signed(_zz_523) + $signed(_zz_524));
  assign _zz_8483 = _zz_8484[15 : 0];
  assign _zz_8484 = fixTo_389_dout;
  assign _zz_8485 = _zz_8486[15 : 0];
  assign _zz_8486 = fixTo_388_dout;
  assign _zz_8487 = _zz_8488;
  assign _zz_8488 = ($signed(_zz_8489) >>> _zz_2441);
  assign _zz_8489 = _zz_8490;
  assign _zz_8490 = ($signed(_zz_515) - $signed(_zz_2438));
  assign _zz_8491 = _zz_8492;
  assign _zz_8492 = ($signed(_zz_8493) >>> _zz_2441);
  assign _zz_8493 = _zz_8494;
  assign _zz_8494 = ($signed(_zz_516) - $signed(_zz_2439));
  assign _zz_8495 = _zz_8496;
  assign _zz_8496 = ($signed(_zz_8497) >>> _zz_2442);
  assign _zz_8497 = _zz_8498;
  assign _zz_8498 = ($signed(_zz_515) + $signed(_zz_2438));
  assign _zz_8499 = _zz_8500;
  assign _zz_8500 = ($signed(_zz_8501) >>> _zz_2442);
  assign _zz_8501 = _zz_8502;
  assign _zz_8502 = ($signed(_zz_516) + $signed(_zz_2439));
  assign _zz_8503 = ($signed(twiddle_factor_table_5_real) + $signed(twiddle_factor_table_5_imag));
  assign _zz_8504 = fixTo_390_dout;
  assign _zz_8505 = ($signed(_zz_526) - $signed(_zz_525));
  assign _zz_8506 = ($signed(_zz_525) + $signed(_zz_526));
  assign _zz_8507 = _zz_8508[15 : 0];
  assign _zz_8508 = fixTo_392_dout;
  assign _zz_8509 = _zz_8510[15 : 0];
  assign _zz_8510 = fixTo_391_dout;
  assign _zz_8511 = _zz_8512;
  assign _zz_8512 = ($signed(_zz_8513) >>> _zz_2446);
  assign _zz_8513 = _zz_8514;
  assign _zz_8514 = ($signed(_zz_517) - $signed(_zz_2443));
  assign _zz_8515 = _zz_8516;
  assign _zz_8516 = ($signed(_zz_8517) >>> _zz_2446);
  assign _zz_8517 = _zz_8518;
  assign _zz_8518 = ($signed(_zz_518) - $signed(_zz_2444));
  assign _zz_8519 = _zz_8520;
  assign _zz_8520 = ($signed(_zz_8521) >>> _zz_2447);
  assign _zz_8521 = _zz_8522;
  assign _zz_8522 = ($signed(_zz_517) + $signed(_zz_2443));
  assign _zz_8523 = _zz_8524;
  assign _zz_8524 = ($signed(_zz_8525) >>> _zz_2447);
  assign _zz_8525 = _zz_8526;
  assign _zz_8526 = ($signed(_zz_518) + $signed(_zz_2444));
  assign _zz_8527 = ($signed(twiddle_factor_table_6_real) + $signed(twiddle_factor_table_6_imag));
  assign _zz_8528 = fixTo_393_dout;
  assign _zz_8529 = ($signed(_zz_528) - $signed(_zz_527));
  assign _zz_8530 = ($signed(_zz_527) + $signed(_zz_528));
  assign _zz_8531 = _zz_8532[15 : 0];
  assign _zz_8532 = fixTo_395_dout;
  assign _zz_8533 = _zz_8534[15 : 0];
  assign _zz_8534 = fixTo_394_dout;
  assign _zz_8535 = _zz_8536;
  assign _zz_8536 = ($signed(_zz_8537) >>> _zz_2451);
  assign _zz_8537 = _zz_8538;
  assign _zz_8538 = ($signed(_zz_519) - $signed(_zz_2448));
  assign _zz_8539 = _zz_8540;
  assign _zz_8540 = ($signed(_zz_8541) >>> _zz_2451);
  assign _zz_8541 = _zz_8542;
  assign _zz_8542 = ($signed(_zz_520) - $signed(_zz_2449));
  assign _zz_8543 = _zz_8544;
  assign _zz_8544 = ($signed(_zz_8545) >>> _zz_2452);
  assign _zz_8545 = _zz_8546;
  assign _zz_8546 = ($signed(_zz_519) + $signed(_zz_2448));
  assign _zz_8547 = _zz_8548;
  assign _zz_8548 = ($signed(_zz_8549) >>> _zz_2452);
  assign _zz_8549 = _zz_8550;
  assign _zz_8550 = ($signed(_zz_520) + $signed(_zz_2449));
  assign _zz_8551 = ($signed(twiddle_factor_table_3_real) + $signed(twiddle_factor_table_3_imag));
  assign _zz_8552 = fixTo_396_dout;
  assign _zz_8553 = ($signed(_zz_538) - $signed(_zz_537));
  assign _zz_8554 = ($signed(_zz_537) + $signed(_zz_538));
  assign _zz_8555 = _zz_8556[15 : 0];
  assign _zz_8556 = fixTo_398_dout;
  assign _zz_8557 = _zz_8558[15 : 0];
  assign _zz_8558 = fixTo_397_dout;
  assign _zz_8559 = _zz_8560;
  assign _zz_8560 = ($signed(_zz_8561) >>> _zz_2456);
  assign _zz_8561 = _zz_8562;
  assign _zz_8562 = ($signed(_zz_529) - $signed(_zz_2453));
  assign _zz_8563 = _zz_8564;
  assign _zz_8564 = ($signed(_zz_8565) >>> _zz_2456);
  assign _zz_8565 = _zz_8566;
  assign _zz_8566 = ($signed(_zz_530) - $signed(_zz_2454));
  assign _zz_8567 = _zz_8568;
  assign _zz_8568 = ($signed(_zz_8569) >>> _zz_2457);
  assign _zz_8569 = _zz_8570;
  assign _zz_8570 = ($signed(_zz_529) + $signed(_zz_2453));
  assign _zz_8571 = _zz_8572;
  assign _zz_8572 = ($signed(_zz_8573) >>> _zz_2457);
  assign _zz_8573 = _zz_8574;
  assign _zz_8574 = ($signed(_zz_530) + $signed(_zz_2454));
  assign _zz_8575 = ($signed(twiddle_factor_table_4_real) + $signed(twiddle_factor_table_4_imag));
  assign _zz_8576 = fixTo_399_dout;
  assign _zz_8577 = ($signed(_zz_540) - $signed(_zz_539));
  assign _zz_8578 = ($signed(_zz_539) + $signed(_zz_540));
  assign _zz_8579 = _zz_8580[15 : 0];
  assign _zz_8580 = fixTo_401_dout;
  assign _zz_8581 = _zz_8582[15 : 0];
  assign _zz_8582 = fixTo_400_dout;
  assign _zz_8583 = _zz_8584;
  assign _zz_8584 = ($signed(_zz_8585) >>> _zz_2461);
  assign _zz_8585 = _zz_8586;
  assign _zz_8586 = ($signed(_zz_531) - $signed(_zz_2458));
  assign _zz_8587 = _zz_8588;
  assign _zz_8588 = ($signed(_zz_8589) >>> _zz_2461);
  assign _zz_8589 = _zz_8590;
  assign _zz_8590 = ($signed(_zz_532) - $signed(_zz_2459));
  assign _zz_8591 = _zz_8592;
  assign _zz_8592 = ($signed(_zz_8593) >>> _zz_2462);
  assign _zz_8593 = _zz_8594;
  assign _zz_8594 = ($signed(_zz_531) + $signed(_zz_2458));
  assign _zz_8595 = _zz_8596;
  assign _zz_8596 = ($signed(_zz_8597) >>> _zz_2462);
  assign _zz_8597 = _zz_8598;
  assign _zz_8598 = ($signed(_zz_532) + $signed(_zz_2459));
  assign _zz_8599 = ($signed(twiddle_factor_table_5_real) + $signed(twiddle_factor_table_5_imag));
  assign _zz_8600 = fixTo_402_dout;
  assign _zz_8601 = ($signed(_zz_542) - $signed(_zz_541));
  assign _zz_8602 = ($signed(_zz_541) + $signed(_zz_542));
  assign _zz_8603 = _zz_8604[15 : 0];
  assign _zz_8604 = fixTo_404_dout;
  assign _zz_8605 = _zz_8606[15 : 0];
  assign _zz_8606 = fixTo_403_dout;
  assign _zz_8607 = _zz_8608;
  assign _zz_8608 = ($signed(_zz_8609) >>> _zz_2466);
  assign _zz_8609 = _zz_8610;
  assign _zz_8610 = ($signed(_zz_533) - $signed(_zz_2463));
  assign _zz_8611 = _zz_8612;
  assign _zz_8612 = ($signed(_zz_8613) >>> _zz_2466);
  assign _zz_8613 = _zz_8614;
  assign _zz_8614 = ($signed(_zz_534) - $signed(_zz_2464));
  assign _zz_8615 = _zz_8616;
  assign _zz_8616 = ($signed(_zz_8617) >>> _zz_2467);
  assign _zz_8617 = _zz_8618;
  assign _zz_8618 = ($signed(_zz_533) + $signed(_zz_2463));
  assign _zz_8619 = _zz_8620;
  assign _zz_8620 = ($signed(_zz_8621) >>> _zz_2467);
  assign _zz_8621 = _zz_8622;
  assign _zz_8622 = ($signed(_zz_534) + $signed(_zz_2464));
  assign _zz_8623 = ($signed(twiddle_factor_table_6_real) + $signed(twiddle_factor_table_6_imag));
  assign _zz_8624 = fixTo_405_dout;
  assign _zz_8625 = ($signed(_zz_544) - $signed(_zz_543));
  assign _zz_8626 = ($signed(_zz_543) + $signed(_zz_544));
  assign _zz_8627 = _zz_8628[15 : 0];
  assign _zz_8628 = fixTo_407_dout;
  assign _zz_8629 = _zz_8630[15 : 0];
  assign _zz_8630 = fixTo_406_dout;
  assign _zz_8631 = _zz_8632;
  assign _zz_8632 = ($signed(_zz_8633) >>> _zz_2471);
  assign _zz_8633 = _zz_8634;
  assign _zz_8634 = ($signed(_zz_535) - $signed(_zz_2468));
  assign _zz_8635 = _zz_8636;
  assign _zz_8636 = ($signed(_zz_8637) >>> _zz_2471);
  assign _zz_8637 = _zz_8638;
  assign _zz_8638 = ($signed(_zz_536) - $signed(_zz_2469));
  assign _zz_8639 = _zz_8640;
  assign _zz_8640 = ($signed(_zz_8641) >>> _zz_2472);
  assign _zz_8641 = _zz_8642;
  assign _zz_8642 = ($signed(_zz_535) + $signed(_zz_2468));
  assign _zz_8643 = _zz_8644;
  assign _zz_8644 = ($signed(_zz_8645) >>> _zz_2472);
  assign _zz_8645 = _zz_8646;
  assign _zz_8646 = ($signed(_zz_536) + $signed(_zz_2469));
  assign _zz_8647 = ($signed(twiddle_factor_table_3_real) + $signed(twiddle_factor_table_3_imag));
  assign _zz_8648 = fixTo_408_dout;
  assign _zz_8649 = ($signed(_zz_554) - $signed(_zz_553));
  assign _zz_8650 = ($signed(_zz_553) + $signed(_zz_554));
  assign _zz_8651 = _zz_8652[15 : 0];
  assign _zz_8652 = fixTo_410_dout;
  assign _zz_8653 = _zz_8654[15 : 0];
  assign _zz_8654 = fixTo_409_dout;
  assign _zz_8655 = _zz_8656;
  assign _zz_8656 = ($signed(_zz_8657) >>> _zz_2476);
  assign _zz_8657 = _zz_8658;
  assign _zz_8658 = ($signed(_zz_545) - $signed(_zz_2473));
  assign _zz_8659 = _zz_8660;
  assign _zz_8660 = ($signed(_zz_8661) >>> _zz_2476);
  assign _zz_8661 = _zz_8662;
  assign _zz_8662 = ($signed(_zz_546) - $signed(_zz_2474));
  assign _zz_8663 = _zz_8664;
  assign _zz_8664 = ($signed(_zz_8665) >>> _zz_2477);
  assign _zz_8665 = _zz_8666;
  assign _zz_8666 = ($signed(_zz_545) + $signed(_zz_2473));
  assign _zz_8667 = _zz_8668;
  assign _zz_8668 = ($signed(_zz_8669) >>> _zz_2477);
  assign _zz_8669 = _zz_8670;
  assign _zz_8670 = ($signed(_zz_546) + $signed(_zz_2474));
  assign _zz_8671 = ($signed(twiddle_factor_table_4_real) + $signed(twiddle_factor_table_4_imag));
  assign _zz_8672 = fixTo_411_dout;
  assign _zz_8673 = ($signed(_zz_556) - $signed(_zz_555));
  assign _zz_8674 = ($signed(_zz_555) + $signed(_zz_556));
  assign _zz_8675 = _zz_8676[15 : 0];
  assign _zz_8676 = fixTo_413_dout;
  assign _zz_8677 = _zz_8678[15 : 0];
  assign _zz_8678 = fixTo_412_dout;
  assign _zz_8679 = _zz_8680;
  assign _zz_8680 = ($signed(_zz_8681) >>> _zz_2481);
  assign _zz_8681 = _zz_8682;
  assign _zz_8682 = ($signed(_zz_547) - $signed(_zz_2478));
  assign _zz_8683 = _zz_8684;
  assign _zz_8684 = ($signed(_zz_8685) >>> _zz_2481);
  assign _zz_8685 = _zz_8686;
  assign _zz_8686 = ($signed(_zz_548) - $signed(_zz_2479));
  assign _zz_8687 = _zz_8688;
  assign _zz_8688 = ($signed(_zz_8689) >>> _zz_2482);
  assign _zz_8689 = _zz_8690;
  assign _zz_8690 = ($signed(_zz_547) + $signed(_zz_2478));
  assign _zz_8691 = _zz_8692;
  assign _zz_8692 = ($signed(_zz_8693) >>> _zz_2482);
  assign _zz_8693 = _zz_8694;
  assign _zz_8694 = ($signed(_zz_548) + $signed(_zz_2479));
  assign _zz_8695 = ($signed(twiddle_factor_table_5_real) + $signed(twiddle_factor_table_5_imag));
  assign _zz_8696 = fixTo_414_dout;
  assign _zz_8697 = ($signed(_zz_558) - $signed(_zz_557));
  assign _zz_8698 = ($signed(_zz_557) + $signed(_zz_558));
  assign _zz_8699 = _zz_8700[15 : 0];
  assign _zz_8700 = fixTo_416_dout;
  assign _zz_8701 = _zz_8702[15 : 0];
  assign _zz_8702 = fixTo_415_dout;
  assign _zz_8703 = _zz_8704;
  assign _zz_8704 = ($signed(_zz_8705) >>> _zz_2486);
  assign _zz_8705 = _zz_8706;
  assign _zz_8706 = ($signed(_zz_549) - $signed(_zz_2483));
  assign _zz_8707 = _zz_8708;
  assign _zz_8708 = ($signed(_zz_8709) >>> _zz_2486);
  assign _zz_8709 = _zz_8710;
  assign _zz_8710 = ($signed(_zz_550) - $signed(_zz_2484));
  assign _zz_8711 = _zz_8712;
  assign _zz_8712 = ($signed(_zz_8713) >>> _zz_2487);
  assign _zz_8713 = _zz_8714;
  assign _zz_8714 = ($signed(_zz_549) + $signed(_zz_2483));
  assign _zz_8715 = _zz_8716;
  assign _zz_8716 = ($signed(_zz_8717) >>> _zz_2487);
  assign _zz_8717 = _zz_8718;
  assign _zz_8718 = ($signed(_zz_550) + $signed(_zz_2484));
  assign _zz_8719 = ($signed(twiddle_factor_table_6_real) + $signed(twiddle_factor_table_6_imag));
  assign _zz_8720 = fixTo_417_dout;
  assign _zz_8721 = ($signed(_zz_560) - $signed(_zz_559));
  assign _zz_8722 = ($signed(_zz_559) + $signed(_zz_560));
  assign _zz_8723 = _zz_8724[15 : 0];
  assign _zz_8724 = fixTo_419_dout;
  assign _zz_8725 = _zz_8726[15 : 0];
  assign _zz_8726 = fixTo_418_dout;
  assign _zz_8727 = _zz_8728;
  assign _zz_8728 = ($signed(_zz_8729) >>> _zz_2491);
  assign _zz_8729 = _zz_8730;
  assign _zz_8730 = ($signed(_zz_551) - $signed(_zz_2488));
  assign _zz_8731 = _zz_8732;
  assign _zz_8732 = ($signed(_zz_8733) >>> _zz_2491);
  assign _zz_8733 = _zz_8734;
  assign _zz_8734 = ($signed(_zz_552) - $signed(_zz_2489));
  assign _zz_8735 = _zz_8736;
  assign _zz_8736 = ($signed(_zz_8737) >>> _zz_2492);
  assign _zz_8737 = _zz_8738;
  assign _zz_8738 = ($signed(_zz_551) + $signed(_zz_2488));
  assign _zz_8739 = _zz_8740;
  assign _zz_8740 = ($signed(_zz_8741) >>> _zz_2492);
  assign _zz_8741 = _zz_8742;
  assign _zz_8742 = ($signed(_zz_552) + $signed(_zz_2489));
  assign _zz_8743 = ($signed(twiddle_factor_table_3_real) + $signed(twiddle_factor_table_3_imag));
  assign _zz_8744 = fixTo_420_dout;
  assign _zz_8745 = ($signed(_zz_570) - $signed(_zz_569));
  assign _zz_8746 = ($signed(_zz_569) + $signed(_zz_570));
  assign _zz_8747 = _zz_8748[15 : 0];
  assign _zz_8748 = fixTo_422_dout;
  assign _zz_8749 = _zz_8750[15 : 0];
  assign _zz_8750 = fixTo_421_dout;
  assign _zz_8751 = _zz_8752;
  assign _zz_8752 = ($signed(_zz_8753) >>> _zz_2496);
  assign _zz_8753 = _zz_8754;
  assign _zz_8754 = ($signed(_zz_561) - $signed(_zz_2493));
  assign _zz_8755 = _zz_8756;
  assign _zz_8756 = ($signed(_zz_8757) >>> _zz_2496);
  assign _zz_8757 = _zz_8758;
  assign _zz_8758 = ($signed(_zz_562) - $signed(_zz_2494));
  assign _zz_8759 = _zz_8760;
  assign _zz_8760 = ($signed(_zz_8761) >>> _zz_2497);
  assign _zz_8761 = _zz_8762;
  assign _zz_8762 = ($signed(_zz_561) + $signed(_zz_2493));
  assign _zz_8763 = _zz_8764;
  assign _zz_8764 = ($signed(_zz_8765) >>> _zz_2497);
  assign _zz_8765 = _zz_8766;
  assign _zz_8766 = ($signed(_zz_562) + $signed(_zz_2494));
  assign _zz_8767 = ($signed(twiddle_factor_table_4_real) + $signed(twiddle_factor_table_4_imag));
  assign _zz_8768 = fixTo_423_dout;
  assign _zz_8769 = ($signed(_zz_572) - $signed(_zz_571));
  assign _zz_8770 = ($signed(_zz_571) + $signed(_zz_572));
  assign _zz_8771 = _zz_8772[15 : 0];
  assign _zz_8772 = fixTo_425_dout;
  assign _zz_8773 = _zz_8774[15 : 0];
  assign _zz_8774 = fixTo_424_dout;
  assign _zz_8775 = _zz_8776;
  assign _zz_8776 = ($signed(_zz_8777) >>> _zz_2501);
  assign _zz_8777 = _zz_8778;
  assign _zz_8778 = ($signed(_zz_563) - $signed(_zz_2498));
  assign _zz_8779 = _zz_8780;
  assign _zz_8780 = ($signed(_zz_8781) >>> _zz_2501);
  assign _zz_8781 = _zz_8782;
  assign _zz_8782 = ($signed(_zz_564) - $signed(_zz_2499));
  assign _zz_8783 = _zz_8784;
  assign _zz_8784 = ($signed(_zz_8785) >>> _zz_2502);
  assign _zz_8785 = _zz_8786;
  assign _zz_8786 = ($signed(_zz_563) + $signed(_zz_2498));
  assign _zz_8787 = _zz_8788;
  assign _zz_8788 = ($signed(_zz_8789) >>> _zz_2502);
  assign _zz_8789 = _zz_8790;
  assign _zz_8790 = ($signed(_zz_564) + $signed(_zz_2499));
  assign _zz_8791 = ($signed(twiddle_factor_table_5_real) + $signed(twiddle_factor_table_5_imag));
  assign _zz_8792 = fixTo_426_dout;
  assign _zz_8793 = ($signed(_zz_574) - $signed(_zz_573));
  assign _zz_8794 = ($signed(_zz_573) + $signed(_zz_574));
  assign _zz_8795 = _zz_8796[15 : 0];
  assign _zz_8796 = fixTo_428_dout;
  assign _zz_8797 = _zz_8798[15 : 0];
  assign _zz_8798 = fixTo_427_dout;
  assign _zz_8799 = _zz_8800;
  assign _zz_8800 = ($signed(_zz_8801) >>> _zz_2506);
  assign _zz_8801 = _zz_8802;
  assign _zz_8802 = ($signed(_zz_565) - $signed(_zz_2503));
  assign _zz_8803 = _zz_8804;
  assign _zz_8804 = ($signed(_zz_8805) >>> _zz_2506);
  assign _zz_8805 = _zz_8806;
  assign _zz_8806 = ($signed(_zz_566) - $signed(_zz_2504));
  assign _zz_8807 = _zz_8808;
  assign _zz_8808 = ($signed(_zz_8809) >>> _zz_2507);
  assign _zz_8809 = _zz_8810;
  assign _zz_8810 = ($signed(_zz_565) + $signed(_zz_2503));
  assign _zz_8811 = _zz_8812;
  assign _zz_8812 = ($signed(_zz_8813) >>> _zz_2507);
  assign _zz_8813 = _zz_8814;
  assign _zz_8814 = ($signed(_zz_566) + $signed(_zz_2504));
  assign _zz_8815 = ($signed(twiddle_factor_table_6_real) + $signed(twiddle_factor_table_6_imag));
  assign _zz_8816 = fixTo_429_dout;
  assign _zz_8817 = ($signed(_zz_576) - $signed(_zz_575));
  assign _zz_8818 = ($signed(_zz_575) + $signed(_zz_576));
  assign _zz_8819 = _zz_8820[15 : 0];
  assign _zz_8820 = fixTo_431_dout;
  assign _zz_8821 = _zz_8822[15 : 0];
  assign _zz_8822 = fixTo_430_dout;
  assign _zz_8823 = _zz_8824;
  assign _zz_8824 = ($signed(_zz_8825) >>> _zz_2511);
  assign _zz_8825 = _zz_8826;
  assign _zz_8826 = ($signed(_zz_567) - $signed(_zz_2508));
  assign _zz_8827 = _zz_8828;
  assign _zz_8828 = ($signed(_zz_8829) >>> _zz_2511);
  assign _zz_8829 = _zz_8830;
  assign _zz_8830 = ($signed(_zz_568) - $signed(_zz_2509));
  assign _zz_8831 = _zz_8832;
  assign _zz_8832 = ($signed(_zz_8833) >>> _zz_2512);
  assign _zz_8833 = _zz_8834;
  assign _zz_8834 = ($signed(_zz_567) + $signed(_zz_2508));
  assign _zz_8835 = _zz_8836;
  assign _zz_8836 = ($signed(_zz_8837) >>> _zz_2512);
  assign _zz_8837 = _zz_8838;
  assign _zz_8838 = ($signed(_zz_568) + $signed(_zz_2509));
  assign _zz_8839 = ($signed(twiddle_factor_table_3_real) + $signed(twiddle_factor_table_3_imag));
  assign _zz_8840 = fixTo_432_dout;
  assign _zz_8841 = ($signed(_zz_586) - $signed(_zz_585));
  assign _zz_8842 = ($signed(_zz_585) + $signed(_zz_586));
  assign _zz_8843 = _zz_8844[15 : 0];
  assign _zz_8844 = fixTo_434_dout;
  assign _zz_8845 = _zz_8846[15 : 0];
  assign _zz_8846 = fixTo_433_dout;
  assign _zz_8847 = _zz_8848;
  assign _zz_8848 = ($signed(_zz_8849) >>> _zz_2516);
  assign _zz_8849 = _zz_8850;
  assign _zz_8850 = ($signed(_zz_577) - $signed(_zz_2513));
  assign _zz_8851 = _zz_8852;
  assign _zz_8852 = ($signed(_zz_8853) >>> _zz_2516);
  assign _zz_8853 = _zz_8854;
  assign _zz_8854 = ($signed(_zz_578) - $signed(_zz_2514));
  assign _zz_8855 = _zz_8856;
  assign _zz_8856 = ($signed(_zz_8857) >>> _zz_2517);
  assign _zz_8857 = _zz_8858;
  assign _zz_8858 = ($signed(_zz_577) + $signed(_zz_2513));
  assign _zz_8859 = _zz_8860;
  assign _zz_8860 = ($signed(_zz_8861) >>> _zz_2517);
  assign _zz_8861 = _zz_8862;
  assign _zz_8862 = ($signed(_zz_578) + $signed(_zz_2514));
  assign _zz_8863 = ($signed(twiddle_factor_table_4_real) + $signed(twiddle_factor_table_4_imag));
  assign _zz_8864 = fixTo_435_dout;
  assign _zz_8865 = ($signed(_zz_588) - $signed(_zz_587));
  assign _zz_8866 = ($signed(_zz_587) + $signed(_zz_588));
  assign _zz_8867 = _zz_8868[15 : 0];
  assign _zz_8868 = fixTo_437_dout;
  assign _zz_8869 = _zz_8870[15 : 0];
  assign _zz_8870 = fixTo_436_dout;
  assign _zz_8871 = _zz_8872;
  assign _zz_8872 = ($signed(_zz_8873) >>> _zz_2521);
  assign _zz_8873 = _zz_8874;
  assign _zz_8874 = ($signed(_zz_579) - $signed(_zz_2518));
  assign _zz_8875 = _zz_8876;
  assign _zz_8876 = ($signed(_zz_8877) >>> _zz_2521);
  assign _zz_8877 = _zz_8878;
  assign _zz_8878 = ($signed(_zz_580) - $signed(_zz_2519));
  assign _zz_8879 = _zz_8880;
  assign _zz_8880 = ($signed(_zz_8881) >>> _zz_2522);
  assign _zz_8881 = _zz_8882;
  assign _zz_8882 = ($signed(_zz_579) + $signed(_zz_2518));
  assign _zz_8883 = _zz_8884;
  assign _zz_8884 = ($signed(_zz_8885) >>> _zz_2522);
  assign _zz_8885 = _zz_8886;
  assign _zz_8886 = ($signed(_zz_580) + $signed(_zz_2519));
  assign _zz_8887 = ($signed(twiddle_factor_table_5_real) + $signed(twiddle_factor_table_5_imag));
  assign _zz_8888 = fixTo_438_dout;
  assign _zz_8889 = ($signed(_zz_590) - $signed(_zz_589));
  assign _zz_8890 = ($signed(_zz_589) + $signed(_zz_590));
  assign _zz_8891 = _zz_8892[15 : 0];
  assign _zz_8892 = fixTo_440_dout;
  assign _zz_8893 = _zz_8894[15 : 0];
  assign _zz_8894 = fixTo_439_dout;
  assign _zz_8895 = _zz_8896;
  assign _zz_8896 = ($signed(_zz_8897) >>> _zz_2526);
  assign _zz_8897 = _zz_8898;
  assign _zz_8898 = ($signed(_zz_581) - $signed(_zz_2523));
  assign _zz_8899 = _zz_8900;
  assign _zz_8900 = ($signed(_zz_8901) >>> _zz_2526);
  assign _zz_8901 = _zz_8902;
  assign _zz_8902 = ($signed(_zz_582) - $signed(_zz_2524));
  assign _zz_8903 = _zz_8904;
  assign _zz_8904 = ($signed(_zz_8905) >>> _zz_2527);
  assign _zz_8905 = _zz_8906;
  assign _zz_8906 = ($signed(_zz_581) + $signed(_zz_2523));
  assign _zz_8907 = _zz_8908;
  assign _zz_8908 = ($signed(_zz_8909) >>> _zz_2527);
  assign _zz_8909 = _zz_8910;
  assign _zz_8910 = ($signed(_zz_582) + $signed(_zz_2524));
  assign _zz_8911 = ($signed(twiddle_factor_table_6_real) + $signed(twiddle_factor_table_6_imag));
  assign _zz_8912 = fixTo_441_dout;
  assign _zz_8913 = ($signed(_zz_592) - $signed(_zz_591));
  assign _zz_8914 = ($signed(_zz_591) + $signed(_zz_592));
  assign _zz_8915 = _zz_8916[15 : 0];
  assign _zz_8916 = fixTo_443_dout;
  assign _zz_8917 = _zz_8918[15 : 0];
  assign _zz_8918 = fixTo_442_dout;
  assign _zz_8919 = _zz_8920;
  assign _zz_8920 = ($signed(_zz_8921) >>> _zz_2531);
  assign _zz_8921 = _zz_8922;
  assign _zz_8922 = ($signed(_zz_583) - $signed(_zz_2528));
  assign _zz_8923 = _zz_8924;
  assign _zz_8924 = ($signed(_zz_8925) >>> _zz_2531);
  assign _zz_8925 = _zz_8926;
  assign _zz_8926 = ($signed(_zz_584) - $signed(_zz_2529));
  assign _zz_8927 = _zz_8928;
  assign _zz_8928 = ($signed(_zz_8929) >>> _zz_2532);
  assign _zz_8929 = _zz_8930;
  assign _zz_8930 = ($signed(_zz_583) + $signed(_zz_2528));
  assign _zz_8931 = _zz_8932;
  assign _zz_8932 = ($signed(_zz_8933) >>> _zz_2532);
  assign _zz_8933 = _zz_8934;
  assign _zz_8934 = ($signed(_zz_584) + $signed(_zz_2529));
  assign _zz_8935 = ($signed(twiddle_factor_table_3_real) + $signed(twiddle_factor_table_3_imag));
  assign _zz_8936 = fixTo_444_dout;
  assign _zz_8937 = ($signed(_zz_602) - $signed(_zz_601));
  assign _zz_8938 = ($signed(_zz_601) + $signed(_zz_602));
  assign _zz_8939 = _zz_8940[15 : 0];
  assign _zz_8940 = fixTo_446_dout;
  assign _zz_8941 = _zz_8942[15 : 0];
  assign _zz_8942 = fixTo_445_dout;
  assign _zz_8943 = _zz_8944;
  assign _zz_8944 = ($signed(_zz_8945) >>> _zz_2536);
  assign _zz_8945 = _zz_8946;
  assign _zz_8946 = ($signed(_zz_593) - $signed(_zz_2533));
  assign _zz_8947 = _zz_8948;
  assign _zz_8948 = ($signed(_zz_8949) >>> _zz_2536);
  assign _zz_8949 = _zz_8950;
  assign _zz_8950 = ($signed(_zz_594) - $signed(_zz_2534));
  assign _zz_8951 = _zz_8952;
  assign _zz_8952 = ($signed(_zz_8953) >>> _zz_2537);
  assign _zz_8953 = _zz_8954;
  assign _zz_8954 = ($signed(_zz_593) + $signed(_zz_2533));
  assign _zz_8955 = _zz_8956;
  assign _zz_8956 = ($signed(_zz_8957) >>> _zz_2537);
  assign _zz_8957 = _zz_8958;
  assign _zz_8958 = ($signed(_zz_594) + $signed(_zz_2534));
  assign _zz_8959 = ($signed(twiddle_factor_table_4_real) + $signed(twiddle_factor_table_4_imag));
  assign _zz_8960 = fixTo_447_dout;
  assign _zz_8961 = ($signed(_zz_604) - $signed(_zz_603));
  assign _zz_8962 = ($signed(_zz_603) + $signed(_zz_604));
  assign _zz_8963 = _zz_8964[15 : 0];
  assign _zz_8964 = fixTo_449_dout;
  assign _zz_8965 = _zz_8966[15 : 0];
  assign _zz_8966 = fixTo_448_dout;
  assign _zz_8967 = _zz_8968;
  assign _zz_8968 = ($signed(_zz_8969) >>> _zz_2541);
  assign _zz_8969 = _zz_8970;
  assign _zz_8970 = ($signed(_zz_595) - $signed(_zz_2538));
  assign _zz_8971 = _zz_8972;
  assign _zz_8972 = ($signed(_zz_8973) >>> _zz_2541);
  assign _zz_8973 = _zz_8974;
  assign _zz_8974 = ($signed(_zz_596) - $signed(_zz_2539));
  assign _zz_8975 = _zz_8976;
  assign _zz_8976 = ($signed(_zz_8977) >>> _zz_2542);
  assign _zz_8977 = _zz_8978;
  assign _zz_8978 = ($signed(_zz_595) + $signed(_zz_2538));
  assign _zz_8979 = _zz_8980;
  assign _zz_8980 = ($signed(_zz_8981) >>> _zz_2542);
  assign _zz_8981 = _zz_8982;
  assign _zz_8982 = ($signed(_zz_596) + $signed(_zz_2539));
  assign _zz_8983 = ($signed(twiddle_factor_table_5_real) + $signed(twiddle_factor_table_5_imag));
  assign _zz_8984 = fixTo_450_dout;
  assign _zz_8985 = ($signed(_zz_606) - $signed(_zz_605));
  assign _zz_8986 = ($signed(_zz_605) + $signed(_zz_606));
  assign _zz_8987 = _zz_8988[15 : 0];
  assign _zz_8988 = fixTo_452_dout;
  assign _zz_8989 = _zz_8990[15 : 0];
  assign _zz_8990 = fixTo_451_dout;
  assign _zz_8991 = _zz_8992;
  assign _zz_8992 = ($signed(_zz_8993) >>> _zz_2546);
  assign _zz_8993 = _zz_8994;
  assign _zz_8994 = ($signed(_zz_597) - $signed(_zz_2543));
  assign _zz_8995 = _zz_8996;
  assign _zz_8996 = ($signed(_zz_8997) >>> _zz_2546);
  assign _zz_8997 = _zz_8998;
  assign _zz_8998 = ($signed(_zz_598) - $signed(_zz_2544));
  assign _zz_8999 = _zz_9000;
  assign _zz_9000 = ($signed(_zz_9001) >>> _zz_2547);
  assign _zz_9001 = _zz_9002;
  assign _zz_9002 = ($signed(_zz_597) + $signed(_zz_2543));
  assign _zz_9003 = _zz_9004;
  assign _zz_9004 = ($signed(_zz_9005) >>> _zz_2547);
  assign _zz_9005 = _zz_9006;
  assign _zz_9006 = ($signed(_zz_598) + $signed(_zz_2544));
  assign _zz_9007 = ($signed(twiddle_factor_table_6_real) + $signed(twiddle_factor_table_6_imag));
  assign _zz_9008 = fixTo_453_dout;
  assign _zz_9009 = ($signed(_zz_608) - $signed(_zz_607));
  assign _zz_9010 = ($signed(_zz_607) + $signed(_zz_608));
  assign _zz_9011 = _zz_9012[15 : 0];
  assign _zz_9012 = fixTo_455_dout;
  assign _zz_9013 = _zz_9014[15 : 0];
  assign _zz_9014 = fixTo_454_dout;
  assign _zz_9015 = _zz_9016;
  assign _zz_9016 = ($signed(_zz_9017) >>> _zz_2551);
  assign _zz_9017 = _zz_9018;
  assign _zz_9018 = ($signed(_zz_599) - $signed(_zz_2548));
  assign _zz_9019 = _zz_9020;
  assign _zz_9020 = ($signed(_zz_9021) >>> _zz_2551);
  assign _zz_9021 = _zz_9022;
  assign _zz_9022 = ($signed(_zz_600) - $signed(_zz_2549));
  assign _zz_9023 = _zz_9024;
  assign _zz_9024 = ($signed(_zz_9025) >>> _zz_2552);
  assign _zz_9025 = _zz_9026;
  assign _zz_9026 = ($signed(_zz_599) + $signed(_zz_2548));
  assign _zz_9027 = _zz_9028;
  assign _zz_9028 = ($signed(_zz_9029) >>> _zz_2552);
  assign _zz_9029 = _zz_9030;
  assign _zz_9030 = ($signed(_zz_600) + $signed(_zz_2549));
  assign _zz_9031 = ($signed(twiddle_factor_table_3_real) + $signed(twiddle_factor_table_3_imag));
  assign _zz_9032 = fixTo_456_dout;
  assign _zz_9033 = ($signed(_zz_618) - $signed(_zz_617));
  assign _zz_9034 = ($signed(_zz_617) + $signed(_zz_618));
  assign _zz_9035 = _zz_9036[15 : 0];
  assign _zz_9036 = fixTo_458_dout;
  assign _zz_9037 = _zz_9038[15 : 0];
  assign _zz_9038 = fixTo_457_dout;
  assign _zz_9039 = _zz_9040;
  assign _zz_9040 = ($signed(_zz_9041) >>> _zz_2556);
  assign _zz_9041 = _zz_9042;
  assign _zz_9042 = ($signed(_zz_609) - $signed(_zz_2553));
  assign _zz_9043 = _zz_9044;
  assign _zz_9044 = ($signed(_zz_9045) >>> _zz_2556);
  assign _zz_9045 = _zz_9046;
  assign _zz_9046 = ($signed(_zz_610) - $signed(_zz_2554));
  assign _zz_9047 = _zz_9048;
  assign _zz_9048 = ($signed(_zz_9049) >>> _zz_2557);
  assign _zz_9049 = _zz_9050;
  assign _zz_9050 = ($signed(_zz_609) + $signed(_zz_2553));
  assign _zz_9051 = _zz_9052;
  assign _zz_9052 = ($signed(_zz_9053) >>> _zz_2557);
  assign _zz_9053 = _zz_9054;
  assign _zz_9054 = ($signed(_zz_610) + $signed(_zz_2554));
  assign _zz_9055 = ($signed(twiddle_factor_table_4_real) + $signed(twiddle_factor_table_4_imag));
  assign _zz_9056 = fixTo_459_dout;
  assign _zz_9057 = ($signed(_zz_620) - $signed(_zz_619));
  assign _zz_9058 = ($signed(_zz_619) + $signed(_zz_620));
  assign _zz_9059 = _zz_9060[15 : 0];
  assign _zz_9060 = fixTo_461_dout;
  assign _zz_9061 = _zz_9062[15 : 0];
  assign _zz_9062 = fixTo_460_dout;
  assign _zz_9063 = _zz_9064;
  assign _zz_9064 = ($signed(_zz_9065) >>> _zz_2561);
  assign _zz_9065 = _zz_9066;
  assign _zz_9066 = ($signed(_zz_611) - $signed(_zz_2558));
  assign _zz_9067 = _zz_9068;
  assign _zz_9068 = ($signed(_zz_9069) >>> _zz_2561);
  assign _zz_9069 = _zz_9070;
  assign _zz_9070 = ($signed(_zz_612) - $signed(_zz_2559));
  assign _zz_9071 = _zz_9072;
  assign _zz_9072 = ($signed(_zz_9073) >>> _zz_2562);
  assign _zz_9073 = _zz_9074;
  assign _zz_9074 = ($signed(_zz_611) + $signed(_zz_2558));
  assign _zz_9075 = _zz_9076;
  assign _zz_9076 = ($signed(_zz_9077) >>> _zz_2562);
  assign _zz_9077 = _zz_9078;
  assign _zz_9078 = ($signed(_zz_612) + $signed(_zz_2559));
  assign _zz_9079 = ($signed(twiddle_factor_table_5_real) + $signed(twiddle_factor_table_5_imag));
  assign _zz_9080 = fixTo_462_dout;
  assign _zz_9081 = ($signed(_zz_622) - $signed(_zz_621));
  assign _zz_9082 = ($signed(_zz_621) + $signed(_zz_622));
  assign _zz_9083 = _zz_9084[15 : 0];
  assign _zz_9084 = fixTo_464_dout;
  assign _zz_9085 = _zz_9086[15 : 0];
  assign _zz_9086 = fixTo_463_dout;
  assign _zz_9087 = _zz_9088;
  assign _zz_9088 = ($signed(_zz_9089) >>> _zz_2566);
  assign _zz_9089 = _zz_9090;
  assign _zz_9090 = ($signed(_zz_613) - $signed(_zz_2563));
  assign _zz_9091 = _zz_9092;
  assign _zz_9092 = ($signed(_zz_9093) >>> _zz_2566);
  assign _zz_9093 = _zz_9094;
  assign _zz_9094 = ($signed(_zz_614) - $signed(_zz_2564));
  assign _zz_9095 = _zz_9096;
  assign _zz_9096 = ($signed(_zz_9097) >>> _zz_2567);
  assign _zz_9097 = _zz_9098;
  assign _zz_9098 = ($signed(_zz_613) + $signed(_zz_2563));
  assign _zz_9099 = _zz_9100;
  assign _zz_9100 = ($signed(_zz_9101) >>> _zz_2567);
  assign _zz_9101 = _zz_9102;
  assign _zz_9102 = ($signed(_zz_614) + $signed(_zz_2564));
  assign _zz_9103 = ($signed(twiddle_factor_table_6_real) + $signed(twiddle_factor_table_6_imag));
  assign _zz_9104 = fixTo_465_dout;
  assign _zz_9105 = ($signed(_zz_624) - $signed(_zz_623));
  assign _zz_9106 = ($signed(_zz_623) + $signed(_zz_624));
  assign _zz_9107 = _zz_9108[15 : 0];
  assign _zz_9108 = fixTo_467_dout;
  assign _zz_9109 = _zz_9110[15 : 0];
  assign _zz_9110 = fixTo_466_dout;
  assign _zz_9111 = _zz_9112;
  assign _zz_9112 = ($signed(_zz_9113) >>> _zz_2571);
  assign _zz_9113 = _zz_9114;
  assign _zz_9114 = ($signed(_zz_615) - $signed(_zz_2568));
  assign _zz_9115 = _zz_9116;
  assign _zz_9116 = ($signed(_zz_9117) >>> _zz_2571);
  assign _zz_9117 = _zz_9118;
  assign _zz_9118 = ($signed(_zz_616) - $signed(_zz_2569));
  assign _zz_9119 = _zz_9120;
  assign _zz_9120 = ($signed(_zz_9121) >>> _zz_2572);
  assign _zz_9121 = _zz_9122;
  assign _zz_9122 = ($signed(_zz_615) + $signed(_zz_2568));
  assign _zz_9123 = _zz_9124;
  assign _zz_9124 = ($signed(_zz_9125) >>> _zz_2572);
  assign _zz_9125 = _zz_9126;
  assign _zz_9126 = ($signed(_zz_616) + $signed(_zz_2569));
  assign _zz_9127 = ($signed(twiddle_factor_table_3_real) + $signed(twiddle_factor_table_3_imag));
  assign _zz_9128 = fixTo_468_dout;
  assign _zz_9129 = ($signed(_zz_634) - $signed(_zz_633));
  assign _zz_9130 = ($signed(_zz_633) + $signed(_zz_634));
  assign _zz_9131 = _zz_9132[15 : 0];
  assign _zz_9132 = fixTo_470_dout;
  assign _zz_9133 = _zz_9134[15 : 0];
  assign _zz_9134 = fixTo_469_dout;
  assign _zz_9135 = _zz_9136;
  assign _zz_9136 = ($signed(_zz_9137) >>> _zz_2576);
  assign _zz_9137 = _zz_9138;
  assign _zz_9138 = ($signed(_zz_625) - $signed(_zz_2573));
  assign _zz_9139 = _zz_9140;
  assign _zz_9140 = ($signed(_zz_9141) >>> _zz_2576);
  assign _zz_9141 = _zz_9142;
  assign _zz_9142 = ($signed(_zz_626) - $signed(_zz_2574));
  assign _zz_9143 = _zz_9144;
  assign _zz_9144 = ($signed(_zz_9145) >>> _zz_2577);
  assign _zz_9145 = _zz_9146;
  assign _zz_9146 = ($signed(_zz_625) + $signed(_zz_2573));
  assign _zz_9147 = _zz_9148;
  assign _zz_9148 = ($signed(_zz_9149) >>> _zz_2577);
  assign _zz_9149 = _zz_9150;
  assign _zz_9150 = ($signed(_zz_626) + $signed(_zz_2574));
  assign _zz_9151 = ($signed(twiddle_factor_table_4_real) + $signed(twiddle_factor_table_4_imag));
  assign _zz_9152 = fixTo_471_dout;
  assign _zz_9153 = ($signed(_zz_636) - $signed(_zz_635));
  assign _zz_9154 = ($signed(_zz_635) + $signed(_zz_636));
  assign _zz_9155 = _zz_9156[15 : 0];
  assign _zz_9156 = fixTo_473_dout;
  assign _zz_9157 = _zz_9158[15 : 0];
  assign _zz_9158 = fixTo_472_dout;
  assign _zz_9159 = _zz_9160;
  assign _zz_9160 = ($signed(_zz_9161) >>> _zz_2581);
  assign _zz_9161 = _zz_9162;
  assign _zz_9162 = ($signed(_zz_627) - $signed(_zz_2578));
  assign _zz_9163 = _zz_9164;
  assign _zz_9164 = ($signed(_zz_9165) >>> _zz_2581);
  assign _zz_9165 = _zz_9166;
  assign _zz_9166 = ($signed(_zz_628) - $signed(_zz_2579));
  assign _zz_9167 = _zz_9168;
  assign _zz_9168 = ($signed(_zz_9169) >>> _zz_2582);
  assign _zz_9169 = _zz_9170;
  assign _zz_9170 = ($signed(_zz_627) + $signed(_zz_2578));
  assign _zz_9171 = _zz_9172;
  assign _zz_9172 = ($signed(_zz_9173) >>> _zz_2582);
  assign _zz_9173 = _zz_9174;
  assign _zz_9174 = ($signed(_zz_628) + $signed(_zz_2579));
  assign _zz_9175 = ($signed(twiddle_factor_table_5_real) + $signed(twiddle_factor_table_5_imag));
  assign _zz_9176 = fixTo_474_dout;
  assign _zz_9177 = ($signed(_zz_638) - $signed(_zz_637));
  assign _zz_9178 = ($signed(_zz_637) + $signed(_zz_638));
  assign _zz_9179 = _zz_9180[15 : 0];
  assign _zz_9180 = fixTo_476_dout;
  assign _zz_9181 = _zz_9182[15 : 0];
  assign _zz_9182 = fixTo_475_dout;
  assign _zz_9183 = _zz_9184;
  assign _zz_9184 = ($signed(_zz_9185) >>> _zz_2586);
  assign _zz_9185 = _zz_9186;
  assign _zz_9186 = ($signed(_zz_629) - $signed(_zz_2583));
  assign _zz_9187 = _zz_9188;
  assign _zz_9188 = ($signed(_zz_9189) >>> _zz_2586);
  assign _zz_9189 = _zz_9190;
  assign _zz_9190 = ($signed(_zz_630) - $signed(_zz_2584));
  assign _zz_9191 = _zz_9192;
  assign _zz_9192 = ($signed(_zz_9193) >>> _zz_2587);
  assign _zz_9193 = _zz_9194;
  assign _zz_9194 = ($signed(_zz_629) + $signed(_zz_2583));
  assign _zz_9195 = _zz_9196;
  assign _zz_9196 = ($signed(_zz_9197) >>> _zz_2587);
  assign _zz_9197 = _zz_9198;
  assign _zz_9198 = ($signed(_zz_630) + $signed(_zz_2584));
  assign _zz_9199 = ($signed(twiddle_factor_table_6_real) + $signed(twiddle_factor_table_6_imag));
  assign _zz_9200 = fixTo_477_dout;
  assign _zz_9201 = ($signed(_zz_640) - $signed(_zz_639));
  assign _zz_9202 = ($signed(_zz_639) + $signed(_zz_640));
  assign _zz_9203 = _zz_9204[15 : 0];
  assign _zz_9204 = fixTo_479_dout;
  assign _zz_9205 = _zz_9206[15 : 0];
  assign _zz_9206 = fixTo_478_dout;
  assign _zz_9207 = _zz_9208;
  assign _zz_9208 = ($signed(_zz_9209) >>> _zz_2591);
  assign _zz_9209 = _zz_9210;
  assign _zz_9210 = ($signed(_zz_631) - $signed(_zz_2588));
  assign _zz_9211 = _zz_9212;
  assign _zz_9212 = ($signed(_zz_9213) >>> _zz_2591);
  assign _zz_9213 = _zz_9214;
  assign _zz_9214 = ($signed(_zz_632) - $signed(_zz_2589));
  assign _zz_9215 = _zz_9216;
  assign _zz_9216 = ($signed(_zz_9217) >>> _zz_2592);
  assign _zz_9217 = _zz_9218;
  assign _zz_9218 = ($signed(_zz_631) + $signed(_zz_2588));
  assign _zz_9219 = _zz_9220;
  assign _zz_9220 = ($signed(_zz_9221) >>> _zz_2592);
  assign _zz_9221 = _zz_9222;
  assign _zz_9222 = ($signed(_zz_632) + $signed(_zz_2589));
  assign _zz_9223 = ($signed(twiddle_factor_table_3_real) + $signed(twiddle_factor_table_3_imag));
  assign _zz_9224 = fixTo_480_dout;
  assign _zz_9225 = ($signed(_zz_650) - $signed(_zz_649));
  assign _zz_9226 = ($signed(_zz_649) + $signed(_zz_650));
  assign _zz_9227 = _zz_9228[15 : 0];
  assign _zz_9228 = fixTo_482_dout;
  assign _zz_9229 = _zz_9230[15 : 0];
  assign _zz_9230 = fixTo_481_dout;
  assign _zz_9231 = _zz_9232;
  assign _zz_9232 = ($signed(_zz_9233) >>> _zz_2596);
  assign _zz_9233 = _zz_9234;
  assign _zz_9234 = ($signed(_zz_641) - $signed(_zz_2593));
  assign _zz_9235 = _zz_9236;
  assign _zz_9236 = ($signed(_zz_9237) >>> _zz_2596);
  assign _zz_9237 = _zz_9238;
  assign _zz_9238 = ($signed(_zz_642) - $signed(_zz_2594));
  assign _zz_9239 = _zz_9240;
  assign _zz_9240 = ($signed(_zz_9241) >>> _zz_2597);
  assign _zz_9241 = _zz_9242;
  assign _zz_9242 = ($signed(_zz_641) + $signed(_zz_2593));
  assign _zz_9243 = _zz_9244;
  assign _zz_9244 = ($signed(_zz_9245) >>> _zz_2597);
  assign _zz_9245 = _zz_9246;
  assign _zz_9246 = ($signed(_zz_642) + $signed(_zz_2594));
  assign _zz_9247 = ($signed(twiddle_factor_table_4_real) + $signed(twiddle_factor_table_4_imag));
  assign _zz_9248 = fixTo_483_dout;
  assign _zz_9249 = ($signed(_zz_652) - $signed(_zz_651));
  assign _zz_9250 = ($signed(_zz_651) + $signed(_zz_652));
  assign _zz_9251 = _zz_9252[15 : 0];
  assign _zz_9252 = fixTo_485_dout;
  assign _zz_9253 = _zz_9254[15 : 0];
  assign _zz_9254 = fixTo_484_dout;
  assign _zz_9255 = _zz_9256;
  assign _zz_9256 = ($signed(_zz_9257) >>> _zz_2601);
  assign _zz_9257 = _zz_9258;
  assign _zz_9258 = ($signed(_zz_643) - $signed(_zz_2598));
  assign _zz_9259 = _zz_9260;
  assign _zz_9260 = ($signed(_zz_9261) >>> _zz_2601);
  assign _zz_9261 = _zz_9262;
  assign _zz_9262 = ($signed(_zz_644) - $signed(_zz_2599));
  assign _zz_9263 = _zz_9264;
  assign _zz_9264 = ($signed(_zz_9265) >>> _zz_2602);
  assign _zz_9265 = _zz_9266;
  assign _zz_9266 = ($signed(_zz_643) + $signed(_zz_2598));
  assign _zz_9267 = _zz_9268;
  assign _zz_9268 = ($signed(_zz_9269) >>> _zz_2602);
  assign _zz_9269 = _zz_9270;
  assign _zz_9270 = ($signed(_zz_644) + $signed(_zz_2599));
  assign _zz_9271 = ($signed(twiddle_factor_table_5_real) + $signed(twiddle_factor_table_5_imag));
  assign _zz_9272 = fixTo_486_dout;
  assign _zz_9273 = ($signed(_zz_654) - $signed(_zz_653));
  assign _zz_9274 = ($signed(_zz_653) + $signed(_zz_654));
  assign _zz_9275 = _zz_9276[15 : 0];
  assign _zz_9276 = fixTo_488_dout;
  assign _zz_9277 = _zz_9278[15 : 0];
  assign _zz_9278 = fixTo_487_dout;
  assign _zz_9279 = _zz_9280;
  assign _zz_9280 = ($signed(_zz_9281) >>> _zz_2606);
  assign _zz_9281 = _zz_9282;
  assign _zz_9282 = ($signed(_zz_645) - $signed(_zz_2603));
  assign _zz_9283 = _zz_9284;
  assign _zz_9284 = ($signed(_zz_9285) >>> _zz_2606);
  assign _zz_9285 = _zz_9286;
  assign _zz_9286 = ($signed(_zz_646) - $signed(_zz_2604));
  assign _zz_9287 = _zz_9288;
  assign _zz_9288 = ($signed(_zz_9289) >>> _zz_2607);
  assign _zz_9289 = _zz_9290;
  assign _zz_9290 = ($signed(_zz_645) + $signed(_zz_2603));
  assign _zz_9291 = _zz_9292;
  assign _zz_9292 = ($signed(_zz_9293) >>> _zz_2607);
  assign _zz_9293 = _zz_9294;
  assign _zz_9294 = ($signed(_zz_646) + $signed(_zz_2604));
  assign _zz_9295 = ($signed(twiddle_factor_table_6_real) + $signed(twiddle_factor_table_6_imag));
  assign _zz_9296 = fixTo_489_dout;
  assign _zz_9297 = ($signed(_zz_656) - $signed(_zz_655));
  assign _zz_9298 = ($signed(_zz_655) + $signed(_zz_656));
  assign _zz_9299 = _zz_9300[15 : 0];
  assign _zz_9300 = fixTo_491_dout;
  assign _zz_9301 = _zz_9302[15 : 0];
  assign _zz_9302 = fixTo_490_dout;
  assign _zz_9303 = _zz_9304;
  assign _zz_9304 = ($signed(_zz_9305) >>> _zz_2611);
  assign _zz_9305 = _zz_9306;
  assign _zz_9306 = ($signed(_zz_647) - $signed(_zz_2608));
  assign _zz_9307 = _zz_9308;
  assign _zz_9308 = ($signed(_zz_9309) >>> _zz_2611);
  assign _zz_9309 = _zz_9310;
  assign _zz_9310 = ($signed(_zz_648) - $signed(_zz_2609));
  assign _zz_9311 = _zz_9312;
  assign _zz_9312 = ($signed(_zz_9313) >>> _zz_2612);
  assign _zz_9313 = _zz_9314;
  assign _zz_9314 = ($signed(_zz_647) + $signed(_zz_2608));
  assign _zz_9315 = _zz_9316;
  assign _zz_9316 = ($signed(_zz_9317) >>> _zz_2612);
  assign _zz_9317 = _zz_9318;
  assign _zz_9318 = ($signed(_zz_648) + $signed(_zz_2609));
  assign _zz_9319 = ($signed(twiddle_factor_table_3_real) + $signed(twiddle_factor_table_3_imag));
  assign _zz_9320 = fixTo_492_dout;
  assign _zz_9321 = ($signed(_zz_666) - $signed(_zz_665));
  assign _zz_9322 = ($signed(_zz_665) + $signed(_zz_666));
  assign _zz_9323 = _zz_9324[15 : 0];
  assign _zz_9324 = fixTo_494_dout;
  assign _zz_9325 = _zz_9326[15 : 0];
  assign _zz_9326 = fixTo_493_dout;
  assign _zz_9327 = _zz_9328;
  assign _zz_9328 = ($signed(_zz_9329) >>> _zz_2616);
  assign _zz_9329 = _zz_9330;
  assign _zz_9330 = ($signed(_zz_657) - $signed(_zz_2613));
  assign _zz_9331 = _zz_9332;
  assign _zz_9332 = ($signed(_zz_9333) >>> _zz_2616);
  assign _zz_9333 = _zz_9334;
  assign _zz_9334 = ($signed(_zz_658) - $signed(_zz_2614));
  assign _zz_9335 = _zz_9336;
  assign _zz_9336 = ($signed(_zz_9337) >>> _zz_2617);
  assign _zz_9337 = _zz_9338;
  assign _zz_9338 = ($signed(_zz_657) + $signed(_zz_2613));
  assign _zz_9339 = _zz_9340;
  assign _zz_9340 = ($signed(_zz_9341) >>> _zz_2617);
  assign _zz_9341 = _zz_9342;
  assign _zz_9342 = ($signed(_zz_658) + $signed(_zz_2614));
  assign _zz_9343 = ($signed(twiddle_factor_table_4_real) + $signed(twiddle_factor_table_4_imag));
  assign _zz_9344 = fixTo_495_dout;
  assign _zz_9345 = ($signed(_zz_668) - $signed(_zz_667));
  assign _zz_9346 = ($signed(_zz_667) + $signed(_zz_668));
  assign _zz_9347 = _zz_9348[15 : 0];
  assign _zz_9348 = fixTo_497_dout;
  assign _zz_9349 = _zz_9350[15 : 0];
  assign _zz_9350 = fixTo_496_dout;
  assign _zz_9351 = _zz_9352;
  assign _zz_9352 = ($signed(_zz_9353) >>> _zz_2621);
  assign _zz_9353 = _zz_9354;
  assign _zz_9354 = ($signed(_zz_659) - $signed(_zz_2618));
  assign _zz_9355 = _zz_9356;
  assign _zz_9356 = ($signed(_zz_9357) >>> _zz_2621);
  assign _zz_9357 = _zz_9358;
  assign _zz_9358 = ($signed(_zz_660) - $signed(_zz_2619));
  assign _zz_9359 = _zz_9360;
  assign _zz_9360 = ($signed(_zz_9361) >>> _zz_2622);
  assign _zz_9361 = _zz_9362;
  assign _zz_9362 = ($signed(_zz_659) + $signed(_zz_2618));
  assign _zz_9363 = _zz_9364;
  assign _zz_9364 = ($signed(_zz_9365) >>> _zz_2622);
  assign _zz_9365 = _zz_9366;
  assign _zz_9366 = ($signed(_zz_660) + $signed(_zz_2619));
  assign _zz_9367 = ($signed(twiddle_factor_table_5_real) + $signed(twiddle_factor_table_5_imag));
  assign _zz_9368 = fixTo_498_dout;
  assign _zz_9369 = ($signed(_zz_670) - $signed(_zz_669));
  assign _zz_9370 = ($signed(_zz_669) + $signed(_zz_670));
  assign _zz_9371 = _zz_9372[15 : 0];
  assign _zz_9372 = fixTo_500_dout;
  assign _zz_9373 = _zz_9374[15 : 0];
  assign _zz_9374 = fixTo_499_dout;
  assign _zz_9375 = _zz_9376;
  assign _zz_9376 = ($signed(_zz_9377) >>> _zz_2626);
  assign _zz_9377 = _zz_9378;
  assign _zz_9378 = ($signed(_zz_661) - $signed(_zz_2623));
  assign _zz_9379 = _zz_9380;
  assign _zz_9380 = ($signed(_zz_9381) >>> _zz_2626);
  assign _zz_9381 = _zz_9382;
  assign _zz_9382 = ($signed(_zz_662) - $signed(_zz_2624));
  assign _zz_9383 = _zz_9384;
  assign _zz_9384 = ($signed(_zz_9385) >>> _zz_2627);
  assign _zz_9385 = _zz_9386;
  assign _zz_9386 = ($signed(_zz_661) + $signed(_zz_2623));
  assign _zz_9387 = _zz_9388;
  assign _zz_9388 = ($signed(_zz_9389) >>> _zz_2627);
  assign _zz_9389 = _zz_9390;
  assign _zz_9390 = ($signed(_zz_662) + $signed(_zz_2624));
  assign _zz_9391 = ($signed(twiddle_factor_table_6_real) + $signed(twiddle_factor_table_6_imag));
  assign _zz_9392 = fixTo_501_dout;
  assign _zz_9393 = ($signed(_zz_672) - $signed(_zz_671));
  assign _zz_9394 = ($signed(_zz_671) + $signed(_zz_672));
  assign _zz_9395 = _zz_9396[15 : 0];
  assign _zz_9396 = fixTo_503_dout;
  assign _zz_9397 = _zz_9398[15 : 0];
  assign _zz_9398 = fixTo_502_dout;
  assign _zz_9399 = _zz_9400;
  assign _zz_9400 = ($signed(_zz_9401) >>> _zz_2631);
  assign _zz_9401 = _zz_9402;
  assign _zz_9402 = ($signed(_zz_663) - $signed(_zz_2628));
  assign _zz_9403 = _zz_9404;
  assign _zz_9404 = ($signed(_zz_9405) >>> _zz_2631);
  assign _zz_9405 = _zz_9406;
  assign _zz_9406 = ($signed(_zz_664) - $signed(_zz_2629));
  assign _zz_9407 = _zz_9408;
  assign _zz_9408 = ($signed(_zz_9409) >>> _zz_2632);
  assign _zz_9409 = _zz_9410;
  assign _zz_9410 = ($signed(_zz_663) + $signed(_zz_2628));
  assign _zz_9411 = _zz_9412;
  assign _zz_9412 = ($signed(_zz_9413) >>> _zz_2632);
  assign _zz_9413 = _zz_9414;
  assign _zz_9414 = ($signed(_zz_664) + $signed(_zz_2629));
  assign _zz_9415 = ($signed(twiddle_factor_table_3_real) + $signed(twiddle_factor_table_3_imag));
  assign _zz_9416 = fixTo_504_dout;
  assign _zz_9417 = ($signed(_zz_682) - $signed(_zz_681));
  assign _zz_9418 = ($signed(_zz_681) + $signed(_zz_682));
  assign _zz_9419 = _zz_9420[15 : 0];
  assign _zz_9420 = fixTo_506_dout;
  assign _zz_9421 = _zz_9422[15 : 0];
  assign _zz_9422 = fixTo_505_dout;
  assign _zz_9423 = _zz_9424;
  assign _zz_9424 = ($signed(_zz_9425) >>> _zz_2636);
  assign _zz_9425 = _zz_9426;
  assign _zz_9426 = ($signed(_zz_673) - $signed(_zz_2633));
  assign _zz_9427 = _zz_9428;
  assign _zz_9428 = ($signed(_zz_9429) >>> _zz_2636);
  assign _zz_9429 = _zz_9430;
  assign _zz_9430 = ($signed(_zz_674) - $signed(_zz_2634));
  assign _zz_9431 = _zz_9432;
  assign _zz_9432 = ($signed(_zz_9433) >>> _zz_2637);
  assign _zz_9433 = _zz_9434;
  assign _zz_9434 = ($signed(_zz_673) + $signed(_zz_2633));
  assign _zz_9435 = _zz_9436;
  assign _zz_9436 = ($signed(_zz_9437) >>> _zz_2637);
  assign _zz_9437 = _zz_9438;
  assign _zz_9438 = ($signed(_zz_674) + $signed(_zz_2634));
  assign _zz_9439 = ($signed(twiddle_factor_table_4_real) + $signed(twiddle_factor_table_4_imag));
  assign _zz_9440 = fixTo_507_dout;
  assign _zz_9441 = ($signed(_zz_684) - $signed(_zz_683));
  assign _zz_9442 = ($signed(_zz_683) + $signed(_zz_684));
  assign _zz_9443 = _zz_9444[15 : 0];
  assign _zz_9444 = fixTo_509_dout;
  assign _zz_9445 = _zz_9446[15 : 0];
  assign _zz_9446 = fixTo_508_dout;
  assign _zz_9447 = _zz_9448;
  assign _zz_9448 = ($signed(_zz_9449) >>> _zz_2641);
  assign _zz_9449 = _zz_9450;
  assign _zz_9450 = ($signed(_zz_675) - $signed(_zz_2638));
  assign _zz_9451 = _zz_9452;
  assign _zz_9452 = ($signed(_zz_9453) >>> _zz_2641);
  assign _zz_9453 = _zz_9454;
  assign _zz_9454 = ($signed(_zz_676) - $signed(_zz_2639));
  assign _zz_9455 = _zz_9456;
  assign _zz_9456 = ($signed(_zz_9457) >>> _zz_2642);
  assign _zz_9457 = _zz_9458;
  assign _zz_9458 = ($signed(_zz_675) + $signed(_zz_2638));
  assign _zz_9459 = _zz_9460;
  assign _zz_9460 = ($signed(_zz_9461) >>> _zz_2642);
  assign _zz_9461 = _zz_9462;
  assign _zz_9462 = ($signed(_zz_676) + $signed(_zz_2639));
  assign _zz_9463 = ($signed(twiddle_factor_table_5_real) + $signed(twiddle_factor_table_5_imag));
  assign _zz_9464 = fixTo_510_dout;
  assign _zz_9465 = ($signed(_zz_686) - $signed(_zz_685));
  assign _zz_9466 = ($signed(_zz_685) + $signed(_zz_686));
  assign _zz_9467 = _zz_9468[15 : 0];
  assign _zz_9468 = fixTo_512_dout;
  assign _zz_9469 = _zz_9470[15 : 0];
  assign _zz_9470 = fixTo_511_dout;
  assign _zz_9471 = _zz_9472;
  assign _zz_9472 = ($signed(_zz_9473) >>> _zz_2646);
  assign _zz_9473 = _zz_9474;
  assign _zz_9474 = ($signed(_zz_677) - $signed(_zz_2643));
  assign _zz_9475 = _zz_9476;
  assign _zz_9476 = ($signed(_zz_9477) >>> _zz_2646);
  assign _zz_9477 = _zz_9478;
  assign _zz_9478 = ($signed(_zz_678) - $signed(_zz_2644));
  assign _zz_9479 = _zz_9480;
  assign _zz_9480 = ($signed(_zz_9481) >>> _zz_2647);
  assign _zz_9481 = _zz_9482;
  assign _zz_9482 = ($signed(_zz_677) + $signed(_zz_2643));
  assign _zz_9483 = _zz_9484;
  assign _zz_9484 = ($signed(_zz_9485) >>> _zz_2647);
  assign _zz_9485 = _zz_9486;
  assign _zz_9486 = ($signed(_zz_678) + $signed(_zz_2644));
  assign _zz_9487 = ($signed(twiddle_factor_table_6_real) + $signed(twiddle_factor_table_6_imag));
  assign _zz_9488 = fixTo_513_dout;
  assign _zz_9489 = ($signed(_zz_688) - $signed(_zz_687));
  assign _zz_9490 = ($signed(_zz_687) + $signed(_zz_688));
  assign _zz_9491 = _zz_9492[15 : 0];
  assign _zz_9492 = fixTo_515_dout;
  assign _zz_9493 = _zz_9494[15 : 0];
  assign _zz_9494 = fixTo_514_dout;
  assign _zz_9495 = _zz_9496;
  assign _zz_9496 = ($signed(_zz_9497) >>> _zz_2651);
  assign _zz_9497 = _zz_9498;
  assign _zz_9498 = ($signed(_zz_679) - $signed(_zz_2648));
  assign _zz_9499 = _zz_9500;
  assign _zz_9500 = ($signed(_zz_9501) >>> _zz_2651);
  assign _zz_9501 = _zz_9502;
  assign _zz_9502 = ($signed(_zz_680) - $signed(_zz_2649));
  assign _zz_9503 = _zz_9504;
  assign _zz_9504 = ($signed(_zz_9505) >>> _zz_2652);
  assign _zz_9505 = _zz_9506;
  assign _zz_9506 = ($signed(_zz_679) + $signed(_zz_2648));
  assign _zz_9507 = _zz_9508;
  assign _zz_9508 = ($signed(_zz_9509) >>> _zz_2652);
  assign _zz_9509 = _zz_9510;
  assign _zz_9510 = ($signed(_zz_680) + $signed(_zz_2649));
  assign _zz_9511 = ($signed(twiddle_factor_table_3_real) + $signed(twiddle_factor_table_3_imag));
  assign _zz_9512 = fixTo_516_dout;
  assign _zz_9513 = ($signed(_zz_698) - $signed(_zz_697));
  assign _zz_9514 = ($signed(_zz_697) + $signed(_zz_698));
  assign _zz_9515 = _zz_9516[15 : 0];
  assign _zz_9516 = fixTo_518_dout;
  assign _zz_9517 = _zz_9518[15 : 0];
  assign _zz_9518 = fixTo_517_dout;
  assign _zz_9519 = _zz_9520;
  assign _zz_9520 = ($signed(_zz_9521) >>> _zz_2656);
  assign _zz_9521 = _zz_9522;
  assign _zz_9522 = ($signed(_zz_689) - $signed(_zz_2653));
  assign _zz_9523 = _zz_9524;
  assign _zz_9524 = ($signed(_zz_9525) >>> _zz_2656);
  assign _zz_9525 = _zz_9526;
  assign _zz_9526 = ($signed(_zz_690) - $signed(_zz_2654));
  assign _zz_9527 = _zz_9528;
  assign _zz_9528 = ($signed(_zz_9529) >>> _zz_2657);
  assign _zz_9529 = _zz_9530;
  assign _zz_9530 = ($signed(_zz_689) + $signed(_zz_2653));
  assign _zz_9531 = _zz_9532;
  assign _zz_9532 = ($signed(_zz_9533) >>> _zz_2657);
  assign _zz_9533 = _zz_9534;
  assign _zz_9534 = ($signed(_zz_690) + $signed(_zz_2654));
  assign _zz_9535 = ($signed(twiddle_factor_table_4_real) + $signed(twiddle_factor_table_4_imag));
  assign _zz_9536 = fixTo_519_dout;
  assign _zz_9537 = ($signed(_zz_700) - $signed(_zz_699));
  assign _zz_9538 = ($signed(_zz_699) + $signed(_zz_700));
  assign _zz_9539 = _zz_9540[15 : 0];
  assign _zz_9540 = fixTo_521_dout;
  assign _zz_9541 = _zz_9542[15 : 0];
  assign _zz_9542 = fixTo_520_dout;
  assign _zz_9543 = _zz_9544;
  assign _zz_9544 = ($signed(_zz_9545) >>> _zz_2661);
  assign _zz_9545 = _zz_9546;
  assign _zz_9546 = ($signed(_zz_691) - $signed(_zz_2658));
  assign _zz_9547 = _zz_9548;
  assign _zz_9548 = ($signed(_zz_9549) >>> _zz_2661);
  assign _zz_9549 = _zz_9550;
  assign _zz_9550 = ($signed(_zz_692) - $signed(_zz_2659));
  assign _zz_9551 = _zz_9552;
  assign _zz_9552 = ($signed(_zz_9553) >>> _zz_2662);
  assign _zz_9553 = _zz_9554;
  assign _zz_9554 = ($signed(_zz_691) + $signed(_zz_2658));
  assign _zz_9555 = _zz_9556;
  assign _zz_9556 = ($signed(_zz_9557) >>> _zz_2662);
  assign _zz_9557 = _zz_9558;
  assign _zz_9558 = ($signed(_zz_692) + $signed(_zz_2659));
  assign _zz_9559 = ($signed(twiddle_factor_table_5_real) + $signed(twiddle_factor_table_5_imag));
  assign _zz_9560 = fixTo_522_dout;
  assign _zz_9561 = ($signed(_zz_702) - $signed(_zz_701));
  assign _zz_9562 = ($signed(_zz_701) + $signed(_zz_702));
  assign _zz_9563 = _zz_9564[15 : 0];
  assign _zz_9564 = fixTo_524_dout;
  assign _zz_9565 = _zz_9566[15 : 0];
  assign _zz_9566 = fixTo_523_dout;
  assign _zz_9567 = _zz_9568;
  assign _zz_9568 = ($signed(_zz_9569) >>> _zz_2666);
  assign _zz_9569 = _zz_9570;
  assign _zz_9570 = ($signed(_zz_693) - $signed(_zz_2663));
  assign _zz_9571 = _zz_9572;
  assign _zz_9572 = ($signed(_zz_9573) >>> _zz_2666);
  assign _zz_9573 = _zz_9574;
  assign _zz_9574 = ($signed(_zz_694) - $signed(_zz_2664));
  assign _zz_9575 = _zz_9576;
  assign _zz_9576 = ($signed(_zz_9577) >>> _zz_2667);
  assign _zz_9577 = _zz_9578;
  assign _zz_9578 = ($signed(_zz_693) + $signed(_zz_2663));
  assign _zz_9579 = _zz_9580;
  assign _zz_9580 = ($signed(_zz_9581) >>> _zz_2667);
  assign _zz_9581 = _zz_9582;
  assign _zz_9582 = ($signed(_zz_694) + $signed(_zz_2664));
  assign _zz_9583 = ($signed(twiddle_factor_table_6_real) + $signed(twiddle_factor_table_6_imag));
  assign _zz_9584 = fixTo_525_dout;
  assign _zz_9585 = ($signed(_zz_704) - $signed(_zz_703));
  assign _zz_9586 = ($signed(_zz_703) + $signed(_zz_704));
  assign _zz_9587 = _zz_9588[15 : 0];
  assign _zz_9588 = fixTo_527_dout;
  assign _zz_9589 = _zz_9590[15 : 0];
  assign _zz_9590 = fixTo_526_dout;
  assign _zz_9591 = _zz_9592;
  assign _zz_9592 = ($signed(_zz_9593) >>> _zz_2671);
  assign _zz_9593 = _zz_9594;
  assign _zz_9594 = ($signed(_zz_695) - $signed(_zz_2668));
  assign _zz_9595 = _zz_9596;
  assign _zz_9596 = ($signed(_zz_9597) >>> _zz_2671);
  assign _zz_9597 = _zz_9598;
  assign _zz_9598 = ($signed(_zz_696) - $signed(_zz_2669));
  assign _zz_9599 = _zz_9600;
  assign _zz_9600 = ($signed(_zz_9601) >>> _zz_2672);
  assign _zz_9601 = _zz_9602;
  assign _zz_9602 = ($signed(_zz_695) + $signed(_zz_2668));
  assign _zz_9603 = _zz_9604;
  assign _zz_9604 = ($signed(_zz_9605) >>> _zz_2672);
  assign _zz_9605 = _zz_9606;
  assign _zz_9606 = ($signed(_zz_696) + $signed(_zz_2669));
  assign _zz_9607 = ($signed(twiddle_factor_table_3_real) + $signed(twiddle_factor_table_3_imag));
  assign _zz_9608 = fixTo_528_dout;
  assign _zz_9609 = ($signed(_zz_714) - $signed(_zz_713));
  assign _zz_9610 = ($signed(_zz_713) + $signed(_zz_714));
  assign _zz_9611 = _zz_9612[15 : 0];
  assign _zz_9612 = fixTo_530_dout;
  assign _zz_9613 = _zz_9614[15 : 0];
  assign _zz_9614 = fixTo_529_dout;
  assign _zz_9615 = _zz_9616;
  assign _zz_9616 = ($signed(_zz_9617) >>> _zz_2676);
  assign _zz_9617 = _zz_9618;
  assign _zz_9618 = ($signed(_zz_705) - $signed(_zz_2673));
  assign _zz_9619 = _zz_9620;
  assign _zz_9620 = ($signed(_zz_9621) >>> _zz_2676);
  assign _zz_9621 = _zz_9622;
  assign _zz_9622 = ($signed(_zz_706) - $signed(_zz_2674));
  assign _zz_9623 = _zz_9624;
  assign _zz_9624 = ($signed(_zz_9625) >>> _zz_2677);
  assign _zz_9625 = _zz_9626;
  assign _zz_9626 = ($signed(_zz_705) + $signed(_zz_2673));
  assign _zz_9627 = _zz_9628;
  assign _zz_9628 = ($signed(_zz_9629) >>> _zz_2677);
  assign _zz_9629 = _zz_9630;
  assign _zz_9630 = ($signed(_zz_706) + $signed(_zz_2674));
  assign _zz_9631 = ($signed(twiddle_factor_table_4_real) + $signed(twiddle_factor_table_4_imag));
  assign _zz_9632 = fixTo_531_dout;
  assign _zz_9633 = ($signed(_zz_716) - $signed(_zz_715));
  assign _zz_9634 = ($signed(_zz_715) + $signed(_zz_716));
  assign _zz_9635 = _zz_9636[15 : 0];
  assign _zz_9636 = fixTo_533_dout;
  assign _zz_9637 = _zz_9638[15 : 0];
  assign _zz_9638 = fixTo_532_dout;
  assign _zz_9639 = _zz_9640;
  assign _zz_9640 = ($signed(_zz_9641) >>> _zz_2681);
  assign _zz_9641 = _zz_9642;
  assign _zz_9642 = ($signed(_zz_707) - $signed(_zz_2678));
  assign _zz_9643 = _zz_9644;
  assign _zz_9644 = ($signed(_zz_9645) >>> _zz_2681);
  assign _zz_9645 = _zz_9646;
  assign _zz_9646 = ($signed(_zz_708) - $signed(_zz_2679));
  assign _zz_9647 = _zz_9648;
  assign _zz_9648 = ($signed(_zz_9649) >>> _zz_2682);
  assign _zz_9649 = _zz_9650;
  assign _zz_9650 = ($signed(_zz_707) + $signed(_zz_2678));
  assign _zz_9651 = _zz_9652;
  assign _zz_9652 = ($signed(_zz_9653) >>> _zz_2682);
  assign _zz_9653 = _zz_9654;
  assign _zz_9654 = ($signed(_zz_708) + $signed(_zz_2679));
  assign _zz_9655 = ($signed(twiddle_factor_table_5_real) + $signed(twiddle_factor_table_5_imag));
  assign _zz_9656 = fixTo_534_dout;
  assign _zz_9657 = ($signed(_zz_718) - $signed(_zz_717));
  assign _zz_9658 = ($signed(_zz_717) + $signed(_zz_718));
  assign _zz_9659 = _zz_9660[15 : 0];
  assign _zz_9660 = fixTo_536_dout;
  assign _zz_9661 = _zz_9662[15 : 0];
  assign _zz_9662 = fixTo_535_dout;
  assign _zz_9663 = _zz_9664;
  assign _zz_9664 = ($signed(_zz_9665) >>> _zz_2686);
  assign _zz_9665 = _zz_9666;
  assign _zz_9666 = ($signed(_zz_709) - $signed(_zz_2683));
  assign _zz_9667 = _zz_9668;
  assign _zz_9668 = ($signed(_zz_9669) >>> _zz_2686);
  assign _zz_9669 = _zz_9670;
  assign _zz_9670 = ($signed(_zz_710) - $signed(_zz_2684));
  assign _zz_9671 = _zz_9672;
  assign _zz_9672 = ($signed(_zz_9673) >>> _zz_2687);
  assign _zz_9673 = _zz_9674;
  assign _zz_9674 = ($signed(_zz_709) + $signed(_zz_2683));
  assign _zz_9675 = _zz_9676;
  assign _zz_9676 = ($signed(_zz_9677) >>> _zz_2687);
  assign _zz_9677 = _zz_9678;
  assign _zz_9678 = ($signed(_zz_710) + $signed(_zz_2684));
  assign _zz_9679 = ($signed(twiddle_factor_table_6_real) + $signed(twiddle_factor_table_6_imag));
  assign _zz_9680 = fixTo_537_dout;
  assign _zz_9681 = ($signed(_zz_720) - $signed(_zz_719));
  assign _zz_9682 = ($signed(_zz_719) + $signed(_zz_720));
  assign _zz_9683 = _zz_9684[15 : 0];
  assign _zz_9684 = fixTo_539_dout;
  assign _zz_9685 = _zz_9686[15 : 0];
  assign _zz_9686 = fixTo_538_dout;
  assign _zz_9687 = _zz_9688;
  assign _zz_9688 = ($signed(_zz_9689) >>> _zz_2691);
  assign _zz_9689 = _zz_9690;
  assign _zz_9690 = ($signed(_zz_711) - $signed(_zz_2688));
  assign _zz_9691 = _zz_9692;
  assign _zz_9692 = ($signed(_zz_9693) >>> _zz_2691);
  assign _zz_9693 = _zz_9694;
  assign _zz_9694 = ($signed(_zz_712) - $signed(_zz_2689));
  assign _zz_9695 = _zz_9696;
  assign _zz_9696 = ($signed(_zz_9697) >>> _zz_2692);
  assign _zz_9697 = _zz_9698;
  assign _zz_9698 = ($signed(_zz_711) + $signed(_zz_2688));
  assign _zz_9699 = _zz_9700;
  assign _zz_9700 = ($signed(_zz_9701) >>> _zz_2692);
  assign _zz_9701 = _zz_9702;
  assign _zz_9702 = ($signed(_zz_712) + $signed(_zz_2689));
  assign _zz_9703 = ($signed(twiddle_factor_table_3_real) + $signed(twiddle_factor_table_3_imag));
  assign _zz_9704 = fixTo_540_dout;
  assign _zz_9705 = ($signed(_zz_730) - $signed(_zz_729));
  assign _zz_9706 = ($signed(_zz_729) + $signed(_zz_730));
  assign _zz_9707 = _zz_9708[15 : 0];
  assign _zz_9708 = fixTo_542_dout;
  assign _zz_9709 = _zz_9710[15 : 0];
  assign _zz_9710 = fixTo_541_dout;
  assign _zz_9711 = _zz_9712;
  assign _zz_9712 = ($signed(_zz_9713) >>> _zz_2696);
  assign _zz_9713 = _zz_9714;
  assign _zz_9714 = ($signed(_zz_721) - $signed(_zz_2693));
  assign _zz_9715 = _zz_9716;
  assign _zz_9716 = ($signed(_zz_9717) >>> _zz_2696);
  assign _zz_9717 = _zz_9718;
  assign _zz_9718 = ($signed(_zz_722) - $signed(_zz_2694));
  assign _zz_9719 = _zz_9720;
  assign _zz_9720 = ($signed(_zz_9721) >>> _zz_2697);
  assign _zz_9721 = _zz_9722;
  assign _zz_9722 = ($signed(_zz_721) + $signed(_zz_2693));
  assign _zz_9723 = _zz_9724;
  assign _zz_9724 = ($signed(_zz_9725) >>> _zz_2697);
  assign _zz_9725 = _zz_9726;
  assign _zz_9726 = ($signed(_zz_722) + $signed(_zz_2694));
  assign _zz_9727 = ($signed(twiddle_factor_table_4_real) + $signed(twiddle_factor_table_4_imag));
  assign _zz_9728 = fixTo_543_dout;
  assign _zz_9729 = ($signed(_zz_732) - $signed(_zz_731));
  assign _zz_9730 = ($signed(_zz_731) + $signed(_zz_732));
  assign _zz_9731 = _zz_9732[15 : 0];
  assign _zz_9732 = fixTo_545_dout;
  assign _zz_9733 = _zz_9734[15 : 0];
  assign _zz_9734 = fixTo_544_dout;
  assign _zz_9735 = _zz_9736;
  assign _zz_9736 = ($signed(_zz_9737) >>> _zz_2701);
  assign _zz_9737 = _zz_9738;
  assign _zz_9738 = ($signed(_zz_723) - $signed(_zz_2698));
  assign _zz_9739 = _zz_9740;
  assign _zz_9740 = ($signed(_zz_9741) >>> _zz_2701);
  assign _zz_9741 = _zz_9742;
  assign _zz_9742 = ($signed(_zz_724) - $signed(_zz_2699));
  assign _zz_9743 = _zz_9744;
  assign _zz_9744 = ($signed(_zz_9745) >>> _zz_2702);
  assign _zz_9745 = _zz_9746;
  assign _zz_9746 = ($signed(_zz_723) + $signed(_zz_2698));
  assign _zz_9747 = _zz_9748;
  assign _zz_9748 = ($signed(_zz_9749) >>> _zz_2702);
  assign _zz_9749 = _zz_9750;
  assign _zz_9750 = ($signed(_zz_724) + $signed(_zz_2699));
  assign _zz_9751 = ($signed(twiddle_factor_table_5_real) + $signed(twiddle_factor_table_5_imag));
  assign _zz_9752 = fixTo_546_dout;
  assign _zz_9753 = ($signed(_zz_734) - $signed(_zz_733));
  assign _zz_9754 = ($signed(_zz_733) + $signed(_zz_734));
  assign _zz_9755 = _zz_9756[15 : 0];
  assign _zz_9756 = fixTo_548_dout;
  assign _zz_9757 = _zz_9758[15 : 0];
  assign _zz_9758 = fixTo_547_dout;
  assign _zz_9759 = _zz_9760;
  assign _zz_9760 = ($signed(_zz_9761) >>> _zz_2706);
  assign _zz_9761 = _zz_9762;
  assign _zz_9762 = ($signed(_zz_725) - $signed(_zz_2703));
  assign _zz_9763 = _zz_9764;
  assign _zz_9764 = ($signed(_zz_9765) >>> _zz_2706);
  assign _zz_9765 = _zz_9766;
  assign _zz_9766 = ($signed(_zz_726) - $signed(_zz_2704));
  assign _zz_9767 = _zz_9768;
  assign _zz_9768 = ($signed(_zz_9769) >>> _zz_2707);
  assign _zz_9769 = _zz_9770;
  assign _zz_9770 = ($signed(_zz_725) + $signed(_zz_2703));
  assign _zz_9771 = _zz_9772;
  assign _zz_9772 = ($signed(_zz_9773) >>> _zz_2707);
  assign _zz_9773 = _zz_9774;
  assign _zz_9774 = ($signed(_zz_726) + $signed(_zz_2704));
  assign _zz_9775 = ($signed(twiddle_factor_table_6_real) + $signed(twiddle_factor_table_6_imag));
  assign _zz_9776 = fixTo_549_dout;
  assign _zz_9777 = ($signed(_zz_736) - $signed(_zz_735));
  assign _zz_9778 = ($signed(_zz_735) + $signed(_zz_736));
  assign _zz_9779 = _zz_9780[15 : 0];
  assign _zz_9780 = fixTo_551_dout;
  assign _zz_9781 = _zz_9782[15 : 0];
  assign _zz_9782 = fixTo_550_dout;
  assign _zz_9783 = _zz_9784;
  assign _zz_9784 = ($signed(_zz_9785) >>> _zz_2711);
  assign _zz_9785 = _zz_9786;
  assign _zz_9786 = ($signed(_zz_727) - $signed(_zz_2708));
  assign _zz_9787 = _zz_9788;
  assign _zz_9788 = ($signed(_zz_9789) >>> _zz_2711);
  assign _zz_9789 = _zz_9790;
  assign _zz_9790 = ($signed(_zz_728) - $signed(_zz_2709));
  assign _zz_9791 = _zz_9792;
  assign _zz_9792 = ($signed(_zz_9793) >>> _zz_2712);
  assign _zz_9793 = _zz_9794;
  assign _zz_9794 = ($signed(_zz_727) + $signed(_zz_2708));
  assign _zz_9795 = _zz_9796;
  assign _zz_9796 = ($signed(_zz_9797) >>> _zz_2712);
  assign _zz_9797 = _zz_9798;
  assign _zz_9798 = ($signed(_zz_728) + $signed(_zz_2709));
  assign _zz_9799 = ($signed(twiddle_factor_table_3_real) + $signed(twiddle_factor_table_3_imag));
  assign _zz_9800 = fixTo_552_dout;
  assign _zz_9801 = ($signed(_zz_746) - $signed(_zz_745));
  assign _zz_9802 = ($signed(_zz_745) + $signed(_zz_746));
  assign _zz_9803 = _zz_9804[15 : 0];
  assign _zz_9804 = fixTo_554_dout;
  assign _zz_9805 = _zz_9806[15 : 0];
  assign _zz_9806 = fixTo_553_dout;
  assign _zz_9807 = _zz_9808;
  assign _zz_9808 = ($signed(_zz_9809) >>> _zz_2716);
  assign _zz_9809 = _zz_9810;
  assign _zz_9810 = ($signed(_zz_737) - $signed(_zz_2713));
  assign _zz_9811 = _zz_9812;
  assign _zz_9812 = ($signed(_zz_9813) >>> _zz_2716);
  assign _zz_9813 = _zz_9814;
  assign _zz_9814 = ($signed(_zz_738) - $signed(_zz_2714));
  assign _zz_9815 = _zz_9816;
  assign _zz_9816 = ($signed(_zz_9817) >>> _zz_2717);
  assign _zz_9817 = _zz_9818;
  assign _zz_9818 = ($signed(_zz_737) + $signed(_zz_2713));
  assign _zz_9819 = _zz_9820;
  assign _zz_9820 = ($signed(_zz_9821) >>> _zz_2717);
  assign _zz_9821 = _zz_9822;
  assign _zz_9822 = ($signed(_zz_738) + $signed(_zz_2714));
  assign _zz_9823 = ($signed(twiddle_factor_table_4_real) + $signed(twiddle_factor_table_4_imag));
  assign _zz_9824 = fixTo_555_dout;
  assign _zz_9825 = ($signed(_zz_748) - $signed(_zz_747));
  assign _zz_9826 = ($signed(_zz_747) + $signed(_zz_748));
  assign _zz_9827 = _zz_9828[15 : 0];
  assign _zz_9828 = fixTo_557_dout;
  assign _zz_9829 = _zz_9830[15 : 0];
  assign _zz_9830 = fixTo_556_dout;
  assign _zz_9831 = _zz_9832;
  assign _zz_9832 = ($signed(_zz_9833) >>> _zz_2721);
  assign _zz_9833 = _zz_9834;
  assign _zz_9834 = ($signed(_zz_739) - $signed(_zz_2718));
  assign _zz_9835 = _zz_9836;
  assign _zz_9836 = ($signed(_zz_9837) >>> _zz_2721);
  assign _zz_9837 = _zz_9838;
  assign _zz_9838 = ($signed(_zz_740) - $signed(_zz_2719));
  assign _zz_9839 = _zz_9840;
  assign _zz_9840 = ($signed(_zz_9841) >>> _zz_2722);
  assign _zz_9841 = _zz_9842;
  assign _zz_9842 = ($signed(_zz_739) + $signed(_zz_2718));
  assign _zz_9843 = _zz_9844;
  assign _zz_9844 = ($signed(_zz_9845) >>> _zz_2722);
  assign _zz_9845 = _zz_9846;
  assign _zz_9846 = ($signed(_zz_740) + $signed(_zz_2719));
  assign _zz_9847 = ($signed(twiddle_factor_table_5_real) + $signed(twiddle_factor_table_5_imag));
  assign _zz_9848 = fixTo_558_dout;
  assign _zz_9849 = ($signed(_zz_750) - $signed(_zz_749));
  assign _zz_9850 = ($signed(_zz_749) + $signed(_zz_750));
  assign _zz_9851 = _zz_9852[15 : 0];
  assign _zz_9852 = fixTo_560_dout;
  assign _zz_9853 = _zz_9854[15 : 0];
  assign _zz_9854 = fixTo_559_dout;
  assign _zz_9855 = _zz_9856;
  assign _zz_9856 = ($signed(_zz_9857) >>> _zz_2726);
  assign _zz_9857 = _zz_9858;
  assign _zz_9858 = ($signed(_zz_741) - $signed(_zz_2723));
  assign _zz_9859 = _zz_9860;
  assign _zz_9860 = ($signed(_zz_9861) >>> _zz_2726);
  assign _zz_9861 = _zz_9862;
  assign _zz_9862 = ($signed(_zz_742) - $signed(_zz_2724));
  assign _zz_9863 = _zz_9864;
  assign _zz_9864 = ($signed(_zz_9865) >>> _zz_2727);
  assign _zz_9865 = _zz_9866;
  assign _zz_9866 = ($signed(_zz_741) + $signed(_zz_2723));
  assign _zz_9867 = _zz_9868;
  assign _zz_9868 = ($signed(_zz_9869) >>> _zz_2727);
  assign _zz_9869 = _zz_9870;
  assign _zz_9870 = ($signed(_zz_742) + $signed(_zz_2724));
  assign _zz_9871 = ($signed(twiddle_factor_table_6_real) + $signed(twiddle_factor_table_6_imag));
  assign _zz_9872 = fixTo_561_dout;
  assign _zz_9873 = ($signed(_zz_752) - $signed(_zz_751));
  assign _zz_9874 = ($signed(_zz_751) + $signed(_zz_752));
  assign _zz_9875 = _zz_9876[15 : 0];
  assign _zz_9876 = fixTo_563_dout;
  assign _zz_9877 = _zz_9878[15 : 0];
  assign _zz_9878 = fixTo_562_dout;
  assign _zz_9879 = _zz_9880;
  assign _zz_9880 = ($signed(_zz_9881) >>> _zz_2731);
  assign _zz_9881 = _zz_9882;
  assign _zz_9882 = ($signed(_zz_743) - $signed(_zz_2728));
  assign _zz_9883 = _zz_9884;
  assign _zz_9884 = ($signed(_zz_9885) >>> _zz_2731);
  assign _zz_9885 = _zz_9886;
  assign _zz_9886 = ($signed(_zz_744) - $signed(_zz_2729));
  assign _zz_9887 = _zz_9888;
  assign _zz_9888 = ($signed(_zz_9889) >>> _zz_2732);
  assign _zz_9889 = _zz_9890;
  assign _zz_9890 = ($signed(_zz_743) + $signed(_zz_2728));
  assign _zz_9891 = _zz_9892;
  assign _zz_9892 = ($signed(_zz_9893) >>> _zz_2732);
  assign _zz_9893 = _zz_9894;
  assign _zz_9894 = ($signed(_zz_744) + $signed(_zz_2729));
  assign _zz_9895 = ($signed(twiddle_factor_table_3_real) + $signed(twiddle_factor_table_3_imag));
  assign _zz_9896 = fixTo_564_dout;
  assign _zz_9897 = ($signed(_zz_762) - $signed(_zz_761));
  assign _zz_9898 = ($signed(_zz_761) + $signed(_zz_762));
  assign _zz_9899 = _zz_9900[15 : 0];
  assign _zz_9900 = fixTo_566_dout;
  assign _zz_9901 = _zz_9902[15 : 0];
  assign _zz_9902 = fixTo_565_dout;
  assign _zz_9903 = _zz_9904;
  assign _zz_9904 = ($signed(_zz_9905) >>> _zz_2736);
  assign _zz_9905 = _zz_9906;
  assign _zz_9906 = ($signed(_zz_753) - $signed(_zz_2733));
  assign _zz_9907 = _zz_9908;
  assign _zz_9908 = ($signed(_zz_9909) >>> _zz_2736);
  assign _zz_9909 = _zz_9910;
  assign _zz_9910 = ($signed(_zz_754) - $signed(_zz_2734));
  assign _zz_9911 = _zz_9912;
  assign _zz_9912 = ($signed(_zz_9913) >>> _zz_2737);
  assign _zz_9913 = _zz_9914;
  assign _zz_9914 = ($signed(_zz_753) + $signed(_zz_2733));
  assign _zz_9915 = _zz_9916;
  assign _zz_9916 = ($signed(_zz_9917) >>> _zz_2737);
  assign _zz_9917 = _zz_9918;
  assign _zz_9918 = ($signed(_zz_754) + $signed(_zz_2734));
  assign _zz_9919 = ($signed(twiddle_factor_table_4_real) + $signed(twiddle_factor_table_4_imag));
  assign _zz_9920 = fixTo_567_dout;
  assign _zz_9921 = ($signed(_zz_764) - $signed(_zz_763));
  assign _zz_9922 = ($signed(_zz_763) + $signed(_zz_764));
  assign _zz_9923 = _zz_9924[15 : 0];
  assign _zz_9924 = fixTo_569_dout;
  assign _zz_9925 = _zz_9926[15 : 0];
  assign _zz_9926 = fixTo_568_dout;
  assign _zz_9927 = _zz_9928;
  assign _zz_9928 = ($signed(_zz_9929) >>> _zz_2741);
  assign _zz_9929 = _zz_9930;
  assign _zz_9930 = ($signed(_zz_755) - $signed(_zz_2738));
  assign _zz_9931 = _zz_9932;
  assign _zz_9932 = ($signed(_zz_9933) >>> _zz_2741);
  assign _zz_9933 = _zz_9934;
  assign _zz_9934 = ($signed(_zz_756) - $signed(_zz_2739));
  assign _zz_9935 = _zz_9936;
  assign _zz_9936 = ($signed(_zz_9937) >>> _zz_2742);
  assign _zz_9937 = _zz_9938;
  assign _zz_9938 = ($signed(_zz_755) + $signed(_zz_2738));
  assign _zz_9939 = _zz_9940;
  assign _zz_9940 = ($signed(_zz_9941) >>> _zz_2742);
  assign _zz_9941 = _zz_9942;
  assign _zz_9942 = ($signed(_zz_756) + $signed(_zz_2739));
  assign _zz_9943 = ($signed(twiddle_factor_table_5_real) + $signed(twiddle_factor_table_5_imag));
  assign _zz_9944 = fixTo_570_dout;
  assign _zz_9945 = ($signed(_zz_766) - $signed(_zz_765));
  assign _zz_9946 = ($signed(_zz_765) + $signed(_zz_766));
  assign _zz_9947 = _zz_9948[15 : 0];
  assign _zz_9948 = fixTo_572_dout;
  assign _zz_9949 = _zz_9950[15 : 0];
  assign _zz_9950 = fixTo_571_dout;
  assign _zz_9951 = _zz_9952;
  assign _zz_9952 = ($signed(_zz_9953) >>> _zz_2746);
  assign _zz_9953 = _zz_9954;
  assign _zz_9954 = ($signed(_zz_757) - $signed(_zz_2743));
  assign _zz_9955 = _zz_9956;
  assign _zz_9956 = ($signed(_zz_9957) >>> _zz_2746);
  assign _zz_9957 = _zz_9958;
  assign _zz_9958 = ($signed(_zz_758) - $signed(_zz_2744));
  assign _zz_9959 = _zz_9960;
  assign _zz_9960 = ($signed(_zz_9961) >>> _zz_2747);
  assign _zz_9961 = _zz_9962;
  assign _zz_9962 = ($signed(_zz_757) + $signed(_zz_2743));
  assign _zz_9963 = _zz_9964;
  assign _zz_9964 = ($signed(_zz_9965) >>> _zz_2747);
  assign _zz_9965 = _zz_9966;
  assign _zz_9966 = ($signed(_zz_758) + $signed(_zz_2744));
  assign _zz_9967 = ($signed(twiddle_factor_table_6_real) + $signed(twiddle_factor_table_6_imag));
  assign _zz_9968 = fixTo_573_dout;
  assign _zz_9969 = ($signed(_zz_768) - $signed(_zz_767));
  assign _zz_9970 = ($signed(_zz_767) + $signed(_zz_768));
  assign _zz_9971 = _zz_9972[15 : 0];
  assign _zz_9972 = fixTo_575_dout;
  assign _zz_9973 = _zz_9974[15 : 0];
  assign _zz_9974 = fixTo_574_dout;
  assign _zz_9975 = _zz_9976;
  assign _zz_9976 = ($signed(_zz_9977) >>> _zz_2751);
  assign _zz_9977 = _zz_9978;
  assign _zz_9978 = ($signed(_zz_759) - $signed(_zz_2748));
  assign _zz_9979 = _zz_9980;
  assign _zz_9980 = ($signed(_zz_9981) >>> _zz_2751);
  assign _zz_9981 = _zz_9982;
  assign _zz_9982 = ($signed(_zz_760) - $signed(_zz_2749));
  assign _zz_9983 = _zz_9984;
  assign _zz_9984 = ($signed(_zz_9985) >>> _zz_2752);
  assign _zz_9985 = _zz_9986;
  assign _zz_9986 = ($signed(_zz_759) + $signed(_zz_2748));
  assign _zz_9987 = _zz_9988;
  assign _zz_9988 = ($signed(_zz_9989) >>> _zz_2752);
  assign _zz_9989 = _zz_9990;
  assign _zz_9990 = ($signed(_zz_760) + $signed(_zz_2749));
  assign _zz_9991 = ($signed(twiddle_factor_table_7_real) + $signed(twiddle_factor_table_7_imag));
  assign _zz_9992 = fixTo_576_dout;
  assign _zz_9993 = ($signed(_zz_786) - $signed(_zz_785));
  assign _zz_9994 = ($signed(_zz_785) + $signed(_zz_786));
  assign _zz_9995 = _zz_9996[15 : 0];
  assign _zz_9996 = fixTo_578_dout;
  assign _zz_9997 = _zz_9998[15 : 0];
  assign _zz_9998 = fixTo_577_dout;
  assign _zz_9999 = _zz_10000;
  assign _zz_10000 = ($signed(_zz_10001) >>> _zz_2756);
  assign _zz_10001 = _zz_10002;
  assign _zz_10002 = ($signed(_zz_769) - $signed(_zz_2753));
  assign _zz_10003 = _zz_10004;
  assign _zz_10004 = ($signed(_zz_10005) >>> _zz_2756);
  assign _zz_10005 = _zz_10006;
  assign _zz_10006 = ($signed(_zz_770) - $signed(_zz_2754));
  assign _zz_10007 = _zz_10008;
  assign _zz_10008 = ($signed(_zz_10009) >>> _zz_2757);
  assign _zz_10009 = _zz_10010;
  assign _zz_10010 = ($signed(_zz_769) + $signed(_zz_2753));
  assign _zz_10011 = _zz_10012;
  assign _zz_10012 = ($signed(_zz_10013) >>> _zz_2757);
  assign _zz_10013 = _zz_10014;
  assign _zz_10014 = ($signed(_zz_770) + $signed(_zz_2754));
  assign _zz_10015 = ($signed(twiddle_factor_table_8_real) + $signed(twiddle_factor_table_8_imag));
  assign _zz_10016 = fixTo_579_dout;
  assign _zz_10017 = ($signed(_zz_788) - $signed(_zz_787));
  assign _zz_10018 = ($signed(_zz_787) + $signed(_zz_788));
  assign _zz_10019 = _zz_10020[15 : 0];
  assign _zz_10020 = fixTo_581_dout;
  assign _zz_10021 = _zz_10022[15 : 0];
  assign _zz_10022 = fixTo_580_dout;
  assign _zz_10023 = _zz_10024;
  assign _zz_10024 = ($signed(_zz_10025) >>> _zz_2761);
  assign _zz_10025 = _zz_10026;
  assign _zz_10026 = ($signed(_zz_771) - $signed(_zz_2758));
  assign _zz_10027 = _zz_10028;
  assign _zz_10028 = ($signed(_zz_10029) >>> _zz_2761);
  assign _zz_10029 = _zz_10030;
  assign _zz_10030 = ($signed(_zz_772) - $signed(_zz_2759));
  assign _zz_10031 = _zz_10032;
  assign _zz_10032 = ($signed(_zz_10033) >>> _zz_2762);
  assign _zz_10033 = _zz_10034;
  assign _zz_10034 = ($signed(_zz_771) + $signed(_zz_2758));
  assign _zz_10035 = _zz_10036;
  assign _zz_10036 = ($signed(_zz_10037) >>> _zz_2762);
  assign _zz_10037 = _zz_10038;
  assign _zz_10038 = ($signed(_zz_772) + $signed(_zz_2759));
  assign _zz_10039 = ($signed(twiddle_factor_table_9_real) + $signed(twiddle_factor_table_9_imag));
  assign _zz_10040 = fixTo_582_dout;
  assign _zz_10041 = ($signed(_zz_790) - $signed(_zz_789));
  assign _zz_10042 = ($signed(_zz_789) + $signed(_zz_790));
  assign _zz_10043 = _zz_10044[15 : 0];
  assign _zz_10044 = fixTo_584_dout;
  assign _zz_10045 = _zz_10046[15 : 0];
  assign _zz_10046 = fixTo_583_dout;
  assign _zz_10047 = _zz_10048;
  assign _zz_10048 = ($signed(_zz_10049) >>> _zz_2766);
  assign _zz_10049 = _zz_10050;
  assign _zz_10050 = ($signed(_zz_773) - $signed(_zz_2763));
  assign _zz_10051 = _zz_10052;
  assign _zz_10052 = ($signed(_zz_10053) >>> _zz_2766);
  assign _zz_10053 = _zz_10054;
  assign _zz_10054 = ($signed(_zz_774) - $signed(_zz_2764));
  assign _zz_10055 = _zz_10056;
  assign _zz_10056 = ($signed(_zz_10057) >>> _zz_2767);
  assign _zz_10057 = _zz_10058;
  assign _zz_10058 = ($signed(_zz_773) + $signed(_zz_2763));
  assign _zz_10059 = _zz_10060;
  assign _zz_10060 = ($signed(_zz_10061) >>> _zz_2767);
  assign _zz_10061 = _zz_10062;
  assign _zz_10062 = ($signed(_zz_774) + $signed(_zz_2764));
  assign _zz_10063 = ($signed(twiddle_factor_table_10_real) + $signed(twiddle_factor_table_10_imag));
  assign _zz_10064 = fixTo_585_dout;
  assign _zz_10065 = ($signed(_zz_792) - $signed(_zz_791));
  assign _zz_10066 = ($signed(_zz_791) + $signed(_zz_792));
  assign _zz_10067 = _zz_10068[15 : 0];
  assign _zz_10068 = fixTo_587_dout;
  assign _zz_10069 = _zz_10070[15 : 0];
  assign _zz_10070 = fixTo_586_dout;
  assign _zz_10071 = _zz_10072;
  assign _zz_10072 = ($signed(_zz_10073) >>> _zz_2771);
  assign _zz_10073 = _zz_10074;
  assign _zz_10074 = ($signed(_zz_775) - $signed(_zz_2768));
  assign _zz_10075 = _zz_10076;
  assign _zz_10076 = ($signed(_zz_10077) >>> _zz_2771);
  assign _zz_10077 = _zz_10078;
  assign _zz_10078 = ($signed(_zz_776) - $signed(_zz_2769));
  assign _zz_10079 = _zz_10080;
  assign _zz_10080 = ($signed(_zz_10081) >>> _zz_2772);
  assign _zz_10081 = _zz_10082;
  assign _zz_10082 = ($signed(_zz_775) + $signed(_zz_2768));
  assign _zz_10083 = _zz_10084;
  assign _zz_10084 = ($signed(_zz_10085) >>> _zz_2772);
  assign _zz_10085 = _zz_10086;
  assign _zz_10086 = ($signed(_zz_776) + $signed(_zz_2769));
  assign _zz_10087 = ($signed(twiddle_factor_table_11_real) + $signed(twiddle_factor_table_11_imag));
  assign _zz_10088 = fixTo_588_dout;
  assign _zz_10089 = ($signed(_zz_794) - $signed(_zz_793));
  assign _zz_10090 = ($signed(_zz_793) + $signed(_zz_794));
  assign _zz_10091 = _zz_10092[15 : 0];
  assign _zz_10092 = fixTo_590_dout;
  assign _zz_10093 = _zz_10094[15 : 0];
  assign _zz_10094 = fixTo_589_dout;
  assign _zz_10095 = _zz_10096;
  assign _zz_10096 = ($signed(_zz_10097) >>> _zz_2776);
  assign _zz_10097 = _zz_10098;
  assign _zz_10098 = ($signed(_zz_777) - $signed(_zz_2773));
  assign _zz_10099 = _zz_10100;
  assign _zz_10100 = ($signed(_zz_10101) >>> _zz_2776);
  assign _zz_10101 = _zz_10102;
  assign _zz_10102 = ($signed(_zz_778) - $signed(_zz_2774));
  assign _zz_10103 = _zz_10104;
  assign _zz_10104 = ($signed(_zz_10105) >>> _zz_2777);
  assign _zz_10105 = _zz_10106;
  assign _zz_10106 = ($signed(_zz_777) + $signed(_zz_2773));
  assign _zz_10107 = _zz_10108;
  assign _zz_10108 = ($signed(_zz_10109) >>> _zz_2777);
  assign _zz_10109 = _zz_10110;
  assign _zz_10110 = ($signed(_zz_778) + $signed(_zz_2774));
  assign _zz_10111 = ($signed(twiddle_factor_table_12_real) + $signed(twiddle_factor_table_12_imag));
  assign _zz_10112 = fixTo_591_dout;
  assign _zz_10113 = ($signed(_zz_796) - $signed(_zz_795));
  assign _zz_10114 = ($signed(_zz_795) + $signed(_zz_796));
  assign _zz_10115 = _zz_10116[15 : 0];
  assign _zz_10116 = fixTo_593_dout;
  assign _zz_10117 = _zz_10118[15 : 0];
  assign _zz_10118 = fixTo_592_dout;
  assign _zz_10119 = _zz_10120;
  assign _zz_10120 = ($signed(_zz_10121) >>> _zz_2781);
  assign _zz_10121 = _zz_10122;
  assign _zz_10122 = ($signed(_zz_779) - $signed(_zz_2778));
  assign _zz_10123 = _zz_10124;
  assign _zz_10124 = ($signed(_zz_10125) >>> _zz_2781);
  assign _zz_10125 = _zz_10126;
  assign _zz_10126 = ($signed(_zz_780) - $signed(_zz_2779));
  assign _zz_10127 = _zz_10128;
  assign _zz_10128 = ($signed(_zz_10129) >>> _zz_2782);
  assign _zz_10129 = _zz_10130;
  assign _zz_10130 = ($signed(_zz_779) + $signed(_zz_2778));
  assign _zz_10131 = _zz_10132;
  assign _zz_10132 = ($signed(_zz_10133) >>> _zz_2782);
  assign _zz_10133 = _zz_10134;
  assign _zz_10134 = ($signed(_zz_780) + $signed(_zz_2779));
  assign _zz_10135 = ($signed(twiddle_factor_table_13_real) + $signed(twiddle_factor_table_13_imag));
  assign _zz_10136 = fixTo_594_dout;
  assign _zz_10137 = ($signed(_zz_798) - $signed(_zz_797));
  assign _zz_10138 = ($signed(_zz_797) + $signed(_zz_798));
  assign _zz_10139 = _zz_10140[15 : 0];
  assign _zz_10140 = fixTo_596_dout;
  assign _zz_10141 = _zz_10142[15 : 0];
  assign _zz_10142 = fixTo_595_dout;
  assign _zz_10143 = _zz_10144;
  assign _zz_10144 = ($signed(_zz_10145) >>> _zz_2786);
  assign _zz_10145 = _zz_10146;
  assign _zz_10146 = ($signed(_zz_781) - $signed(_zz_2783));
  assign _zz_10147 = _zz_10148;
  assign _zz_10148 = ($signed(_zz_10149) >>> _zz_2786);
  assign _zz_10149 = _zz_10150;
  assign _zz_10150 = ($signed(_zz_782) - $signed(_zz_2784));
  assign _zz_10151 = _zz_10152;
  assign _zz_10152 = ($signed(_zz_10153) >>> _zz_2787);
  assign _zz_10153 = _zz_10154;
  assign _zz_10154 = ($signed(_zz_781) + $signed(_zz_2783));
  assign _zz_10155 = _zz_10156;
  assign _zz_10156 = ($signed(_zz_10157) >>> _zz_2787);
  assign _zz_10157 = _zz_10158;
  assign _zz_10158 = ($signed(_zz_782) + $signed(_zz_2784));
  assign _zz_10159 = ($signed(twiddle_factor_table_14_real) + $signed(twiddle_factor_table_14_imag));
  assign _zz_10160 = fixTo_597_dout;
  assign _zz_10161 = ($signed(_zz_800) - $signed(_zz_799));
  assign _zz_10162 = ($signed(_zz_799) + $signed(_zz_800));
  assign _zz_10163 = _zz_10164[15 : 0];
  assign _zz_10164 = fixTo_599_dout;
  assign _zz_10165 = _zz_10166[15 : 0];
  assign _zz_10166 = fixTo_598_dout;
  assign _zz_10167 = _zz_10168;
  assign _zz_10168 = ($signed(_zz_10169) >>> _zz_2791);
  assign _zz_10169 = _zz_10170;
  assign _zz_10170 = ($signed(_zz_783) - $signed(_zz_2788));
  assign _zz_10171 = _zz_10172;
  assign _zz_10172 = ($signed(_zz_10173) >>> _zz_2791);
  assign _zz_10173 = _zz_10174;
  assign _zz_10174 = ($signed(_zz_784) - $signed(_zz_2789));
  assign _zz_10175 = _zz_10176;
  assign _zz_10176 = ($signed(_zz_10177) >>> _zz_2792);
  assign _zz_10177 = _zz_10178;
  assign _zz_10178 = ($signed(_zz_783) + $signed(_zz_2788));
  assign _zz_10179 = _zz_10180;
  assign _zz_10180 = ($signed(_zz_10181) >>> _zz_2792);
  assign _zz_10181 = _zz_10182;
  assign _zz_10182 = ($signed(_zz_784) + $signed(_zz_2789));
  assign _zz_10183 = ($signed(twiddle_factor_table_7_real) + $signed(twiddle_factor_table_7_imag));
  assign _zz_10184 = fixTo_600_dout;
  assign _zz_10185 = ($signed(_zz_818) - $signed(_zz_817));
  assign _zz_10186 = ($signed(_zz_817) + $signed(_zz_818));
  assign _zz_10187 = _zz_10188[15 : 0];
  assign _zz_10188 = fixTo_602_dout;
  assign _zz_10189 = _zz_10190[15 : 0];
  assign _zz_10190 = fixTo_601_dout;
  assign _zz_10191 = _zz_10192;
  assign _zz_10192 = ($signed(_zz_10193) >>> _zz_2796);
  assign _zz_10193 = _zz_10194;
  assign _zz_10194 = ($signed(_zz_801) - $signed(_zz_2793));
  assign _zz_10195 = _zz_10196;
  assign _zz_10196 = ($signed(_zz_10197) >>> _zz_2796);
  assign _zz_10197 = _zz_10198;
  assign _zz_10198 = ($signed(_zz_802) - $signed(_zz_2794));
  assign _zz_10199 = _zz_10200;
  assign _zz_10200 = ($signed(_zz_10201) >>> _zz_2797);
  assign _zz_10201 = _zz_10202;
  assign _zz_10202 = ($signed(_zz_801) + $signed(_zz_2793));
  assign _zz_10203 = _zz_10204;
  assign _zz_10204 = ($signed(_zz_10205) >>> _zz_2797);
  assign _zz_10205 = _zz_10206;
  assign _zz_10206 = ($signed(_zz_802) + $signed(_zz_2794));
  assign _zz_10207 = ($signed(twiddle_factor_table_8_real) + $signed(twiddle_factor_table_8_imag));
  assign _zz_10208 = fixTo_603_dout;
  assign _zz_10209 = ($signed(_zz_820) - $signed(_zz_819));
  assign _zz_10210 = ($signed(_zz_819) + $signed(_zz_820));
  assign _zz_10211 = _zz_10212[15 : 0];
  assign _zz_10212 = fixTo_605_dout;
  assign _zz_10213 = _zz_10214[15 : 0];
  assign _zz_10214 = fixTo_604_dout;
  assign _zz_10215 = _zz_10216;
  assign _zz_10216 = ($signed(_zz_10217) >>> _zz_2801);
  assign _zz_10217 = _zz_10218;
  assign _zz_10218 = ($signed(_zz_803) - $signed(_zz_2798));
  assign _zz_10219 = _zz_10220;
  assign _zz_10220 = ($signed(_zz_10221) >>> _zz_2801);
  assign _zz_10221 = _zz_10222;
  assign _zz_10222 = ($signed(_zz_804) - $signed(_zz_2799));
  assign _zz_10223 = _zz_10224;
  assign _zz_10224 = ($signed(_zz_10225) >>> _zz_2802);
  assign _zz_10225 = _zz_10226;
  assign _zz_10226 = ($signed(_zz_803) + $signed(_zz_2798));
  assign _zz_10227 = _zz_10228;
  assign _zz_10228 = ($signed(_zz_10229) >>> _zz_2802);
  assign _zz_10229 = _zz_10230;
  assign _zz_10230 = ($signed(_zz_804) + $signed(_zz_2799));
  assign _zz_10231 = ($signed(twiddle_factor_table_9_real) + $signed(twiddle_factor_table_9_imag));
  assign _zz_10232 = fixTo_606_dout;
  assign _zz_10233 = ($signed(_zz_822) - $signed(_zz_821));
  assign _zz_10234 = ($signed(_zz_821) + $signed(_zz_822));
  assign _zz_10235 = _zz_10236[15 : 0];
  assign _zz_10236 = fixTo_608_dout;
  assign _zz_10237 = _zz_10238[15 : 0];
  assign _zz_10238 = fixTo_607_dout;
  assign _zz_10239 = _zz_10240;
  assign _zz_10240 = ($signed(_zz_10241) >>> _zz_2806);
  assign _zz_10241 = _zz_10242;
  assign _zz_10242 = ($signed(_zz_805) - $signed(_zz_2803));
  assign _zz_10243 = _zz_10244;
  assign _zz_10244 = ($signed(_zz_10245) >>> _zz_2806);
  assign _zz_10245 = _zz_10246;
  assign _zz_10246 = ($signed(_zz_806) - $signed(_zz_2804));
  assign _zz_10247 = _zz_10248;
  assign _zz_10248 = ($signed(_zz_10249) >>> _zz_2807);
  assign _zz_10249 = _zz_10250;
  assign _zz_10250 = ($signed(_zz_805) + $signed(_zz_2803));
  assign _zz_10251 = _zz_10252;
  assign _zz_10252 = ($signed(_zz_10253) >>> _zz_2807);
  assign _zz_10253 = _zz_10254;
  assign _zz_10254 = ($signed(_zz_806) + $signed(_zz_2804));
  assign _zz_10255 = ($signed(twiddle_factor_table_10_real) + $signed(twiddle_factor_table_10_imag));
  assign _zz_10256 = fixTo_609_dout;
  assign _zz_10257 = ($signed(_zz_824) - $signed(_zz_823));
  assign _zz_10258 = ($signed(_zz_823) + $signed(_zz_824));
  assign _zz_10259 = _zz_10260[15 : 0];
  assign _zz_10260 = fixTo_611_dout;
  assign _zz_10261 = _zz_10262[15 : 0];
  assign _zz_10262 = fixTo_610_dout;
  assign _zz_10263 = _zz_10264;
  assign _zz_10264 = ($signed(_zz_10265) >>> _zz_2811);
  assign _zz_10265 = _zz_10266;
  assign _zz_10266 = ($signed(_zz_807) - $signed(_zz_2808));
  assign _zz_10267 = _zz_10268;
  assign _zz_10268 = ($signed(_zz_10269) >>> _zz_2811);
  assign _zz_10269 = _zz_10270;
  assign _zz_10270 = ($signed(_zz_808) - $signed(_zz_2809));
  assign _zz_10271 = _zz_10272;
  assign _zz_10272 = ($signed(_zz_10273) >>> _zz_2812);
  assign _zz_10273 = _zz_10274;
  assign _zz_10274 = ($signed(_zz_807) + $signed(_zz_2808));
  assign _zz_10275 = _zz_10276;
  assign _zz_10276 = ($signed(_zz_10277) >>> _zz_2812);
  assign _zz_10277 = _zz_10278;
  assign _zz_10278 = ($signed(_zz_808) + $signed(_zz_2809));
  assign _zz_10279 = ($signed(twiddle_factor_table_11_real) + $signed(twiddle_factor_table_11_imag));
  assign _zz_10280 = fixTo_612_dout;
  assign _zz_10281 = ($signed(_zz_826) - $signed(_zz_825));
  assign _zz_10282 = ($signed(_zz_825) + $signed(_zz_826));
  assign _zz_10283 = _zz_10284[15 : 0];
  assign _zz_10284 = fixTo_614_dout;
  assign _zz_10285 = _zz_10286[15 : 0];
  assign _zz_10286 = fixTo_613_dout;
  assign _zz_10287 = _zz_10288;
  assign _zz_10288 = ($signed(_zz_10289) >>> _zz_2816);
  assign _zz_10289 = _zz_10290;
  assign _zz_10290 = ($signed(_zz_809) - $signed(_zz_2813));
  assign _zz_10291 = _zz_10292;
  assign _zz_10292 = ($signed(_zz_10293) >>> _zz_2816);
  assign _zz_10293 = _zz_10294;
  assign _zz_10294 = ($signed(_zz_810) - $signed(_zz_2814));
  assign _zz_10295 = _zz_10296;
  assign _zz_10296 = ($signed(_zz_10297) >>> _zz_2817);
  assign _zz_10297 = _zz_10298;
  assign _zz_10298 = ($signed(_zz_809) + $signed(_zz_2813));
  assign _zz_10299 = _zz_10300;
  assign _zz_10300 = ($signed(_zz_10301) >>> _zz_2817);
  assign _zz_10301 = _zz_10302;
  assign _zz_10302 = ($signed(_zz_810) + $signed(_zz_2814));
  assign _zz_10303 = ($signed(twiddle_factor_table_12_real) + $signed(twiddle_factor_table_12_imag));
  assign _zz_10304 = fixTo_615_dout;
  assign _zz_10305 = ($signed(_zz_828) - $signed(_zz_827));
  assign _zz_10306 = ($signed(_zz_827) + $signed(_zz_828));
  assign _zz_10307 = _zz_10308[15 : 0];
  assign _zz_10308 = fixTo_617_dout;
  assign _zz_10309 = _zz_10310[15 : 0];
  assign _zz_10310 = fixTo_616_dout;
  assign _zz_10311 = _zz_10312;
  assign _zz_10312 = ($signed(_zz_10313) >>> _zz_2821);
  assign _zz_10313 = _zz_10314;
  assign _zz_10314 = ($signed(_zz_811) - $signed(_zz_2818));
  assign _zz_10315 = _zz_10316;
  assign _zz_10316 = ($signed(_zz_10317) >>> _zz_2821);
  assign _zz_10317 = _zz_10318;
  assign _zz_10318 = ($signed(_zz_812) - $signed(_zz_2819));
  assign _zz_10319 = _zz_10320;
  assign _zz_10320 = ($signed(_zz_10321) >>> _zz_2822);
  assign _zz_10321 = _zz_10322;
  assign _zz_10322 = ($signed(_zz_811) + $signed(_zz_2818));
  assign _zz_10323 = _zz_10324;
  assign _zz_10324 = ($signed(_zz_10325) >>> _zz_2822);
  assign _zz_10325 = _zz_10326;
  assign _zz_10326 = ($signed(_zz_812) + $signed(_zz_2819));
  assign _zz_10327 = ($signed(twiddle_factor_table_13_real) + $signed(twiddle_factor_table_13_imag));
  assign _zz_10328 = fixTo_618_dout;
  assign _zz_10329 = ($signed(_zz_830) - $signed(_zz_829));
  assign _zz_10330 = ($signed(_zz_829) + $signed(_zz_830));
  assign _zz_10331 = _zz_10332[15 : 0];
  assign _zz_10332 = fixTo_620_dout;
  assign _zz_10333 = _zz_10334[15 : 0];
  assign _zz_10334 = fixTo_619_dout;
  assign _zz_10335 = _zz_10336;
  assign _zz_10336 = ($signed(_zz_10337) >>> _zz_2826);
  assign _zz_10337 = _zz_10338;
  assign _zz_10338 = ($signed(_zz_813) - $signed(_zz_2823));
  assign _zz_10339 = _zz_10340;
  assign _zz_10340 = ($signed(_zz_10341) >>> _zz_2826);
  assign _zz_10341 = _zz_10342;
  assign _zz_10342 = ($signed(_zz_814) - $signed(_zz_2824));
  assign _zz_10343 = _zz_10344;
  assign _zz_10344 = ($signed(_zz_10345) >>> _zz_2827);
  assign _zz_10345 = _zz_10346;
  assign _zz_10346 = ($signed(_zz_813) + $signed(_zz_2823));
  assign _zz_10347 = _zz_10348;
  assign _zz_10348 = ($signed(_zz_10349) >>> _zz_2827);
  assign _zz_10349 = _zz_10350;
  assign _zz_10350 = ($signed(_zz_814) + $signed(_zz_2824));
  assign _zz_10351 = ($signed(twiddle_factor_table_14_real) + $signed(twiddle_factor_table_14_imag));
  assign _zz_10352 = fixTo_621_dout;
  assign _zz_10353 = ($signed(_zz_832) - $signed(_zz_831));
  assign _zz_10354 = ($signed(_zz_831) + $signed(_zz_832));
  assign _zz_10355 = _zz_10356[15 : 0];
  assign _zz_10356 = fixTo_623_dout;
  assign _zz_10357 = _zz_10358[15 : 0];
  assign _zz_10358 = fixTo_622_dout;
  assign _zz_10359 = _zz_10360;
  assign _zz_10360 = ($signed(_zz_10361) >>> _zz_2831);
  assign _zz_10361 = _zz_10362;
  assign _zz_10362 = ($signed(_zz_815) - $signed(_zz_2828));
  assign _zz_10363 = _zz_10364;
  assign _zz_10364 = ($signed(_zz_10365) >>> _zz_2831);
  assign _zz_10365 = _zz_10366;
  assign _zz_10366 = ($signed(_zz_816) - $signed(_zz_2829));
  assign _zz_10367 = _zz_10368;
  assign _zz_10368 = ($signed(_zz_10369) >>> _zz_2832);
  assign _zz_10369 = _zz_10370;
  assign _zz_10370 = ($signed(_zz_815) + $signed(_zz_2828));
  assign _zz_10371 = _zz_10372;
  assign _zz_10372 = ($signed(_zz_10373) >>> _zz_2832);
  assign _zz_10373 = _zz_10374;
  assign _zz_10374 = ($signed(_zz_816) + $signed(_zz_2829));
  assign _zz_10375 = ($signed(twiddle_factor_table_7_real) + $signed(twiddle_factor_table_7_imag));
  assign _zz_10376 = fixTo_624_dout;
  assign _zz_10377 = ($signed(_zz_850) - $signed(_zz_849));
  assign _zz_10378 = ($signed(_zz_849) + $signed(_zz_850));
  assign _zz_10379 = _zz_10380[15 : 0];
  assign _zz_10380 = fixTo_626_dout;
  assign _zz_10381 = _zz_10382[15 : 0];
  assign _zz_10382 = fixTo_625_dout;
  assign _zz_10383 = _zz_10384;
  assign _zz_10384 = ($signed(_zz_10385) >>> _zz_2836);
  assign _zz_10385 = _zz_10386;
  assign _zz_10386 = ($signed(_zz_833) - $signed(_zz_2833));
  assign _zz_10387 = _zz_10388;
  assign _zz_10388 = ($signed(_zz_10389) >>> _zz_2836);
  assign _zz_10389 = _zz_10390;
  assign _zz_10390 = ($signed(_zz_834) - $signed(_zz_2834));
  assign _zz_10391 = _zz_10392;
  assign _zz_10392 = ($signed(_zz_10393) >>> _zz_2837);
  assign _zz_10393 = _zz_10394;
  assign _zz_10394 = ($signed(_zz_833) + $signed(_zz_2833));
  assign _zz_10395 = _zz_10396;
  assign _zz_10396 = ($signed(_zz_10397) >>> _zz_2837);
  assign _zz_10397 = _zz_10398;
  assign _zz_10398 = ($signed(_zz_834) + $signed(_zz_2834));
  assign _zz_10399 = ($signed(twiddle_factor_table_8_real) + $signed(twiddle_factor_table_8_imag));
  assign _zz_10400 = fixTo_627_dout;
  assign _zz_10401 = ($signed(_zz_852) - $signed(_zz_851));
  assign _zz_10402 = ($signed(_zz_851) + $signed(_zz_852));
  assign _zz_10403 = _zz_10404[15 : 0];
  assign _zz_10404 = fixTo_629_dout;
  assign _zz_10405 = _zz_10406[15 : 0];
  assign _zz_10406 = fixTo_628_dout;
  assign _zz_10407 = _zz_10408;
  assign _zz_10408 = ($signed(_zz_10409) >>> _zz_2841);
  assign _zz_10409 = _zz_10410;
  assign _zz_10410 = ($signed(_zz_835) - $signed(_zz_2838));
  assign _zz_10411 = _zz_10412;
  assign _zz_10412 = ($signed(_zz_10413) >>> _zz_2841);
  assign _zz_10413 = _zz_10414;
  assign _zz_10414 = ($signed(_zz_836) - $signed(_zz_2839));
  assign _zz_10415 = _zz_10416;
  assign _zz_10416 = ($signed(_zz_10417) >>> _zz_2842);
  assign _zz_10417 = _zz_10418;
  assign _zz_10418 = ($signed(_zz_835) + $signed(_zz_2838));
  assign _zz_10419 = _zz_10420;
  assign _zz_10420 = ($signed(_zz_10421) >>> _zz_2842);
  assign _zz_10421 = _zz_10422;
  assign _zz_10422 = ($signed(_zz_836) + $signed(_zz_2839));
  assign _zz_10423 = ($signed(twiddle_factor_table_9_real) + $signed(twiddle_factor_table_9_imag));
  assign _zz_10424 = fixTo_630_dout;
  assign _zz_10425 = ($signed(_zz_854) - $signed(_zz_853));
  assign _zz_10426 = ($signed(_zz_853) + $signed(_zz_854));
  assign _zz_10427 = _zz_10428[15 : 0];
  assign _zz_10428 = fixTo_632_dout;
  assign _zz_10429 = _zz_10430[15 : 0];
  assign _zz_10430 = fixTo_631_dout;
  assign _zz_10431 = _zz_10432;
  assign _zz_10432 = ($signed(_zz_10433) >>> _zz_2846);
  assign _zz_10433 = _zz_10434;
  assign _zz_10434 = ($signed(_zz_837) - $signed(_zz_2843));
  assign _zz_10435 = _zz_10436;
  assign _zz_10436 = ($signed(_zz_10437) >>> _zz_2846);
  assign _zz_10437 = _zz_10438;
  assign _zz_10438 = ($signed(_zz_838) - $signed(_zz_2844));
  assign _zz_10439 = _zz_10440;
  assign _zz_10440 = ($signed(_zz_10441) >>> _zz_2847);
  assign _zz_10441 = _zz_10442;
  assign _zz_10442 = ($signed(_zz_837) + $signed(_zz_2843));
  assign _zz_10443 = _zz_10444;
  assign _zz_10444 = ($signed(_zz_10445) >>> _zz_2847);
  assign _zz_10445 = _zz_10446;
  assign _zz_10446 = ($signed(_zz_838) + $signed(_zz_2844));
  assign _zz_10447 = ($signed(twiddle_factor_table_10_real) + $signed(twiddle_factor_table_10_imag));
  assign _zz_10448 = fixTo_633_dout;
  assign _zz_10449 = ($signed(_zz_856) - $signed(_zz_855));
  assign _zz_10450 = ($signed(_zz_855) + $signed(_zz_856));
  assign _zz_10451 = _zz_10452[15 : 0];
  assign _zz_10452 = fixTo_635_dout;
  assign _zz_10453 = _zz_10454[15 : 0];
  assign _zz_10454 = fixTo_634_dout;
  assign _zz_10455 = _zz_10456;
  assign _zz_10456 = ($signed(_zz_10457) >>> _zz_2851);
  assign _zz_10457 = _zz_10458;
  assign _zz_10458 = ($signed(_zz_839) - $signed(_zz_2848));
  assign _zz_10459 = _zz_10460;
  assign _zz_10460 = ($signed(_zz_10461) >>> _zz_2851);
  assign _zz_10461 = _zz_10462;
  assign _zz_10462 = ($signed(_zz_840) - $signed(_zz_2849));
  assign _zz_10463 = _zz_10464;
  assign _zz_10464 = ($signed(_zz_10465) >>> _zz_2852);
  assign _zz_10465 = _zz_10466;
  assign _zz_10466 = ($signed(_zz_839) + $signed(_zz_2848));
  assign _zz_10467 = _zz_10468;
  assign _zz_10468 = ($signed(_zz_10469) >>> _zz_2852);
  assign _zz_10469 = _zz_10470;
  assign _zz_10470 = ($signed(_zz_840) + $signed(_zz_2849));
  assign _zz_10471 = ($signed(twiddle_factor_table_11_real) + $signed(twiddle_factor_table_11_imag));
  assign _zz_10472 = fixTo_636_dout;
  assign _zz_10473 = ($signed(_zz_858) - $signed(_zz_857));
  assign _zz_10474 = ($signed(_zz_857) + $signed(_zz_858));
  assign _zz_10475 = _zz_10476[15 : 0];
  assign _zz_10476 = fixTo_638_dout;
  assign _zz_10477 = _zz_10478[15 : 0];
  assign _zz_10478 = fixTo_637_dout;
  assign _zz_10479 = _zz_10480;
  assign _zz_10480 = ($signed(_zz_10481) >>> _zz_2856);
  assign _zz_10481 = _zz_10482;
  assign _zz_10482 = ($signed(_zz_841) - $signed(_zz_2853));
  assign _zz_10483 = _zz_10484;
  assign _zz_10484 = ($signed(_zz_10485) >>> _zz_2856);
  assign _zz_10485 = _zz_10486;
  assign _zz_10486 = ($signed(_zz_842) - $signed(_zz_2854));
  assign _zz_10487 = _zz_10488;
  assign _zz_10488 = ($signed(_zz_10489) >>> _zz_2857);
  assign _zz_10489 = _zz_10490;
  assign _zz_10490 = ($signed(_zz_841) + $signed(_zz_2853));
  assign _zz_10491 = _zz_10492;
  assign _zz_10492 = ($signed(_zz_10493) >>> _zz_2857);
  assign _zz_10493 = _zz_10494;
  assign _zz_10494 = ($signed(_zz_842) + $signed(_zz_2854));
  assign _zz_10495 = ($signed(twiddle_factor_table_12_real) + $signed(twiddle_factor_table_12_imag));
  assign _zz_10496 = fixTo_639_dout;
  assign _zz_10497 = ($signed(_zz_860) - $signed(_zz_859));
  assign _zz_10498 = ($signed(_zz_859) + $signed(_zz_860));
  assign _zz_10499 = _zz_10500[15 : 0];
  assign _zz_10500 = fixTo_641_dout;
  assign _zz_10501 = _zz_10502[15 : 0];
  assign _zz_10502 = fixTo_640_dout;
  assign _zz_10503 = _zz_10504;
  assign _zz_10504 = ($signed(_zz_10505) >>> _zz_2861);
  assign _zz_10505 = _zz_10506;
  assign _zz_10506 = ($signed(_zz_843) - $signed(_zz_2858));
  assign _zz_10507 = _zz_10508;
  assign _zz_10508 = ($signed(_zz_10509) >>> _zz_2861);
  assign _zz_10509 = _zz_10510;
  assign _zz_10510 = ($signed(_zz_844) - $signed(_zz_2859));
  assign _zz_10511 = _zz_10512;
  assign _zz_10512 = ($signed(_zz_10513) >>> _zz_2862);
  assign _zz_10513 = _zz_10514;
  assign _zz_10514 = ($signed(_zz_843) + $signed(_zz_2858));
  assign _zz_10515 = _zz_10516;
  assign _zz_10516 = ($signed(_zz_10517) >>> _zz_2862);
  assign _zz_10517 = _zz_10518;
  assign _zz_10518 = ($signed(_zz_844) + $signed(_zz_2859));
  assign _zz_10519 = ($signed(twiddle_factor_table_13_real) + $signed(twiddle_factor_table_13_imag));
  assign _zz_10520 = fixTo_642_dout;
  assign _zz_10521 = ($signed(_zz_862) - $signed(_zz_861));
  assign _zz_10522 = ($signed(_zz_861) + $signed(_zz_862));
  assign _zz_10523 = _zz_10524[15 : 0];
  assign _zz_10524 = fixTo_644_dout;
  assign _zz_10525 = _zz_10526[15 : 0];
  assign _zz_10526 = fixTo_643_dout;
  assign _zz_10527 = _zz_10528;
  assign _zz_10528 = ($signed(_zz_10529) >>> _zz_2866);
  assign _zz_10529 = _zz_10530;
  assign _zz_10530 = ($signed(_zz_845) - $signed(_zz_2863));
  assign _zz_10531 = _zz_10532;
  assign _zz_10532 = ($signed(_zz_10533) >>> _zz_2866);
  assign _zz_10533 = _zz_10534;
  assign _zz_10534 = ($signed(_zz_846) - $signed(_zz_2864));
  assign _zz_10535 = _zz_10536;
  assign _zz_10536 = ($signed(_zz_10537) >>> _zz_2867);
  assign _zz_10537 = _zz_10538;
  assign _zz_10538 = ($signed(_zz_845) + $signed(_zz_2863));
  assign _zz_10539 = _zz_10540;
  assign _zz_10540 = ($signed(_zz_10541) >>> _zz_2867);
  assign _zz_10541 = _zz_10542;
  assign _zz_10542 = ($signed(_zz_846) + $signed(_zz_2864));
  assign _zz_10543 = ($signed(twiddle_factor_table_14_real) + $signed(twiddle_factor_table_14_imag));
  assign _zz_10544 = fixTo_645_dout;
  assign _zz_10545 = ($signed(_zz_864) - $signed(_zz_863));
  assign _zz_10546 = ($signed(_zz_863) + $signed(_zz_864));
  assign _zz_10547 = _zz_10548[15 : 0];
  assign _zz_10548 = fixTo_647_dout;
  assign _zz_10549 = _zz_10550[15 : 0];
  assign _zz_10550 = fixTo_646_dout;
  assign _zz_10551 = _zz_10552;
  assign _zz_10552 = ($signed(_zz_10553) >>> _zz_2871);
  assign _zz_10553 = _zz_10554;
  assign _zz_10554 = ($signed(_zz_847) - $signed(_zz_2868));
  assign _zz_10555 = _zz_10556;
  assign _zz_10556 = ($signed(_zz_10557) >>> _zz_2871);
  assign _zz_10557 = _zz_10558;
  assign _zz_10558 = ($signed(_zz_848) - $signed(_zz_2869));
  assign _zz_10559 = _zz_10560;
  assign _zz_10560 = ($signed(_zz_10561) >>> _zz_2872);
  assign _zz_10561 = _zz_10562;
  assign _zz_10562 = ($signed(_zz_847) + $signed(_zz_2868));
  assign _zz_10563 = _zz_10564;
  assign _zz_10564 = ($signed(_zz_10565) >>> _zz_2872);
  assign _zz_10565 = _zz_10566;
  assign _zz_10566 = ($signed(_zz_848) + $signed(_zz_2869));
  assign _zz_10567 = ($signed(twiddle_factor_table_7_real) + $signed(twiddle_factor_table_7_imag));
  assign _zz_10568 = fixTo_648_dout;
  assign _zz_10569 = ($signed(_zz_882) - $signed(_zz_881));
  assign _zz_10570 = ($signed(_zz_881) + $signed(_zz_882));
  assign _zz_10571 = _zz_10572[15 : 0];
  assign _zz_10572 = fixTo_650_dout;
  assign _zz_10573 = _zz_10574[15 : 0];
  assign _zz_10574 = fixTo_649_dout;
  assign _zz_10575 = _zz_10576;
  assign _zz_10576 = ($signed(_zz_10577) >>> _zz_2876);
  assign _zz_10577 = _zz_10578;
  assign _zz_10578 = ($signed(_zz_865) - $signed(_zz_2873));
  assign _zz_10579 = _zz_10580;
  assign _zz_10580 = ($signed(_zz_10581) >>> _zz_2876);
  assign _zz_10581 = _zz_10582;
  assign _zz_10582 = ($signed(_zz_866) - $signed(_zz_2874));
  assign _zz_10583 = _zz_10584;
  assign _zz_10584 = ($signed(_zz_10585) >>> _zz_2877);
  assign _zz_10585 = _zz_10586;
  assign _zz_10586 = ($signed(_zz_865) + $signed(_zz_2873));
  assign _zz_10587 = _zz_10588;
  assign _zz_10588 = ($signed(_zz_10589) >>> _zz_2877);
  assign _zz_10589 = _zz_10590;
  assign _zz_10590 = ($signed(_zz_866) + $signed(_zz_2874));
  assign _zz_10591 = ($signed(twiddle_factor_table_8_real) + $signed(twiddle_factor_table_8_imag));
  assign _zz_10592 = fixTo_651_dout;
  assign _zz_10593 = ($signed(_zz_884) - $signed(_zz_883));
  assign _zz_10594 = ($signed(_zz_883) + $signed(_zz_884));
  assign _zz_10595 = _zz_10596[15 : 0];
  assign _zz_10596 = fixTo_653_dout;
  assign _zz_10597 = _zz_10598[15 : 0];
  assign _zz_10598 = fixTo_652_dout;
  assign _zz_10599 = _zz_10600;
  assign _zz_10600 = ($signed(_zz_10601) >>> _zz_2881);
  assign _zz_10601 = _zz_10602;
  assign _zz_10602 = ($signed(_zz_867) - $signed(_zz_2878));
  assign _zz_10603 = _zz_10604;
  assign _zz_10604 = ($signed(_zz_10605) >>> _zz_2881);
  assign _zz_10605 = _zz_10606;
  assign _zz_10606 = ($signed(_zz_868) - $signed(_zz_2879));
  assign _zz_10607 = _zz_10608;
  assign _zz_10608 = ($signed(_zz_10609) >>> _zz_2882);
  assign _zz_10609 = _zz_10610;
  assign _zz_10610 = ($signed(_zz_867) + $signed(_zz_2878));
  assign _zz_10611 = _zz_10612;
  assign _zz_10612 = ($signed(_zz_10613) >>> _zz_2882);
  assign _zz_10613 = _zz_10614;
  assign _zz_10614 = ($signed(_zz_868) + $signed(_zz_2879));
  assign _zz_10615 = ($signed(twiddle_factor_table_9_real) + $signed(twiddle_factor_table_9_imag));
  assign _zz_10616 = fixTo_654_dout;
  assign _zz_10617 = ($signed(_zz_886) - $signed(_zz_885));
  assign _zz_10618 = ($signed(_zz_885) + $signed(_zz_886));
  assign _zz_10619 = _zz_10620[15 : 0];
  assign _zz_10620 = fixTo_656_dout;
  assign _zz_10621 = _zz_10622[15 : 0];
  assign _zz_10622 = fixTo_655_dout;
  assign _zz_10623 = _zz_10624;
  assign _zz_10624 = ($signed(_zz_10625) >>> _zz_2886);
  assign _zz_10625 = _zz_10626;
  assign _zz_10626 = ($signed(_zz_869) - $signed(_zz_2883));
  assign _zz_10627 = _zz_10628;
  assign _zz_10628 = ($signed(_zz_10629) >>> _zz_2886);
  assign _zz_10629 = _zz_10630;
  assign _zz_10630 = ($signed(_zz_870) - $signed(_zz_2884));
  assign _zz_10631 = _zz_10632;
  assign _zz_10632 = ($signed(_zz_10633) >>> _zz_2887);
  assign _zz_10633 = _zz_10634;
  assign _zz_10634 = ($signed(_zz_869) + $signed(_zz_2883));
  assign _zz_10635 = _zz_10636;
  assign _zz_10636 = ($signed(_zz_10637) >>> _zz_2887);
  assign _zz_10637 = _zz_10638;
  assign _zz_10638 = ($signed(_zz_870) + $signed(_zz_2884));
  assign _zz_10639 = ($signed(twiddle_factor_table_10_real) + $signed(twiddle_factor_table_10_imag));
  assign _zz_10640 = fixTo_657_dout;
  assign _zz_10641 = ($signed(_zz_888) - $signed(_zz_887));
  assign _zz_10642 = ($signed(_zz_887) + $signed(_zz_888));
  assign _zz_10643 = _zz_10644[15 : 0];
  assign _zz_10644 = fixTo_659_dout;
  assign _zz_10645 = _zz_10646[15 : 0];
  assign _zz_10646 = fixTo_658_dout;
  assign _zz_10647 = _zz_10648;
  assign _zz_10648 = ($signed(_zz_10649) >>> _zz_2891);
  assign _zz_10649 = _zz_10650;
  assign _zz_10650 = ($signed(_zz_871) - $signed(_zz_2888));
  assign _zz_10651 = _zz_10652;
  assign _zz_10652 = ($signed(_zz_10653) >>> _zz_2891);
  assign _zz_10653 = _zz_10654;
  assign _zz_10654 = ($signed(_zz_872) - $signed(_zz_2889));
  assign _zz_10655 = _zz_10656;
  assign _zz_10656 = ($signed(_zz_10657) >>> _zz_2892);
  assign _zz_10657 = _zz_10658;
  assign _zz_10658 = ($signed(_zz_871) + $signed(_zz_2888));
  assign _zz_10659 = _zz_10660;
  assign _zz_10660 = ($signed(_zz_10661) >>> _zz_2892);
  assign _zz_10661 = _zz_10662;
  assign _zz_10662 = ($signed(_zz_872) + $signed(_zz_2889));
  assign _zz_10663 = ($signed(twiddle_factor_table_11_real) + $signed(twiddle_factor_table_11_imag));
  assign _zz_10664 = fixTo_660_dout;
  assign _zz_10665 = ($signed(_zz_890) - $signed(_zz_889));
  assign _zz_10666 = ($signed(_zz_889) + $signed(_zz_890));
  assign _zz_10667 = _zz_10668[15 : 0];
  assign _zz_10668 = fixTo_662_dout;
  assign _zz_10669 = _zz_10670[15 : 0];
  assign _zz_10670 = fixTo_661_dout;
  assign _zz_10671 = _zz_10672;
  assign _zz_10672 = ($signed(_zz_10673) >>> _zz_2896);
  assign _zz_10673 = _zz_10674;
  assign _zz_10674 = ($signed(_zz_873) - $signed(_zz_2893));
  assign _zz_10675 = _zz_10676;
  assign _zz_10676 = ($signed(_zz_10677) >>> _zz_2896);
  assign _zz_10677 = _zz_10678;
  assign _zz_10678 = ($signed(_zz_874) - $signed(_zz_2894));
  assign _zz_10679 = _zz_10680;
  assign _zz_10680 = ($signed(_zz_10681) >>> _zz_2897);
  assign _zz_10681 = _zz_10682;
  assign _zz_10682 = ($signed(_zz_873) + $signed(_zz_2893));
  assign _zz_10683 = _zz_10684;
  assign _zz_10684 = ($signed(_zz_10685) >>> _zz_2897);
  assign _zz_10685 = _zz_10686;
  assign _zz_10686 = ($signed(_zz_874) + $signed(_zz_2894));
  assign _zz_10687 = ($signed(twiddle_factor_table_12_real) + $signed(twiddle_factor_table_12_imag));
  assign _zz_10688 = fixTo_663_dout;
  assign _zz_10689 = ($signed(_zz_892) - $signed(_zz_891));
  assign _zz_10690 = ($signed(_zz_891) + $signed(_zz_892));
  assign _zz_10691 = _zz_10692[15 : 0];
  assign _zz_10692 = fixTo_665_dout;
  assign _zz_10693 = _zz_10694[15 : 0];
  assign _zz_10694 = fixTo_664_dout;
  assign _zz_10695 = _zz_10696;
  assign _zz_10696 = ($signed(_zz_10697) >>> _zz_2901);
  assign _zz_10697 = _zz_10698;
  assign _zz_10698 = ($signed(_zz_875) - $signed(_zz_2898));
  assign _zz_10699 = _zz_10700;
  assign _zz_10700 = ($signed(_zz_10701) >>> _zz_2901);
  assign _zz_10701 = _zz_10702;
  assign _zz_10702 = ($signed(_zz_876) - $signed(_zz_2899));
  assign _zz_10703 = _zz_10704;
  assign _zz_10704 = ($signed(_zz_10705) >>> _zz_2902);
  assign _zz_10705 = _zz_10706;
  assign _zz_10706 = ($signed(_zz_875) + $signed(_zz_2898));
  assign _zz_10707 = _zz_10708;
  assign _zz_10708 = ($signed(_zz_10709) >>> _zz_2902);
  assign _zz_10709 = _zz_10710;
  assign _zz_10710 = ($signed(_zz_876) + $signed(_zz_2899));
  assign _zz_10711 = ($signed(twiddle_factor_table_13_real) + $signed(twiddle_factor_table_13_imag));
  assign _zz_10712 = fixTo_666_dout;
  assign _zz_10713 = ($signed(_zz_894) - $signed(_zz_893));
  assign _zz_10714 = ($signed(_zz_893) + $signed(_zz_894));
  assign _zz_10715 = _zz_10716[15 : 0];
  assign _zz_10716 = fixTo_668_dout;
  assign _zz_10717 = _zz_10718[15 : 0];
  assign _zz_10718 = fixTo_667_dout;
  assign _zz_10719 = _zz_10720;
  assign _zz_10720 = ($signed(_zz_10721) >>> _zz_2906);
  assign _zz_10721 = _zz_10722;
  assign _zz_10722 = ($signed(_zz_877) - $signed(_zz_2903));
  assign _zz_10723 = _zz_10724;
  assign _zz_10724 = ($signed(_zz_10725) >>> _zz_2906);
  assign _zz_10725 = _zz_10726;
  assign _zz_10726 = ($signed(_zz_878) - $signed(_zz_2904));
  assign _zz_10727 = _zz_10728;
  assign _zz_10728 = ($signed(_zz_10729) >>> _zz_2907);
  assign _zz_10729 = _zz_10730;
  assign _zz_10730 = ($signed(_zz_877) + $signed(_zz_2903));
  assign _zz_10731 = _zz_10732;
  assign _zz_10732 = ($signed(_zz_10733) >>> _zz_2907);
  assign _zz_10733 = _zz_10734;
  assign _zz_10734 = ($signed(_zz_878) + $signed(_zz_2904));
  assign _zz_10735 = ($signed(twiddle_factor_table_14_real) + $signed(twiddle_factor_table_14_imag));
  assign _zz_10736 = fixTo_669_dout;
  assign _zz_10737 = ($signed(_zz_896) - $signed(_zz_895));
  assign _zz_10738 = ($signed(_zz_895) + $signed(_zz_896));
  assign _zz_10739 = _zz_10740[15 : 0];
  assign _zz_10740 = fixTo_671_dout;
  assign _zz_10741 = _zz_10742[15 : 0];
  assign _zz_10742 = fixTo_670_dout;
  assign _zz_10743 = _zz_10744;
  assign _zz_10744 = ($signed(_zz_10745) >>> _zz_2911);
  assign _zz_10745 = _zz_10746;
  assign _zz_10746 = ($signed(_zz_879) - $signed(_zz_2908));
  assign _zz_10747 = _zz_10748;
  assign _zz_10748 = ($signed(_zz_10749) >>> _zz_2911);
  assign _zz_10749 = _zz_10750;
  assign _zz_10750 = ($signed(_zz_880) - $signed(_zz_2909));
  assign _zz_10751 = _zz_10752;
  assign _zz_10752 = ($signed(_zz_10753) >>> _zz_2912);
  assign _zz_10753 = _zz_10754;
  assign _zz_10754 = ($signed(_zz_879) + $signed(_zz_2908));
  assign _zz_10755 = _zz_10756;
  assign _zz_10756 = ($signed(_zz_10757) >>> _zz_2912);
  assign _zz_10757 = _zz_10758;
  assign _zz_10758 = ($signed(_zz_880) + $signed(_zz_2909));
  assign _zz_10759 = ($signed(twiddle_factor_table_7_real) + $signed(twiddle_factor_table_7_imag));
  assign _zz_10760 = fixTo_672_dout;
  assign _zz_10761 = ($signed(_zz_914) - $signed(_zz_913));
  assign _zz_10762 = ($signed(_zz_913) + $signed(_zz_914));
  assign _zz_10763 = _zz_10764[15 : 0];
  assign _zz_10764 = fixTo_674_dout;
  assign _zz_10765 = _zz_10766[15 : 0];
  assign _zz_10766 = fixTo_673_dout;
  assign _zz_10767 = _zz_10768;
  assign _zz_10768 = ($signed(_zz_10769) >>> _zz_2916);
  assign _zz_10769 = _zz_10770;
  assign _zz_10770 = ($signed(_zz_897) - $signed(_zz_2913));
  assign _zz_10771 = _zz_10772;
  assign _zz_10772 = ($signed(_zz_10773) >>> _zz_2916);
  assign _zz_10773 = _zz_10774;
  assign _zz_10774 = ($signed(_zz_898) - $signed(_zz_2914));
  assign _zz_10775 = _zz_10776;
  assign _zz_10776 = ($signed(_zz_10777) >>> _zz_2917);
  assign _zz_10777 = _zz_10778;
  assign _zz_10778 = ($signed(_zz_897) + $signed(_zz_2913));
  assign _zz_10779 = _zz_10780;
  assign _zz_10780 = ($signed(_zz_10781) >>> _zz_2917);
  assign _zz_10781 = _zz_10782;
  assign _zz_10782 = ($signed(_zz_898) + $signed(_zz_2914));
  assign _zz_10783 = ($signed(twiddle_factor_table_8_real) + $signed(twiddle_factor_table_8_imag));
  assign _zz_10784 = fixTo_675_dout;
  assign _zz_10785 = ($signed(_zz_916) - $signed(_zz_915));
  assign _zz_10786 = ($signed(_zz_915) + $signed(_zz_916));
  assign _zz_10787 = _zz_10788[15 : 0];
  assign _zz_10788 = fixTo_677_dout;
  assign _zz_10789 = _zz_10790[15 : 0];
  assign _zz_10790 = fixTo_676_dout;
  assign _zz_10791 = _zz_10792;
  assign _zz_10792 = ($signed(_zz_10793) >>> _zz_2921);
  assign _zz_10793 = _zz_10794;
  assign _zz_10794 = ($signed(_zz_899) - $signed(_zz_2918));
  assign _zz_10795 = _zz_10796;
  assign _zz_10796 = ($signed(_zz_10797) >>> _zz_2921);
  assign _zz_10797 = _zz_10798;
  assign _zz_10798 = ($signed(_zz_900) - $signed(_zz_2919));
  assign _zz_10799 = _zz_10800;
  assign _zz_10800 = ($signed(_zz_10801) >>> _zz_2922);
  assign _zz_10801 = _zz_10802;
  assign _zz_10802 = ($signed(_zz_899) + $signed(_zz_2918));
  assign _zz_10803 = _zz_10804;
  assign _zz_10804 = ($signed(_zz_10805) >>> _zz_2922);
  assign _zz_10805 = _zz_10806;
  assign _zz_10806 = ($signed(_zz_900) + $signed(_zz_2919));
  assign _zz_10807 = ($signed(twiddle_factor_table_9_real) + $signed(twiddle_factor_table_9_imag));
  assign _zz_10808 = fixTo_678_dout;
  assign _zz_10809 = ($signed(_zz_918) - $signed(_zz_917));
  assign _zz_10810 = ($signed(_zz_917) + $signed(_zz_918));
  assign _zz_10811 = _zz_10812[15 : 0];
  assign _zz_10812 = fixTo_680_dout;
  assign _zz_10813 = _zz_10814[15 : 0];
  assign _zz_10814 = fixTo_679_dout;
  assign _zz_10815 = _zz_10816;
  assign _zz_10816 = ($signed(_zz_10817) >>> _zz_2926);
  assign _zz_10817 = _zz_10818;
  assign _zz_10818 = ($signed(_zz_901) - $signed(_zz_2923));
  assign _zz_10819 = _zz_10820;
  assign _zz_10820 = ($signed(_zz_10821) >>> _zz_2926);
  assign _zz_10821 = _zz_10822;
  assign _zz_10822 = ($signed(_zz_902) - $signed(_zz_2924));
  assign _zz_10823 = _zz_10824;
  assign _zz_10824 = ($signed(_zz_10825) >>> _zz_2927);
  assign _zz_10825 = _zz_10826;
  assign _zz_10826 = ($signed(_zz_901) + $signed(_zz_2923));
  assign _zz_10827 = _zz_10828;
  assign _zz_10828 = ($signed(_zz_10829) >>> _zz_2927);
  assign _zz_10829 = _zz_10830;
  assign _zz_10830 = ($signed(_zz_902) + $signed(_zz_2924));
  assign _zz_10831 = ($signed(twiddle_factor_table_10_real) + $signed(twiddle_factor_table_10_imag));
  assign _zz_10832 = fixTo_681_dout;
  assign _zz_10833 = ($signed(_zz_920) - $signed(_zz_919));
  assign _zz_10834 = ($signed(_zz_919) + $signed(_zz_920));
  assign _zz_10835 = _zz_10836[15 : 0];
  assign _zz_10836 = fixTo_683_dout;
  assign _zz_10837 = _zz_10838[15 : 0];
  assign _zz_10838 = fixTo_682_dout;
  assign _zz_10839 = _zz_10840;
  assign _zz_10840 = ($signed(_zz_10841) >>> _zz_2931);
  assign _zz_10841 = _zz_10842;
  assign _zz_10842 = ($signed(_zz_903) - $signed(_zz_2928));
  assign _zz_10843 = _zz_10844;
  assign _zz_10844 = ($signed(_zz_10845) >>> _zz_2931);
  assign _zz_10845 = _zz_10846;
  assign _zz_10846 = ($signed(_zz_904) - $signed(_zz_2929));
  assign _zz_10847 = _zz_10848;
  assign _zz_10848 = ($signed(_zz_10849) >>> _zz_2932);
  assign _zz_10849 = _zz_10850;
  assign _zz_10850 = ($signed(_zz_903) + $signed(_zz_2928));
  assign _zz_10851 = _zz_10852;
  assign _zz_10852 = ($signed(_zz_10853) >>> _zz_2932);
  assign _zz_10853 = _zz_10854;
  assign _zz_10854 = ($signed(_zz_904) + $signed(_zz_2929));
  assign _zz_10855 = ($signed(twiddle_factor_table_11_real) + $signed(twiddle_factor_table_11_imag));
  assign _zz_10856 = fixTo_684_dout;
  assign _zz_10857 = ($signed(_zz_922) - $signed(_zz_921));
  assign _zz_10858 = ($signed(_zz_921) + $signed(_zz_922));
  assign _zz_10859 = _zz_10860[15 : 0];
  assign _zz_10860 = fixTo_686_dout;
  assign _zz_10861 = _zz_10862[15 : 0];
  assign _zz_10862 = fixTo_685_dout;
  assign _zz_10863 = _zz_10864;
  assign _zz_10864 = ($signed(_zz_10865) >>> _zz_2936);
  assign _zz_10865 = _zz_10866;
  assign _zz_10866 = ($signed(_zz_905) - $signed(_zz_2933));
  assign _zz_10867 = _zz_10868;
  assign _zz_10868 = ($signed(_zz_10869) >>> _zz_2936);
  assign _zz_10869 = _zz_10870;
  assign _zz_10870 = ($signed(_zz_906) - $signed(_zz_2934));
  assign _zz_10871 = _zz_10872;
  assign _zz_10872 = ($signed(_zz_10873) >>> _zz_2937);
  assign _zz_10873 = _zz_10874;
  assign _zz_10874 = ($signed(_zz_905) + $signed(_zz_2933));
  assign _zz_10875 = _zz_10876;
  assign _zz_10876 = ($signed(_zz_10877) >>> _zz_2937);
  assign _zz_10877 = _zz_10878;
  assign _zz_10878 = ($signed(_zz_906) + $signed(_zz_2934));
  assign _zz_10879 = ($signed(twiddle_factor_table_12_real) + $signed(twiddle_factor_table_12_imag));
  assign _zz_10880 = fixTo_687_dout;
  assign _zz_10881 = ($signed(_zz_924) - $signed(_zz_923));
  assign _zz_10882 = ($signed(_zz_923) + $signed(_zz_924));
  assign _zz_10883 = _zz_10884[15 : 0];
  assign _zz_10884 = fixTo_689_dout;
  assign _zz_10885 = _zz_10886[15 : 0];
  assign _zz_10886 = fixTo_688_dout;
  assign _zz_10887 = _zz_10888;
  assign _zz_10888 = ($signed(_zz_10889) >>> _zz_2941);
  assign _zz_10889 = _zz_10890;
  assign _zz_10890 = ($signed(_zz_907) - $signed(_zz_2938));
  assign _zz_10891 = _zz_10892;
  assign _zz_10892 = ($signed(_zz_10893) >>> _zz_2941);
  assign _zz_10893 = _zz_10894;
  assign _zz_10894 = ($signed(_zz_908) - $signed(_zz_2939));
  assign _zz_10895 = _zz_10896;
  assign _zz_10896 = ($signed(_zz_10897) >>> _zz_2942);
  assign _zz_10897 = _zz_10898;
  assign _zz_10898 = ($signed(_zz_907) + $signed(_zz_2938));
  assign _zz_10899 = _zz_10900;
  assign _zz_10900 = ($signed(_zz_10901) >>> _zz_2942);
  assign _zz_10901 = _zz_10902;
  assign _zz_10902 = ($signed(_zz_908) + $signed(_zz_2939));
  assign _zz_10903 = ($signed(twiddle_factor_table_13_real) + $signed(twiddle_factor_table_13_imag));
  assign _zz_10904 = fixTo_690_dout;
  assign _zz_10905 = ($signed(_zz_926) - $signed(_zz_925));
  assign _zz_10906 = ($signed(_zz_925) + $signed(_zz_926));
  assign _zz_10907 = _zz_10908[15 : 0];
  assign _zz_10908 = fixTo_692_dout;
  assign _zz_10909 = _zz_10910[15 : 0];
  assign _zz_10910 = fixTo_691_dout;
  assign _zz_10911 = _zz_10912;
  assign _zz_10912 = ($signed(_zz_10913) >>> _zz_2946);
  assign _zz_10913 = _zz_10914;
  assign _zz_10914 = ($signed(_zz_909) - $signed(_zz_2943));
  assign _zz_10915 = _zz_10916;
  assign _zz_10916 = ($signed(_zz_10917) >>> _zz_2946);
  assign _zz_10917 = _zz_10918;
  assign _zz_10918 = ($signed(_zz_910) - $signed(_zz_2944));
  assign _zz_10919 = _zz_10920;
  assign _zz_10920 = ($signed(_zz_10921) >>> _zz_2947);
  assign _zz_10921 = _zz_10922;
  assign _zz_10922 = ($signed(_zz_909) + $signed(_zz_2943));
  assign _zz_10923 = _zz_10924;
  assign _zz_10924 = ($signed(_zz_10925) >>> _zz_2947);
  assign _zz_10925 = _zz_10926;
  assign _zz_10926 = ($signed(_zz_910) + $signed(_zz_2944));
  assign _zz_10927 = ($signed(twiddle_factor_table_14_real) + $signed(twiddle_factor_table_14_imag));
  assign _zz_10928 = fixTo_693_dout;
  assign _zz_10929 = ($signed(_zz_928) - $signed(_zz_927));
  assign _zz_10930 = ($signed(_zz_927) + $signed(_zz_928));
  assign _zz_10931 = _zz_10932[15 : 0];
  assign _zz_10932 = fixTo_695_dout;
  assign _zz_10933 = _zz_10934[15 : 0];
  assign _zz_10934 = fixTo_694_dout;
  assign _zz_10935 = _zz_10936;
  assign _zz_10936 = ($signed(_zz_10937) >>> _zz_2951);
  assign _zz_10937 = _zz_10938;
  assign _zz_10938 = ($signed(_zz_911) - $signed(_zz_2948));
  assign _zz_10939 = _zz_10940;
  assign _zz_10940 = ($signed(_zz_10941) >>> _zz_2951);
  assign _zz_10941 = _zz_10942;
  assign _zz_10942 = ($signed(_zz_912) - $signed(_zz_2949));
  assign _zz_10943 = _zz_10944;
  assign _zz_10944 = ($signed(_zz_10945) >>> _zz_2952);
  assign _zz_10945 = _zz_10946;
  assign _zz_10946 = ($signed(_zz_911) + $signed(_zz_2948));
  assign _zz_10947 = _zz_10948;
  assign _zz_10948 = ($signed(_zz_10949) >>> _zz_2952);
  assign _zz_10949 = _zz_10950;
  assign _zz_10950 = ($signed(_zz_912) + $signed(_zz_2949));
  assign _zz_10951 = ($signed(twiddle_factor_table_7_real) + $signed(twiddle_factor_table_7_imag));
  assign _zz_10952 = fixTo_696_dout;
  assign _zz_10953 = ($signed(_zz_946) - $signed(_zz_945));
  assign _zz_10954 = ($signed(_zz_945) + $signed(_zz_946));
  assign _zz_10955 = _zz_10956[15 : 0];
  assign _zz_10956 = fixTo_698_dout;
  assign _zz_10957 = _zz_10958[15 : 0];
  assign _zz_10958 = fixTo_697_dout;
  assign _zz_10959 = _zz_10960;
  assign _zz_10960 = ($signed(_zz_10961) >>> _zz_2956);
  assign _zz_10961 = _zz_10962;
  assign _zz_10962 = ($signed(_zz_929) - $signed(_zz_2953));
  assign _zz_10963 = _zz_10964;
  assign _zz_10964 = ($signed(_zz_10965) >>> _zz_2956);
  assign _zz_10965 = _zz_10966;
  assign _zz_10966 = ($signed(_zz_930) - $signed(_zz_2954));
  assign _zz_10967 = _zz_10968;
  assign _zz_10968 = ($signed(_zz_10969) >>> _zz_2957);
  assign _zz_10969 = _zz_10970;
  assign _zz_10970 = ($signed(_zz_929) + $signed(_zz_2953));
  assign _zz_10971 = _zz_10972;
  assign _zz_10972 = ($signed(_zz_10973) >>> _zz_2957);
  assign _zz_10973 = _zz_10974;
  assign _zz_10974 = ($signed(_zz_930) + $signed(_zz_2954));
  assign _zz_10975 = ($signed(twiddle_factor_table_8_real) + $signed(twiddle_factor_table_8_imag));
  assign _zz_10976 = fixTo_699_dout;
  assign _zz_10977 = ($signed(_zz_948) - $signed(_zz_947));
  assign _zz_10978 = ($signed(_zz_947) + $signed(_zz_948));
  assign _zz_10979 = _zz_10980[15 : 0];
  assign _zz_10980 = fixTo_701_dout;
  assign _zz_10981 = _zz_10982[15 : 0];
  assign _zz_10982 = fixTo_700_dout;
  assign _zz_10983 = _zz_10984;
  assign _zz_10984 = ($signed(_zz_10985) >>> _zz_2961);
  assign _zz_10985 = _zz_10986;
  assign _zz_10986 = ($signed(_zz_931) - $signed(_zz_2958));
  assign _zz_10987 = _zz_10988;
  assign _zz_10988 = ($signed(_zz_10989) >>> _zz_2961);
  assign _zz_10989 = _zz_10990;
  assign _zz_10990 = ($signed(_zz_932) - $signed(_zz_2959));
  assign _zz_10991 = _zz_10992;
  assign _zz_10992 = ($signed(_zz_10993) >>> _zz_2962);
  assign _zz_10993 = _zz_10994;
  assign _zz_10994 = ($signed(_zz_931) + $signed(_zz_2958));
  assign _zz_10995 = _zz_10996;
  assign _zz_10996 = ($signed(_zz_10997) >>> _zz_2962);
  assign _zz_10997 = _zz_10998;
  assign _zz_10998 = ($signed(_zz_932) + $signed(_zz_2959));
  assign _zz_10999 = ($signed(twiddle_factor_table_9_real) + $signed(twiddle_factor_table_9_imag));
  assign _zz_11000 = fixTo_702_dout;
  assign _zz_11001 = ($signed(_zz_950) - $signed(_zz_949));
  assign _zz_11002 = ($signed(_zz_949) + $signed(_zz_950));
  assign _zz_11003 = _zz_11004[15 : 0];
  assign _zz_11004 = fixTo_704_dout;
  assign _zz_11005 = _zz_11006[15 : 0];
  assign _zz_11006 = fixTo_703_dout;
  assign _zz_11007 = _zz_11008;
  assign _zz_11008 = ($signed(_zz_11009) >>> _zz_2966);
  assign _zz_11009 = _zz_11010;
  assign _zz_11010 = ($signed(_zz_933) - $signed(_zz_2963));
  assign _zz_11011 = _zz_11012;
  assign _zz_11012 = ($signed(_zz_11013) >>> _zz_2966);
  assign _zz_11013 = _zz_11014;
  assign _zz_11014 = ($signed(_zz_934) - $signed(_zz_2964));
  assign _zz_11015 = _zz_11016;
  assign _zz_11016 = ($signed(_zz_11017) >>> _zz_2967);
  assign _zz_11017 = _zz_11018;
  assign _zz_11018 = ($signed(_zz_933) + $signed(_zz_2963));
  assign _zz_11019 = _zz_11020;
  assign _zz_11020 = ($signed(_zz_11021) >>> _zz_2967);
  assign _zz_11021 = _zz_11022;
  assign _zz_11022 = ($signed(_zz_934) + $signed(_zz_2964));
  assign _zz_11023 = ($signed(twiddle_factor_table_10_real) + $signed(twiddle_factor_table_10_imag));
  assign _zz_11024 = fixTo_705_dout;
  assign _zz_11025 = ($signed(_zz_952) - $signed(_zz_951));
  assign _zz_11026 = ($signed(_zz_951) + $signed(_zz_952));
  assign _zz_11027 = _zz_11028[15 : 0];
  assign _zz_11028 = fixTo_707_dout;
  assign _zz_11029 = _zz_11030[15 : 0];
  assign _zz_11030 = fixTo_706_dout;
  assign _zz_11031 = _zz_11032;
  assign _zz_11032 = ($signed(_zz_11033) >>> _zz_2971);
  assign _zz_11033 = _zz_11034;
  assign _zz_11034 = ($signed(_zz_935) - $signed(_zz_2968));
  assign _zz_11035 = _zz_11036;
  assign _zz_11036 = ($signed(_zz_11037) >>> _zz_2971);
  assign _zz_11037 = _zz_11038;
  assign _zz_11038 = ($signed(_zz_936) - $signed(_zz_2969));
  assign _zz_11039 = _zz_11040;
  assign _zz_11040 = ($signed(_zz_11041) >>> _zz_2972);
  assign _zz_11041 = _zz_11042;
  assign _zz_11042 = ($signed(_zz_935) + $signed(_zz_2968));
  assign _zz_11043 = _zz_11044;
  assign _zz_11044 = ($signed(_zz_11045) >>> _zz_2972);
  assign _zz_11045 = _zz_11046;
  assign _zz_11046 = ($signed(_zz_936) + $signed(_zz_2969));
  assign _zz_11047 = ($signed(twiddle_factor_table_11_real) + $signed(twiddle_factor_table_11_imag));
  assign _zz_11048 = fixTo_708_dout;
  assign _zz_11049 = ($signed(_zz_954) - $signed(_zz_953));
  assign _zz_11050 = ($signed(_zz_953) + $signed(_zz_954));
  assign _zz_11051 = _zz_11052[15 : 0];
  assign _zz_11052 = fixTo_710_dout;
  assign _zz_11053 = _zz_11054[15 : 0];
  assign _zz_11054 = fixTo_709_dout;
  assign _zz_11055 = _zz_11056;
  assign _zz_11056 = ($signed(_zz_11057) >>> _zz_2976);
  assign _zz_11057 = _zz_11058;
  assign _zz_11058 = ($signed(_zz_937) - $signed(_zz_2973));
  assign _zz_11059 = _zz_11060;
  assign _zz_11060 = ($signed(_zz_11061) >>> _zz_2976);
  assign _zz_11061 = _zz_11062;
  assign _zz_11062 = ($signed(_zz_938) - $signed(_zz_2974));
  assign _zz_11063 = _zz_11064;
  assign _zz_11064 = ($signed(_zz_11065) >>> _zz_2977);
  assign _zz_11065 = _zz_11066;
  assign _zz_11066 = ($signed(_zz_937) + $signed(_zz_2973));
  assign _zz_11067 = _zz_11068;
  assign _zz_11068 = ($signed(_zz_11069) >>> _zz_2977);
  assign _zz_11069 = _zz_11070;
  assign _zz_11070 = ($signed(_zz_938) + $signed(_zz_2974));
  assign _zz_11071 = ($signed(twiddle_factor_table_12_real) + $signed(twiddle_factor_table_12_imag));
  assign _zz_11072 = fixTo_711_dout;
  assign _zz_11073 = ($signed(_zz_956) - $signed(_zz_955));
  assign _zz_11074 = ($signed(_zz_955) + $signed(_zz_956));
  assign _zz_11075 = _zz_11076[15 : 0];
  assign _zz_11076 = fixTo_713_dout;
  assign _zz_11077 = _zz_11078[15 : 0];
  assign _zz_11078 = fixTo_712_dout;
  assign _zz_11079 = _zz_11080;
  assign _zz_11080 = ($signed(_zz_11081) >>> _zz_2981);
  assign _zz_11081 = _zz_11082;
  assign _zz_11082 = ($signed(_zz_939) - $signed(_zz_2978));
  assign _zz_11083 = _zz_11084;
  assign _zz_11084 = ($signed(_zz_11085) >>> _zz_2981);
  assign _zz_11085 = _zz_11086;
  assign _zz_11086 = ($signed(_zz_940) - $signed(_zz_2979));
  assign _zz_11087 = _zz_11088;
  assign _zz_11088 = ($signed(_zz_11089) >>> _zz_2982);
  assign _zz_11089 = _zz_11090;
  assign _zz_11090 = ($signed(_zz_939) + $signed(_zz_2978));
  assign _zz_11091 = _zz_11092;
  assign _zz_11092 = ($signed(_zz_11093) >>> _zz_2982);
  assign _zz_11093 = _zz_11094;
  assign _zz_11094 = ($signed(_zz_940) + $signed(_zz_2979));
  assign _zz_11095 = ($signed(twiddle_factor_table_13_real) + $signed(twiddle_factor_table_13_imag));
  assign _zz_11096 = fixTo_714_dout;
  assign _zz_11097 = ($signed(_zz_958) - $signed(_zz_957));
  assign _zz_11098 = ($signed(_zz_957) + $signed(_zz_958));
  assign _zz_11099 = _zz_11100[15 : 0];
  assign _zz_11100 = fixTo_716_dout;
  assign _zz_11101 = _zz_11102[15 : 0];
  assign _zz_11102 = fixTo_715_dout;
  assign _zz_11103 = _zz_11104;
  assign _zz_11104 = ($signed(_zz_11105) >>> _zz_2986);
  assign _zz_11105 = _zz_11106;
  assign _zz_11106 = ($signed(_zz_941) - $signed(_zz_2983));
  assign _zz_11107 = _zz_11108;
  assign _zz_11108 = ($signed(_zz_11109) >>> _zz_2986);
  assign _zz_11109 = _zz_11110;
  assign _zz_11110 = ($signed(_zz_942) - $signed(_zz_2984));
  assign _zz_11111 = _zz_11112;
  assign _zz_11112 = ($signed(_zz_11113) >>> _zz_2987);
  assign _zz_11113 = _zz_11114;
  assign _zz_11114 = ($signed(_zz_941) + $signed(_zz_2983));
  assign _zz_11115 = _zz_11116;
  assign _zz_11116 = ($signed(_zz_11117) >>> _zz_2987);
  assign _zz_11117 = _zz_11118;
  assign _zz_11118 = ($signed(_zz_942) + $signed(_zz_2984));
  assign _zz_11119 = ($signed(twiddle_factor_table_14_real) + $signed(twiddle_factor_table_14_imag));
  assign _zz_11120 = fixTo_717_dout;
  assign _zz_11121 = ($signed(_zz_960) - $signed(_zz_959));
  assign _zz_11122 = ($signed(_zz_959) + $signed(_zz_960));
  assign _zz_11123 = _zz_11124[15 : 0];
  assign _zz_11124 = fixTo_719_dout;
  assign _zz_11125 = _zz_11126[15 : 0];
  assign _zz_11126 = fixTo_718_dout;
  assign _zz_11127 = _zz_11128;
  assign _zz_11128 = ($signed(_zz_11129) >>> _zz_2991);
  assign _zz_11129 = _zz_11130;
  assign _zz_11130 = ($signed(_zz_943) - $signed(_zz_2988));
  assign _zz_11131 = _zz_11132;
  assign _zz_11132 = ($signed(_zz_11133) >>> _zz_2991);
  assign _zz_11133 = _zz_11134;
  assign _zz_11134 = ($signed(_zz_944) - $signed(_zz_2989));
  assign _zz_11135 = _zz_11136;
  assign _zz_11136 = ($signed(_zz_11137) >>> _zz_2992);
  assign _zz_11137 = _zz_11138;
  assign _zz_11138 = ($signed(_zz_943) + $signed(_zz_2988));
  assign _zz_11139 = _zz_11140;
  assign _zz_11140 = ($signed(_zz_11141) >>> _zz_2992);
  assign _zz_11141 = _zz_11142;
  assign _zz_11142 = ($signed(_zz_944) + $signed(_zz_2989));
  assign _zz_11143 = ($signed(twiddle_factor_table_7_real) + $signed(twiddle_factor_table_7_imag));
  assign _zz_11144 = fixTo_720_dout;
  assign _zz_11145 = ($signed(_zz_978) - $signed(_zz_977));
  assign _zz_11146 = ($signed(_zz_977) + $signed(_zz_978));
  assign _zz_11147 = _zz_11148[15 : 0];
  assign _zz_11148 = fixTo_722_dout;
  assign _zz_11149 = _zz_11150[15 : 0];
  assign _zz_11150 = fixTo_721_dout;
  assign _zz_11151 = _zz_11152;
  assign _zz_11152 = ($signed(_zz_11153) >>> _zz_2996);
  assign _zz_11153 = _zz_11154;
  assign _zz_11154 = ($signed(_zz_961) - $signed(_zz_2993));
  assign _zz_11155 = _zz_11156;
  assign _zz_11156 = ($signed(_zz_11157) >>> _zz_2996);
  assign _zz_11157 = _zz_11158;
  assign _zz_11158 = ($signed(_zz_962) - $signed(_zz_2994));
  assign _zz_11159 = _zz_11160;
  assign _zz_11160 = ($signed(_zz_11161) >>> _zz_2997);
  assign _zz_11161 = _zz_11162;
  assign _zz_11162 = ($signed(_zz_961) + $signed(_zz_2993));
  assign _zz_11163 = _zz_11164;
  assign _zz_11164 = ($signed(_zz_11165) >>> _zz_2997);
  assign _zz_11165 = _zz_11166;
  assign _zz_11166 = ($signed(_zz_962) + $signed(_zz_2994));
  assign _zz_11167 = ($signed(twiddle_factor_table_8_real) + $signed(twiddle_factor_table_8_imag));
  assign _zz_11168 = fixTo_723_dout;
  assign _zz_11169 = ($signed(_zz_980) - $signed(_zz_979));
  assign _zz_11170 = ($signed(_zz_979) + $signed(_zz_980));
  assign _zz_11171 = _zz_11172[15 : 0];
  assign _zz_11172 = fixTo_725_dout;
  assign _zz_11173 = _zz_11174[15 : 0];
  assign _zz_11174 = fixTo_724_dout;
  assign _zz_11175 = _zz_11176;
  assign _zz_11176 = ($signed(_zz_11177) >>> _zz_3001);
  assign _zz_11177 = _zz_11178;
  assign _zz_11178 = ($signed(_zz_963) - $signed(_zz_2998));
  assign _zz_11179 = _zz_11180;
  assign _zz_11180 = ($signed(_zz_11181) >>> _zz_3001);
  assign _zz_11181 = _zz_11182;
  assign _zz_11182 = ($signed(_zz_964) - $signed(_zz_2999));
  assign _zz_11183 = _zz_11184;
  assign _zz_11184 = ($signed(_zz_11185) >>> _zz_3002);
  assign _zz_11185 = _zz_11186;
  assign _zz_11186 = ($signed(_zz_963) + $signed(_zz_2998));
  assign _zz_11187 = _zz_11188;
  assign _zz_11188 = ($signed(_zz_11189) >>> _zz_3002);
  assign _zz_11189 = _zz_11190;
  assign _zz_11190 = ($signed(_zz_964) + $signed(_zz_2999));
  assign _zz_11191 = ($signed(twiddle_factor_table_9_real) + $signed(twiddle_factor_table_9_imag));
  assign _zz_11192 = fixTo_726_dout;
  assign _zz_11193 = ($signed(_zz_982) - $signed(_zz_981));
  assign _zz_11194 = ($signed(_zz_981) + $signed(_zz_982));
  assign _zz_11195 = _zz_11196[15 : 0];
  assign _zz_11196 = fixTo_728_dout;
  assign _zz_11197 = _zz_11198[15 : 0];
  assign _zz_11198 = fixTo_727_dout;
  assign _zz_11199 = _zz_11200;
  assign _zz_11200 = ($signed(_zz_11201) >>> _zz_3006);
  assign _zz_11201 = _zz_11202;
  assign _zz_11202 = ($signed(_zz_965) - $signed(_zz_3003));
  assign _zz_11203 = _zz_11204;
  assign _zz_11204 = ($signed(_zz_11205) >>> _zz_3006);
  assign _zz_11205 = _zz_11206;
  assign _zz_11206 = ($signed(_zz_966) - $signed(_zz_3004));
  assign _zz_11207 = _zz_11208;
  assign _zz_11208 = ($signed(_zz_11209) >>> _zz_3007);
  assign _zz_11209 = _zz_11210;
  assign _zz_11210 = ($signed(_zz_965) + $signed(_zz_3003));
  assign _zz_11211 = _zz_11212;
  assign _zz_11212 = ($signed(_zz_11213) >>> _zz_3007);
  assign _zz_11213 = _zz_11214;
  assign _zz_11214 = ($signed(_zz_966) + $signed(_zz_3004));
  assign _zz_11215 = ($signed(twiddle_factor_table_10_real) + $signed(twiddle_factor_table_10_imag));
  assign _zz_11216 = fixTo_729_dout;
  assign _zz_11217 = ($signed(_zz_984) - $signed(_zz_983));
  assign _zz_11218 = ($signed(_zz_983) + $signed(_zz_984));
  assign _zz_11219 = _zz_11220[15 : 0];
  assign _zz_11220 = fixTo_731_dout;
  assign _zz_11221 = _zz_11222[15 : 0];
  assign _zz_11222 = fixTo_730_dout;
  assign _zz_11223 = _zz_11224;
  assign _zz_11224 = ($signed(_zz_11225) >>> _zz_3011);
  assign _zz_11225 = _zz_11226;
  assign _zz_11226 = ($signed(_zz_967) - $signed(_zz_3008));
  assign _zz_11227 = _zz_11228;
  assign _zz_11228 = ($signed(_zz_11229) >>> _zz_3011);
  assign _zz_11229 = _zz_11230;
  assign _zz_11230 = ($signed(_zz_968) - $signed(_zz_3009));
  assign _zz_11231 = _zz_11232;
  assign _zz_11232 = ($signed(_zz_11233) >>> _zz_3012);
  assign _zz_11233 = _zz_11234;
  assign _zz_11234 = ($signed(_zz_967) + $signed(_zz_3008));
  assign _zz_11235 = _zz_11236;
  assign _zz_11236 = ($signed(_zz_11237) >>> _zz_3012);
  assign _zz_11237 = _zz_11238;
  assign _zz_11238 = ($signed(_zz_968) + $signed(_zz_3009));
  assign _zz_11239 = ($signed(twiddle_factor_table_11_real) + $signed(twiddle_factor_table_11_imag));
  assign _zz_11240 = fixTo_732_dout;
  assign _zz_11241 = ($signed(_zz_986) - $signed(_zz_985));
  assign _zz_11242 = ($signed(_zz_985) + $signed(_zz_986));
  assign _zz_11243 = _zz_11244[15 : 0];
  assign _zz_11244 = fixTo_734_dout;
  assign _zz_11245 = _zz_11246[15 : 0];
  assign _zz_11246 = fixTo_733_dout;
  assign _zz_11247 = _zz_11248;
  assign _zz_11248 = ($signed(_zz_11249) >>> _zz_3016);
  assign _zz_11249 = _zz_11250;
  assign _zz_11250 = ($signed(_zz_969) - $signed(_zz_3013));
  assign _zz_11251 = _zz_11252;
  assign _zz_11252 = ($signed(_zz_11253) >>> _zz_3016);
  assign _zz_11253 = _zz_11254;
  assign _zz_11254 = ($signed(_zz_970) - $signed(_zz_3014));
  assign _zz_11255 = _zz_11256;
  assign _zz_11256 = ($signed(_zz_11257) >>> _zz_3017);
  assign _zz_11257 = _zz_11258;
  assign _zz_11258 = ($signed(_zz_969) + $signed(_zz_3013));
  assign _zz_11259 = _zz_11260;
  assign _zz_11260 = ($signed(_zz_11261) >>> _zz_3017);
  assign _zz_11261 = _zz_11262;
  assign _zz_11262 = ($signed(_zz_970) + $signed(_zz_3014));
  assign _zz_11263 = ($signed(twiddle_factor_table_12_real) + $signed(twiddle_factor_table_12_imag));
  assign _zz_11264 = fixTo_735_dout;
  assign _zz_11265 = ($signed(_zz_988) - $signed(_zz_987));
  assign _zz_11266 = ($signed(_zz_987) + $signed(_zz_988));
  assign _zz_11267 = _zz_11268[15 : 0];
  assign _zz_11268 = fixTo_737_dout;
  assign _zz_11269 = _zz_11270[15 : 0];
  assign _zz_11270 = fixTo_736_dout;
  assign _zz_11271 = _zz_11272;
  assign _zz_11272 = ($signed(_zz_11273) >>> _zz_3021);
  assign _zz_11273 = _zz_11274;
  assign _zz_11274 = ($signed(_zz_971) - $signed(_zz_3018));
  assign _zz_11275 = _zz_11276;
  assign _zz_11276 = ($signed(_zz_11277) >>> _zz_3021);
  assign _zz_11277 = _zz_11278;
  assign _zz_11278 = ($signed(_zz_972) - $signed(_zz_3019));
  assign _zz_11279 = _zz_11280;
  assign _zz_11280 = ($signed(_zz_11281) >>> _zz_3022);
  assign _zz_11281 = _zz_11282;
  assign _zz_11282 = ($signed(_zz_971) + $signed(_zz_3018));
  assign _zz_11283 = _zz_11284;
  assign _zz_11284 = ($signed(_zz_11285) >>> _zz_3022);
  assign _zz_11285 = _zz_11286;
  assign _zz_11286 = ($signed(_zz_972) + $signed(_zz_3019));
  assign _zz_11287 = ($signed(twiddle_factor_table_13_real) + $signed(twiddle_factor_table_13_imag));
  assign _zz_11288 = fixTo_738_dout;
  assign _zz_11289 = ($signed(_zz_990) - $signed(_zz_989));
  assign _zz_11290 = ($signed(_zz_989) + $signed(_zz_990));
  assign _zz_11291 = _zz_11292[15 : 0];
  assign _zz_11292 = fixTo_740_dout;
  assign _zz_11293 = _zz_11294[15 : 0];
  assign _zz_11294 = fixTo_739_dout;
  assign _zz_11295 = _zz_11296;
  assign _zz_11296 = ($signed(_zz_11297) >>> _zz_3026);
  assign _zz_11297 = _zz_11298;
  assign _zz_11298 = ($signed(_zz_973) - $signed(_zz_3023));
  assign _zz_11299 = _zz_11300;
  assign _zz_11300 = ($signed(_zz_11301) >>> _zz_3026);
  assign _zz_11301 = _zz_11302;
  assign _zz_11302 = ($signed(_zz_974) - $signed(_zz_3024));
  assign _zz_11303 = _zz_11304;
  assign _zz_11304 = ($signed(_zz_11305) >>> _zz_3027);
  assign _zz_11305 = _zz_11306;
  assign _zz_11306 = ($signed(_zz_973) + $signed(_zz_3023));
  assign _zz_11307 = _zz_11308;
  assign _zz_11308 = ($signed(_zz_11309) >>> _zz_3027);
  assign _zz_11309 = _zz_11310;
  assign _zz_11310 = ($signed(_zz_974) + $signed(_zz_3024));
  assign _zz_11311 = ($signed(twiddle_factor_table_14_real) + $signed(twiddle_factor_table_14_imag));
  assign _zz_11312 = fixTo_741_dout;
  assign _zz_11313 = ($signed(_zz_992) - $signed(_zz_991));
  assign _zz_11314 = ($signed(_zz_991) + $signed(_zz_992));
  assign _zz_11315 = _zz_11316[15 : 0];
  assign _zz_11316 = fixTo_743_dout;
  assign _zz_11317 = _zz_11318[15 : 0];
  assign _zz_11318 = fixTo_742_dout;
  assign _zz_11319 = _zz_11320;
  assign _zz_11320 = ($signed(_zz_11321) >>> _zz_3031);
  assign _zz_11321 = _zz_11322;
  assign _zz_11322 = ($signed(_zz_975) - $signed(_zz_3028));
  assign _zz_11323 = _zz_11324;
  assign _zz_11324 = ($signed(_zz_11325) >>> _zz_3031);
  assign _zz_11325 = _zz_11326;
  assign _zz_11326 = ($signed(_zz_976) - $signed(_zz_3029));
  assign _zz_11327 = _zz_11328;
  assign _zz_11328 = ($signed(_zz_11329) >>> _zz_3032);
  assign _zz_11329 = _zz_11330;
  assign _zz_11330 = ($signed(_zz_975) + $signed(_zz_3028));
  assign _zz_11331 = _zz_11332;
  assign _zz_11332 = ($signed(_zz_11333) >>> _zz_3032);
  assign _zz_11333 = _zz_11334;
  assign _zz_11334 = ($signed(_zz_976) + $signed(_zz_3029));
  assign _zz_11335 = ($signed(twiddle_factor_table_7_real) + $signed(twiddle_factor_table_7_imag));
  assign _zz_11336 = fixTo_744_dout;
  assign _zz_11337 = ($signed(_zz_1010) - $signed(_zz_1009));
  assign _zz_11338 = ($signed(_zz_1009) + $signed(_zz_1010));
  assign _zz_11339 = _zz_11340[15 : 0];
  assign _zz_11340 = fixTo_746_dout;
  assign _zz_11341 = _zz_11342[15 : 0];
  assign _zz_11342 = fixTo_745_dout;
  assign _zz_11343 = _zz_11344;
  assign _zz_11344 = ($signed(_zz_11345) >>> _zz_3036);
  assign _zz_11345 = _zz_11346;
  assign _zz_11346 = ($signed(_zz_993) - $signed(_zz_3033));
  assign _zz_11347 = _zz_11348;
  assign _zz_11348 = ($signed(_zz_11349) >>> _zz_3036);
  assign _zz_11349 = _zz_11350;
  assign _zz_11350 = ($signed(_zz_994) - $signed(_zz_3034));
  assign _zz_11351 = _zz_11352;
  assign _zz_11352 = ($signed(_zz_11353) >>> _zz_3037);
  assign _zz_11353 = _zz_11354;
  assign _zz_11354 = ($signed(_zz_993) + $signed(_zz_3033));
  assign _zz_11355 = _zz_11356;
  assign _zz_11356 = ($signed(_zz_11357) >>> _zz_3037);
  assign _zz_11357 = _zz_11358;
  assign _zz_11358 = ($signed(_zz_994) + $signed(_zz_3034));
  assign _zz_11359 = ($signed(twiddle_factor_table_8_real) + $signed(twiddle_factor_table_8_imag));
  assign _zz_11360 = fixTo_747_dout;
  assign _zz_11361 = ($signed(_zz_1012) - $signed(_zz_1011));
  assign _zz_11362 = ($signed(_zz_1011) + $signed(_zz_1012));
  assign _zz_11363 = _zz_11364[15 : 0];
  assign _zz_11364 = fixTo_749_dout;
  assign _zz_11365 = _zz_11366[15 : 0];
  assign _zz_11366 = fixTo_748_dout;
  assign _zz_11367 = _zz_11368;
  assign _zz_11368 = ($signed(_zz_11369) >>> _zz_3041);
  assign _zz_11369 = _zz_11370;
  assign _zz_11370 = ($signed(_zz_995) - $signed(_zz_3038));
  assign _zz_11371 = _zz_11372;
  assign _zz_11372 = ($signed(_zz_11373) >>> _zz_3041);
  assign _zz_11373 = _zz_11374;
  assign _zz_11374 = ($signed(_zz_996) - $signed(_zz_3039));
  assign _zz_11375 = _zz_11376;
  assign _zz_11376 = ($signed(_zz_11377) >>> _zz_3042);
  assign _zz_11377 = _zz_11378;
  assign _zz_11378 = ($signed(_zz_995) + $signed(_zz_3038));
  assign _zz_11379 = _zz_11380;
  assign _zz_11380 = ($signed(_zz_11381) >>> _zz_3042);
  assign _zz_11381 = _zz_11382;
  assign _zz_11382 = ($signed(_zz_996) + $signed(_zz_3039));
  assign _zz_11383 = ($signed(twiddle_factor_table_9_real) + $signed(twiddle_factor_table_9_imag));
  assign _zz_11384 = fixTo_750_dout;
  assign _zz_11385 = ($signed(_zz_1014) - $signed(_zz_1013));
  assign _zz_11386 = ($signed(_zz_1013) + $signed(_zz_1014));
  assign _zz_11387 = _zz_11388[15 : 0];
  assign _zz_11388 = fixTo_752_dout;
  assign _zz_11389 = _zz_11390[15 : 0];
  assign _zz_11390 = fixTo_751_dout;
  assign _zz_11391 = _zz_11392;
  assign _zz_11392 = ($signed(_zz_11393) >>> _zz_3046);
  assign _zz_11393 = _zz_11394;
  assign _zz_11394 = ($signed(_zz_997) - $signed(_zz_3043));
  assign _zz_11395 = _zz_11396;
  assign _zz_11396 = ($signed(_zz_11397) >>> _zz_3046);
  assign _zz_11397 = _zz_11398;
  assign _zz_11398 = ($signed(_zz_998) - $signed(_zz_3044));
  assign _zz_11399 = _zz_11400;
  assign _zz_11400 = ($signed(_zz_11401) >>> _zz_3047);
  assign _zz_11401 = _zz_11402;
  assign _zz_11402 = ($signed(_zz_997) + $signed(_zz_3043));
  assign _zz_11403 = _zz_11404;
  assign _zz_11404 = ($signed(_zz_11405) >>> _zz_3047);
  assign _zz_11405 = _zz_11406;
  assign _zz_11406 = ($signed(_zz_998) + $signed(_zz_3044));
  assign _zz_11407 = ($signed(twiddle_factor_table_10_real) + $signed(twiddle_factor_table_10_imag));
  assign _zz_11408 = fixTo_753_dout;
  assign _zz_11409 = ($signed(_zz_1016) - $signed(_zz_1015));
  assign _zz_11410 = ($signed(_zz_1015) + $signed(_zz_1016));
  assign _zz_11411 = _zz_11412[15 : 0];
  assign _zz_11412 = fixTo_755_dout;
  assign _zz_11413 = _zz_11414[15 : 0];
  assign _zz_11414 = fixTo_754_dout;
  assign _zz_11415 = _zz_11416;
  assign _zz_11416 = ($signed(_zz_11417) >>> _zz_3051);
  assign _zz_11417 = _zz_11418;
  assign _zz_11418 = ($signed(_zz_999) - $signed(_zz_3048));
  assign _zz_11419 = _zz_11420;
  assign _zz_11420 = ($signed(_zz_11421) >>> _zz_3051);
  assign _zz_11421 = _zz_11422;
  assign _zz_11422 = ($signed(_zz_1000) - $signed(_zz_3049));
  assign _zz_11423 = _zz_11424;
  assign _zz_11424 = ($signed(_zz_11425) >>> _zz_3052);
  assign _zz_11425 = _zz_11426;
  assign _zz_11426 = ($signed(_zz_999) + $signed(_zz_3048));
  assign _zz_11427 = _zz_11428;
  assign _zz_11428 = ($signed(_zz_11429) >>> _zz_3052);
  assign _zz_11429 = _zz_11430;
  assign _zz_11430 = ($signed(_zz_1000) + $signed(_zz_3049));
  assign _zz_11431 = ($signed(twiddle_factor_table_11_real) + $signed(twiddle_factor_table_11_imag));
  assign _zz_11432 = fixTo_756_dout;
  assign _zz_11433 = ($signed(_zz_1018) - $signed(_zz_1017));
  assign _zz_11434 = ($signed(_zz_1017) + $signed(_zz_1018));
  assign _zz_11435 = _zz_11436[15 : 0];
  assign _zz_11436 = fixTo_758_dout;
  assign _zz_11437 = _zz_11438[15 : 0];
  assign _zz_11438 = fixTo_757_dout;
  assign _zz_11439 = _zz_11440;
  assign _zz_11440 = ($signed(_zz_11441) >>> _zz_3056);
  assign _zz_11441 = _zz_11442;
  assign _zz_11442 = ($signed(_zz_1001) - $signed(_zz_3053));
  assign _zz_11443 = _zz_11444;
  assign _zz_11444 = ($signed(_zz_11445) >>> _zz_3056);
  assign _zz_11445 = _zz_11446;
  assign _zz_11446 = ($signed(_zz_1002) - $signed(_zz_3054));
  assign _zz_11447 = _zz_11448;
  assign _zz_11448 = ($signed(_zz_11449) >>> _zz_3057);
  assign _zz_11449 = _zz_11450;
  assign _zz_11450 = ($signed(_zz_1001) + $signed(_zz_3053));
  assign _zz_11451 = _zz_11452;
  assign _zz_11452 = ($signed(_zz_11453) >>> _zz_3057);
  assign _zz_11453 = _zz_11454;
  assign _zz_11454 = ($signed(_zz_1002) + $signed(_zz_3054));
  assign _zz_11455 = ($signed(twiddle_factor_table_12_real) + $signed(twiddle_factor_table_12_imag));
  assign _zz_11456 = fixTo_759_dout;
  assign _zz_11457 = ($signed(_zz_1020) - $signed(_zz_1019));
  assign _zz_11458 = ($signed(_zz_1019) + $signed(_zz_1020));
  assign _zz_11459 = _zz_11460[15 : 0];
  assign _zz_11460 = fixTo_761_dout;
  assign _zz_11461 = _zz_11462[15 : 0];
  assign _zz_11462 = fixTo_760_dout;
  assign _zz_11463 = _zz_11464;
  assign _zz_11464 = ($signed(_zz_11465) >>> _zz_3061);
  assign _zz_11465 = _zz_11466;
  assign _zz_11466 = ($signed(_zz_1003) - $signed(_zz_3058));
  assign _zz_11467 = _zz_11468;
  assign _zz_11468 = ($signed(_zz_11469) >>> _zz_3061);
  assign _zz_11469 = _zz_11470;
  assign _zz_11470 = ($signed(_zz_1004) - $signed(_zz_3059));
  assign _zz_11471 = _zz_11472;
  assign _zz_11472 = ($signed(_zz_11473) >>> _zz_3062);
  assign _zz_11473 = _zz_11474;
  assign _zz_11474 = ($signed(_zz_1003) + $signed(_zz_3058));
  assign _zz_11475 = _zz_11476;
  assign _zz_11476 = ($signed(_zz_11477) >>> _zz_3062);
  assign _zz_11477 = _zz_11478;
  assign _zz_11478 = ($signed(_zz_1004) + $signed(_zz_3059));
  assign _zz_11479 = ($signed(twiddle_factor_table_13_real) + $signed(twiddle_factor_table_13_imag));
  assign _zz_11480 = fixTo_762_dout;
  assign _zz_11481 = ($signed(_zz_1022) - $signed(_zz_1021));
  assign _zz_11482 = ($signed(_zz_1021) + $signed(_zz_1022));
  assign _zz_11483 = _zz_11484[15 : 0];
  assign _zz_11484 = fixTo_764_dout;
  assign _zz_11485 = _zz_11486[15 : 0];
  assign _zz_11486 = fixTo_763_dout;
  assign _zz_11487 = _zz_11488;
  assign _zz_11488 = ($signed(_zz_11489) >>> _zz_3066);
  assign _zz_11489 = _zz_11490;
  assign _zz_11490 = ($signed(_zz_1005) - $signed(_zz_3063));
  assign _zz_11491 = _zz_11492;
  assign _zz_11492 = ($signed(_zz_11493) >>> _zz_3066);
  assign _zz_11493 = _zz_11494;
  assign _zz_11494 = ($signed(_zz_1006) - $signed(_zz_3064));
  assign _zz_11495 = _zz_11496;
  assign _zz_11496 = ($signed(_zz_11497) >>> _zz_3067);
  assign _zz_11497 = _zz_11498;
  assign _zz_11498 = ($signed(_zz_1005) + $signed(_zz_3063));
  assign _zz_11499 = _zz_11500;
  assign _zz_11500 = ($signed(_zz_11501) >>> _zz_3067);
  assign _zz_11501 = _zz_11502;
  assign _zz_11502 = ($signed(_zz_1006) + $signed(_zz_3064));
  assign _zz_11503 = ($signed(twiddle_factor_table_14_real) + $signed(twiddle_factor_table_14_imag));
  assign _zz_11504 = fixTo_765_dout;
  assign _zz_11505 = ($signed(_zz_1024) - $signed(_zz_1023));
  assign _zz_11506 = ($signed(_zz_1023) + $signed(_zz_1024));
  assign _zz_11507 = _zz_11508[15 : 0];
  assign _zz_11508 = fixTo_767_dout;
  assign _zz_11509 = _zz_11510[15 : 0];
  assign _zz_11510 = fixTo_766_dout;
  assign _zz_11511 = _zz_11512;
  assign _zz_11512 = ($signed(_zz_11513) >>> _zz_3071);
  assign _zz_11513 = _zz_11514;
  assign _zz_11514 = ($signed(_zz_1007) - $signed(_zz_3068));
  assign _zz_11515 = _zz_11516;
  assign _zz_11516 = ($signed(_zz_11517) >>> _zz_3071);
  assign _zz_11517 = _zz_11518;
  assign _zz_11518 = ($signed(_zz_1008) - $signed(_zz_3069));
  assign _zz_11519 = _zz_11520;
  assign _zz_11520 = ($signed(_zz_11521) >>> _zz_3072);
  assign _zz_11521 = _zz_11522;
  assign _zz_11522 = ($signed(_zz_1007) + $signed(_zz_3068));
  assign _zz_11523 = _zz_11524;
  assign _zz_11524 = ($signed(_zz_11525) >>> _zz_3072);
  assign _zz_11525 = _zz_11526;
  assign _zz_11526 = ($signed(_zz_1008) + $signed(_zz_3069));
  assign _zz_11527 = ($signed(twiddle_factor_table_15_real) + $signed(twiddle_factor_table_15_imag));
  assign _zz_11528 = fixTo_768_dout;
  assign _zz_11529 = ($signed(_zz_1058) - $signed(_zz_1057));
  assign _zz_11530 = ($signed(_zz_1057) + $signed(_zz_1058));
  assign _zz_11531 = _zz_11532[15 : 0];
  assign _zz_11532 = fixTo_770_dout;
  assign _zz_11533 = _zz_11534[15 : 0];
  assign _zz_11534 = fixTo_769_dout;
  assign _zz_11535 = _zz_11536;
  assign _zz_11536 = ($signed(_zz_11537) >>> _zz_3076);
  assign _zz_11537 = _zz_11538;
  assign _zz_11538 = ($signed(_zz_1025) - $signed(_zz_3073));
  assign _zz_11539 = _zz_11540;
  assign _zz_11540 = ($signed(_zz_11541) >>> _zz_3076);
  assign _zz_11541 = _zz_11542;
  assign _zz_11542 = ($signed(_zz_1026) - $signed(_zz_3074));
  assign _zz_11543 = _zz_11544;
  assign _zz_11544 = ($signed(_zz_11545) >>> _zz_3077);
  assign _zz_11545 = _zz_11546;
  assign _zz_11546 = ($signed(_zz_1025) + $signed(_zz_3073));
  assign _zz_11547 = _zz_11548;
  assign _zz_11548 = ($signed(_zz_11549) >>> _zz_3077);
  assign _zz_11549 = _zz_11550;
  assign _zz_11550 = ($signed(_zz_1026) + $signed(_zz_3074));
  assign _zz_11551 = ($signed(twiddle_factor_table_16_real) + $signed(twiddle_factor_table_16_imag));
  assign _zz_11552 = fixTo_771_dout;
  assign _zz_11553 = ($signed(_zz_1060) - $signed(_zz_1059));
  assign _zz_11554 = ($signed(_zz_1059) + $signed(_zz_1060));
  assign _zz_11555 = _zz_11556[15 : 0];
  assign _zz_11556 = fixTo_773_dout;
  assign _zz_11557 = _zz_11558[15 : 0];
  assign _zz_11558 = fixTo_772_dout;
  assign _zz_11559 = _zz_11560;
  assign _zz_11560 = ($signed(_zz_11561) >>> _zz_3081);
  assign _zz_11561 = _zz_11562;
  assign _zz_11562 = ($signed(_zz_1027) - $signed(_zz_3078));
  assign _zz_11563 = _zz_11564;
  assign _zz_11564 = ($signed(_zz_11565) >>> _zz_3081);
  assign _zz_11565 = _zz_11566;
  assign _zz_11566 = ($signed(_zz_1028) - $signed(_zz_3079));
  assign _zz_11567 = _zz_11568;
  assign _zz_11568 = ($signed(_zz_11569) >>> _zz_3082);
  assign _zz_11569 = _zz_11570;
  assign _zz_11570 = ($signed(_zz_1027) + $signed(_zz_3078));
  assign _zz_11571 = _zz_11572;
  assign _zz_11572 = ($signed(_zz_11573) >>> _zz_3082);
  assign _zz_11573 = _zz_11574;
  assign _zz_11574 = ($signed(_zz_1028) + $signed(_zz_3079));
  assign _zz_11575 = ($signed(twiddle_factor_table_17_real) + $signed(twiddle_factor_table_17_imag));
  assign _zz_11576 = fixTo_774_dout;
  assign _zz_11577 = ($signed(_zz_1062) - $signed(_zz_1061));
  assign _zz_11578 = ($signed(_zz_1061) + $signed(_zz_1062));
  assign _zz_11579 = _zz_11580[15 : 0];
  assign _zz_11580 = fixTo_776_dout;
  assign _zz_11581 = _zz_11582[15 : 0];
  assign _zz_11582 = fixTo_775_dout;
  assign _zz_11583 = _zz_11584;
  assign _zz_11584 = ($signed(_zz_11585) >>> _zz_3086);
  assign _zz_11585 = _zz_11586;
  assign _zz_11586 = ($signed(_zz_1029) - $signed(_zz_3083));
  assign _zz_11587 = _zz_11588;
  assign _zz_11588 = ($signed(_zz_11589) >>> _zz_3086);
  assign _zz_11589 = _zz_11590;
  assign _zz_11590 = ($signed(_zz_1030) - $signed(_zz_3084));
  assign _zz_11591 = _zz_11592;
  assign _zz_11592 = ($signed(_zz_11593) >>> _zz_3087);
  assign _zz_11593 = _zz_11594;
  assign _zz_11594 = ($signed(_zz_1029) + $signed(_zz_3083));
  assign _zz_11595 = _zz_11596;
  assign _zz_11596 = ($signed(_zz_11597) >>> _zz_3087);
  assign _zz_11597 = _zz_11598;
  assign _zz_11598 = ($signed(_zz_1030) + $signed(_zz_3084));
  assign _zz_11599 = ($signed(twiddle_factor_table_18_real) + $signed(twiddle_factor_table_18_imag));
  assign _zz_11600 = fixTo_777_dout;
  assign _zz_11601 = ($signed(_zz_1064) - $signed(_zz_1063));
  assign _zz_11602 = ($signed(_zz_1063) + $signed(_zz_1064));
  assign _zz_11603 = _zz_11604[15 : 0];
  assign _zz_11604 = fixTo_779_dout;
  assign _zz_11605 = _zz_11606[15 : 0];
  assign _zz_11606 = fixTo_778_dout;
  assign _zz_11607 = _zz_11608;
  assign _zz_11608 = ($signed(_zz_11609) >>> _zz_3091);
  assign _zz_11609 = _zz_11610;
  assign _zz_11610 = ($signed(_zz_1031) - $signed(_zz_3088));
  assign _zz_11611 = _zz_11612;
  assign _zz_11612 = ($signed(_zz_11613) >>> _zz_3091);
  assign _zz_11613 = _zz_11614;
  assign _zz_11614 = ($signed(_zz_1032) - $signed(_zz_3089));
  assign _zz_11615 = _zz_11616;
  assign _zz_11616 = ($signed(_zz_11617) >>> _zz_3092);
  assign _zz_11617 = _zz_11618;
  assign _zz_11618 = ($signed(_zz_1031) + $signed(_zz_3088));
  assign _zz_11619 = _zz_11620;
  assign _zz_11620 = ($signed(_zz_11621) >>> _zz_3092);
  assign _zz_11621 = _zz_11622;
  assign _zz_11622 = ($signed(_zz_1032) + $signed(_zz_3089));
  assign _zz_11623 = ($signed(twiddle_factor_table_19_real) + $signed(twiddle_factor_table_19_imag));
  assign _zz_11624 = fixTo_780_dout;
  assign _zz_11625 = ($signed(_zz_1066) - $signed(_zz_1065));
  assign _zz_11626 = ($signed(_zz_1065) + $signed(_zz_1066));
  assign _zz_11627 = _zz_11628[15 : 0];
  assign _zz_11628 = fixTo_782_dout;
  assign _zz_11629 = _zz_11630[15 : 0];
  assign _zz_11630 = fixTo_781_dout;
  assign _zz_11631 = _zz_11632;
  assign _zz_11632 = ($signed(_zz_11633) >>> _zz_3096);
  assign _zz_11633 = _zz_11634;
  assign _zz_11634 = ($signed(_zz_1033) - $signed(_zz_3093));
  assign _zz_11635 = _zz_11636;
  assign _zz_11636 = ($signed(_zz_11637) >>> _zz_3096);
  assign _zz_11637 = _zz_11638;
  assign _zz_11638 = ($signed(_zz_1034) - $signed(_zz_3094));
  assign _zz_11639 = _zz_11640;
  assign _zz_11640 = ($signed(_zz_11641) >>> _zz_3097);
  assign _zz_11641 = _zz_11642;
  assign _zz_11642 = ($signed(_zz_1033) + $signed(_zz_3093));
  assign _zz_11643 = _zz_11644;
  assign _zz_11644 = ($signed(_zz_11645) >>> _zz_3097);
  assign _zz_11645 = _zz_11646;
  assign _zz_11646 = ($signed(_zz_1034) + $signed(_zz_3094));
  assign _zz_11647 = ($signed(twiddle_factor_table_20_real) + $signed(twiddle_factor_table_20_imag));
  assign _zz_11648 = fixTo_783_dout;
  assign _zz_11649 = ($signed(_zz_1068) - $signed(_zz_1067));
  assign _zz_11650 = ($signed(_zz_1067) + $signed(_zz_1068));
  assign _zz_11651 = _zz_11652[15 : 0];
  assign _zz_11652 = fixTo_785_dout;
  assign _zz_11653 = _zz_11654[15 : 0];
  assign _zz_11654 = fixTo_784_dout;
  assign _zz_11655 = _zz_11656;
  assign _zz_11656 = ($signed(_zz_11657) >>> _zz_3101);
  assign _zz_11657 = _zz_11658;
  assign _zz_11658 = ($signed(_zz_1035) - $signed(_zz_3098));
  assign _zz_11659 = _zz_11660;
  assign _zz_11660 = ($signed(_zz_11661) >>> _zz_3101);
  assign _zz_11661 = _zz_11662;
  assign _zz_11662 = ($signed(_zz_1036) - $signed(_zz_3099));
  assign _zz_11663 = _zz_11664;
  assign _zz_11664 = ($signed(_zz_11665) >>> _zz_3102);
  assign _zz_11665 = _zz_11666;
  assign _zz_11666 = ($signed(_zz_1035) + $signed(_zz_3098));
  assign _zz_11667 = _zz_11668;
  assign _zz_11668 = ($signed(_zz_11669) >>> _zz_3102);
  assign _zz_11669 = _zz_11670;
  assign _zz_11670 = ($signed(_zz_1036) + $signed(_zz_3099));
  assign _zz_11671 = ($signed(twiddle_factor_table_21_real) + $signed(twiddle_factor_table_21_imag));
  assign _zz_11672 = fixTo_786_dout;
  assign _zz_11673 = ($signed(_zz_1070) - $signed(_zz_1069));
  assign _zz_11674 = ($signed(_zz_1069) + $signed(_zz_1070));
  assign _zz_11675 = _zz_11676[15 : 0];
  assign _zz_11676 = fixTo_788_dout;
  assign _zz_11677 = _zz_11678[15 : 0];
  assign _zz_11678 = fixTo_787_dout;
  assign _zz_11679 = _zz_11680;
  assign _zz_11680 = ($signed(_zz_11681) >>> _zz_3106);
  assign _zz_11681 = _zz_11682;
  assign _zz_11682 = ($signed(_zz_1037) - $signed(_zz_3103));
  assign _zz_11683 = _zz_11684;
  assign _zz_11684 = ($signed(_zz_11685) >>> _zz_3106);
  assign _zz_11685 = _zz_11686;
  assign _zz_11686 = ($signed(_zz_1038) - $signed(_zz_3104));
  assign _zz_11687 = _zz_11688;
  assign _zz_11688 = ($signed(_zz_11689) >>> _zz_3107);
  assign _zz_11689 = _zz_11690;
  assign _zz_11690 = ($signed(_zz_1037) + $signed(_zz_3103));
  assign _zz_11691 = _zz_11692;
  assign _zz_11692 = ($signed(_zz_11693) >>> _zz_3107);
  assign _zz_11693 = _zz_11694;
  assign _zz_11694 = ($signed(_zz_1038) + $signed(_zz_3104));
  assign _zz_11695 = ($signed(twiddle_factor_table_22_real) + $signed(twiddle_factor_table_22_imag));
  assign _zz_11696 = fixTo_789_dout;
  assign _zz_11697 = ($signed(_zz_1072) - $signed(_zz_1071));
  assign _zz_11698 = ($signed(_zz_1071) + $signed(_zz_1072));
  assign _zz_11699 = _zz_11700[15 : 0];
  assign _zz_11700 = fixTo_791_dout;
  assign _zz_11701 = _zz_11702[15 : 0];
  assign _zz_11702 = fixTo_790_dout;
  assign _zz_11703 = _zz_11704;
  assign _zz_11704 = ($signed(_zz_11705) >>> _zz_3111);
  assign _zz_11705 = _zz_11706;
  assign _zz_11706 = ($signed(_zz_1039) - $signed(_zz_3108));
  assign _zz_11707 = _zz_11708;
  assign _zz_11708 = ($signed(_zz_11709) >>> _zz_3111);
  assign _zz_11709 = _zz_11710;
  assign _zz_11710 = ($signed(_zz_1040) - $signed(_zz_3109));
  assign _zz_11711 = _zz_11712;
  assign _zz_11712 = ($signed(_zz_11713) >>> _zz_3112);
  assign _zz_11713 = _zz_11714;
  assign _zz_11714 = ($signed(_zz_1039) + $signed(_zz_3108));
  assign _zz_11715 = _zz_11716;
  assign _zz_11716 = ($signed(_zz_11717) >>> _zz_3112);
  assign _zz_11717 = _zz_11718;
  assign _zz_11718 = ($signed(_zz_1040) + $signed(_zz_3109));
  assign _zz_11719 = ($signed(twiddle_factor_table_23_real) + $signed(twiddle_factor_table_23_imag));
  assign _zz_11720 = fixTo_792_dout;
  assign _zz_11721 = ($signed(_zz_1074) - $signed(_zz_1073));
  assign _zz_11722 = ($signed(_zz_1073) + $signed(_zz_1074));
  assign _zz_11723 = _zz_11724[15 : 0];
  assign _zz_11724 = fixTo_794_dout;
  assign _zz_11725 = _zz_11726[15 : 0];
  assign _zz_11726 = fixTo_793_dout;
  assign _zz_11727 = _zz_11728;
  assign _zz_11728 = ($signed(_zz_11729) >>> _zz_3116);
  assign _zz_11729 = _zz_11730;
  assign _zz_11730 = ($signed(_zz_1041) - $signed(_zz_3113));
  assign _zz_11731 = _zz_11732;
  assign _zz_11732 = ($signed(_zz_11733) >>> _zz_3116);
  assign _zz_11733 = _zz_11734;
  assign _zz_11734 = ($signed(_zz_1042) - $signed(_zz_3114));
  assign _zz_11735 = _zz_11736;
  assign _zz_11736 = ($signed(_zz_11737) >>> _zz_3117);
  assign _zz_11737 = _zz_11738;
  assign _zz_11738 = ($signed(_zz_1041) + $signed(_zz_3113));
  assign _zz_11739 = _zz_11740;
  assign _zz_11740 = ($signed(_zz_11741) >>> _zz_3117);
  assign _zz_11741 = _zz_11742;
  assign _zz_11742 = ($signed(_zz_1042) + $signed(_zz_3114));
  assign _zz_11743 = ($signed(twiddle_factor_table_24_real) + $signed(twiddle_factor_table_24_imag));
  assign _zz_11744 = fixTo_795_dout;
  assign _zz_11745 = ($signed(_zz_1076) - $signed(_zz_1075));
  assign _zz_11746 = ($signed(_zz_1075) + $signed(_zz_1076));
  assign _zz_11747 = _zz_11748[15 : 0];
  assign _zz_11748 = fixTo_797_dout;
  assign _zz_11749 = _zz_11750[15 : 0];
  assign _zz_11750 = fixTo_796_dout;
  assign _zz_11751 = _zz_11752;
  assign _zz_11752 = ($signed(_zz_11753) >>> _zz_3121);
  assign _zz_11753 = _zz_11754;
  assign _zz_11754 = ($signed(_zz_1043) - $signed(_zz_3118));
  assign _zz_11755 = _zz_11756;
  assign _zz_11756 = ($signed(_zz_11757) >>> _zz_3121);
  assign _zz_11757 = _zz_11758;
  assign _zz_11758 = ($signed(_zz_1044) - $signed(_zz_3119));
  assign _zz_11759 = _zz_11760;
  assign _zz_11760 = ($signed(_zz_11761) >>> _zz_3122);
  assign _zz_11761 = _zz_11762;
  assign _zz_11762 = ($signed(_zz_1043) + $signed(_zz_3118));
  assign _zz_11763 = _zz_11764;
  assign _zz_11764 = ($signed(_zz_11765) >>> _zz_3122);
  assign _zz_11765 = _zz_11766;
  assign _zz_11766 = ($signed(_zz_1044) + $signed(_zz_3119));
  assign _zz_11767 = ($signed(twiddle_factor_table_25_real) + $signed(twiddle_factor_table_25_imag));
  assign _zz_11768 = fixTo_798_dout;
  assign _zz_11769 = ($signed(_zz_1078) - $signed(_zz_1077));
  assign _zz_11770 = ($signed(_zz_1077) + $signed(_zz_1078));
  assign _zz_11771 = _zz_11772[15 : 0];
  assign _zz_11772 = fixTo_800_dout;
  assign _zz_11773 = _zz_11774[15 : 0];
  assign _zz_11774 = fixTo_799_dout;
  assign _zz_11775 = _zz_11776;
  assign _zz_11776 = ($signed(_zz_11777) >>> _zz_3126);
  assign _zz_11777 = _zz_11778;
  assign _zz_11778 = ($signed(_zz_1045) - $signed(_zz_3123));
  assign _zz_11779 = _zz_11780;
  assign _zz_11780 = ($signed(_zz_11781) >>> _zz_3126);
  assign _zz_11781 = _zz_11782;
  assign _zz_11782 = ($signed(_zz_1046) - $signed(_zz_3124));
  assign _zz_11783 = _zz_11784;
  assign _zz_11784 = ($signed(_zz_11785) >>> _zz_3127);
  assign _zz_11785 = _zz_11786;
  assign _zz_11786 = ($signed(_zz_1045) + $signed(_zz_3123));
  assign _zz_11787 = _zz_11788;
  assign _zz_11788 = ($signed(_zz_11789) >>> _zz_3127);
  assign _zz_11789 = _zz_11790;
  assign _zz_11790 = ($signed(_zz_1046) + $signed(_zz_3124));
  assign _zz_11791 = ($signed(twiddle_factor_table_26_real) + $signed(twiddle_factor_table_26_imag));
  assign _zz_11792 = fixTo_801_dout;
  assign _zz_11793 = ($signed(_zz_1080) - $signed(_zz_1079));
  assign _zz_11794 = ($signed(_zz_1079) + $signed(_zz_1080));
  assign _zz_11795 = _zz_11796[15 : 0];
  assign _zz_11796 = fixTo_803_dout;
  assign _zz_11797 = _zz_11798[15 : 0];
  assign _zz_11798 = fixTo_802_dout;
  assign _zz_11799 = _zz_11800;
  assign _zz_11800 = ($signed(_zz_11801) >>> _zz_3131);
  assign _zz_11801 = _zz_11802;
  assign _zz_11802 = ($signed(_zz_1047) - $signed(_zz_3128));
  assign _zz_11803 = _zz_11804;
  assign _zz_11804 = ($signed(_zz_11805) >>> _zz_3131);
  assign _zz_11805 = _zz_11806;
  assign _zz_11806 = ($signed(_zz_1048) - $signed(_zz_3129));
  assign _zz_11807 = _zz_11808;
  assign _zz_11808 = ($signed(_zz_11809) >>> _zz_3132);
  assign _zz_11809 = _zz_11810;
  assign _zz_11810 = ($signed(_zz_1047) + $signed(_zz_3128));
  assign _zz_11811 = _zz_11812;
  assign _zz_11812 = ($signed(_zz_11813) >>> _zz_3132);
  assign _zz_11813 = _zz_11814;
  assign _zz_11814 = ($signed(_zz_1048) + $signed(_zz_3129));
  assign _zz_11815 = ($signed(twiddle_factor_table_27_real) + $signed(twiddle_factor_table_27_imag));
  assign _zz_11816 = fixTo_804_dout;
  assign _zz_11817 = ($signed(_zz_1082) - $signed(_zz_1081));
  assign _zz_11818 = ($signed(_zz_1081) + $signed(_zz_1082));
  assign _zz_11819 = _zz_11820[15 : 0];
  assign _zz_11820 = fixTo_806_dout;
  assign _zz_11821 = _zz_11822[15 : 0];
  assign _zz_11822 = fixTo_805_dout;
  assign _zz_11823 = _zz_11824;
  assign _zz_11824 = ($signed(_zz_11825) >>> _zz_3136);
  assign _zz_11825 = _zz_11826;
  assign _zz_11826 = ($signed(_zz_1049) - $signed(_zz_3133));
  assign _zz_11827 = _zz_11828;
  assign _zz_11828 = ($signed(_zz_11829) >>> _zz_3136);
  assign _zz_11829 = _zz_11830;
  assign _zz_11830 = ($signed(_zz_1050) - $signed(_zz_3134));
  assign _zz_11831 = _zz_11832;
  assign _zz_11832 = ($signed(_zz_11833) >>> _zz_3137);
  assign _zz_11833 = _zz_11834;
  assign _zz_11834 = ($signed(_zz_1049) + $signed(_zz_3133));
  assign _zz_11835 = _zz_11836;
  assign _zz_11836 = ($signed(_zz_11837) >>> _zz_3137);
  assign _zz_11837 = _zz_11838;
  assign _zz_11838 = ($signed(_zz_1050) + $signed(_zz_3134));
  assign _zz_11839 = ($signed(twiddle_factor_table_28_real) + $signed(twiddle_factor_table_28_imag));
  assign _zz_11840 = fixTo_807_dout;
  assign _zz_11841 = ($signed(_zz_1084) - $signed(_zz_1083));
  assign _zz_11842 = ($signed(_zz_1083) + $signed(_zz_1084));
  assign _zz_11843 = _zz_11844[15 : 0];
  assign _zz_11844 = fixTo_809_dout;
  assign _zz_11845 = _zz_11846[15 : 0];
  assign _zz_11846 = fixTo_808_dout;
  assign _zz_11847 = _zz_11848;
  assign _zz_11848 = ($signed(_zz_11849) >>> _zz_3141);
  assign _zz_11849 = _zz_11850;
  assign _zz_11850 = ($signed(_zz_1051) - $signed(_zz_3138));
  assign _zz_11851 = _zz_11852;
  assign _zz_11852 = ($signed(_zz_11853) >>> _zz_3141);
  assign _zz_11853 = _zz_11854;
  assign _zz_11854 = ($signed(_zz_1052) - $signed(_zz_3139));
  assign _zz_11855 = _zz_11856;
  assign _zz_11856 = ($signed(_zz_11857) >>> _zz_3142);
  assign _zz_11857 = _zz_11858;
  assign _zz_11858 = ($signed(_zz_1051) + $signed(_zz_3138));
  assign _zz_11859 = _zz_11860;
  assign _zz_11860 = ($signed(_zz_11861) >>> _zz_3142);
  assign _zz_11861 = _zz_11862;
  assign _zz_11862 = ($signed(_zz_1052) + $signed(_zz_3139));
  assign _zz_11863 = ($signed(twiddle_factor_table_29_real) + $signed(twiddle_factor_table_29_imag));
  assign _zz_11864 = fixTo_810_dout;
  assign _zz_11865 = ($signed(_zz_1086) - $signed(_zz_1085));
  assign _zz_11866 = ($signed(_zz_1085) + $signed(_zz_1086));
  assign _zz_11867 = _zz_11868[15 : 0];
  assign _zz_11868 = fixTo_812_dout;
  assign _zz_11869 = _zz_11870[15 : 0];
  assign _zz_11870 = fixTo_811_dout;
  assign _zz_11871 = _zz_11872;
  assign _zz_11872 = ($signed(_zz_11873) >>> _zz_3146);
  assign _zz_11873 = _zz_11874;
  assign _zz_11874 = ($signed(_zz_1053) - $signed(_zz_3143));
  assign _zz_11875 = _zz_11876;
  assign _zz_11876 = ($signed(_zz_11877) >>> _zz_3146);
  assign _zz_11877 = _zz_11878;
  assign _zz_11878 = ($signed(_zz_1054) - $signed(_zz_3144));
  assign _zz_11879 = _zz_11880;
  assign _zz_11880 = ($signed(_zz_11881) >>> _zz_3147);
  assign _zz_11881 = _zz_11882;
  assign _zz_11882 = ($signed(_zz_1053) + $signed(_zz_3143));
  assign _zz_11883 = _zz_11884;
  assign _zz_11884 = ($signed(_zz_11885) >>> _zz_3147);
  assign _zz_11885 = _zz_11886;
  assign _zz_11886 = ($signed(_zz_1054) + $signed(_zz_3144));
  assign _zz_11887 = ($signed(twiddle_factor_table_30_real) + $signed(twiddle_factor_table_30_imag));
  assign _zz_11888 = fixTo_813_dout;
  assign _zz_11889 = ($signed(_zz_1088) - $signed(_zz_1087));
  assign _zz_11890 = ($signed(_zz_1087) + $signed(_zz_1088));
  assign _zz_11891 = _zz_11892[15 : 0];
  assign _zz_11892 = fixTo_815_dout;
  assign _zz_11893 = _zz_11894[15 : 0];
  assign _zz_11894 = fixTo_814_dout;
  assign _zz_11895 = _zz_11896;
  assign _zz_11896 = ($signed(_zz_11897) >>> _zz_3151);
  assign _zz_11897 = _zz_11898;
  assign _zz_11898 = ($signed(_zz_1055) - $signed(_zz_3148));
  assign _zz_11899 = _zz_11900;
  assign _zz_11900 = ($signed(_zz_11901) >>> _zz_3151);
  assign _zz_11901 = _zz_11902;
  assign _zz_11902 = ($signed(_zz_1056) - $signed(_zz_3149));
  assign _zz_11903 = _zz_11904;
  assign _zz_11904 = ($signed(_zz_11905) >>> _zz_3152);
  assign _zz_11905 = _zz_11906;
  assign _zz_11906 = ($signed(_zz_1055) + $signed(_zz_3148));
  assign _zz_11907 = _zz_11908;
  assign _zz_11908 = ($signed(_zz_11909) >>> _zz_3152);
  assign _zz_11909 = _zz_11910;
  assign _zz_11910 = ($signed(_zz_1056) + $signed(_zz_3149));
  assign _zz_11911 = ($signed(twiddle_factor_table_15_real) + $signed(twiddle_factor_table_15_imag));
  assign _zz_11912 = fixTo_816_dout;
  assign _zz_11913 = ($signed(_zz_1122) - $signed(_zz_1121));
  assign _zz_11914 = ($signed(_zz_1121) + $signed(_zz_1122));
  assign _zz_11915 = _zz_11916[15 : 0];
  assign _zz_11916 = fixTo_818_dout;
  assign _zz_11917 = _zz_11918[15 : 0];
  assign _zz_11918 = fixTo_817_dout;
  assign _zz_11919 = _zz_11920;
  assign _zz_11920 = ($signed(_zz_11921) >>> _zz_3156);
  assign _zz_11921 = _zz_11922;
  assign _zz_11922 = ($signed(_zz_1089) - $signed(_zz_3153));
  assign _zz_11923 = _zz_11924;
  assign _zz_11924 = ($signed(_zz_11925) >>> _zz_3156);
  assign _zz_11925 = _zz_11926;
  assign _zz_11926 = ($signed(_zz_1090) - $signed(_zz_3154));
  assign _zz_11927 = _zz_11928;
  assign _zz_11928 = ($signed(_zz_11929) >>> _zz_3157);
  assign _zz_11929 = _zz_11930;
  assign _zz_11930 = ($signed(_zz_1089) + $signed(_zz_3153));
  assign _zz_11931 = _zz_11932;
  assign _zz_11932 = ($signed(_zz_11933) >>> _zz_3157);
  assign _zz_11933 = _zz_11934;
  assign _zz_11934 = ($signed(_zz_1090) + $signed(_zz_3154));
  assign _zz_11935 = ($signed(twiddle_factor_table_16_real) + $signed(twiddle_factor_table_16_imag));
  assign _zz_11936 = fixTo_819_dout;
  assign _zz_11937 = ($signed(_zz_1124) - $signed(_zz_1123));
  assign _zz_11938 = ($signed(_zz_1123) + $signed(_zz_1124));
  assign _zz_11939 = _zz_11940[15 : 0];
  assign _zz_11940 = fixTo_821_dout;
  assign _zz_11941 = _zz_11942[15 : 0];
  assign _zz_11942 = fixTo_820_dout;
  assign _zz_11943 = _zz_11944;
  assign _zz_11944 = ($signed(_zz_11945) >>> _zz_3161);
  assign _zz_11945 = _zz_11946;
  assign _zz_11946 = ($signed(_zz_1091) - $signed(_zz_3158));
  assign _zz_11947 = _zz_11948;
  assign _zz_11948 = ($signed(_zz_11949) >>> _zz_3161);
  assign _zz_11949 = _zz_11950;
  assign _zz_11950 = ($signed(_zz_1092) - $signed(_zz_3159));
  assign _zz_11951 = _zz_11952;
  assign _zz_11952 = ($signed(_zz_11953) >>> _zz_3162);
  assign _zz_11953 = _zz_11954;
  assign _zz_11954 = ($signed(_zz_1091) + $signed(_zz_3158));
  assign _zz_11955 = _zz_11956;
  assign _zz_11956 = ($signed(_zz_11957) >>> _zz_3162);
  assign _zz_11957 = _zz_11958;
  assign _zz_11958 = ($signed(_zz_1092) + $signed(_zz_3159));
  assign _zz_11959 = ($signed(twiddle_factor_table_17_real) + $signed(twiddle_factor_table_17_imag));
  assign _zz_11960 = fixTo_822_dout;
  assign _zz_11961 = ($signed(_zz_1126) - $signed(_zz_1125));
  assign _zz_11962 = ($signed(_zz_1125) + $signed(_zz_1126));
  assign _zz_11963 = _zz_11964[15 : 0];
  assign _zz_11964 = fixTo_824_dout;
  assign _zz_11965 = _zz_11966[15 : 0];
  assign _zz_11966 = fixTo_823_dout;
  assign _zz_11967 = _zz_11968;
  assign _zz_11968 = ($signed(_zz_11969) >>> _zz_3166);
  assign _zz_11969 = _zz_11970;
  assign _zz_11970 = ($signed(_zz_1093) - $signed(_zz_3163));
  assign _zz_11971 = _zz_11972;
  assign _zz_11972 = ($signed(_zz_11973) >>> _zz_3166);
  assign _zz_11973 = _zz_11974;
  assign _zz_11974 = ($signed(_zz_1094) - $signed(_zz_3164));
  assign _zz_11975 = _zz_11976;
  assign _zz_11976 = ($signed(_zz_11977) >>> _zz_3167);
  assign _zz_11977 = _zz_11978;
  assign _zz_11978 = ($signed(_zz_1093) + $signed(_zz_3163));
  assign _zz_11979 = _zz_11980;
  assign _zz_11980 = ($signed(_zz_11981) >>> _zz_3167);
  assign _zz_11981 = _zz_11982;
  assign _zz_11982 = ($signed(_zz_1094) + $signed(_zz_3164));
  assign _zz_11983 = ($signed(twiddle_factor_table_18_real) + $signed(twiddle_factor_table_18_imag));
  assign _zz_11984 = fixTo_825_dout;
  assign _zz_11985 = ($signed(_zz_1128) - $signed(_zz_1127));
  assign _zz_11986 = ($signed(_zz_1127) + $signed(_zz_1128));
  assign _zz_11987 = _zz_11988[15 : 0];
  assign _zz_11988 = fixTo_827_dout;
  assign _zz_11989 = _zz_11990[15 : 0];
  assign _zz_11990 = fixTo_826_dout;
  assign _zz_11991 = _zz_11992;
  assign _zz_11992 = ($signed(_zz_11993) >>> _zz_3171);
  assign _zz_11993 = _zz_11994;
  assign _zz_11994 = ($signed(_zz_1095) - $signed(_zz_3168));
  assign _zz_11995 = _zz_11996;
  assign _zz_11996 = ($signed(_zz_11997) >>> _zz_3171);
  assign _zz_11997 = _zz_11998;
  assign _zz_11998 = ($signed(_zz_1096) - $signed(_zz_3169));
  assign _zz_11999 = _zz_12000;
  assign _zz_12000 = ($signed(_zz_12001) >>> _zz_3172);
  assign _zz_12001 = _zz_12002;
  assign _zz_12002 = ($signed(_zz_1095) + $signed(_zz_3168));
  assign _zz_12003 = _zz_12004;
  assign _zz_12004 = ($signed(_zz_12005) >>> _zz_3172);
  assign _zz_12005 = _zz_12006;
  assign _zz_12006 = ($signed(_zz_1096) + $signed(_zz_3169));
  assign _zz_12007 = ($signed(twiddle_factor_table_19_real) + $signed(twiddle_factor_table_19_imag));
  assign _zz_12008 = fixTo_828_dout;
  assign _zz_12009 = ($signed(_zz_1130) - $signed(_zz_1129));
  assign _zz_12010 = ($signed(_zz_1129) + $signed(_zz_1130));
  assign _zz_12011 = _zz_12012[15 : 0];
  assign _zz_12012 = fixTo_830_dout;
  assign _zz_12013 = _zz_12014[15 : 0];
  assign _zz_12014 = fixTo_829_dout;
  assign _zz_12015 = _zz_12016;
  assign _zz_12016 = ($signed(_zz_12017) >>> _zz_3176);
  assign _zz_12017 = _zz_12018;
  assign _zz_12018 = ($signed(_zz_1097) - $signed(_zz_3173));
  assign _zz_12019 = _zz_12020;
  assign _zz_12020 = ($signed(_zz_12021) >>> _zz_3176);
  assign _zz_12021 = _zz_12022;
  assign _zz_12022 = ($signed(_zz_1098) - $signed(_zz_3174));
  assign _zz_12023 = _zz_12024;
  assign _zz_12024 = ($signed(_zz_12025) >>> _zz_3177);
  assign _zz_12025 = _zz_12026;
  assign _zz_12026 = ($signed(_zz_1097) + $signed(_zz_3173));
  assign _zz_12027 = _zz_12028;
  assign _zz_12028 = ($signed(_zz_12029) >>> _zz_3177);
  assign _zz_12029 = _zz_12030;
  assign _zz_12030 = ($signed(_zz_1098) + $signed(_zz_3174));
  assign _zz_12031 = ($signed(twiddle_factor_table_20_real) + $signed(twiddle_factor_table_20_imag));
  assign _zz_12032 = fixTo_831_dout;
  assign _zz_12033 = ($signed(_zz_1132) - $signed(_zz_1131));
  assign _zz_12034 = ($signed(_zz_1131) + $signed(_zz_1132));
  assign _zz_12035 = _zz_12036[15 : 0];
  assign _zz_12036 = fixTo_833_dout;
  assign _zz_12037 = _zz_12038[15 : 0];
  assign _zz_12038 = fixTo_832_dout;
  assign _zz_12039 = _zz_12040;
  assign _zz_12040 = ($signed(_zz_12041) >>> _zz_3181);
  assign _zz_12041 = _zz_12042;
  assign _zz_12042 = ($signed(_zz_1099) - $signed(_zz_3178));
  assign _zz_12043 = _zz_12044;
  assign _zz_12044 = ($signed(_zz_12045) >>> _zz_3181);
  assign _zz_12045 = _zz_12046;
  assign _zz_12046 = ($signed(_zz_1100) - $signed(_zz_3179));
  assign _zz_12047 = _zz_12048;
  assign _zz_12048 = ($signed(_zz_12049) >>> _zz_3182);
  assign _zz_12049 = _zz_12050;
  assign _zz_12050 = ($signed(_zz_1099) + $signed(_zz_3178));
  assign _zz_12051 = _zz_12052;
  assign _zz_12052 = ($signed(_zz_12053) >>> _zz_3182);
  assign _zz_12053 = _zz_12054;
  assign _zz_12054 = ($signed(_zz_1100) + $signed(_zz_3179));
  assign _zz_12055 = ($signed(twiddle_factor_table_21_real) + $signed(twiddle_factor_table_21_imag));
  assign _zz_12056 = fixTo_834_dout;
  assign _zz_12057 = ($signed(_zz_1134) - $signed(_zz_1133));
  assign _zz_12058 = ($signed(_zz_1133) + $signed(_zz_1134));
  assign _zz_12059 = _zz_12060[15 : 0];
  assign _zz_12060 = fixTo_836_dout;
  assign _zz_12061 = _zz_12062[15 : 0];
  assign _zz_12062 = fixTo_835_dout;
  assign _zz_12063 = _zz_12064;
  assign _zz_12064 = ($signed(_zz_12065) >>> _zz_3186);
  assign _zz_12065 = _zz_12066;
  assign _zz_12066 = ($signed(_zz_1101) - $signed(_zz_3183));
  assign _zz_12067 = _zz_12068;
  assign _zz_12068 = ($signed(_zz_12069) >>> _zz_3186);
  assign _zz_12069 = _zz_12070;
  assign _zz_12070 = ($signed(_zz_1102) - $signed(_zz_3184));
  assign _zz_12071 = _zz_12072;
  assign _zz_12072 = ($signed(_zz_12073) >>> _zz_3187);
  assign _zz_12073 = _zz_12074;
  assign _zz_12074 = ($signed(_zz_1101) + $signed(_zz_3183));
  assign _zz_12075 = _zz_12076;
  assign _zz_12076 = ($signed(_zz_12077) >>> _zz_3187);
  assign _zz_12077 = _zz_12078;
  assign _zz_12078 = ($signed(_zz_1102) + $signed(_zz_3184));
  assign _zz_12079 = ($signed(twiddle_factor_table_22_real) + $signed(twiddle_factor_table_22_imag));
  assign _zz_12080 = fixTo_837_dout;
  assign _zz_12081 = ($signed(_zz_1136) - $signed(_zz_1135));
  assign _zz_12082 = ($signed(_zz_1135) + $signed(_zz_1136));
  assign _zz_12083 = _zz_12084[15 : 0];
  assign _zz_12084 = fixTo_839_dout;
  assign _zz_12085 = _zz_12086[15 : 0];
  assign _zz_12086 = fixTo_838_dout;
  assign _zz_12087 = _zz_12088;
  assign _zz_12088 = ($signed(_zz_12089) >>> _zz_3191);
  assign _zz_12089 = _zz_12090;
  assign _zz_12090 = ($signed(_zz_1103) - $signed(_zz_3188));
  assign _zz_12091 = _zz_12092;
  assign _zz_12092 = ($signed(_zz_12093) >>> _zz_3191);
  assign _zz_12093 = _zz_12094;
  assign _zz_12094 = ($signed(_zz_1104) - $signed(_zz_3189));
  assign _zz_12095 = _zz_12096;
  assign _zz_12096 = ($signed(_zz_12097) >>> _zz_3192);
  assign _zz_12097 = _zz_12098;
  assign _zz_12098 = ($signed(_zz_1103) + $signed(_zz_3188));
  assign _zz_12099 = _zz_12100;
  assign _zz_12100 = ($signed(_zz_12101) >>> _zz_3192);
  assign _zz_12101 = _zz_12102;
  assign _zz_12102 = ($signed(_zz_1104) + $signed(_zz_3189));
  assign _zz_12103 = ($signed(twiddle_factor_table_23_real) + $signed(twiddle_factor_table_23_imag));
  assign _zz_12104 = fixTo_840_dout;
  assign _zz_12105 = ($signed(_zz_1138) - $signed(_zz_1137));
  assign _zz_12106 = ($signed(_zz_1137) + $signed(_zz_1138));
  assign _zz_12107 = _zz_12108[15 : 0];
  assign _zz_12108 = fixTo_842_dout;
  assign _zz_12109 = _zz_12110[15 : 0];
  assign _zz_12110 = fixTo_841_dout;
  assign _zz_12111 = _zz_12112;
  assign _zz_12112 = ($signed(_zz_12113) >>> _zz_3196);
  assign _zz_12113 = _zz_12114;
  assign _zz_12114 = ($signed(_zz_1105) - $signed(_zz_3193));
  assign _zz_12115 = _zz_12116;
  assign _zz_12116 = ($signed(_zz_12117) >>> _zz_3196);
  assign _zz_12117 = _zz_12118;
  assign _zz_12118 = ($signed(_zz_1106) - $signed(_zz_3194));
  assign _zz_12119 = _zz_12120;
  assign _zz_12120 = ($signed(_zz_12121) >>> _zz_3197);
  assign _zz_12121 = _zz_12122;
  assign _zz_12122 = ($signed(_zz_1105) + $signed(_zz_3193));
  assign _zz_12123 = _zz_12124;
  assign _zz_12124 = ($signed(_zz_12125) >>> _zz_3197);
  assign _zz_12125 = _zz_12126;
  assign _zz_12126 = ($signed(_zz_1106) + $signed(_zz_3194));
  assign _zz_12127 = ($signed(twiddle_factor_table_24_real) + $signed(twiddle_factor_table_24_imag));
  assign _zz_12128 = fixTo_843_dout;
  assign _zz_12129 = ($signed(_zz_1140) - $signed(_zz_1139));
  assign _zz_12130 = ($signed(_zz_1139) + $signed(_zz_1140));
  assign _zz_12131 = _zz_12132[15 : 0];
  assign _zz_12132 = fixTo_845_dout;
  assign _zz_12133 = _zz_12134[15 : 0];
  assign _zz_12134 = fixTo_844_dout;
  assign _zz_12135 = _zz_12136;
  assign _zz_12136 = ($signed(_zz_12137) >>> _zz_3201);
  assign _zz_12137 = _zz_12138;
  assign _zz_12138 = ($signed(_zz_1107) - $signed(_zz_3198));
  assign _zz_12139 = _zz_12140;
  assign _zz_12140 = ($signed(_zz_12141) >>> _zz_3201);
  assign _zz_12141 = _zz_12142;
  assign _zz_12142 = ($signed(_zz_1108) - $signed(_zz_3199));
  assign _zz_12143 = _zz_12144;
  assign _zz_12144 = ($signed(_zz_12145) >>> _zz_3202);
  assign _zz_12145 = _zz_12146;
  assign _zz_12146 = ($signed(_zz_1107) + $signed(_zz_3198));
  assign _zz_12147 = _zz_12148;
  assign _zz_12148 = ($signed(_zz_12149) >>> _zz_3202);
  assign _zz_12149 = _zz_12150;
  assign _zz_12150 = ($signed(_zz_1108) + $signed(_zz_3199));
  assign _zz_12151 = ($signed(twiddle_factor_table_25_real) + $signed(twiddle_factor_table_25_imag));
  assign _zz_12152 = fixTo_846_dout;
  assign _zz_12153 = ($signed(_zz_1142) - $signed(_zz_1141));
  assign _zz_12154 = ($signed(_zz_1141) + $signed(_zz_1142));
  assign _zz_12155 = _zz_12156[15 : 0];
  assign _zz_12156 = fixTo_848_dout;
  assign _zz_12157 = _zz_12158[15 : 0];
  assign _zz_12158 = fixTo_847_dout;
  assign _zz_12159 = _zz_12160;
  assign _zz_12160 = ($signed(_zz_12161) >>> _zz_3206);
  assign _zz_12161 = _zz_12162;
  assign _zz_12162 = ($signed(_zz_1109) - $signed(_zz_3203));
  assign _zz_12163 = _zz_12164;
  assign _zz_12164 = ($signed(_zz_12165) >>> _zz_3206);
  assign _zz_12165 = _zz_12166;
  assign _zz_12166 = ($signed(_zz_1110) - $signed(_zz_3204));
  assign _zz_12167 = _zz_12168;
  assign _zz_12168 = ($signed(_zz_12169) >>> _zz_3207);
  assign _zz_12169 = _zz_12170;
  assign _zz_12170 = ($signed(_zz_1109) + $signed(_zz_3203));
  assign _zz_12171 = _zz_12172;
  assign _zz_12172 = ($signed(_zz_12173) >>> _zz_3207);
  assign _zz_12173 = _zz_12174;
  assign _zz_12174 = ($signed(_zz_1110) + $signed(_zz_3204));
  assign _zz_12175 = ($signed(twiddle_factor_table_26_real) + $signed(twiddle_factor_table_26_imag));
  assign _zz_12176 = fixTo_849_dout;
  assign _zz_12177 = ($signed(_zz_1144) - $signed(_zz_1143));
  assign _zz_12178 = ($signed(_zz_1143) + $signed(_zz_1144));
  assign _zz_12179 = _zz_12180[15 : 0];
  assign _zz_12180 = fixTo_851_dout;
  assign _zz_12181 = _zz_12182[15 : 0];
  assign _zz_12182 = fixTo_850_dout;
  assign _zz_12183 = _zz_12184;
  assign _zz_12184 = ($signed(_zz_12185) >>> _zz_3211);
  assign _zz_12185 = _zz_12186;
  assign _zz_12186 = ($signed(_zz_1111) - $signed(_zz_3208));
  assign _zz_12187 = _zz_12188;
  assign _zz_12188 = ($signed(_zz_12189) >>> _zz_3211);
  assign _zz_12189 = _zz_12190;
  assign _zz_12190 = ($signed(_zz_1112) - $signed(_zz_3209));
  assign _zz_12191 = _zz_12192;
  assign _zz_12192 = ($signed(_zz_12193) >>> _zz_3212);
  assign _zz_12193 = _zz_12194;
  assign _zz_12194 = ($signed(_zz_1111) + $signed(_zz_3208));
  assign _zz_12195 = _zz_12196;
  assign _zz_12196 = ($signed(_zz_12197) >>> _zz_3212);
  assign _zz_12197 = _zz_12198;
  assign _zz_12198 = ($signed(_zz_1112) + $signed(_zz_3209));
  assign _zz_12199 = ($signed(twiddle_factor_table_27_real) + $signed(twiddle_factor_table_27_imag));
  assign _zz_12200 = fixTo_852_dout;
  assign _zz_12201 = ($signed(_zz_1146) - $signed(_zz_1145));
  assign _zz_12202 = ($signed(_zz_1145) + $signed(_zz_1146));
  assign _zz_12203 = _zz_12204[15 : 0];
  assign _zz_12204 = fixTo_854_dout;
  assign _zz_12205 = _zz_12206[15 : 0];
  assign _zz_12206 = fixTo_853_dout;
  assign _zz_12207 = _zz_12208;
  assign _zz_12208 = ($signed(_zz_12209) >>> _zz_3216);
  assign _zz_12209 = _zz_12210;
  assign _zz_12210 = ($signed(_zz_1113) - $signed(_zz_3213));
  assign _zz_12211 = _zz_12212;
  assign _zz_12212 = ($signed(_zz_12213) >>> _zz_3216);
  assign _zz_12213 = _zz_12214;
  assign _zz_12214 = ($signed(_zz_1114) - $signed(_zz_3214));
  assign _zz_12215 = _zz_12216;
  assign _zz_12216 = ($signed(_zz_12217) >>> _zz_3217);
  assign _zz_12217 = _zz_12218;
  assign _zz_12218 = ($signed(_zz_1113) + $signed(_zz_3213));
  assign _zz_12219 = _zz_12220;
  assign _zz_12220 = ($signed(_zz_12221) >>> _zz_3217);
  assign _zz_12221 = _zz_12222;
  assign _zz_12222 = ($signed(_zz_1114) + $signed(_zz_3214));
  assign _zz_12223 = ($signed(twiddle_factor_table_28_real) + $signed(twiddle_factor_table_28_imag));
  assign _zz_12224 = fixTo_855_dout;
  assign _zz_12225 = ($signed(_zz_1148) - $signed(_zz_1147));
  assign _zz_12226 = ($signed(_zz_1147) + $signed(_zz_1148));
  assign _zz_12227 = _zz_12228[15 : 0];
  assign _zz_12228 = fixTo_857_dout;
  assign _zz_12229 = _zz_12230[15 : 0];
  assign _zz_12230 = fixTo_856_dout;
  assign _zz_12231 = _zz_12232;
  assign _zz_12232 = ($signed(_zz_12233) >>> _zz_3221);
  assign _zz_12233 = _zz_12234;
  assign _zz_12234 = ($signed(_zz_1115) - $signed(_zz_3218));
  assign _zz_12235 = _zz_12236;
  assign _zz_12236 = ($signed(_zz_12237) >>> _zz_3221);
  assign _zz_12237 = _zz_12238;
  assign _zz_12238 = ($signed(_zz_1116) - $signed(_zz_3219));
  assign _zz_12239 = _zz_12240;
  assign _zz_12240 = ($signed(_zz_12241) >>> _zz_3222);
  assign _zz_12241 = _zz_12242;
  assign _zz_12242 = ($signed(_zz_1115) + $signed(_zz_3218));
  assign _zz_12243 = _zz_12244;
  assign _zz_12244 = ($signed(_zz_12245) >>> _zz_3222);
  assign _zz_12245 = _zz_12246;
  assign _zz_12246 = ($signed(_zz_1116) + $signed(_zz_3219));
  assign _zz_12247 = ($signed(twiddle_factor_table_29_real) + $signed(twiddle_factor_table_29_imag));
  assign _zz_12248 = fixTo_858_dout;
  assign _zz_12249 = ($signed(_zz_1150) - $signed(_zz_1149));
  assign _zz_12250 = ($signed(_zz_1149) + $signed(_zz_1150));
  assign _zz_12251 = _zz_12252[15 : 0];
  assign _zz_12252 = fixTo_860_dout;
  assign _zz_12253 = _zz_12254[15 : 0];
  assign _zz_12254 = fixTo_859_dout;
  assign _zz_12255 = _zz_12256;
  assign _zz_12256 = ($signed(_zz_12257) >>> _zz_3226);
  assign _zz_12257 = _zz_12258;
  assign _zz_12258 = ($signed(_zz_1117) - $signed(_zz_3223));
  assign _zz_12259 = _zz_12260;
  assign _zz_12260 = ($signed(_zz_12261) >>> _zz_3226);
  assign _zz_12261 = _zz_12262;
  assign _zz_12262 = ($signed(_zz_1118) - $signed(_zz_3224));
  assign _zz_12263 = _zz_12264;
  assign _zz_12264 = ($signed(_zz_12265) >>> _zz_3227);
  assign _zz_12265 = _zz_12266;
  assign _zz_12266 = ($signed(_zz_1117) + $signed(_zz_3223));
  assign _zz_12267 = _zz_12268;
  assign _zz_12268 = ($signed(_zz_12269) >>> _zz_3227);
  assign _zz_12269 = _zz_12270;
  assign _zz_12270 = ($signed(_zz_1118) + $signed(_zz_3224));
  assign _zz_12271 = ($signed(twiddle_factor_table_30_real) + $signed(twiddle_factor_table_30_imag));
  assign _zz_12272 = fixTo_861_dout;
  assign _zz_12273 = ($signed(_zz_1152) - $signed(_zz_1151));
  assign _zz_12274 = ($signed(_zz_1151) + $signed(_zz_1152));
  assign _zz_12275 = _zz_12276[15 : 0];
  assign _zz_12276 = fixTo_863_dout;
  assign _zz_12277 = _zz_12278[15 : 0];
  assign _zz_12278 = fixTo_862_dout;
  assign _zz_12279 = _zz_12280;
  assign _zz_12280 = ($signed(_zz_12281) >>> _zz_3231);
  assign _zz_12281 = _zz_12282;
  assign _zz_12282 = ($signed(_zz_1119) - $signed(_zz_3228));
  assign _zz_12283 = _zz_12284;
  assign _zz_12284 = ($signed(_zz_12285) >>> _zz_3231);
  assign _zz_12285 = _zz_12286;
  assign _zz_12286 = ($signed(_zz_1120) - $signed(_zz_3229));
  assign _zz_12287 = _zz_12288;
  assign _zz_12288 = ($signed(_zz_12289) >>> _zz_3232);
  assign _zz_12289 = _zz_12290;
  assign _zz_12290 = ($signed(_zz_1119) + $signed(_zz_3228));
  assign _zz_12291 = _zz_12292;
  assign _zz_12292 = ($signed(_zz_12293) >>> _zz_3232);
  assign _zz_12293 = _zz_12294;
  assign _zz_12294 = ($signed(_zz_1120) + $signed(_zz_3229));
  assign _zz_12295 = ($signed(twiddle_factor_table_15_real) + $signed(twiddle_factor_table_15_imag));
  assign _zz_12296 = fixTo_864_dout;
  assign _zz_12297 = ($signed(_zz_1186) - $signed(_zz_1185));
  assign _zz_12298 = ($signed(_zz_1185) + $signed(_zz_1186));
  assign _zz_12299 = _zz_12300[15 : 0];
  assign _zz_12300 = fixTo_866_dout;
  assign _zz_12301 = _zz_12302[15 : 0];
  assign _zz_12302 = fixTo_865_dout;
  assign _zz_12303 = _zz_12304;
  assign _zz_12304 = ($signed(_zz_12305) >>> _zz_3236);
  assign _zz_12305 = _zz_12306;
  assign _zz_12306 = ($signed(_zz_1153) - $signed(_zz_3233));
  assign _zz_12307 = _zz_12308;
  assign _zz_12308 = ($signed(_zz_12309) >>> _zz_3236);
  assign _zz_12309 = _zz_12310;
  assign _zz_12310 = ($signed(_zz_1154) - $signed(_zz_3234));
  assign _zz_12311 = _zz_12312;
  assign _zz_12312 = ($signed(_zz_12313) >>> _zz_3237);
  assign _zz_12313 = _zz_12314;
  assign _zz_12314 = ($signed(_zz_1153) + $signed(_zz_3233));
  assign _zz_12315 = _zz_12316;
  assign _zz_12316 = ($signed(_zz_12317) >>> _zz_3237);
  assign _zz_12317 = _zz_12318;
  assign _zz_12318 = ($signed(_zz_1154) + $signed(_zz_3234));
  assign _zz_12319 = ($signed(twiddle_factor_table_16_real) + $signed(twiddle_factor_table_16_imag));
  assign _zz_12320 = fixTo_867_dout;
  assign _zz_12321 = ($signed(_zz_1188) - $signed(_zz_1187));
  assign _zz_12322 = ($signed(_zz_1187) + $signed(_zz_1188));
  assign _zz_12323 = _zz_12324[15 : 0];
  assign _zz_12324 = fixTo_869_dout;
  assign _zz_12325 = _zz_12326[15 : 0];
  assign _zz_12326 = fixTo_868_dout;
  assign _zz_12327 = _zz_12328;
  assign _zz_12328 = ($signed(_zz_12329) >>> _zz_3241);
  assign _zz_12329 = _zz_12330;
  assign _zz_12330 = ($signed(_zz_1155) - $signed(_zz_3238));
  assign _zz_12331 = _zz_12332;
  assign _zz_12332 = ($signed(_zz_12333) >>> _zz_3241);
  assign _zz_12333 = _zz_12334;
  assign _zz_12334 = ($signed(_zz_1156) - $signed(_zz_3239));
  assign _zz_12335 = _zz_12336;
  assign _zz_12336 = ($signed(_zz_12337) >>> _zz_3242);
  assign _zz_12337 = _zz_12338;
  assign _zz_12338 = ($signed(_zz_1155) + $signed(_zz_3238));
  assign _zz_12339 = _zz_12340;
  assign _zz_12340 = ($signed(_zz_12341) >>> _zz_3242);
  assign _zz_12341 = _zz_12342;
  assign _zz_12342 = ($signed(_zz_1156) + $signed(_zz_3239));
  assign _zz_12343 = ($signed(twiddle_factor_table_17_real) + $signed(twiddle_factor_table_17_imag));
  assign _zz_12344 = fixTo_870_dout;
  assign _zz_12345 = ($signed(_zz_1190) - $signed(_zz_1189));
  assign _zz_12346 = ($signed(_zz_1189) + $signed(_zz_1190));
  assign _zz_12347 = _zz_12348[15 : 0];
  assign _zz_12348 = fixTo_872_dout;
  assign _zz_12349 = _zz_12350[15 : 0];
  assign _zz_12350 = fixTo_871_dout;
  assign _zz_12351 = _zz_12352;
  assign _zz_12352 = ($signed(_zz_12353) >>> _zz_3246);
  assign _zz_12353 = _zz_12354;
  assign _zz_12354 = ($signed(_zz_1157) - $signed(_zz_3243));
  assign _zz_12355 = _zz_12356;
  assign _zz_12356 = ($signed(_zz_12357) >>> _zz_3246);
  assign _zz_12357 = _zz_12358;
  assign _zz_12358 = ($signed(_zz_1158) - $signed(_zz_3244));
  assign _zz_12359 = _zz_12360;
  assign _zz_12360 = ($signed(_zz_12361) >>> _zz_3247);
  assign _zz_12361 = _zz_12362;
  assign _zz_12362 = ($signed(_zz_1157) + $signed(_zz_3243));
  assign _zz_12363 = _zz_12364;
  assign _zz_12364 = ($signed(_zz_12365) >>> _zz_3247);
  assign _zz_12365 = _zz_12366;
  assign _zz_12366 = ($signed(_zz_1158) + $signed(_zz_3244));
  assign _zz_12367 = ($signed(twiddle_factor_table_18_real) + $signed(twiddle_factor_table_18_imag));
  assign _zz_12368 = fixTo_873_dout;
  assign _zz_12369 = ($signed(_zz_1192) - $signed(_zz_1191));
  assign _zz_12370 = ($signed(_zz_1191) + $signed(_zz_1192));
  assign _zz_12371 = _zz_12372[15 : 0];
  assign _zz_12372 = fixTo_875_dout;
  assign _zz_12373 = _zz_12374[15 : 0];
  assign _zz_12374 = fixTo_874_dout;
  assign _zz_12375 = _zz_12376;
  assign _zz_12376 = ($signed(_zz_12377) >>> _zz_3251);
  assign _zz_12377 = _zz_12378;
  assign _zz_12378 = ($signed(_zz_1159) - $signed(_zz_3248));
  assign _zz_12379 = _zz_12380;
  assign _zz_12380 = ($signed(_zz_12381) >>> _zz_3251);
  assign _zz_12381 = _zz_12382;
  assign _zz_12382 = ($signed(_zz_1160) - $signed(_zz_3249));
  assign _zz_12383 = _zz_12384;
  assign _zz_12384 = ($signed(_zz_12385) >>> _zz_3252);
  assign _zz_12385 = _zz_12386;
  assign _zz_12386 = ($signed(_zz_1159) + $signed(_zz_3248));
  assign _zz_12387 = _zz_12388;
  assign _zz_12388 = ($signed(_zz_12389) >>> _zz_3252);
  assign _zz_12389 = _zz_12390;
  assign _zz_12390 = ($signed(_zz_1160) + $signed(_zz_3249));
  assign _zz_12391 = ($signed(twiddle_factor_table_19_real) + $signed(twiddle_factor_table_19_imag));
  assign _zz_12392 = fixTo_876_dout;
  assign _zz_12393 = ($signed(_zz_1194) - $signed(_zz_1193));
  assign _zz_12394 = ($signed(_zz_1193) + $signed(_zz_1194));
  assign _zz_12395 = _zz_12396[15 : 0];
  assign _zz_12396 = fixTo_878_dout;
  assign _zz_12397 = _zz_12398[15 : 0];
  assign _zz_12398 = fixTo_877_dout;
  assign _zz_12399 = _zz_12400;
  assign _zz_12400 = ($signed(_zz_12401) >>> _zz_3256);
  assign _zz_12401 = _zz_12402;
  assign _zz_12402 = ($signed(_zz_1161) - $signed(_zz_3253));
  assign _zz_12403 = _zz_12404;
  assign _zz_12404 = ($signed(_zz_12405) >>> _zz_3256);
  assign _zz_12405 = _zz_12406;
  assign _zz_12406 = ($signed(_zz_1162) - $signed(_zz_3254));
  assign _zz_12407 = _zz_12408;
  assign _zz_12408 = ($signed(_zz_12409) >>> _zz_3257);
  assign _zz_12409 = _zz_12410;
  assign _zz_12410 = ($signed(_zz_1161) + $signed(_zz_3253));
  assign _zz_12411 = _zz_12412;
  assign _zz_12412 = ($signed(_zz_12413) >>> _zz_3257);
  assign _zz_12413 = _zz_12414;
  assign _zz_12414 = ($signed(_zz_1162) + $signed(_zz_3254));
  assign _zz_12415 = ($signed(twiddle_factor_table_20_real) + $signed(twiddle_factor_table_20_imag));
  assign _zz_12416 = fixTo_879_dout;
  assign _zz_12417 = ($signed(_zz_1196) - $signed(_zz_1195));
  assign _zz_12418 = ($signed(_zz_1195) + $signed(_zz_1196));
  assign _zz_12419 = _zz_12420[15 : 0];
  assign _zz_12420 = fixTo_881_dout;
  assign _zz_12421 = _zz_12422[15 : 0];
  assign _zz_12422 = fixTo_880_dout;
  assign _zz_12423 = _zz_12424;
  assign _zz_12424 = ($signed(_zz_12425) >>> _zz_3261);
  assign _zz_12425 = _zz_12426;
  assign _zz_12426 = ($signed(_zz_1163) - $signed(_zz_3258));
  assign _zz_12427 = _zz_12428;
  assign _zz_12428 = ($signed(_zz_12429) >>> _zz_3261);
  assign _zz_12429 = _zz_12430;
  assign _zz_12430 = ($signed(_zz_1164) - $signed(_zz_3259));
  assign _zz_12431 = _zz_12432;
  assign _zz_12432 = ($signed(_zz_12433) >>> _zz_3262);
  assign _zz_12433 = _zz_12434;
  assign _zz_12434 = ($signed(_zz_1163) + $signed(_zz_3258));
  assign _zz_12435 = _zz_12436;
  assign _zz_12436 = ($signed(_zz_12437) >>> _zz_3262);
  assign _zz_12437 = _zz_12438;
  assign _zz_12438 = ($signed(_zz_1164) + $signed(_zz_3259));
  assign _zz_12439 = ($signed(twiddle_factor_table_21_real) + $signed(twiddle_factor_table_21_imag));
  assign _zz_12440 = fixTo_882_dout;
  assign _zz_12441 = ($signed(_zz_1198) - $signed(_zz_1197));
  assign _zz_12442 = ($signed(_zz_1197) + $signed(_zz_1198));
  assign _zz_12443 = _zz_12444[15 : 0];
  assign _zz_12444 = fixTo_884_dout;
  assign _zz_12445 = _zz_12446[15 : 0];
  assign _zz_12446 = fixTo_883_dout;
  assign _zz_12447 = _zz_12448;
  assign _zz_12448 = ($signed(_zz_12449) >>> _zz_3266);
  assign _zz_12449 = _zz_12450;
  assign _zz_12450 = ($signed(_zz_1165) - $signed(_zz_3263));
  assign _zz_12451 = _zz_12452;
  assign _zz_12452 = ($signed(_zz_12453) >>> _zz_3266);
  assign _zz_12453 = _zz_12454;
  assign _zz_12454 = ($signed(_zz_1166) - $signed(_zz_3264));
  assign _zz_12455 = _zz_12456;
  assign _zz_12456 = ($signed(_zz_12457) >>> _zz_3267);
  assign _zz_12457 = _zz_12458;
  assign _zz_12458 = ($signed(_zz_1165) + $signed(_zz_3263));
  assign _zz_12459 = _zz_12460;
  assign _zz_12460 = ($signed(_zz_12461) >>> _zz_3267);
  assign _zz_12461 = _zz_12462;
  assign _zz_12462 = ($signed(_zz_1166) + $signed(_zz_3264));
  assign _zz_12463 = ($signed(twiddle_factor_table_22_real) + $signed(twiddle_factor_table_22_imag));
  assign _zz_12464 = fixTo_885_dout;
  assign _zz_12465 = ($signed(_zz_1200) - $signed(_zz_1199));
  assign _zz_12466 = ($signed(_zz_1199) + $signed(_zz_1200));
  assign _zz_12467 = _zz_12468[15 : 0];
  assign _zz_12468 = fixTo_887_dout;
  assign _zz_12469 = _zz_12470[15 : 0];
  assign _zz_12470 = fixTo_886_dout;
  assign _zz_12471 = _zz_12472;
  assign _zz_12472 = ($signed(_zz_12473) >>> _zz_3271);
  assign _zz_12473 = _zz_12474;
  assign _zz_12474 = ($signed(_zz_1167) - $signed(_zz_3268));
  assign _zz_12475 = _zz_12476;
  assign _zz_12476 = ($signed(_zz_12477) >>> _zz_3271);
  assign _zz_12477 = _zz_12478;
  assign _zz_12478 = ($signed(_zz_1168) - $signed(_zz_3269));
  assign _zz_12479 = _zz_12480;
  assign _zz_12480 = ($signed(_zz_12481) >>> _zz_3272);
  assign _zz_12481 = _zz_12482;
  assign _zz_12482 = ($signed(_zz_1167) + $signed(_zz_3268));
  assign _zz_12483 = _zz_12484;
  assign _zz_12484 = ($signed(_zz_12485) >>> _zz_3272);
  assign _zz_12485 = _zz_12486;
  assign _zz_12486 = ($signed(_zz_1168) + $signed(_zz_3269));
  assign _zz_12487 = ($signed(twiddle_factor_table_23_real) + $signed(twiddle_factor_table_23_imag));
  assign _zz_12488 = fixTo_888_dout;
  assign _zz_12489 = ($signed(_zz_1202) - $signed(_zz_1201));
  assign _zz_12490 = ($signed(_zz_1201) + $signed(_zz_1202));
  assign _zz_12491 = _zz_12492[15 : 0];
  assign _zz_12492 = fixTo_890_dout;
  assign _zz_12493 = _zz_12494[15 : 0];
  assign _zz_12494 = fixTo_889_dout;
  assign _zz_12495 = _zz_12496;
  assign _zz_12496 = ($signed(_zz_12497) >>> _zz_3276);
  assign _zz_12497 = _zz_12498;
  assign _zz_12498 = ($signed(_zz_1169) - $signed(_zz_3273));
  assign _zz_12499 = _zz_12500;
  assign _zz_12500 = ($signed(_zz_12501) >>> _zz_3276);
  assign _zz_12501 = _zz_12502;
  assign _zz_12502 = ($signed(_zz_1170) - $signed(_zz_3274));
  assign _zz_12503 = _zz_12504;
  assign _zz_12504 = ($signed(_zz_12505) >>> _zz_3277);
  assign _zz_12505 = _zz_12506;
  assign _zz_12506 = ($signed(_zz_1169) + $signed(_zz_3273));
  assign _zz_12507 = _zz_12508;
  assign _zz_12508 = ($signed(_zz_12509) >>> _zz_3277);
  assign _zz_12509 = _zz_12510;
  assign _zz_12510 = ($signed(_zz_1170) + $signed(_zz_3274));
  assign _zz_12511 = ($signed(twiddle_factor_table_24_real) + $signed(twiddle_factor_table_24_imag));
  assign _zz_12512 = fixTo_891_dout;
  assign _zz_12513 = ($signed(_zz_1204) - $signed(_zz_1203));
  assign _zz_12514 = ($signed(_zz_1203) + $signed(_zz_1204));
  assign _zz_12515 = _zz_12516[15 : 0];
  assign _zz_12516 = fixTo_893_dout;
  assign _zz_12517 = _zz_12518[15 : 0];
  assign _zz_12518 = fixTo_892_dout;
  assign _zz_12519 = _zz_12520;
  assign _zz_12520 = ($signed(_zz_12521) >>> _zz_3281);
  assign _zz_12521 = _zz_12522;
  assign _zz_12522 = ($signed(_zz_1171) - $signed(_zz_3278));
  assign _zz_12523 = _zz_12524;
  assign _zz_12524 = ($signed(_zz_12525) >>> _zz_3281);
  assign _zz_12525 = _zz_12526;
  assign _zz_12526 = ($signed(_zz_1172) - $signed(_zz_3279));
  assign _zz_12527 = _zz_12528;
  assign _zz_12528 = ($signed(_zz_12529) >>> _zz_3282);
  assign _zz_12529 = _zz_12530;
  assign _zz_12530 = ($signed(_zz_1171) + $signed(_zz_3278));
  assign _zz_12531 = _zz_12532;
  assign _zz_12532 = ($signed(_zz_12533) >>> _zz_3282);
  assign _zz_12533 = _zz_12534;
  assign _zz_12534 = ($signed(_zz_1172) + $signed(_zz_3279));
  assign _zz_12535 = ($signed(twiddle_factor_table_25_real) + $signed(twiddle_factor_table_25_imag));
  assign _zz_12536 = fixTo_894_dout;
  assign _zz_12537 = ($signed(_zz_1206) - $signed(_zz_1205));
  assign _zz_12538 = ($signed(_zz_1205) + $signed(_zz_1206));
  assign _zz_12539 = _zz_12540[15 : 0];
  assign _zz_12540 = fixTo_896_dout;
  assign _zz_12541 = _zz_12542[15 : 0];
  assign _zz_12542 = fixTo_895_dout;
  assign _zz_12543 = _zz_12544;
  assign _zz_12544 = ($signed(_zz_12545) >>> _zz_3286);
  assign _zz_12545 = _zz_12546;
  assign _zz_12546 = ($signed(_zz_1173) - $signed(_zz_3283));
  assign _zz_12547 = _zz_12548;
  assign _zz_12548 = ($signed(_zz_12549) >>> _zz_3286);
  assign _zz_12549 = _zz_12550;
  assign _zz_12550 = ($signed(_zz_1174) - $signed(_zz_3284));
  assign _zz_12551 = _zz_12552;
  assign _zz_12552 = ($signed(_zz_12553) >>> _zz_3287);
  assign _zz_12553 = _zz_12554;
  assign _zz_12554 = ($signed(_zz_1173) + $signed(_zz_3283));
  assign _zz_12555 = _zz_12556;
  assign _zz_12556 = ($signed(_zz_12557) >>> _zz_3287);
  assign _zz_12557 = _zz_12558;
  assign _zz_12558 = ($signed(_zz_1174) + $signed(_zz_3284));
  assign _zz_12559 = ($signed(twiddle_factor_table_26_real) + $signed(twiddle_factor_table_26_imag));
  assign _zz_12560 = fixTo_897_dout;
  assign _zz_12561 = ($signed(_zz_1208) - $signed(_zz_1207));
  assign _zz_12562 = ($signed(_zz_1207) + $signed(_zz_1208));
  assign _zz_12563 = _zz_12564[15 : 0];
  assign _zz_12564 = fixTo_899_dout;
  assign _zz_12565 = _zz_12566[15 : 0];
  assign _zz_12566 = fixTo_898_dout;
  assign _zz_12567 = _zz_12568;
  assign _zz_12568 = ($signed(_zz_12569) >>> _zz_3291);
  assign _zz_12569 = _zz_12570;
  assign _zz_12570 = ($signed(_zz_1175) - $signed(_zz_3288));
  assign _zz_12571 = _zz_12572;
  assign _zz_12572 = ($signed(_zz_12573) >>> _zz_3291);
  assign _zz_12573 = _zz_12574;
  assign _zz_12574 = ($signed(_zz_1176) - $signed(_zz_3289));
  assign _zz_12575 = _zz_12576;
  assign _zz_12576 = ($signed(_zz_12577) >>> _zz_3292);
  assign _zz_12577 = _zz_12578;
  assign _zz_12578 = ($signed(_zz_1175) + $signed(_zz_3288));
  assign _zz_12579 = _zz_12580;
  assign _zz_12580 = ($signed(_zz_12581) >>> _zz_3292);
  assign _zz_12581 = _zz_12582;
  assign _zz_12582 = ($signed(_zz_1176) + $signed(_zz_3289));
  assign _zz_12583 = ($signed(twiddle_factor_table_27_real) + $signed(twiddle_factor_table_27_imag));
  assign _zz_12584 = fixTo_900_dout;
  assign _zz_12585 = ($signed(_zz_1210) - $signed(_zz_1209));
  assign _zz_12586 = ($signed(_zz_1209) + $signed(_zz_1210));
  assign _zz_12587 = _zz_12588[15 : 0];
  assign _zz_12588 = fixTo_902_dout;
  assign _zz_12589 = _zz_12590[15 : 0];
  assign _zz_12590 = fixTo_901_dout;
  assign _zz_12591 = _zz_12592;
  assign _zz_12592 = ($signed(_zz_12593) >>> _zz_3296);
  assign _zz_12593 = _zz_12594;
  assign _zz_12594 = ($signed(_zz_1177) - $signed(_zz_3293));
  assign _zz_12595 = _zz_12596;
  assign _zz_12596 = ($signed(_zz_12597) >>> _zz_3296);
  assign _zz_12597 = _zz_12598;
  assign _zz_12598 = ($signed(_zz_1178) - $signed(_zz_3294));
  assign _zz_12599 = _zz_12600;
  assign _zz_12600 = ($signed(_zz_12601) >>> _zz_3297);
  assign _zz_12601 = _zz_12602;
  assign _zz_12602 = ($signed(_zz_1177) + $signed(_zz_3293));
  assign _zz_12603 = _zz_12604;
  assign _zz_12604 = ($signed(_zz_12605) >>> _zz_3297);
  assign _zz_12605 = _zz_12606;
  assign _zz_12606 = ($signed(_zz_1178) + $signed(_zz_3294));
  assign _zz_12607 = ($signed(twiddle_factor_table_28_real) + $signed(twiddle_factor_table_28_imag));
  assign _zz_12608 = fixTo_903_dout;
  assign _zz_12609 = ($signed(_zz_1212) - $signed(_zz_1211));
  assign _zz_12610 = ($signed(_zz_1211) + $signed(_zz_1212));
  assign _zz_12611 = _zz_12612[15 : 0];
  assign _zz_12612 = fixTo_905_dout;
  assign _zz_12613 = _zz_12614[15 : 0];
  assign _zz_12614 = fixTo_904_dout;
  assign _zz_12615 = _zz_12616;
  assign _zz_12616 = ($signed(_zz_12617) >>> _zz_3301);
  assign _zz_12617 = _zz_12618;
  assign _zz_12618 = ($signed(_zz_1179) - $signed(_zz_3298));
  assign _zz_12619 = _zz_12620;
  assign _zz_12620 = ($signed(_zz_12621) >>> _zz_3301);
  assign _zz_12621 = _zz_12622;
  assign _zz_12622 = ($signed(_zz_1180) - $signed(_zz_3299));
  assign _zz_12623 = _zz_12624;
  assign _zz_12624 = ($signed(_zz_12625) >>> _zz_3302);
  assign _zz_12625 = _zz_12626;
  assign _zz_12626 = ($signed(_zz_1179) + $signed(_zz_3298));
  assign _zz_12627 = _zz_12628;
  assign _zz_12628 = ($signed(_zz_12629) >>> _zz_3302);
  assign _zz_12629 = _zz_12630;
  assign _zz_12630 = ($signed(_zz_1180) + $signed(_zz_3299));
  assign _zz_12631 = ($signed(twiddle_factor_table_29_real) + $signed(twiddle_factor_table_29_imag));
  assign _zz_12632 = fixTo_906_dout;
  assign _zz_12633 = ($signed(_zz_1214) - $signed(_zz_1213));
  assign _zz_12634 = ($signed(_zz_1213) + $signed(_zz_1214));
  assign _zz_12635 = _zz_12636[15 : 0];
  assign _zz_12636 = fixTo_908_dout;
  assign _zz_12637 = _zz_12638[15 : 0];
  assign _zz_12638 = fixTo_907_dout;
  assign _zz_12639 = _zz_12640;
  assign _zz_12640 = ($signed(_zz_12641) >>> _zz_3306);
  assign _zz_12641 = _zz_12642;
  assign _zz_12642 = ($signed(_zz_1181) - $signed(_zz_3303));
  assign _zz_12643 = _zz_12644;
  assign _zz_12644 = ($signed(_zz_12645) >>> _zz_3306);
  assign _zz_12645 = _zz_12646;
  assign _zz_12646 = ($signed(_zz_1182) - $signed(_zz_3304));
  assign _zz_12647 = _zz_12648;
  assign _zz_12648 = ($signed(_zz_12649) >>> _zz_3307);
  assign _zz_12649 = _zz_12650;
  assign _zz_12650 = ($signed(_zz_1181) + $signed(_zz_3303));
  assign _zz_12651 = _zz_12652;
  assign _zz_12652 = ($signed(_zz_12653) >>> _zz_3307);
  assign _zz_12653 = _zz_12654;
  assign _zz_12654 = ($signed(_zz_1182) + $signed(_zz_3304));
  assign _zz_12655 = ($signed(twiddle_factor_table_30_real) + $signed(twiddle_factor_table_30_imag));
  assign _zz_12656 = fixTo_909_dout;
  assign _zz_12657 = ($signed(_zz_1216) - $signed(_zz_1215));
  assign _zz_12658 = ($signed(_zz_1215) + $signed(_zz_1216));
  assign _zz_12659 = _zz_12660[15 : 0];
  assign _zz_12660 = fixTo_911_dout;
  assign _zz_12661 = _zz_12662[15 : 0];
  assign _zz_12662 = fixTo_910_dout;
  assign _zz_12663 = _zz_12664;
  assign _zz_12664 = ($signed(_zz_12665) >>> _zz_3311);
  assign _zz_12665 = _zz_12666;
  assign _zz_12666 = ($signed(_zz_1183) - $signed(_zz_3308));
  assign _zz_12667 = _zz_12668;
  assign _zz_12668 = ($signed(_zz_12669) >>> _zz_3311);
  assign _zz_12669 = _zz_12670;
  assign _zz_12670 = ($signed(_zz_1184) - $signed(_zz_3309));
  assign _zz_12671 = _zz_12672;
  assign _zz_12672 = ($signed(_zz_12673) >>> _zz_3312);
  assign _zz_12673 = _zz_12674;
  assign _zz_12674 = ($signed(_zz_1183) + $signed(_zz_3308));
  assign _zz_12675 = _zz_12676;
  assign _zz_12676 = ($signed(_zz_12677) >>> _zz_3312);
  assign _zz_12677 = _zz_12678;
  assign _zz_12678 = ($signed(_zz_1184) + $signed(_zz_3309));
  assign _zz_12679 = ($signed(twiddle_factor_table_15_real) + $signed(twiddle_factor_table_15_imag));
  assign _zz_12680 = fixTo_912_dout;
  assign _zz_12681 = ($signed(_zz_1250) - $signed(_zz_1249));
  assign _zz_12682 = ($signed(_zz_1249) + $signed(_zz_1250));
  assign _zz_12683 = _zz_12684[15 : 0];
  assign _zz_12684 = fixTo_914_dout;
  assign _zz_12685 = _zz_12686[15 : 0];
  assign _zz_12686 = fixTo_913_dout;
  assign _zz_12687 = _zz_12688;
  assign _zz_12688 = ($signed(_zz_12689) >>> _zz_3316);
  assign _zz_12689 = _zz_12690;
  assign _zz_12690 = ($signed(_zz_1217) - $signed(_zz_3313));
  assign _zz_12691 = _zz_12692;
  assign _zz_12692 = ($signed(_zz_12693) >>> _zz_3316);
  assign _zz_12693 = _zz_12694;
  assign _zz_12694 = ($signed(_zz_1218) - $signed(_zz_3314));
  assign _zz_12695 = _zz_12696;
  assign _zz_12696 = ($signed(_zz_12697) >>> _zz_3317);
  assign _zz_12697 = _zz_12698;
  assign _zz_12698 = ($signed(_zz_1217) + $signed(_zz_3313));
  assign _zz_12699 = _zz_12700;
  assign _zz_12700 = ($signed(_zz_12701) >>> _zz_3317);
  assign _zz_12701 = _zz_12702;
  assign _zz_12702 = ($signed(_zz_1218) + $signed(_zz_3314));
  assign _zz_12703 = ($signed(twiddle_factor_table_16_real) + $signed(twiddle_factor_table_16_imag));
  assign _zz_12704 = fixTo_915_dout;
  assign _zz_12705 = ($signed(_zz_1252) - $signed(_zz_1251));
  assign _zz_12706 = ($signed(_zz_1251) + $signed(_zz_1252));
  assign _zz_12707 = _zz_12708[15 : 0];
  assign _zz_12708 = fixTo_917_dout;
  assign _zz_12709 = _zz_12710[15 : 0];
  assign _zz_12710 = fixTo_916_dout;
  assign _zz_12711 = _zz_12712;
  assign _zz_12712 = ($signed(_zz_12713) >>> _zz_3321);
  assign _zz_12713 = _zz_12714;
  assign _zz_12714 = ($signed(_zz_1219) - $signed(_zz_3318));
  assign _zz_12715 = _zz_12716;
  assign _zz_12716 = ($signed(_zz_12717) >>> _zz_3321);
  assign _zz_12717 = _zz_12718;
  assign _zz_12718 = ($signed(_zz_1220) - $signed(_zz_3319));
  assign _zz_12719 = _zz_12720;
  assign _zz_12720 = ($signed(_zz_12721) >>> _zz_3322);
  assign _zz_12721 = _zz_12722;
  assign _zz_12722 = ($signed(_zz_1219) + $signed(_zz_3318));
  assign _zz_12723 = _zz_12724;
  assign _zz_12724 = ($signed(_zz_12725) >>> _zz_3322);
  assign _zz_12725 = _zz_12726;
  assign _zz_12726 = ($signed(_zz_1220) + $signed(_zz_3319));
  assign _zz_12727 = ($signed(twiddle_factor_table_17_real) + $signed(twiddle_factor_table_17_imag));
  assign _zz_12728 = fixTo_918_dout;
  assign _zz_12729 = ($signed(_zz_1254) - $signed(_zz_1253));
  assign _zz_12730 = ($signed(_zz_1253) + $signed(_zz_1254));
  assign _zz_12731 = _zz_12732[15 : 0];
  assign _zz_12732 = fixTo_920_dout;
  assign _zz_12733 = _zz_12734[15 : 0];
  assign _zz_12734 = fixTo_919_dout;
  assign _zz_12735 = _zz_12736;
  assign _zz_12736 = ($signed(_zz_12737) >>> _zz_3326);
  assign _zz_12737 = _zz_12738;
  assign _zz_12738 = ($signed(_zz_1221) - $signed(_zz_3323));
  assign _zz_12739 = _zz_12740;
  assign _zz_12740 = ($signed(_zz_12741) >>> _zz_3326);
  assign _zz_12741 = _zz_12742;
  assign _zz_12742 = ($signed(_zz_1222) - $signed(_zz_3324));
  assign _zz_12743 = _zz_12744;
  assign _zz_12744 = ($signed(_zz_12745) >>> _zz_3327);
  assign _zz_12745 = _zz_12746;
  assign _zz_12746 = ($signed(_zz_1221) + $signed(_zz_3323));
  assign _zz_12747 = _zz_12748;
  assign _zz_12748 = ($signed(_zz_12749) >>> _zz_3327);
  assign _zz_12749 = _zz_12750;
  assign _zz_12750 = ($signed(_zz_1222) + $signed(_zz_3324));
  assign _zz_12751 = ($signed(twiddle_factor_table_18_real) + $signed(twiddle_factor_table_18_imag));
  assign _zz_12752 = fixTo_921_dout;
  assign _zz_12753 = ($signed(_zz_1256) - $signed(_zz_1255));
  assign _zz_12754 = ($signed(_zz_1255) + $signed(_zz_1256));
  assign _zz_12755 = _zz_12756[15 : 0];
  assign _zz_12756 = fixTo_923_dout;
  assign _zz_12757 = _zz_12758[15 : 0];
  assign _zz_12758 = fixTo_922_dout;
  assign _zz_12759 = _zz_12760;
  assign _zz_12760 = ($signed(_zz_12761) >>> _zz_3331);
  assign _zz_12761 = _zz_12762;
  assign _zz_12762 = ($signed(_zz_1223) - $signed(_zz_3328));
  assign _zz_12763 = _zz_12764;
  assign _zz_12764 = ($signed(_zz_12765) >>> _zz_3331);
  assign _zz_12765 = _zz_12766;
  assign _zz_12766 = ($signed(_zz_1224) - $signed(_zz_3329));
  assign _zz_12767 = _zz_12768;
  assign _zz_12768 = ($signed(_zz_12769) >>> _zz_3332);
  assign _zz_12769 = _zz_12770;
  assign _zz_12770 = ($signed(_zz_1223) + $signed(_zz_3328));
  assign _zz_12771 = _zz_12772;
  assign _zz_12772 = ($signed(_zz_12773) >>> _zz_3332);
  assign _zz_12773 = _zz_12774;
  assign _zz_12774 = ($signed(_zz_1224) + $signed(_zz_3329));
  assign _zz_12775 = ($signed(twiddle_factor_table_19_real) + $signed(twiddle_factor_table_19_imag));
  assign _zz_12776 = fixTo_924_dout;
  assign _zz_12777 = ($signed(_zz_1258) - $signed(_zz_1257));
  assign _zz_12778 = ($signed(_zz_1257) + $signed(_zz_1258));
  assign _zz_12779 = _zz_12780[15 : 0];
  assign _zz_12780 = fixTo_926_dout;
  assign _zz_12781 = _zz_12782[15 : 0];
  assign _zz_12782 = fixTo_925_dout;
  assign _zz_12783 = _zz_12784;
  assign _zz_12784 = ($signed(_zz_12785) >>> _zz_3336);
  assign _zz_12785 = _zz_12786;
  assign _zz_12786 = ($signed(_zz_1225) - $signed(_zz_3333));
  assign _zz_12787 = _zz_12788;
  assign _zz_12788 = ($signed(_zz_12789) >>> _zz_3336);
  assign _zz_12789 = _zz_12790;
  assign _zz_12790 = ($signed(_zz_1226) - $signed(_zz_3334));
  assign _zz_12791 = _zz_12792;
  assign _zz_12792 = ($signed(_zz_12793) >>> _zz_3337);
  assign _zz_12793 = _zz_12794;
  assign _zz_12794 = ($signed(_zz_1225) + $signed(_zz_3333));
  assign _zz_12795 = _zz_12796;
  assign _zz_12796 = ($signed(_zz_12797) >>> _zz_3337);
  assign _zz_12797 = _zz_12798;
  assign _zz_12798 = ($signed(_zz_1226) + $signed(_zz_3334));
  assign _zz_12799 = ($signed(twiddle_factor_table_20_real) + $signed(twiddle_factor_table_20_imag));
  assign _zz_12800 = fixTo_927_dout;
  assign _zz_12801 = ($signed(_zz_1260) - $signed(_zz_1259));
  assign _zz_12802 = ($signed(_zz_1259) + $signed(_zz_1260));
  assign _zz_12803 = _zz_12804[15 : 0];
  assign _zz_12804 = fixTo_929_dout;
  assign _zz_12805 = _zz_12806[15 : 0];
  assign _zz_12806 = fixTo_928_dout;
  assign _zz_12807 = _zz_12808;
  assign _zz_12808 = ($signed(_zz_12809) >>> _zz_3341);
  assign _zz_12809 = _zz_12810;
  assign _zz_12810 = ($signed(_zz_1227) - $signed(_zz_3338));
  assign _zz_12811 = _zz_12812;
  assign _zz_12812 = ($signed(_zz_12813) >>> _zz_3341);
  assign _zz_12813 = _zz_12814;
  assign _zz_12814 = ($signed(_zz_1228) - $signed(_zz_3339));
  assign _zz_12815 = _zz_12816;
  assign _zz_12816 = ($signed(_zz_12817) >>> _zz_3342);
  assign _zz_12817 = _zz_12818;
  assign _zz_12818 = ($signed(_zz_1227) + $signed(_zz_3338));
  assign _zz_12819 = _zz_12820;
  assign _zz_12820 = ($signed(_zz_12821) >>> _zz_3342);
  assign _zz_12821 = _zz_12822;
  assign _zz_12822 = ($signed(_zz_1228) + $signed(_zz_3339));
  assign _zz_12823 = ($signed(twiddle_factor_table_21_real) + $signed(twiddle_factor_table_21_imag));
  assign _zz_12824 = fixTo_930_dout;
  assign _zz_12825 = ($signed(_zz_1262) - $signed(_zz_1261));
  assign _zz_12826 = ($signed(_zz_1261) + $signed(_zz_1262));
  assign _zz_12827 = _zz_12828[15 : 0];
  assign _zz_12828 = fixTo_932_dout;
  assign _zz_12829 = _zz_12830[15 : 0];
  assign _zz_12830 = fixTo_931_dout;
  assign _zz_12831 = _zz_12832;
  assign _zz_12832 = ($signed(_zz_12833) >>> _zz_3346);
  assign _zz_12833 = _zz_12834;
  assign _zz_12834 = ($signed(_zz_1229) - $signed(_zz_3343));
  assign _zz_12835 = _zz_12836;
  assign _zz_12836 = ($signed(_zz_12837) >>> _zz_3346);
  assign _zz_12837 = _zz_12838;
  assign _zz_12838 = ($signed(_zz_1230) - $signed(_zz_3344));
  assign _zz_12839 = _zz_12840;
  assign _zz_12840 = ($signed(_zz_12841) >>> _zz_3347);
  assign _zz_12841 = _zz_12842;
  assign _zz_12842 = ($signed(_zz_1229) + $signed(_zz_3343));
  assign _zz_12843 = _zz_12844;
  assign _zz_12844 = ($signed(_zz_12845) >>> _zz_3347);
  assign _zz_12845 = _zz_12846;
  assign _zz_12846 = ($signed(_zz_1230) + $signed(_zz_3344));
  assign _zz_12847 = ($signed(twiddle_factor_table_22_real) + $signed(twiddle_factor_table_22_imag));
  assign _zz_12848 = fixTo_933_dout;
  assign _zz_12849 = ($signed(_zz_1264) - $signed(_zz_1263));
  assign _zz_12850 = ($signed(_zz_1263) + $signed(_zz_1264));
  assign _zz_12851 = _zz_12852[15 : 0];
  assign _zz_12852 = fixTo_935_dout;
  assign _zz_12853 = _zz_12854[15 : 0];
  assign _zz_12854 = fixTo_934_dout;
  assign _zz_12855 = _zz_12856;
  assign _zz_12856 = ($signed(_zz_12857) >>> _zz_3351);
  assign _zz_12857 = _zz_12858;
  assign _zz_12858 = ($signed(_zz_1231) - $signed(_zz_3348));
  assign _zz_12859 = _zz_12860;
  assign _zz_12860 = ($signed(_zz_12861) >>> _zz_3351);
  assign _zz_12861 = _zz_12862;
  assign _zz_12862 = ($signed(_zz_1232) - $signed(_zz_3349));
  assign _zz_12863 = _zz_12864;
  assign _zz_12864 = ($signed(_zz_12865) >>> _zz_3352);
  assign _zz_12865 = _zz_12866;
  assign _zz_12866 = ($signed(_zz_1231) + $signed(_zz_3348));
  assign _zz_12867 = _zz_12868;
  assign _zz_12868 = ($signed(_zz_12869) >>> _zz_3352);
  assign _zz_12869 = _zz_12870;
  assign _zz_12870 = ($signed(_zz_1232) + $signed(_zz_3349));
  assign _zz_12871 = ($signed(twiddle_factor_table_23_real) + $signed(twiddle_factor_table_23_imag));
  assign _zz_12872 = fixTo_936_dout;
  assign _zz_12873 = ($signed(_zz_1266) - $signed(_zz_1265));
  assign _zz_12874 = ($signed(_zz_1265) + $signed(_zz_1266));
  assign _zz_12875 = _zz_12876[15 : 0];
  assign _zz_12876 = fixTo_938_dout;
  assign _zz_12877 = _zz_12878[15 : 0];
  assign _zz_12878 = fixTo_937_dout;
  assign _zz_12879 = _zz_12880;
  assign _zz_12880 = ($signed(_zz_12881) >>> _zz_3356);
  assign _zz_12881 = _zz_12882;
  assign _zz_12882 = ($signed(_zz_1233) - $signed(_zz_3353));
  assign _zz_12883 = _zz_12884;
  assign _zz_12884 = ($signed(_zz_12885) >>> _zz_3356);
  assign _zz_12885 = _zz_12886;
  assign _zz_12886 = ($signed(_zz_1234) - $signed(_zz_3354));
  assign _zz_12887 = _zz_12888;
  assign _zz_12888 = ($signed(_zz_12889) >>> _zz_3357);
  assign _zz_12889 = _zz_12890;
  assign _zz_12890 = ($signed(_zz_1233) + $signed(_zz_3353));
  assign _zz_12891 = _zz_12892;
  assign _zz_12892 = ($signed(_zz_12893) >>> _zz_3357);
  assign _zz_12893 = _zz_12894;
  assign _zz_12894 = ($signed(_zz_1234) + $signed(_zz_3354));
  assign _zz_12895 = ($signed(twiddle_factor_table_24_real) + $signed(twiddle_factor_table_24_imag));
  assign _zz_12896 = fixTo_939_dout;
  assign _zz_12897 = ($signed(_zz_1268) - $signed(_zz_1267));
  assign _zz_12898 = ($signed(_zz_1267) + $signed(_zz_1268));
  assign _zz_12899 = _zz_12900[15 : 0];
  assign _zz_12900 = fixTo_941_dout;
  assign _zz_12901 = _zz_12902[15 : 0];
  assign _zz_12902 = fixTo_940_dout;
  assign _zz_12903 = _zz_12904;
  assign _zz_12904 = ($signed(_zz_12905) >>> _zz_3361);
  assign _zz_12905 = _zz_12906;
  assign _zz_12906 = ($signed(_zz_1235) - $signed(_zz_3358));
  assign _zz_12907 = _zz_12908;
  assign _zz_12908 = ($signed(_zz_12909) >>> _zz_3361);
  assign _zz_12909 = _zz_12910;
  assign _zz_12910 = ($signed(_zz_1236) - $signed(_zz_3359));
  assign _zz_12911 = _zz_12912;
  assign _zz_12912 = ($signed(_zz_12913) >>> _zz_3362);
  assign _zz_12913 = _zz_12914;
  assign _zz_12914 = ($signed(_zz_1235) + $signed(_zz_3358));
  assign _zz_12915 = _zz_12916;
  assign _zz_12916 = ($signed(_zz_12917) >>> _zz_3362);
  assign _zz_12917 = _zz_12918;
  assign _zz_12918 = ($signed(_zz_1236) + $signed(_zz_3359));
  assign _zz_12919 = ($signed(twiddle_factor_table_25_real) + $signed(twiddle_factor_table_25_imag));
  assign _zz_12920 = fixTo_942_dout;
  assign _zz_12921 = ($signed(_zz_1270) - $signed(_zz_1269));
  assign _zz_12922 = ($signed(_zz_1269) + $signed(_zz_1270));
  assign _zz_12923 = _zz_12924[15 : 0];
  assign _zz_12924 = fixTo_944_dout;
  assign _zz_12925 = _zz_12926[15 : 0];
  assign _zz_12926 = fixTo_943_dout;
  assign _zz_12927 = _zz_12928;
  assign _zz_12928 = ($signed(_zz_12929) >>> _zz_3366);
  assign _zz_12929 = _zz_12930;
  assign _zz_12930 = ($signed(_zz_1237) - $signed(_zz_3363));
  assign _zz_12931 = _zz_12932;
  assign _zz_12932 = ($signed(_zz_12933) >>> _zz_3366);
  assign _zz_12933 = _zz_12934;
  assign _zz_12934 = ($signed(_zz_1238) - $signed(_zz_3364));
  assign _zz_12935 = _zz_12936;
  assign _zz_12936 = ($signed(_zz_12937) >>> _zz_3367);
  assign _zz_12937 = _zz_12938;
  assign _zz_12938 = ($signed(_zz_1237) + $signed(_zz_3363));
  assign _zz_12939 = _zz_12940;
  assign _zz_12940 = ($signed(_zz_12941) >>> _zz_3367);
  assign _zz_12941 = _zz_12942;
  assign _zz_12942 = ($signed(_zz_1238) + $signed(_zz_3364));
  assign _zz_12943 = ($signed(twiddle_factor_table_26_real) + $signed(twiddle_factor_table_26_imag));
  assign _zz_12944 = fixTo_945_dout;
  assign _zz_12945 = ($signed(_zz_1272) - $signed(_zz_1271));
  assign _zz_12946 = ($signed(_zz_1271) + $signed(_zz_1272));
  assign _zz_12947 = _zz_12948[15 : 0];
  assign _zz_12948 = fixTo_947_dout;
  assign _zz_12949 = _zz_12950[15 : 0];
  assign _zz_12950 = fixTo_946_dout;
  assign _zz_12951 = _zz_12952;
  assign _zz_12952 = ($signed(_zz_12953) >>> _zz_3371);
  assign _zz_12953 = _zz_12954;
  assign _zz_12954 = ($signed(_zz_1239) - $signed(_zz_3368));
  assign _zz_12955 = _zz_12956;
  assign _zz_12956 = ($signed(_zz_12957) >>> _zz_3371);
  assign _zz_12957 = _zz_12958;
  assign _zz_12958 = ($signed(_zz_1240) - $signed(_zz_3369));
  assign _zz_12959 = _zz_12960;
  assign _zz_12960 = ($signed(_zz_12961) >>> _zz_3372);
  assign _zz_12961 = _zz_12962;
  assign _zz_12962 = ($signed(_zz_1239) + $signed(_zz_3368));
  assign _zz_12963 = _zz_12964;
  assign _zz_12964 = ($signed(_zz_12965) >>> _zz_3372);
  assign _zz_12965 = _zz_12966;
  assign _zz_12966 = ($signed(_zz_1240) + $signed(_zz_3369));
  assign _zz_12967 = ($signed(twiddle_factor_table_27_real) + $signed(twiddle_factor_table_27_imag));
  assign _zz_12968 = fixTo_948_dout;
  assign _zz_12969 = ($signed(_zz_1274) - $signed(_zz_1273));
  assign _zz_12970 = ($signed(_zz_1273) + $signed(_zz_1274));
  assign _zz_12971 = _zz_12972[15 : 0];
  assign _zz_12972 = fixTo_950_dout;
  assign _zz_12973 = _zz_12974[15 : 0];
  assign _zz_12974 = fixTo_949_dout;
  assign _zz_12975 = _zz_12976;
  assign _zz_12976 = ($signed(_zz_12977) >>> _zz_3376);
  assign _zz_12977 = _zz_12978;
  assign _zz_12978 = ($signed(_zz_1241) - $signed(_zz_3373));
  assign _zz_12979 = _zz_12980;
  assign _zz_12980 = ($signed(_zz_12981) >>> _zz_3376);
  assign _zz_12981 = _zz_12982;
  assign _zz_12982 = ($signed(_zz_1242) - $signed(_zz_3374));
  assign _zz_12983 = _zz_12984;
  assign _zz_12984 = ($signed(_zz_12985) >>> _zz_3377);
  assign _zz_12985 = _zz_12986;
  assign _zz_12986 = ($signed(_zz_1241) + $signed(_zz_3373));
  assign _zz_12987 = _zz_12988;
  assign _zz_12988 = ($signed(_zz_12989) >>> _zz_3377);
  assign _zz_12989 = _zz_12990;
  assign _zz_12990 = ($signed(_zz_1242) + $signed(_zz_3374));
  assign _zz_12991 = ($signed(twiddle_factor_table_28_real) + $signed(twiddle_factor_table_28_imag));
  assign _zz_12992 = fixTo_951_dout;
  assign _zz_12993 = ($signed(_zz_1276) - $signed(_zz_1275));
  assign _zz_12994 = ($signed(_zz_1275) + $signed(_zz_1276));
  assign _zz_12995 = _zz_12996[15 : 0];
  assign _zz_12996 = fixTo_953_dout;
  assign _zz_12997 = _zz_12998[15 : 0];
  assign _zz_12998 = fixTo_952_dout;
  assign _zz_12999 = _zz_13000;
  assign _zz_13000 = ($signed(_zz_13001) >>> _zz_3381);
  assign _zz_13001 = _zz_13002;
  assign _zz_13002 = ($signed(_zz_1243) - $signed(_zz_3378));
  assign _zz_13003 = _zz_13004;
  assign _zz_13004 = ($signed(_zz_13005) >>> _zz_3381);
  assign _zz_13005 = _zz_13006;
  assign _zz_13006 = ($signed(_zz_1244) - $signed(_zz_3379));
  assign _zz_13007 = _zz_13008;
  assign _zz_13008 = ($signed(_zz_13009) >>> _zz_3382);
  assign _zz_13009 = _zz_13010;
  assign _zz_13010 = ($signed(_zz_1243) + $signed(_zz_3378));
  assign _zz_13011 = _zz_13012;
  assign _zz_13012 = ($signed(_zz_13013) >>> _zz_3382);
  assign _zz_13013 = _zz_13014;
  assign _zz_13014 = ($signed(_zz_1244) + $signed(_zz_3379));
  assign _zz_13015 = ($signed(twiddle_factor_table_29_real) + $signed(twiddle_factor_table_29_imag));
  assign _zz_13016 = fixTo_954_dout;
  assign _zz_13017 = ($signed(_zz_1278) - $signed(_zz_1277));
  assign _zz_13018 = ($signed(_zz_1277) + $signed(_zz_1278));
  assign _zz_13019 = _zz_13020[15 : 0];
  assign _zz_13020 = fixTo_956_dout;
  assign _zz_13021 = _zz_13022[15 : 0];
  assign _zz_13022 = fixTo_955_dout;
  assign _zz_13023 = _zz_13024;
  assign _zz_13024 = ($signed(_zz_13025) >>> _zz_3386);
  assign _zz_13025 = _zz_13026;
  assign _zz_13026 = ($signed(_zz_1245) - $signed(_zz_3383));
  assign _zz_13027 = _zz_13028;
  assign _zz_13028 = ($signed(_zz_13029) >>> _zz_3386);
  assign _zz_13029 = _zz_13030;
  assign _zz_13030 = ($signed(_zz_1246) - $signed(_zz_3384));
  assign _zz_13031 = _zz_13032;
  assign _zz_13032 = ($signed(_zz_13033) >>> _zz_3387);
  assign _zz_13033 = _zz_13034;
  assign _zz_13034 = ($signed(_zz_1245) + $signed(_zz_3383));
  assign _zz_13035 = _zz_13036;
  assign _zz_13036 = ($signed(_zz_13037) >>> _zz_3387);
  assign _zz_13037 = _zz_13038;
  assign _zz_13038 = ($signed(_zz_1246) + $signed(_zz_3384));
  assign _zz_13039 = ($signed(twiddle_factor_table_30_real) + $signed(twiddle_factor_table_30_imag));
  assign _zz_13040 = fixTo_957_dout;
  assign _zz_13041 = ($signed(_zz_1280) - $signed(_zz_1279));
  assign _zz_13042 = ($signed(_zz_1279) + $signed(_zz_1280));
  assign _zz_13043 = _zz_13044[15 : 0];
  assign _zz_13044 = fixTo_959_dout;
  assign _zz_13045 = _zz_13046[15 : 0];
  assign _zz_13046 = fixTo_958_dout;
  assign _zz_13047 = _zz_13048;
  assign _zz_13048 = ($signed(_zz_13049) >>> _zz_3391);
  assign _zz_13049 = _zz_13050;
  assign _zz_13050 = ($signed(_zz_1247) - $signed(_zz_3388));
  assign _zz_13051 = _zz_13052;
  assign _zz_13052 = ($signed(_zz_13053) >>> _zz_3391);
  assign _zz_13053 = _zz_13054;
  assign _zz_13054 = ($signed(_zz_1248) - $signed(_zz_3389));
  assign _zz_13055 = _zz_13056;
  assign _zz_13056 = ($signed(_zz_13057) >>> _zz_3392);
  assign _zz_13057 = _zz_13058;
  assign _zz_13058 = ($signed(_zz_1247) + $signed(_zz_3388));
  assign _zz_13059 = _zz_13060;
  assign _zz_13060 = ($signed(_zz_13061) >>> _zz_3392);
  assign _zz_13061 = _zz_13062;
  assign _zz_13062 = ($signed(_zz_1248) + $signed(_zz_3389));
  assign _zz_13063 = ($signed(twiddle_factor_table_31_real) + $signed(twiddle_factor_table_31_imag));
  assign _zz_13064 = fixTo_960_dout;
  assign _zz_13065 = ($signed(_zz_1346) - $signed(_zz_1345));
  assign _zz_13066 = ($signed(_zz_1345) + $signed(_zz_1346));
  assign _zz_13067 = _zz_13068[15 : 0];
  assign _zz_13068 = fixTo_962_dout;
  assign _zz_13069 = _zz_13070[15 : 0];
  assign _zz_13070 = fixTo_961_dout;
  assign _zz_13071 = _zz_13072;
  assign _zz_13072 = ($signed(_zz_13073) >>> _zz_3396);
  assign _zz_13073 = _zz_13074;
  assign _zz_13074 = ($signed(_zz_1281) - $signed(_zz_3393));
  assign _zz_13075 = _zz_13076;
  assign _zz_13076 = ($signed(_zz_13077) >>> _zz_3396);
  assign _zz_13077 = _zz_13078;
  assign _zz_13078 = ($signed(_zz_1282) - $signed(_zz_3394));
  assign _zz_13079 = _zz_13080;
  assign _zz_13080 = ($signed(_zz_13081) >>> _zz_3397);
  assign _zz_13081 = _zz_13082;
  assign _zz_13082 = ($signed(_zz_1281) + $signed(_zz_3393));
  assign _zz_13083 = _zz_13084;
  assign _zz_13084 = ($signed(_zz_13085) >>> _zz_3397);
  assign _zz_13085 = _zz_13086;
  assign _zz_13086 = ($signed(_zz_1282) + $signed(_zz_3394));
  assign _zz_13087 = ($signed(twiddle_factor_table_32_real) + $signed(twiddle_factor_table_32_imag));
  assign _zz_13088 = fixTo_963_dout;
  assign _zz_13089 = ($signed(_zz_1348) - $signed(_zz_1347));
  assign _zz_13090 = ($signed(_zz_1347) + $signed(_zz_1348));
  assign _zz_13091 = _zz_13092[15 : 0];
  assign _zz_13092 = fixTo_965_dout;
  assign _zz_13093 = _zz_13094[15 : 0];
  assign _zz_13094 = fixTo_964_dout;
  assign _zz_13095 = _zz_13096;
  assign _zz_13096 = ($signed(_zz_13097) >>> _zz_3401);
  assign _zz_13097 = _zz_13098;
  assign _zz_13098 = ($signed(_zz_1283) - $signed(_zz_3398));
  assign _zz_13099 = _zz_13100;
  assign _zz_13100 = ($signed(_zz_13101) >>> _zz_3401);
  assign _zz_13101 = _zz_13102;
  assign _zz_13102 = ($signed(_zz_1284) - $signed(_zz_3399));
  assign _zz_13103 = _zz_13104;
  assign _zz_13104 = ($signed(_zz_13105) >>> _zz_3402);
  assign _zz_13105 = _zz_13106;
  assign _zz_13106 = ($signed(_zz_1283) + $signed(_zz_3398));
  assign _zz_13107 = _zz_13108;
  assign _zz_13108 = ($signed(_zz_13109) >>> _zz_3402);
  assign _zz_13109 = _zz_13110;
  assign _zz_13110 = ($signed(_zz_1284) + $signed(_zz_3399));
  assign _zz_13111 = ($signed(twiddle_factor_table_33_real) + $signed(twiddle_factor_table_33_imag));
  assign _zz_13112 = fixTo_966_dout;
  assign _zz_13113 = ($signed(_zz_1350) - $signed(_zz_1349));
  assign _zz_13114 = ($signed(_zz_1349) + $signed(_zz_1350));
  assign _zz_13115 = _zz_13116[15 : 0];
  assign _zz_13116 = fixTo_968_dout;
  assign _zz_13117 = _zz_13118[15 : 0];
  assign _zz_13118 = fixTo_967_dout;
  assign _zz_13119 = _zz_13120;
  assign _zz_13120 = ($signed(_zz_13121) >>> _zz_3406);
  assign _zz_13121 = _zz_13122;
  assign _zz_13122 = ($signed(_zz_1285) - $signed(_zz_3403));
  assign _zz_13123 = _zz_13124;
  assign _zz_13124 = ($signed(_zz_13125) >>> _zz_3406);
  assign _zz_13125 = _zz_13126;
  assign _zz_13126 = ($signed(_zz_1286) - $signed(_zz_3404));
  assign _zz_13127 = _zz_13128;
  assign _zz_13128 = ($signed(_zz_13129) >>> _zz_3407);
  assign _zz_13129 = _zz_13130;
  assign _zz_13130 = ($signed(_zz_1285) + $signed(_zz_3403));
  assign _zz_13131 = _zz_13132;
  assign _zz_13132 = ($signed(_zz_13133) >>> _zz_3407);
  assign _zz_13133 = _zz_13134;
  assign _zz_13134 = ($signed(_zz_1286) + $signed(_zz_3404));
  assign _zz_13135 = ($signed(twiddle_factor_table_34_real) + $signed(twiddle_factor_table_34_imag));
  assign _zz_13136 = fixTo_969_dout;
  assign _zz_13137 = ($signed(_zz_1352) - $signed(_zz_1351));
  assign _zz_13138 = ($signed(_zz_1351) + $signed(_zz_1352));
  assign _zz_13139 = _zz_13140[15 : 0];
  assign _zz_13140 = fixTo_971_dout;
  assign _zz_13141 = _zz_13142[15 : 0];
  assign _zz_13142 = fixTo_970_dout;
  assign _zz_13143 = _zz_13144;
  assign _zz_13144 = ($signed(_zz_13145) >>> _zz_3411);
  assign _zz_13145 = _zz_13146;
  assign _zz_13146 = ($signed(_zz_1287) - $signed(_zz_3408));
  assign _zz_13147 = _zz_13148;
  assign _zz_13148 = ($signed(_zz_13149) >>> _zz_3411);
  assign _zz_13149 = _zz_13150;
  assign _zz_13150 = ($signed(_zz_1288) - $signed(_zz_3409));
  assign _zz_13151 = _zz_13152;
  assign _zz_13152 = ($signed(_zz_13153) >>> _zz_3412);
  assign _zz_13153 = _zz_13154;
  assign _zz_13154 = ($signed(_zz_1287) + $signed(_zz_3408));
  assign _zz_13155 = _zz_13156;
  assign _zz_13156 = ($signed(_zz_13157) >>> _zz_3412);
  assign _zz_13157 = _zz_13158;
  assign _zz_13158 = ($signed(_zz_1288) + $signed(_zz_3409));
  assign _zz_13159 = ($signed(twiddle_factor_table_35_real) + $signed(twiddle_factor_table_35_imag));
  assign _zz_13160 = fixTo_972_dout;
  assign _zz_13161 = ($signed(_zz_1354) - $signed(_zz_1353));
  assign _zz_13162 = ($signed(_zz_1353) + $signed(_zz_1354));
  assign _zz_13163 = _zz_13164[15 : 0];
  assign _zz_13164 = fixTo_974_dout;
  assign _zz_13165 = _zz_13166[15 : 0];
  assign _zz_13166 = fixTo_973_dout;
  assign _zz_13167 = _zz_13168;
  assign _zz_13168 = ($signed(_zz_13169) >>> _zz_3416);
  assign _zz_13169 = _zz_13170;
  assign _zz_13170 = ($signed(_zz_1289) - $signed(_zz_3413));
  assign _zz_13171 = _zz_13172;
  assign _zz_13172 = ($signed(_zz_13173) >>> _zz_3416);
  assign _zz_13173 = _zz_13174;
  assign _zz_13174 = ($signed(_zz_1290) - $signed(_zz_3414));
  assign _zz_13175 = _zz_13176;
  assign _zz_13176 = ($signed(_zz_13177) >>> _zz_3417);
  assign _zz_13177 = _zz_13178;
  assign _zz_13178 = ($signed(_zz_1289) + $signed(_zz_3413));
  assign _zz_13179 = _zz_13180;
  assign _zz_13180 = ($signed(_zz_13181) >>> _zz_3417);
  assign _zz_13181 = _zz_13182;
  assign _zz_13182 = ($signed(_zz_1290) + $signed(_zz_3414));
  assign _zz_13183 = ($signed(twiddle_factor_table_36_real) + $signed(twiddle_factor_table_36_imag));
  assign _zz_13184 = fixTo_975_dout;
  assign _zz_13185 = ($signed(_zz_1356) - $signed(_zz_1355));
  assign _zz_13186 = ($signed(_zz_1355) + $signed(_zz_1356));
  assign _zz_13187 = _zz_13188[15 : 0];
  assign _zz_13188 = fixTo_977_dout;
  assign _zz_13189 = _zz_13190[15 : 0];
  assign _zz_13190 = fixTo_976_dout;
  assign _zz_13191 = _zz_13192;
  assign _zz_13192 = ($signed(_zz_13193) >>> _zz_3421);
  assign _zz_13193 = _zz_13194;
  assign _zz_13194 = ($signed(_zz_1291) - $signed(_zz_3418));
  assign _zz_13195 = _zz_13196;
  assign _zz_13196 = ($signed(_zz_13197) >>> _zz_3421);
  assign _zz_13197 = _zz_13198;
  assign _zz_13198 = ($signed(_zz_1292) - $signed(_zz_3419));
  assign _zz_13199 = _zz_13200;
  assign _zz_13200 = ($signed(_zz_13201) >>> _zz_3422);
  assign _zz_13201 = _zz_13202;
  assign _zz_13202 = ($signed(_zz_1291) + $signed(_zz_3418));
  assign _zz_13203 = _zz_13204;
  assign _zz_13204 = ($signed(_zz_13205) >>> _zz_3422);
  assign _zz_13205 = _zz_13206;
  assign _zz_13206 = ($signed(_zz_1292) + $signed(_zz_3419));
  assign _zz_13207 = ($signed(twiddle_factor_table_37_real) + $signed(twiddle_factor_table_37_imag));
  assign _zz_13208 = fixTo_978_dout;
  assign _zz_13209 = ($signed(_zz_1358) - $signed(_zz_1357));
  assign _zz_13210 = ($signed(_zz_1357) + $signed(_zz_1358));
  assign _zz_13211 = _zz_13212[15 : 0];
  assign _zz_13212 = fixTo_980_dout;
  assign _zz_13213 = _zz_13214[15 : 0];
  assign _zz_13214 = fixTo_979_dout;
  assign _zz_13215 = _zz_13216;
  assign _zz_13216 = ($signed(_zz_13217) >>> _zz_3426);
  assign _zz_13217 = _zz_13218;
  assign _zz_13218 = ($signed(_zz_1293) - $signed(_zz_3423));
  assign _zz_13219 = _zz_13220;
  assign _zz_13220 = ($signed(_zz_13221) >>> _zz_3426);
  assign _zz_13221 = _zz_13222;
  assign _zz_13222 = ($signed(_zz_1294) - $signed(_zz_3424));
  assign _zz_13223 = _zz_13224;
  assign _zz_13224 = ($signed(_zz_13225) >>> _zz_3427);
  assign _zz_13225 = _zz_13226;
  assign _zz_13226 = ($signed(_zz_1293) + $signed(_zz_3423));
  assign _zz_13227 = _zz_13228;
  assign _zz_13228 = ($signed(_zz_13229) >>> _zz_3427);
  assign _zz_13229 = _zz_13230;
  assign _zz_13230 = ($signed(_zz_1294) + $signed(_zz_3424));
  assign _zz_13231 = ($signed(twiddle_factor_table_38_real) + $signed(twiddle_factor_table_38_imag));
  assign _zz_13232 = fixTo_981_dout;
  assign _zz_13233 = ($signed(_zz_1360) - $signed(_zz_1359));
  assign _zz_13234 = ($signed(_zz_1359) + $signed(_zz_1360));
  assign _zz_13235 = _zz_13236[15 : 0];
  assign _zz_13236 = fixTo_983_dout;
  assign _zz_13237 = _zz_13238[15 : 0];
  assign _zz_13238 = fixTo_982_dout;
  assign _zz_13239 = _zz_13240;
  assign _zz_13240 = ($signed(_zz_13241) >>> _zz_3431);
  assign _zz_13241 = _zz_13242;
  assign _zz_13242 = ($signed(_zz_1295) - $signed(_zz_3428));
  assign _zz_13243 = _zz_13244;
  assign _zz_13244 = ($signed(_zz_13245) >>> _zz_3431);
  assign _zz_13245 = _zz_13246;
  assign _zz_13246 = ($signed(_zz_1296) - $signed(_zz_3429));
  assign _zz_13247 = _zz_13248;
  assign _zz_13248 = ($signed(_zz_13249) >>> _zz_3432);
  assign _zz_13249 = _zz_13250;
  assign _zz_13250 = ($signed(_zz_1295) + $signed(_zz_3428));
  assign _zz_13251 = _zz_13252;
  assign _zz_13252 = ($signed(_zz_13253) >>> _zz_3432);
  assign _zz_13253 = _zz_13254;
  assign _zz_13254 = ($signed(_zz_1296) + $signed(_zz_3429));
  assign _zz_13255 = ($signed(twiddle_factor_table_39_real) + $signed(twiddle_factor_table_39_imag));
  assign _zz_13256 = fixTo_984_dout;
  assign _zz_13257 = ($signed(_zz_1362) - $signed(_zz_1361));
  assign _zz_13258 = ($signed(_zz_1361) + $signed(_zz_1362));
  assign _zz_13259 = _zz_13260[15 : 0];
  assign _zz_13260 = fixTo_986_dout;
  assign _zz_13261 = _zz_13262[15 : 0];
  assign _zz_13262 = fixTo_985_dout;
  assign _zz_13263 = _zz_13264;
  assign _zz_13264 = ($signed(_zz_13265) >>> _zz_3436);
  assign _zz_13265 = _zz_13266;
  assign _zz_13266 = ($signed(_zz_1297) - $signed(_zz_3433));
  assign _zz_13267 = _zz_13268;
  assign _zz_13268 = ($signed(_zz_13269) >>> _zz_3436);
  assign _zz_13269 = _zz_13270;
  assign _zz_13270 = ($signed(_zz_1298) - $signed(_zz_3434));
  assign _zz_13271 = _zz_13272;
  assign _zz_13272 = ($signed(_zz_13273) >>> _zz_3437);
  assign _zz_13273 = _zz_13274;
  assign _zz_13274 = ($signed(_zz_1297) + $signed(_zz_3433));
  assign _zz_13275 = _zz_13276;
  assign _zz_13276 = ($signed(_zz_13277) >>> _zz_3437);
  assign _zz_13277 = _zz_13278;
  assign _zz_13278 = ($signed(_zz_1298) + $signed(_zz_3434));
  assign _zz_13279 = ($signed(twiddle_factor_table_40_real) + $signed(twiddle_factor_table_40_imag));
  assign _zz_13280 = fixTo_987_dout;
  assign _zz_13281 = ($signed(_zz_1364) - $signed(_zz_1363));
  assign _zz_13282 = ($signed(_zz_1363) + $signed(_zz_1364));
  assign _zz_13283 = _zz_13284[15 : 0];
  assign _zz_13284 = fixTo_989_dout;
  assign _zz_13285 = _zz_13286[15 : 0];
  assign _zz_13286 = fixTo_988_dout;
  assign _zz_13287 = _zz_13288;
  assign _zz_13288 = ($signed(_zz_13289) >>> _zz_3441);
  assign _zz_13289 = _zz_13290;
  assign _zz_13290 = ($signed(_zz_1299) - $signed(_zz_3438));
  assign _zz_13291 = _zz_13292;
  assign _zz_13292 = ($signed(_zz_13293) >>> _zz_3441);
  assign _zz_13293 = _zz_13294;
  assign _zz_13294 = ($signed(_zz_1300) - $signed(_zz_3439));
  assign _zz_13295 = _zz_13296;
  assign _zz_13296 = ($signed(_zz_13297) >>> _zz_3442);
  assign _zz_13297 = _zz_13298;
  assign _zz_13298 = ($signed(_zz_1299) + $signed(_zz_3438));
  assign _zz_13299 = _zz_13300;
  assign _zz_13300 = ($signed(_zz_13301) >>> _zz_3442);
  assign _zz_13301 = _zz_13302;
  assign _zz_13302 = ($signed(_zz_1300) + $signed(_zz_3439));
  assign _zz_13303 = ($signed(twiddle_factor_table_41_real) + $signed(twiddle_factor_table_41_imag));
  assign _zz_13304 = fixTo_990_dout;
  assign _zz_13305 = ($signed(_zz_1366) - $signed(_zz_1365));
  assign _zz_13306 = ($signed(_zz_1365) + $signed(_zz_1366));
  assign _zz_13307 = _zz_13308[15 : 0];
  assign _zz_13308 = fixTo_992_dout;
  assign _zz_13309 = _zz_13310[15 : 0];
  assign _zz_13310 = fixTo_991_dout;
  assign _zz_13311 = _zz_13312;
  assign _zz_13312 = ($signed(_zz_13313) >>> _zz_3446);
  assign _zz_13313 = _zz_13314;
  assign _zz_13314 = ($signed(_zz_1301) - $signed(_zz_3443));
  assign _zz_13315 = _zz_13316;
  assign _zz_13316 = ($signed(_zz_13317) >>> _zz_3446);
  assign _zz_13317 = _zz_13318;
  assign _zz_13318 = ($signed(_zz_1302) - $signed(_zz_3444));
  assign _zz_13319 = _zz_13320;
  assign _zz_13320 = ($signed(_zz_13321) >>> _zz_3447);
  assign _zz_13321 = _zz_13322;
  assign _zz_13322 = ($signed(_zz_1301) + $signed(_zz_3443));
  assign _zz_13323 = _zz_13324;
  assign _zz_13324 = ($signed(_zz_13325) >>> _zz_3447);
  assign _zz_13325 = _zz_13326;
  assign _zz_13326 = ($signed(_zz_1302) + $signed(_zz_3444));
  assign _zz_13327 = ($signed(twiddle_factor_table_42_real) + $signed(twiddle_factor_table_42_imag));
  assign _zz_13328 = fixTo_993_dout;
  assign _zz_13329 = ($signed(_zz_1368) - $signed(_zz_1367));
  assign _zz_13330 = ($signed(_zz_1367) + $signed(_zz_1368));
  assign _zz_13331 = _zz_13332[15 : 0];
  assign _zz_13332 = fixTo_995_dout;
  assign _zz_13333 = _zz_13334[15 : 0];
  assign _zz_13334 = fixTo_994_dout;
  assign _zz_13335 = _zz_13336;
  assign _zz_13336 = ($signed(_zz_13337) >>> _zz_3451);
  assign _zz_13337 = _zz_13338;
  assign _zz_13338 = ($signed(_zz_1303) - $signed(_zz_3448));
  assign _zz_13339 = _zz_13340;
  assign _zz_13340 = ($signed(_zz_13341) >>> _zz_3451);
  assign _zz_13341 = _zz_13342;
  assign _zz_13342 = ($signed(_zz_1304) - $signed(_zz_3449));
  assign _zz_13343 = _zz_13344;
  assign _zz_13344 = ($signed(_zz_13345) >>> _zz_3452);
  assign _zz_13345 = _zz_13346;
  assign _zz_13346 = ($signed(_zz_1303) + $signed(_zz_3448));
  assign _zz_13347 = _zz_13348;
  assign _zz_13348 = ($signed(_zz_13349) >>> _zz_3452);
  assign _zz_13349 = _zz_13350;
  assign _zz_13350 = ($signed(_zz_1304) + $signed(_zz_3449));
  assign _zz_13351 = ($signed(twiddle_factor_table_43_real) + $signed(twiddle_factor_table_43_imag));
  assign _zz_13352 = fixTo_996_dout;
  assign _zz_13353 = ($signed(_zz_1370) - $signed(_zz_1369));
  assign _zz_13354 = ($signed(_zz_1369) + $signed(_zz_1370));
  assign _zz_13355 = _zz_13356[15 : 0];
  assign _zz_13356 = fixTo_998_dout;
  assign _zz_13357 = _zz_13358[15 : 0];
  assign _zz_13358 = fixTo_997_dout;
  assign _zz_13359 = _zz_13360;
  assign _zz_13360 = ($signed(_zz_13361) >>> _zz_3456);
  assign _zz_13361 = _zz_13362;
  assign _zz_13362 = ($signed(_zz_1305) - $signed(_zz_3453));
  assign _zz_13363 = _zz_13364;
  assign _zz_13364 = ($signed(_zz_13365) >>> _zz_3456);
  assign _zz_13365 = _zz_13366;
  assign _zz_13366 = ($signed(_zz_1306) - $signed(_zz_3454));
  assign _zz_13367 = _zz_13368;
  assign _zz_13368 = ($signed(_zz_13369) >>> _zz_3457);
  assign _zz_13369 = _zz_13370;
  assign _zz_13370 = ($signed(_zz_1305) + $signed(_zz_3453));
  assign _zz_13371 = _zz_13372;
  assign _zz_13372 = ($signed(_zz_13373) >>> _zz_3457);
  assign _zz_13373 = _zz_13374;
  assign _zz_13374 = ($signed(_zz_1306) + $signed(_zz_3454));
  assign _zz_13375 = ($signed(twiddle_factor_table_44_real) + $signed(twiddle_factor_table_44_imag));
  assign _zz_13376 = fixTo_999_dout;
  assign _zz_13377 = ($signed(_zz_1372) - $signed(_zz_1371));
  assign _zz_13378 = ($signed(_zz_1371) + $signed(_zz_1372));
  assign _zz_13379 = _zz_13380[15 : 0];
  assign _zz_13380 = fixTo_1001_dout;
  assign _zz_13381 = _zz_13382[15 : 0];
  assign _zz_13382 = fixTo_1000_dout;
  assign _zz_13383 = _zz_13384;
  assign _zz_13384 = ($signed(_zz_13385) >>> _zz_3461);
  assign _zz_13385 = _zz_13386;
  assign _zz_13386 = ($signed(_zz_1307) - $signed(_zz_3458));
  assign _zz_13387 = _zz_13388;
  assign _zz_13388 = ($signed(_zz_13389) >>> _zz_3461);
  assign _zz_13389 = _zz_13390;
  assign _zz_13390 = ($signed(_zz_1308) - $signed(_zz_3459));
  assign _zz_13391 = _zz_13392;
  assign _zz_13392 = ($signed(_zz_13393) >>> _zz_3462);
  assign _zz_13393 = _zz_13394;
  assign _zz_13394 = ($signed(_zz_1307) + $signed(_zz_3458));
  assign _zz_13395 = _zz_13396;
  assign _zz_13396 = ($signed(_zz_13397) >>> _zz_3462);
  assign _zz_13397 = _zz_13398;
  assign _zz_13398 = ($signed(_zz_1308) + $signed(_zz_3459));
  assign _zz_13399 = ($signed(twiddle_factor_table_45_real) + $signed(twiddle_factor_table_45_imag));
  assign _zz_13400 = fixTo_1002_dout;
  assign _zz_13401 = ($signed(_zz_1374) - $signed(_zz_1373));
  assign _zz_13402 = ($signed(_zz_1373) + $signed(_zz_1374));
  assign _zz_13403 = _zz_13404[15 : 0];
  assign _zz_13404 = fixTo_1004_dout;
  assign _zz_13405 = _zz_13406[15 : 0];
  assign _zz_13406 = fixTo_1003_dout;
  assign _zz_13407 = _zz_13408;
  assign _zz_13408 = ($signed(_zz_13409) >>> _zz_3466);
  assign _zz_13409 = _zz_13410;
  assign _zz_13410 = ($signed(_zz_1309) - $signed(_zz_3463));
  assign _zz_13411 = _zz_13412;
  assign _zz_13412 = ($signed(_zz_13413) >>> _zz_3466);
  assign _zz_13413 = _zz_13414;
  assign _zz_13414 = ($signed(_zz_1310) - $signed(_zz_3464));
  assign _zz_13415 = _zz_13416;
  assign _zz_13416 = ($signed(_zz_13417) >>> _zz_3467);
  assign _zz_13417 = _zz_13418;
  assign _zz_13418 = ($signed(_zz_1309) + $signed(_zz_3463));
  assign _zz_13419 = _zz_13420;
  assign _zz_13420 = ($signed(_zz_13421) >>> _zz_3467);
  assign _zz_13421 = _zz_13422;
  assign _zz_13422 = ($signed(_zz_1310) + $signed(_zz_3464));
  assign _zz_13423 = ($signed(twiddle_factor_table_46_real) + $signed(twiddle_factor_table_46_imag));
  assign _zz_13424 = fixTo_1005_dout;
  assign _zz_13425 = ($signed(_zz_1376) - $signed(_zz_1375));
  assign _zz_13426 = ($signed(_zz_1375) + $signed(_zz_1376));
  assign _zz_13427 = _zz_13428[15 : 0];
  assign _zz_13428 = fixTo_1007_dout;
  assign _zz_13429 = _zz_13430[15 : 0];
  assign _zz_13430 = fixTo_1006_dout;
  assign _zz_13431 = _zz_13432;
  assign _zz_13432 = ($signed(_zz_13433) >>> _zz_3471);
  assign _zz_13433 = _zz_13434;
  assign _zz_13434 = ($signed(_zz_1311) - $signed(_zz_3468));
  assign _zz_13435 = _zz_13436;
  assign _zz_13436 = ($signed(_zz_13437) >>> _zz_3471);
  assign _zz_13437 = _zz_13438;
  assign _zz_13438 = ($signed(_zz_1312) - $signed(_zz_3469));
  assign _zz_13439 = _zz_13440;
  assign _zz_13440 = ($signed(_zz_13441) >>> _zz_3472);
  assign _zz_13441 = _zz_13442;
  assign _zz_13442 = ($signed(_zz_1311) + $signed(_zz_3468));
  assign _zz_13443 = _zz_13444;
  assign _zz_13444 = ($signed(_zz_13445) >>> _zz_3472);
  assign _zz_13445 = _zz_13446;
  assign _zz_13446 = ($signed(_zz_1312) + $signed(_zz_3469));
  assign _zz_13447 = ($signed(twiddle_factor_table_47_real) + $signed(twiddle_factor_table_47_imag));
  assign _zz_13448 = fixTo_1008_dout;
  assign _zz_13449 = ($signed(_zz_1378) - $signed(_zz_1377));
  assign _zz_13450 = ($signed(_zz_1377) + $signed(_zz_1378));
  assign _zz_13451 = _zz_13452[15 : 0];
  assign _zz_13452 = fixTo_1010_dout;
  assign _zz_13453 = _zz_13454[15 : 0];
  assign _zz_13454 = fixTo_1009_dout;
  assign _zz_13455 = _zz_13456;
  assign _zz_13456 = ($signed(_zz_13457) >>> _zz_3476);
  assign _zz_13457 = _zz_13458;
  assign _zz_13458 = ($signed(_zz_1313) - $signed(_zz_3473));
  assign _zz_13459 = _zz_13460;
  assign _zz_13460 = ($signed(_zz_13461) >>> _zz_3476);
  assign _zz_13461 = _zz_13462;
  assign _zz_13462 = ($signed(_zz_1314) - $signed(_zz_3474));
  assign _zz_13463 = _zz_13464;
  assign _zz_13464 = ($signed(_zz_13465) >>> _zz_3477);
  assign _zz_13465 = _zz_13466;
  assign _zz_13466 = ($signed(_zz_1313) + $signed(_zz_3473));
  assign _zz_13467 = _zz_13468;
  assign _zz_13468 = ($signed(_zz_13469) >>> _zz_3477);
  assign _zz_13469 = _zz_13470;
  assign _zz_13470 = ($signed(_zz_1314) + $signed(_zz_3474));
  assign _zz_13471 = ($signed(twiddle_factor_table_48_real) + $signed(twiddle_factor_table_48_imag));
  assign _zz_13472 = fixTo_1011_dout;
  assign _zz_13473 = ($signed(_zz_1380) - $signed(_zz_1379));
  assign _zz_13474 = ($signed(_zz_1379) + $signed(_zz_1380));
  assign _zz_13475 = _zz_13476[15 : 0];
  assign _zz_13476 = fixTo_1013_dout;
  assign _zz_13477 = _zz_13478[15 : 0];
  assign _zz_13478 = fixTo_1012_dout;
  assign _zz_13479 = _zz_13480;
  assign _zz_13480 = ($signed(_zz_13481) >>> _zz_3481);
  assign _zz_13481 = _zz_13482;
  assign _zz_13482 = ($signed(_zz_1315) - $signed(_zz_3478));
  assign _zz_13483 = _zz_13484;
  assign _zz_13484 = ($signed(_zz_13485) >>> _zz_3481);
  assign _zz_13485 = _zz_13486;
  assign _zz_13486 = ($signed(_zz_1316) - $signed(_zz_3479));
  assign _zz_13487 = _zz_13488;
  assign _zz_13488 = ($signed(_zz_13489) >>> _zz_3482);
  assign _zz_13489 = _zz_13490;
  assign _zz_13490 = ($signed(_zz_1315) + $signed(_zz_3478));
  assign _zz_13491 = _zz_13492;
  assign _zz_13492 = ($signed(_zz_13493) >>> _zz_3482);
  assign _zz_13493 = _zz_13494;
  assign _zz_13494 = ($signed(_zz_1316) + $signed(_zz_3479));
  assign _zz_13495 = ($signed(twiddle_factor_table_49_real) + $signed(twiddle_factor_table_49_imag));
  assign _zz_13496 = fixTo_1014_dout;
  assign _zz_13497 = ($signed(_zz_1382) - $signed(_zz_1381));
  assign _zz_13498 = ($signed(_zz_1381) + $signed(_zz_1382));
  assign _zz_13499 = _zz_13500[15 : 0];
  assign _zz_13500 = fixTo_1016_dout;
  assign _zz_13501 = _zz_13502[15 : 0];
  assign _zz_13502 = fixTo_1015_dout;
  assign _zz_13503 = _zz_13504;
  assign _zz_13504 = ($signed(_zz_13505) >>> _zz_3486);
  assign _zz_13505 = _zz_13506;
  assign _zz_13506 = ($signed(_zz_1317) - $signed(_zz_3483));
  assign _zz_13507 = _zz_13508;
  assign _zz_13508 = ($signed(_zz_13509) >>> _zz_3486);
  assign _zz_13509 = _zz_13510;
  assign _zz_13510 = ($signed(_zz_1318) - $signed(_zz_3484));
  assign _zz_13511 = _zz_13512;
  assign _zz_13512 = ($signed(_zz_13513) >>> _zz_3487);
  assign _zz_13513 = _zz_13514;
  assign _zz_13514 = ($signed(_zz_1317) + $signed(_zz_3483));
  assign _zz_13515 = _zz_13516;
  assign _zz_13516 = ($signed(_zz_13517) >>> _zz_3487);
  assign _zz_13517 = _zz_13518;
  assign _zz_13518 = ($signed(_zz_1318) + $signed(_zz_3484));
  assign _zz_13519 = ($signed(twiddle_factor_table_50_real) + $signed(twiddle_factor_table_50_imag));
  assign _zz_13520 = fixTo_1017_dout;
  assign _zz_13521 = ($signed(_zz_1384) - $signed(_zz_1383));
  assign _zz_13522 = ($signed(_zz_1383) + $signed(_zz_1384));
  assign _zz_13523 = _zz_13524[15 : 0];
  assign _zz_13524 = fixTo_1019_dout;
  assign _zz_13525 = _zz_13526[15 : 0];
  assign _zz_13526 = fixTo_1018_dout;
  assign _zz_13527 = _zz_13528;
  assign _zz_13528 = ($signed(_zz_13529) >>> _zz_3491);
  assign _zz_13529 = _zz_13530;
  assign _zz_13530 = ($signed(_zz_1319) - $signed(_zz_3488));
  assign _zz_13531 = _zz_13532;
  assign _zz_13532 = ($signed(_zz_13533) >>> _zz_3491);
  assign _zz_13533 = _zz_13534;
  assign _zz_13534 = ($signed(_zz_1320) - $signed(_zz_3489));
  assign _zz_13535 = _zz_13536;
  assign _zz_13536 = ($signed(_zz_13537) >>> _zz_3492);
  assign _zz_13537 = _zz_13538;
  assign _zz_13538 = ($signed(_zz_1319) + $signed(_zz_3488));
  assign _zz_13539 = _zz_13540;
  assign _zz_13540 = ($signed(_zz_13541) >>> _zz_3492);
  assign _zz_13541 = _zz_13542;
  assign _zz_13542 = ($signed(_zz_1320) + $signed(_zz_3489));
  assign _zz_13543 = ($signed(twiddle_factor_table_51_real) + $signed(twiddle_factor_table_51_imag));
  assign _zz_13544 = fixTo_1020_dout;
  assign _zz_13545 = ($signed(_zz_1386) - $signed(_zz_1385));
  assign _zz_13546 = ($signed(_zz_1385) + $signed(_zz_1386));
  assign _zz_13547 = _zz_13548[15 : 0];
  assign _zz_13548 = fixTo_1022_dout;
  assign _zz_13549 = _zz_13550[15 : 0];
  assign _zz_13550 = fixTo_1021_dout;
  assign _zz_13551 = _zz_13552;
  assign _zz_13552 = ($signed(_zz_13553) >>> _zz_3496);
  assign _zz_13553 = _zz_13554;
  assign _zz_13554 = ($signed(_zz_1321) - $signed(_zz_3493));
  assign _zz_13555 = _zz_13556;
  assign _zz_13556 = ($signed(_zz_13557) >>> _zz_3496);
  assign _zz_13557 = _zz_13558;
  assign _zz_13558 = ($signed(_zz_1322) - $signed(_zz_3494));
  assign _zz_13559 = _zz_13560;
  assign _zz_13560 = ($signed(_zz_13561) >>> _zz_3497);
  assign _zz_13561 = _zz_13562;
  assign _zz_13562 = ($signed(_zz_1321) + $signed(_zz_3493));
  assign _zz_13563 = _zz_13564;
  assign _zz_13564 = ($signed(_zz_13565) >>> _zz_3497);
  assign _zz_13565 = _zz_13566;
  assign _zz_13566 = ($signed(_zz_1322) + $signed(_zz_3494));
  assign _zz_13567 = ($signed(twiddle_factor_table_52_real) + $signed(twiddle_factor_table_52_imag));
  assign _zz_13568 = fixTo_1023_dout;
  assign _zz_13569 = ($signed(_zz_1388) - $signed(_zz_1387));
  assign _zz_13570 = ($signed(_zz_1387) + $signed(_zz_1388));
  assign _zz_13571 = _zz_13572[15 : 0];
  assign _zz_13572 = fixTo_1025_dout;
  assign _zz_13573 = _zz_13574[15 : 0];
  assign _zz_13574 = fixTo_1024_dout;
  assign _zz_13575 = _zz_13576;
  assign _zz_13576 = ($signed(_zz_13577) >>> _zz_3501);
  assign _zz_13577 = _zz_13578;
  assign _zz_13578 = ($signed(_zz_1323) - $signed(_zz_3498));
  assign _zz_13579 = _zz_13580;
  assign _zz_13580 = ($signed(_zz_13581) >>> _zz_3501);
  assign _zz_13581 = _zz_13582;
  assign _zz_13582 = ($signed(_zz_1324) - $signed(_zz_3499));
  assign _zz_13583 = _zz_13584;
  assign _zz_13584 = ($signed(_zz_13585) >>> _zz_3502);
  assign _zz_13585 = _zz_13586;
  assign _zz_13586 = ($signed(_zz_1323) + $signed(_zz_3498));
  assign _zz_13587 = _zz_13588;
  assign _zz_13588 = ($signed(_zz_13589) >>> _zz_3502);
  assign _zz_13589 = _zz_13590;
  assign _zz_13590 = ($signed(_zz_1324) + $signed(_zz_3499));
  assign _zz_13591 = ($signed(twiddle_factor_table_53_real) + $signed(twiddle_factor_table_53_imag));
  assign _zz_13592 = fixTo_1026_dout;
  assign _zz_13593 = ($signed(_zz_1390) - $signed(_zz_1389));
  assign _zz_13594 = ($signed(_zz_1389) + $signed(_zz_1390));
  assign _zz_13595 = _zz_13596[15 : 0];
  assign _zz_13596 = fixTo_1028_dout;
  assign _zz_13597 = _zz_13598[15 : 0];
  assign _zz_13598 = fixTo_1027_dout;
  assign _zz_13599 = _zz_13600;
  assign _zz_13600 = ($signed(_zz_13601) >>> _zz_3506);
  assign _zz_13601 = _zz_13602;
  assign _zz_13602 = ($signed(_zz_1325) - $signed(_zz_3503));
  assign _zz_13603 = _zz_13604;
  assign _zz_13604 = ($signed(_zz_13605) >>> _zz_3506);
  assign _zz_13605 = _zz_13606;
  assign _zz_13606 = ($signed(_zz_1326) - $signed(_zz_3504));
  assign _zz_13607 = _zz_13608;
  assign _zz_13608 = ($signed(_zz_13609) >>> _zz_3507);
  assign _zz_13609 = _zz_13610;
  assign _zz_13610 = ($signed(_zz_1325) + $signed(_zz_3503));
  assign _zz_13611 = _zz_13612;
  assign _zz_13612 = ($signed(_zz_13613) >>> _zz_3507);
  assign _zz_13613 = _zz_13614;
  assign _zz_13614 = ($signed(_zz_1326) + $signed(_zz_3504));
  assign _zz_13615 = ($signed(twiddle_factor_table_54_real) + $signed(twiddle_factor_table_54_imag));
  assign _zz_13616 = fixTo_1029_dout;
  assign _zz_13617 = ($signed(_zz_1392) - $signed(_zz_1391));
  assign _zz_13618 = ($signed(_zz_1391) + $signed(_zz_1392));
  assign _zz_13619 = _zz_13620[15 : 0];
  assign _zz_13620 = fixTo_1031_dout;
  assign _zz_13621 = _zz_13622[15 : 0];
  assign _zz_13622 = fixTo_1030_dout;
  assign _zz_13623 = _zz_13624;
  assign _zz_13624 = ($signed(_zz_13625) >>> _zz_3511);
  assign _zz_13625 = _zz_13626;
  assign _zz_13626 = ($signed(_zz_1327) - $signed(_zz_3508));
  assign _zz_13627 = _zz_13628;
  assign _zz_13628 = ($signed(_zz_13629) >>> _zz_3511);
  assign _zz_13629 = _zz_13630;
  assign _zz_13630 = ($signed(_zz_1328) - $signed(_zz_3509));
  assign _zz_13631 = _zz_13632;
  assign _zz_13632 = ($signed(_zz_13633) >>> _zz_3512);
  assign _zz_13633 = _zz_13634;
  assign _zz_13634 = ($signed(_zz_1327) + $signed(_zz_3508));
  assign _zz_13635 = _zz_13636;
  assign _zz_13636 = ($signed(_zz_13637) >>> _zz_3512);
  assign _zz_13637 = _zz_13638;
  assign _zz_13638 = ($signed(_zz_1328) + $signed(_zz_3509));
  assign _zz_13639 = ($signed(twiddle_factor_table_55_real) + $signed(twiddle_factor_table_55_imag));
  assign _zz_13640 = fixTo_1032_dout;
  assign _zz_13641 = ($signed(_zz_1394) - $signed(_zz_1393));
  assign _zz_13642 = ($signed(_zz_1393) + $signed(_zz_1394));
  assign _zz_13643 = _zz_13644[15 : 0];
  assign _zz_13644 = fixTo_1034_dout;
  assign _zz_13645 = _zz_13646[15 : 0];
  assign _zz_13646 = fixTo_1033_dout;
  assign _zz_13647 = _zz_13648;
  assign _zz_13648 = ($signed(_zz_13649) >>> _zz_3516);
  assign _zz_13649 = _zz_13650;
  assign _zz_13650 = ($signed(_zz_1329) - $signed(_zz_3513));
  assign _zz_13651 = _zz_13652;
  assign _zz_13652 = ($signed(_zz_13653) >>> _zz_3516);
  assign _zz_13653 = _zz_13654;
  assign _zz_13654 = ($signed(_zz_1330) - $signed(_zz_3514));
  assign _zz_13655 = _zz_13656;
  assign _zz_13656 = ($signed(_zz_13657) >>> _zz_3517);
  assign _zz_13657 = _zz_13658;
  assign _zz_13658 = ($signed(_zz_1329) + $signed(_zz_3513));
  assign _zz_13659 = _zz_13660;
  assign _zz_13660 = ($signed(_zz_13661) >>> _zz_3517);
  assign _zz_13661 = _zz_13662;
  assign _zz_13662 = ($signed(_zz_1330) + $signed(_zz_3514));
  assign _zz_13663 = ($signed(twiddle_factor_table_56_real) + $signed(twiddle_factor_table_56_imag));
  assign _zz_13664 = fixTo_1035_dout;
  assign _zz_13665 = ($signed(_zz_1396) - $signed(_zz_1395));
  assign _zz_13666 = ($signed(_zz_1395) + $signed(_zz_1396));
  assign _zz_13667 = _zz_13668[15 : 0];
  assign _zz_13668 = fixTo_1037_dout;
  assign _zz_13669 = _zz_13670[15 : 0];
  assign _zz_13670 = fixTo_1036_dout;
  assign _zz_13671 = _zz_13672;
  assign _zz_13672 = ($signed(_zz_13673) >>> _zz_3521);
  assign _zz_13673 = _zz_13674;
  assign _zz_13674 = ($signed(_zz_1331) - $signed(_zz_3518));
  assign _zz_13675 = _zz_13676;
  assign _zz_13676 = ($signed(_zz_13677) >>> _zz_3521);
  assign _zz_13677 = _zz_13678;
  assign _zz_13678 = ($signed(_zz_1332) - $signed(_zz_3519));
  assign _zz_13679 = _zz_13680;
  assign _zz_13680 = ($signed(_zz_13681) >>> _zz_3522);
  assign _zz_13681 = _zz_13682;
  assign _zz_13682 = ($signed(_zz_1331) + $signed(_zz_3518));
  assign _zz_13683 = _zz_13684;
  assign _zz_13684 = ($signed(_zz_13685) >>> _zz_3522);
  assign _zz_13685 = _zz_13686;
  assign _zz_13686 = ($signed(_zz_1332) + $signed(_zz_3519));
  assign _zz_13687 = ($signed(twiddle_factor_table_57_real) + $signed(twiddle_factor_table_57_imag));
  assign _zz_13688 = fixTo_1038_dout;
  assign _zz_13689 = ($signed(_zz_1398) - $signed(_zz_1397));
  assign _zz_13690 = ($signed(_zz_1397) + $signed(_zz_1398));
  assign _zz_13691 = _zz_13692[15 : 0];
  assign _zz_13692 = fixTo_1040_dout;
  assign _zz_13693 = _zz_13694[15 : 0];
  assign _zz_13694 = fixTo_1039_dout;
  assign _zz_13695 = _zz_13696;
  assign _zz_13696 = ($signed(_zz_13697) >>> _zz_3526);
  assign _zz_13697 = _zz_13698;
  assign _zz_13698 = ($signed(_zz_1333) - $signed(_zz_3523));
  assign _zz_13699 = _zz_13700;
  assign _zz_13700 = ($signed(_zz_13701) >>> _zz_3526);
  assign _zz_13701 = _zz_13702;
  assign _zz_13702 = ($signed(_zz_1334) - $signed(_zz_3524));
  assign _zz_13703 = _zz_13704;
  assign _zz_13704 = ($signed(_zz_13705) >>> _zz_3527);
  assign _zz_13705 = _zz_13706;
  assign _zz_13706 = ($signed(_zz_1333) + $signed(_zz_3523));
  assign _zz_13707 = _zz_13708;
  assign _zz_13708 = ($signed(_zz_13709) >>> _zz_3527);
  assign _zz_13709 = _zz_13710;
  assign _zz_13710 = ($signed(_zz_1334) + $signed(_zz_3524));
  assign _zz_13711 = ($signed(twiddle_factor_table_58_real) + $signed(twiddle_factor_table_58_imag));
  assign _zz_13712 = fixTo_1041_dout;
  assign _zz_13713 = ($signed(_zz_1400) - $signed(_zz_1399));
  assign _zz_13714 = ($signed(_zz_1399) + $signed(_zz_1400));
  assign _zz_13715 = _zz_13716[15 : 0];
  assign _zz_13716 = fixTo_1043_dout;
  assign _zz_13717 = _zz_13718[15 : 0];
  assign _zz_13718 = fixTo_1042_dout;
  assign _zz_13719 = _zz_13720;
  assign _zz_13720 = ($signed(_zz_13721) >>> _zz_3531);
  assign _zz_13721 = _zz_13722;
  assign _zz_13722 = ($signed(_zz_1335) - $signed(_zz_3528));
  assign _zz_13723 = _zz_13724;
  assign _zz_13724 = ($signed(_zz_13725) >>> _zz_3531);
  assign _zz_13725 = _zz_13726;
  assign _zz_13726 = ($signed(_zz_1336) - $signed(_zz_3529));
  assign _zz_13727 = _zz_13728;
  assign _zz_13728 = ($signed(_zz_13729) >>> _zz_3532);
  assign _zz_13729 = _zz_13730;
  assign _zz_13730 = ($signed(_zz_1335) + $signed(_zz_3528));
  assign _zz_13731 = _zz_13732;
  assign _zz_13732 = ($signed(_zz_13733) >>> _zz_3532);
  assign _zz_13733 = _zz_13734;
  assign _zz_13734 = ($signed(_zz_1336) + $signed(_zz_3529));
  assign _zz_13735 = ($signed(twiddle_factor_table_59_real) + $signed(twiddle_factor_table_59_imag));
  assign _zz_13736 = fixTo_1044_dout;
  assign _zz_13737 = ($signed(_zz_1402) - $signed(_zz_1401));
  assign _zz_13738 = ($signed(_zz_1401) + $signed(_zz_1402));
  assign _zz_13739 = _zz_13740[15 : 0];
  assign _zz_13740 = fixTo_1046_dout;
  assign _zz_13741 = _zz_13742[15 : 0];
  assign _zz_13742 = fixTo_1045_dout;
  assign _zz_13743 = _zz_13744;
  assign _zz_13744 = ($signed(_zz_13745) >>> _zz_3536);
  assign _zz_13745 = _zz_13746;
  assign _zz_13746 = ($signed(_zz_1337) - $signed(_zz_3533));
  assign _zz_13747 = _zz_13748;
  assign _zz_13748 = ($signed(_zz_13749) >>> _zz_3536);
  assign _zz_13749 = _zz_13750;
  assign _zz_13750 = ($signed(_zz_1338) - $signed(_zz_3534));
  assign _zz_13751 = _zz_13752;
  assign _zz_13752 = ($signed(_zz_13753) >>> _zz_3537);
  assign _zz_13753 = _zz_13754;
  assign _zz_13754 = ($signed(_zz_1337) + $signed(_zz_3533));
  assign _zz_13755 = _zz_13756;
  assign _zz_13756 = ($signed(_zz_13757) >>> _zz_3537);
  assign _zz_13757 = _zz_13758;
  assign _zz_13758 = ($signed(_zz_1338) + $signed(_zz_3534));
  assign _zz_13759 = ($signed(twiddle_factor_table_60_real) + $signed(twiddle_factor_table_60_imag));
  assign _zz_13760 = fixTo_1047_dout;
  assign _zz_13761 = ($signed(_zz_1404) - $signed(_zz_1403));
  assign _zz_13762 = ($signed(_zz_1403) + $signed(_zz_1404));
  assign _zz_13763 = _zz_13764[15 : 0];
  assign _zz_13764 = fixTo_1049_dout;
  assign _zz_13765 = _zz_13766[15 : 0];
  assign _zz_13766 = fixTo_1048_dout;
  assign _zz_13767 = _zz_13768;
  assign _zz_13768 = ($signed(_zz_13769) >>> _zz_3541);
  assign _zz_13769 = _zz_13770;
  assign _zz_13770 = ($signed(_zz_1339) - $signed(_zz_3538));
  assign _zz_13771 = _zz_13772;
  assign _zz_13772 = ($signed(_zz_13773) >>> _zz_3541);
  assign _zz_13773 = _zz_13774;
  assign _zz_13774 = ($signed(_zz_1340) - $signed(_zz_3539));
  assign _zz_13775 = _zz_13776;
  assign _zz_13776 = ($signed(_zz_13777) >>> _zz_3542);
  assign _zz_13777 = _zz_13778;
  assign _zz_13778 = ($signed(_zz_1339) + $signed(_zz_3538));
  assign _zz_13779 = _zz_13780;
  assign _zz_13780 = ($signed(_zz_13781) >>> _zz_3542);
  assign _zz_13781 = _zz_13782;
  assign _zz_13782 = ($signed(_zz_1340) + $signed(_zz_3539));
  assign _zz_13783 = ($signed(twiddle_factor_table_61_real) + $signed(twiddle_factor_table_61_imag));
  assign _zz_13784 = fixTo_1050_dout;
  assign _zz_13785 = ($signed(_zz_1406) - $signed(_zz_1405));
  assign _zz_13786 = ($signed(_zz_1405) + $signed(_zz_1406));
  assign _zz_13787 = _zz_13788[15 : 0];
  assign _zz_13788 = fixTo_1052_dout;
  assign _zz_13789 = _zz_13790[15 : 0];
  assign _zz_13790 = fixTo_1051_dout;
  assign _zz_13791 = _zz_13792;
  assign _zz_13792 = ($signed(_zz_13793) >>> _zz_3546);
  assign _zz_13793 = _zz_13794;
  assign _zz_13794 = ($signed(_zz_1341) - $signed(_zz_3543));
  assign _zz_13795 = _zz_13796;
  assign _zz_13796 = ($signed(_zz_13797) >>> _zz_3546);
  assign _zz_13797 = _zz_13798;
  assign _zz_13798 = ($signed(_zz_1342) - $signed(_zz_3544));
  assign _zz_13799 = _zz_13800;
  assign _zz_13800 = ($signed(_zz_13801) >>> _zz_3547);
  assign _zz_13801 = _zz_13802;
  assign _zz_13802 = ($signed(_zz_1341) + $signed(_zz_3543));
  assign _zz_13803 = _zz_13804;
  assign _zz_13804 = ($signed(_zz_13805) >>> _zz_3547);
  assign _zz_13805 = _zz_13806;
  assign _zz_13806 = ($signed(_zz_1342) + $signed(_zz_3544));
  assign _zz_13807 = ($signed(twiddle_factor_table_62_real) + $signed(twiddle_factor_table_62_imag));
  assign _zz_13808 = fixTo_1053_dout;
  assign _zz_13809 = ($signed(_zz_1408) - $signed(_zz_1407));
  assign _zz_13810 = ($signed(_zz_1407) + $signed(_zz_1408));
  assign _zz_13811 = _zz_13812[15 : 0];
  assign _zz_13812 = fixTo_1055_dout;
  assign _zz_13813 = _zz_13814[15 : 0];
  assign _zz_13814 = fixTo_1054_dout;
  assign _zz_13815 = _zz_13816;
  assign _zz_13816 = ($signed(_zz_13817) >>> _zz_3551);
  assign _zz_13817 = _zz_13818;
  assign _zz_13818 = ($signed(_zz_1343) - $signed(_zz_3548));
  assign _zz_13819 = _zz_13820;
  assign _zz_13820 = ($signed(_zz_13821) >>> _zz_3551);
  assign _zz_13821 = _zz_13822;
  assign _zz_13822 = ($signed(_zz_1344) - $signed(_zz_3549));
  assign _zz_13823 = _zz_13824;
  assign _zz_13824 = ($signed(_zz_13825) >>> _zz_3552);
  assign _zz_13825 = _zz_13826;
  assign _zz_13826 = ($signed(_zz_1343) + $signed(_zz_3548));
  assign _zz_13827 = _zz_13828;
  assign _zz_13828 = ($signed(_zz_13829) >>> _zz_3552);
  assign _zz_13829 = _zz_13830;
  assign _zz_13830 = ($signed(_zz_1344) + $signed(_zz_3549));
  assign _zz_13831 = ($signed(twiddle_factor_table_31_real) + $signed(twiddle_factor_table_31_imag));
  assign _zz_13832 = fixTo_1056_dout;
  assign _zz_13833 = ($signed(_zz_1474) - $signed(_zz_1473));
  assign _zz_13834 = ($signed(_zz_1473) + $signed(_zz_1474));
  assign _zz_13835 = _zz_13836[15 : 0];
  assign _zz_13836 = fixTo_1058_dout;
  assign _zz_13837 = _zz_13838[15 : 0];
  assign _zz_13838 = fixTo_1057_dout;
  assign _zz_13839 = _zz_13840;
  assign _zz_13840 = ($signed(_zz_13841) >>> _zz_3556);
  assign _zz_13841 = _zz_13842;
  assign _zz_13842 = ($signed(_zz_1409) - $signed(_zz_3553));
  assign _zz_13843 = _zz_13844;
  assign _zz_13844 = ($signed(_zz_13845) >>> _zz_3556);
  assign _zz_13845 = _zz_13846;
  assign _zz_13846 = ($signed(_zz_1410) - $signed(_zz_3554));
  assign _zz_13847 = _zz_13848;
  assign _zz_13848 = ($signed(_zz_13849) >>> _zz_3557);
  assign _zz_13849 = _zz_13850;
  assign _zz_13850 = ($signed(_zz_1409) + $signed(_zz_3553));
  assign _zz_13851 = _zz_13852;
  assign _zz_13852 = ($signed(_zz_13853) >>> _zz_3557);
  assign _zz_13853 = _zz_13854;
  assign _zz_13854 = ($signed(_zz_1410) + $signed(_zz_3554));
  assign _zz_13855 = ($signed(twiddle_factor_table_32_real) + $signed(twiddle_factor_table_32_imag));
  assign _zz_13856 = fixTo_1059_dout;
  assign _zz_13857 = ($signed(_zz_1476) - $signed(_zz_1475));
  assign _zz_13858 = ($signed(_zz_1475) + $signed(_zz_1476));
  assign _zz_13859 = _zz_13860[15 : 0];
  assign _zz_13860 = fixTo_1061_dout;
  assign _zz_13861 = _zz_13862[15 : 0];
  assign _zz_13862 = fixTo_1060_dout;
  assign _zz_13863 = _zz_13864;
  assign _zz_13864 = ($signed(_zz_13865) >>> _zz_3561);
  assign _zz_13865 = _zz_13866;
  assign _zz_13866 = ($signed(_zz_1411) - $signed(_zz_3558));
  assign _zz_13867 = _zz_13868;
  assign _zz_13868 = ($signed(_zz_13869) >>> _zz_3561);
  assign _zz_13869 = _zz_13870;
  assign _zz_13870 = ($signed(_zz_1412) - $signed(_zz_3559));
  assign _zz_13871 = _zz_13872;
  assign _zz_13872 = ($signed(_zz_13873) >>> _zz_3562);
  assign _zz_13873 = _zz_13874;
  assign _zz_13874 = ($signed(_zz_1411) + $signed(_zz_3558));
  assign _zz_13875 = _zz_13876;
  assign _zz_13876 = ($signed(_zz_13877) >>> _zz_3562);
  assign _zz_13877 = _zz_13878;
  assign _zz_13878 = ($signed(_zz_1412) + $signed(_zz_3559));
  assign _zz_13879 = ($signed(twiddle_factor_table_33_real) + $signed(twiddle_factor_table_33_imag));
  assign _zz_13880 = fixTo_1062_dout;
  assign _zz_13881 = ($signed(_zz_1478) - $signed(_zz_1477));
  assign _zz_13882 = ($signed(_zz_1477) + $signed(_zz_1478));
  assign _zz_13883 = _zz_13884[15 : 0];
  assign _zz_13884 = fixTo_1064_dout;
  assign _zz_13885 = _zz_13886[15 : 0];
  assign _zz_13886 = fixTo_1063_dout;
  assign _zz_13887 = _zz_13888;
  assign _zz_13888 = ($signed(_zz_13889) >>> _zz_3566);
  assign _zz_13889 = _zz_13890;
  assign _zz_13890 = ($signed(_zz_1413) - $signed(_zz_3563));
  assign _zz_13891 = _zz_13892;
  assign _zz_13892 = ($signed(_zz_13893) >>> _zz_3566);
  assign _zz_13893 = _zz_13894;
  assign _zz_13894 = ($signed(_zz_1414) - $signed(_zz_3564));
  assign _zz_13895 = _zz_13896;
  assign _zz_13896 = ($signed(_zz_13897) >>> _zz_3567);
  assign _zz_13897 = _zz_13898;
  assign _zz_13898 = ($signed(_zz_1413) + $signed(_zz_3563));
  assign _zz_13899 = _zz_13900;
  assign _zz_13900 = ($signed(_zz_13901) >>> _zz_3567);
  assign _zz_13901 = _zz_13902;
  assign _zz_13902 = ($signed(_zz_1414) + $signed(_zz_3564));
  assign _zz_13903 = ($signed(twiddle_factor_table_34_real) + $signed(twiddle_factor_table_34_imag));
  assign _zz_13904 = fixTo_1065_dout;
  assign _zz_13905 = ($signed(_zz_1480) - $signed(_zz_1479));
  assign _zz_13906 = ($signed(_zz_1479) + $signed(_zz_1480));
  assign _zz_13907 = _zz_13908[15 : 0];
  assign _zz_13908 = fixTo_1067_dout;
  assign _zz_13909 = _zz_13910[15 : 0];
  assign _zz_13910 = fixTo_1066_dout;
  assign _zz_13911 = _zz_13912;
  assign _zz_13912 = ($signed(_zz_13913) >>> _zz_3571);
  assign _zz_13913 = _zz_13914;
  assign _zz_13914 = ($signed(_zz_1415) - $signed(_zz_3568));
  assign _zz_13915 = _zz_13916;
  assign _zz_13916 = ($signed(_zz_13917) >>> _zz_3571);
  assign _zz_13917 = _zz_13918;
  assign _zz_13918 = ($signed(_zz_1416) - $signed(_zz_3569));
  assign _zz_13919 = _zz_13920;
  assign _zz_13920 = ($signed(_zz_13921) >>> _zz_3572);
  assign _zz_13921 = _zz_13922;
  assign _zz_13922 = ($signed(_zz_1415) + $signed(_zz_3568));
  assign _zz_13923 = _zz_13924;
  assign _zz_13924 = ($signed(_zz_13925) >>> _zz_3572);
  assign _zz_13925 = _zz_13926;
  assign _zz_13926 = ($signed(_zz_1416) + $signed(_zz_3569));
  assign _zz_13927 = ($signed(twiddle_factor_table_35_real) + $signed(twiddle_factor_table_35_imag));
  assign _zz_13928 = fixTo_1068_dout;
  assign _zz_13929 = ($signed(_zz_1482) - $signed(_zz_1481));
  assign _zz_13930 = ($signed(_zz_1481) + $signed(_zz_1482));
  assign _zz_13931 = _zz_13932[15 : 0];
  assign _zz_13932 = fixTo_1070_dout;
  assign _zz_13933 = _zz_13934[15 : 0];
  assign _zz_13934 = fixTo_1069_dout;
  assign _zz_13935 = _zz_13936;
  assign _zz_13936 = ($signed(_zz_13937) >>> _zz_3576);
  assign _zz_13937 = _zz_13938;
  assign _zz_13938 = ($signed(_zz_1417) - $signed(_zz_3573));
  assign _zz_13939 = _zz_13940;
  assign _zz_13940 = ($signed(_zz_13941) >>> _zz_3576);
  assign _zz_13941 = _zz_13942;
  assign _zz_13942 = ($signed(_zz_1418) - $signed(_zz_3574));
  assign _zz_13943 = _zz_13944;
  assign _zz_13944 = ($signed(_zz_13945) >>> _zz_3577);
  assign _zz_13945 = _zz_13946;
  assign _zz_13946 = ($signed(_zz_1417) + $signed(_zz_3573));
  assign _zz_13947 = _zz_13948;
  assign _zz_13948 = ($signed(_zz_13949) >>> _zz_3577);
  assign _zz_13949 = _zz_13950;
  assign _zz_13950 = ($signed(_zz_1418) + $signed(_zz_3574));
  assign _zz_13951 = ($signed(twiddle_factor_table_36_real) + $signed(twiddle_factor_table_36_imag));
  assign _zz_13952 = fixTo_1071_dout;
  assign _zz_13953 = ($signed(_zz_1484) - $signed(_zz_1483));
  assign _zz_13954 = ($signed(_zz_1483) + $signed(_zz_1484));
  assign _zz_13955 = _zz_13956[15 : 0];
  assign _zz_13956 = fixTo_1073_dout;
  assign _zz_13957 = _zz_13958[15 : 0];
  assign _zz_13958 = fixTo_1072_dout;
  assign _zz_13959 = _zz_13960;
  assign _zz_13960 = ($signed(_zz_13961) >>> _zz_3581);
  assign _zz_13961 = _zz_13962;
  assign _zz_13962 = ($signed(_zz_1419) - $signed(_zz_3578));
  assign _zz_13963 = _zz_13964;
  assign _zz_13964 = ($signed(_zz_13965) >>> _zz_3581);
  assign _zz_13965 = _zz_13966;
  assign _zz_13966 = ($signed(_zz_1420) - $signed(_zz_3579));
  assign _zz_13967 = _zz_13968;
  assign _zz_13968 = ($signed(_zz_13969) >>> _zz_3582);
  assign _zz_13969 = _zz_13970;
  assign _zz_13970 = ($signed(_zz_1419) + $signed(_zz_3578));
  assign _zz_13971 = _zz_13972;
  assign _zz_13972 = ($signed(_zz_13973) >>> _zz_3582);
  assign _zz_13973 = _zz_13974;
  assign _zz_13974 = ($signed(_zz_1420) + $signed(_zz_3579));
  assign _zz_13975 = ($signed(twiddle_factor_table_37_real) + $signed(twiddle_factor_table_37_imag));
  assign _zz_13976 = fixTo_1074_dout;
  assign _zz_13977 = ($signed(_zz_1486) - $signed(_zz_1485));
  assign _zz_13978 = ($signed(_zz_1485) + $signed(_zz_1486));
  assign _zz_13979 = _zz_13980[15 : 0];
  assign _zz_13980 = fixTo_1076_dout;
  assign _zz_13981 = _zz_13982[15 : 0];
  assign _zz_13982 = fixTo_1075_dout;
  assign _zz_13983 = _zz_13984;
  assign _zz_13984 = ($signed(_zz_13985) >>> _zz_3586);
  assign _zz_13985 = _zz_13986;
  assign _zz_13986 = ($signed(_zz_1421) - $signed(_zz_3583));
  assign _zz_13987 = _zz_13988;
  assign _zz_13988 = ($signed(_zz_13989) >>> _zz_3586);
  assign _zz_13989 = _zz_13990;
  assign _zz_13990 = ($signed(_zz_1422) - $signed(_zz_3584));
  assign _zz_13991 = _zz_13992;
  assign _zz_13992 = ($signed(_zz_13993) >>> _zz_3587);
  assign _zz_13993 = _zz_13994;
  assign _zz_13994 = ($signed(_zz_1421) + $signed(_zz_3583));
  assign _zz_13995 = _zz_13996;
  assign _zz_13996 = ($signed(_zz_13997) >>> _zz_3587);
  assign _zz_13997 = _zz_13998;
  assign _zz_13998 = ($signed(_zz_1422) + $signed(_zz_3584));
  assign _zz_13999 = ($signed(twiddle_factor_table_38_real) + $signed(twiddle_factor_table_38_imag));
  assign _zz_14000 = fixTo_1077_dout;
  assign _zz_14001 = ($signed(_zz_1488) - $signed(_zz_1487));
  assign _zz_14002 = ($signed(_zz_1487) + $signed(_zz_1488));
  assign _zz_14003 = _zz_14004[15 : 0];
  assign _zz_14004 = fixTo_1079_dout;
  assign _zz_14005 = _zz_14006[15 : 0];
  assign _zz_14006 = fixTo_1078_dout;
  assign _zz_14007 = _zz_14008;
  assign _zz_14008 = ($signed(_zz_14009) >>> _zz_3591);
  assign _zz_14009 = _zz_14010;
  assign _zz_14010 = ($signed(_zz_1423) - $signed(_zz_3588));
  assign _zz_14011 = _zz_14012;
  assign _zz_14012 = ($signed(_zz_14013) >>> _zz_3591);
  assign _zz_14013 = _zz_14014;
  assign _zz_14014 = ($signed(_zz_1424) - $signed(_zz_3589));
  assign _zz_14015 = _zz_14016;
  assign _zz_14016 = ($signed(_zz_14017) >>> _zz_3592);
  assign _zz_14017 = _zz_14018;
  assign _zz_14018 = ($signed(_zz_1423) + $signed(_zz_3588));
  assign _zz_14019 = _zz_14020;
  assign _zz_14020 = ($signed(_zz_14021) >>> _zz_3592);
  assign _zz_14021 = _zz_14022;
  assign _zz_14022 = ($signed(_zz_1424) + $signed(_zz_3589));
  assign _zz_14023 = ($signed(twiddle_factor_table_39_real) + $signed(twiddle_factor_table_39_imag));
  assign _zz_14024 = fixTo_1080_dout;
  assign _zz_14025 = ($signed(_zz_1490) - $signed(_zz_1489));
  assign _zz_14026 = ($signed(_zz_1489) + $signed(_zz_1490));
  assign _zz_14027 = _zz_14028[15 : 0];
  assign _zz_14028 = fixTo_1082_dout;
  assign _zz_14029 = _zz_14030[15 : 0];
  assign _zz_14030 = fixTo_1081_dout;
  assign _zz_14031 = _zz_14032;
  assign _zz_14032 = ($signed(_zz_14033) >>> _zz_3596);
  assign _zz_14033 = _zz_14034;
  assign _zz_14034 = ($signed(_zz_1425) - $signed(_zz_3593));
  assign _zz_14035 = _zz_14036;
  assign _zz_14036 = ($signed(_zz_14037) >>> _zz_3596);
  assign _zz_14037 = _zz_14038;
  assign _zz_14038 = ($signed(_zz_1426) - $signed(_zz_3594));
  assign _zz_14039 = _zz_14040;
  assign _zz_14040 = ($signed(_zz_14041) >>> _zz_3597);
  assign _zz_14041 = _zz_14042;
  assign _zz_14042 = ($signed(_zz_1425) + $signed(_zz_3593));
  assign _zz_14043 = _zz_14044;
  assign _zz_14044 = ($signed(_zz_14045) >>> _zz_3597);
  assign _zz_14045 = _zz_14046;
  assign _zz_14046 = ($signed(_zz_1426) + $signed(_zz_3594));
  assign _zz_14047 = ($signed(twiddle_factor_table_40_real) + $signed(twiddle_factor_table_40_imag));
  assign _zz_14048 = fixTo_1083_dout;
  assign _zz_14049 = ($signed(_zz_1492) - $signed(_zz_1491));
  assign _zz_14050 = ($signed(_zz_1491) + $signed(_zz_1492));
  assign _zz_14051 = _zz_14052[15 : 0];
  assign _zz_14052 = fixTo_1085_dout;
  assign _zz_14053 = _zz_14054[15 : 0];
  assign _zz_14054 = fixTo_1084_dout;
  assign _zz_14055 = _zz_14056;
  assign _zz_14056 = ($signed(_zz_14057) >>> _zz_3601);
  assign _zz_14057 = _zz_14058;
  assign _zz_14058 = ($signed(_zz_1427) - $signed(_zz_3598));
  assign _zz_14059 = _zz_14060;
  assign _zz_14060 = ($signed(_zz_14061) >>> _zz_3601);
  assign _zz_14061 = _zz_14062;
  assign _zz_14062 = ($signed(_zz_1428) - $signed(_zz_3599));
  assign _zz_14063 = _zz_14064;
  assign _zz_14064 = ($signed(_zz_14065) >>> _zz_3602);
  assign _zz_14065 = _zz_14066;
  assign _zz_14066 = ($signed(_zz_1427) + $signed(_zz_3598));
  assign _zz_14067 = _zz_14068;
  assign _zz_14068 = ($signed(_zz_14069) >>> _zz_3602);
  assign _zz_14069 = _zz_14070;
  assign _zz_14070 = ($signed(_zz_1428) + $signed(_zz_3599));
  assign _zz_14071 = ($signed(twiddle_factor_table_41_real) + $signed(twiddle_factor_table_41_imag));
  assign _zz_14072 = fixTo_1086_dout;
  assign _zz_14073 = ($signed(_zz_1494) - $signed(_zz_1493));
  assign _zz_14074 = ($signed(_zz_1493) + $signed(_zz_1494));
  assign _zz_14075 = _zz_14076[15 : 0];
  assign _zz_14076 = fixTo_1088_dout;
  assign _zz_14077 = _zz_14078[15 : 0];
  assign _zz_14078 = fixTo_1087_dout;
  assign _zz_14079 = _zz_14080;
  assign _zz_14080 = ($signed(_zz_14081) >>> _zz_3606);
  assign _zz_14081 = _zz_14082;
  assign _zz_14082 = ($signed(_zz_1429) - $signed(_zz_3603));
  assign _zz_14083 = _zz_14084;
  assign _zz_14084 = ($signed(_zz_14085) >>> _zz_3606);
  assign _zz_14085 = _zz_14086;
  assign _zz_14086 = ($signed(_zz_1430) - $signed(_zz_3604));
  assign _zz_14087 = _zz_14088;
  assign _zz_14088 = ($signed(_zz_14089) >>> _zz_3607);
  assign _zz_14089 = _zz_14090;
  assign _zz_14090 = ($signed(_zz_1429) + $signed(_zz_3603));
  assign _zz_14091 = _zz_14092;
  assign _zz_14092 = ($signed(_zz_14093) >>> _zz_3607);
  assign _zz_14093 = _zz_14094;
  assign _zz_14094 = ($signed(_zz_1430) + $signed(_zz_3604));
  assign _zz_14095 = ($signed(twiddle_factor_table_42_real) + $signed(twiddle_factor_table_42_imag));
  assign _zz_14096 = fixTo_1089_dout;
  assign _zz_14097 = ($signed(_zz_1496) - $signed(_zz_1495));
  assign _zz_14098 = ($signed(_zz_1495) + $signed(_zz_1496));
  assign _zz_14099 = _zz_14100[15 : 0];
  assign _zz_14100 = fixTo_1091_dout;
  assign _zz_14101 = _zz_14102[15 : 0];
  assign _zz_14102 = fixTo_1090_dout;
  assign _zz_14103 = _zz_14104;
  assign _zz_14104 = ($signed(_zz_14105) >>> _zz_3611);
  assign _zz_14105 = _zz_14106;
  assign _zz_14106 = ($signed(_zz_1431) - $signed(_zz_3608));
  assign _zz_14107 = _zz_14108;
  assign _zz_14108 = ($signed(_zz_14109) >>> _zz_3611);
  assign _zz_14109 = _zz_14110;
  assign _zz_14110 = ($signed(_zz_1432) - $signed(_zz_3609));
  assign _zz_14111 = _zz_14112;
  assign _zz_14112 = ($signed(_zz_14113) >>> _zz_3612);
  assign _zz_14113 = _zz_14114;
  assign _zz_14114 = ($signed(_zz_1431) + $signed(_zz_3608));
  assign _zz_14115 = _zz_14116;
  assign _zz_14116 = ($signed(_zz_14117) >>> _zz_3612);
  assign _zz_14117 = _zz_14118;
  assign _zz_14118 = ($signed(_zz_1432) + $signed(_zz_3609));
  assign _zz_14119 = ($signed(twiddle_factor_table_43_real) + $signed(twiddle_factor_table_43_imag));
  assign _zz_14120 = fixTo_1092_dout;
  assign _zz_14121 = ($signed(_zz_1498) - $signed(_zz_1497));
  assign _zz_14122 = ($signed(_zz_1497) + $signed(_zz_1498));
  assign _zz_14123 = _zz_14124[15 : 0];
  assign _zz_14124 = fixTo_1094_dout;
  assign _zz_14125 = _zz_14126[15 : 0];
  assign _zz_14126 = fixTo_1093_dout;
  assign _zz_14127 = _zz_14128;
  assign _zz_14128 = ($signed(_zz_14129) >>> _zz_3616);
  assign _zz_14129 = _zz_14130;
  assign _zz_14130 = ($signed(_zz_1433) - $signed(_zz_3613));
  assign _zz_14131 = _zz_14132;
  assign _zz_14132 = ($signed(_zz_14133) >>> _zz_3616);
  assign _zz_14133 = _zz_14134;
  assign _zz_14134 = ($signed(_zz_1434) - $signed(_zz_3614));
  assign _zz_14135 = _zz_14136;
  assign _zz_14136 = ($signed(_zz_14137) >>> _zz_3617);
  assign _zz_14137 = _zz_14138;
  assign _zz_14138 = ($signed(_zz_1433) + $signed(_zz_3613));
  assign _zz_14139 = _zz_14140;
  assign _zz_14140 = ($signed(_zz_14141) >>> _zz_3617);
  assign _zz_14141 = _zz_14142;
  assign _zz_14142 = ($signed(_zz_1434) + $signed(_zz_3614));
  assign _zz_14143 = ($signed(twiddle_factor_table_44_real) + $signed(twiddle_factor_table_44_imag));
  assign _zz_14144 = fixTo_1095_dout;
  assign _zz_14145 = ($signed(_zz_1500) - $signed(_zz_1499));
  assign _zz_14146 = ($signed(_zz_1499) + $signed(_zz_1500));
  assign _zz_14147 = _zz_14148[15 : 0];
  assign _zz_14148 = fixTo_1097_dout;
  assign _zz_14149 = _zz_14150[15 : 0];
  assign _zz_14150 = fixTo_1096_dout;
  assign _zz_14151 = _zz_14152;
  assign _zz_14152 = ($signed(_zz_14153) >>> _zz_3621);
  assign _zz_14153 = _zz_14154;
  assign _zz_14154 = ($signed(_zz_1435) - $signed(_zz_3618));
  assign _zz_14155 = _zz_14156;
  assign _zz_14156 = ($signed(_zz_14157) >>> _zz_3621);
  assign _zz_14157 = _zz_14158;
  assign _zz_14158 = ($signed(_zz_1436) - $signed(_zz_3619));
  assign _zz_14159 = _zz_14160;
  assign _zz_14160 = ($signed(_zz_14161) >>> _zz_3622);
  assign _zz_14161 = _zz_14162;
  assign _zz_14162 = ($signed(_zz_1435) + $signed(_zz_3618));
  assign _zz_14163 = _zz_14164;
  assign _zz_14164 = ($signed(_zz_14165) >>> _zz_3622);
  assign _zz_14165 = _zz_14166;
  assign _zz_14166 = ($signed(_zz_1436) + $signed(_zz_3619));
  assign _zz_14167 = ($signed(twiddle_factor_table_45_real) + $signed(twiddle_factor_table_45_imag));
  assign _zz_14168 = fixTo_1098_dout;
  assign _zz_14169 = ($signed(_zz_1502) - $signed(_zz_1501));
  assign _zz_14170 = ($signed(_zz_1501) + $signed(_zz_1502));
  assign _zz_14171 = _zz_14172[15 : 0];
  assign _zz_14172 = fixTo_1100_dout;
  assign _zz_14173 = _zz_14174[15 : 0];
  assign _zz_14174 = fixTo_1099_dout;
  assign _zz_14175 = _zz_14176;
  assign _zz_14176 = ($signed(_zz_14177) >>> _zz_3626);
  assign _zz_14177 = _zz_14178;
  assign _zz_14178 = ($signed(_zz_1437) - $signed(_zz_3623));
  assign _zz_14179 = _zz_14180;
  assign _zz_14180 = ($signed(_zz_14181) >>> _zz_3626);
  assign _zz_14181 = _zz_14182;
  assign _zz_14182 = ($signed(_zz_1438) - $signed(_zz_3624));
  assign _zz_14183 = _zz_14184;
  assign _zz_14184 = ($signed(_zz_14185) >>> _zz_3627);
  assign _zz_14185 = _zz_14186;
  assign _zz_14186 = ($signed(_zz_1437) + $signed(_zz_3623));
  assign _zz_14187 = _zz_14188;
  assign _zz_14188 = ($signed(_zz_14189) >>> _zz_3627);
  assign _zz_14189 = _zz_14190;
  assign _zz_14190 = ($signed(_zz_1438) + $signed(_zz_3624));
  assign _zz_14191 = ($signed(twiddle_factor_table_46_real) + $signed(twiddle_factor_table_46_imag));
  assign _zz_14192 = fixTo_1101_dout;
  assign _zz_14193 = ($signed(_zz_1504) - $signed(_zz_1503));
  assign _zz_14194 = ($signed(_zz_1503) + $signed(_zz_1504));
  assign _zz_14195 = _zz_14196[15 : 0];
  assign _zz_14196 = fixTo_1103_dout;
  assign _zz_14197 = _zz_14198[15 : 0];
  assign _zz_14198 = fixTo_1102_dout;
  assign _zz_14199 = _zz_14200;
  assign _zz_14200 = ($signed(_zz_14201) >>> _zz_3631);
  assign _zz_14201 = _zz_14202;
  assign _zz_14202 = ($signed(_zz_1439) - $signed(_zz_3628));
  assign _zz_14203 = _zz_14204;
  assign _zz_14204 = ($signed(_zz_14205) >>> _zz_3631);
  assign _zz_14205 = _zz_14206;
  assign _zz_14206 = ($signed(_zz_1440) - $signed(_zz_3629));
  assign _zz_14207 = _zz_14208;
  assign _zz_14208 = ($signed(_zz_14209) >>> _zz_3632);
  assign _zz_14209 = _zz_14210;
  assign _zz_14210 = ($signed(_zz_1439) + $signed(_zz_3628));
  assign _zz_14211 = _zz_14212;
  assign _zz_14212 = ($signed(_zz_14213) >>> _zz_3632);
  assign _zz_14213 = _zz_14214;
  assign _zz_14214 = ($signed(_zz_1440) + $signed(_zz_3629));
  assign _zz_14215 = ($signed(twiddle_factor_table_47_real) + $signed(twiddle_factor_table_47_imag));
  assign _zz_14216 = fixTo_1104_dout;
  assign _zz_14217 = ($signed(_zz_1506) - $signed(_zz_1505));
  assign _zz_14218 = ($signed(_zz_1505) + $signed(_zz_1506));
  assign _zz_14219 = _zz_14220[15 : 0];
  assign _zz_14220 = fixTo_1106_dout;
  assign _zz_14221 = _zz_14222[15 : 0];
  assign _zz_14222 = fixTo_1105_dout;
  assign _zz_14223 = _zz_14224;
  assign _zz_14224 = ($signed(_zz_14225) >>> _zz_3636);
  assign _zz_14225 = _zz_14226;
  assign _zz_14226 = ($signed(_zz_1441) - $signed(_zz_3633));
  assign _zz_14227 = _zz_14228;
  assign _zz_14228 = ($signed(_zz_14229) >>> _zz_3636);
  assign _zz_14229 = _zz_14230;
  assign _zz_14230 = ($signed(_zz_1442) - $signed(_zz_3634));
  assign _zz_14231 = _zz_14232;
  assign _zz_14232 = ($signed(_zz_14233) >>> _zz_3637);
  assign _zz_14233 = _zz_14234;
  assign _zz_14234 = ($signed(_zz_1441) + $signed(_zz_3633));
  assign _zz_14235 = _zz_14236;
  assign _zz_14236 = ($signed(_zz_14237) >>> _zz_3637);
  assign _zz_14237 = _zz_14238;
  assign _zz_14238 = ($signed(_zz_1442) + $signed(_zz_3634));
  assign _zz_14239 = ($signed(twiddle_factor_table_48_real) + $signed(twiddle_factor_table_48_imag));
  assign _zz_14240 = fixTo_1107_dout;
  assign _zz_14241 = ($signed(_zz_1508) - $signed(_zz_1507));
  assign _zz_14242 = ($signed(_zz_1507) + $signed(_zz_1508));
  assign _zz_14243 = _zz_14244[15 : 0];
  assign _zz_14244 = fixTo_1109_dout;
  assign _zz_14245 = _zz_14246[15 : 0];
  assign _zz_14246 = fixTo_1108_dout;
  assign _zz_14247 = _zz_14248;
  assign _zz_14248 = ($signed(_zz_14249) >>> _zz_3641);
  assign _zz_14249 = _zz_14250;
  assign _zz_14250 = ($signed(_zz_1443) - $signed(_zz_3638));
  assign _zz_14251 = _zz_14252;
  assign _zz_14252 = ($signed(_zz_14253) >>> _zz_3641);
  assign _zz_14253 = _zz_14254;
  assign _zz_14254 = ($signed(_zz_1444) - $signed(_zz_3639));
  assign _zz_14255 = _zz_14256;
  assign _zz_14256 = ($signed(_zz_14257) >>> _zz_3642);
  assign _zz_14257 = _zz_14258;
  assign _zz_14258 = ($signed(_zz_1443) + $signed(_zz_3638));
  assign _zz_14259 = _zz_14260;
  assign _zz_14260 = ($signed(_zz_14261) >>> _zz_3642);
  assign _zz_14261 = _zz_14262;
  assign _zz_14262 = ($signed(_zz_1444) + $signed(_zz_3639));
  assign _zz_14263 = ($signed(twiddle_factor_table_49_real) + $signed(twiddle_factor_table_49_imag));
  assign _zz_14264 = fixTo_1110_dout;
  assign _zz_14265 = ($signed(_zz_1510) - $signed(_zz_1509));
  assign _zz_14266 = ($signed(_zz_1509) + $signed(_zz_1510));
  assign _zz_14267 = _zz_14268[15 : 0];
  assign _zz_14268 = fixTo_1112_dout;
  assign _zz_14269 = _zz_14270[15 : 0];
  assign _zz_14270 = fixTo_1111_dout;
  assign _zz_14271 = _zz_14272;
  assign _zz_14272 = ($signed(_zz_14273) >>> _zz_3646);
  assign _zz_14273 = _zz_14274;
  assign _zz_14274 = ($signed(_zz_1445) - $signed(_zz_3643));
  assign _zz_14275 = _zz_14276;
  assign _zz_14276 = ($signed(_zz_14277) >>> _zz_3646);
  assign _zz_14277 = _zz_14278;
  assign _zz_14278 = ($signed(_zz_1446) - $signed(_zz_3644));
  assign _zz_14279 = _zz_14280;
  assign _zz_14280 = ($signed(_zz_14281) >>> _zz_3647);
  assign _zz_14281 = _zz_14282;
  assign _zz_14282 = ($signed(_zz_1445) + $signed(_zz_3643));
  assign _zz_14283 = _zz_14284;
  assign _zz_14284 = ($signed(_zz_14285) >>> _zz_3647);
  assign _zz_14285 = _zz_14286;
  assign _zz_14286 = ($signed(_zz_1446) + $signed(_zz_3644));
  assign _zz_14287 = ($signed(twiddle_factor_table_50_real) + $signed(twiddle_factor_table_50_imag));
  assign _zz_14288 = fixTo_1113_dout;
  assign _zz_14289 = ($signed(_zz_1512) - $signed(_zz_1511));
  assign _zz_14290 = ($signed(_zz_1511) + $signed(_zz_1512));
  assign _zz_14291 = _zz_14292[15 : 0];
  assign _zz_14292 = fixTo_1115_dout;
  assign _zz_14293 = _zz_14294[15 : 0];
  assign _zz_14294 = fixTo_1114_dout;
  assign _zz_14295 = _zz_14296;
  assign _zz_14296 = ($signed(_zz_14297) >>> _zz_3651);
  assign _zz_14297 = _zz_14298;
  assign _zz_14298 = ($signed(_zz_1447) - $signed(_zz_3648));
  assign _zz_14299 = _zz_14300;
  assign _zz_14300 = ($signed(_zz_14301) >>> _zz_3651);
  assign _zz_14301 = _zz_14302;
  assign _zz_14302 = ($signed(_zz_1448) - $signed(_zz_3649));
  assign _zz_14303 = _zz_14304;
  assign _zz_14304 = ($signed(_zz_14305) >>> _zz_3652);
  assign _zz_14305 = _zz_14306;
  assign _zz_14306 = ($signed(_zz_1447) + $signed(_zz_3648));
  assign _zz_14307 = _zz_14308;
  assign _zz_14308 = ($signed(_zz_14309) >>> _zz_3652);
  assign _zz_14309 = _zz_14310;
  assign _zz_14310 = ($signed(_zz_1448) + $signed(_zz_3649));
  assign _zz_14311 = ($signed(twiddle_factor_table_51_real) + $signed(twiddle_factor_table_51_imag));
  assign _zz_14312 = fixTo_1116_dout;
  assign _zz_14313 = ($signed(_zz_1514) - $signed(_zz_1513));
  assign _zz_14314 = ($signed(_zz_1513) + $signed(_zz_1514));
  assign _zz_14315 = _zz_14316[15 : 0];
  assign _zz_14316 = fixTo_1118_dout;
  assign _zz_14317 = _zz_14318[15 : 0];
  assign _zz_14318 = fixTo_1117_dout;
  assign _zz_14319 = _zz_14320;
  assign _zz_14320 = ($signed(_zz_14321) >>> _zz_3656);
  assign _zz_14321 = _zz_14322;
  assign _zz_14322 = ($signed(_zz_1449) - $signed(_zz_3653));
  assign _zz_14323 = _zz_14324;
  assign _zz_14324 = ($signed(_zz_14325) >>> _zz_3656);
  assign _zz_14325 = _zz_14326;
  assign _zz_14326 = ($signed(_zz_1450) - $signed(_zz_3654));
  assign _zz_14327 = _zz_14328;
  assign _zz_14328 = ($signed(_zz_14329) >>> _zz_3657);
  assign _zz_14329 = _zz_14330;
  assign _zz_14330 = ($signed(_zz_1449) + $signed(_zz_3653));
  assign _zz_14331 = _zz_14332;
  assign _zz_14332 = ($signed(_zz_14333) >>> _zz_3657);
  assign _zz_14333 = _zz_14334;
  assign _zz_14334 = ($signed(_zz_1450) + $signed(_zz_3654));
  assign _zz_14335 = ($signed(twiddle_factor_table_52_real) + $signed(twiddle_factor_table_52_imag));
  assign _zz_14336 = fixTo_1119_dout;
  assign _zz_14337 = ($signed(_zz_1516) - $signed(_zz_1515));
  assign _zz_14338 = ($signed(_zz_1515) + $signed(_zz_1516));
  assign _zz_14339 = _zz_14340[15 : 0];
  assign _zz_14340 = fixTo_1121_dout;
  assign _zz_14341 = _zz_14342[15 : 0];
  assign _zz_14342 = fixTo_1120_dout;
  assign _zz_14343 = _zz_14344;
  assign _zz_14344 = ($signed(_zz_14345) >>> _zz_3661);
  assign _zz_14345 = _zz_14346;
  assign _zz_14346 = ($signed(_zz_1451) - $signed(_zz_3658));
  assign _zz_14347 = _zz_14348;
  assign _zz_14348 = ($signed(_zz_14349) >>> _zz_3661);
  assign _zz_14349 = _zz_14350;
  assign _zz_14350 = ($signed(_zz_1452) - $signed(_zz_3659));
  assign _zz_14351 = _zz_14352;
  assign _zz_14352 = ($signed(_zz_14353) >>> _zz_3662);
  assign _zz_14353 = _zz_14354;
  assign _zz_14354 = ($signed(_zz_1451) + $signed(_zz_3658));
  assign _zz_14355 = _zz_14356;
  assign _zz_14356 = ($signed(_zz_14357) >>> _zz_3662);
  assign _zz_14357 = _zz_14358;
  assign _zz_14358 = ($signed(_zz_1452) + $signed(_zz_3659));
  assign _zz_14359 = ($signed(twiddle_factor_table_53_real) + $signed(twiddle_factor_table_53_imag));
  assign _zz_14360 = fixTo_1122_dout;
  assign _zz_14361 = ($signed(_zz_1518) - $signed(_zz_1517));
  assign _zz_14362 = ($signed(_zz_1517) + $signed(_zz_1518));
  assign _zz_14363 = _zz_14364[15 : 0];
  assign _zz_14364 = fixTo_1124_dout;
  assign _zz_14365 = _zz_14366[15 : 0];
  assign _zz_14366 = fixTo_1123_dout;
  assign _zz_14367 = _zz_14368;
  assign _zz_14368 = ($signed(_zz_14369) >>> _zz_3666);
  assign _zz_14369 = _zz_14370;
  assign _zz_14370 = ($signed(_zz_1453) - $signed(_zz_3663));
  assign _zz_14371 = _zz_14372;
  assign _zz_14372 = ($signed(_zz_14373) >>> _zz_3666);
  assign _zz_14373 = _zz_14374;
  assign _zz_14374 = ($signed(_zz_1454) - $signed(_zz_3664));
  assign _zz_14375 = _zz_14376;
  assign _zz_14376 = ($signed(_zz_14377) >>> _zz_3667);
  assign _zz_14377 = _zz_14378;
  assign _zz_14378 = ($signed(_zz_1453) + $signed(_zz_3663));
  assign _zz_14379 = _zz_14380;
  assign _zz_14380 = ($signed(_zz_14381) >>> _zz_3667);
  assign _zz_14381 = _zz_14382;
  assign _zz_14382 = ($signed(_zz_1454) + $signed(_zz_3664));
  assign _zz_14383 = ($signed(twiddle_factor_table_54_real) + $signed(twiddle_factor_table_54_imag));
  assign _zz_14384 = fixTo_1125_dout;
  assign _zz_14385 = ($signed(_zz_1520) - $signed(_zz_1519));
  assign _zz_14386 = ($signed(_zz_1519) + $signed(_zz_1520));
  assign _zz_14387 = _zz_14388[15 : 0];
  assign _zz_14388 = fixTo_1127_dout;
  assign _zz_14389 = _zz_14390[15 : 0];
  assign _zz_14390 = fixTo_1126_dout;
  assign _zz_14391 = _zz_14392;
  assign _zz_14392 = ($signed(_zz_14393) >>> _zz_3671);
  assign _zz_14393 = _zz_14394;
  assign _zz_14394 = ($signed(_zz_1455) - $signed(_zz_3668));
  assign _zz_14395 = _zz_14396;
  assign _zz_14396 = ($signed(_zz_14397) >>> _zz_3671);
  assign _zz_14397 = _zz_14398;
  assign _zz_14398 = ($signed(_zz_1456) - $signed(_zz_3669));
  assign _zz_14399 = _zz_14400;
  assign _zz_14400 = ($signed(_zz_14401) >>> _zz_3672);
  assign _zz_14401 = _zz_14402;
  assign _zz_14402 = ($signed(_zz_1455) + $signed(_zz_3668));
  assign _zz_14403 = _zz_14404;
  assign _zz_14404 = ($signed(_zz_14405) >>> _zz_3672);
  assign _zz_14405 = _zz_14406;
  assign _zz_14406 = ($signed(_zz_1456) + $signed(_zz_3669));
  assign _zz_14407 = ($signed(twiddle_factor_table_55_real) + $signed(twiddle_factor_table_55_imag));
  assign _zz_14408 = fixTo_1128_dout;
  assign _zz_14409 = ($signed(_zz_1522) - $signed(_zz_1521));
  assign _zz_14410 = ($signed(_zz_1521) + $signed(_zz_1522));
  assign _zz_14411 = _zz_14412[15 : 0];
  assign _zz_14412 = fixTo_1130_dout;
  assign _zz_14413 = _zz_14414[15 : 0];
  assign _zz_14414 = fixTo_1129_dout;
  assign _zz_14415 = _zz_14416;
  assign _zz_14416 = ($signed(_zz_14417) >>> _zz_3676);
  assign _zz_14417 = _zz_14418;
  assign _zz_14418 = ($signed(_zz_1457) - $signed(_zz_3673));
  assign _zz_14419 = _zz_14420;
  assign _zz_14420 = ($signed(_zz_14421) >>> _zz_3676);
  assign _zz_14421 = _zz_14422;
  assign _zz_14422 = ($signed(_zz_1458) - $signed(_zz_3674));
  assign _zz_14423 = _zz_14424;
  assign _zz_14424 = ($signed(_zz_14425) >>> _zz_3677);
  assign _zz_14425 = _zz_14426;
  assign _zz_14426 = ($signed(_zz_1457) + $signed(_zz_3673));
  assign _zz_14427 = _zz_14428;
  assign _zz_14428 = ($signed(_zz_14429) >>> _zz_3677);
  assign _zz_14429 = _zz_14430;
  assign _zz_14430 = ($signed(_zz_1458) + $signed(_zz_3674));
  assign _zz_14431 = ($signed(twiddle_factor_table_56_real) + $signed(twiddle_factor_table_56_imag));
  assign _zz_14432 = fixTo_1131_dout;
  assign _zz_14433 = ($signed(_zz_1524) - $signed(_zz_1523));
  assign _zz_14434 = ($signed(_zz_1523) + $signed(_zz_1524));
  assign _zz_14435 = _zz_14436[15 : 0];
  assign _zz_14436 = fixTo_1133_dout;
  assign _zz_14437 = _zz_14438[15 : 0];
  assign _zz_14438 = fixTo_1132_dout;
  assign _zz_14439 = _zz_14440;
  assign _zz_14440 = ($signed(_zz_14441) >>> _zz_3681);
  assign _zz_14441 = _zz_14442;
  assign _zz_14442 = ($signed(_zz_1459) - $signed(_zz_3678));
  assign _zz_14443 = _zz_14444;
  assign _zz_14444 = ($signed(_zz_14445) >>> _zz_3681);
  assign _zz_14445 = _zz_14446;
  assign _zz_14446 = ($signed(_zz_1460) - $signed(_zz_3679));
  assign _zz_14447 = _zz_14448;
  assign _zz_14448 = ($signed(_zz_14449) >>> _zz_3682);
  assign _zz_14449 = _zz_14450;
  assign _zz_14450 = ($signed(_zz_1459) + $signed(_zz_3678));
  assign _zz_14451 = _zz_14452;
  assign _zz_14452 = ($signed(_zz_14453) >>> _zz_3682);
  assign _zz_14453 = _zz_14454;
  assign _zz_14454 = ($signed(_zz_1460) + $signed(_zz_3679));
  assign _zz_14455 = ($signed(twiddle_factor_table_57_real) + $signed(twiddle_factor_table_57_imag));
  assign _zz_14456 = fixTo_1134_dout;
  assign _zz_14457 = ($signed(_zz_1526) - $signed(_zz_1525));
  assign _zz_14458 = ($signed(_zz_1525) + $signed(_zz_1526));
  assign _zz_14459 = _zz_14460[15 : 0];
  assign _zz_14460 = fixTo_1136_dout;
  assign _zz_14461 = _zz_14462[15 : 0];
  assign _zz_14462 = fixTo_1135_dout;
  assign _zz_14463 = _zz_14464;
  assign _zz_14464 = ($signed(_zz_14465) >>> _zz_3686);
  assign _zz_14465 = _zz_14466;
  assign _zz_14466 = ($signed(_zz_1461) - $signed(_zz_3683));
  assign _zz_14467 = _zz_14468;
  assign _zz_14468 = ($signed(_zz_14469) >>> _zz_3686);
  assign _zz_14469 = _zz_14470;
  assign _zz_14470 = ($signed(_zz_1462) - $signed(_zz_3684));
  assign _zz_14471 = _zz_14472;
  assign _zz_14472 = ($signed(_zz_14473) >>> _zz_3687);
  assign _zz_14473 = _zz_14474;
  assign _zz_14474 = ($signed(_zz_1461) + $signed(_zz_3683));
  assign _zz_14475 = _zz_14476;
  assign _zz_14476 = ($signed(_zz_14477) >>> _zz_3687);
  assign _zz_14477 = _zz_14478;
  assign _zz_14478 = ($signed(_zz_1462) + $signed(_zz_3684));
  assign _zz_14479 = ($signed(twiddle_factor_table_58_real) + $signed(twiddle_factor_table_58_imag));
  assign _zz_14480 = fixTo_1137_dout;
  assign _zz_14481 = ($signed(_zz_1528) - $signed(_zz_1527));
  assign _zz_14482 = ($signed(_zz_1527) + $signed(_zz_1528));
  assign _zz_14483 = _zz_14484[15 : 0];
  assign _zz_14484 = fixTo_1139_dout;
  assign _zz_14485 = _zz_14486[15 : 0];
  assign _zz_14486 = fixTo_1138_dout;
  assign _zz_14487 = _zz_14488;
  assign _zz_14488 = ($signed(_zz_14489) >>> _zz_3691);
  assign _zz_14489 = _zz_14490;
  assign _zz_14490 = ($signed(_zz_1463) - $signed(_zz_3688));
  assign _zz_14491 = _zz_14492;
  assign _zz_14492 = ($signed(_zz_14493) >>> _zz_3691);
  assign _zz_14493 = _zz_14494;
  assign _zz_14494 = ($signed(_zz_1464) - $signed(_zz_3689));
  assign _zz_14495 = _zz_14496;
  assign _zz_14496 = ($signed(_zz_14497) >>> _zz_3692);
  assign _zz_14497 = _zz_14498;
  assign _zz_14498 = ($signed(_zz_1463) + $signed(_zz_3688));
  assign _zz_14499 = _zz_14500;
  assign _zz_14500 = ($signed(_zz_14501) >>> _zz_3692);
  assign _zz_14501 = _zz_14502;
  assign _zz_14502 = ($signed(_zz_1464) + $signed(_zz_3689));
  assign _zz_14503 = ($signed(twiddle_factor_table_59_real) + $signed(twiddle_factor_table_59_imag));
  assign _zz_14504 = fixTo_1140_dout;
  assign _zz_14505 = ($signed(_zz_1530) - $signed(_zz_1529));
  assign _zz_14506 = ($signed(_zz_1529) + $signed(_zz_1530));
  assign _zz_14507 = _zz_14508[15 : 0];
  assign _zz_14508 = fixTo_1142_dout;
  assign _zz_14509 = _zz_14510[15 : 0];
  assign _zz_14510 = fixTo_1141_dout;
  assign _zz_14511 = _zz_14512;
  assign _zz_14512 = ($signed(_zz_14513) >>> _zz_3696);
  assign _zz_14513 = _zz_14514;
  assign _zz_14514 = ($signed(_zz_1465) - $signed(_zz_3693));
  assign _zz_14515 = _zz_14516;
  assign _zz_14516 = ($signed(_zz_14517) >>> _zz_3696);
  assign _zz_14517 = _zz_14518;
  assign _zz_14518 = ($signed(_zz_1466) - $signed(_zz_3694));
  assign _zz_14519 = _zz_14520;
  assign _zz_14520 = ($signed(_zz_14521) >>> _zz_3697);
  assign _zz_14521 = _zz_14522;
  assign _zz_14522 = ($signed(_zz_1465) + $signed(_zz_3693));
  assign _zz_14523 = _zz_14524;
  assign _zz_14524 = ($signed(_zz_14525) >>> _zz_3697);
  assign _zz_14525 = _zz_14526;
  assign _zz_14526 = ($signed(_zz_1466) + $signed(_zz_3694));
  assign _zz_14527 = ($signed(twiddle_factor_table_60_real) + $signed(twiddle_factor_table_60_imag));
  assign _zz_14528 = fixTo_1143_dout;
  assign _zz_14529 = ($signed(_zz_1532) - $signed(_zz_1531));
  assign _zz_14530 = ($signed(_zz_1531) + $signed(_zz_1532));
  assign _zz_14531 = _zz_14532[15 : 0];
  assign _zz_14532 = fixTo_1145_dout;
  assign _zz_14533 = _zz_14534[15 : 0];
  assign _zz_14534 = fixTo_1144_dout;
  assign _zz_14535 = _zz_14536;
  assign _zz_14536 = ($signed(_zz_14537) >>> _zz_3701);
  assign _zz_14537 = _zz_14538;
  assign _zz_14538 = ($signed(_zz_1467) - $signed(_zz_3698));
  assign _zz_14539 = _zz_14540;
  assign _zz_14540 = ($signed(_zz_14541) >>> _zz_3701);
  assign _zz_14541 = _zz_14542;
  assign _zz_14542 = ($signed(_zz_1468) - $signed(_zz_3699));
  assign _zz_14543 = _zz_14544;
  assign _zz_14544 = ($signed(_zz_14545) >>> _zz_3702);
  assign _zz_14545 = _zz_14546;
  assign _zz_14546 = ($signed(_zz_1467) + $signed(_zz_3698));
  assign _zz_14547 = _zz_14548;
  assign _zz_14548 = ($signed(_zz_14549) >>> _zz_3702);
  assign _zz_14549 = _zz_14550;
  assign _zz_14550 = ($signed(_zz_1468) + $signed(_zz_3699));
  assign _zz_14551 = ($signed(twiddle_factor_table_61_real) + $signed(twiddle_factor_table_61_imag));
  assign _zz_14552 = fixTo_1146_dout;
  assign _zz_14553 = ($signed(_zz_1534) - $signed(_zz_1533));
  assign _zz_14554 = ($signed(_zz_1533) + $signed(_zz_1534));
  assign _zz_14555 = _zz_14556[15 : 0];
  assign _zz_14556 = fixTo_1148_dout;
  assign _zz_14557 = _zz_14558[15 : 0];
  assign _zz_14558 = fixTo_1147_dout;
  assign _zz_14559 = _zz_14560;
  assign _zz_14560 = ($signed(_zz_14561) >>> _zz_3706);
  assign _zz_14561 = _zz_14562;
  assign _zz_14562 = ($signed(_zz_1469) - $signed(_zz_3703));
  assign _zz_14563 = _zz_14564;
  assign _zz_14564 = ($signed(_zz_14565) >>> _zz_3706);
  assign _zz_14565 = _zz_14566;
  assign _zz_14566 = ($signed(_zz_1470) - $signed(_zz_3704));
  assign _zz_14567 = _zz_14568;
  assign _zz_14568 = ($signed(_zz_14569) >>> _zz_3707);
  assign _zz_14569 = _zz_14570;
  assign _zz_14570 = ($signed(_zz_1469) + $signed(_zz_3703));
  assign _zz_14571 = _zz_14572;
  assign _zz_14572 = ($signed(_zz_14573) >>> _zz_3707);
  assign _zz_14573 = _zz_14574;
  assign _zz_14574 = ($signed(_zz_1470) + $signed(_zz_3704));
  assign _zz_14575 = ($signed(twiddle_factor_table_62_real) + $signed(twiddle_factor_table_62_imag));
  assign _zz_14576 = fixTo_1149_dout;
  assign _zz_14577 = ($signed(_zz_1536) - $signed(_zz_1535));
  assign _zz_14578 = ($signed(_zz_1535) + $signed(_zz_1536));
  assign _zz_14579 = _zz_14580[15 : 0];
  assign _zz_14580 = fixTo_1151_dout;
  assign _zz_14581 = _zz_14582[15 : 0];
  assign _zz_14582 = fixTo_1150_dout;
  assign _zz_14583 = _zz_14584;
  assign _zz_14584 = ($signed(_zz_14585) >>> _zz_3711);
  assign _zz_14585 = _zz_14586;
  assign _zz_14586 = ($signed(_zz_1471) - $signed(_zz_3708));
  assign _zz_14587 = _zz_14588;
  assign _zz_14588 = ($signed(_zz_14589) >>> _zz_3711);
  assign _zz_14589 = _zz_14590;
  assign _zz_14590 = ($signed(_zz_1472) - $signed(_zz_3709));
  assign _zz_14591 = _zz_14592;
  assign _zz_14592 = ($signed(_zz_14593) >>> _zz_3712);
  assign _zz_14593 = _zz_14594;
  assign _zz_14594 = ($signed(_zz_1471) + $signed(_zz_3708));
  assign _zz_14595 = _zz_14596;
  assign _zz_14596 = ($signed(_zz_14597) >>> _zz_3712);
  assign _zz_14597 = _zz_14598;
  assign _zz_14598 = ($signed(_zz_1472) + $signed(_zz_3709));
  assign _zz_14599 = ($signed(twiddle_factor_table_63_real) + $signed(twiddle_factor_table_63_imag));
  assign _zz_14600 = fixTo_1152_dout;
  assign _zz_14601 = ($signed(_zz_1666) - $signed(_zz_1665));
  assign _zz_14602 = ($signed(_zz_1665) + $signed(_zz_1666));
  assign _zz_14603 = _zz_14604[15 : 0];
  assign _zz_14604 = fixTo_1154_dout;
  assign _zz_14605 = _zz_14606[15 : 0];
  assign _zz_14606 = fixTo_1153_dout;
  assign _zz_14607 = _zz_14608;
  assign _zz_14608 = ($signed(_zz_14609) >>> _zz_3716);
  assign _zz_14609 = _zz_14610;
  assign _zz_14610 = ($signed(_zz_1537) - $signed(_zz_3713));
  assign _zz_14611 = _zz_14612;
  assign _zz_14612 = ($signed(_zz_14613) >>> _zz_3716);
  assign _zz_14613 = _zz_14614;
  assign _zz_14614 = ($signed(_zz_1538) - $signed(_zz_3714));
  assign _zz_14615 = _zz_14616;
  assign _zz_14616 = ($signed(_zz_14617) >>> _zz_3717);
  assign _zz_14617 = _zz_14618;
  assign _zz_14618 = ($signed(_zz_1537) + $signed(_zz_3713));
  assign _zz_14619 = _zz_14620;
  assign _zz_14620 = ($signed(_zz_14621) >>> _zz_3717);
  assign _zz_14621 = _zz_14622;
  assign _zz_14622 = ($signed(_zz_1538) + $signed(_zz_3714));
  assign _zz_14623 = ($signed(twiddle_factor_table_64_real) + $signed(twiddle_factor_table_64_imag));
  assign _zz_14624 = fixTo_1155_dout;
  assign _zz_14625 = ($signed(_zz_1668) - $signed(_zz_1667));
  assign _zz_14626 = ($signed(_zz_1667) + $signed(_zz_1668));
  assign _zz_14627 = _zz_14628[15 : 0];
  assign _zz_14628 = fixTo_1157_dout;
  assign _zz_14629 = _zz_14630[15 : 0];
  assign _zz_14630 = fixTo_1156_dout;
  assign _zz_14631 = _zz_14632;
  assign _zz_14632 = ($signed(_zz_14633) >>> _zz_3721);
  assign _zz_14633 = _zz_14634;
  assign _zz_14634 = ($signed(_zz_1539) - $signed(_zz_3718));
  assign _zz_14635 = _zz_14636;
  assign _zz_14636 = ($signed(_zz_14637) >>> _zz_3721);
  assign _zz_14637 = _zz_14638;
  assign _zz_14638 = ($signed(_zz_1540) - $signed(_zz_3719));
  assign _zz_14639 = _zz_14640;
  assign _zz_14640 = ($signed(_zz_14641) >>> _zz_3722);
  assign _zz_14641 = _zz_14642;
  assign _zz_14642 = ($signed(_zz_1539) + $signed(_zz_3718));
  assign _zz_14643 = _zz_14644;
  assign _zz_14644 = ($signed(_zz_14645) >>> _zz_3722);
  assign _zz_14645 = _zz_14646;
  assign _zz_14646 = ($signed(_zz_1540) + $signed(_zz_3719));
  assign _zz_14647 = ($signed(twiddle_factor_table_65_real) + $signed(twiddle_factor_table_65_imag));
  assign _zz_14648 = fixTo_1158_dout;
  assign _zz_14649 = ($signed(_zz_1670) - $signed(_zz_1669));
  assign _zz_14650 = ($signed(_zz_1669) + $signed(_zz_1670));
  assign _zz_14651 = _zz_14652[15 : 0];
  assign _zz_14652 = fixTo_1160_dout;
  assign _zz_14653 = _zz_14654[15 : 0];
  assign _zz_14654 = fixTo_1159_dout;
  assign _zz_14655 = _zz_14656;
  assign _zz_14656 = ($signed(_zz_14657) >>> _zz_3726);
  assign _zz_14657 = _zz_14658;
  assign _zz_14658 = ($signed(_zz_1541) - $signed(_zz_3723));
  assign _zz_14659 = _zz_14660;
  assign _zz_14660 = ($signed(_zz_14661) >>> _zz_3726);
  assign _zz_14661 = _zz_14662;
  assign _zz_14662 = ($signed(_zz_1542) - $signed(_zz_3724));
  assign _zz_14663 = _zz_14664;
  assign _zz_14664 = ($signed(_zz_14665) >>> _zz_3727);
  assign _zz_14665 = _zz_14666;
  assign _zz_14666 = ($signed(_zz_1541) + $signed(_zz_3723));
  assign _zz_14667 = _zz_14668;
  assign _zz_14668 = ($signed(_zz_14669) >>> _zz_3727);
  assign _zz_14669 = _zz_14670;
  assign _zz_14670 = ($signed(_zz_1542) + $signed(_zz_3724));
  assign _zz_14671 = ($signed(twiddle_factor_table_66_real) + $signed(twiddle_factor_table_66_imag));
  assign _zz_14672 = fixTo_1161_dout;
  assign _zz_14673 = ($signed(_zz_1672) - $signed(_zz_1671));
  assign _zz_14674 = ($signed(_zz_1671) + $signed(_zz_1672));
  assign _zz_14675 = _zz_14676[15 : 0];
  assign _zz_14676 = fixTo_1163_dout;
  assign _zz_14677 = _zz_14678[15 : 0];
  assign _zz_14678 = fixTo_1162_dout;
  assign _zz_14679 = _zz_14680;
  assign _zz_14680 = ($signed(_zz_14681) >>> _zz_3731);
  assign _zz_14681 = _zz_14682;
  assign _zz_14682 = ($signed(_zz_1543) - $signed(_zz_3728));
  assign _zz_14683 = _zz_14684;
  assign _zz_14684 = ($signed(_zz_14685) >>> _zz_3731);
  assign _zz_14685 = _zz_14686;
  assign _zz_14686 = ($signed(_zz_1544) - $signed(_zz_3729));
  assign _zz_14687 = _zz_14688;
  assign _zz_14688 = ($signed(_zz_14689) >>> _zz_3732);
  assign _zz_14689 = _zz_14690;
  assign _zz_14690 = ($signed(_zz_1543) + $signed(_zz_3728));
  assign _zz_14691 = _zz_14692;
  assign _zz_14692 = ($signed(_zz_14693) >>> _zz_3732);
  assign _zz_14693 = _zz_14694;
  assign _zz_14694 = ($signed(_zz_1544) + $signed(_zz_3729));
  assign _zz_14695 = ($signed(twiddle_factor_table_67_real) + $signed(twiddle_factor_table_67_imag));
  assign _zz_14696 = fixTo_1164_dout;
  assign _zz_14697 = ($signed(_zz_1674) - $signed(_zz_1673));
  assign _zz_14698 = ($signed(_zz_1673) + $signed(_zz_1674));
  assign _zz_14699 = _zz_14700[15 : 0];
  assign _zz_14700 = fixTo_1166_dout;
  assign _zz_14701 = _zz_14702[15 : 0];
  assign _zz_14702 = fixTo_1165_dout;
  assign _zz_14703 = _zz_14704;
  assign _zz_14704 = ($signed(_zz_14705) >>> _zz_3736);
  assign _zz_14705 = _zz_14706;
  assign _zz_14706 = ($signed(_zz_1545) - $signed(_zz_3733));
  assign _zz_14707 = _zz_14708;
  assign _zz_14708 = ($signed(_zz_14709) >>> _zz_3736);
  assign _zz_14709 = _zz_14710;
  assign _zz_14710 = ($signed(_zz_1546) - $signed(_zz_3734));
  assign _zz_14711 = _zz_14712;
  assign _zz_14712 = ($signed(_zz_14713) >>> _zz_3737);
  assign _zz_14713 = _zz_14714;
  assign _zz_14714 = ($signed(_zz_1545) + $signed(_zz_3733));
  assign _zz_14715 = _zz_14716;
  assign _zz_14716 = ($signed(_zz_14717) >>> _zz_3737);
  assign _zz_14717 = _zz_14718;
  assign _zz_14718 = ($signed(_zz_1546) + $signed(_zz_3734));
  assign _zz_14719 = ($signed(twiddle_factor_table_68_real) + $signed(twiddle_factor_table_68_imag));
  assign _zz_14720 = fixTo_1167_dout;
  assign _zz_14721 = ($signed(_zz_1676) - $signed(_zz_1675));
  assign _zz_14722 = ($signed(_zz_1675) + $signed(_zz_1676));
  assign _zz_14723 = _zz_14724[15 : 0];
  assign _zz_14724 = fixTo_1169_dout;
  assign _zz_14725 = _zz_14726[15 : 0];
  assign _zz_14726 = fixTo_1168_dout;
  assign _zz_14727 = _zz_14728;
  assign _zz_14728 = ($signed(_zz_14729) >>> _zz_3741);
  assign _zz_14729 = _zz_14730;
  assign _zz_14730 = ($signed(_zz_1547) - $signed(_zz_3738));
  assign _zz_14731 = _zz_14732;
  assign _zz_14732 = ($signed(_zz_14733) >>> _zz_3741);
  assign _zz_14733 = _zz_14734;
  assign _zz_14734 = ($signed(_zz_1548) - $signed(_zz_3739));
  assign _zz_14735 = _zz_14736;
  assign _zz_14736 = ($signed(_zz_14737) >>> _zz_3742);
  assign _zz_14737 = _zz_14738;
  assign _zz_14738 = ($signed(_zz_1547) + $signed(_zz_3738));
  assign _zz_14739 = _zz_14740;
  assign _zz_14740 = ($signed(_zz_14741) >>> _zz_3742);
  assign _zz_14741 = _zz_14742;
  assign _zz_14742 = ($signed(_zz_1548) + $signed(_zz_3739));
  assign _zz_14743 = ($signed(twiddle_factor_table_69_real) + $signed(twiddle_factor_table_69_imag));
  assign _zz_14744 = fixTo_1170_dout;
  assign _zz_14745 = ($signed(_zz_1678) - $signed(_zz_1677));
  assign _zz_14746 = ($signed(_zz_1677) + $signed(_zz_1678));
  assign _zz_14747 = _zz_14748[15 : 0];
  assign _zz_14748 = fixTo_1172_dout;
  assign _zz_14749 = _zz_14750[15 : 0];
  assign _zz_14750 = fixTo_1171_dout;
  assign _zz_14751 = _zz_14752;
  assign _zz_14752 = ($signed(_zz_14753) >>> _zz_3746);
  assign _zz_14753 = _zz_14754;
  assign _zz_14754 = ($signed(_zz_1549) - $signed(_zz_3743));
  assign _zz_14755 = _zz_14756;
  assign _zz_14756 = ($signed(_zz_14757) >>> _zz_3746);
  assign _zz_14757 = _zz_14758;
  assign _zz_14758 = ($signed(_zz_1550) - $signed(_zz_3744));
  assign _zz_14759 = _zz_14760;
  assign _zz_14760 = ($signed(_zz_14761) >>> _zz_3747);
  assign _zz_14761 = _zz_14762;
  assign _zz_14762 = ($signed(_zz_1549) + $signed(_zz_3743));
  assign _zz_14763 = _zz_14764;
  assign _zz_14764 = ($signed(_zz_14765) >>> _zz_3747);
  assign _zz_14765 = _zz_14766;
  assign _zz_14766 = ($signed(_zz_1550) + $signed(_zz_3744));
  assign _zz_14767 = ($signed(twiddle_factor_table_70_real) + $signed(twiddle_factor_table_70_imag));
  assign _zz_14768 = fixTo_1173_dout;
  assign _zz_14769 = ($signed(_zz_1680) - $signed(_zz_1679));
  assign _zz_14770 = ($signed(_zz_1679) + $signed(_zz_1680));
  assign _zz_14771 = _zz_14772[15 : 0];
  assign _zz_14772 = fixTo_1175_dout;
  assign _zz_14773 = _zz_14774[15 : 0];
  assign _zz_14774 = fixTo_1174_dout;
  assign _zz_14775 = _zz_14776;
  assign _zz_14776 = ($signed(_zz_14777) >>> _zz_3751);
  assign _zz_14777 = _zz_14778;
  assign _zz_14778 = ($signed(_zz_1551) - $signed(_zz_3748));
  assign _zz_14779 = _zz_14780;
  assign _zz_14780 = ($signed(_zz_14781) >>> _zz_3751);
  assign _zz_14781 = _zz_14782;
  assign _zz_14782 = ($signed(_zz_1552) - $signed(_zz_3749));
  assign _zz_14783 = _zz_14784;
  assign _zz_14784 = ($signed(_zz_14785) >>> _zz_3752);
  assign _zz_14785 = _zz_14786;
  assign _zz_14786 = ($signed(_zz_1551) + $signed(_zz_3748));
  assign _zz_14787 = _zz_14788;
  assign _zz_14788 = ($signed(_zz_14789) >>> _zz_3752);
  assign _zz_14789 = _zz_14790;
  assign _zz_14790 = ($signed(_zz_1552) + $signed(_zz_3749));
  assign _zz_14791 = ($signed(twiddle_factor_table_71_real) + $signed(twiddle_factor_table_71_imag));
  assign _zz_14792 = fixTo_1176_dout;
  assign _zz_14793 = ($signed(_zz_1682) - $signed(_zz_1681));
  assign _zz_14794 = ($signed(_zz_1681) + $signed(_zz_1682));
  assign _zz_14795 = _zz_14796[15 : 0];
  assign _zz_14796 = fixTo_1178_dout;
  assign _zz_14797 = _zz_14798[15 : 0];
  assign _zz_14798 = fixTo_1177_dout;
  assign _zz_14799 = _zz_14800;
  assign _zz_14800 = ($signed(_zz_14801) >>> _zz_3756);
  assign _zz_14801 = _zz_14802;
  assign _zz_14802 = ($signed(_zz_1553) - $signed(_zz_3753));
  assign _zz_14803 = _zz_14804;
  assign _zz_14804 = ($signed(_zz_14805) >>> _zz_3756);
  assign _zz_14805 = _zz_14806;
  assign _zz_14806 = ($signed(_zz_1554) - $signed(_zz_3754));
  assign _zz_14807 = _zz_14808;
  assign _zz_14808 = ($signed(_zz_14809) >>> _zz_3757);
  assign _zz_14809 = _zz_14810;
  assign _zz_14810 = ($signed(_zz_1553) + $signed(_zz_3753));
  assign _zz_14811 = _zz_14812;
  assign _zz_14812 = ($signed(_zz_14813) >>> _zz_3757);
  assign _zz_14813 = _zz_14814;
  assign _zz_14814 = ($signed(_zz_1554) + $signed(_zz_3754));
  assign _zz_14815 = ($signed(twiddle_factor_table_72_real) + $signed(twiddle_factor_table_72_imag));
  assign _zz_14816 = fixTo_1179_dout;
  assign _zz_14817 = ($signed(_zz_1684) - $signed(_zz_1683));
  assign _zz_14818 = ($signed(_zz_1683) + $signed(_zz_1684));
  assign _zz_14819 = _zz_14820[15 : 0];
  assign _zz_14820 = fixTo_1181_dout;
  assign _zz_14821 = _zz_14822[15 : 0];
  assign _zz_14822 = fixTo_1180_dout;
  assign _zz_14823 = _zz_14824;
  assign _zz_14824 = ($signed(_zz_14825) >>> _zz_3761);
  assign _zz_14825 = _zz_14826;
  assign _zz_14826 = ($signed(_zz_1555) - $signed(_zz_3758));
  assign _zz_14827 = _zz_14828;
  assign _zz_14828 = ($signed(_zz_14829) >>> _zz_3761);
  assign _zz_14829 = _zz_14830;
  assign _zz_14830 = ($signed(_zz_1556) - $signed(_zz_3759));
  assign _zz_14831 = _zz_14832;
  assign _zz_14832 = ($signed(_zz_14833) >>> _zz_3762);
  assign _zz_14833 = _zz_14834;
  assign _zz_14834 = ($signed(_zz_1555) + $signed(_zz_3758));
  assign _zz_14835 = _zz_14836;
  assign _zz_14836 = ($signed(_zz_14837) >>> _zz_3762);
  assign _zz_14837 = _zz_14838;
  assign _zz_14838 = ($signed(_zz_1556) + $signed(_zz_3759));
  assign _zz_14839 = ($signed(twiddle_factor_table_73_real) + $signed(twiddle_factor_table_73_imag));
  assign _zz_14840 = fixTo_1182_dout;
  assign _zz_14841 = ($signed(_zz_1686) - $signed(_zz_1685));
  assign _zz_14842 = ($signed(_zz_1685) + $signed(_zz_1686));
  assign _zz_14843 = _zz_14844[15 : 0];
  assign _zz_14844 = fixTo_1184_dout;
  assign _zz_14845 = _zz_14846[15 : 0];
  assign _zz_14846 = fixTo_1183_dout;
  assign _zz_14847 = _zz_14848;
  assign _zz_14848 = ($signed(_zz_14849) >>> _zz_3766);
  assign _zz_14849 = _zz_14850;
  assign _zz_14850 = ($signed(_zz_1557) - $signed(_zz_3763));
  assign _zz_14851 = _zz_14852;
  assign _zz_14852 = ($signed(_zz_14853) >>> _zz_3766);
  assign _zz_14853 = _zz_14854;
  assign _zz_14854 = ($signed(_zz_1558) - $signed(_zz_3764));
  assign _zz_14855 = _zz_14856;
  assign _zz_14856 = ($signed(_zz_14857) >>> _zz_3767);
  assign _zz_14857 = _zz_14858;
  assign _zz_14858 = ($signed(_zz_1557) + $signed(_zz_3763));
  assign _zz_14859 = _zz_14860;
  assign _zz_14860 = ($signed(_zz_14861) >>> _zz_3767);
  assign _zz_14861 = _zz_14862;
  assign _zz_14862 = ($signed(_zz_1558) + $signed(_zz_3764));
  assign _zz_14863 = ($signed(twiddle_factor_table_74_real) + $signed(twiddle_factor_table_74_imag));
  assign _zz_14864 = fixTo_1185_dout;
  assign _zz_14865 = ($signed(_zz_1688) - $signed(_zz_1687));
  assign _zz_14866 = ($signed(_zz_1687) + $signed(_zz_1688));
  assign _zz_14867 = _zz_14868[15 : 0];
  assign _zz_14868 = fixTo_1187_dout;
  assign _zz_14869 = _zz_14870[15 : 0];
  assign _zz_14870 = fixTo_1186_dout;
  assign _zz_14871 = _zz_14872;
  assign _zz_14872 = ($signed(_zz_14873) >>> _zz_3771);
  assign _zz_14873 = _zz_14874;
  assign _zz_14874 = ($signed(_zz_1559) - $signed(_zz_3768));
  assign _zz_14875 = _zz_14876;
  assign _zz_14876 = ($signed(_zz_14877) >>> _zz_3771);
  assign _zz_14877 = _zz_14878;
  assign _zz_14878 = ($signed(_zz_1560) - $signed(_zz_3769));
  assign _zz_14879 = _zz_14880;
  assign _zz_14880 = ($signed(_zz_14881) >>> _zz_3772);
  assign _zz_14881 = _zz_14882;
  assign _zz_14882 = ($signed(_zz_1559) + $signed(_zz_3768));
  assign _zz_14883 = _zz_14884;
  assign _zz_14884 = ($signed(_zz_14885) >>> _zz_3772);
  assign _zz_14885 = _zz_14886;
  assign _zz_14886 = ($signed(_zz_1560) + $signed(_zz_3769));
  assign _zz_14887 = ($signed(twiddle_factor_table_75_real) + $signed(twiddle_factor_table_75_imag));
  assign _zz_14888 = fixTo_1188_dout;
  assign _zz_14889 = ($signed(_zz_1690) - $signed(_zz_1689));
  assign _zz_14890 = ($signed(_zz_1689) + $signed(_zz_1690));
  assign _zz_14891 = _zz_14892[15 : 0];
  assign _zz_14892 = fixTo_1190_dout;
  assign _zz_14893 = _zz_14894[15 : 0];
  assign _zz_14894 = fixTo_1189_dout;
  assign _zz_14895 = _zz_14896;
  assign _zz_14896 = ($signed(_zz_14897) >>> _zz_3776);
  assign _zz_14897 = _zz_14898;
  assign _zz_14898 = ($signed(_zz_1561) - $signed(_zz_3773));
  assign _zz_14899 = _zz_14900;
  assign _zz_14900 = ($signed(_zz_14901) >>> _zz_3776);
  assign _zz_14901 = _zz_14902;
  assign _zz_14902 = ($signed(_zz_1562) - $signed(_zz_3774));
  assign _zz_14903 = _zz_14904;
  assign _zz_14904 = ($signed(_zz_14905) >>> _zz_3777);
  assign _zz_14905 = _zz_14906;
  assign _zz_14906 = ($signed(_zz_1561) + $signed(_zz_3773));
  assign _zz_14907 = _zz_14908;
  assign _zz_14908 = ($signed(_zz_14909) >>> _zz_3777);
  assign _zz_14909 = _zz_14910;
  assign _zz_14910 = ($signed(_zz_1562) + $signed(_zz_3774));
  assign _zz_14911 = ($signed(twiddle_factor_table_76_real) + $signed(twiddle_factor_table_76_imag));
  assign _zz_14912 = fixTo_1191_dout;
  assign _zz_14913 = ($signed(_zz_1692) - $signed(_zz_1691));
  assign _zz_14914 = ($signed(_zz_1691) + $signed(_zz_1692));
  assign _zz_14915 = _zz_14916[15 : 0];
  assign _zz_14916 = fixTo_1193_dout;
  assign _zz_14917 = _zz_14918[15 : 0];
  assign _zz_14918 = fixTo_1192_dout;
  assign _zz_14919 = _zz_14920;
  assign _zz_14920 = ($signed(_zz_14921) >>> _zz_3781);
  assign _zz_14921 = _zz_14922;
  assign _zz_14922 = ($signed(_zz_1563) - $signed(_zz_3778));
  assign _zz_14923 = _zz_14924;
  assign _zz_14924 = ($signed(_zz_14925) >>> _zz_3781);
  assign _zz_14925 = _zz_14926;
  assign _zz_14926 = ($signed(_zz_1564) - $signed(_zz_3779));
  assign _zz_14927 = _zz_14928;
  assign _zz_14928 = ($signed(_zz_14929) >>> _zz_3782);
  assign _zz_14929 = _zz_14930;
  assign _zz_14930 = ($signed(_zz_1563) + $signed(_zz_3778));
  assign _zz_14931 = _zz_14932;
  assign _zz_14932 = ($signed(_zz_14933) >>> _zz_3782);
  assign _zz_14933 = _zz_14934;
  assign _zz_14934 = ($signed(_zz_1564) + $signed(_zz_3779));
  assign _zz_14935 = ($signed(twiddle_factor_table_77_real) + $signed(twiddle_factor_table_77_imag));
  assign _zz_14936 = fixTo_1194_dout;
  assign _zz_14937 = ($signed(_zz_1694) - $signed(_zz_1693));
  assign _zz_14938 = ($signed(_zz_1693) + $signed(_zz_1694));
  assign _zz_14939 = _zz_14940[15 : 0];
  assign _zz_14940 = fixTo_1196_dout;
  assign _zz_14941 = _zz_14942[15 : 0];
  assign _zz_14942 = fixTo_1195_dout;
  assign _zz_14943 = _zz_14944;
  assign _zz_14944 = ($signed(_zz_14945) >>> _zz_3786);
  assign _zz_14945 = _zz_14946;
  assign _zz_14946 = ($signed(_zz_1565) - $signed(_zz_3783));
  assign _zz_14947 = _zz_14948;
  assign _zz_14948 = ($signed(_zz_14949) >>> _zz_3786);
  assign _zz_14949 = _zz_14950;
  assign _zz_14950 = ($signed(_zz_1566) - $signed(_zz_3784));
  assign _zz_14951 = _zz_14952;
  assign _zz_14952 = ($signed(_zz_14953) >>> _zz_3787);
  assign _zz_14953 = _zz_14954;
  assign _zz_14954 = ($signed(_zz_1565) + $signed(_zz_3783));
  assign _zz_14955 = _zz_14956;
  assign _zz_14956 = ($signed(_zz_14957) >>> _zz_3787);
  assign _zz_14957 = _zz_14958;
  assign _zz_14958 = ($signed(_zz_1566) + $signed(_zz_3784));
  assign _zz_14959 = ($signed(twiddle_factor_table_78_real) + $signed(twiddle_factor_table_78_imag));
  assign _zz_14960 = fixTo_1197_dout;
  assign _zz_14961 = ($signed(_zz_1696) - $signed(_zz_1695));
  assign _zz_14962 = ($signed(_zz_1695) + $signed(_zz_1696));
  assign _zz_14963 = _zz_14964[15 : 0];
  assign _zz_14964 = fixTo_1199_dout;
  assign _zz_14965 = _zz_14966[15 : 0];
  assign _zz_14966 = fixTo_1198_dout;
  assign _zz_14967 = _zz_14968;
  assign _zz_14968 = ($signed(_zz_14969) >>> _zz_3791);
  assign _zz_14969 = _zz_14970;
  assign _zz_14970 = ($signed(_zz_1567) - $signed(_zz_3788));
  assign _zz_14971 = _zz_14972;
  assign _zz_14972 = ($signed(_zz_14973) >>> _zz_3791);
  assign _zz_14973 = _zz_14974;
  assign _zz_14974 = ($signed(_zz_1568) - $signed(_zz_3789));
  assign _zz_14975 = _zz_14976;
  assign _zz_14976 = ($signed(_zz_14977) >>> _zz_3792);
  assign _zz_14977 = _zz_14978;
  assign _zz_14978 = ($signed(_zz_1567) + $signed(_zz_3788));
  assign _zz_14979 = _zz_14980;
  assign _zz_14980 = ($signed(_zz_14981) >>> _zz_3792);
  assign _zz_14981 = _zz_14982;
  assign _zz_14982 = ($signed(_zz_1568) + $signed(_zz_3789));
  assign _zz_14983 = ($signed(twiddle_factor_table_79_real) + $signed(twiddle_factor_table_79_imag));
  assign _zz_14984 = fixTo_1200_dout;
  assign _zz_14985 = ($signed(_zz_1698) - $signed(_zz_1697));
  assign _zz_14986 = ($signed(_zz_1697) + $signed(_zz_1698));
  assign _zz_14987 = _zz_14988[15 : 0];
  assign _zz_14988 = fixTo_1202_dout;
  assign _zz_14989 = _zz_14990[15 : 0];
  assign _zz_14990 = fixTo_1201_dout;
  assign _zz_14991 = _zz_14992;
  assign _zz_14992 = ($signed(_zz_14993) >>> _zz_3796);
  assign _zz_14993 = _zz_14994;
  assign _zz_14994 = ($signed(_zz_1569) - $signed(_zz_3793));
  assign _zz_14995 = _zz_14996;
  assign _zz_14996 = ($signed(_zz_14997) >>> _zz_3796);
  assign _zz_14997 = _zz_14998;
  assign _zz_14998 = ($signed(_zz_1570) - $signed(_zz_3794));
  assign _zz_14999 = _zz_15000;
  assign _zz_15000 = ($signed(_zz_15001) >>> _zz_3797);
  assign _zz_15001 = _zz_15002;
  assign _zz_15002 = ($signed(_zz_1569) + $signed(_zz_3793));
  assign _zz_15003 = _zz_15004;
  assign _zz_15004 = ($signed(_zz_15005) >>> _zz_3797);
  assign _zz_15005 = _zz_15006;
  assign _zz_15006 = ($signed(_zz_1570) + $signed(_zz_3794));
  assign _zz_15007 = ($signed(twiddle_factor_table_80_real) + $signed(twiddle_factor_table_80_imag));
  assign _zz_15008 = fixTo_1203_dout;
  assign _zz_15009 = ($signed(_zz_1700) - $signed(_zz_1699));
  assign _zz_15010 = ($signed(_zz_1699) + $signed(_zz_1700));
  assign _zz_15011 = _zz_15012[15 : 0];
  assign _zz_15012 = fixTo_1205_dout;
  assign _zz_15013 = _zz_15014[15 : 0];
  assign _zz_15014 = fixTo_1204_dout;
  assign _zz_15015 = _zz_15016;
  assign _zz_15016 = ($signed(_zz_15017) >>> _zz_3801);
  assign _zz_15017 = _zz_15018;
  assign _zz_15018 = ($signed(_zz_1571) - $signed(_zz_3798));
  assign _zz_15019 = _zz_15020;
  assign _zz_15020 = ($signed(_zz_15021) >>> _zz_3801);
  assign _zz_15021 = _zz_15022;
  assign _zz_15022 = ($signed(_zz_1572) - $signed(_zz_3799));
  assign _zz_15023 = _zz_15024;
  assign _zz_15024 = ($signed(_zz_15025) >>> _zz_3802);
  assign _zz_15025 = _zz_15026;
  assign _zz_15026 = ($signed(_zz_1571) + $signed(_zz_3798));
  assign _zz_15027 = _zz_15028;
  assign _zz_15028 = ($signed(_zz_15029) >>> _zz_3802);
  assign _zz_15029 = _zz_15030;
  assign _zz_15030 = ($signed(_zz_1572) + $signed(_zz_3799));
  assign _zz_15031 = ($signed(twiddle_factor_table_81_real) + $signed(twiddle_factor_table_81_imag));
  assign _zz_15032 = fixTo_1206_dout;
  assign _zz_15033 = ($signed(_zz_1702) - $signed(_zz_1701));
  assign _zz_15034 = ($signed(_zz_1701) + $signed(_zz_1702));
  assign _zz_15035 = _zz_15036[15 : 0];
  assign _zz_15036 = fixTo_1208_dout;
  assign _zz_15037 = _zz_15038[15 : 0];
  assign _zz_15038 = fixTo_1207_dout;
  assign _zz_15039 = _zz_15040;
  assign _zz_15040 = ($signed(_zz_15041) >>> _zz_3806);
  assign _zz_15041 = _zz_15042;
  assign _zz_15042 = ($signed(_zz_1573) - $signed(_zz_3803));
  assign _zz_15043 = _zz_15044;
  assign _zz_15044 = ($signed(_zz_15045) >>> _zz_3806);
  assign _zz_15045 = _zz_15046;
  assign _zz_15046 = ($signed(_zz_1574) - $signed(_zz_3804));
  assign _zz_15047 = _zz_15048;
  assign _zz_15048 = ($signed(_zz_15049) >>> _zz_3807);
  assign _zz_15049 = _zz_15050;
  assign _zz_15050 = ($signed(_zz_1573) + $signed(_zz_3803));
  assign _zz_15051 = _zz_15052;
  assign _zz_15052 = ($signed(_zz_15053) >>> _zz_3807);
  assign _zz_15053 = _zz_15054;
  assign _zz_15054 = ($signed(_zz_1574) + $signed(_zz_3804));
  assign _zz_15055 = ($signed(twiddle_factor_table_82_real) + $signed(twiddle_factor_table_82_imag));
  assign _zz_15056 = fixTo_1209_dout;
  assign _zz_15057 = ($signed(_zz_1704) - $signed(_zz_1703));
  assign _zz_15058 = ($signed(_zz_1703) + $signed(_zz_1704));
  assign _zz_15059 = _zz_15060[15 : 0];
  assign _zz_15060 = fixTo_1211_dout;
  assign _zz_15061 = _zz_15062[15 : 0];
  assign _zz_15062 = fixTo_1210_dout;
  assign _zz_15063 = _zz_15064;
  assign _zz_15064 = ($signed(_zz_15065) >>> _zz_3811);
  assign _zz_15065 = _zz_15066;
  assign _zz_15066 = ($signed(_zz_1575) - $signed(_zz_3808));
  assign _zz_15067 = _zz_15068;
  assign _zz_15068 = ($signed(_zz_15069) >>> _zz_3811);
  assign _zz_15069 = _zz_15070;
  assign _zz_15070 = ($signed(_zz_1576) - $signed(_zz_3809));
  assign _zz_15071 = _zz_15072;
  assign _zz_15072 = ($signed(_zz_15073) >>> _zz_3812);
  assign _zz_15073 = _zz_15074;
  assign _zz_15074 = ($signed(_zz_1575) + $signed(_zz_3808));
  assign _zz_15075 = _zz_15076;
  assign _zz_15076 = ($signed(_zz_15077) >>> _zz_3812);
  assign _zz_15077 = _zz_15078;
  assign _zz_15078 = ($signed(_zz_1576) + $signed(_zz_3809));
  assign _zz_15079 = ($signed(twiddle_factor_table_83_real) + $signed(twiddle_factor_table_83_imag));
  assign _zz_15080 = fixTo_1212_dout;
  assign _zz_15081 = ($signed(_zz_1706) - $signed(_zz_1705));
  assign _zz_15082 = ($signed(_zz_1705) + $signed(_zz_1706));
  assign _zz_15083 = _zz_15084[15 : 0];
  assign _zz_15084 = fixTo_1214_dout;
  assign _zz_15085 = _zz_15086[15 : 0];
  assign _zz_15086 = fixTo_1213_dout;
  assign _zz_15087 = _zz_15088;
  assign _zz_15088 = ($signed(_zz_15089) >>> _zz_3816);
  assign _zz_15089 = _zz_15090;
  assign _zz_15090 = ($signed(_zz_1577) - $signed(_zz_3813));
  assign _zz_15091 = _zz_15092;
  assign _zz_15092 = ($signed(_zz_15093) >>> _zz_3816);
  assign _zz_15093 = _zz_15094;
  assign _zz_15094 = ($signed(_zz_1578) - $signed(_zz_3814));
  assign _zz_15095 = _zz_15096;
  assign _zz_15096 = ($signed(_zz_15097) >>> _zz_3817);
  assign _zz_15097 = _zz_15098;
  assign _zz_15098 = ($signed(_zz_1577) + $signed(_zz_3813));
  assign _zz_15099 = _zz_15100;
  assign _zz_15100 = ($signed(_zz_15101) >>> _zz_3817);
  assign _zz_15101 = _zz_15102;
  assign _zz_15102 = ($signed(_zz_1578) + $signed(_zz_3814));
  assign _zz_15103 = ($signed(twiddle_factor_table_84_real) + $signed(twiddle_factor_table_84_imag));
  assign _zz_15104 = fixTo_1215_dout;
  assign _zz_15105 = ($signed(_zz_1708) - $signed(_zz_1707));
  assign _zz_15106 = ($signed(_zz_1707) + $signed(_zz_1708));
  assign _zz_15107 = _zz_15108[15 : 0];
  assign _zz_15108 = fixTo_1217_dout;
  assign _zz_15109 = _zz_15110[15 : 0];
  assign _zz_15110 = fixTo_1216_dout;
  assign _zz_15111 = _zz_15112;
  assign _zz_15112 = ($signed(_zz_15113) >>> _zz_3821);
  assign _zz_15113 = _zz_15114;
  assign _zz_15114 = ($signed(_zz_1579) - $signed(_zz_3818));
  assign _zz_15115 = _zz_15116;
  assign _zz_15116 = ($signed(_zz_15117) >>> _zz_3821);
  assign _zz_15117 = _zz_15118;
  assign _zz_15118 = ($signed(_zz_1580) - $signed(_zz_3819));
  assign _zz_15119 = _zz_15120;
  assign _zz_15120 = ($signed(_zz_15121) >>> _zz_3822);
  assign _zz_15121 = _zz_15122;
  assign _zz_15122 = ($signed(_zz_1579) + $signed(_zz_3818));
  assign _zz_15123 = _zz_15124;
  assign _zz_15124 = ($signed(_zz_15125) >>> _zz_3822);
  assign _zz_15125 = _zz_15126;
  assign _zz_15126 = ($signed(_zz_1580) + $signed(_zz_3819));
  assign _zz_15127 = ($signed(twiddle_factor_table_85_real) + $signed(twiddle_factor_table_85_imag));
  assign _zz_15128 = fixTo_1218_dout;
  assign _zz_15129 = ($signed(_zz_1710) - $signed(_zz_1709));
  assign _zz_15130 = ($signed(_zz_1709) + $signed(_zz_1710));
  assign _zz_15131 = _zz_15132[15 : 0];
  assign _zz_15132 = fixTo_1220_dout;
  assign _zz_15133 = _zz_15134[15 : 0];
  assign _zz_15134 = fixTo_1219_dout;
  assign _zz_15135 = _zz_15136;
  assign _zz_15136 = ($signed(_zz_15137) >>> _zz_3826);
  assign _zz_15137 = _zz_15138;
  assign _zz_15138 = ($signed(_zz_1581) - $signed(_zz_3823));
  assign _zz_15139 = _zz_15140;
  assign _zz_15140 = ($signed(_zz_15141) >>> _zz_3826);
  assign _zz_15141 = _zz_15142;
  assign _zz_15142 = ($signed(_zz_1582) - $signed(_zz_3824));
  assign _zz_15143 = _zz_15144;
  assign _zz_15144 = ($signed(_zz_15145) >>> _zz_3827);
  assign _zz_15145 = _zz_15146;
  assign _zz_15146 = ($signed(_zz_1581) + $signed(_zz_3823));
  assign _zz_15147 = _zz_15148;
  assign _zz_15148 = ($signed(_zz_15149) >>> _zz_3827);
  assign _zz_15149 = _zz_15150;
  assign _zz_15150 = ($signed(_zz_1582) + $signed(_zz_3824));
  assign _zz_15151 = ($signed(twiddle_factor_table_86_real) + $signed(twiddle_factor_table_86_imag));
  assign _zz_15152 = fixTo_1221_dout;
  assign _zz_15153 = ($signed(_zz_1712) - $signed(_zz_1711));
  assign _zz_15154 = ($signed(_zz_1711) + $signed(_zz_1712));
  assign _zz_15155 = _zz_15156[15 : 0];
  assign _zz_15156 = fixTo_1223_dout;
  assign _zz_15157 = _zz_15158[15 : 0];
  assign _zz_15158 = fixTo_1222_dout;
  assign _zz_15159 = _zz_15160;
  assign _zz_15160 = ($signed(_zz_15161) >>> _zz_3831);
  assign _zz_15161 = _zz_15162;
  assign _zz_15162 = ($signed(_zz_1583) - $signed(_zz_3828));
  assign _zz_15163 = _zz_15164;
  assign _zz_15164 = ($signed(_zz_15165) >>> _zz_3831);
  assign _zz_15165 = _zz_15166;
  assign _zz_15166 = ($signed(_zz_1584) - $signed(_zz_3829));
  assign _zz_15167 = _zz_15168;
  assign _zz_15168 = ($signed(_zz_15169) >>> _zz_3832);
  assign _zz_15169 = _zz_15170;
  assign _zz_15170 = ($signed(_zz_1583) + $signed(_zz_3828));
  assign _zz_15171 = _zz_15172;
  assign _zz_15172 = ($signed(_zz_15173) >>> _zz_3832);
  assign _zz_15173 = _zz_15174;
  assign _zz_15174 = ($signed(_zz_1584) + $signed(_zz_3829));
  assign _zz_15175 = ($signed(twiddle_factor_table_87_real) + $signed(twiddle_factor_table_87_imag));
  assign _zz_15176 = fixTo_1224_dout;
  assign _zz_15177 = ($signed(_zz_1714) - $signed(_zz_1713));
  assign _zz_15178 = ($signed(_zz_1713) + $signed(_zz_1714));
  assign _zz_15179 = _zz_15180[15 : 0];
  assign _zz_15180 = fixTo_1226_dout;
  assign _zz_15181 = _zz_15182[15 : 0];
  assign _zz_15182 = fixTo_1225_dout;
  assign _zz_15183 = _zz_15184;
  assign _zz_15184 = ($signed(_zz_15185) >>> _zz_3836);
  assign _zz_15185 = _zz_15186;
  assign _zz_15186 = ($signed(_zz_1585) - $signed(_zz_3833));
  assign _zz_15187 = _zz_15188;
  assign _zz_15188 = ($signed(_zz_15189) >>> _zz_3836);
  assign _zz_15189 = _zz_15190;
  assign _zz_15190 = ($signed(_zz_1586) - $signed(_zz_3834));
  assign _zz_15191 = _zz_15192;
  assign _zz_15192 = ($signed(_zz_15193) >>> _zz_3837);
  assign _zz_15193 = _zz_15194;
  assign _zz_15194 = ($signed(_zz_1585) + $signed(_zz_3833));
  assign _zz_15195 = _zz_15196;
  assign _zz_15196 = ($signed(_zz_15197) >>> _zz_3837);
  assign _zz_15197 = _zz_15198;
  assign _zz_15198 = ($signed(_zz_1586) + $signed(_zz_3834));
  assign _zz_15199 = ($signed(twiddle_factor_table_88_real) + $signed(twiddle_factor_table_88_imag));
  assign _zz_15200 = fixTo_1227_dout;
  assign _zz_15201 = ($signed(_zz_1716) - $signed(_zz_1715));
  assign _zz_15202 = ($signed(_zz_1715) + $signed(_zz_1716));
  assign _zz_15203 = _zz_15204[15 : 0];
  assign _zz_15204 = fixTo_1229_dout;
  assign _zz_15205 = _zz_15206[15 : 0];
  assign _zz_15206 = fixTo_1228_dout;
  assign _zz_15207 = _zz_15208;
  assign _zz_15208 = ($signed(_zz_15209) >>> _zz_3841);
  assign _zz_15209 = _zz_15210;
  assign _zz_15210 = ($signed(_zz_1587) - $signed(_zz_3838));
  assign _zz_15211 = _zz_15212;
  assign _zz_15212 = ($signed(_zz_15213) >>> _zz_3841);
  assign _zz_15213 = _zz_15214;
  assign _zz_15214 = ($signed(_zz_1588) - $signed(_zz_3839));
  assign _zz_15215 = _zz_15216;
  assign _zz_15216 = ($signed(_zz_15217) >>> _zz_3842);
  assign _zz_15217 = _zz_15218;
  assign _zz_15218 = ($signed(_zz_1587) + $signed(_zz_3838));
  assign _zz_15219 = _zz_15220;
  assign _zz_15220 = ($signed(_zz_15221) >>> _zz_3842);
  assign _zz_15221 = _zz_15222;
  assign _zz_15222 = ($signed(_zz_1588) + $signed(_zz_3839));
  assign _zz_15223 = ($signed(twiddle_factor_table_89_real) + $signed(twiddle_factor_table_89_imag));
  assign _zz_15224 = fixTo_1230_dout;
  assign _zz_15225 = ($signed(_zz_1718) - $signed(_zz_1717));
  assign _zz_15226 = ($signed(_zz_1717) + $signed(_zz_1718));
  assign _zz_15227 = _zz_15228[15 : 0];
  assign _zz_15228 = fixTo_1232_dout;
  assign _zz_15229 = _zz_15230[15 : 0];
  assign _zz_15230 = fixTo_1231_dout;
  assign _zz_15231 = _zz_15232;
  assign _zz_15232 = ($signed(_zz_15233) >>> _zz_3846);
  assign _zz_15233 = _zz_15234;
  assign _zz_15234 = ($signed(_zz_1589) - $signed(_zz_3843));
  assign _zz_15235 = _zz_15236;
  assign _zz_15236 = ($signed(_zz_15237) >>> _zz_3846);
  assign _zz_15237 = _zz_15238;
  assign _zz_15238 = ($signed(_zz_1590) - $signed(_zz_3844));
  assign _zz_15239 = _zz_15240;
  assign _zz_15240 = ($signed(_zz_15241) >>> _zz_3847);
  assign _zz_15241 = _zz_15242;
  assign _zz_15242 = ($signed(_zz_1589) + $signed(_zz_3843));
  assign _zz_15243 = _zz_15244;
  assign _zz_15244 = ($signed(_zz_15245) >>> _zz_3847);
  assign _zz_15245 = _zz_15246;
  assign _zz_15246 = ($signed(_zz_1590) + $signed(_zz_3844));
  assign _zz_15247 = ($signed(twiddle_factor_table_90_real) + $signed(twiddle_factor_table_90_imag));
  assign _zz_15248 = fixTo_1233_dout;
  assign _zz_15249 = ($signed(_zz_1720) - $signed(_zz_1719));
  assign _zz_15250 = ($signed(_zz_1719) + $signed(_zz_1720));
  assign _zz_15251 = _zz_15252[15 : 0];
  assign _zz_15252 = fixTo_1235_dout;
  assign _zz_15253 = _zz_15254[15 : 0];
  assign _zz_15254 = fixTo_1234_dout;
  assign _zz_15255 = _zz_15256;
  assign _zz_15256 = ($signed(_zz_15257) >>> _zz_3851);
  assign _zz_15257 = _zz_15258;
  assign _zz_15258 = ($signed(_zz_1591) - $signed(_zz_3848));
  assign _zz_15259 = _zz_15260;
  assign _zz_15260 = ($signed(_zz_15261) >>> _zz_3851);
  assign _zz_15261 = _zz_15262;
  assign _zz_15262 = ($signed(_zz_1592) - $signed(_zz_3849));
  assign _zz_15263 = _zz_15264;
  assign _zz_15264 = ($signed(_zz_15265) >>> _zz_3852);
  assign _zz_15265 = _zz_15266;
  assign _zz_15266 = ($signed(_zz_1591) + $signed(_zz_3848));
  assign _zz_15267 = _zz_15268;
  assign _zz_15268 = ($signed(_zz_15269) >>> _zz_3852);
  assign _zz_15269 = _zz_15270;
  assign _zz_15270 = ($signed(_zz_1592) + $signed(_zz_3849));
  assign _zz_15271 = ($signed(twiddle_factor_table_91_real) + $signed(twiddle_factor_table_91_imag));
  assign _zz_15272 = fixTo_1236_dout;
  assign _zz_15273 = ($signed(_zz_1722) - $signed(_zz_1721));
  assign _zz_15274 = ($signed(_zz_1721) + $signed(_zz_1722));
  assign _zz_15275 = _zz_15276[15 : 0];
  assign _zz_15276 = fixTo_1238_dout;
  assign _zz_15277 = _zz_15278[15 : 0];
  assign _zz_15278 = fixTo_1237_dout;
  assign _zz_15279 = _zz_15280;
  assign _zz_15280 = ($signed(_zz_15281) >>> _zz_3856);
  assign _zz_15281 = _zz_15282;
  assign _zz_15282 = ($signed(_zz_1593) - $signed(_zz_3853));
  assign _zz_15283 = _zz_15284;
  assign _zz_15284 = ($signed(_zz_15285) >>> _zz_3856);
  assign _zz_15285 = _zz_15286;
  assign _zz_15286 = ($signed(_zz_1594) - $signed(_zz_3854));
  assign _zz_15287 = _zz_15288;
  assign _zz_15288 = ($signed(_zz_15289) >>> _zz_3857);
  assign _zz_15289 = _zz_15290;
  assign _zz_15290 = ($signed(_zz_1593) + $signed(_zz_3853));
  assign _zz_15291 = _zz_15292;
  assign _zz_15292 = ($signed(_zz_15293) >>> _zz_3857);
  assign _zz_15293 = _zz_15294;
  assign _zz_15294 = ($signed(_zz_1594) + $signed(_zz_3854));
  assign _zz_15295 = ($signed(twiddle_factor_table_92_real) + $signed(twiddle_factor_table_92_imag));
  assign _zz_15296 = fixTo_1239_dout;
  assign _zz_15297 = ($signed(_zz_1724) - $signed(_zz_1723));
  assign _zz_15298 = ($signed(_zz_1723) + $signed(_zz_1724));
  assign _zz_15299 = _zz_15300[15 : 0];
  assign _zz_15300 = fixTo_1241_dout;
  assign _zz_15301 = _zz_15302[15 : 0];
  assign _zz_15302 = fixTo_1240_dout;
  assign _zz_15303 = _zz_15304;
  assign _zz_15304 = ($signed(_zz_15305) >>> _zz_3861);
  assign _zz_15305 = _zz_15306;
  assign _zz_15306 = ($signed(_zz_1595) - $signed(_zz_3858));
  assign _zz_15307 = _zz_15308;
  assign _zz_15308 = ($signed(_zz_15309) >>> _zz_3861);
  assign _zz_15309 = _zz_15310;
  assign _zz_15310 = ($signed(_zz_1596) - $signed(_zz_3859));
  assign _zz_15311 = _zz_15312;
  assign _zz_15312 = ($signed(_zz_15313) >>> _zz_3862);
  assign _zz_15313 = _zz_15314;
  assign _zz_15314 = ($signed(_zz_1595) + $signed(_zz_3858));
  assign _zz_15315 = _zz_15316;
  assign _zz_15316 = ($signed(_zz_15317) >>> _zz_3862);
  assign _zz_15317 = _zz_15318;
  assign _zz_15318 = ($signed(_zz_1596) + $signed(_zz_3859));
  assign _zz_15319 = ($signed(twiddle_factor_table_93_real) + $signed(twiddle_factor_table_93_imag));
  assign _zz_15320 = fixTo_1242_dout;
  assign _zz_15321 = ($signed(_zz_1726) - $signed(_zz_1725));
  assign _zz_15322 = ($signed(_zz_1725) + $signed(_zz_1726));
  assign _zz_15323 = _zz_15324[15 : 0];
  assign _zz_15324 = fixTo_1244_dout;
  assign _zz_15325 = _zz_15326[15 : 0];
  assign _zz_15326 = fixTo_1243_dout;
  assign _zz_15327 = _zz_15328;
  assign _zz_15328 = ($signed(_zz_15329) >>> _zz_3866);
  assign _zz_15329 = _zz_15330;
  assign _zz_15330 = ($signed(_zz_1597) - $signed(_zz_3863));
  assign _zz_15331 = _zz_15332;
  assign _zz_15332 = ($signed(_zz_15333) >>> _zz_3866);
  assign _zz_15333 = _zz_15334;
  assign _zz_15334 = ($signed(_zz_1598) - $signed(_zz_3864));
  assign _zz_15335 = _zz_15336;
  assign _zz_15336 = ($signed(_zz_15337) >>> _zz_3867);
  assign _zz_15337 = _zz_15338;
  assign _zz_15338 = ($signed(_zz_1597) + $signed(_zz_3863));
  assign _zz_15339 = _zz_15340;
  assign _zz_15340 = ($signed(_zz_15341) >>> _zz_3867);
  assign _zz_15341 = _zz_15342;
  assign _zz_15342 = ($signed(_zz_1598) + $signed(_zz_3864));
  assign _zz_15343 = ($signed(twiddle_factor_table_94_real) + $signed(twiddle_factor_table_94_imag));
  assign _zz_15344 = fixTo_1245_dout;
  assign _zz_15345 = ($signed(_zz_1728) - $signed(_zz_1727));
  assign _zz_15346 = ($signed(_zz_1727) + $signed(_zz_1728));
  assign _zz_15347 = _zz_15348[15 : 0];
  assign _zz_15348 = fixTo_1247_dout;
  assign _zz_15349 = _zz_15350[15 : 0];
  assign _zz_15350 = fixTo_1246_dout;
  assign _zz_15351 = _zz_15352;
  assign _zz_15352 = ($signed(_zz_15353) >>> _zz_3871);
  assign _zz_15353 = _zz_15354;
  assign _zz_15354 = ($signed(_zz_1599) - $signed(_zz_3868));
  assign _zz_15355 = _zz_15356;
  assign _zz_15356 = ($signed(_zz_15357) >>> _zz_3871);
  assign _zz_15357 = _zz_15358;
  assign _zz_15358 = ($signed(_zz_1600) - $signed(_zz_3869));
  assign _zz_15359 = _zz_15360;
  assign _zz_15360 = ($signed(_zz_15361) >>> _zz_3872);
  assign _zz_15361 = _zz_15362;
  assign _zz_15362 = ($signed(_zz_1599) + $signed(_zz_3868));
  assign _zz_15363 = _zz_15364;
  assign _zz_15364 = ($signed(_zz_15365) >>> _zz_3872);
  assign _zz_15365 = _zz_15366;
  assign _zz_15366 = ($signed(_zz_1600) + $signed(_zz_3869));
  assign _zz_15367 = ($signed(twiddle_factor_table_95_real) + $signed(twiddle_factor_table_95_imag));
  assign _zz_15368 = fixTo_1248_dout;
  assign _zz_15369 = ($signed(_zz_1730) - $signed(_zz_1729));
  assign _zz_15370 = ($signed(_zz_1729) + $signed(_zz_1730));
  assign _zz_15371 = _zz_15372[15 : 0];
  assign _zz_15372 = fixTo_1250_dout;
  assign _zz_15373 = _zz_15374[15 : 0];
  assign _zz_15374 = fixTo_1249_dout;
  assign _zz_15375 = _zz_15376;
  assign _zz_15376 = ($signed(_zz_15377) >>> _zz_3876);
  assign _zz_15377 = _zz_15378;
  assign _zz_15378 = ($signed(_zz_1601) - $signed(_zz_3873));
  assign _zz_15379 = _zz_15380;
  assign _zz_15380 = ($signed(_zz_15381) >>> _zz_3876);
  assign _zz_15381 = _zz_15382;
  assign _zz_15382 = ($signed(_zz_1602) - $signed(_zz_3874));
  assign _zz_15383 = _zz_15384;
  assign _zz_15384 = ($signed(_zz_15385) >>> _zz_3877);
  assign _zz_15385 = _zz_15386;
  assign _zz_15386 = ($signed(_zz_1601) + $signed(_zz_3873));
  assign _zz_15387 = _zz_15388;
  assign _zz_15388 = ($signed(_zz_15389) >>> _zz_3877);
  assign _zz_15389 = _zz_15390;
  assign _zz_15390 = ($signed(_zz_1602) + $signed(_zz_3874));
  assign _zz_15391 = ($signed(twiddle_factor_table_96_real) + $signed(twiddle_factor_table_96_imag));
  assign _zz_15392 = fixTo_1251_dout;
  assign _zz_15393 = ($signed(_zz_1732) - $signed(_zz_1731));
  assign _zz_15394 = ($signed(_zz_1731) + $signed(_zz_1732));
  assign _zz_15395 = _zz_15396[15 : 0];
  assign _zz_15396 = fixTo_1253_dout;
  assign _zz_15397 = _zz_15398[15 : 0];
  assign _zz_15398 = fixTo_1252_dout;
  assign _zz_15399 = _zz_15400;
  assign _zz_15400 = ($signed(_zz_15401) >>> _zz_3881);
  assign _zz_15401 = _zz_15402;
  assign _zz_15402 = ($signed(_zz_1603) - $signed(_zz_3878));
  assign _zz_15403 = _zz_15404;
  assign _zz_15404 = ($signed(_zz_15405) >>> _zz_3881);
  assign _zz_15405 = _zz_15406;
  assign _zz_15406 = ($signed(_zz_1604) - $signed(_zz_3879));
  assign _zz_15407 = _zz_15408;
  assign _zz_15408 = ($signed(_zz_15409) >>> _zz_3882);
  assign _zz_15409 = _zz_15410;
  assign _zz_15410 = ($signed(_zz_1603) + $signed(_zz_3878));
  assign _zz_15411 = _zz_15412;
  assign _zz_15412 = ($signed(_zz_15413) >>> _zz_3882);
  assign _zz_15413 = _zz_15414;
  assign _zz_15414 = ($signed(_zz_1604) + $signed(_zz_3879));
  assign _zz_15415 = ($signed(twiddle_factor_table_97_real) + $signed(twiddle_factor_table_97_imag));
  assign _zz_15416 = fixTo_1254_dout;
  assign _zz_15417 = ($signed(_zz_1734) - $signed(_zz_1733));
  assign _zz_15418 = ($signed(_zz_1733) + $signed(_zz_1734));
  assign _zz_15419 = _zz_15420[15 : 0];
  assign _zz_15420 = fixTo_1256_dout;
  assign _zz_15421 = _zz_15422[15 : 0];
  assign _zz_15422 = fixTo_1255_dout;
  assign _zz_15423 = _zz_15424;
  assign _zz_15424 = ($signed(_zz_15425) >>> _zz_3886);
  assign _zz_15425 = _zz_15426;
  assign _zz_15426 = ($signed(_zz_1605) - $signed(_zz_3883));
  assign _zz_15427 = _zz_15428;
  assign _zz_15428 = ($signed(_zz_15429) >>> _zz_3886);
  assign _zz_15429 = _zz_15430;
  assign _zz_15430 = ($signed(_zz_1606) - $signed(_zz_3884));
  assign _zz_15431 = _zz_15432;
  assign _zz_15432 = ($signed(_zz_15433) >>> _zz_3887);
  assign _zz_15433 = _zz_15434;
  assign _zz_15434 = ($signed(_zz_1605) + $signed(_zz_3883));
  assign _zz_15435 = _zz_15436;
  assign _zz_15436 = ($signed(_zz_15437) >>> _zz_3887);
  assign _zz_15437 = _zz_15438;
  assign _zz_15438 = ($signed(_zz_1606) + $signed(_zz_3884));
  assign _zz_15439 = ($signed(twiddle_factor_table_98_real) + $signed(twiddle_factor_table_98_imag));
  assign _zz_15440 = fixTo_1257_dout;
  assign _zz_15441 = ($signed(_zz_1736) - $signed(_zz_1735));
  assign _zz_15442 = ($signed(_zz_1735) + $signed(_zz_1736));
  assign _zz_15443 = _zz_15444[15 : 0];
  assign _zz_15444 = fixTo_1259_dout;
  assign _zz_15445 = _zz_15446[15 : 0];
  assign _zz_15446 = fixTo_1258_dout;
  assign _zz_15447 = _zz_15448;
  assign _zz_15448 = ($signed(_zz_15449) >>> _zz_3891);
  assign _zz_15449 = _zz_15450;
  assign _zz_15450 = ($signed(_zz_1607) - $signed(_zz_3888));
  assign _zz_15451 = _zz_15452;
  assign _zz_15452 = ($signed(_zz_15453) >>> _zz_3891);
  assign _zz_15453 = _zz_15454;
  assign _zz_15454 = ($signed(_zz_1608) - $signed(_zz_3889));
  assign _zz_15455 = _zz_15456;
  assign _zz_15456 = ($signed(_zz_15457) >>> _zz_3892);
  assign _zz_15457 = _zz_15458;
  assign _zz_15458 = ($signed(_zz_1607) + $signed(_zz_3888));
  assign _zz_15459 = _zz_15460;
  assign _zz_15460 = ($signed(_zz_15461) >>> _zz_3892);
  assign _zz_15461 = _zz_15462;
  assign _zz_15462 = ($signed(_zz_1608) + $signed(_zz_3889));
  assign _zz_15463 = ($signed(twiddle_factor_table_99_real) + $signed(twiddle_factor_table_99_imag));
  assign _zz_15464 = fixTo_1260_dout;
  assign _zz_15465 = ($signed(_zz_1738) - $signed(_zz_1737));
  assign _zz_15466 = ($signed(_zz_1737) + $signed(_zz_1738));
  assign _zz_15467 = _zz_15468[15 : 0];
  assign _zz_15468 = fixTo_1262_dout;
  assign _zz_15469 = _zz_15470[15 : 0];
  assign _zz_15470 = fixTo_1261_dout;
  assign _zz_15471 = _zz_15472;
  assign _zz_15472 = ($signed(_zz_15473) >>> _zz_3896);
  assign _zz_15473 = _zz_15474;
  assign _zz_15474 = ($signed(_zz_1609) - $signed(_zz_3893));
  assign _zz_15475 = _zz_15476;
  assign _zz_15476 = ($signed(_zz_15477) >>> _zz_3896);
  assign _zz_15477 = _zz_15478;
  assign _zz_15478 = ($signed(_zz_1610) - $signed(_zz_3894));
  assign _zz_15479 = _zz_15480;
  assign _zz_15480 = ($signed(_zz_15481) >>> _zz_3897);
  assign _zz_15481 = _zz_15482;
  assign _zz_15482 = ($signed(_zz_1609) + $signed(_zz_3893));
  assign _zz_15483 = _zz_15484;
  assign _zz_15484 = ($signed(_zz_15485) >>> _zz_3897);
  assign _zz_15485 = _zz_15486;
  assign _zz_15486 = ($signed(_zz_1610) + $signed(_zz_3894));
  assign _zz_15487 = ($signed(twiddle_factor_table_100_real) + $signed(twiddle_factor_table_100_imag));
  assign _zz_15488 = fixTo_1263_dout;
  assign _zz_15489 = ($signed(_zz_1740) - $signed(_zz_1739));
  assign _zz_15490 = ($signed(_zz_1739) + $signed(_zz_1740));
  assign _zz_15491 = _zz_15492[15 : 0];
  assign _zz_15492 = fixTo_1265_dout;
  assign _zz_15493 = _zz_15494[15 : 0];
  assign _zz_15494 = fixTo_1264_dout;
  assign _zz_15495 = _zz_15496;
  assign _zz_15496 = ($signed(_zz_15497) >>> _zz_3901);
  assign _zz_15497 = _zz_15498;
  assign _zz_15498 = ($signed(_zz_1611) - $signed(_zz_3898));
  assign _zz_15499 = _zz_15500;
  assign _zz_15500 = ($signed(_zz_15501) >>> _zz_3901);
  assign _zz_15501 = _zz_15502;
  assign _zz_15502 = ($signed(_zz_1612) - $signed(_zz_3899));
  assign _zz_15503 = _zz_15504;
  assign _zz_15504 = ($signed(_zz_15505) >>> _zz_3902);
  assign _zz_15505 = _zz_15506;
  assign _zz_15506 = ($signed(_zz_1611) + $signed(_zz_3898));
  assign _zz_15507 = _zz_15508;
  assign _zz_15508 = ($signed(_zz_15509) >>> _zz_3902);
  assign _zz_15509 = _zz_15510;
  assign _zz_15510 = ($signed(_zz_1612) + $signed(_zz_3899));
  assign _zz_15511 = ($signed(twiddle_factor_table_101_real) + $signed(twiddle_factor_table_101_imag));
  assign _zz_15512 = fixTo_1266_dout;
  assign _zz_15513 = ($signed(_zz_1742) - $signed(_zz_1741));
  assign _zz_15514 = ($signed(_zz_1741) + $signed(_zz_1742));
  assign _zz_15515 = _zz_15516[15 : 0];
  assign _zz_15516 = fixTo_1268_dout;
  assign _zz_15517 = _zz_15518[15 : 0];
  assign _zz_15518 = fixTo_1267_dout;
  assign _zz_15519 = _zz_15520;
  assign _zz_15520 = ($signed(_zz_15521) >>> _zz_3906);
  assign _zz_15521 = _zz_15522;
  assign _zz_15522 = ($signed(_zz_1613) - $signed(_zz_3903));
  assign _zz_15523 = _zz_15524;
  assign _zz_15524 = ($signed(_zz_15525) >>> _zz_3906);
  assign _zz_15525 = _zz_15526;
  assign _zz_15526 = ($signed(_zz_1614) - $signed(_zz_3904));
  assign _zz_15527 = _zz_15528;
  assign _zz_15528 = ($signed(_zz_15529) >>> _zz_3907);
  assign _zz_15529 = _zz_15530;
  assign _zz_15530 = ($signed(_zz_1613) + $signed(_zz_3903));
  assign _zz_15531 = _zz_15532;
  assign _zz_15532 = ($signed(_zz_15533) >>> _zz_3907);
  assign _zz_15533 = _zz_15534;
  assign _zz_15534 = ($signed(_zz_1614) + $signed(_zz_3904));
  assign _zz_15535 = ($signed(twiddle_factor_table_102_real) + $signed(twiddle_factor_table_102_imag));
  assign _zz_15536 = fixTo_1269_dout;
  assign _zz_15537 = ($signed(_zz_1744) - $signed(_zz_1743));
  assign _zz_15538 = ($signed(_zz_1743) + $signed(_zz_1744));
  assign _zz_15539 = _zz_15540[15 : 0];
  assign _zz_15540 = fixTo_1271_dout;
  assign _zz_15541 = _zz_15542[15 : 0];
  assign _zz_15542 = fixTo_1270_dout;
  assign _zz_15543 = _zz_15544;
  assign _zz_15544 = ($signed(_zz_15545) >>> _zz_3911);
  assign _zz_15545 = _zz_15546;
  assign _zz_15546 = ($signed(_zz_1615) - $signed(_zz_3908));
  assign _zz_15547 = _zz_15548;
  assign _zz_15548 = ($signed(_zz_15549) >>> _zz_3911);
  assign _zz_15549 = _zz_15550;
  assign _zz_15550 = ($signed(_zz_1616) - $signed(_zz_3909));
  assign _zz_15551 = _zz_15552;
  assign _zz_15552 = ($signed(_zz_15553) >>> _zz_3912);
  assign _zz_15553 = _zz_15554;
  assign _zz_15554 = ($signed(_zz_1615) + $signed(_zz_3908));
  assign _zz_15555 = _zz_15556;
  assign _zz_15556 = ($signed(_zz_15557) >>> _zz_3912);
  assign _zz_15557 = _zz_15558;
  assign _zz_15558 = ($signed(_zz_1616) + $signed(_zz_3909));
  assign _zz_15559 = ($signed(twiddle_factor_table_103_real) + $signed(twiddle_factor_table_103_imag));
  assign _zz_15560 = fixTo_1272_dout;
  assign _zz_15561 = ($signed(_zz_1746) - $signed(_zz_1745));
  assign _zz_15562 = ($signed(_zz_1745) + $signed(_zz_1746));
  assign _zz_15563 = _zz_15564[15 : 0];
  assign _zz_15564 = fixTo_1274_dout;
  assign _zz_15565 = _zz_15566[15 : 0];
  assign _zz_15566 = fixTo_1273_dout;
  assign _zz_15567 = _zz_15568;
  assign _zz_15568 = ($signed(_zz_15569) >>> _zz_3916);
  assign _zz_15569 = _zz_15570;
  assign _zz_15570 = ($signed(_zz_1617) - $signed(_zz_3913));
  assign _zz_15571 = _zz_15572;
  assign _zz_15572 = ($signed(_zz_15573) >>> _zz_3916);
  assign _zz_15573 = _zz_15574;
  assign _zz_15574 = ($signed(_zz_1618) - $signed(_zz_3914));
  assign _zz_15575 = _zz_15576;
  assign _zz_15576 = ($signed(_zz_15577) >>> _zz_3917);
  assign _zz_15577 = _zz_15578;
  assign _zz_15578 = ($signed(_zz_1617) + $signed(_zz_3913));
  assign _zz_15579 = _zz_15580;
  assign _zz_15580 = ($signed(_zz_15581) >>> _zz_3917);
  assign _zz_15581 = _zz_15582;
  assign _zz_15582 = ($signed(_zz_1618) + $signed(_zz_3914));
  assign _zz_15583 = ($signed(twiddle_factor_table_104_real) + $signed(twiddle_factor_table_104_imag));
  assign _zz_15584 = fixTo_1275_dout;
  assign _zz_15585 = ($signed(_zz_1748) - $signed(_zz_1747));
  assign _zz_15586 = ($signed(_zz_1747) + $signed(_zz_1748));
  assign _zz_15587 = _zz_15588[15 : 0];
  assign _zz_15588 = fixTo_1277_dout;
  assign _zz_15589 = _zz_15590[15 : 0];
  assign _zz_15590 = fixTo_1276_dout;
  assign _zz_15591 = _zz_15592;
  assign _zz_15592 = ($signed(_zz_15593) >>> _zz_3921);
  assign _zz_15593 = _zz_15594;
  assign _zz_15594 = ($signed(_zz_1619) - $signed(_zz_3918));
  assign _zz_15595 = _zz_15596;
  assign _zz_15596 = ($signed(_zz_15597) >>> _zz_3921);
  assign _zz_15597 = _zz_15598;
  assign _zz_15598 = ($signed(_zz_1620) - $signed(_zz_3919));
  assign _zz_15599 = _zz_15600;
  assign _zz_15600 = ($signed(_zz_15601) >>> _zz_3922);
  assign _zz_15601 = _zz_15602;
  assign _zz_15602 = ($signed(_zz_1619) + $signed(_zz_3918));
  assign _zz_15603 = _zz_15604;
  assign _zz_15604 = ($signed(_zz_15605) >>> _zz_3922);
  assign _zz_15605 = _zz_15606;
  assign _zz_15606 = ($signed(_zz_1620) + $signed(_zz_3919));
  assign _zz_15607 = ($signed(twiddle_factor_table_105_real) + $signed(twiddle_factor_table_105_imag));
  assign _zz_15608 = fixTo_1278_dout;
  assign _zz_15609 = ($signed(_zz_1750) - $signed(_zz_1749));
  assign _zz_15610 = ($signed(_zz_1749) + $signed(_zz_1750));
  assign _zz_15611 = _zz_15612[15 : 0];
  assign _zz_15612 = fixTo_1280_dout;
  assign _zz_15613 = _zz_15614[15 : 0];
  assign _zz_15614 = fixTo_1279_dout;
  assign _zz_15615 = _zz_15616;
  assign _zz_15616 = ($signed(_zz_15617) >>> _zz_3926);
  assign _zz_15617 = _zz_15618;
  assign _zz_15618 = ($signed(_zz_1621) - $signed(_zz_3923));
  assign _zz_15619 = _zz_15620;
  assign _zz_15620 = ($signed(_zz_15621) >>> _zz_3926);
  assign _zz_15621 = _zz_15622;
  assign _zz_15622 = ($signed(_zz_1622) - $signed(_zz_3924));
  assign _zz_15623 = _zz_15624;
  assign _zz_15624 = ($signed(_zz_15625) >>> _zz_3927);
  assign _zz_15625 = _zz_15626;
  assign _zz_15626 = ($signed(_zz_1621) + $signed(_zz_3923));
  assign _zz_15627 = _zz_15628;
  assign _zz_15628 = ($signed(_zz_15629) >>> _zz_3927);
  assign _zz_15629 = _zz_15630;
  assign _zz_15630 = ($signed(_zz_1622) + $signed(_zz_3924));
  assign _zz_15631 = ($signed(twiddle_factor_table_106_real) + $signed(twiddle_factor_table_106_imag));
  assign _zz_15632 = fixTo_1281_dout;
  assign _zz_15633 = ($signed(_zz_1752) - $signed(_zz_1751));
  assign _zz_15634 = ($signed(_zz_1751) + $signed(_zz_1752));
  assign _zz_15635 = _zz_15636[15 : 0];
  assign _zz_15636 = fixTo_1283_dout;
  assign _zz_15637 = _zz_15638[15 : 0];
  assign _zz_15638 = fixTo_1282_dout;
  assign _zz_15639 = _zz_15640;
  assign _zz_15640 = ($signed(_zz_15641) >>> _zz_3931);
  assign _zz_15641 = _zz_15642;
  assign _zz_15642 = ($signed(_zz_1623) - $signed(_zz_3928));
  assign _zz_15643 = _zz_15644;
  assign _zz_15644 = ($signed(_zz_15645) >>> _zz_3931);
  assign _zz_15645 = _zz_15646;
  assign _zz_15646 = ($signed(_zz_1624) - $signed(_zz_3929));
  assign _zz_15647 = _zz_15648;
  assign _zz_15648 = ($signed(_zz_15649) >>> _zz_3932);
  assign _zz_15649 = _zz_15650;
  assign _zz_15650 = ($signed(_zz_1623) + $signed(_zz_3928));
  assign _zz_15651 = _zz_15652;
  assign _zz_15652 = ($signed(_zz_15653) >>> _zz_3932);
  assign _zz_15653 = _zz_15654;
  assign _zz_15654 = ($signed(_zz_1624) + $signed(_zz_3929));
  assign _zz_15655 = ($signed(twiddle_factor_table_107_real) + $signed(twiddle_factor_table_107_imag));
  assign _zz_15656 = fixTo_1284_dout;
  assign _zz_15657 = ($signed(_zz_1754) - $signed(_zz_1753));
  assign _zz_15658 = ($signed(_zz_1753) + $signed(_zz_1754));
  assign _zz_15659 = _zz_15660[15 : 0];
  assign _zz_15660 = fixTo_1286_dout;
  assign _zz_15661 = _zz_15662[15 : 0];
  assign _zz_15662 = fixTo_1285_dout;
  assign _zz_15663 = _zz_15664;
  assign _zz_15664 = ($signed(_zz_15665) >>> _zz_3936);
  assign _zz_15665 = _zz_15666;
  assign _zz_15666 = ($signed(_zz_1625) - $signed(_zz_3933));
  assign _zz_15667 = _zz_15668;
  assign _zz_15668 = ($signed(_zz_15669) >>> _zz_3936);
  assign _zz_15669 = _zz_15670;
  assign _zz_15670 = ($signed(_zz_1626) - $signed(_zz_3934));
  assign _zz_15671 = _zz_15672;
  assign _zz_15672 = ($signed(_zz_15673) >>> _zz_3937);
  assign _zz_15673 = _zz_15674;
  assign _zz_15674 = ($signed(_zz_1625) + $signed(_zz_3933));
  assign _zz_15675 = _zz_15676;
  assign _zz_15676 = ($signed(_zz_15677) >>> _zz_3937);
  assign _zz_15677 = _zz_15678;
  assign _zz_15678 = ($signed(_zz_1626) + $signed(_zz_3934));
  assign _zz_15679 = ($signed(twiddle_factor_table_108_real) + $signed(twiddle_factor_table_108_imag));
  assign _zz_15680 = fixTo_1287_dout;
  assign _zz_15681 = ($signed(_zz_1756) - $signed(_zz_1755));
  assign _zz_15682 = ($signed(_zz_1755) + $signed(_zz_1756));
  assign _zz_15683 = _zz_15684[15 : 0];
  assign _zz_15684 = fixTo_1289_dout;
  assign _zz_15685 = _zz_15686[15 : 0];
  assign _zz_15686 = fixTo_1288_dout;
  assign _zz_15687 = _zz_15688;
  assign _zz_15688 = ($signed(_zz_15689) >>> _zz_3941);
  assign _zz_15689 = _zz_15690;
  assign _zz_15690 = ($signed(_zz_1627) - $signed(_zz_3938));
  assign _zz_15691 = _zz_15692;
  assign _zz_15692 = ($signed(_zz_15693) >>> _zz_3941);
  assign _zz_15693 = _zz_15694;
  assign _zz_15694 = ($signed(_zz_1628) - $signed(_zz_3939));
  assign _zz_15695 = _zz_15696;
  assign _zz_15696 = ($signed(_zz_15697) >>> _zz_3942);
  assign _zz_15697 = _zz_15698;
  assign _zz_15698 = ($signed(_zz_1627) + $signed(_zz_3938));
  assign _zz_15699 = _zz_15700;
  assign _zz_15700 = ($signed(_zz_15701) >>> _zz_3942);
  assign _zz_15701 = _zz_15702;
  assign _zz_15702 = ($signed(_zz_1628) + $signed(_zz_3939));
  assign _zz_15703 = ($signed(twiddle_factor_table_109_real) + $signed(twiddle_factor_table_109_imag));
  assign _zz_15704 = fixTo_1290_dout;
  assign _zz_15705 = ($signed(_zz_1758) - $signed(_zz_1757));
  assign _zz_15706 = ($signed(_zz_1757) + $signed(_zz_1758));
  assign _zz_15707 = _zz_15708[15 : 0];
  assign _zz_15708 = fixTo_1292_dout;
  assign _zz_15709 = _zz_15710[15 : 0];
  assign _zz_15710 = fixTo_1291_dout;
  assign _zz_15711 = _zz_15712;
  assign _zz_15712 = ($signed(_zz_15713) >>> _zz_3946);
  assign _zz_15713 = _zz_15714;
  assign _zz_15714 = ($signed(_zz_1629) - $signed(_zz_3943));
  assign _zz_15715 = _zz_15716;
  assign _zz_15716 = ($signed(_zz_15717) >>> _zz_3946);
  assign _zz_15717 = _zz_15718;
  assign _zz_15718 = ($signed(_zz_1630) - $signed(_zz_3944));
  assign _zz_15719 = _zz_15720;
  assign _zz_15720 = ($signed(_zz_15721) >>> _zz_3947);
  assign _zz_15721 = _zz_15722;
  assign _zz_15722 = ($signed(_zz_1629) + $signed(_zz_3943));
  assign _zz_15723 = _zz_15724;
  assign _zz_15724 = ($signed(_zz_15725) >>> _zz_3947);
  assign _zz_15725 = _zz_15726;
  assign _zz_15726 = ($signed(_zz_1630) + $signed(_zz_3944));
  assign _zz_15727 = ($signed(twiddle_factor_table_110_real) + $signed(twiddle_factor_table_110_imag));
  assign _zz_15728 = fixTo_1293_dout;
  assign _zz_15729 = ($signed(_zz_1760) - $signed(_zz_1759));
  assign _zz_15730 = ($signed(_zz_1759) + $signed(_zz_1760));
  assign _zz_15731 = _zz_15732[15 : 0];
  assign _zz_15732 = fixTo_1295_dout;
  assign _zz_15733 = _zz_15734[15 : 0];
  assign _zz_15734 = fixTo_1294_dout;
  assign _zz_15735 = _zz_15736;
  assign _zz_15736 = ($signed(_zz_15737) >>> _zz_3951);
  assign _zz_15737 = _zz_15738;
  assign _zz_15738 = ($signed(_zz_1631) - $signed(_zz_3948));
  assign _zz_15739 = _zz_15740;
  assign _zz_15740 = ($signed(_zz_15741) >>> _zz_3951);
  assign _zz_15741 = _zz_15742;
  assign _zz_15742 = ($signed(_zz_1632) - $signed(_zz_3949));
  assign _zz_15743 = _zz_15744;
  assign _zz_15744 = ($signed(_zz_15745) >>> _zz_3952);
  assign _zz_15745 = _zz_15746;
  assign _zz_15746 = ($signed(_zz_1631) + $signed(_zz_3948));
  assign _zz_15747 = _zz_15748;
  assign _zz_15748 = ($signed(_zz_15749) >>> _zz_3952);
  assign _zz_15749 = _zz_15750;
  assign _zz_15750 = ($signed(_zz_1632) + $signed(_zz_3949));
  assign _zz_15751 = ($signed(twiddle_factor_table_111_real) + $signed(twiddle_factor_table_111_imag));
  assign _zz_15752 = fixTo_1296_dout;
  assign _zz_15753 = ($signed(_zz_1762) - $signed(_zz_1761));
  assign _zz_15754 = ($signed(_zz_1761) + $signed(_zz_1762));
  assign _zz_15755 = _zz_15756[15 : 0];
  assign _zz_15756 = fixTo_1298_dout;
  assign _zz_15757 = _zz_15758[15 : 0];
  assign _zz_15758 = fixTo_1297_dout;
  assign _zz_15759 = _zz_15760;
  assign _zz_15760 = ($signed(_zz_15761) >>> _zz_3956);
  assign _zz_15761 = _zz_15762;
  assign _zz_15762 = ($signed(_zz_1633) - $signed(_zz_3953));
  assign _zz_15763 = _zz_15764;
  assign _zz_15764 = ($signed(_zz_15765) >>> _zz_3956);
  assign _zz_15765 = _zz_15766;
  assign _zz_15766 = ($signed(_zz_1634) - $signed(_zz_3954));
  assign _zz_15767 = _zz_15768;
  assign _zz_15768 = ($signed(_zz_15769) >>> _zz_3957);
  assign _zz_15769 = _zz_15770;
  assign _zz_15770 = ($signed(_zz_1633) + $signed(_zz_3953));
  assign _zz_15771 = _zz_15772;
  assign _zz_15772 = ($signed(_zz_15773) >>> _zz_3957);
  assign _zz_15773 = _zz_15774;
  assign _zz_15774 = ($signed(_zz_1634) + $signed(_zz_3954));
  assign _zz_15775 = ($signed(twiddle_factor_table_112_real) + $signed(twiddle_factor_table_112_imag));
  assign _zz_15776 = fixTo_1299_dout;
  assign _zz_15777 = ($signed(_zz_1764) - $signed(_zz_1763));
  assign _zz_15778 = ($signed(_zz_1763) + $signed(_zz_1764));
  assign _zz_15779 = _zz_15780[15 : 0];
  assign _zz_15780 = fixTo_1301_dout;
  assign _zz_15781 = _zz_15782[15 : 0];
  assign _zz_15782 = fixTo_1300_dout;
  assign _zz_15783 = _zz_15784;
  assign _zz_15784 = ($signed(_zz_15785) >>> _zz_3961);
  assign _zz_15785 = _zz_15786;
  assign _zz_15786 = ($signed(_zz_1635) - $signed(_zz_3958));
  assign _zz_15787 = _zz_15788;
  assign _zz_15788 = ($signed(_zz_15789) >>> _zz_3961);
  assign _zz_15789 = _zz_15790;
  assign _zz_15790 = ($signed(_zz_1636) - $signed(_zz_3959));
  assign _zz_15791 = _zz_15792;
  assign _zz_15792 = ($signed(_zz_15793) >>> _zz_3962);
  assign _zz_15793 = _zz_15794;
  assign _zz_15794 = ($signed(_zz_1635) + $signed(_zz_3958));
  assign _zz_15795 = _zz_15796;
  assign _zz_15796 = ($signed(_zz_15797) >>> _zz_3962);
  assign _zz_15797 = _zz_15798;
  assign _zz_15798 = ($signed(_zz_1636) + $signed(_zz_3959));
  assign _zz_15799 = ($signed(twiddle_factor_table_113_real) + $signed(twiddle_factor_table_113_imag));
  assign _zz_15800 = fixTo_1302_dout;
  assign _zz_15801 = ($signed(_zz_1766) - $signed(_zz_1765));
  assign _zz_15802 = ($signed(_zz_1765) + $signed(_zz_1766));
  assign _zz_15803 = _zz_15804[15 : 0];
  assign _zz_15804 = fixTo_1304_dout;
  assign _zz_15805 = _zz_15806[15 : 0];
  assign _zz_15806 = fixTo_1303_dout;
  assign _zz_15807 = _zz_15808;
  assign _zz_15808 = ($signed(_zz_15809) >>> _zz_3966);
  assign _zz_15809 = _zz_15810;
  assign _zz_15810 = ($signed(_zz_1637) - $signed(_zz_3963));
  assign _zz_15811 = _zz_15812;
  assign _zz_15812 = ($signed(_zz_15813) >>> _zz_3966);
  assign _zz_15813 = _zz_15814;
  assign _zz_15814 = ($signed(_zz_1638) - $signed(_zz_3964));
  assign _zz_15815 = _zz_15816;
  assign _zz_15816 = ($signed(_zz_15817) >>> _zz_3967);
  assign _zz_15817 = _zz_15818;
  assign _zz_15818 = ($signed(_zz_1637) + $signed(_zz_3963));
  assign _zz_15819 = _zz_15820;
  assign _zz_15820 = ($signed(_zz_15821) >>> _zz_3967);
  assign _zz_15821 = _zz_15822;
  assign _zz_15822 = ($signed(_zz_1638) + $signed(_zz_3964));
  assign _zz_15823 = ($signed(twiddle_factor_table_114_real) + $signed(twiddle_factor_table_114_imag));
  assign _zz_15824 = fixTo_1305_dout;
  assign _zz_15825 = ($signed(_zz_1768) - $signed(_zz_1767));
  assign _zz_15826 = ($signed(_zz_1767) + $signed(_zz_1768));
  assign _zz_15827 = _zz_15828[15 : 0];
  assign _zz_15828 = fixTo_1307_dout;
  assign _zz_15829 = _zz_15830[15 : 0];
  assign _zz_15830 = fixTo_1306_dout;
  assign _zz_15831 = _zz_15832;
  assign _zz_15832 = ($signed(_zz_15833) >>> _zz_3971);
  assign _zz_15833 = _zz_15834;
  assign _zz_15834 = ($signed(_zz_1639) - $signed(_zz_3968));
  assign _zz_15835 = _zz_15836;
  assign _zz_15836 = ($signed(_zz_15837) >>> _zz_3971);
  assign _zz_15837 = _zz_15838;
  assign _zz_15838 = ($signed(_zz_1640) - $signed(_zz_3969));
  assign _zz_15839 = _zz_15840;
  assign _zz_15840 = ($signed(_zz_15841) >>> _zz_3972);
  assign _zz_15841 = _zz_15842;
  assign _zz_15842 = ($signed(_zz_1639) + $signed(_zz_3968));
  assign _zz_15843 = _zz_15844;
  assign _zz_15844 = ($signed(_zz_15845) >>> _zz_3972);
  assign _zz_15845 = _zz_15846;
  assign _zz_15846 = ($signed(_zz_1640) + $signed(_zz_3969));
  assign _zz_15847 = ($signed(twiddle_factor_table_115_real) + $signed(twiddle_factor_table_115_imag));
  assign _zz_15848 = fixTo_1308_dout;
  assign _zz_15849 = ($signed(_zz_1770) - $signed(_zz_1769));
  assign _zz_15850 = ($signed(_zz_1769) + $signed(_zz_1770));
  assign _zz_15851 = _zz_15852[15 : 0];
  assign _zz_15852 = fixTo_1310_dout;
  assign _zz_15853 = _zz_15854[15 : 0];
  assign _zz_15854 = fixTo_1309_dout;
  assign _zz_15855 = _zz_15856;
  assign _zz_15856 = ($signed(_zz_15857) >>> _zz_3976);
  assign _zz_15857 = _zz_15858;
  assign _zz_15858 = ($signed(_zz_1641) - $signed(_zz_3973));
  assign _zz_15859 = _zz_15860;
  assign _zz_15860 = ($signed(_zz_15861) >>> _zz_3976);
  assign _zz_15861 = _zz_15862;
  assign _zz_15862 = ($signed(_zz_1642) - $signed(_zz_3974));
  assign _zz_15863 = _zz_15864;
  assign _zz_15864 = ($signed(_zz_15865) >>> _zz_3977);
  assign _zz_15865 = _zz_15866;
  assign _zz_15866 = ($signed(_zz_1641) + $signed(_zz_3973));
  assign _zz_15867 = _zz_15868;
  assign _zz_15868 = ($signed(_zz_15869) >>> _zz_3977);
  assign _zz_15869 = _zz_15870;
  assign _zz_15870 = ($signed(_zz_1642) + $signed(_zz_3974));
  assign _zz_15871 = ($signed(twiddle_factor_table_116_real) + $signed(twiddle_factor_table_116_imag));
  assign _zz_15872 = fixTo_1311_dout;
  assign _zz_15873 = ($signed(_zz_1772) - $signed(_zz_1771));
  assign _zz_15874 = ($signed(_zz_1771) + $signed(_zz_1772));
  assign _zz_15875 = _zz_15876[15 : 0];
  assign _zz_15876 = fixTo_1313_dout;
  assign _zz_15877 = _zz_15878[15 : 0];
  assign _zz_15878 = fixTo_1312_dout;
  assign _zz_15879 = _zz_15880;
  assign _zz_15880 = ($signed(_zz_15881) >>> _zz_3981);
  assign _zz_15881 = _zz_15882;
  assign _zz_15882 = ($signed(_zz_1643) - $signed(_zz_3978));
  assign _zz_15883 = _zz_15884;
  assign _zz_15884 = ($signed(_zz_15885) >>> _zz_3981);
  assign _zz_15885 = _zz_15886;
  assign _zz_15886 = ($signed(_zz_1644) - $signed(_zz_3979));
  assign _zz_15887 = _zz_15888;
  assign _zz_15888 = ($signed(_zz_15889) >>> _zz_3982);
  assign _zz_15889 = _zz_15890;
  assign _zz_15890 = ($signed(_zz_1643) + $signed(_zz_3978));
  assign _zz_15891 = _zz_15892;
  assign _zz_15892 = ($signed(_zz_15893) >>> _zz_3982);
  assign _zz_15893 = _zz_15894;
  assign _zz_15894 = ($signed(_zz_1644) + $signed(_zz_3979));
  assign _zz_15895 = ($signed(twiddle_factor_table_117_real) + $signed(twiddle_factor_table_117_imag));
  assign _zz_15896 = fixTo_1314_dout;
  assign _zz_15897 = ($signed(_zz_1774) - $signed(_zz_1773));
  assign _zz_15898 = ($signed(_zz_1773) + $signed(_zz_1774));
  assign _zz_15899 = _zz_15900[15 : 0];
  assign _zz_15900 = fixTo_1316_dout;
  assign _zz_15901 = _zz_15902[15 : 0];
  assign _zz_15902 = fixTo_1315_dout;
  assign _zz_15903 = _zz_15904;
  assign _zz_15904 = ($signed(_zz_15905) >>> _zz_3986);
  assign _zz_15905 = _zz_15906;
  assign _zz_15906 = ($signed(_zz_1645) - $signed(_zz_3983));
  assign _zz_15907 = _zz_15908;
  assign _zz_15908 = ($signed(_zz_15909) >>> _zz_3986);
  assign _zz_15909 = _zz_15910;
  assign _zz_15910 = ($signed(_zz_1646) - $signed(_zz_3984));
  assign _zz_15911 = _zz_15912;
  assign _zz_15912 = ($signed(_zz_15913) >>> _zz_3987);
  assign _zz_15913 = _zz_15914;
  assign _zz_15914 = ($signed(_zz_1645) + $signed(_zz_3983));
  assign _zz_15915 = _zz_15916;
  assign _zz_15916 = ($signed(_zz_15917) >>> _zz_3987);
  assign _zz_15917 = _zz_15918;
  assign _zz_15918 = ($signed(_zz_1646) + $signed(_zz_3984));
  assign _zz_15919 = ($signed(twiddle_factor_table_118_real) + $signed(twiddle_factor_table_118_imag));
  assign _zz_15920 = fixTo_1317_dout;
  assign _zz_15921 = ($signed(_zz_1776) - $signed(_zz_1775));
  assign _zz_15922 = ($signed(_zz_1775) + $signed(_zz_1776));
  assign _zz_15923 = _zz_15924[15 : 0];
  assign _zz_15924 = fixTo_1319_dout;
  assign _zz_15925 = _zz_15926[15 : 0];
  assign _zz_15926 = fixTo_1318_dout;
  assign _zz_15927 = _zz_15928;
  assign _zz_15928 = ($signed(_zz_15929) >>> _zz_3991);
  assign _zz_15929 = _zz_15930;
  assign _zz_15930 = ($signed(_zz_1647) - $signed(_zz_3988));
  assign _zz_15931 = _zz_15932;
  assign _zz_15932 = ($signed(_zz_15933) >>> _zz_3991);
  assign _zz_15933 = _zz_15934;
  assign _zz_15934 = ($signed(_zz_1648) - $signed(_zz_3989));
  assign _zz_15935 = _zz_15936;
  assign _zz_15936 = ($signed(_zz_15937) >>> _zz_3992);
  assign _zz_15937 = _zz_15938;
  assign _zz_15938 = ($signed(_zz_1647) + $signed(_zz_3988));
  assign _zz_15939 = _zz_15940;
  assign _zz_15940 = ($signed(_zz_15941) >>> _zz_3992);
  assign _zz_15941 = _zz_15942;
  assign _zz_15942 = ($signed(_zz_1648) + $signed(_zz_3989));
  assign _zz_15943 = ($signed(twiddle_factor_table_119_real) + $signed(twiddle_factor_table_119_imag));
  assign _zz_15944 = fixTo_1320_dout;
  assign _zz_15945 = ($signed(_zz_1778) - $signed(_zz_1777));
  assign _zz_15946 = ($signed(_zz_1777) + $signed(_zz_1778));
  assign _zz_15947 = _zz_15948[15 : 0];
  assign _zz_15948 = fixTo_1322_dout;
  assign _zz_15949 = _zz_15950[15 : 0];
  assign _zz_15950 = fixTo_1321_dout;
  assign _zz_15951 = _zz_15952;
  assign _zz_15952 = ($signed(_zz_15953) >>> _zz_3996);
  assign _zz_15953 = _zz_15954;
  assign _zz_15954 = ($signed(_zz_1649) - $signed(_zz_3993));
  assign _zz_15955 = _zz_15956;
  assign _zz_15956 = ($signed(_zz_15957) >>> _zz_3996);
  assign _zz_15957 = _zz_15958;
  assign _zz_15958 = ($signed(_zz_1650) - $signed(_zz_3994));
  assign _zz_15959 = _zz_15960;
  assign _zz_15960 = ($signed(_zz_15961) >>> _zz_3997);
  assign _zz_15961 = _zz_15962;
  assign _zz_15962 = ($signed(_zz_1649) + $signed(_zz_3993));
  assign _zz_15963 = _zz_15964;
  assign _zz_15964 = ($signed(_zz_15965) >>> _zz_3997);
  assign _zz_15965 = _zz_15966;
  assign _zz_15966 = ($signed(_zz_1650) + $signed(_zz_3994));
  assign _zz_15967 = ($signed(twiddle_factor_table_120_real) + $signed(twiddle_factor_table_120_imag));
  assign _zz_15968 = fixTo_1323_dout;
  assign _zz_15969 = ($signed(_zz_1780) - $signed(_zz_1779));
  assign _zz_15970 = ($signed(_zz_1779) + $signed(_zz_1780));
  assign _zz_15971 = _zz_15972[15 : 0];
  assign _zz_15972 = fixTo_1325_dout;
  assign _zz_15973 = _zz_15974[15 : 0];
  assign _zz_15974 = fixTo_1324_dout;
  assign _zz_15975 = _zz_15976;
  assign _zz_15976 = ($signed(_zz_15977) >>> _zz_4001);
  assign _zz_15977 = _zz_15978;
  assign _zz_15978 = ($signed(_zz_1651) - $signed(_zz_3998));
  assign _zz_15979 = _zz_15980;
  assign _zz_15980 = ($signed(_zz_15981) >>> _zz_4001);
  assign _zz_15981 = _zz_15982;
  assign _zz_15982 = ($signed(_zz_1652) - $signed(_zz_3999));
  assign _zz_15983 = _zz_15984;
  assign _zz_15984 = ($signed(_zz_15985) >>> _zz_4002);
  assign _zz_15985 = _zz_15986;
  assign _zz_15986 = ($signed(_zz_1651) + $signed(_zz_3998));
  assign _zz_15987 = _zz_15988;
  assign _zz_15988 = ($signed(_zz_15989) >>> _zz_4002);
  assign _zz_15989 = _zz_15990;
  assign _zz_15990 = ($signed(_zz_1652) + $signed(_zz_3999));
  assign _zz_15991 = ($signed(twiddle_factor_table_121_real) + $signed(twiddle_factor_table_121_imag));
  assign _zz_15992 = fixTo_1326_dout;
  assign _zz_15993 = ($signed(_zz_1782) - $signed(_zz_1781));
  assign _zz_15994 = ($signed(_zz_1781) + $signed(_zz_1782));
  assign _zz_15995 = _zz_15996[15 : 0];
  assign _zz_15996 = fixTo_1328_dout;
  assign _zz_15997 = _zz_15998[15 : 0];
  assign _zz_15998 = fixTo_1327_dout;
  assign _zz_15999 = _zz_16000;
  assign _zz_16000 = ($signed(_zz_16001) >>> _zz_4006);
  assign _zz_16001 = _zz_16002;
  assign _zz_16002 = ($signed(_zz_1653) - $signed(_zz_4003));
  assign _zz_16003 = _zz_16004;
  assign _zz_16004 = ($signed(_zz_16005) >>> _zz_4006);
  assign _zz_16005 = _zz_16006;
  assign _zz_16006 = ($signed(_zz_1654) - $signed(_zz_4004));
  assign _zz_16007 = _zz_16008;
  assign _zz_16008 = ($signed(_zz_16009) >>> _zz_4007);
  assign _zz_16009 = _zz_16010;
  assign _zz_16010 = ($signed(_zz_1653) + $signed(_zz_4003));
  assign _zz_16011 = _zz_16012;
  assign _zz_16012 = ($signed(_zz_16013) >>> _zz_4007);
  assign _zz_16013 = _zz_16014;
  assign _zz_16014 = ($signed(_zz_1654) + $signed(_zz_4004));
  assign _zz_16015 = ($signed(twiddle_factor_table_122_real) + $signed(twiddle_factor_table_122_imag));
  assign _zz_16016 = fixTo_1329_dout;
  assign _zz_16017 = ($signed(_zz_1784) - $signed(_zz_1783));
  assign _zz_16018 = ($signed(_zz_1783) + $signed(_zz_1784));
  assign _zz_16019 = _zz_16020[15 : 0];
  assign _zz_16020 = fixTo_1331_dout;
  assign _zz_16021 = _zz_16022[15 : 0];
  assign _zz_16022 = fixTo_1330_dout;
  assign _zz_16023 = _zz_16024;
  assign _zz_16024 = ($signed(_zz_16025) >>> _zz_4011);
  assign _zz_16025 = _zz_16026;
  assign _zz_16026 = ($signed(_zz_1655) - $signed(_zz_4008));
  assign _zz_16027 = _zz_16028;
  assign _zz_16028 = ($signed(_zz_16029) >>> _zz_4011);
  assign _zz_16029 = _zz_16030;
  assign _zz_16030 = ($signed(_zz_1656) - $signed(_zz_4009));
  assign _zz_16031 = _zz_16032;
  assign _zz_16032 = ($signed(_zz_16033) >>> _zz_4012);
  assign _zz_16033 = _zz_16034;
  assign _zz_16034 = ($signed(_zz_1655) + $signed(_zz_4008));
  assign _zz_16035 = _zz_16036;
  assign _zz_16036 = ($signed(_zz_16037) >>> _zz_4012);
  assign _zz_16037 = _zz_16038;
  assign _zz_16038 = ($signed(_zz_1656) + $signed(_zz_4009));
  assign _zz_16039 = ($signed(twiddle_factor_table_123_real) + $signed(twiddle_factor_table_123_imag));
  assign _zz_16040 = fixTo_1332_dout;
  assign _zz_16041 = ($signed(_zz_1786) - $signed(_zz_1785));
  assign _zz_16042 = ($signed(_zz_1785) + $signed(_zz_1786));
  assign _zz_16043 = _zz_16044[15 : 0];
  assign _zz_16044 = fixTo_1334_dout;
  assign _zz_16045 = _zz_16046[15 : 0];
  assign _zz_16046 = fixTo_1333_dout;
  assign _zz_16047 = _zz_16048;
  assign _zz_16048 = ($signed(_zz_16049) >>> _zz_4016);
  assign _zz_16049 = _zz_16050;
  assign _zz_16050 = ($signed(_zz_1657) - $signed(_zz_4013));
  assign _zz_16051 = _zz_16052;
  assign _zz_16052 = ($signed(_zz_16053) >>> _zz_4016);
  assign _zz_16053 = _zz_16054;
  assign _zz_16054 = ($signed(_zz_1658) - $signed(_zz_4014));
  assign _zz_16055 = _zz_16056;
  assign _zz_16056 = ($signed(_zz_16057) >>> _zz_4017);
  assign _zz_16057 = _zz_16058;
  assign _zz_16058 = ($signed(_zz_1657) + $signed(_zz_4013));
  assign _zz_16059 = _zz_16060;
  assign _zz_16060 = ($signed(_zz_16061) >>> _zz_4017);
  assign _zz_16061 = _zz_16062;
  assign _zz_16062 = ($signed(_zz_1658) + $signed(_zz_4014));
  assign _zz_16063 = ($signed(twiddle_factor_table_124_real) + $signed(twiddle_factor_table_124_imag));
  assign _zz_16064 = fixTo_1335_dout;
  assign _zz_16065 = ($signed(_zz_1788) - $signed(_zz_1787));
  assign _zz_16066 = ($signed(_zz_1787) + $signed(_zz_1788));
  assign _zz_16067 = _zz_16068[15 : 0];
  assign _zz_16068 = fixTo_1337_dout;
  assign _zz_16069 = _zz_16070[15 : 0];
  assign _zz_16070 = fixTo_1336_dout;
  assign _zz_16071 = _zz_16072;
  assign _zz_16072 = ($signed(_zz_16073) >>> _zz_4021);
  assign _zz_16073 = _zz_16074;
  assign _zz_16074 = ($signed(_zz_1659) - $signed(_zz_4018));
  assign _zz_16075 = _zz_16076;
  assign _zz_16076 = ($signed(_zz_16077) >>> _zz_4021);
  assign _zz_16077 = _zz_16078;
  assign _zz_16078 = ($signed(_zz_1660) - $signed(_zz_4019));
  assign _zz_16079 = _zz_16080;
  assign _zz_16080 = ($signed(_zz_16081) >>> _zz_4022);
  assign _zz_16081 = _zz_16082;
  assign _zz_16082 = ($signed(_zz_1659) + $signed(_zz_4018));
  assign _zz_16083 = _zz_16084;
  assign _zz_16084 = ($signed(_zz_16085) >>> _zz_4022);
  assign _zz_16085 = _zz_16086;
  assign _zz_16086 = ($signed(_zz_1660) + $signed(_zz_4019));
  assign _zz_16087 = ($signed(twiddle_factor_table_125_real) + $signed(twiddle_factor_table_125_imag));
  assign _zz_16088 = fixTo_1338_dout;
  assign _zz_16089 = ($signed(_zz_1790) - $signed(_zz_1789));
  assign _zz_16090 = ($signed(_zz_1789) + $signed(_zz_1790));
  assign _zz_16091 = _zz_16092[15 : 0];
  assign _zz_16092 = fixTo_1340_dout;
  assign _zz_16093 = _zz_16094[15 : 0];
  assign _zz_16094 = fixTo_1339_dout;
  assign _zz_16095 = _zz_16096;
  assign _zz_16096 = ($signed(_zz_16097) >>> _zz_4026);
  assign _zz_16097 = _zz_16098;
  assign _zz_16098 = ($signed(_zz_1661) - $signed(_zz_4023));
  assign _zz_16099 = _zz_16100;
  assign _zz_16100 = ($signed(_zz_16101) >>> _zz_4026);
  assign _zz_16101 = _zz_16102;
  assign _zz_16102 = ($signed(_zz_1662) - $signed(_zz_4024));
  assign _zz_16103 = _zz_16104;
  assign _zz_16104 = ($signed(_zz_16105) >>> _zz_4027);
  assign _zz_16105 = _zz_16106;
  assign _zz_16106 = ($signed(_zz_1661) + $signed(_zz_4023));
  assign _zz_16107 = _zz_16108;
  assign _zz_16108 = ($signed(_zz_16109) >>> _zz_4027);
  assign _zz_16109 = _zz_16110;
  assign _zz_16110 = ($signed(_zz_1662) + $signed(_zz_4024));
  assign _zz_16111 = ($signed(twiddle_factor_table_126_real) + $signed(twiddle_factor_table_126_imag));
  assign _zz_16112 = fixTo_1341_dout;
  assign _zz_16113 = ($signed(_zz_1792) - $signed(_zz_1791));
  assign _zz_16114 = ($signed(_zz_1791) + $signed(_zz_1792));
  assign _zz_16115 = _zz_16116[15 : 0];
  assign _zz_16116 = fixTo_1343_dout;
  assign _zz_16117 = _zz_16118[15 : 0];
  assign _zz_16118 = fixTo_1342_dout;
  assign _zz_16119 = _zz_16120;
  assign _zz_16120 = ($signed(_zz_16121) >>> _zz_4031);
  assign _zz_16121 = _zz_16122;
  assign _zz_16122 = ($signed(_zz_1663) - $signed(_zz_4028));
  assign _zz_16123 = _zz_16124;
  assign _zz_16124 = ($signed(_zz_16125) >>> _zz_4031);
  assign _zz_16125 = _zz_16126;
  assign _zz_16126 = ($signed(_zz_1664) - $signed(_zz_4029));
  assign _zz_16127 = _zz_16128;
  assign _zz_16128 = ($signed(_zz_16129) >>> _zz_4032);
  assign _zz_16129 = _zz_16130;
  assign _zz_16130 = ($signed(_zz_1663) + $signed(_zz_4028));
  assign _zz_16131 = _zz_16132;
  assign _zz_16132 = ($signed(_zz_16133) >>> _zz_4032);
  assign _zz_16133 = _zz_16134;
  assign _zz_16134 = ($signed(_zz_1664) + $signed(_zz_4029));
  assign _zz_16135 = _zz_4033;
  assign _zz_16136 = {3'd0, _zz_16135};
  SInt32fixTo23_8_ROUNDTOINF fixTo (
    .din     (_zz_4039[31:0]    ), //i
    .dout    (fixTo_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1 (
    .din     (_zz_4040[31:0]      ), //i
    .dout    (fixTo_1_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_2 (
    .din     (_zz_4041[31:0]      ), //i
    .dout    (fixTo_2_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_3 (
    .din     (_zz_4042[31:0]      ), //i
    .dout    (fixTo_3_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_4 (
    .din     (_zz_4043[31:0]      ), //i
    .dout    (fixTo_4_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_5 (
    .din     (_zz_4044[31:0]      ), //i
    .dout    (fixTo_5_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_6 (
    .din     (_zz_4045[31:0]      ), //i
    .dout    (fixTo_6_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_7 (
    .din     (_zz_4046[31:0]      ), //i
    .dout    (fixTo_7_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_8 (
    .din     (_zz_4047[31:0]      ), //i
    .dout    (fixTo_8_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_9 (
    .din     (_zz_4048[31:0]      ), //i
    .dout    (fixTo_9_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_10 (
    .din     (_zz_4049[31:0]       ), //i
    .dout    (fixTo_10_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_11 (
    .din     (_zz_4050[31:0]       ), //i
    .dout    (fixTo_11_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_12 (
    .din     (_zz_4051[31:0]       ), //i
    .dout    (fixTo_12_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_13 (
    .din     (_zz_4052[31:0]       ), //i
    .dout    (fixTo_13_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_14 (
    .din     (_zz_4053[31:0]       ), //i
    .dout    (fixTo_14_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_15 (
    .din     (_zz_4054[31:0]       ), //i
    .dout    (fixTo_15_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_16 (
    .din     (_zz_4055[31:0]       ), //i
    .dout    (fixTo_16_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_17 (
    .din     (_zz_4056[31:0]       ), //i
    .dout    (fixTo_17_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_18 (
    .din     (_zz_4057[31:0]       ), //i
    .dout    (fixTo_18_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_19 (
    .din     (_zz_4058[31:0]       ), //i
    .dout    (fixTo_19_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_20 (
    .din     (_zz_4059[31:0]       ), //i
    .dout    (fixTo_20_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_21 (
    .din     (_zz_4060[31:0]       ), //i
    .dout    (fixTo_21_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_22 (
    .din     (_zz_4061[31:0]       ), //i
    .dout    (fixTo_22_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_23 (
    .din     (_zz_4062[31:0]       ), //i
    .dout    (fixTo_23_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_24 (
    .din     (_zz_4063[31:0]       ), //i
    .dout    (fixTo_24_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_25 (
    .din     (_zz_4064[31:0]       ), //i
    .dout    (fixTo_25_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_26 (
    .din     (_zz_4065[31:0]       ), //i
    .dout    (fixTo_26_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_27 (
    .din     (_zz_4066[31:0]       ), //i
    .dout    (fixTo_27_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_28 (
    .din     (_zz_4067[31:0]       ), //i
    .dout    (fixTo_28_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_29 (
    .din     (_zz_4068[31:0]       ), //i
    .dout    (fixTo_29_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_30 (
    .din     (_zz_4069[31:0]       ), //i
    .dout    (fixTo_30_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_31 (
    .din     (_zz_4070[31:0]       ), //i
    .dout    (fixTo_31_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_32 (
    .din     (_zz_4071[31:0]       ), //i
    .dout    (fixTo_32_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_33 (
    .din     (_zz_4072[31:0]       ), //i
    .dout    (fixTo_33_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_34 (
    .din     (_zz_4073[31:0]       ), //i
    .dout    (fixTo_34_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_35 (
    .din     (_zz_4074[31:0]       ), //i
    .dout    (fixTo_35_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_36 (
    .din     (_zz_4075[31:0]       ), //i
    .dout    (fixTo_36_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_37 (
    .din     (_zz_4076[31:0]       ), //i
    .dout    (fixTo_37_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_38 (
    .din     (_zz_4077[31:0]       ), //i
    .dout    (fixTo_38_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_39 (
    .din     (_zz_4078[31:0]       ), //i
    .dout    (fixTo_39_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_40 (
    .din     (_zz_4079[31:0]       ), //i
    .dout    (fixTo_40_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_41 (
    .din     (_zz_4080[31:0]       ), //i
    .dout    (fixTo_41_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_42 (
    .din     (_zz_4081[31:0]       ), //i
    .dout    (fixTo_42_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_43 (
    .din     (_zz_4082[31:0]       ), //i
    .dout    (fixTo_43_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_44 (
    .din     (_zz_4083[31:0]       ), //i
    .dout    (fixTo_44_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_45 (
    .din     (_zz_4084[31:0]       ), //i
    .dout    (fixTo_45_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_46 (
    .din     (_zz_4085[31:0]       ), //i
    .dout    (fixTo_46_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_47 (
    .din     (_zz_4086[31:0]       ), //i
    .dout    (fixTo_47_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_48 (
    .din     (_zz_4087[31:0]       ), //i
    .dout    (fixTo_48_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_49 (
    .din     (_zz_4088[31:0]       ), //i
    .dout    (fixTo_49_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_50 (
    .din     (_zz_4089[31:0]       ), //i
    .dout    (fixTo_50_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_51 (
    .din     (_zz_4090[31:0]       ), //i
    .dout    (fixTo_51_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_52 (
    .din     (_zz_4091[31:0]       ), //i
    .dout    (fixTo_52_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_53 (
    .din     (_zz_4092[31:0]       ), //i
    .dout    (fixTo_53_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_54 (
    .din     (_zz_4093[31:0]       ), //i
    .dout    (fixTo_54_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_55 (
    .din     (_zz_4094[31:0]       ), //i
    .dout    (fixTo_55_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_56 (
    .din     (_zz_4095[31:0]       ), //i
    .dout    (fixTo_56_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_57 (
    .din     (_zz_4096[31:0]       ), //i
    .dout    (fixTo_57_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_58 (
    .din     (_zz_4097[31:0]       ), //i
    .dout    (fixTo_58_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_59 (
    .din     (_zz_4098[31:0]       ), //i
    .dout    (fixTo_59_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_60 (
    .din     (_zz_4099[31:0]       ), //i
    .dout    (fixTo_60_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_61 (
    .din     (_zz_4100[31:0]       ), //i
    .dout    (fixTo_61_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_62 (
    .din     (_zz_4101[31:0]       ), //i
    .dout    (fixTo_62_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_63 (
    .din     (_zz_4102[31:0]       ), //i
    .dout    (fixTo_63_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_64 (
    .din     (_zz_4103[31:0]       ), //i
    .dout    (fixTo_64_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_65 (
    .din     (_zz_4104[31:0]       ), //i
    .dout    (fixTo_65_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_66 (
    .din     (_zz_4105[31:0]       ), //i
    .dout    (fixTo_66_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_67 (
    .din     (_zz_4106[31:0]       ), //i
    .dout    (fixTo_67_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_68 (
    .din     (_zz_4107[31:0]       ), //i
    .dout    (fixTo_68_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_69 (
    .din     (_zz_4108[31:0]       ), //i
    .dout    (fixTo_69_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_70 (
    .din     (_zz_4109[31:0]       ), //i
    .dout    (fixTo_70_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_71 (
    .din     (_zz_4110[31:0]       ), //i
    .dout    (fixTo_71_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_72 (
    .din     (_zz_4111[31:0]       ), //i
    .dout    (fixTo_72_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_73 (
    .din     (_zz_4112[31:0]       ), //i
    .dout    (fixTo_73_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_74 (
    .din     (_zz_4113[31:0]       ), //i
    .dout    (fixTo_74_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_75 (
    .din     (_zz_4114[31:0]       ), //i
    .dout    (fixTo_75_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_76 (
    .din     (_zz_4115[31:0]       ), //i
    .dout    (fixTo_76_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_77 (
    .din     (_zz_4116[31:0]       ), //i
    .dout    (fixTo_77_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_78 (
    .din     (_zz_4117[31:0]       ), //i
    .dout    (fixTo_78_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_79 (
    .din     (_zz_4118[31:0]       ), //i
    .dout    (fixTo_79_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_80 (
    .din     (_zz_4119[31:0]       ), //i
    .dout    (fixTo_80_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_81 (
    .din     (_zz_4120[31:0]       ), //i
    .dout    (fixTo_81_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_82 (
    .din     (_zz_4121[31:0]       ), //i
    .dout    (fixTo_82_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_83 (
    .din     (_zz_4122[31:0]       ), //i
    .dout    (fixTo_83_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_84 (
    .din     (_zz_4123[31:0]       ), //i
    .dout    (fixTo_84_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_85 (
    .din     (_zz_4124[31:0]       ), //i
    .dout    (fixTo_85_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_86 (
    .din     (_zz_4125[31:0]       ), //i
    .dout    (fixTo_86_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_87 (
    .din     (_zz_4126[31:0]       ), //i
    .dout    (fixTo_87_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_88 (
    .din     (_zz_4127[31:0]       ), //i
    .dout    (fixTo_88_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_89 (
    .din     (_zz_4128[31:0]       ), //i
    .dout    (fixTo_89_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_90 (
    .din     (_zz_4129[31:0]       ), //i
    .dout    (fixTo_90_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_91 (
    .din     (_zz_4130[31:0]       ), //i
    .dout    (fixTo_91_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_92 (
    .din     (_zz_4131[31:0]       ), //i
    .dout    (fixTo_92_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_93 (
    .din     (_zz_4132[31:0]       ), //i
    .dout    (fixTo_93_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_94 (
    .din     (_zz_4133[31:0]       ), //i
    .dout    (fixTo_94_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_95 (
    .din     (_zz_4134[31:0]       ), //i
    .dout    (fixTo_95_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_96 (
    .din     (_zz_4135[31:0]       ), //i
    .dout    (fixTo_96_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_97 (
    .din     (_zz_4136[31:0]       ), //i
    .dout    (fixTo_97_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_98 (
    .din     (_zz_4137[31:0]       ), //i
    .dout    (fixTo_98_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_99 (
    .din     (_zz_4138[31:0]       ), //i
    .dout    (fixTo_99_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_100 (
    .din     (_zz_4139[31:0]        ), //i
    .dout    (fixTo_100_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_101 (
    .din     (_zz_4140[31:0]        ), //i
    .dout    (fixTo_101_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_102 (
    .din     (_zz_4141[31:0]        ), //i
    .dout    (fixTo_102_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_103 (
    .din     (_zz_4142[31:0]        ), //i
    .dout    (fixTo_103_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_104 (
    .din     (_zz_4143[31:0]        ), //i
    .dout    (fixTo_104_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_105 (
    .din     (_zz_4144[31:0]        ), //i
    .dout    (fixTo_105_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_106 (
    .din     (_zz_4145[31:0]        ), //i
    .dout    (fixTo_106_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_107 (
    .din     (_zz_4146[31:0]        ), //i
    .dout    (fixTo_107_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_108 (
    .din     (_zz_4147[31:0]        ), //i
    .dout    (fixTo_108_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_109 (
    .din     (_zz_4148[31:0]        ), //i
    .dout    (fixTo_109_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_110 (
    .din     (_zz_4149[31:0]        ), //i
    .dout    (fixTo_110_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_111 (
    .din     (_zz_4150[31:0]        ), //i
    .dout    (fixTo_111_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_112 (
    .din     (_zz_4151[31:0]        ), //i
    .dout    (fixTo_112_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_113 (
    .din     (_zz_4152[31:0]        ), //i
    .dout    (fixTo_113_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_114 (
    .din     (_zz_4153[31:0]        ), //i
    .dout    (fixTo_114_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_115 (
    .din     (_zz_4154[31:0]        ), //i
    .dout    (fixTo_115_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_116 (
    .din     (_zz_4155[31:0]        ), //i
    .dout    (fixTo_116_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_117 (
    .din     (_zz_4156[31:0]        ), //i
    .dout    (fixTo_117_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_118 (
    .din     (_zz_4157[31:0]        ), //i
    .dout    (fixTo_118_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_119 (
    .din     (_zz_4158[31:0]        ), //i
    .dout    (fixTo_119_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_120 (
    .din     (_zz_4159[31:0]        ), //i
    .dout    (fixTo_120_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_121 (
    .din     (_zz_4160[31:0]        ), //i
    .dout    (fixTo_121_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_122 (
    .din     (_zz_4161[31:0]        ), //i
    .dout    (fixTo_122_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_123 (
    .din     (_zz_4162[31:0]        ), //i
    .dout    (fixTo_123_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_124 (
    .din     (_zz_4163[31:0]        ), //i
    .dout    (fixTo_124_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_125 (
    .din     (_zz_4164[31:0]        ), //i
    .dout    (fixTo_125_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_126 (
    .din     (_zz_4165[31:0]        ), //i
    .dout    (fixTo_126_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_127 (
    .din     (_zz_4166[31:0]        ), //i
    .dout    (fixTo_127_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_128 (
    .din     (_zz_4167[31:0]        ), //i
    .dout    (fixTo_128_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_129 (
    .din     (_zz_4168[31:0]        ), //i
    .dout    (fixTo_129_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_130 (
    .din     (_zz_4169[31:0]        ), //i
    .dout    (fixTo_130_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_131 (
    .din     (_zz_4170[31:0]        ), //i
    .dout    (fixTo_131_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_132 (
    .din     (_zz_4171[31:0]        ), //i
    .dout    (fixTo_132_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_133 (
    .din     (_zz_4172[31:0]        ), //i
    .dout    (fixTo_133_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_134 (
    .din     (_zz_4173[31:0]        ), //i
    .dout    (fixTo_134_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_135 (
    .din     (_zz_4174[31:0]        ), //i
    .dout    (fixTo_135_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_136 (
    .din     (_zz_4175[31:0]        ), //i
    .dout    (fixTo_136_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_137 (
    .din     (_zz_4176[31:0]        ), //i
    .dout    (fixTo_137_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_138 (
    .din     (_zz_4177[31:0]        ), //i
    .dout    (fixTo_138_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_139 (
    .din     (_zz_4178[31:0]        ), //i
    .dout    (fixTo_139_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_140 (
    .din     (_zz_4179[31:0]        ), //i
    .dout    (fixTo_140_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_141 (
    .din     (_zz_4180[31:0]        ), //i
    .dout    (fixTo_141_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_142 (
    .din     (_zz_4181[31:0]        ), //i
    .dout    (fixTo_142_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_143 (
    .din     (_zz_4182[31:0]        ), //i
    .dout    (fixTo_143_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_144 (
    .din     (_zz_4183[31:0]        ), //i
    .dout    (fixTo_144_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_145 (
    .din     (_zz_4184[31:0]        ), //i
    .dout    (fixTo_145_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_146 (
    .din     (_zz_4185[31:0]        ), //i
    .dout    (fixTo_146_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_147 (
    .din     (_zz_4186[31:0]        ), //i
    .dout    (fixTo_147_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_148 (
    .din     (_zz_4187[31:0]        ), //i
    .dout    (fixTo_148_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_149 (
    .din     (_zz_4188[31:0]        ), //i
    .dout    (fixTo_149_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_150 (
    .din     (_zz_4189[31:0]        ), //i
    .dout    (fixTo_150_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_151 (
    .din     (_zz_4190[31:0]        ), //i
    .dout    (fixTo_151_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_152 (
    .din     (_zz_4191[31:0]        ), //i
    .dout    (fixTo_152_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_153 (
    .din     (_zz_4192[31:0]        ), //i
    .dout    (fixTo_153_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_154 (
    .din     (_zz_4193[31:0]        ), //i
    .dout    (fixTo_154_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_155 (
    .din     (_zz_4194[31:0]        ), //i
    .dout    (fixTo_155_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_156 (
    .din     (_zz_4195[31:0]        ), //i
    .dout    (fixTo_156_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_157 (
    .din     (_zz_4196[31:0]        ), //i
    .dout    (fixTo_157_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_158 (
    .din     (_zz_4197[31:0]        ), //i
    .dout    (fixTo_158_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_159 (
    .din     (_zz_4198[31:0]        ), //i
    .dout    (fixTo_159_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_160 (
    .din     (_zz_4199[31:0]        ), //i
    .dout    (fixTo_160_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_161 (
    .din     (_zz_4200[31:0]        ), //i
    .dout    (fixTo_161_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_162 (
    .din     (_zz_4201[31:0]        ), //i
    .dout    (fixTo_162_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_163 (
    .din     (_zz_4202[31:0]        ), //i
    .dout    (fixTo_163_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_164 (
    .din     (_zz_4203[31:0]        ), //i
    .dout    (fixTo_164_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_165 (
    .din     (_zz_4204[31:0]        ), //i
    .dout    (fixTo_165_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_166 (
    .din     (_zz_4205[31:0]        ), //i
    .dout    (fixTo_166_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_167 (
    .din     (_zz_4206[31:0]        ), //i
    .dout    (fixTo_167_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_168 (
    .din     (_zz_4207[31:0]        ), //i
    .dout    (fixTo_168_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_169 (
    .din     (_zz_4208[31:0]        ), //i
    .dout    (fixTo_169_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_170 (
    .din     (_zz_4209[31:0]        ), //i
    .dout    (fixTo_170_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_171 (
    .din     (_zz_4210[31:0]        ), //i
    .dout    (fixTo_171_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_172 (
    .din     (_zz_4211[31:0]        ), //i
    .dout    (fixTo_172_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_173 (
    .din     (_zz_4212[31:0]        ), //i
    .dout    (fixTo_173_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_174 (
    .din     (_zz_4213[31:0]        ), //i
    .dout    (fixTo_174_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_175 (
    .din     (_zz_4214[31:0]        ), //i
    .dout    (fixTo_175_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_176 (
    .din     (_zz_4215[31:0]        ), //i
    .dout    (fixTo_176_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_177 (
    .din     (_zz_4216[31:0]        ), //i
    .dout    (fixTo_177_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_178 (
    .din     (_zz_4217[31:0]        ), //i
    .dout    (fixTo_178_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_179 (
    .din     (_zz_4218[31:0]        ), //i
    .dout    (fixTo_179_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_180 (
    .din     (_zz_4219[31:0]        ), //i
    .dout    (fixTo_180_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_181 (
    .din     (_zz_4220[31:0]        ), //i
    .dout    (fixTo_181_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_182 (
    .din     (_zz_4221[31:0]        ), //i
    .dout    (fixTo_182_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_183 (
    .din     (_zz_4222[31:0]        ), //i
    .dout    (fixTo_183_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_184 (
    .din     (_zz_4223[31:0]        ), //i
    .dout    (fixTo_184_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_185 (
    .din     (_zz_4224[31:0]        ), //i
    .dout    (fixTo_185_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_186 (
    .din     (_zz_4225[31:0]        ), //i
    .dout    (fixTo_186_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_187 (
    .din     (_zz_4226[31:0]        ), //i
    .dout    (fixTo_187_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_188 (
    .din     (_zz_4227[31:0]        ), //i
    .dout    (fixTo_188_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_189 (
    .din     (_zz_4228[31:0]        ), //i
    .dout    (fixTo_189_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_190 (
    .din     (_zz_4229[31:0]        ), //i
    .dout    (fixTo_190_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_191 (
    .din     (_zz_4230[31:0]        ), //i
    .dout    (fixTo_191_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_192 (
    .din     (_zz_4231[31:0]        ), //i
    .dout    (fixTo_192_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_193 (
    .din     (_zz_4232[31:0]        ), //i
    .dout    (fixTo_193_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_194 (
    .din     (_zz_4233[31:0]        ), //i
    .dout    (fixTo_194_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_195 (
    .din     (_zz_4234[31:0]        ), //i
    .dout    (fixTo_195_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_196 (
    .din     (_zz_4235[31:0]        ), //i
    .dout    (fixTo_196_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_197 (
    .din     (_zz_4236[31:0]        ), //i
    .dout    (fixTo_197_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_198 (
    .din     (_zz_4237[31:0]        ), //i
    .dout    (fixTo_198_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_199 (
    .din     (_zz_4238[31:0]        ), //i
    .dout    (fixTo_199_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_200 (
    .din     (_zz_4239[31:0]        ), //i
    .dout    (fixTo_200_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_201 (
    .din     (_zz_4240[31:0]        ), //i
    .dout    (fixTo_201_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_202 (
    .din     (_zz_4241[31:0]        ), //i
    .dout    (fixTo_202_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_203 (
    .din     (_zz_4242[31:0]        ), //i
    .dout    (fixTo_203_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_204 (
    .din     (_zz_4243[31:0]        ), //i
    .dout    (fixTo_204_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_205 (
    .din     (_zz_4244[31:0]        ), //i
    .dout    (fixTo_205_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_206 (
    .din     (_zz_4245[31:0]        ), //i
    .dout    (fixTo_206_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_207 (
    .din     (_zz_4246[31:0]        ), //i
    .dout    (fixTo_207_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_208 (
    .din     (_zz_4247[31:0]        ), //i
    .dout    (fixTo_208_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_209 (
    .din     (_zz_4248[31:0]        ), //i
    .dout    (fixTo_209_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_210 (
    .din     (_zz_4249[31:0]        ), //i
    .dout    (fixTo_210_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_211 (
    .din     (_zz_4250[31:0]        ), //i
    .dout    (fixTo_211_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_212 (
    .din     (_zz_4251[31:0]        ), //i
    .dout    (fixTo_212_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_213 (
    .din     (_zz_4252[31:0]        ), //i
    .dout    (fixTo_213_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_214 (
    .din     (_zz_4253[31:0]        ), //i
    .dout    (fixTo_214_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_215 (
    .din     (_zz_4254[31:0]        ), //i
    .dout    (fixTo_215_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_216 (
    .din     (_zz_4255[31:0]        ), //i
    .dout    (fixTo_216_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_217 (
    .din     (_zz_4256[31:0]        ), //i
    .dout    (fixTo_217_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_218 (
    .din     (_zz_4257[31:0]        ), //i
    .dout    (fixTo_218_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_219 (
    .din     (_zz_4258[31:0]        ), //i
    .dout    (fixTo_219_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_220 (
    .din     (_zz_4259[31:0]        ), //i
    .dout    (fixTo_220_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_221 (
    .din     (_zz_4260[31:0]        ), //i
    .dout    (fixTo_221_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_222 (
    .din     (_zz_4261[31:0]        ), //i
    .dout    (fixTo_222_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_223 (
    .din     (_zz_4262[31:0]        ), //i
    .dout    (fixTo_223_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_224 (
    .din     (_zz_4263[31:0]        ), //i
    .dout    (fixTo_224_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_225 (
    .din     (_zz_4264[31:0]        ), //i
    .dout    (fixTo_225_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_226 (
    .din     (_zz_4265[31:0]        ), //i
    .dout    (fixTo_226_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_227 (
    .din     (_zz_4266[31:0]        ), //i
    .dout    (fixTo_227_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_228 (
    .din     (_zz_4267[31:0]        ), //i
    .dout    (fixTo_228_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_229 (
    .din     (_zz_4268[31:0]        ), //i
    .dout    (fixTo_229_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_230 (
    .din     (_zz_4269[31:0]        ), //i
    .dout    (fixTo_230_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_231 (
    .din     (_zz_4270[31:0]        ), //i
    .dout    (fixTo_231_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_232 (
    .din     (_zz_4271[31:0]        ), //i
    .dout    (fixTo_232_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_233 (
    .din     (_zz_4272[31:0]        ), //i
    .dout    (fixTo_233_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_234 (
    .din     (_zz_4273[31:0]        ), //i
    .dout    (fixTo_234_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_235 (
    .din     (_zz_4274[31:0]        ), //i
    .dout    (fixTo_235_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_236 (
    .din     (_zz_4275[31:0]        ), //i
    .dout    (fixTo_236_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_237 (
    .din     (_zz_4276[31:0]        ), //i
    .dout    (fixTo_237_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_238 (
    .din     (_zz_4277[31:0]        ), //i
    .dout    (fixTo_238_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_239 (
    .din     (_zz_4278[31:0]        ), //i
    .dout    (fixTo_239_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_240 (
    .din     (_zz_4279[31:0]        ), //i
    .dout    (fixTo_240_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_241 (
    .din     (_zz_4280[31:0]        ), //i
    .dout    (fixTo_241_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_242 (
    .din     (_zz_4281[31:0]        ), //i
    .dout    (fixTo_242_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_243 (
    .din     (_zz_4282[31:0]        ), //i
    .dout    (fixTo_243_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_244 (
    .din     (_zz_4283[31:0]        ), //i
    .dout    (fixTo_244_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_245 (
    .din     (_zz_4284[31:0]        ), //i
    .dout    (fixTo_245_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_246 (
    .din     (_zz_4285[31:0]        ), //i
    .dout    (fixTo_246_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_247 (
    .din     (_zz_4286[31:0]        ), //i
    .dout    (fixTo_247_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_248 (
    .din     (_zz_4287[31:0]        ), //i
    .dout    (fixTo_248_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_249 (
    .din     (_zz_4288[31:0]        ), //i
    .dout    (fixTo_249_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_250 (
    .din     (_zz_4289[31:0]        ), //i
    .dout    (fixTo_250_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_251 (
    .din     (_zz_4290[31:0]        ), //i
    .dout    (fixTo_251_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_252 (
    .din     (_zz_4291[31:0]        ), //i
    .dout    (fixTo_252_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_253 (
    .din     (_zz_4292[31:0]        ), //i
    .dout    (fixTo_253_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_254 (
    .din     (_zz_4293[31:0]        ), //i
    .dout    (fixTo_254_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_255 (
    .din     (_zz_4294[31:0]        ), //i
    .dout    (fixTo_255_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_256 (
    .din     (_zz_4295[31:0]        ), //i
    .dout    (fixTo_256_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_257 (
    .din     (_zz_4296[31:0]        ), //i
    .dout    (fixTo_257_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_258 (
    .din     (_zz_4297[31:0]        ), //i
    .dout    (fixTo_258_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_259 (
    .din     (_zz_4298[31:0]        ), //i
    .dout    (fixTo_259_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_260 (
    .din     (_zz_4299[31:0]        ), //i
    .dout    (fixTo_260_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_261 (
    .din     (_zz_4300[31:0]        ), //i
    .dout    (fixTo_261_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_262 (
    .din     (_zz_4301[31:0]        ), //i
    .dout    (fixTo_262_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_263 (
    .din     (_zz_4302[31:0]        ), //i
    .dout    (fixTo_263_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_264 (
    .din     (_zz_4303[31:0]        ), //i
    .dout    (fixTo_264_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_265 (
    .din     (_zz_4304[31:0]        ), //i
    .dout    (fixTo_265_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_266 (
    .din     (_zz_4305[31:0]        ), //i
    .dout    (fixTo_266_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_267 (
    .din     (_zz_4306[31:0]        ), //i
    .dout    (fixTo_267_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_268 (
    .din     (_zz_4307[31:0]        ), //i
    .dout    (fixTo_268_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_269 (
    .din     (_zz_4308[31:0]        ), //i
    .dout    (fixTo_269_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_270 (
    .din     (_zz_4309[31:0]        ), //i
    .dout    (fixTo_270_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_271 (
    .din     (_zz_4310[31:0]        ), //i
    .dout    (fixTo_271_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_272 (
    .din     (_zz_4311[31:0]        ), //i
    .dout    (fixTo_272_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_273 (
    .din     (_zz_4312[31:0]        ), //i
    .dout    (fixTo_273_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_274 (
    .din     (_zz_4313[31:0]        ), //i
    .dout    (fixTo_274_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_275 (
    .din     (_zz_4314[31:0]        ), //i
    .dout    (fixTo_275_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_276 (
    .din     (_zz_4315[31:0]        ), //i
    .dout    (fixTo_276_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_277 (
    .din     (_zz_4316[31:0]        ), //i
    .dout    (fixTo_277_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_278 (
    .din     (_zz_4317[31:0]        ), //i
    .dout    (fixTo_278_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_279 (
    .din     (_zz_4318[31:0]        ), //i
    .dout    (fixTo_279_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_280 (
    .din     (_zz_4319[31:0]        ), //i
    .dout    (fixTo_280_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_281 (
    .din     (_zz_4320[31:0]        ), //i
    .dout    (fixTo_281_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_282 (
    .din     (_zz_4321[31:0]        ), //i
    .dout    (fixTo_282_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_283 (
    .din     (_zz_4322[31:0]        ), //i
    .dout    (fixTo_283_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_284 (
    .din     (_zz_4323[31:0]        ), //i
    .dout    (fixTo_284_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_285 (
    .din     (_zz_4324[31:0]        ), //i
    .dout    (fixTo_285_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_286 (
    .din     (_zz_4325[31:0]        ), //i
    .dout    (fixTo_286_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_287 (
    .din     (_zz_4326[31:0]        ), //i
    .dout    (fixTo_287_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_288 (
    .din     (_zz_4327[31:0]        ), //i
    .dout    (fixTo_288_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_289 (
    .din     (_zz_4328[31:0]        ), //i
    .dout    (fixTo_289_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_290 (
    .din     (_zz_4329[31:0]        ), //i
    .dout    (fixTo_290_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_291 (
    .din     (_zz_4330[31:0]        ), //i
    .dout    (fixTo_291_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_292 (
    .din     (_zz_4331[31:0]        ), //i
    .dout    (fixTo_292_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_293 (
    .din     (_zz_4332[31:0]        ), //i
    .dout    (fixTo_293_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_294 (
    .din     (_zz_4333[31:0]        ), //i
    .dout    (fixTo_294_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_295 (
    .din     (_zz_4334[31:0]        ), //i
    .dout    (fixTo_295_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_296 (
    .din     (_zz_4335[31:0]        ), //i
    .dout    (fixTo_296_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_297 (
    .din     (_zz_4336[31:0]        ), //i
    .dout    (fixTo_297_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_298 (
    .din     (_zz_4337[31:0]        ), //i
    .dout    (fixTo_298_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_299 (
    .din     (_zz_4338[31:0]        ), //i
    .dout    (fixTo_299_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_300 (
    .din     (_zz_4339[31:0]        ), //i
    .dout    (fixTo_300_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_301 (
    .din     (_zz_4340[31:0]        ), //i
    .dout    (fixTo_301_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_302 (
    .din     (_zz_4341[31:0]        ), //i
    .dout    (fixTo_302_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_303 (
    .din     (_zz_4342[31:0]        ), //i
    .dout    (fixTo_303_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_304 (
    .din     (_zz_4343[31:0]        ), //i
    .dout    (fixTo_304_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_305 (
    .din     (_zz_4344[31:0]        ), //i
    .dout    (fixTo_305_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_306 (
    .din     (_zz_4345[31:0]        ), //i
    .dout    (fixTo_306_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_307 (
    .din     (_zz_4346[31:0]        ), //i
    .dout    (fixTo_307_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_308 (
    .din     (_zz_4347[31:0]        ), //i
    .dout    (fixTo_308_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_309 (
    .din     (_zz_4348[31:0]        ), //i
    .dout    (fixTo_309_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_310 (
    .din     (_zz_4349[31:0]        ), //i
    .dout    (fixTo_310_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_311 (
    .din     (_zz_4350[31:0]        ), //i
    .dout    (fixTo_311_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_312 (
    .din     (_zz_4351[31:0]        ), //i
    .dout    (fixTo_312_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_313 (
    .din     (_zz_4352[31:0]        ), //i
    .dout    (fixTo_313_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_314 (
    .din     (_zz_4353[31:0]        ), //i
    .dout    (fixTo_314_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_315 (
    .din     (_zz_4354[31:0]        ), //i
    .dout    (fixTo_315_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_316 (
    .din     (_zz_4355[31:0]        ), //i
    .dout    (fixTo_316_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_317 (
    .din     (_zz_4356[31:0]        ), //i
    .dout    (fixTo_317_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_318 (
    .din     (_zz_4357[31:0]        ), //i
    .dout    (fixTo_318_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_319 (
    .din     (_zz_4358[31:0]        ), //i
    .dout    (fixTo_319_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_320 (
    .din     (_zz_4359[31:0]        ), //i
    .dout    (fixTo_320_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_321 (
    .din     (_zz_4360[31:0]        ), //i
    .dout    (fixTo_321_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_322 (
    .din     (_zz_4361[31:0]        ), //i
    .dout    (fixTo_322_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_323 (
    .din     (_zz_4362[31:0]        ), //i
    .dout    (fixTo_323_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_324 (
    .din     (_zz_4363[31:0]        ), //i
    .dout    (fixTo_324_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_325 (
    .din     (_zz_4364[31:0]        ), //i
    .dout    (fixTo_325_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_326 (
    .din     (_zz_4365[31:0]        ), //i
    .dout    (fixTo_326_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_327 (
    .din     (_zz_4366[31:0]        ), //i
    .dout    (fixTo_327_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_328 (
    .din     (_zz_4367[31:0]        ), //i
    .dout    (fixTo_328_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_329 (
    .din     (_zz_4368[31:0]        ), //i
    .dout    (fixTo_329_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_330 (
    .din     (_zz_4369[31:0]        ), //i
    .dout    (fixTo_330_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_331 (
    .din     (_zz_4370[31:0]        ), //i
    .dout    (fixTo_331_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_332 (
    .din     (_zz_4371[31:0]        ), //i
    .dout    (fixTo_332_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_333 (
    .din     (_zz_4372[31:0]        ), //i
    .dout    (fixTo_333_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_334 (
    .din     (_zz_4373[31:0]        ), //i
    .dout    (fixTo_334_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_335 (
    .din     (_zz_4374[31:0]        ), //i
    .dout    (fixTo_335_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_336 (
    .din     (_zz_4375[31:0]        ), //i
    .dout    (fixTo_336_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_337 (
    .din     (_zz_4376[31:0]        ), //i
    .dout    (fixTo_337_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_338 (
    .din     (_zz_4377[31:0]        ), //i
    .dout    (fixTo_338_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_339 (
    .din     (_zz_4378[31:0]        ), //i
    .dout    (fixTo_339_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_340 (
    .din     (_zz_4379[31:0]        ), //i
    .dout    (fixTo_340_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_341 (
    .din     (_zz_4380[31:0]        ), //i
    .dout    (fixTo_341_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_342 (
    .din     (_zz_4381[31:0]        ), //i
    .dout    (fixTo_342_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_343 (
    .din     (_zz_4382[31:0]        ), //i
    .dout    (fixTo_343_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_344 (
    .din     (_zz_4383[31:0]        ), //i
    .dout    (fixTo_344_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_345 (
    .din     (_zz_4384[31:0]        ), //i
    .dout    (fixTo_345_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_346 (
    .din     (_zz_4385[31:0]        ), //i
    .dout    (fixTo_346_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_347 (
    .din     (_zz_4386[31:0]        ), //i
    .dout    (fixTo_347_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_348 (
    .din     (_zz_4387[31:0]        ), //i
    .dout    (fixTo_348_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_349 (
    .din     (_zz_4388[31:0]        ), //i
    .dout    (fixTo_349_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_350 (
    .din     (_zz_4389[31:0]        ), //i
    .dout    (fixTo_350_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_351 (
    .din     (_zz_4390[31:0]        ), //i
    .dout    (fixTo_351_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_352 (
    .din     (_zz_4391[31:0]        ), //i
    .dout    (fixTo_352_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_353 (
    .din     (_zz_4392[31:0]        ), //i
    .dout    (fixTo_353_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_354 (
    .din     (_zz_4393[31:0]        ), //i
    .dout    (fixTo_354_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_355 (
    .din     (_zz_4394[31:0]        ), //i
    .dout    (fixTo_355_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_356 (
    .din     (_zz_4395[31:0]        ), //i
    .dout    (fixTo_356_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_357 (
    .din     (_zz_4396[31:0]        ), //i
    .dout    (fixTo_357_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_358 (
    .din     (_zz_4397[31:0]        ), //i
    .dout    (fixTo_358_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_359 (
    .din     (_zz_4398[31:0]        ), //i
    .dout    (fixTo_359_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_360 (
    .din     (_zz_4399[31:0]        ), //i
    .dout    (fixTo_360_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_361 (
    .din     (_zz_4400[31:0]        ), //i
    .dout    (fixTo_361_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_362 (
    .din     (_zz_4401[31:0]        ), //i
    .dout    (fixTo_362_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_363 (
    .din     (_zz_4402[31:0]        ), //i
    .dout    (fixTo_363_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_364 (
    .din     (_zz_4403[31:0]        ), //i
    .dout    (fixTo_364_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_365 (
    .din     (_zz_4404[31:0]        ), //i
    .dout    (fixTo_365_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_366 (
    .din     (_zz_4405[31:0]        ), //i
    .dout    (fixTo_366_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_367 (
    .din     (_zz_4406[31:0]        ), //i
    .dout    (fixTo_367_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_368 (
    .din     (_zz_4407[31:0]        ), //i
    .dout    (fixTo_368_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_369 (
    .din     (_zz_4408[31:0]        ), //i
    .dout    (fixTo_369_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_370 (
    .din     (_zz_4409[31:0]        ), //i
    .dout    (fixTo_370_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_371 (
    .din     (_zz_4410[31:0]        ), //i
    .dout    (fixTo_371_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_372 (
    .din     (_zz_4411[31:0]        ), //i
    .dout    (fixTo_372_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_373 (
    .din     (_zz_4412[31:0]        ), //i
    .dout    (fixTo_373_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_374 (
    .din     (_zz_4413[31:0]        ), //i
    .dout    (fixTo_374_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_375 (
    .din     (_zz_4414[31:0]        ), //i
    .dout    (fixTo_375_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_376 (
    .din     (_zz_4415[31:0]        ), //i
    .dout    (fixTo_376_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_377 (
    .din     (_zz_4416[31:0]        ), //i
    .dout    (fixTo_377_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_378 (
    .din     (_zz_4417[31:0]        ), //i
    .dout    (fixTo_378_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_379 (
    .din     (_zz_4418[31:0]        ), //i
    .dout    (fixTo_379_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_380 (
    .din     (_zz_4419[31:0]        ), //i
    .dout    (fixTo_380_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_381 (
    .din     (_zz_4420[31:0]        ), //i
    .dout    (fixTo_381_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_382 (
    .din     (_zz_4421[31:0]        ), //i
    .dout    (fixTo_382_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_383 (
    .din     (_zz_4422[31:0]        ), //i
    .dout    (fixTo_383_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_384 (
    .din     (_zz_4423[31:0]        ), //i
    .dout    (fixTo_384_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_385 (
    .din     (_zz_4424[31:0]        ), //i
    .dout    (fixTo_385_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_386 (
    .din     (_zz_4425[31:0]        ), //i
    .dout    (fixTo_386_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_387 (
    .din     (_zz_4426[31:0]        ), //i
    .dout    (fixTo_387_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_388 (
    .din     (_zz_4427[31:0]        ), //i
    .dout    (fixTo_388_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_389 (
    .din     (_zz_4428[31:0]        ), //i
    .dout    (fixTo_389_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_390 (
    .din     (_zz_4429[31:0]        ), //i
    .dout    (fixTo_390_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_391 (
    .din     (_zz_4430[31:0]        ), //i
    .dout    (fixTo_391_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_392 (
    .din     (_zz_4431[31:0]        ), //i
    .dout    (fixTo_392_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_393 (
    .din     (_zz_4432[31:0]        ), //i
    .dout    (fixTo_393_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_394 (
    .din     (_zz_4433[31:0]        ), //i
    .dout    (fixTo_394_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_395 (
    .din     (_zz_4434[31:0]        ), //i
    .dout    (fixTo_395_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_396 (
    .din     (_zz_4435[31:0]        ), //i
    .dout    (fixTo_396_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_397 (
    .din     (_zz_4436[31:0]        ), //i
    .dout    (fixTo_397_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_398 (
    .din     (_zz_4437[31:0]        ), //i
    .dout    (fixTo_398_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_399 (
    .din     (_zz_4438[31:0]        ), //i
    .dout    (fixTo_399_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_400 (
    .din     (_zz_4439[31:0]        ), //i
    .dout    (fixTo_400_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_401 (
    .din     (_zz_4440[31:0]        ), //i
    .dout    (fixTo_401_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_402 (
    .din     (_zz_4441[31:0]        ), //i
    .dout    (fixTo_402_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_403 (
    .din     (_zz_4442[31:0]        ), //i
    .dout    (fixTo_403_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_404 (
    .din     (_zz_4443[31:0]        ), //i
    .dout    (fixTo_404_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_405 (
    .din     (_zz_4444[31:0]        ), //i
    .dout    (fixTo_405_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_406 (
    .din     (_zz_4445[31:0]        ), //i
    .dout    (fixTo_406_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_407 (
    .din     (_zz_4446[31:0]        ), //i
    .dout    (fixTo_407_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_408 (
    .din     (_zz_4447[31:0]        ), //i
    .dout    (fixTo_408_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_409 (
    .din     (_zz_4448[31:0]        ), //i
    .dout    (fixTo_409_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_410 (
    .din     (_zz_4449[31:0]        ), //i
    .dout    (fixTo_410_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_411 (
    .din     (_zz_4450[31:0]        ), //i
    .dout    (fixTo_411_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_412 (
    .din     (_zz_4451[31:0]        ), //i
    .dout    (fixTo_412_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_413 (
    .din     (_zz_4452[31:0]        ), //i
    .dout    (fixTo_413_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_414 (
    .din     (_zz_4453[31:0]        ), //i
    .dout    (fixTo_414_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_415 (
    .din     (_zz_4454[31:0]        ), //i
    .dout    (fixTo_415_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_416 (
    .din     (_zz_4455[31:0]        ), //i
    .dout    (fixTo_416_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_417 (
    .din     (_zz_4456[31:0]        ), //i
    .dout    (fixTo_417_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_418 (
    .din     (_zz_4457[31:0]        ), //i
    .dout    (fixTo_418_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_419 (
    .din     (_zz_4458[31:0]        ), //i
    .dout    (fixTo_419_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_420 (
    .din     (_zz_4459[31:0]        ), //i
    .dout    (fixTo_420_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_421 (
    .din     (_zz_4460[31:0]        ), //i
    .dout    (fixTo_421_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_422 (
    .din     (_zz_4461[31:0]        ), //i
    .dout    (fixTo_422_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_423 (
    .din     (_zz_4462[31:0]        ), //i
    .dout    (fixTo_423_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_424 (
    .din     (_zz_4463[31:0]        ), //i
    .dout    (fixTo_424_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_425 (
    .din     (_zz_4464[31:0]        ), //i
    .dout    (fixTo_425_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_426 (
    .din     (_zz_4465[31:0]        ), //i
    .dout    (fixTo_426_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_427 (
    .din     (_zz_4466[31:0]        ), //i
    .dout    (fixTo_427_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_428 (
    .din     (_zz_4467[31:0]        ), //i
    .dout    (fixTo_428_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_429 (
    .din     (_zz_4468[31:0]        ), //i
    .dout    (fixTo_429_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_430 (
    .din     (_zz_4469[31:0]        ), //i
    .dout    (fixTo_430_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_431 (
    .din     (_zz_4470[31:0]        ), //i
    .dout    (fixTo_431_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_432 (
    .din     (_zz_4471[31:0]        ), //i
    .dout    (fixTo_432_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_433 (
    .din     (_zz_4472[31:0]        ), //i
    .dout    (fixTo_433_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_434 (
    .din     (_zz_4473[31:0]        ), //i
    .dout    (fixTo_434_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_435 (
    .din     (_zz_4474[31:0]        ), //i
    .dout    (fixTo_435_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_436 (
    .din     (_zz_4475[31:0]        ), //i
    .dout    (fixTo_436_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_437 (
    .din     (_zz_4476[31:0]        ), //i
    .dout    (fixTo_437_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_438 (
    .din     (_zz_4477[31:0]        ), //i
    .dout    (fixTo_438_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_439 (
    .din     (_zz_4478[31:0]        ), //i
    .dout    (fixTo_439_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_440 (
    .din     (_zz_4479[31:0]        ), //i
    .dout    (fixTo_440_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_441 (
    .din     (_zz_4480[31:0]        ), //i
    .dout    (fixTo_441_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_442 (
    .din     (_zz_4481[31:0]        ), //i
    .dout    (fixTo_442_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_443 (
    .din     (_zz_4482[31:0]        ), //i
    .dout    (fixTo_443_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_444 (
    .din     (_zz_4483[31:0]        ), //i
    .dout    (fixTo_444_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_445 (
    .din     (_zz_4484[31:0]        ), //i
    .dout    (fixTo_445_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_446 (
    .din     (_zz_4485[31:0]        ), //i
    .dout    (fixTo_446_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_447 (
    .din     (_zz_4486[31:0]        ), //i
    .dout    (fixTo_447_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_448 (
    .din     (_zz_4487[31:0]        ), //i
    .dout    (fixTo_448_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_449 (
    .din     (_zz_4488[31:0]        ), //i
    .dout    (fixTo_449_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_450 (
    .din     (_zz_4489[31:0]        ), //i
    .dout    (fixTo_450_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_451 (
    .din     (_zz_4490[31:0]        ), //i
    .dout    (fixTo_451_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_452 (
    .din     (_zz_4491[31:0]        ), //i
    .dout    (fixTo_452_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_453 (
    .din     (_zz_4492[31:0]        ), //i
    .dout    (fixTo_453_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_454 (
    .din     (_zz_4493[31:0]        ), //i
    .dout    (fixTo_454_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_455 (
    .din     (_zz_4494[31:0]        ), //i
    .dout    (fixTo_455_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_456 (
    .din     (_zz_4495[31:0]        ), //i
    .dout    (fixTo_456_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_457 (
    .din     (_zz_4496[31:0]        ), //i
    .dout    (fixTo_457_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_458 (
    .din     (_zz_4497[31:0]        ), //i
    .dout    (fixTo_458_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_459 (
    .din     (_zz_4498[31:0]        ), //i
    .dout    (fixTo_459_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_460 (
    .din     (_zz_4499[31:0]        ), //i
    .dout    (fixTo_460_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_461 (
    .din     (_zz_4500[31:0]        ), //i
    .dout    (fixTo_461_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_462 (
    .din     (_zz_4501[31:0]        ), //i
    .dout    (fixTo_462_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_463 (
    .din     (_zz_4502[31:0]        ), //i
    .dout    (fixTo_463_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_464 (
    .din     (_zz_4503[31:0]        ), //i
    .dout    (fixTo_464_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_465 (
    .din     (_zz_4504[31:0]        ), //i
    .dout    (fixTo_465_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_466 (
    .din     (_zz_4505[31:0]        ), //i
    .dout    (fixTo_466_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_467 (
    .din     (_zz_4506[31:0]        ), //i
    .dout    (fixTo_467_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_468 (
    .din     (_zz_4507[31:0]        ), //i
    .dout    (fixTo_468_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_469 (
    .din     (_zz_4508[31:0]        ), //i
    .dout    (fixTo_469_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_470 (
    .din     (_zz_4509[31:0]        ), //i
    .dout    (fixTo_470_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_471 (
    .din     (_zz_4510[31:0]        ), //i
    .dout    (fixTo_471_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_472 (
    .din     (_zz_4511[31:0]        ), //i
    .dout    (fixTo_472_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_473 (
    .din     (_zz_4512[31:0]        ), //i
    .dout    (fixTo_473_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_474 (
    .din     (_zz_4513[31:0]        ), //i
    .dout    (fixTo_474_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_475 (
    .din     (_zz_4514[31:0]        ), //i
    .dout    (fixTo_475_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_476 (
    .din     (_zz_4515[31:0]        ), //i
    .dout    (fixTo_476_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_477 (
    .din     (_zz_4516[31:0]        ), //i
    .dout    (fixTo_477_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_478 (
    .din     (_zz_4517[31:0]        ), //i
    .dout    (fixTo_478_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_479 (
    .din     (_zz_4518[31:0]        ), //i
    .dout    (fixTo_479_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_480 (
    .din     (_zz_4519[31:0]        ), //i
    .dout    (fixTo_480_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_481 (
    .din     (_zz_4520[31:0]        ), //i
    .dout    (fixTo_481_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_482 (
    .din     (_zz_4521[31:0]        ), //i
    .dout    (fixTo_482_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_483 (
    .din     (_zz_4522[31:0]        ), //i
    .dout    (fixTo_483_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_484 (
    .din     (_zz_4523[31:0]        ), //i
    .dout    (fixTo_484_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_485 (
    .din     (_zz_4524[31:0]        ), //i
    .dout    (fixTo_485_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_486 (
    .din     (_zz_4525[31:0]        ), //i
    .dout    (fixTo_486_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_487 (
    .din     (_zz_4526[31:0]        ), //i
    .dout    (fixTo_487_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_488 (
    .din     (_zz_4527[31:0]        ), //i
    .dout    (fixTo_488_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_489 (
    .din     (_zz_4528[31:0]        ), //i
    .dout    (fixTo_489_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_490 (
    .din     (_zz_4529[31:0]        ), //i
    .dout    (fixTo_490_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_491 (
    .din     (_zz_4530[31:0]        ), //i
    .dout    (fixTo_491_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_492 (
    .din     (_zz_4531[31:0]        ), //i
    .dout    (fixTo_492_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_493 (
    .din     (_zz_4532[31:0]        ), //i
    .dout    (fixTo_493_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_494 (
    .din     (_zz_4533[31:0]        ), //i
    .dout    (fixTo_494_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_495 (
    .din     (_zz_4534[31:0]        ), //i
    .dout    (fixTo_495_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_496 (
    .din     (_zz_4535[31:0]        ), //i
    .dout    (fixTo_496_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_497 (
    .din     (_zz_4536[31:0]        ), //i
    .dout    (fixTo_497_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_498 (
    .din     (_zz_4537[31:0]        ), //i
    .dout    (fixTo_498_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_499 (
    .din     (_zz_4538[31:0]        ), //i
    .dout    (fixTo_499_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_500 (
    .din     (_zz_4539[31:0]        ), //i
    .dout    (fixTo_500_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_501 (
    .din     (_zz_4540[31:0]        ), //i
    .dout    (fixTo_501_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_502 (
    .din     (_zz_4541[31:0]        ), //i
    .dout    (fixTo_502_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_503 (
    .din     (_zz_4542[31:0]        ), //i
    .dout    (fixTo_503_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_504 (
    .din     (_zz_4543[31:0]        ), //i
    .dout    (fixTo_504_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_505 (
    .din     (_zz_4544[31:0]        ), //i
    .dout    (fixTo_505_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_506 (
    .din     (_zz_4545[31:0]        ), //i
    .dout    (fixTo_506_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_507 (
    .din     (_zz_4546[31:0]        ), //i
    .dout    (fixTo_507_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_508 (
    .din     (_zz_4547[31:0]        ), //i
    .dout    (fixTo_508_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_509 (
    .din     (_zz_4548[31:0]        ), //i
    .dout    (fixTo_509_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_510 (
    .din     (_zz_4549[31:0]        ), //i
    .dout    (fixTo_510_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_511 (
    .din     (_zz_4550[31:0]        ), //i
    .dout    (fixTo_511_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_512 (
    .din     (_zz_4551[31:0]        ), //i
    .dout    (fixTo_512_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_513 (
    .din     (_zz_4552[31:0]        ), //i
    .dout    (fixTo_513_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_514 (
    .din     (_zz_4553[31:0]        ), //i
    .dout    (fixTo_514_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_515 (
    .din     (_zz_4554[31:0]        ), //i
    .dout    (fixTo_515_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_516 (
    .din     (_zz_4555[31:0]        ), //i
    .dout    (fixTo_516_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_517 (
    .din     (_zz_4556[31:0]        ), //i
    .dout    (fixTo_517_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_518 (
    .din     (_zz_4557[31:0]        ), //i
    .dout    (fixTo_518_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_519 (
    .din     (_zz_4558[31:0]        ), //i
    .dout    (fixTo_519_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_520 (
    .din     (_zz_4559[31:0]        ), //i
    .dout    (fixTo_520_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_521 (
    .din     (_zz_4560[31:0]        ), //i
    .dout    (fixTo_521_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_522 (
    .din     (_zz_4561[31:0]        ), //i
    .dout    (fixTo_522_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_523 (
    .din     (_zz_4562[31:0]        ), //i
    .dout    (fixTo_523_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_524 (
    .din     (_zz_4563[31:0]        ), //i
    .dout    (fixTo_524_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_525 (
    .din     (_zz_4564[31:0]        ), //i
    .dout    (fixTo_525_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_526 (
    .din     (_zz_4565[31:0]        ), //i
    .dout    (fixTo_526_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_527 (
    .din     (_zz_4566[31:0]        ), //i
    .dout    (fixTo_527_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_528 (
    .din     (_zz_4567[31:0]        ), //i
    .dout    (fixTo_528_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_529 (
    .din     (_zz_4568[31:0]        ), //i
    .dout    (fixTo_529_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_530 (
    .din     (_zz_4569[31:0]        ), //i
    .dout    (fixTo_530_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_531 (
    .din     (_zz_4570[31:0]        ), //i
    .dout    (fixTo_531_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_532 (
    .din     (_zz_4571[31:0]        ), //i
    .dout    (fixTo_532_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_533 (
    .din     (_zz_4572[31:0]        ), //i
    .dout    (fixTo_533_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_534 (
    .din     (_zz_4573[31:0]        ), //i
    .dout    (fixTo_534_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_535 (
    .din     (_zz_4574[31:0]        ), //i
    .dout    (fixTo_535_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_536 (
    .din     (_zz_4575[31:0]        ), //i
    .dout    (fixTo_536_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_537 (
    .din     (_zz_4576[31:0]        ), //i
    .dout    (fixTo_537_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_538 (
    .din     (_zz_4577[31:0]        ), //i
    .dout    (fixTo_538_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_539 (
    .din     (_zz_4578[31:0]        ), //i
    .dout    (fixTo_539_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_540 (
    .din     (_zz_4579[31:0]        ), //i
    .dout    (fixTo_540_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_541 (
    .din     (_zz_4580[31:0]        ), //i
    .dout    (fixTo_541_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_542 (
    .din     (_zz_4581[31:0]        ), //i
    .dout    (fixTo_542_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_543 (
    .din     (_zz_4582[31:0]        ), //i
    .dout    (fixTo_543_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_544 (
    .din     (_zz_4583[31:0]        ), //i
    .dout    (fixTo_544_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_545 (
    .din     (_zz_4584[31:0]        ), //i
    .dout    (fixTo_545_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_546 (
    .din     (_zz_4585[31:0]        ), //i
    .dout    (fixTo_546_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_547 (
    .din     (_zz_4586[31:0]        ), //i
    .dout    (fixTo_547_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_548 (
    .din     (_zz_4587[31:0]        ), //i
    .dout    (fixTo_548_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_549 (
    .din     (_zz_4588[31:0]        ), //i
    .dout    (fixTo_549_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_550 (
    .din     (_zz_4589[31:0]        ), //i
    .dout    (fixTo_550_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_551 (
    .din     (_zz_4590[31:0]        ), //i
    .dout    (fixTo_551_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_552 (
    .din     (_zz_4591[31:0]        ), //i
    .dout    (fixTo_552_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_553 (
    .din     (_zz_4592[31:0]        ), //i
    .dout    (fixTo_553_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_554 (
    .din     (_zz_4593[31:0]        ), //i
    .dout    (fixTo_554_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_555 (
    .din     (_zz_4594[31:0]        ), //i
    .dout    (fixTo_555_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_556 (
    .din     (_zz_4595[31:0]        ), //i
    .dout    (fixTo_556_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_557 (
    .din     (_zz_4596[31:0]        ), //i
    .dout    (fixTo_557_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_558 (
    .din     (_zz_4597[31:0]        ), //i
    .dout    (fixTo_558_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_559 (
    .din     (_zz_4598[31:0]        ), //i
    .dout    (fixTo_559_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_560 (
    .din     (_zz_4599[31:0]        ), //i
    .dout    (fixTo_560_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_561 (
    .din     (_zz_4600[31:0]        ), //i
    .dout    (fixTo_561_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_562 (
    .din     (_zz_4601[31:0]        ), //i
    .dout    (fixTo_562_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_563 (
    .din     (_zz_4602[31:0]        ), //i
    .dout    (fixTo_563_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_564 (
    .din     (_zz_4603[31:0]        ), //i
    .dout    (fixTo_564_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_565 (
    .din     (_zz_4604[31:0]        ), //i
    .dout    (fixTo_565_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_566 (
    .din     (_zz_4605[31:0]        ), //i
    .dout    (fixTo_566_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_567 (
    .din     (_zz_4606[31:0]        ), //i
    .dout    (fixTo_567_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_568 (
    .din     (_zz_4607[31:0]        ), //i
    .dout    (fixTo_568_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_569 (
    .din     (_zz_4608[31:0]        ), //i
    .dout    (fixTo_569_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_570 (
    .din     (_zz_4609[31:0]        ), //i
    .dout    (fixTo_570_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_571 (
    .din     (_zz_4610[31:0]        ), //i
    .dout    (fixTo_571_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_572 (
    .din     (_zz_4611[31:0]        ), //i
    .dout    (fixTo_572_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_573 (
    .din     (_zz_4612[31:0]        ), //i
    .dout    (fixTo_573_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_574 (
    .din     (_zz_4613[31:0]        ), //i
    .dout    (fixTo_574_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_575 (
    .din     (_zz_4614[31:0]        ), //i
    .dout    (fixTo_575_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_576 (
    .din     (_zz_4615[31:0]        ), //i
    .dout    (fixTo_576_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_577 (
    .din     (_zz_4616[31:0]        ), //i
    .dout    (fixTo_577_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_578 (
    .din     (_zz_4617[31:0]        ), //i
    .dout    (fixTo_578_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_579 (
    .din     (_zz_4618[31:0]        ), //i
    .dout    (fixTo_579_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_580 (
    .din     (_zz_4619[31:0]        ), //i
    .dout    (fixTo_580_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_581 (
    .din     (_zz_4620[31:0]        ), //i
    .dout    (fixTo_581_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_582 (
    .din     (_zz_4621[31:0]        ), //i
    .dout    (fixTo_582_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_583 (
    .din     (_zz_4622[31:0]        ), //i
    .dout    (fixTo_583_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_584 (
    .din     (_zz_4623[31:0]        ), //i
    .dout    (fixTo_584_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_585 (
    .din     (_zz_4624[31:0]        ), //i
    .dout    (fixTo_585_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_586 (
    .din     (_zz_4625[31:0]        ), //i
    .dout    (fixTo_586_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_587 (
    .din     (_zz_4626[31:0]        ), //i
    .dout    (fixTo_587_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_588 (
    .din     (_zz_4627[31:0]        ), //i
    .dout    (fixTo_588_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_589 (
    .din     (_zz_4628[31:0]        ), //i
    .dout    (fixTo_589_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_590 (
    .din     (_zz_4629[31:0]        ), //i
    .dout    (fixTo_590_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_591 (
    .din     (_zz_4630[31:0]        ), //i
    .dout    (fixTo_591_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_592 (
    .din     (_zz_4631[31:0]        ), //i
    .dout    (fixTo_592_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_593 (
    .din     (_zz_4632[31:0]        ), //i
    .dout    (fixTo_593_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_594 (
    .din     (_zz_4633[31:0]        ), //i
    .dout    (fixTo_594_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_595 (
    .din     (_zz_4634[31:0]        ), //i
    .dout    (fixTo_595_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_596 (
    .din     (_zz_4635[31:0]        ), //i
    .dout    (fixTo_596_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_597 (
    .din     (_zz_4636[31:0]        ), //i
    .dout    (fixTo_597_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_598 (
    .din     (_zz_4637[31:0]        ), //i
    .dout    (fixTo_598_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_599 (
    .din     (_zz_4638[31:0]        ), //i
    .dout    (fixTo_599_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_600 (
    .din     (_zz_4639[31:0]        ), //i
    .dout    (fixTo_600_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_601 (
    .din     (_zz_4640[31:0]        ), //i
    .dout    (fixTo_601_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_602 (
    .din     (_zz_4641[31:0]        ), //i
    .dout    (fixTo_602_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_603 (
    .din     (_zz_4642[31:0]        ), //i
    .dout    (fixTo_603_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_604 (
    .din     (_zz_4643[31:0]        ), //i
    .dout    (fixTo_604_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_605 (
    .din     (_zz_4644[31:0]        ), //i
    .dout    (fixTo_605_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_606 (
    .din     (_zz_4645[31:0]        ), //i
    .dout    (fixTo_606_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_607 (
    .din     (_zz_4646[31:0]        ), //i
    .dout    (fixTo_607_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_608 (
    .din     (_zz_4647[31:0]        ), //i
    .dout    (fixTo_608_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_609 (
    .din     (_zz_4648[31:0]        ), //i
    .dout    (fixTo_609_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_610 (
    .din     (_zz_4649[31:0]        ), //i
    .dout    (fixTo_610_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_611 (
    .din     (_zz_4650[31:0]        ), //i
    .dout    (fixTo_611_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_612 (
    .din     (_zz_4651[31:0]        ), //i
    .dout    (fixTo_612_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_613 (
    .din     (_zz_4652[31:0]        ), //i
    .dout    (fixTo_613_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_614 (
    .din     (_zz_4653[31:0]        ), //i
    .dout    (fixTo_614_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_615 (
    .din     (_zz_4654[31:0]        ), //i
    .dout    (fixTo_615_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_616 (
    .din     (_zz_4655[31:0]        ), //i
    .dout    (fixTo_616_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_617 (
    .din     (_zz_4656[31:0]        ), //i
    .dout    (fixTo_617_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_618 (
    .din     (_zz_4657[31:0]        ), //i
    .dout    (fixTo_618_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_619 (
    .din     (_zz_4658[31:0]        ), //i
    .dout    (fixTo_619_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_620 (
    .din     (_zz_4659[31:0]        ), //i
    .dout    (fixTo_620_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_621 (
    .din     (_zz_4660[31:0]        ), //i
    .dout    (fixTo_621_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_622 (
    .din     (_zz_4661[31:0]        ), //i
    .dout    (fixTo_622_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_623 (
    .din     (_zz_4662[31:0]        ), //i
    .dout    (fixTo_623_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_624 (
    .din     (_zz_4663[31:0]        ), //i
    .dout    (fixTo_624_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_625 (
    .din     (_zz_4664[31:0]        ), //i
    .dout    (fixTo_625_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_626 (
    .din     (_zz_4665[31:0]        ), //i
    .dout    (fixTo_626_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_627 (
    .din     (_zz_4666[31:0]        ), //i
    .dout    (fixTo_627_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_628 (
    .din     (_zz_4667[31:0]        ), //i
    .dout    (fixTo_628_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_629 (
    .din     (_zz_4668[31:0]        ), //i
    .dout    (fixTo_629_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_630 (
    .din     (_zz_4669[31:0]        ), //i
    .dout    (fixTo_630_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_631 (
    .din     (_zz_4670[31:0]        ), //i
    .dout    (fixTo_631_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_632 (
    .din     (_zz_4671[31:0]        ), //i
    .dout    (fixTo_632_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_633 (
    .din     (_zz_4672[31:0]        ), //i
    .dout    (fixTo_633_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_634 (
    .din     (_zz_4673[31:0]        ), //i
    .dout    (fixTo_634_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_635 (
    .din     (_zz_4674[31:0]        ), //i
    .dout    (fixTo_635_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_636 (
    .din     (_zz_4675[31:0]        ), //i
    .dout    (fixTo_636_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_637 (
    .din     (_zz_4676[31:0]        ), //i
    .dout    (fixTo_637_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_638 (
    .din     (_zz_4677[31:0]        ), //i
    .dout    (fixTo_638_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_639 (
    .din     (_zz_4678[31:0]        ), //i
    .dout    (fixTo_639_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_640 (
    .din     (_zz_4679[31:0]        ), //i
    .dout    (fixTo_640_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_641 (
    .din     (_zz_4680[31:0]        ), //i
    .dout    (fixTo_641_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_642 (
    .din     (_zz_4681[31:0]        ), //i
    .dout    (fixTo_642_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_643 (
    .din     (_zz_4682[31:0]        ), //i
    .dout    (fixTo_643_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_644 (
    .din     (_zz_4683[31:0]        ), //i
    .dout    (fixTo_644_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_645 (
    .din     (_zz_4684[31:0]        ), //i
    .dout    (fixTo_645_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_646 (
    .din     (_zz_4685[31:0]        ), //i
    .dout    (fixTo_646_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_647 (
    .din     (_zz_4686[31:0]        ), //i
    .dout    (fixTo_647_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_648 (
    .din     (_zz_4687[31:0]        ), //i
    .dout    (fixTo_648_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_649 (
    .din     (_zz_4688[31:0]        ), //i
    .dout    (fixTo_649_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_650 (
    .din     (_zz_4689[31:0]        ), //i
    .dout    (fixTo_650_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_651 (
    .din     (_zz_4690[31:0]        ), //i
    .dout    (fixTo_651_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_652 (
    .din     (_zz_4691[31:0]        ), //i
    .dout    (fixTo_652_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_653 (
    .din     (_zz_4692[31:0]        ), //i
    .dout    (fixTo_653_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_654 (
    .din     (_zz_4693[31:0]        ), //i
    .dout    (fixTo_654_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_655 (
    .din     (_zz_4694[31:0]        ), //i
    .dout    (fixTo_655_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_656 (
    .din     (_zz_4695[31:0]        ), //i
    .dout    (fixTo_656_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_657 (
    .din     (_zz_4696[31:0]        ), //i
    .dout    (fixTo_657_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_658 (
    .din     (_zz_4697[31:0]        ), //i
    .dout    (fixTo_658_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_659 (
    .din     (_zz_4698[31:0]        ), //i
    .dout    (fixTo_659_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_660 (
    .din     (_zz_4699[31:0]        ), //i
    .dout    (fixTo_660_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_661 (
    .din     (_zz_4700[31:0]        ), //i
    .dout    (fixTo_661_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_662 (
    .din     (_zz_4701[31:0]        ), //i
    .dout    (fixTo_662_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_663 (
    .din     (_zz_4702[31:0]        ), //i
    .dout    (fixTo_663_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_664 (
    .din     (_zz_4703[31:0]        ), //i
    .dout    (fixTo_664_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_665 (
    .din     (_zz_4704[31:0]        ), //i
    .dout    (fixTo_665_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_666 (
    .din     (_zz_4705[31:0]        ), //i
    .dout    (fixTo_666_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_667 (
    .din     (_zz_4706[31:0]        ), //i
    .dout    (fixTo_667_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_668 (
    .din     (_zz_4707[31:0]        ), //i
    .dout    (fixTo_668_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_669 (
    .din     (_zz_4708[31:0]        ), //i
    .dout    (fixTo_669_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_670 (
    .din     (_zz_4709[31:0]        ), //i
    .dout    (fixTo_670_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_671 (
    .din     (_zz_4710[31:0]        ), //i
    .dout    (fixTo_671_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_672 (
    .din     (_zz_4711[31:0]        ), //i
    .dout    (fixTo_672_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_673 (
    .din     (_zz_4712[31:0]        ), //i
    .dout    (fixTo_673_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_674 (
    .din     (_zz_4713[31:0]        ), //i
    .dout    (fixTo_674_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_675 (
    .din     (_zz_4714[31:0]        ), //i
    .dout    (fixTo_675_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_676 (
    .din     (_zz_4715[31:0]        ), //i
    .dout    (fixTo_676_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_677 (
    .din     (_zz_4716[31:0]        ), //i
    .dout    (fixTo_677_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_678 (
    .din     (_zz_4717[31:0]        ), //i
    .dout    (fixTo_678_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_679 (
    .din     (_zz_4718[31:0]        ), //i
    .dout    (fixTo_679_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_680 (
    .din     (_zz_4719[31:0]        ), //i
    .dout    (fixTo_680_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_681 (
    .din     (_zz_4720[31:0]        ), //i
    .dout    (fixTo_681_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_682 (
    .din     (_zz_4721[31:0]        ), //i
    .dout    (fixTo_682_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_683 (
    .din     (_zz_4722[31:0]        ), //i
    .dout    (fixTo_683_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_684 (
    .din     (_zz_4723[31:0]        ), //i
    .dout    (fixTo_684_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_685 (
    .din     (_zz_4724[31:0]        ), //i
    .dout    (fixTo_685_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_686 (
    .din     (_zz_4725[31:0]        ), //i
    .dout    (fixTo_686_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_687 (
    .din     (_zz_4726[31:0]        ), //i
    .dout    (fixTo_687_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_688 (
    .din     (_zz_4727[31:0]        ), //i
    .dout    (fixTo_688_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_689 (
    .din     (_zz_4728[31:0]        ), //i
    .dout    (fixTo_689_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_690 (
    .din     (_zz_4729[31:0]        ), //i
    .dout    (fixTo_690_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_691 (
    .din     (_zz_4730[31:0]        ), //i
    .dout    (fixTo_691_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_692 (
    .din     (_zz_4731[31:0]        ), //i
    .dout    (fixTo_692_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_693 (
    .din     (_zz_4732[31:0]        ), //i
    .dout    (fixTo_693_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_694 (
    .din     (_zz_4733[31:0]        ), //i
    .dout    (fixTo_694_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_695 (
    .din     (_zz_4734[31:0]        ), //i
    .dout    (fixTo_695_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_696 (
    .din     (_zz_4735[31:0]        ), //i
    .dout    (fixTo_696_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_697 (
    .din     (_zz_4736[31:0]        ), //i
    .dout    (fixTo_697_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_698 (
    .din     (_zz_4737[31:0]        ), //i
    .dout    (fixTo_698_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_699 (
    .din     (_zz_4738[31:0]        ), //i
    .dout    (fixTo_699_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_700 (
    .din     (_zz_4739[31:0]        ), //i
    .dout    (fixTo_700_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_701 (
    .din     (_zz_4740[31:0]        ), //i
    .dout    (fixTo_701_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_702 (
    .din     (_zz_4741[31:0]        ), //i
    .dout    (fixTo_702_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_703 (
    .din     (_zz_4742[31:0]        ), //i
    .dout    (fixTo_703_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_704 (
    .din     (_zz_4743[31:0]        ), //i
    .dout    (fixTo_704_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_705 (
    .din     (_zz_4744[31:0]        ), //i
    .dout    (fixTo_705_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_706 (
    .din     (_zz_4745[31:0]        ), //i
    .dout    (fixTo_706_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_707 (
    .din     (_zz_4746[31:0]        ), //i
    .dout    (fixTo_707_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_708 (
    .din     (_zz_4747[31:0]        ), //i
    .dout    (fixTo_708_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_709 (
    .din     (_zz_4748[31:0]        ), //i
    .dout    (fixTo_709_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_710 (
    .din     (_zz_4749[31:0]        ), //i
    .dout    (fixTo_710_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_711 (
    .din     (_zz_4750[31:0]        ), //i
    .dout    (fixTo_711_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_712 (
    .din     (_zz_4751[31:0]        ), //i
    .dout    (fixTo_712_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_713 (
    .din     (_zz_4752[31:0]        ), //i
    .dout    (fixTo_713_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_714 (
    .din     (_zz_4753[31:0]        ), //i
    .dout    (fixTo_714_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_715 (
    .din     (_zz_4754[31:0]        ), //i
    .dout    (fixTo_715_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_716 (
    .din     (_zz_4755[31:0]        ), //i
    .dout    (fixTo_716_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_717 (
    .din     (_zz_4756[31:0]        ), //i
    .dout    (fixTo_717_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_718 (
    .din     (_zz_4757[31:0]        ), //i
    .dout    (fixTo_718_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_719 (
    .din     (_zz_4758[31:0]        ), //i
    .dout    (fixTo_719_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_720 (
    .din     (_zz_4759[31:0]        ), //i
    .dout    (fixTo_720_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_721 (
    .din     (_zz_4760[31:0]        ), //i
    .dout    (fixTo_721_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_722 (
    .din     (_zz_4761[31:0]        ), //i
    .dout    (fixTo_722_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_723 (
    .din     (_zz_4762[31:0]        ), //i
    .dout    (fixTo_723_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_724 (
    .din     (_zz_4763[31:0]        ), //i
    .dout    (fixTo_724_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_725 (
    .din     (_zz_4764[31:0]        ), //i
    .dout    (fixTo_725_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_726 (
    .din     (_zz_4765[31:0]        ), //i
    .dout    (fixTo_726_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_727 (
    .din     (_zz_4766[31:0]        ), //i
    .dout    (fixTo_727_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_728 (
    .din     (_zz_4767[31:0]        ), //i
    .dout    (fixTo_728_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_729 (
    .din     (_zz_4768[31:0]        ), //i
    .dout    (fixTo_729_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_730 (
    .din     (_zz_4769[31:0]        ), //i
    .dout    (fixTo_730_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_731 (
    .din     (_zz_4770[31:0]        ), //i
    .dout    (fixTo_731_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_732 (
    .din     (_zz_4771[31:0]        ), //i
    .dout    (fixTo_732_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_733 (
    .din     (_zz_4772[31:0]        ), //i
    .dout    (fixTo_733_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_734 (
    .din     (_zz_4773[31:0]        ), //i
    .dout    (fixTo_734_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_735 (
    .din     (_zz_4774[31:0]        ), //i
    .dout    (fixTo_735_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_736 (
    .din     (_zz_4775[31:0]        ), //i
    .dout    (fixTo_736_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_737 (
    .din     (_zz_4776[31:0]        ), //i
    .dout    (fixTo_737_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_738 (
    .din     (_zz_4777[31:0]        ), //i
    .dout    (fixTo_738_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_739 (
    .din     (_zz_4778[31:0]        ), //i
    .dout    (fixTo_739_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_740 (
    .din     (_zz_4779[31:0]        ), //i
    .dout    (fixTo_740_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_741 (
    .din     (_zz_4780[31:0]        ), //i
    .dout    (fixTo_741_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_742 (
    .din     (_zz_4781[31:0]        ), //i
    .dout    (fixTo_742_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_743 (
    .din     (_zz_4782[31:0]        ), //i
    .dout    (fixTo_743_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_744 (
    .din     (_zz_4783[31:0]        ), //i
    .dout    (fixTo_744_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_745 (
    .din     (_zz_4784[31:0]        ), //i
    .dout    (fixTo_745_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_746 (
    .din     (_zz_4785[31:0]        ), //i
    .dout    (fixTo_746_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_747 (
    .din     (_zz_4786[31:0]        ), //i
    .dout    (fixTo_747_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_748 (
    .din     (_zz_4787[31:0]        ), //i
    .dout    (fixTo_748_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_749 (
    .din     (_zz_4788[31:0]        ), //i
    .dout    (fixTo_749_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_750 (
    .din     (_zz_4789[31:0]        ), //i
    .dout    (fixTo_750_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_751 (
    .din     (_zz_4790[31:0]        ), //i
    .dout    (fixTo_751_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_752 (
    .din     (_zz_4791[31:0]        ), //i
    .dout    (fixTo_752_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_753 (
    .din     (_zz_4792[31:0]        ), //i
    .dout    (fixTo_753_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_754 (
    .din     (_zz_4793[31:0]        ), //i
    .dout    (fixTo_754_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_755 (
    .din     (_zz_4794[31:0]        ), //i
    .dout    (fixTo_755_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_756 (
    .din     (_zz_4795[31:0]        ), //i
    .dout    (fixTo_756_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_757 (
    .din     (_zz_4796[31:0]        ), //i
    .dout    (fixTo_757_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_758 (
    .din     (_zz_4797[31:0]        ), //i
    .dout    (fixTo_758_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_759 (
    .din     (_zz_4798[31:0]        ), //i
    .dout    (fixTo_759_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_760 (
    .din     (_zz_4799[31:0]        ), //i
    .dout    (fixTo_760_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_761 (
    .din     (_zz_4800[31:0]        ), //i
    .dout    (fixTo_761_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_762 (
    .din     (_zz_4801[31:0]        ), //i
    .dout    (fixTo_762_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_763 (
    .din     (_zz_4802[31:0]        ), //i
    .dout    (fixTo_763_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_764 (
    .din     (_zz_4803[31:0]        ), //i
    .dout    (fixTo_764_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_765 (
    .din     (_zz_4804[31:0]        ), //i
    .dout    (fixTo_765_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_766 (
    .din     (_zz_4805[31:0]        ), //i
    .dout    (fixTo_766_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_767 (
    .din     (_zz_4806[31:0]        ), //i
    .dout    (fixTo_767_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_768 (
    .din     (_zz_4807[31:0]        ), //i
    .dout    (fixTo_768_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_769 (
    .din     (_zz_4808[31:0]        ), //i
    .dout    (fixTo_769_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_770 (
    .din     (_zz_4809[31:0]        ), //i
    .dout    (fixTo_770_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_771 (
    .din     (_zz_4810[31:0]        ), //i
    .dout    (fixTo_771_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_772 (
    .din     (_zz_4811[31:0]        ), //i
    .dout    (fixTo_772_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_773 (
    .din     (_zz_4812[31:0]        ), //i
    .dout    (fixTo_773_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_774 (
    .din     (_zz_4813[31:0]        ), //i
    .dout    (fixTo_774_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_775 (
    .din     (_zz_4814[31:0]        ), //i
    .dout    (fixTo_775_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_776 (
    .din     (_zz_4815[31:0]        ), //i
    .dout    (fixTo_776_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_777 (
    .din     (_zz_4816[31:0]        ), //i
    .dout    (fixTo_777_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_778 (
    .din     (_zz_4817[31:0]        ), //i
    .dout    (fixTo_778_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_779 (
    .din     (_zz_4818[31:0]        ), //i
    .dout    (fixTo_779_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_780 (
    .din     (_zz_4819[31:0]        ), //i
    .dout    (fixTo_780_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_781 (
    .din     (_zz_4820[31:0]        ), //i
    .dout    (fixTo_781_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_782 (
    .din     (_zz_4821[31:0]        ), //i
    .dout    (fixTo_782_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_783 (
    .din     (_zz_4822[31:0]        ), //i
    .dout    (fixTo_783_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_784 (
    .din     (_zz_4823[31:0]        ), //i
    .dout    (fixTo_784_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_785 (
    .din     (_zz_4824[31:0]        ), //i
    .dout    (fixTo_785_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_786 (
    .din     (_zz_4825[31:0]        ), //i
    .dout    (fixTo_786_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_787 (
    .din     (_zz_4826[31:0]        ), //i
    .dout    (fixTo_787_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_788 (
    .din     (_zz_4827[31:0]        ), //i
    .dout    (fixTo_788_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_789 (
    .din     (_zz_4828[31:0]        ), //i
    .dout    (fixTo_789_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_790 (
    .din     (_zz_4829[31:0]        ), //i
    .dout    (fixTo_790_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_791 (
    .din     (_zz_4830[31:0]        ), //i
    .dout    (fixTo_791_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_792 (
    .din     (_zz_4831[31:0]        ), //i
    .dout    (fixTo_792_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_793 (
    .din     (_zz_4832[31:0]        ), //i
    .dout    (fixTo_793_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_794 (
    .din     (_zz_4833[31:0]        ), //i
    .dout    (fixTo_794_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_795 (
    .din     (_zz_4834[31:0]        ), //i
    .dout    (fixTo_795_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_796 (
    .din     (_zz_4835[31:0]        ), //i
    .dout    (fixTo_796_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_797 (
    .din     (_zz_4836[31:0]        ), //i
    .dout    (fixTo_797_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_798 (
    .din     (_zz_4837[31:0]        ), //i
    .dout    (fixTo_798_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_799 (
    .din     (_zz_4838[31:0]        ), //i
    .dout    (fixTo_799_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_800 (
    .din     (_zz_4839[31:0]        ), //i
    .dout    (fixTo_800_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_801 (
    .din     (_zz_4840[31:0]        ), //i
    .dout    (fixTo_801_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_802 (
    .din     (_zz_4841[31:0]        ), //i
    .dout    (fixTo_802_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_803 (
    .din     (_zz_4842[31:0]        ), //i
    .dout    (fixTo_803_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_804 (
    .din     (_zz_4843[31:0]        ), //i
    .dout    (fixTo_804_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_805 (
    .din     (_zz_4844[31:0]        ), //i
    .dout    (fixTo_805_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_806 (
    .din     (_zz_4845[31:0]        ), //i
    .dout    (fixTo_806_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_807 (
    .din     (_zz_4846[31:0]        ), //i
    .dout    (fixTo_807_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_808 (
    .din     (_zz_4847[31:0]        ), //i
    .dout    (fixTo_808_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_809 (
    .din     (_zz_4848[31:0]        ), //i
    .dout    (fixTo_809_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_810 (
    .din     (_zz_4849[31:0]        ), //i
    .dout    (fixTo_810_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_811 (
    .din     (_zz_4850[31:0]        ), //i
    .dout    (fixTo_811_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_812 (
    .din     (_zz_4851[31:0]        ), //i
    .dout    (fixTo_812_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_813 (
    .din     (_zz_4852[31:0]        ), //i
    .dout    (fixTo_813_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_814 (
    .din     (_zz_4853[31:0]        ), //i
    .dout    (fixTo_814_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_815 (
    .din     (_zz_4854[31:0]        ), //i
    .dout    (fixTo_815_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_816 (
    .din     (_zz_4855[31:0]        ), //i
    .dout    (fixTo_816_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_817 (
    .din     (_zz_4856[31:0]        ), //i
    .dout    (fixTo_817_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_818 (
    .din     (_zz_4857[31:0]        ), //i
    .dout    (fixTo_818_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_819 (
    .din     (_zz_4858[31:0]        ), //i
    .dout    (fixTo_819_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_820 (
    .din     (_zz_4859[31:0]        ), //i
    .dout    (fixTo_820_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_821 (
    .din     (_zz_4860[31:0]        ), //i
    .dout    (fixTo_821_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_822 (
    .din     (_zz_4861[31:0]        ), //i
    .dout    (fixTo_822_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_823 (
    .din     (_zz_4862[31:0]        ), //i
    .dout    (fixTo_823_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_824 (
    .din     (_zz_4863[31:0]        ), //i
    .dout    (fixTo_824_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_825 (
    .din     (_zz_4864[31:0]        ), //i
    .dout    (fixTo_825_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_826 (
    .din     (_zz_4865[31:0]        ), //i
    .dout    (fixTo_826_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_827 (
    .din     (_zz_4866[31:0]        ), //i
    .dout    (fixTo_827_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_828 (
    .din     (_zz_4867[31:0]        ), //i
    .dout    (fixTo_828_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_829 (
    .din     (_zz_4868[31:0]        ), //i
    .dout    (fixTo_829_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_830 (
    .din     (_zz_4869[31:0]        ), //i
    .dout    (fixTo_830_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_831 (
    .din     (_zz_4870[31:0]        ), //i
    .dout    (fixTo_831_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_832 (
    .din     (_zz_4871[31:0]        ), //i
    .dout    (fixTo_832_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_833 (
    .din     (_zz_4872[31:0]        ), //i
    .dout    (fixTo_833_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_834 (
    .din     (_zz_4873[31:0]        ), //i
    .dout    (fixTo_834_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_835 (
    .din     (_zz_4874[31:0]        ), //i
    .dout    (fixTo_835_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_836 (
    .din     (_zz_4875[31:0]        ), //i
    .dout    (fixTo_836_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_837 (
    .din     (_zz_4876[31:0]        ), //i
    .dout    (fixTo_837_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_838 (
    .din     (_zz_4877[31:0]        ), //i
    .dout    (fixTo_838_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_839 (
    .din     (_zz_4878[31:0]        ), //i
    .dout    (fixTo_839_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_840 (
    .din     (_zz_4879[31:0]        ), //i
    .dout    (fixTo_840_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_841 (
    .din     (_zz_4880[31:0]        ), //i
    .dout    (fixTo_841_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_842 (
    .din     (_zz_4881[31:0]        ), //i
    .dout    (fixTo_842_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_843 (
    .din     (_zz_4882[31:0]        ), //i
    .dout    (fixTo_843_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_844 (
    .din     (_zz_4883[31:0]        ), //i
    .dout    (fixTo_844_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_845 (
    .din     (_zz_4884[31:0]        ), //i
    .dout    (fixTo_845_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_846 (
    .din     (_zz_4885[31:0]        ), //i
    .dout    (fixTo_846_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_847 (
    .din     (_zz_4886[31:0]        ), //i
    .dout    (fixTo_847_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_848 (
    .din     (_zz_4887[31:0]        ), //i
    .dout    (fixTo_848_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_849 (
    .din     (_zz_4888[31:0]        ), //i
    .dout    (fixTo_849_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_850 (
    .din     (_zz_4889[31:0]        ), //i
    .dout    (fixTo_850_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_851 (
    .din     (_zz_4890[31:0]        ), //i
    .dout    (fixTo_851_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_852 (
    .din     (_zz_4891[31:0]        ), //i
    .dout    (fixTo_852_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_853 (
    .din     (_zz_4892[31:0]        ), //i
    .dout    (fixTo_853_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_854 (
    .din     (_zz_4893[31:0]        ), //i
    .dout    (fixTo_854_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_855 (
    .din     (_zz_4894[31:0]        ), //i
    .dout    (fixTo_855_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_856 (
    .din     (_zz_4895[31:0]        ), //i
    .dout    (fixTo_856_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_857 (
    .din     (_zz_4896[31:0]        ), //i
    .dout    (fixTo_857_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_858 (
    .din     (_zz_4897[31:0]        ), //i
    .dout    (fixTo_858_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_859 (
    .din     (_zz_4898[31:0]        ), //i
    .dout    (fixTo_859_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_860 (
    .din     (_zz_4899[31:0]        ), //i
    .dout    (fixTo_860_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_861 (
    .din     (_zz_4900[31:0]        ), //i
    .dout    (fixTo_861_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_862 (
    .din     (_zz_4901[31:0]        ), //i
    .dout    (fixTo_862_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_863 (
    .din     (_zz_4902[31:0]        ), //i
    .dout    (fixTo_863_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_864 (
    .din     (_zz_4903[31:0]        ), //i
    .dout    (fixTo_864_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_865 (
    .din     (_zz_4904[31:0]        ), //i
    .dout    (fixTo_865_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_866 (
    .din     (_zz_4905[31:0]        ), //i
    .dout    (fixTo_866_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_867 (
    .din     (_zz_4906[31:0]        ), //i
    .dout    (fixTo_867_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_868 (
    .din     (_zz_4907[31:0]        ), //i
    .dout    (fixTo_868_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_869 (
    .din     (_zz_4908[31:0]        ), //i
    .dout    (fixTo_869_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_870 (
    .din     (_zz_4909[31:0]        ), //i
    .dout    (fixTo_870_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_871 (
    .din     (_zz_4910[31:0]        ), //i
    .dout    (fixTo_871_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_872 (
    .din     (_zz_4911[31:0]        ), //i
    .dout    (fixTo_872_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_873 (
    .din     (_zz_4912[31:0]        ), //i
    .dout    (fixTo_873_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_874 (
    .din     (_zz_4913[31:0]        ), //i
    .dout    (fixTo_874_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_875 (
    .din     (_zz_4914[31:0]        ), //i
    .dout    (fixTo_875_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_876 (
    .din     (_zz_4915[31:0]        ), //i
    .dout    (fixTo_876_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_877 (
    .din     (_zz_4916[31:0]        ), //i
    .dout    (fixTo_877_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_878 (
    .din     (_zz_4917[31:0]        ), //i
    .dout    (fixTo_878_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_879 (
    .din     (_zz_4918[31:0]        ), //i
    .dout    (fixTo_879_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_880 (
    .din     (_zz_4919[31:0]        ), //i
    .dout    (fixTo_880_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_881 (
    .din     (_zz_4920[31:0]        ), //i
    .dout    (fixTo_881_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_882 (
    .din     (_zz_4921[31:0]        ), //i
    .dout    (fixTo_882_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_883 (
    .din     (_zz_4922[31:0]        ), //i
    .dout    (fixTo_883_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_884 (
    .din     (_zz_4923[31:0]        ), //i
    .dout    (fixTo_884_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_885 (
    .din     (_zz_4924[31:0]        ), //i
    .dout    (fixTo_885_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_886 (
    .din     (_zz_4925[31:0]        ), //i
    .dout    (fixTo_886_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_887 (
    .din     (_zz_4926[31:0]        ), //i
    .dout    (fixTo_887_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_888 (
    .din     (_zz_4927[31:0]        ), //i
    .dout    (fixTo_888_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_889 (
    .din     (_zz_4928[31:0]        ), //i
    .dout    (fixTo_889_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_890 (
    .din     (_zz_4929[31:0]        ), //i
    .dout    (fixTo_890_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_891 (
    .din     (_zz_4930[31:0]        ), //i
    .dout    (fixTo_891_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_892 (
    .din     (_zz_4931[31:0]        ), //i
    .dout    (fixTo_892_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_893 (
    .din     (_zz_4932[31:0]        ), //i
    .dout    (fixTo_893_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_894 (
    .din     (_zz_4933[31:0]        ), //i
    .dout    (fixTo_894_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_895 (
    .din     (_zz_4934[31:0]        ), //i
    .dout    (fixTo_895_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_896 (
    .din     (_zz_4935[31:0]        ), //i
    .dout    (fixTo_896_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_897 (
    .din     (_zz_4936[31:0]        ), //i
    .dout    (fixTo_897_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_898 (
    .din     (_zz_4937[31:0]        ), //i
    .dout    (fixTo_898_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_899 (
    .din     (_zz_4938[31:0]        ), //i
    .dout    (fixTo_899_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_900 (
    .din     (_zz_4939[31:0]        ), //i
    .dout    (fixTo_900_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_901 (
    .din     (_zz_4940[31:0]        ), //i
    .dout    (fixTo_901_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_902 (
    .din     (_zz_4941[31:0]        ), //i
    .dout    (fixTo_902_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_903 (
    .din     (_zz_4942[31:0]        ), //i
    .dout    (fixTo_903_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_904 (
    .din     (_zz_4943[31:0]        ), //i
    .dout    (fixTo_904_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_905 (
    .din     (_zz_4944[31:0]        ), //i
    .dout    (fixTo_905_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_906 (
    .din     (_zz_4945[31:0]        ), //i
    .dout    (fixTo_906_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_907 (
    .din     (_zz_4946[31:0]        ), //i
    .dout    (fixTo_907_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_908 (
    .din     (_zz_4947[31:0]        ), //i
    .dout    (fixTo_908_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_909 (
    .din     (_zz_4948[31:0]        ), //i
    .dout    (fixTo_909_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_910 (
    .din     (_zz_4949[31:0]        ), //i
    .dout    (fixTo_910_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_911 (
    .din     (_zz_4950[31:0]        ), //i
    .dout    (fixTo_911_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_912 (
    .din     (_zz_4951[31:0]        ), //i
    .dout    (fixTo_912_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_913 (
    .din     (_zz_4952[31:0]        ), //i
    .dout    (fixTo_913_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_914 (
    .din     (_zz_4953[31:0]        ), //i
    .dout    (fixTo_914_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_915 (
    .din     (_zz_4954[31:0]        ), //i
    .dout    (fixTo_915_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_916 (
    .din     (_zz_4955[31:0]        ), //i
    .dout    (fixTo_916_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_917 (
    .din     (_zz_4956[31:0]        ), //i
    .dout    (fixTo_917_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_918 (
    .din     (_zz_4957[31:0]        ), //i
    .dout    (fixTo_918_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_919 (
    .din     (_zz_4958[31:0]        ), //i
    .dout    (fixTo_919_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_920 (
    .din     (_zz_4959[31:0]        ), //i
    .dout    (fixTo_920_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_921 (
    .din     (_zz_4960[31:0]        ), //i
    .dout    (fixTo_921_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_922 (
    .din     (_zz_4961[31:0]        ), //i
    .dout    (fixTo_922_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_923 (
    .din     (_zz_4962[31:0]        ), //i
    .dout    (fixTo_923_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_924 (
    .din     (_zz_4963[31:0]        ), //i
    .dout    (fixTo_924_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_925 (
    .din     (_zz_4964[31:0]        ), //i
    .dout    (fixTo_925_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_926 (
    .din     (_zz_4965[31:0]        ), //i
    .dout    (fixTo_926_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_927 (
    .din     (_zz_4966[31:0]        ), //i
    .dout    (fixTo_927_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_928 (
    .din     (_zz_4967[31:0]        ), //i
    .dout    (fixTo_928_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_929 (
    .din     (_zz_4968[31:0]        ), //i
    .dout    (fixTo_929_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_930 (
    .din     (_zz_4969[31:0]        ), //i
    .dout    (fixTo_930_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_931 (
    .din     (_zz_4970[31:0]        ), //i
    .dout    (fixTo_931_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_932 (
    .din     (_zz_4971[31:0]        ), //i
    .dout    (fixTo_932_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_933 (
    .din     (_zz_4972[31:0]        ), //i
    .dout    (fixTo_933_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_934 (
    .din     (_zz_4973[31:0]        ), //i
    .dout    (fixTo_934_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_935 (
    .din     (_zz_4974[31:0]        ), //i
    .dout    (fixTo_935_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_936 (
    .din     (_zz_4975[31:0]        ), //i
    .dout    (fixTo_936_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_937 (
    .din     (_zz_4976[31:0]        ), //i
    .dout    (fixTo_937_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_938 (
    .din     (_zz_4977[31:0]        ), //i
    .dout    (fixTo_938_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_939 (
    .din     (_zz_4978[31:0]        ), //i
    .dout    (fixTo_939_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_940 (
    .din     (_zz_4979[31:0]        ), //i
    .dout    (fixTo_940_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_941 (
    .din     (_zz_4980[31:0]        ), //i
    .dout    (fixTo_941_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_942 (
    .din     (_zz_4981[31:0]        ), //i
    .dout    (fixTo_942_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_943 (
    .din     (_zz_4982[31:0]        ), //i
    .dout    (fixTo_943_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_944 (
    .din     (_zz_4983[31:0]        ), //i
    .dout    (fixTo_944_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_945 (
    .din     (_zz_4984[31:0]        ), //i
    .dout    (fixTo_945_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_946 (
    .din     (_zz_4985[31:0]        ), //i
    .dout    (fixTo_946_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_947 (
    .din     (_zz_4986[31:0]        ), //i
    .dout    (fixTo_947_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_948 (
    .din     (_zz_4987[31:0]        ), //i
    .dout    (fixTo_948_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_949 (
    .din     (_zz_4988[31:0]        ), //i
    .dout    (fixTo_949_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_950 (
    .din     (_zz_4989[31:0]        ), //i
    .dout    (fixTo_950_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_951 (
    .din     (_zz_4990[31:0]        ), //i
    .dout    (fixTo_951_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_952 (
    .din     (_zz_4991[31:0]        ), //i
    .dout    (fixTo_952_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_953 (
    .din     (_zz_4992[31:0]        ), //i
    .dout    (fixTo_953_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_954 (
    .din     (_zz_4993[31:0]        ), //i
    .dout    (fixTo_954_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_955 (
    .din     (_zz_4994[31:0]        ), //i
    .dout    (fixTo_955_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_956 (
    .din     (_zz_4995[31:0]        ), //i
    .dout    (fixTo_956_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_957 (
    .din     (_zz_4996[31:0]        ), //i
    .dout    (fixTo_957_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_958 (
    .din     (_zz_4997[31:0]        ), //i
    .dout    (fixTo_958_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_959 (
    .din     (_zz_4998[31:0]        ), //i
    .dout    (fixTo_959_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_960 (
    .din     (_zz_4999[31:0]        ), //i
    .dout    (fixTo_960_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_961 (
    .din     (_zz_5000[31:0]        ), //i
    .dout    (fixTo_961_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_962 (
    .din     (_zz_5001[31:0]        ), //i
    .dout    (fixTo_962_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_963 (
    .din     (_zz_5002[31:0]        ), //i
    .dout    (fixTo_963_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_964 (
    .din     (_zz_5003[31:0]        ), //i
    .dout    (fixTo_964_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_965 (
    .din     (_zz_5004[31:0]        ), //i
    .dout    (fixTo_965_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_966 (
    .din     (_zz_5005[31:0]        ), //i
    .dout    (fixTo_966_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_967 (
    .din     (_zz_5006[31:0]        ), //i
    .dout    (fixTo_967_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_968 (
    .din     (_zz_5007[31:0]        ), //i
    .dout    (fixTo_968_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_969 (
    .din     (_zz_5008[31:0]        ), //i
    .dout    (fixTo_969_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_970 (
    .din     (_zz_5009[31:0]        ), //i
    .dout    (fixTo_970_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_971 (
    .din     (_zz_5010[31:0]        ), //i
    .dout    (fixTo_971_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_972 (
    .din     (_zz_5011[31:0]        ), //i
    .dout    (fixTo_972_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_973 (
    .din     (_zz_5012[31:0]        ), //i
    .dout    (fixTo_973_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_974 (
    .din     (_zz_5013[31:0]        ), //i
    .dout    (fixTo_974_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_975 (
    .din     (_zz_5014[31:0]        ), //i
    .dout    (fixTo_975_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_976 (
    .din     (_zz_5015[31:0]        ), //i
    .dout    (fixTo_976_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_977 (
    .din     (_zz_5016[31:0]        ), //i
    .dout    (fixTo_977_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_978 (
    .din     (_zz_5017[31:0]        ), //i
    .dout    (fixTo_978_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_979 (
    .din     (_zz_5018[31:0]        ), //i
    .dout    (fixTo_979_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_980 (
    .din     (_zz_5019[31:0]        ), //i
    .dout    (fixTo_980_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_981 (
    .din     (_zz_5020[31:0]        ), //i
    .dout    (fixTo_981_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_982 (
    .din     (_zz_5021[31:0]        ), //i
    .dout    (fixTo_982_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_983 (
    .din     (_zz_5022[31:0]        ), //i
    .dout    (fixTo_983_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_984 (
    .din     (_zz_5023[31:0]        ), //i
    .dout    (fixTo_984_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_985 (
    .din     (_zz_5024[31:0]        ), //i
    .dout    (fixTo_985_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_986 (
    .din     (_zz_5025[31:0]        ), //i
    .dout    (fixTo_986_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_987 (
    .din     (_zz_5026[31:0]        ), //i
    .dout    (fixTo_987_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_988 (
    .din     (_zz_5027[31:0]        ), //i
    .dout    (fixTo_988_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_989 (
    .din     (_zz_5028[31:0]        ), //i
    .dout    (fixTo_989_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_990 (
    .din     (_zz_5029[31:0]        ), //i
    .dout    (fixTo_990_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_991 (
    .din     (_zz_5030[31:0]        ), //i
    .dout    (fixTo_991_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_992 (
    .din     (_zz_5031[31:0]        ), //i
    .dout    (fixTo_992_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_993 (
    .din     (_zz_5032[31:0]        ), //i
    .dout    (fixTo_993_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_994 (
    .din     (_zz_5033[31:0]        ), //i
    .dout    (fixTo_994_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_995 (
    .din     (_zz_5034[31:0]        ), //i
    .dout    (fixTo_995_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_996 (
    .din     (_zz_5035[31:0]        ), //i
    .dout    (fixTo_996_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_997 (
    .din     (_zz_5036[31:0]        ), //i
    .dout    (fixTo_997_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_998 (
    .din     (_zz_5037[31:0]        ), //i
    .dout    (fixTo_998_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_999 (
    .din     (_zz_5038[31:0]        ), //i
    .dout    (fixTo_999_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1000 (
    .din     (_zz_5039[31:0]         ), //i
    .dout    (fixTo_1000_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1001 (
    .din     (_zz_5040[31:0]         ), //i
    .dout    (fixTo_1001_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1002 (
    .din     (_zz_5041[31:0]         ), //i
    .dout    (fixTo_1002_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1003 (
    .din     (_zz_5042[31:0]         ), //i
    .dout    (fixTo_1003_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1004 (
    .din     (_zz_5043[31:0]         ), //i
    .dout    (fixTo_1004_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1005 (
    .din     (_zz_5044[31:0]         ), //i
    .dout    (fixTo_1005_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1006 (
    .din     (_zz_5045[31:0]         ), //i
    .dout    (fixTo_1006_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1007 (
    .din     (_zz_5046[31:0]         ), //i
    .dout    (fixTo_1007_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1008 (
    .din     (_zz_5047[31:0]         ), //i
    .dout    (fixTo_1008_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1009 (
    .din     (_zz_5048[31:0]         ), //i
    .dout    (fixTo_1009_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1010 (
    .din     (_zz_5049[31:0]         ), //i
    .dout    (fixTo_1010_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1011 (
    .din     (_zz_5050[31:0]         ), //i
    .dout    (fixTo_1011_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1012 (
    .din     (_zz_5051[31:0]         ), //i
    .dout    (fixTo_1012_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1013 (
    .din     (_zz_5052[31:0]         ), //i
    .dout    (fixTo_1013_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1014 (
    .din     (_zz_5053[31:0]         ), //i
    .dout    (fixTo_1014_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1015 (
    .din     (_zz_5054[31:0]         ), //i
    .dout    (fixTo_1015_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1016 (
    .din     (_zz_5055[31:0]         ), //i
    .dout    (fixTo_1016_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1017 (
    .din     (_zz_5056[31:0]         ), //i
    .dout    (fixTo_1017_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1018 (
    .din     (_zz_5057[31:0]         ), //i
    .dout    (fixTo_1018_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1019 (
    .din     (_zz_5058[31:0]         ), //i
    .dout    (fixTo_1019_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1020 (
    .din     (_zz_5059[31:0]         ), //i
    .dout    (fixTo_1020_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1021 (
    .din     (_zz_5060[31:0]         ), //i
    .dout    (fixTo_1021_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1022 (
    .din     (_zz_5061[31:0]         ), //i
    .dout    (fixTo_1022_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1023 (
    .din     (_zz_5062[31:0]         ), //i
    .dout    (fixTo_1023_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1024 (
    .din     (_zz_5063[31:0]         ), //i
    .dout    (fixTo_1024_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1025 (
    .din     (_zz_5064[31:0]         ), //i
    .dout    (fixTo_1025_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1026 (
    .din     (_zz_5065[31:0]         ), //i
    .dout    (fixTo_1026_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1027 (
    .din     (_zz_5066[31:0]         ), //i
    .dout    (fixTo_1027_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1028 (
    .din     (_zz_5067[31:0]         ), //i
    .dout    (fixTo_1028_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1029 (
    .din     (_zz_5068[31:0]         ), //i
    .dout    (fixTo_1029_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1030 (
    .din     (_zz_5069[31:0]         ), //i
    .dout    (fixTo_1030_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1031 (
    .din     (_zz_5070[31:0]         ), //i
    .dout    (fixTo_1031_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1032 (
    .din     (_zz_5071[31:0]         ), //i
    .dout    (fixTo_1032_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1033 (
    .din     (_zz_5072[31:0]         ), //i
    .dout    (fixTo_1033_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1034 (
    .din     (_zz_5073[31:0]         ), //i
    .dout    (fixTo_1034_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1035 (
    .din     (_zz_5074[31:0]         ), //i
    .dout    (fixTo_1035_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1036 (
    .din     (_zz_5075[31:0]         ), //i
    .dout    (fixTo_1036_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1037 (
    .din     (_zz_5076[31:0]         ), //i
    .dout    (fixTo_1037_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1038 (
    .din     (_zz_5077[31:0]         ), //i
    .dout    (fixTo_1038_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1039 (
    .din     (_zz_5078[31:0]         ), //i
    .dout    (fixTo_1039_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1040 (
    .din     (_zz_5079[31:0]         ), //i
    .dout    (fixTo_1040_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1041 (
    .din     (_zz_5080[31:0]         ), //i
    .dout    (fixTo_1041_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1042 (
    .din     (_zz_5081[31:0]         ), //i
    .dout    (fixTo_1042_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1043 (
    .din     (_zz_5082[31:0]         ), //i
    .dout    (fixTo_1043_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1044 (
    .din     (_zz_5083[31:0]         ), //i
    .dout    (fixTo_1044_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1045 (
    .din     (_zz_5084[31:0]         ), //i
    .dout    (fixTo_1045_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1046 (
    .din     (_zz_5085[31:0]         ), //i
    .dout    (fixTo_1046_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1047 (
    .din     (_zz_5086[31:0]         ), //i
    .dout    (fixTo_1047_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1048 (
    .din     (_zz_5087[31:0]         ), //i
    .dout    (fixTo_1048_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1049 (
    .din     (_zz_5088[31:0]         ), //i
    .dout    (fixTo_1049_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1050 (
    .din     (_zz_5089[31:0]         ), //i
    .dout    (fixTo_1050_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1051 (
    .din     (_zz_5090[31:0]         ), //i
    .dout    (fixTo_1051_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1052 (
    .din     (_zz_5091[31:0]         ), //i
    .dout    (fixTo_1052_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1053 (
    .din     (_zz_5092[31:0]         ), //i
    .dout    (fixTo_1053_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1054 (
    .din     (_zz_5093[31:0]         ), //i
    .dout    (fixTo_1054_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1055 (
    .din     (_zz_5094[31:0]         ), //i
    .dout    (fixTo_1055_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1056 (
    .din     (_zz_5095[31:0]         ), //i
    .dout    (fixTo_1056_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1057 (
    .din     (_zz_5096[31:0]         ), //i
    .dout    (fixTo_1057_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1058 (
    .din     (_zz_5097[31:0]         ), //i
    .dout    (fixTo_1058_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1059 (
    .din     (_zz_5098[31:0]         ), //i
    .dout    (fixTo_1059_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1060 (
    .din     (_zz_5099[31:0]         ), //i
    .dout    (fixTo_1060_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1061 (
    .din     (_zz_5100[31:0]         ), //i
    .dout    (fixTo_1061_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1062 (
    .din     (_zz_5101[31:0]         ), //i
    .dout    (fixTo_1062_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1063 (
    .din     (_zz_5102[31:0]         ), //i
    .dout    (fixTo_1063_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1064 (
    .din     (_zz_5103[31:0]         ), //i
    .dout    (fixTo_1064_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1065 (
    .din     (_zz_5104[31:0]         ), //i
    .dout    (fixTo_1065_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1066 (
    .din     (_zz_5105[31:0]         ), //i
    .dout    (fixTo_1066_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1067 (
    .din     (_zz_5106[31:0]         ), //i
    .dout    (fixTo_1067_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1068 (
    .din     (_zz_5107[31:0]         ), //i
    .dout    (fixTo_1068_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1069 (
    .din     (_zz_5108[31:0]         ), //i
    .dout    (fixTo_1069_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1070 (
    .din     (_zz_5109[31:0]         ), //i
    .dout    (fixTo_1070_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1071 (
    .din     (_zz_5110[31:0]         ), //i
    .dout    (fixTo_1071_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1072 (
    .din     (_zz_5111[31:0]         ), //i
    .dout    (fixTo_1072_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1073 (
    .din     (_zz_5112[31:0]         ), //i
    .dout    (fixTo_1073_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1074 (
    .din     (_zz_5113[31:0]         ), //i
    .dout    (fixTo_1074_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1075 (
    .din     (_zz_5114[31:0]         ), //i
    .dout    (fixTo_1075_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1076 (
    .din     (_zz_5115[31:0]         ), //i
    .dout    (fixTo_1076_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1077 (
    .din     (_zz_5116[31:0]         ), //i
    .dout    (fixTo_1077_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1078 (
    .din     (_zz_5117[31:0]         ), //i
    .dout    (fixTo_1078_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1079 (
    .din     (_zz_5118[31:0]         ), //i
    .dout    (fixTo_1079_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1080 (
    .din     (_zz_5119[31:0]         ), //i
    .dout    (fixTo_1080_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1081 (
    .din     (_zz_5120[31:0]         ), //i
    .dout    (fixTo_1081_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1082 (
    .din     (_zz_5121[31:0]         ), //i
    .dout    (fixTo_1082_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1083 (
    .din     (_zz_5122[31:0]         ), //i
    .dout    (fixTo_1083_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1084 (
    .din     (_zz_5123[31:0]         ), //i
    .dout    (fixTo_1084_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1085 (
    .din     (_zz_5124[31:0]         ), //i
    .dout    (fixTo_1085_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1086 (
    .din     (_zz_5125[31:0]         ), //i
    .dout    (fixTo_1086_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1087 (
    .din     (_zz_5126[31:0]         ), //i
    .dout    (fixTo_1087_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1088 (
    .din     (_zz_5127[31:0]         ), //i
    .dout    (fixTo_1088_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1089 (
    .din     (_zz_5128[31:0]         ), //i
    .dout    (fixTo_1089_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1090 (
    .din     (_zz_5129[31:0]         ), //i
    .dout    (fixTo_1090_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1091 (
    .din     (_zz_5130[31:0]         ), //i
    .dout    (fixTo_1091_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1092 (
    .din     (_zz_5131[31:0]         ), //i
    .dout    (fixTo_1092_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1093 (
    .din     (_zz_5132[31:0]         ), //i
    .dout    (fixTo_1093_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1094 (
    .din     (_zz_5133[31:0]         ), //i
    .dout    (fixTo_1094_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1095 (
    .din     (_zz_5134[31:0]         ), //i
    .dout    (fixTo_1095_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1096 (
    .din     (_zz_5135[31:0]         ), //i
    .dout    (fixTo_1096_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1097 (
    .din     (_zz_5136[31:0]         ), //i
    .dout    (fixTo_1097_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1098 (
    .din     (_zz_5137[31:0]         ), //i
    .dout    (fixTo_1098_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1099 (
    .din     (_zz_5138[31:0]         ), //i
    .dout    (fixTo_1099_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1100 (
    .din     (_zz_5139[31:0]         ), //i
    .dout    (fixTo_1100_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1101 (
    .din     (_zz_5140[31:0]         ), //i
    .dout    (fixTo_1101_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1102 (
    .din     (_zz_5141[31:0]         ), //i
    .dout    (fixTo_1102_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1103 (
    .din     (_zz_5142[31:0]         ), //i
    .dout    (fixTo_1103_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1104 (
    .din     (_zz_5143[31:0]         ), //i
    .dout    (fixTo_1104_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1105 (
    .din     (_zz_5144[31:0]         ), //i
    .dout    (fixTo_1105_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1106 (
    .din     (_zz_5145[31:0]         ), //i
    .dout    (fixTo_1106_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1107 (
    .din     (_zz_5146[31:0]         ), //i
    .dout    (fixTo_1107_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1108 (
    .din     (_zz_5147[31:0]         ), //i
    .dout    (fixTo_1108_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1109 (
    .din     (_zz_5148[31:0]         ), //i
    .dout    (fixTo_1109_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1110 (
    .din     (_zz_5149[31:0]         ), //i
    .dout    (fixTo_1110_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1111 (
    .din     (_zz_5150[31:0]         ), //i
    .dout    (fixTo_1111_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1112 (
    .din     (_zz_5151[31:0]         ), //i
    .dout    (fixTo_1112_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1113 (
    .din     (_zz_5152[31:0]         ), //i
    .dout    (fixTo_1113_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1114 (
    .din     (_zz_5153[31:0]         ), //i
    .dout    (fixTo_1114_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1115 (
    .din     (_zz_5154[31:0]         ), //i
    .dout    (fixTo_1115_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1116 (
    .din     (_zz_5155[31:0]         ), //i
    .dout    (fixTo_1116_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1117 (
    .din     (_zz_5156[31:0]         ), //i
    .dout    (fixTo_1117_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1118 (
    .din     (_zz_5157[31:0]         ), //i
    .dout    (fixTo_1118_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1119 (
    .din     (_zz_5158[31:0]         ), //i
    .dout    (fixTo_1119_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1120 (
    .din     (_zz_5159[31:0]         ), //i
    .dout    (fixTo_1120_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1121 (
    .din     (_zz_5160[31:0]         ), //i
    .dout    (fixTo_1121_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1122 (
    .din     (_zz_5161[31:0]         ), //i
    .dout    (fixTo_1122_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1123 (
    .din     (_zz_5162[31:0]         ), //i
    .dout    (fixTo_1123_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1124 (
    .din     (_zz_5163[31:0]         ), //i
    .dout    (fixTo_1124_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1125 (
    .din     (_zz_5164[31:0]         ), //i
    .dout    (fixTo_1125_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1126 (
    .din     (_zz_5165[31:0]         ), //i
    .dout    (fixTo_1126_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1127 (
    .din     (_zz_5166[31:0]         ), //i
    .dout    (fixTo_1127_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1128 (
    .din     (_zz_5167[31:0]         ), //i
    .dout    (fixTo_1128_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1129 (
    .din     (_zz_5168[31:0]         ), //i
    .dout    (fixTo_1129_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1130 (
    .din     (_zz_5169[31:0]         ), //i
    .dout    (fixTo_1130_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1131 (
    .din     (_zz_5170[31:0]         ), //i
    .dout    (fixTo_1131_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1132 (
    .din     (_zz_5171[31:0]         ), //i
    .dout    (fixTo_1132_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1133 (
    .din     (_zz_5172[31:0]         ), //i
    .dout    (fixTo_1133_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1134 (
    .din     (_zz_5173[31:0]         ), //i
    .dout    (fixTo_1134_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1135 (
    .din     (_zz_5174[31:0]         ), //i
    .dout    (fixTo_1135_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1136 (
    .din     (_zz_5175[31:0]         ), //i
    .dout    (fixTo_1136_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1137 (
    .din     (_zz_5176[31:0]         ), //i
    .dout    (fixTo_1137_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1138 (
    .din     (_zz_5177[31:0]         ), //i
    .dout    (fixTo_1138_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1139 (
    .din     (_zz_5178[31:0]         ), //i
    .dout    (fixTo_1139_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1140 (
    .din     (_zz_5179[31:0]         ), //i
    .dout    (fixTo_1140_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1141 (
    .din     (_zz_5180[31:0]         ), //i
    .dout    (fixTo_1141_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1142 (
    .din     (_zz_5181[31:0]         ), //i
    .dout    (fixTo_1142_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1143 (
    .din     (_zz_5182[31:0]         ), //i
    .dout    (fixTo_1143_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1144 (
    .din     (_zz_5183[31:0]         ), //i
    .dout    (fixTo_1144_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1145 (
    .din     (_zz_5184[31:0]         ), //i
    .dout    (fixTo_1145_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1146 (
    .din     (_zz_5185[31:0]         ), //i
    .dout    (fixTo_1146_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1147 (
    .din     (_zz_5186[31:0]         ), //i
    .dout    (fixTo_1147_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1148 (
    .din     (_zz_5187[31:0]         ), //i
    .dout    (fixTo_1148_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1149 (
    .din     (_zz_5188[31:0]         ), //i
    .dout    (fixTo_1149_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1150 (
    .din     (_zz_5189[31:0]         ), //i
    .dout    (fixTo_1150_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1151 (
    .din     (_zz_5190[31:0]         ), //i
    .dout    (fixTo_1151_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1152 (
    .din     (_zz_5191[31:0]         ), //i
    .dout    (fixTo_1152_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1153 (
    .din     (_zz_5192[31:0]         ), //i
    .dout    (fixTo_1153_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1154 (
    .din     (_zz_5193[31:0]         ), //i
    .dout    (fixTo_1154_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1155 (
    .din     (_zz_5194[31:0]         ), //i
    .dout    (fixTo_1155_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1156 (
    .din     (_zz_5195[31:0]         ), //i
    .dout    (fixTo_1156_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1157 (
    .din     (_zz_5196[31:0]         ), //i
    .dout    (fixTo_1157_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1158 (
    .din     (_zz_5197[31:0]         ), //i
    .dout    (fixTo_1158_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1159 (
    .din     (_zz_5198[31:0]         ), //i
    .dout    (fixTo_1159_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1160 (
    .din     (_zz_5199[31:0]         ), //i
    .dout    (fixTo_1160_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1161 (
    .din     (_zz_5200[31:0]         ), //i
    .dout    (fixTo_1161_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1162 (
    .din     (_zz_5201[31:0]         ), //i
    .dout    (fixTo_1162_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1163 (
    .din     (_zz_5202[31:0]         ), //i
    .dout    (fixTo_1163_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1164 (
    .din     (_zz_5203[31:0]         ), //i
    .dout    (fixTo_1164_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1165 (
    .din     (_zz_5204[31:0]         ), //i
    .dout    (fixTo_1165_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1166 (
    .din     (_zz_5205[31:0]         ), //i
    .dout    (fixTo_1166_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1167 (
    .din     (_zz_5206[31:0]         ), //i
    .dout    (fixTo_1167_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1168 (
    .din     (_zz_5207[31:0]         ), //i
    .dout    (fixTo_1168_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1169 (
    .din     (_zz_5208[31:0]         ), //i
    .dout    (fixTo_1169_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1170 (
    .din     (_zz_5209[31:0]         ), //i
    .dout    (fixTo_1170_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1171 (
    .din     (_zz_5210[31:0]         ), //i
    .dout    (fixTo_1171_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1172 (
    .din     (_zz_5211[31:0]         ), //i
    .dout    (fixTo_1172_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1173 (
    .din     (_zz_5212[31:0]         ), //i
    .dout    (fixTo_1173_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1174 (
    .din     (_zz_5213[31:0]         ), //i
    .dout    (fixTo_1174_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1175 (
    .din     (_zz_5214[31:0]         ), //i
    .dout    (fixTo_1175_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1176 (
    .din     (_zz_5215[31:0]         ), //i
    .dout    (fixTo_1176_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1177 (
    .din     (_zz_5216[31:0]         ), //i
    .dout    (fixTo_1177_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1178 (
    .din     (_zz_5217[31:0]         ), //i
    .dout    (fixTo_1178_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1179 (
    .din     (_zz_5218[31:0]         ), //i
    .dout    (fixTo_1179_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1180 (
    .din     (_zz_5219[31:0]         ), //i
    .dout    (fixTo_1180_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1181 (
    .din     (_zz_5220[31:0]         ), //i
    .dout    (fixTo_1181_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1182 (
    .din     (_zz_5221[31:0]         ), //i
    .dout    (fixTo_1182_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1183 (
    .din     (_zz_5222[31:0]         ), //i
    .dout    (fixTo_1183_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1184 (
    .din     (_zz_5223[31:0]         ), //i
    .dout    (fixTo_1184_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1185 (
    .din     (_zz_5224[31:0]         ), //i
    .dout    (fixTo_1185_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1186 (
    .din     (_zz_5225[31:0]         ), //i
    .dout    (fixTo_1186_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1187 (
    .din     (_zz_5226[31:0]         ), //i
    .dout    (fixTo_1187_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1188 (
    .din     (_zz_5227[31:0]         ), //i
    .dout    (fixTo_1188_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1189 (
    .din     (_zz_5228[31:0]         ), //i
    .dout    (fixTo_1189_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1190 (
    .din     (_zz_5229[31:0]         ), //i
    .dout    (fixTo_1190_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1191 (
    .din     (_zz_5230[31:0]         ), //i
    .dout    (fixTo_1191_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1192 (
    .din     (_zz_5231[31:0]         ), //i
    .dout    (fixTo_1192_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1193 (
    .din     (_zz_5232[31:0]         ), //i
    .dout    (fixTo_1193_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1194 (
    .din     (_zz_5233[31:0]         ), //i
    .dout    (fixTo_1194_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1195 (
    .din     (_zz_5234[31:0]         ), //i
    .dout    (fixTo_1195_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1196 (
    .din     (_zz_5235[31:0]         ), //i
    .dout    (fixTo_1196_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1197 (
    .din     (_zz_5236[31:0]         ), //i
    .dout    (fixTo_1197_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1198 (
    .din     (_zz_5237[31:0]         ), //i
    .dout    (fixTo_1198_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1199 (
    .din     (_zz_5238[31:0]         ), //i
    .dout    (fixTo_1199_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1200 (
    .din     (_zz_5239[31:0]         ), //i
    .dout    (fixTo_1200_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1201 (
    .din     (_zz_5240[31:0]         ), //i
    .dout    (fixTo_1201_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1202 (
    .din     (_zz_5241[31:0]         ), //i
    .dout    (fixTo_1202_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1203 (
    .din     (_zz_5242[31:0]         ), //i
    .dout    (fixTo_1203_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1204 (
    .din     (_zz_5243[31:0]         ), //i
    .dout    (fixTo_1204_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1205 (
    .din     (_zz_5244[31:0]         ), //i
    .dout    (fixTo_1205_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1206 (
    .din     (_zz_5245[31:0]         ), //i
    .dout    (fixTo_1206_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1207 (
    .din     (_zz_5246[31:0]         ), //i
    .dout    (fixTo_1207_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1208 (
    .din     (_zz_5247[31:0]         ), //i
    .dout    (fixTo_1208_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1209 (
    .din     (_zz_5248[31:0]         ), //i
    .dout    (fixTo_1209_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1210 (
    .din     (_zz_5249[31:0]         ), //i
    .dout    (fixTo_1210_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1211 (
    .din     (_zz_5250[31:0]         ), //i
    .dout    (fixTo_1211_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1212 (
    .din     (_zz_5251[31:0]         ), //i
    .dout    (fixTo_1212_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1213 (
    .din     (_zz_5252[31:0]         ), //i
    .dout    (fixTo_1213_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1214 (
    .din     (_zz_5253[31:0]         ), //i
    .dout    (fixTo_1214_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1215 (
    .din     (_zz_5254[31:0]         ), //i
    .dout    (fixTo_1215_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1216 (
    .din     (_zz_5255[31:0]         ), //i
    .dout    (fixTo_1216_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1217 (
    .din     (_zz_5256[31:0]         ), //i
    .dout    (fixTo_1217_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1218 (
    .din     (_zz_5257[31:0]         ), //i
    .dout    (fixTo_1218_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1219 (
    .din     (_zz_5258[31:0]         ), //i
    .dout    (fixTo_1219_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1220 (
    .din     (_zz_5259[31:0]         ), //i
    .dout    (fixTo_1220_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1221 (
    .din     (_zz_5260[31:0]         ), //i
    .dout    (fixTo_1221_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1222 (
    .din     (_zz_5261[31:0]         ), //i
    .dout    (fixTo_1222_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1223 (
    .din     (_zz_5262[31:0]         ), //i
    .dout    (fixTo_1223_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1224 (
    .din     (_zz_5263[31:0]         ), //i
    .dout    (fixTo_1224_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1225 (
    .din     (_zz_5264[31:0]         ), //i
    .dout    (fixTo_1225_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1226 (
    .din     (_zz_5265[31:0]         ), //i
    .dout    (fixTo_1226_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1227 (
    .din     (_zz_5266[31:0]         ), //i
    .dout    (fixTo_1227_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1228 (
    .din     (_zz_5267[31:0]         ), //i
    .dout    (fixTo_1228_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1229 (
    .din     (_zz_5268[31:0]         ), //i
    .dout    (fixTo_1229_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1230 (
    .din     (_zz_5269[31:0]         ), //i
    .dout    (fixTo_1230_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1231 (
    .din     (_zz_5270[31:0]         ), //i
    .dout    (fixTo_1231_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1232 (
    .din     (_zz_5271[31:0]         ), //i
    .dout    (fixTo_1232_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1233 (
    .din     (_zz_5272[31:0]         ), //i
    .dout    (fixTo_1233_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1234 (
    .din     (_zz_5273[31:0]         ), //i
    .dout    (fixTo_1234_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1235 (
    .din     (_zz_5274[31:0]         ), //i
    .dout    (fixTo_1235_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1236 (
    .din     (_zz_5275[31:0]         ), //i
    .dout    (fixTo_1236_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1237 (
    .din     (_zz_5276[31:0]         ), //i
    .dout    (fixTo_1237_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1238 (
    .din     (_zz_5277[31:0]         ), //i
    .dout    (fixTo_1238_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1239 (
    .din     (_zz_5278[31:0]         ), //i
    .dout    (fixTo_1239_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1240 (
    .din     (_zz_5279[31:0]         ), //i
    .dout    (fixTo_1240_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1241 (
    .din     (_zz_5280[31:0]         ), //i
    .dout    (fixTo_1241_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1242 (
    .din     (_zz_5281[31:0]         ), //i
    .dout    (fixTo_1242_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1243 (
    .din     (_zz_5282[31:0]         ), //i
    .dout    (fixTo_1243_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1244 (
    .din     (_zz_5283[31:0]         ), //i
    .dout    (fixTo_1244_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1245 (
    .din     (_zz_5284[31:0]         ), //i
    .dout    (fixTo_1245_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1246 (
    .din     (_zz_5285[31:0]         ), //i
    .dout    (fixTo_1246_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1247 (
    .din     (_zz_5286[31:0]         ), //i
    .dout    (fixTo_1247_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1248 (
    .din     (_zz_5287[31:0]         ), //i
    .dout    (fixTo_1248_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1249 (
    .din     (_zz_5288[31:0]         ), //i
    .dout    (fixTo_1249_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1250 (
    .din     (_zz_5289[31:0]         ), //i
    .dout    (fixTo_1250_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1251 (
    .din     (_zz_5290[31:0]         ), //i
    .dout    (fixTo_1251_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1252 (
    .din     (_zz_5291[31:0]         ), //i
    .dout    (fixTo_1252_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1253 (
    .din     (_zz_5292[31:0]         ), //i
    .dout    (fixTo_1253_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1254 (
    .din     (_zz_5293[31:0]         ), //i
    .dout    (fixTo_1254_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1255 (
    .din     (_zz_5294[31:0]         ), //i
    .dout    (fixTo_1255_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1256 (
    .din     (_zz_5295[31:0]         ), //i
    .dout    (fixTo_1256_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1257 (
    .din     (_zz_5296[31:0]         ), //i
    .dout    (fixTo_1257_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1258 (
    .din     (_zz_5297[31:0]         ), //i
    .dout    (fixTo_1258_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1259 (
    .din     (_zz_5298[31:0]         ), //i
    .dout    (fixTo_1259_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1260 (
    .din     (_zz_5299[31:0]         ), //i
    .dout    (fixTo_1260_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1261 (
    .din     (_zz_5300[31:0]         ), //i
    .dout    (fixTo_1261_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1262 (
    .din     (_zz_5301[31:0]         ), //i
    .dout    (fixTo_1262_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1263 (
    .din     (_zz_5302[31:0]         ), //i
    .dout    (fixTo_1263_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1264 (
    .din     (_zz_5303[31:0]         ), //i
    .dout    (fixTo_1264_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1265 (
    .din     (_zz_5304[31:0]         ), //i
    .dout    (fixTo_1265_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1266 (
    .din     (_zz_5305[31:0]         ), //i
    .dout    (fixTo_1266_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1267 (
    .din     (_zz_5306[31:0]         ), //i
    .dout    (fixTo_1267_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1268 (
    .din     (_zz_5307[31:0]         ), //i
    .dout    (fixTo_1268_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1269 (
    .din     (_zz_5308[31:0]         ), //i
    .dout    (fixTo_1269_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1270 (
    .din     (_zz_5309[31:0]         ), //i
    .dout    (fixTo_1270_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1271 (
    .din     (_zz_5310[31:0]         ), //i
    .dout    (fixTo_1271_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1272 (
    .din     (_zz_5311[31:0]         ), //i
    .dout    (fixTo_1272_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1273 (
    .din     (_zz_5312[31:0]         ), //i
    .dout    (fixTo_1273_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1274 (
    .din     (_zz_5313[31:0]         ), //i
    .dout    (fixTo_1274_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1275 (
    .din     (_zz_5314[31:0]         ), //i
    .dout    (fixTo_1275_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1276 (
    .din     (_zz_5315[31:0]         ), //i
    .dout    (fixTo_1276_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1277 (
    .din     (_zz_5316[31:0]         ), //i
    .dout    (fixTo_1277_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1278 (
    .din     (_zz_5317[31:0]         ), //i
    .dout    (fixTo_1278_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1279 (
    .din     (_zz_5318[31:0]         ), //i
    .dout    (fixTo_1279_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1280 (
    .din     (_zz_5319[31:0]         ), //i
    .dout    (fixTo_1280_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1281 (
    .din     (_zz_5320[31:0]         ), //i
    .dout    (fixTo_1281_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1282 (
    .din     (_zz_5321[31:0]         ), //i
    .dout    (fixTo_1282_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1283 (
    .din     (_zz_5322[31:0]         ), //i
    .dout    (fixTo_1283_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1284 (
    .din     (_zz_5323[31:0]         ), //i
    .dout    (fixTo_1284_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1285 (
    .din     (_zz_5324[31:0]         ), //i
    .dout    (fixTo_1285_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1286 (
    .din     (_zz_5325[31:0]         ), //i
    .dout    (fixTo_1286_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1287 (
    .din     (_zz_5326[31:0]         ), //i
    .dout    (fixTo_1287_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1288 (
    .din     (_zz_5327[31:0]         ), //i
    .dout    (fixTo_1288_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1289 (
    .din     (_zz_5328[31:0]         ), //i
    .dout    (fixTo_1289_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1290 (
    .din     (_zz_5329[31:0]         ), //i
    .dout    (fixTo_1290_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1291 (
    .din     (_zz_5330[31:0]         ), //i
    .dout    (fixTo_1291_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1292 (
    .din     (_zz_5331[31:0]         ), //i
    .dout    (fixTo_1292_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1293 (
    .din     (_zz_5332[31:0]         ), //i
    .dout    (fixTo_1293_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1294 (
    .din     (_zz_5333[31:0]         ), //i
    .dout    (fixTo_1294_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1295 (
    .din     (_zz_5334[31:0]         ), //i
    .dout    (fixTo_1295_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1296 (
    .din     (_zz_5335[31:0]         ), //i
    .dout    (fixTo_1296_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1297 (
    .din     (_zz_5336[31:0]         ), //i
    .dout    (fixTo_1297_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1298 (
    .din     (_zz_5337[31:0]         ), //i
    .dout    (fixTo_1298_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1299 (
    .din     (_zz_5338[31:0]         ), //i
    .dout    (fixTo_1299_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1300 (
    .din     (_zz_5339[31:0]         ), //i
    .dout    (fixTo_1300_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1301 (
    .din     (_zz_5340[31:0]         ), //i
    .dout    (fixTo_1301_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1302 (
    .din     (_zz_5341[31:0]         ), //i
    .dout    (fixTo_1302_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1303 (
    .din     (_zz_5342[31:0]         ), //i
    .dout    (fixTo_1303_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1304 (
    .din     (_zz_5343[31:0]         ), //i
    .dout    (fixTo_1304_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1305 (
    .din     (_zz_5344[31:0]         ), //i
    .dout    (fixTo_1305_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1306 (
    .din     (_zz_5345[31:0]         ), //i
    .dout    (fixTo_1306_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1307 (
    .din     (_zz_5346[31:0]         ), //i
    .dout    (fixTo_1307_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1308 (
    .din     (_zz_5347[31:0]         ), //i
    .dout    (fixTo_1308_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1309 (
    .din     (_zz_5348[31:0]         ), //i
    .dout    (fixTo_1309_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1310 (
    .din     (_zz_5349[31:0]         ), //i
    .dout    (fixTo_1310_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1311 (
    .din     (_zz_5350[31:0]         ), //i
    .dout    (fixTo_1311_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1312 (
    .din     (_zz_5351[31:0]         ), //i
    .dout    (fixTo_1312_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1313 (
    .din     (_zz_5352[31:0]         ), //i
    .dout    (fixTo_1313_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1314 (
    .din     (_zz_5353[31:0]         ), //i
    .dout    (fixTo_1314_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1315 (
    .din     (_zz_5354[31:0]         ), //i
    .dout    (fixTo_1315_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1316 (
    .din     (_zz_5355[31:0]         ), //i
    .dout    (fixTo_1316_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1317 (
    .din     (_zz_5356[31:0]         ), //i
    .dout    (fixTo_1317_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1318 (
    .din     (_zz_5357[31:0]         ), //i
    .dout    (fixTo_1318_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1319 (
    .din     (_zz_5358[31:0]         ), //i
    .dout    (fixTo_1319_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1320 (
    .din     (_zz_5359[31:0]         ), //i
    .dout    (fixTo_1320_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1321 (
    .din     (_zz_5360[31:0]         ), //i
    .dout    (fixTo_1321_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1322 (
    .din     (_zz_5361[31:0]         ), //i
    .dout    (fixTo_1322_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1323 (
    .din     (_zz_5362[31:0]         ), //i
    .dout    (fixTo_1323_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1324 (
    .din     (_zz_5363[31:0]         ), //i
    .dout    (fixTo_1324_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1325 (
    .din     (_zz_5364[31:0]         ), //i
    .dout    (fixTo_1325_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1326 (
    .din     (_zz_5365[31:0]         ), //i
    .dout    (fixTo_1326_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1327 (
    .din     (_zz_5366[31:0]         ), //i
    .dout    (fixTo_1327_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1328 (
    .din     (_zz_5367[31:0]         ), //i
    .dout    (fixTo_1328_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1329 (
    .din     (_zz_5368[31:0]         ), //i
    .dout    (fixTo_1329_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1330 (
    .din     (_zz_5369[31:0]         ), //i
    .dout    (fixTo_1330_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1331 (
    .din     (_zz_5370[31:0]         ), //i
    .dout    (fixTo_1331_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1332 (
    .din     (_zz_5371[31:0]         ), //i
    .dout    (fixTo_1332_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1333 (
    .din     (_zz_5372[31:0]         ), //i
    .dout    (fixTo_1333_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1334 (
    .din     (_zz_5373[31:0]         ), //i
    .dout    (fixTo_1334_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1335 (
    .din     (_zz_5374[31:0]         ), //i
    .dout    (fixTo_1335_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1336 (
    .din     (_zz_5375[31:0]         ), //i
    .dout    (fixTo_1336_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1337 (
    .din     (_zz_5376[31:0]         ), //i
    .dout    (fixTo_1337_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1338 (
    .din     (_zz_5377[31:0]         ), //i
    .dout    (fixTo_1338_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1339 (
    .din     (_zz_5378[31:0]         ), //i
    .dout    (fixTo_1339_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1340 (
    .din     (_zz_5379[31:0]         ), //i
    .dout    (fixTo_1340_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1341 (
    .din     (_zz_5380[31:0]         ), //i
    .dout    (fixTo_1341_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1342 (
    .din     (_zz_5381[31:0]         ), //i
    .dout    (fixTo_1342_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1343 (
    .din     (_zz_5382[31:0]         ), //i
    .dout    (fixTo_1343_dout[15:0]  )  //o
  );
  assign twiddle_factor_table_0_real = 16'h0100;
  assign twiddle_factor_table_0_imag = 16'h0;
  assign twiddle_factor_table_1_real = 16'h0100;
  assign twiddle_factor_table_1_imag = 16'h0;
  assign twiddle_factor_table_2_real = 16'h0;
  assign twiddle_factor_table_2_imag = 16'hff00;
  assign twiddle_factor_table_3_real = 16'h0100;
  assign twiddle_factor_table_3_imag = 16'h0;
  assign twiddle_factor_table_4_real = 16'h00b5;
  assign twiddle_factor_table_4_imag = 16'hff4b;
  assign twiddle_factor_table_5_real = 16'h0;
  assign twiddle_factor_table_5_imag = 16'hff00;
  assign twiddle_factor_table_6_real = 16'hff4b;
  assign twiddle_factor_table_6_imag = 16'hff4b;
  assign twiddle_factor_table_7_real = 16'h0100;
  assign twiddle_factor_table_7_imag = 16'h0;
  assign twiddle_factor_table_8_real = 16'h00ec;
  assign twiddle_factor_table_8_imag = 16'hff9f;
  assign twiddle_factor_table_9_real = 16'h00b5;
  assign twiddle_factor_table_9_imag = 16'hff4b;
  assign twiddle_factor_table_10_real = 16'h0061;
  assign twiddle_factor_table_10_imag = 16'hff14;
  assign twiddle_factor_table_11_real = 16'h0;
  assign twiddle_factor_table_11_imag = 16'hff00;
  assign twiddle_factor_table_12_real = 16'hff9f;
  assign twiddle_factor_table_12_imag = 16'hff14;
  assign twiddle_factor_table_13_real = 16'hff4b;
  assign twiddle_factor_table_13_imag = 16'hff4b;
  assign twiddle_factor_table_14_real = 16'hff14;
  assign twiddle_factor_table_14_imag = 16'hff9f;
  assign twiddle_factor_table_15_real = 16'h0100;
  assign twiddle_factor_table_15_imag = 16'h0;
  assign twiddle_factor_table_16_real = 16'h00fb;
  assign twiddle_factor_table_16_imag = 16'hffcf;
  assign twiddle_factor_table_17_real = 16'h00ec;
  assign twiddle_factor_table_17_imag = 16'hff9f;
  assign twiddle_factor_table_18_real = 16'h00d4;
  assign twiddle_factor_table_18_imag = 16'hff72;
  assign twiddle_factor_table_19_real = 16'h00b5;
  assign twiddle_factor_table_19_imag = 16'hff4b;
  assign twiddle_factor_table_20_real = 16'h008e;
  assign twiddle_factor_table_20_imag = 16'hff2c;
  assign twiddle_factor_table_21_real = 16'h0061;
  assign twiddle_factor_table_21_imag = 16'hff14;
  assign twiddle_factor_table_22_real = 16'h0031;
  assign twiddle_factor_table_22_imag = 16'hff05;
  assign twiddle_factor_table_23_real = 16'h0;
  assign twiddle_factor_table_23_imag = 16'hff00;
  assign twiddle_factor_table_24_real = 16'hffcf;
  assign twiddle_factor_table_24_imag = 16'hff05;
  assign twiddle_factor_table_25_real = 16'hff9f;
  assign twiddle_factor_table_25_imag = 16'hff14;
  assign twiddle_factor_table_26_real = 16'hff72;
  assign twiddle_factor_table_26_imag = 16'hff2c;
  assign twiddle_factor_table_27_real = 16'hff4b;
  assign twiddle_factor_table_27_imag = 16'hff4b;
  assign twiddle_factor_table_28_real = 16'hff2c;
  assign twiddle_factor_table_28_imag = 16'hff72;
  assign twiddle_factor_table_29_real = 16'hff14;
  assign twiddle_factor_table_29_imag = 16'hff9f;
  assign twiddle_factor_table_30_real = 16'hff05;
  assign twiddle_factor_table_30_imag = 16'hffcf;
  assign twiddle_factor_table_31_real = 16'h0100;
  assign twiddle_factor_table_31_imag = 16'h0;
  assign twiddle_factor_table_32_real = 16'h00fe;
  assign twiddle_factor_table_32_imag = 16'hffe7;
  assign twiddle_factor_table_33_real = 16'h00fb;
  assign twiddle_factor_table_33_imag = 16'hffcf;
  assign twiddle_factor_table_34_real = 16'h00f4;
  assign twiddle_factor_table_34_imag = 16'hffb6;
  assign twiddle_factor_table_35_real = 16'h00ec;
  assign twiddle_factor_table_35_imag = 16'hff9f;
  assign twiddle_factor_table_36_real = 16'h00e1;
  assign twiddle_factor_table_36_imag = 16'hff88;
  assign twiddle_factor_table_37_real = 16'h00d4;
  assign twiddle_factor_table_37_imag = 16'hff72;
  assign twiddle_factor_table_38_real = 16'h00c5;
  assign twiddle_factor_table_38_imag = 16'hff5e;
  assign twiddle_factor_table_39_real = 16'h00b5;
  assign twiddle_factor_table_39_imag = 16'hff4b;
  assign twiddle_factor_table_40_real = 16'h00a2;
  assign twiddle_factor_table_40_imag = 16'hff3b;
  assign twiddle_factor_table_41_real = 16'h008e;
  assign twiddle_factor_table_41_imag = 16'hff2c;
  assign twiddle_factor_table_42_real = 16'h0078;
  assign twiddle_factor_table_42_imag = 16'hff1f;
  assign twiddle_factor_table_43_real = 16'h0061;
  assign twiddle_factor_table_43_imag = 16'hff14;
  assign twiddle_factor_table_44_real = 16'h004a;
  assign twiddle_factor_table_44_imag = 16'hff0c;
  assign twiddle_factor_table_45_real = 16'h0031;
  assign twiddle_factor_table_45_imag = 16'hff05;
  assign twiddle_factor_table_46_real = 16'h0019;
  assign twiddle_factor_table_46_imag = 16'hff02;
  assign twiddle_factor_table_47_real = 16'h0;
  assign twiddle_factor_table_47_imag = 16'hff00;
  assign twiddle_factor_table_48_real = 16'hffe7;
  assign twiddle_factor_table_48_imag = 16'hff02;
  assign twiddle_factor_table_49_real = 16'hffcf;
  assign twiddle_factor_table_49_imag = 16'hff05;
  assign twiddle_factor_table_50_real = 16'hffb6;
  assign twiddle_factor_table_50_imag = 16'hff0c;
  assign twiddle_factor_table_51_real = 16'hff9f;
  assign twiddle_factor_table_51_imag = 16'hff14;
  assign twiddle_factor_table_52_real = 16'hff88;
  assign twiddle_factor_table_52_imag = 16'hff1f;
  assign twiddle_factor_table_53_real = 16'hff72;
  assign twiddle_factor_table_53_imag = 16'hff2c;
  assign twiddle_factor_table_54_real = 16'hff5e;
  assign twiddle_factor_table_54_imag = 16'hff3b;
  assign twiddle_factor_table_55_real = 16'hff4b;
  assign twiddle_factor_table_55_imag = 16'hff4b;
  assign twiddle_factor_table_56_real = 16'hff3b;
  assign twiddle_factor_table_56_imag = 16'hff5e;
  assign twiddle_factor_table_57_real = 16'hff2c;
  assign twiddle_factor_table_57_imag = 16'hff72;
  assign twiddle_factor_table_58_real = 16'hff1f;
  assign twiddle_factor_table_58_imag = 16'hff88;
  assign twiddle_factor_table_59_real = 16'hff14;
  assign twiddle_factor_table_59_imag = 16'hff9f;
  assign twiddle_factor_table_60_real = 16'hff0c;
  assign twiddle_factor_table_60_imag = 16'hffb6;
  assign twiddle_factor_table_61_real = 16'hff05;
  assign twiddle_factor_table_61_imag = 16'hffcf;
  assign twiddle_factor_table_62_real = 16'hff02;
  assign twiddle_factor_table_62_imag = 16'hffe7;
  assign twiddle_factor_table_63_real = 16'h0100;
  assign twiddle_factor_table_63_imag = 16'h0;
  assign twiddle_factor_table_64_real = 16'h00ff;
  assign twiddle_factor_table_64_imag = 16'hfff4;
  assign twiddle_factor_table_65_real = 16'h00fe;
  assign twiddle_factor_table_65_imag = 16'hffe7;
  assign twiddle_factor_table_66_real = 16'h00fd;
  assign twiddle_factor_table_66_imag = 16'hffdb;
  assign twiddle_factor_table_67_real = 16'h00fb;
  assign twiddle_factor_table_67_imag = 16'hffcf;
  assign twiddle_factor_table_68_real = 16'h00f8;
  assign twiddle_factor_table_68_imag = 16'hffc2;
  assign twiddle_factor_table_69_real = 16'h00f4;
  assign twiddle_factor_table_69_imag = 16'hffb6;
  assign twiddle_factor_table_70_real = 16'h00f1;
  assign twiddle_factor_table_70_imag = 16'hffaa;
  assign twiddle_factor_table_71_real = 16'h00ec;
  assign twiddle_factor_table_71_imag = 16'hff9f;
  assign twiddle_factor_table_72_real = 16'h00e7;
  assign twiddle_factor_table_72_imag = 16'hff93;
  assign twiddle_factor_table_73_real = 16'h00e1;
  assign twiddle_factor_table_73_imag = 16'hff88;
  assign twiddle_factor_table_74_real = 16'h00db;
  assign twiddle_factor_table_74_imag = 16'hff7d;
  assign twiddle_factor_table_75_real = 16'h00d4;
  assign twiddle_factor_table_75_imag = 16'hff72;
  assign twiddle_factor_table_76_real = 16'h00cd;
  assign twiddle_factor_table_76_imag = 16'hff68;
  assign twiddle_factor_table_77_real = 16'h00c5;
  assign twiddle_factor_table_77_imag = 16'hff5e;
  assign twiddle_factor_table_78_real = 16'h00bd;
  assign twiddle_factor_table_78_imag = 16'hff55;
  assign twiddle_factor_table_79_real = 16'h00b5;
  assign twiddle_factor_table_79_imag = 16'hff4b;
  assign twiddle_factor_table_80_real = 16'h00ab;
  assign twiddle_factor_table_80_imag = 16'hff43;
  assign twiddle_factor_table_81_real = 16'h00a2;
  assign twiddle_factor_table_81_imag = 16'hff3b;
  assign twiddle_factor_table_82_real = 16'h0098;
  assign twiddle_factor_table_82_imag = 16'hff33;
  assign twiddle_factor_table_83_real = 16'h008e;
  assign twiddle_factor_table_83_imag = 16'hff2c;
  assign twiddle_factor_table_84_real = 16'h0083;
  assign twiddle_factor_table_84_imag = 16'hff25;
  assign twiddle_factor_table_85_real = 16'h0078;
  assign twiddle_factor_table_85_imag = 16'hff1f;
  assign twiddle_factor_table_86_real = 16'h006d;
  assign twiddle_factor_table_86_imag = 16'hff19;
  assign twiddle_factor_table_87_real = 16'h0061;
  assign twiddle_factor_table_87_imag = 16'hff14;
  assign twiddle_factor_table_88_real = 16'h0056;
  assign twiddle_factor_table_88_imag = 16'hff0f;
  assign twiddle_factor_table_89_real = 16'h004a;
  assign twiddle_factor_table_89_imag = 16'hff0c;
  assign twiddle_factor_table_90_real = 16'h003e;
  assign twiddle_factor_table_90_imag = 16'hff08;
  assign twiddle_factor_table_91_real = 16'h0031;
  assign twiddle_factor_table_91_imag = 16'hff05;
  assign twiddle_factor_table_92_real = 16'h0025;
  assign twiddle_factor_table_92_imag = 16'hff03;
  assign twiddle_factor_table_93_real = 16'h0019;
  assign twiddle_factor_table_93_imag = 16'hff02;
  assign twiddle_factor_table_94_real = 16'h000c;
  assign twiddle_factor_table_94_imag = 16'hff01;
  assign twiddle_factor_table_95_real = 16'h0;
  assign twiddle_factor_table_95_imag = 16'hff00;
  assign twiddle_factor_table_96_real = 16'hfff4;
  assign twiddle_factor_table_96_imag = 16'hff01;
  assign twiddle_factor_table_97_real = 16'hffe7;
  assign twiddle_factor_table_97_imag = 16'hff02;
  assign twiddle_factor_table_98_real = 16'hffdb;
  assign twiddle_factor_table_98_imag = 16'hff03;
  assign twiddle_factor_table_99_real = 16'hffcf;
  assign twiddle_factor_table_99_imag = 16'hff05;
  assign twiddle_factor_table_100_real = 16'hffc2;
  assign twiddle_factor_table_100_imag = 16'hff08;
  assign twiddle_factor_table_101_real = 16'hffb6;
  assign twiddle_factor_table_101_imag = 16'hff0c;
  assign twiddle_factor_table_102_real = 16'hffaa;
  assign twiddle_factor_table_102_imag = 16'hff0f;
  assign twiddle_factor_table_103_real = 16'hff9f;
  assign twiddle_factor_table_103_imag = 16'hff14;
  assign twiddle_factor_table_104_real = 16'hff93;
  assign twiddle_factor_table_104_imag = 16'hff19;
  assign twiddle_factor_table_105_real = 16'hff88;
  assign twiddle_factor_table_105_imag = 16'hff1f;
  assign twiddle_factor_table_106_real = 16'hff7d;
  assign twiddle_factor_table_106_imag = 16'hff25;
  assign twiddle_factor_table_107_real = 16'hff72;
  assign twiddle_factor_table_107_imag = 16'hff2c;
  assign twiddle_factor_table_108_real = 16'hff68;
  assign twiddle_factor_table_108_imag = 16'hff33;
  assign twiddle_factor_table_109_real = 16'hff5e;
  assign twiddle_factor_table_109_imag = 16'hff3b;
  assign twiddle_factor_table_110_real = 16'hff55;
  assign twiddle_factor_table_110_imag = 16'hff43;
  assign twiddle_factor_table_111_real = 16'hff4b;
  assign twiddle_factor_table_111_imag = 16'hff4b;
  assign twiddle_factor_table_112_real = 16'hff43;
  assign twiddle_factor_table_112_imag = 16'hff55;
  assign twiddle_factor_table_113_real = 16'hff3b;
  assign twiddle_factor_table_113_imag = 16'hff5e;
  assign twiddle_factor_table_114_real = 16'hff33;
  assign twiddle_factor_table_114_imag = 16'hff68;
  assign twiddle_factor_table_115_real = 16'hff2c;
  assign twiddle_factor_table_115_imag = 16'hff72;
  assign twiddle_factor_table_116_real = 16'hff25;
  assign twiddle_factor_table_116_imag = 16'hff7d;
  assign twiddle_factor_table_117_real = 16'hff1f;
  assign twiddle_factor_table_117_imag = 16'hff88;
  assign twiddle_factor_table_118_real = 16'hff19;
  assign twiddle_factor_table_118_imag = 16'hff93;
  assign twiddle_factor_table_119_real = 16'hff14;
  assign twiddle_factor_table_119_imag = 16'hff9f;
  assign twiddle_factor_table_120_real = 16'hff0f;
  assign twiddle_factor_table_120_imag = 16'hffaa;
  assign twiddle_factor_table_121_real = 16'hff0c;
  assign twiddle_factor_table_121_imag = 16'hffb6;
  assign twiddle_factor_table_122_real = 16'hff08;
  assign twiddle_factor_table_122_imag = 16'hffc2;
  assign twiddle_factor_table_123_real = 16'hff05;
  assign twiddle_factor_table_123_imag = 16'hffcf;
  assign twiddle_factor_table_124_real = 16'hff03;
  assign twiddle_factor_table_124_imag = 16'hffdb;
  assign twiddle_factor_table_125_real = 16'hff02;
  assign twiddle_factor_table_125_imag = 16'hffe7;
  assign twiddle_factor_table_126_real = 16'hff01;
  assign twiddle_factor_table_126_imag = 16'hfff4;
  assign data_reorder_0_real = data_in_0_real;
  assign data_reorder_0_imag = data_in_0_imag;
  assign data_reorder_64_real = data_in_1_real;
  assign data_reorder_64_imag = data_in_1_imag;
  assign data_reorder_32_real = data_in_2_real;
  assign data_reorder_32_imag = data_in_2_imag;
  assign data_reorder_96_real = data_in_3_real;
  assign data_reorder_96_imag = data_in_3_imag;
  assign data_reorder_16_real = data_in_4_real;
  assign data_reorder_16_imag = data_in_4_imag;
  assign data_reorder_80_real = data_in_5_real;
  assign data_reorder_80_imag = data_in_5_imag;
  assign data_reorder_48_real = data_in_6_real;
  assign data_reorder_48_imag = data_in_6_imag;
  assign data_reorder_112_real = data_in_7_real;
  assign data_reorder_112_imag = data_in_7_imag;
  assign data_reorder_8_real = data_in_8_real;
  assign data_reorder_8_imag = data_in_8_imag;
  assign data_reorder_72_real = data_in_9_real;
  assign data_reorder_72_imag = data_in_9_imag;
  assign data_reorder_40_real = data_in_10_real;
  assign data_reorder_40_imag = data_in_10_imag;
  assign data_reorder_104_real = data_in_11_real;
  assign data_reorder_104_imag = data_in_11_imag;
  assign data_reorder_24_real = data_in_12_real;
  assign data_reorder_24_imag = data_in_12_imag;
  assign data_reorder_88_real = data_in_13_real;
  assign data_reorder_88_imag = data_in_13_imag;
  assign data_reorder_56_real = data_in_14_real;
  assign data_reorder_56_imag = data_in_14_imag;
  assign data_reorder_120_real = data_in_15_real;
  assign data_reorder_120_imag = data_in_15_imag;
  assign data_reorder_4_real = data_in_16_real;
  assign data_reorder_4_imag = data_in_16_imag;
  assign data_reorder_68_real = data_in_17_real;
  assign data_reorder_68_imag = data_in_17_imag;
  assign data_reorder_36_real = data_in_18_real;
  assign data_reorder_36_imag = data_in_18_imag;
  assign data_reorder_100_real = data_in_19_real;
  assign data_reorder_100_imag = data_in_19_imag;
  assign data_reorder_20_real = data_in_20_real;
  assign data_reorder_20_imag = data_in_20_imag;
  assign data_reorder_84_real = data_in_21_real;
  assign data_reorder_84_imag = data_in_21_imag;
  assign data_reorder_52_real = data_in_22_real;
  assign data_reorder_52_imag = data_in_22_imag;
  assign data_reorder_116_real = data_in_23_real;
  assign data_reorder_116_imag = data_in_23_imag;
  assign data_reorder_12_real = data_in_24_real;
  assign data_reorder_12_imag = data_in_24_imag;
  assign data_reorder_76_real = data_in_25_real;
  assign data_reorder_76_imag = data_in_25_imag;
  assign data_reorder_44_real = data_in_26_real;
  assign data_reorder_44_imag = data_in_26_imag;
  assign data_reorder_108_real = data_in_27_real;
  assign data_reorder_108_imag = data_in_27_imag;
  assign data_reorder_28_real = data_in_28_real;
  assign data_reorder_28_imag = data_in_28_imag;
  assign data_reorder_92_real = data_in_29_real;
  assign data_reorder_92_imag = data_in_29_imag;
  assign data_reorder_60_real = data_in_30_real;
  assign data_reorder_60_imag = data_in_30_imag;
  assign data_reorder_124_real = data_in_31_real;
  assign data_reorder_124_imag = data_in_31_imag;
  assign data_reorder_2_real = data_in_32_real;
  assign data_reorder_2_imag = data_in_32_imag;
  assign data_reorder_66_real = data_in_33_real;
  assign data_reorder_66_imag = data_in_33_imag;
  assign data_reorder_34_real = data_in_34_real;
  assign data_reorder_34_imag = data_in_34_imag;
  assign data_reorder_98_real = data_in_35_real;
  assign data_reorder_98_imag = data_in_35_imag;
  assign data_reorder_18_real = data_in_36_real;
  assign data_reorder_18_imag = data_in_36_imag;
  assign data_reorder_82_real = data_in_37_real;
  assign data_reorder_82_imag = data_in_37_imag;
  assign data_reorder_50_real = data_in_38_real;
  assign data_reorder_50_imag = data_in_38_imag;
  assign data_reorder_114_real = data_in_39_real;
  assign data_reorder_114_imag = data_in_39_imag;
  assign data_reorder_10_real = data_in_40_real;
  assign data_reorder_10_imag = data_in_40_imag;
  assign data_reorder_74_real = data_in_41_real;
  assign data_reorder_74_imag = data_in_41_imag;
  assign data_reorder_42_real = data_in_42_real;
  assign data_reorder_42_imag = data_in_42_imag;
  assign data_reorder_106_real = data_in_43_real;
  assign data_reorder_106_imag = data_in_43_imag;
  assign data_reorder_26_real = data_in_44_real;
  assign data_reorder_26_imag = data_in_44_imag;
  assign data_reorder_90_real = data_in_45_real;
  assign data_reorder_90_imag = data_in_45_imag;
  assign data_reorder_58_real = data_in_46_real;
  assign data_reorder_58_imag = data_in_46_imag;
  assign data_reorder_122_real = data_in_47_real;
  assign data_reorder_122_imag = data_in_47_imag;
  assign data_reorder_6_real = data_in_48_real;
  assign data_reorder_6_imag = data_in_48_imag;
  assign data_reorder_70_real = data_in_49_real;
  assign data_reorder_70_imag = data_in_49_imag;
  assign data_reorder_38_real = data_in_50_real;
  assign data_reorder_38_imag = data_in_50_imag;
  assign data_reorder_102_real = data_in_51_real;
  assign data_reorder_102_imag = data_in_51_imag;
  assign data_reorder_22_real = data_in_52_real;
  assign data_reorder_22_imag = data_in_52_imag;
  assign data_reorder_86_real = data_in_53_real;
  assign data_reorder_86_imag = data_in_53_imag;
  assign data_reorder_54_real = data_in_54_real;
  assign data_reorder_54_imag = data_in_54_imag;
  assign data_reorder_118_real = data_in_55_real;
  assign data_reorder_118_imag = data_in_55_imag;
  assign data_reorder_14_real = data_in_56_real;
  assign data_reorder_14_imag = data_in_56_imag;
  assign data_reorder_78_real = data_in_57_real;
  assign data_reorder_78_imag = data_in_57_imag;
  assign data_reorder_46_real = data_in_58_real;
  assign data_reorder_46_imag = data_in_58_imag;
  assign data_reorder_110_real = data_in_59_real;
  assign data_reorder_110_imag = data_in_59_imag;
  assign data_reorder_30_real = data_in_60_real;
  assign data_reorder_30_imag = data_in_60_imag;
  assign data_reorder_94_real = data_in_61_real;
  assign data_reorder_94_imag = data_in_61_imag;
  assign data_reorder_62_real = data_in_62_real;
  assign data_reorder_62_imag = data_in_62_imag;
  assign data_reorder_126_real = data_in_63_real;
  assign data_reorder_126_imag = data_in_63_imag;
  assign data_reorder_1_real = data_in_64_real;
  assign data_reorder_1_imag = data_in_64_imag;
  assign data_reorder_65_real = data_in_65_real;
  assign data_reorder_65_imag = data_in_65_imag;
  assign data_reorder_33_real = data_in_66_real;
  assign data_reorder_33_imag = data_in_66_imag;
  assign data_reorder_97_real = data_in_67_real;
  assign data_reorder_97_imag = data_in_67_imag;
  assign data_reorder_17_real = data_in_68_real;
  assign data_reorder_17_imag = data_in_68_imag;
  assign data_reorder_81_real = data_in_69_real;
  assign data_reorder_81_imag = data_in_69_imag;
  assign data_reorder_49_real = data_in_70_real;
  assign data_reorder_49_imag = data_in_70_imag;
  assign data_reorder_113_real = data_in_71_real;
  assign data_reorder_113_imag = data_in_71_imag;
  assign data_reorder_9_real = data_in_72_real;
  assign data_reorder_9_imag = data_in_72_imag;
  assign data_reorder_73_real = data_in_73_real;
  assign data_reorder_73_imag = data_in_73_imag;
  assign data_reorder_41_real = data_in_74_real;
  assign data_reorder_41_imag = data_in_74_imag;
  assign data_reorder_105_real = data_in_75_real;
  assign data_reorder_105_imag = data_in_75_imag;
  assign data_reorder_25_real = data_in_76_real;
  assign data_reorder_25_imag = data_in_76_imag;
  assign data_reorder_89_real = data_in_77_real;
  assign data_reorder_89_imag = data_in_77_imag;
  assign data_reorder_57_real = data_in_78_real;
  assign data_reorder_57_imag = data_in_78_imag;
  assign data_reorder_121_real = data_in_79_real;
  assign data_reorder_121_imag = data_in_79_imag;
  assign data_reorder_5_real = data_in_80_real;
  assign data_reorder_5_imag = data_in_80_imag;
  assign data_reorder_69_real = data_in_81_real;
  assign data_reorder_69_imag = data_in_81_imag;
  assign data_reorder_37_real = data_in_82_real;
  assign data_reorder_37_imag = data_in_82_imag;
  assign data_reorder_101_real = data_in_83_real;
  assign data_reorder_101_imag = data_in_83_imag;
  assign data_reorder_21_real = data_in_84_real;
  assign data_reorder_21_imag = data_in_84_imag;
  assign data_reorder_85_real = data_in_85_real;
  assign data_reorder_85_imag = data_in_85_imag;
  assign data_reorder_53_real = data_in_86_real;
  assign data_reorder_53_imag = data_in_86_imag;
  assign data_reorder_117_real = data_in_87_real;
  assign data_reorder_117_imag = data_in_87_imag;
  assign data_reorder_13_real = data_in_88_real;
  assign data_reorder_13_imag = data_in_88_imag;
  assign data_reorder_77_real = data_in_89_real;
  assign data_reorder_77_imag = data_in_89_imag;
  assign data_reorder_45_real = data_in_90_real;
  assign data_reorder_45_imag = data_in_90_imag;
  assign data_reorder_109_real = data_in_91_real;
  assign data_reorder_109_imag = data_in_91_imag;
  assign data_reorder_29_real = data_in_92_real;
  assign data_reorder_29_imag = data_in_92_imag;
  assign data_reorder_93_real = data_in_93_real;
  assign data_reorder_93_imag = data_in_93_imag;
  assign data_reorder_61_real = data_in_94_real;
  assign data_reorder_61_imag = data_in_94_imag;
  assign data_reorder_125_real = data_in_95_real;
  assign data_reorder_125_imag = data_in_95_imag;
  assign data_reorder_3_real = data_in_96_real;
  assign data_reorder_3_imag = data_in_96_imag;
  assign data_reorder_67_real = data_in_97_real;
  assign data_reorder_67_imag = data_in_97_imag;
  assign data_reorder_35_real = data_in_98_real;
  assign data_reorder_35_imag = data_in_98_imag;
  assign data_reorder_99_real = data_in_99_real;
  assign data_reorder_99_imag = data_in_99_imag;
  assign data_reorder_19_real = data_in_100_real;
  assign data_reorder_19_imag = data_in_100_imag;
  assign data_reorder_83_real = data_in_101_real;
  assign data_reorder_83_imag = data_in_101_imag;
  assign data_reorder_51_real = data_in_102_real;
  assign data_reorder_51_imag = data_in_102_imag;
  assign data_reorder_115_real = data_in_103_real;
  assign data_reorder_115_imag = data_in_103_imag;
  assign data_reorder_11_real = data_in_104_real;
  assign data_reorder_11_imag = data_in_104_imag;
  assign data_reorder_75_real = data_in_105_real;
  assign data_reorder_75_imag = data_in_105_imag;
  assign data_reorder_43_real = data_in_106_real;
  assign data_reorder_43_imag = data_in_106_imag;
  assign data_reorder_107_real = data_in_107_real;
  assign data_reorder_107_imag = data_in_107_imag;
  assign data_reorder_27_real = data_in_108_real;
  assign data_reorder_27_imag = data_in_108_imag;
  assign data_reorder_91_real = data_in_109_real;
  assign data_reorder_91_imag = data_in_109_imag;
  assign data_reorder_59_real = data_in_110_real;
  assign data_reorder_59_imag = data_in_110_imag;
  assign data_reorder_123_real = data_in_111_real;
  assign data_reorder_123_imag = data_in_111_imag;
  assign data_reorder_7_real = data_in_112_real;
  assign data_reorder_7_imag = data_in_112_imag;
  assign data_reorder_71_real = data_in_113_real;
  assign data_reorder_71_imag = data_in_113_imag;
  assign data_reorder_39_real = data_in_114_real;
  assign data_reorder_39_imag = data_in_114_imag;
  assign data_reorder_103_real = data_in_115_real;
  assign data_reorder_103_imag = data_in_115_imag;
  assign data_reorder_23_real = data_in_116_real;
  assign data_reorder_23_imag = data_in_116_imag;
  assign data_reorder_87_real = data_in_117_real;
  assign data_reorder_87_imag = data_in_117_imag;
  assign data_reorder_55_real = data_in_118_real;
  assign data_reorder_55_imag = data_in_118_imag;
  assign data_reorder_119_real = data_in_119_real;
  assign data_reorder_119_imag = data_in_119_imag;
  assign data_reorder_15_real = data_in_120_real;
  assign data_reorder_15_imag = data_in_120_imag;
  assign data_reorder_79_real = data_in_121_real;
  assign data_reorder_79_imag = data_in_121_imag;
  assign data_reorder_47_real = data_in_122_real;
  assign data_reorder_47_imag = data_in_122_imag;
  assign data_reorder_111_real = data_in_123_real;
  assign data_reorder_111_imag = data_in_123_imag;
  assign data_reorder_31_real = data_in_124_real;
  assign data_reorder_31_imag = data_in_124_imag;
  assign data_reorder_95_real = data_in_125_real;
  assign data_reorder_95_imag = data_in_125_imag;
  assign data_reorder_63_real = data_in_126_real;
  assign data_reorder_63_imag = data_in_126_imag;
  assign data_reorder_127_real = data_in_127_real;
  assign data_reorder_127_imag = data_in_127_imag;
  assign _zz_4039 = ($signed(_zz_5383) * $signed(_zz_3));
  assign _zz_1795 = _zz_5384[15 : 0];
  assign _zz_4040 = ($signed(_zz_5385) * $signed(twiddle_factor_table_0_real));
  assign _zz_4041 = ($signed(_zz_5386) * $signed(twiddle_factor_table_0_imag));
  assign _zz_1793 = ($signed(_zz_1795) - $signed(_zz_5387));
  assign _zz_1794 = ($signed(_zz_1795) + $signed(_zz_5389));
  assign _zz_1796 = 1'b1;
  assign _zz_1797 = 1'b1;
  assign _zz_4042 = ($signed(_zz_5407) * $signed(_zz_7));
  assign _zz_1800 = _zz_5408[15 : 0];
  assign _zz_4043 = ($signed(_zz_5409) * $signed(twiddle_factor_table_0_real));
  assign _zz_4044 = ($signed(_zz_5410) * $signed(twiddle_factor_table_0_imag));
  assign _zz_1798 = ($signed(_zz_1800) - $signed(_zz_5411));
  assign _zz_1799 = ($signed(_zz_1800) + $signed(_zz_5413));
  assign _zz_1801 = 1'b1;
  assign _zz_1802 = 1'b1;
  assign _zz_4045 = ($signed(_zz_5431) * $signed(_zz_11));
  assign _zz_1805 = _zz_5432[15 : 0];
  assign _zz_4046 = ($signed(_zz_5433) * $signed(twiddle_factor_table_0_real));
  assign _zz_4047 = ($signed(_zz_5434) * $signed(twiddle_factor_table_0_imag));
  assign _zz_1803 = ($signed(_zz_1805) - $signed(_zz_5435));
  assign _zz_1804 = ($signed(_zz_1805) + $signed(_zz_5437));
  assign _zz_1806 = 1'b1;
  assign _zz_1807 = 1'b1;
  assign _zz_4048 = ($signed(_zz_5455) * $signed(_zz_15));
  assign _zz_1810 = _zz_5456[15 : 0];
  assign _zz_4049 = ($signed(_zz_5457) * $signed(twiddle_factor_table_0_real));
  assign _zz_4050 = ($signed(_zz_5458) * $signed(twiddle_factor_table_0_imag));
  assign _zz_1808 = ($signed(_zz_1810) - $signed(_zz_5459));
  assign _zz_1809 = ($signed(_zz_1810) + $signed(_zz_5461));
  assign _zz_1811 = 1'b1;
  assign _zz_1812 = 1'b1;
  assign _zz_4051 = ($signed(_zz_5479) * $signed(_zz_19));
  assign _zz_1815 = _zz_5480[15 : 0];
  assign _zz_4052 = ($signed(_zz_5481) * $signed(twiddle_factor_table_0_real));
  assign _zz_4053 = ($signed(_zz_5482) * $signed(twiddle_factor_table_0_imag));
  assign _zz_1813 = ($signed(_zz_1815) - $signed(_zz_5483));
  assign _zz_1814 = ($signed(_zz_1815) + $signed(_zz_5485));
  assign _zz_1816 = 1'b1;
  assign _zz_1817 = 1'b1;
  assign _zz_4054 = ($signed(_zz_5503) * $signed(_zz_23));
  assign _zz_1820 = _zz_5504[15 : 0];
  assign _zz_4055 = ($signed(_zz_5505) * $signed(twiddle_factor_table_0_real));
  assign _zz_4056 = ($signed(_zz_5506) * $signed(twiddle_factor_table_0_imag));
  assign _zz_1818 = ($signed(_zz_1820) - $signed(_zz_5507));
  assign _zz_1819 = ($signed(_zz_1820) + $signed(_zz_5509));
  assign _zz_1821 = 1'b1;
  assign _zz_1822 = 1'b1;
  assign _zz_4057 = ($signed(_zz_5527) * $signed(_zz_27));
  assign _zz_1825 = _zz_5528[15 : 0];
  assign _zz_4058 = ($signed(_zz_5529) * $signed(twiddle_factor_table_0_real));
  assign _zz_4059 = ($signed(_zz_5530) * $signed(twiddle_factor_table_0_imag));
  assign _zz_1823 = ($signed(_zz_1825) - $signed(_zz_5531));
  assign _zz_1824 = ($signed(_zz_1825) + $signed(_zz_5533));
  assign _zz_1826 = 1'b1;
  assign _zz_1827 = 1'b1;
  assign _zz_4060 = ($signed(_zz_5551) * $signed(_zz_31));
  assign _zz_1830 = _zz_5552[15 : 0];
  assign _zz_4061 = ($signed(_zz_5553) * $signed(twiddle_factor_table_0_real));
  assign _zz_4062 = ($signed(_zz_5554) * $signed(twiddle_factor_table_0_imag));
  assign _zz_1828 = ($signed(_zz_1830) - $signed(_zz_5555));
  assign _zz_1829 = ($signed(_zz_1830) + $signed(_zz_5557));
  assign _zz_1831 = 1'b1;
  assign _zz_1832 = 1'b1;
  assign _zz_4063 = ($signed(_zz_5575) * $signed(_zz_35));
  assign _zz_1835 = _zz_5576[15 : 0];
  assign _zz_4064 = ($signed(_zz_5577) * $signed(twiddle_factor_table_0_real));
  assign _zz_4065 = ($signed(_zz_5578) * $signed(twiddle_factor_table_0_imag));
  assign _zz_1833 = ($signed(_zz_1835) - $signed(_zz_5579));
  assign _zz_1834 = ($signed(_zz_1835) + $signed(_zz_5581));
  assign _zz_1836 = 1'b1;
  assign _zz_1837 = 1'b1;
  assign _zz_4066 = ($signed(_zz_5599) * $signed(_zz_39));
  assign _zz_1840 = _zz_5600[15 : 0];
  assign _zz_4067 = ($signed(_zz_5601) * $signed(twiddle_factor_table_0_real));
  assign _zz_4068 = ($signed(_zz_5602) * $signed(twiddle_factor_table_0_imag));
  assign _zz_1838 = ($signed(_zz_1840) - $signed(_zz_5603));
  assign _zz_1839 = ($signed(_zz_1840) + $signed(_zz_5605));
  assign _zz_1841 = 1'b1;
  assign _zz_1842 = 1'b1;
  assign _zz_4069 = ($signed(_zz_5623) * $signed(_zz_43));
  assign _zz_1845 = _zz_5624[15 : 0];
  assign _zz_4070 = ($signed(_zz_5625) * $signed(twiddle_factor_table_0_real));
  assign _zz_4071 = ($signed(_zz_5626) * $signed(twiddle_factor_table_0_imag));
  assign _zz_1843 = ($signed(_zz_1845) - $signed(_zz_5627));
  assign _zz_1844 = ($signed(_zz_1845) + $signed(_zz_5629));
  assign _zz_1846 = 1'b1;
  assign _zz_1847 = 1'b1;
  assign _zz_4072 = ($signed(_zz_5647) * $signed(_zz_47));
  assign _zz_1850 = _zz_5648[15 : 0];
  assign _zz_4073 = ($signed(_zz_5649) * $signed(twiddle_factor_table_0_real));
  assign _zz_4074 = ($signed(_zz_5650) * $signed(twiddle_factor_table_0_imag));
  assign _zz_1848 = ($signed(_zz_1850) - $signed(_zz_5651));
  assign _zz_1849 = ($signed(_zz_1850) + $signed(_zz_5653));
  assign _zz_1851 = 1'b1;
  assign _zz_1852 = 1'b1;
  assign _zz_4075 = ($signed(_zz_5671) * $signed(_zz_51));
  assign _zz_1855 = _zz_5672[15 : 0];
  assign _zz_4076 = ($signed(_zz_5673) * $signed(twiddle_factor_table_0_real));
  assign _zz_4077 = ($signed(_zz_5674) * $signed(twiddle_factor_table_0_imag));
  assign _zz_1853 = ($signed(_zz_1855) - $signed(_zz_5675));
  assign _zz_1854 = ($signed(_zz_1855) + $signed(_zz_5677));
  assign _zz_1856 = 1'b1;
  assign _zz_1857 = 1'b1;
  assign _zz_4078 = ($signed(_zz_5695) * $signed(_zz_55));
  assign _zz_1860 = _zz_5696[15 : 0];
  assign _zz_4079 = ($signed(_zz_5697) * $signed(twiddle_factor_table_0_real));
  assign _zz_4080 = ($signed(_zz_5698) * $signed(twiddle_factor_table_0_imag));
  assign _zz_1858 = ($signed(_zz_1860) - $signed(_zz_5699));
  assign _zz_1859 = ($signed(_zz_1860) + $signed(_zz_5701));
  assign _zz_1861 = 1'b1;
  assign _zz_1862 = 1'b1;
  assign _zz_4081 = ($signed(_zz_5719) * $signed(_zz_59));
  assign _zz_1865 = _zz_5720[15 : 0];
  assign _zz_4082 = ($signed(_zz_5721) * $signed(twiddle_factor_table_0_real));
  assign _zz_4083 = ($signed(_zz_5722) * $signed(twiddle_factor_table_0_imag));
  assign _zz_1863 = ($signed(_zz_1865) - $signed(_zz_5723));
  assign _zz_1864 = ($signed(_zz_1865) + $signed(_zz_5725));
  assign _zz_1866 = 1'b1;
  assign _zz_1867 = 1'b1;
  assign _zz_4084 = ($signed(_zz_5743) * $signed(_zz_63));
  assign _zz_1870 = _zz_5744[15 : 0];
  assign _zz_4085 = ($signed(_zz_5745) * $signed(twiddle_factor_table_0_real));
  assign _zz_4086 = ($signed(_zz_5746) * $signed(twiddle_factor_table_0_imag));
  assign _zz_1868 = ($signed(_zz_1870) - $signed(_zz_5747));
  assign _zz_1869 = ($signed(_zz_1870) + $signed(_zz_5749));
  assign _zz_1871 = 1'b1;
  assign _zz_1872 = 1'b1;
  assign _zz_4087 = ($signed(_zz_5767) * $signed(_zz_67));
  assign _zz_1875 = _zz_5768[15 : 0];
  assign _zz_4088 = ($signed(_zz_5769) * $signed(twiddle_factor_table_0_real));
  assign _zz_4089 = ($signed(_zz_5770) * $signed(twiddle_factor_table_0_imag));
  assign _zz_1873 = ($signed(_zz_1875) - $signed(_zz_5771));
  assign _zz_1874 = ($signed(_zz_1875) + $signed(_zz_5773));
  assign _zz_1876 = 1'b1;
  assign _zz_1877 = 1'b1;
  assign _zz_4090 = ($signed(_zz_5791) * $signed(_zz_71));
  assign _zz_1880 = _zz_5792[15 : 0];
  assign _zz_4091 = ($signed(_zz_5793) * $signed(twiddle_factor_table_0_real));
  assign _zz_4092 = ($signed(_zz_5794) * $signed(twiddle_factor_table_0_imag));
  assign _zz_1878 = ($signed(_zz_1880) - $signed(_zz_5795));
  assign _zz_1879 = ($signed(_zz_1880) + $signed(_zz_5797));
  assign _zz_1881 = 1'b1;
  assign _zz_1882 = 1'b1;
  assign _zz_4093 = ($signed(_zz_5815) * $signed(_zz_75));
  assign _zz_1885 = _zz_5816[15 : 0];
  assign _zz_4094 = ($signed(_zz_5817) * $signed(twiddle_factor_table_0_real));
  assign _zz_4095 = ($signed(_zz_5818) * $signed(twiddle_factor_table_0_imag));
  assign _zz_1883 = ($signed(_zz_1885) - $signed(_zz_5819));
  assign _zz_1884 = ($signed(_zz_1885) + $signed(_zz_5821));
  assign _zz_1886 = 1'b1;
  assign _zz_1887 = 1'b1;
  assign _zz_4096 = ($signed(_zz_5839) * $signed(_zz_79));
  assign _zz_1890 = _zz_5840[15 : 0];
  assign _zz_4097 = ($signed(_zz_5841) * $signed(twiddle_factor_table_0_real));
  assign _zz_4098 = ($signed(_zz_5842) * $signed(twiddle_factor_table_0_imag));
  assign _zz_1888 = ($signed(_zz_1890) - $signed(_zz_5843));
  assign _zz_1889 = ($signed(_zz_1890) + $signed(_zz_5845));
  assign _zz_1891 = 1'b1;
  assign _zz_1892 = 1'b1;
  assign _zz_4099 = ($signed(_zz_5863) * $signed(_zz_83));
  assign _zz_1895 = _zz_5864[15 : 0];
  assign _zz_4100 = ($signed(_zz_5865) * $signed(twiddle_factor_table_0_real));
  assign _zz_4101 = ($signed(_zz_5866) * $signed(twiddle_factor_table_0_imag));
  assign _zz_1893 = ($signed(_zz_1895) - $signed(_zz_5867));
  assign _zz_1894 = ($signed(_zz_1895) + $signed(_zz_5869));
  assign _zz_1896 = 1'b1;
  assign _zz_1897 = 1'b1;
  assign _zz_4102 = ($signed(_zz_5887) * $signed(_zz_87));
  assign _zz_1900 = _zz_5888[15 : 0];
  assign _zz_4103 = ($signed(_zz_5889) * $signed(twiddle_factor_table_0_real));
  assign _zz_4104 = ($signed(_zz_5890) * $signed(twiddle_factor_table_0_imag));
  assign _zz_1898 = ($signed(_zz_1900) - $signed(_zz_5891));
  assign _zz_1899 = ($signed(_zz_1900) + $signed(_zz_5893));
  assign _zz_1901 = 1'b1;
  assign _zz_1902 = 1'b1;
  assign _zz_4105 = ($signed(_zz_5911) * $signed(_zz_91));
  assign _zz_1905 = _zz_5912[15 : 0];
  assign _zz_4106 = ($signed(_zz_5913) * $signed(twiddle_factor_table_0_real));
  assign _zz_4107 = ($signed(_zz_5914) * $signed(twiddle_factor_table_0_imag));
  assign _zz_1903 = ($signed(_zz_1905) - $signed(_zz_5915));
  assign _zz_1904 = ($signed(_zz_1905) + $signed(_zz_5917));
  assign _zz_1906 = 1'b1;
  assign _zz_1907 = 1'b1;
  assign _zz_4108 = ($signed(_zz_5935) * $signed(_zz_95));
  assign _zz_1910 = _zz_5936[15 : 0];
  assign _zz_4109 = ($signed(_zz_5937) * $signed(twiddle_factor_table_0_real));
  assign _zz_4110 = ($signed(_zz_5938) * $signed(twiddle_factor_table_0_imag));
  assign _zz_1908 = ($signed(_zz_1910) - $signed(_zz_5939));
  assign _zz_1909 = ($signed(_zz_1910) + $signed(_zz_5941));
  assign _zz_1911 = 1'b1;
  assign _zz_1912 = 1'b1;
  assign _zz_4111 = ($signed(_zz_5959) * $signed(_zz_99));
  assign _zz_1915 = _zz_5960[15 : 0];
  assign _zz_4112 = ($signed(_zz_5961) * $signed(twiddle_factor_table_0_real));
  assign _zz_4113 = ($signed(_zz_5962) * $signed(twiddle_factor_table_0_imag));
  assign _zz_1913 = ($signed(_zz_1915) - $signed(_zz_5963));
  assign _zz_1914 = ($signed(_zz_1915) + $signed(_zz_5965));
  assign _zz_1916 = 1'b1;
  assign _zz_1917 = 1'b1;
  assign _zz_4114 = ($signed(_zz_5983) * $signed(_zz_103));
  assign _zz_1920 = _zz_5984[15 : 0];
  assign _zz_4115 = ($signed(_zz_5985) * $signed(twiddle_factor_table_0_real));
  assign _zz_4116 = ($signed(_zz_5986) * $signed(twiddle_factor_table_0_imag));
  assign _zz_1918 = ($signed(_zz_1920) - $signed(_zz_5987));
  assign _zz_1919 = ($signed(_zz_1920) + $signed(_zz_5989));
  assign _zz_1921 = 1'b1;
  assign _zz_1922 = 1'b1;
  assign _zz_4117 = ($signed(_zz_6007) * $signed(_zz_107));
  assign _zz_1925 = _zz_6008[15 : 0];
  assign _zz_4118 = ($signed(_zz_6009) * $signed(twiddle_factor_table_0_real));
  assign _zz_4119 = ($signed(_zz_6010) * $signed(twiddle_factor_table_0_imag));
  assign _zz_1923 = ($signed(_zz_1925) - $signed(_zz_6011));
  assign _zz_1924 = ($signed(_zz_1925) + $signed(_zz_6013));
  assign _zz_1926 = 1'b1;
  assign _zz_1927 = 1'b1;
  assign _zz_4120 = ($signed(_zz_6031) * $signed(_zz_111));
  assign _zz_1930 = _zz_6032[15 : 0];
  assign _zz_4121 = ($signed(_zz_6033) * $signed(twiddle_factor_table_0_real));
  assign _zz_4122 = ($signed(_zz_6034) * $signed(twiddle_factor_table_0_imag));
  assign _zz_1928 = ($signed(_zz_1930) - $signed(_zz_6035));
  assign _zz_1929 = ($signed(_zz_1930) + $signed(_zz_6037));
  assign _zz_1931 = 1'b1;
  assign _zz_1932 = 1'b1;
  assign _zz_4123 = ($signed(_zz_6055) * $signed(_zz_115));
  assign _zz_1935 = _zz_6056[15 : 0];
  assign _zz_4124 = ($signed(_zz_6057) * $signed(twiddle_factor_table_0_real));
  assign _zz_4125 = ($signed(_zz_6058) * $signed(twiddle_factor_table_0_imag));
  assign _zz_1933 = ($signed(_zz_1935) - $signed(_zz_6059));
  assign _zz_1934 = ($signed(_zz_1935) + $signed(_zz_6061));
  assign _zz_1936 = 1'b1;
  assign _zz_1937 = 1'b1;
  assign _zz_4126 = ($signed(_zz_6079) * $signed(_zz_119));
  assign _zz_1940 = _zz_6080[15 : 0];
  assign _zz_4127 = ($signed(_zz_6081) * $signed(twiddle_factor_table_0_real));
  assign _zz_4128 = ($signed(_zz_6082) * $signed(twiddle_factor_table_0_imag));
  assign _zz_1938 = ($signed(_zz_1940) - $signed(_zz_6083));
  assign _zz_1939 = ($signed(_zz_1940) + $signed(_zz_6085));
  assign _zz_1941 = 1'b1;
  assign _zz_1942 = 1'b1;
  assign _zz_4129 = ($signed(_zz_6103) * $signed(_zz_123));
  assign _zz_1945 = _zz_6104[15 : 0];
  assign _zz_4130 = ($signed(_zz_6105) * $signed(twiddle_factor_table_0_real));
  assign _zz_4131 = ($signed(_zz_6106) * $signed(twiddle_factor_table_0_imag));
  assign _zz_1943 = ($signed(_zz_1945) - $signed(_zz_6107));
  assign _zz_1944 = ($signed(_zz_1945) + $signed(_zz_6109));
  assign _zz_1946 = 1'b1;
  assign _zz_1947 = 1'b1;
  assign _zz_4132 = ($signed(_zz_6127) * $signed(_zz_127));
  assign _zz_1950 = _zz_6128[15 : 0];
  assign _zz_4133 = ($signed(_zz_6129) * $signed(twiddle_factor_table_0_real));
  assign _zz_4134 = ($signed(_zz_6130) * $signed(twiddle_factor_table_0_imag));
  assign _zz_1948 = ($signed(_zz_1950) - $signed(_zz_6131));
  assign _zz_1949 = ($signed(_zz_1950) + $signed(_zz_6133));
  assign _zz_1951 = 1'b1;
  assign _zz_1952 = 1'b1;
  assign _zz_4135 = ($signed(_zz_6151) * $signed(_zz_131));
  assign _zz_1955 = _zz_6152[15 : 0];
  assign _zz_4136 = ($signed(_zz_6153) * $signed(twiddle_factor_table_0_real));
  assign _zz_4137 = ($signed(_zz_6154) * $signed(twiddle_factor_table_0_imag));
  assign _zz_1953 = ($signed(_zz_1955) - $signed(_zz_6155));
  assign _zz_1954 = ($signed(_zz_1955) + $signed(_zz_6157));
  assign _zz_1956 = 1'b1;
  assign _zz_1957 = 1'b1;
  assign _zz_4138 = ($signed(_zz_6175) * $signed(_zz_135));
  assign _zz_1960 = _zz_6176[15 : 0];
  assign _zz_4139 = ($signed(_zz_6177) * $signed(twiddle_factor_table_0_real));
  assign _zz_4140 = ($signed(_zz_6178) * $signed(twiddle_factor_table_0_imag));
  assign _zz_1958 = ($signed(_zz_1960) - $signed(_zz_6179));
  assign _zz_1959 = ($signed(_zz_1960) + $signed(_zz_6181));
  assign _zz_1961 = 1'b1;
  assign _zz_1962 = 1'b1;
  assign _zz_4141 = ($signed(_zz_6199) * $signed(_zz_139));
  assign _zz_1965 = _zz_6200[15 : 0];
  assign _zz_4142 = ($signed(_zz_6201) * $signed(twiddle_factor_table_0_real));
  assign _zz_4143 = ($signed(_zz_6202) * $signed(twiddle_factor_table_0_imag));
  assign _zz_1963 = ($signed(_zz_1965) - $signed(_zz_6203));
  assign _zz_1964 = ($signed(_zz_1965) + $signed(_zz_6205));
  assign _zz_1966 = 1'b1;
  assign _zz_1967 = 1'b1;
  assign _zz_4144 = ($signed(_zz_6223) * $signed(_zz_143));
  assign _zz_1970 = _zz_6224[15 : 0];
  assign _zz_4145 = ($signed(_zz_6225) * $signed(twiddle_factor_table_0_real));
  assign _zz_4146 = ($signed(_zz_6226) * $signed(twiddle_factor_table_0_imag));
  assign _zz_1968 = ($signed(_zz_1970) - $signed(_zz_6227));
  assign _zz_1969 = ($signed(_zz_1970) + $signed(_zz_6229));
  assign _zz_1971 = 1'b1;
  assign _zz_1972 = 1'b1;
  assign _zz_4147 = ($signed(_zz_6247) * $signed(_zz_147));
  assign _zz_1975 = _zz_6248[15 : 0];
  assign _zz_4148 = ($signed(_zz_6249) * $signed(twiddle_factor_table_0_real));
  assign _zz_4149 = ($signed(_zz_6250) * $signed(twiddle_factor_table_0_imag));
  assign _zz_1973 = ($signed(_zz_1975) - $signed(_zz_6251));
  assign _zz_1974 = ($signed(_zz_1975) + $signed(_zz_6253));
  assign _zz_1976 = 1'b1;
  assign _zz_1977 = 1'b1;
  assign _zz_4150 = ($signed(_zz_6271) * $signed(_zz_151));
  assign _zz_1980 = _zz_6272[15 : 0];
  assign _zz_4151 = ($signed(_zz_6273) * $signed(twiddle_factor_table_0_real));
  assign _zz_4152 = ($signed(_zz_6274) * $signed(twiddle_factor_table_0_imag));
  assign _zz_1978 = ($signed(_zz_1980) - $signed(_zz_6275));
  assign _zz_1979 = ($signed(_zz_1980) + $signed(_zz_6277));
  assign _zz_1981 = 1'b1;
  assign _zz_1982 = 1'b1;
  assign _zz_4153 = ($signed(_zz_6295) * $signed(_zz_155));
  assign _zz_1985 = _zz_6296[15 : 0];
  assign _zz_4154 = ($signed(_zz_6297) * $signed(twiddle_factor_table_0_real));
  assign _zz_4155 = ($signed(_zz_6298) * $signed(twiddle_factor_table_0_imag));
  assign _zz_1983 = ($signed(_zz_1985) - $signed(_zz_6299));
  assign _zz_1984 = ($signed(_zz_1985) + $signed(_zz_6301));
  assign _zz_1986 = 1'b1;
  assign _zz_1987 = 1'b1;
  assign _zz_4156 = ($signed(_zz_6319) * $signed(_zz_159));
  assign _zz_1990 = _zz_6320[15 : 0];
  assign _zz_4157 = ($signed(_zz_6321) * $signed(twiddle_factor_table_0_real));
  assign _zz_4158 = ($signed(_zz_6322) * $signed(twiddle_factor_table_0_imag));
  assign _zz_1988 = ($signed(_zz_1990) - $signed(_zz_6323));
  assign _zz_1989 = ($signed(_zz_1990) + $signed(_zz_6325));
  assign _zz_1991 = 1'b1;
  assign _zz_1992 = 1'b1;
  assign _zz_4159 = ($signed(_zz_6343) * $signed(_zz_163));
  assign _zz_1995 = _zz_6344[15 : 0];
  assign _zz_4160 = ($signed(_zz_6345) * $signed(twiddle_factor_table_0_real));
  assign _zz_4161 = ($signed(_zz_6346) * $signed(twiddle_factor_table_0_imag));
  assign _zz_1993 = ($signed(_zz_1995) - $signed(_zz_6347));
  assign _zz_1994 = ($signed(_zz_1995) + $signed(_zz_6349));
  assign _zz_1996 = 1'b1;
  assign _zz_1997 = 1'b1;
  assign _zz_4162 = ($signed(_zz_6367) * $signed(_zz_167));
  assign _zz_2000 = _zz_6368[15 : 0];
  assign _zz_4163 = ($signed(_zz_6369) * $signed(twiddle_factor_table_0_real));
  assign _zz_4164 = ($signed(_zz_6370) * $signed(twiddle_factor_table_0_imag));
  assign _zz_1998 = ($signed(_zz_2000) - $signed(_zz_6371));
  assign _zz_1999 = ($signed(_zz_2000) + $signed(_zz_6373));
  assign _zz_2001 = 1'b1;
  assign _zz_2002 = 1'b1;
  assign _zz_4165 = ($signed(_zz_6391) * $signed(_zz_171));
  assign _zz_2005 = _zz_6392[15 : 0];
  assign _zz_4166 = ($signed(_zz_6393) * $signed(twiddle_factor_table_0_real));
  assign _zz_4167 = ($signed(_zz_6394) * $signed(twiddle_factor_table_0_imag));
  assign _zz_2003 = ($signed(_zz_2005) - $signed(_zz_6395));
  assign _zz_2004 = ($signed(_zz_2005) + $signed(_zz_6397));
  assign _zz_2006 = 1'b1;
  assign _zz_2007 = 1'b1;
  assign _zz_4168 = ($signed(_zz_6415) * $signed(_zz_175));
  assign _zz_2010 = _zz_6416[15 : 0];
  assign _zz_4169 = ($signed(_zz_6417) * $signed(twiddle_factor_table_0_real));
  assign _zz_4170 = ($signed(_zz_6418) * $signed(twiddle_factor_table_0_imag));
  assign _zz_2008 = ($signed(_zz_2010) - $signed(_zz_6419));
  assign _zz_2009 = ($signed(_zz_2010) + $signed(_zz_6421));
  assign _zz_2011 = 1'b1;
  assign _zz_2012 = 1'b1;
  assign _zz_4171 = ($signed(_zz_6439) * $signed(_zz_179));
  assign _zz_2015 = _zz_6440[15 : 0];
  assign _zz_4172 = ($signed(_zz_6441) * $signed(twiddle_factor_table_0_real));
  assign _zz_4173 = ($signed(_zz_6442) * $signed(twiddle_factor_table_0_imag));
  assign _zz_2013 = ($signed(_zz_2015) - $signed(_zz_6443));
  assign _zz_2014 = ($signed(_zz_2015) + $signed(_zz_6445));
  assign _zz_2016 = 1'b1;
  assign _zz_2017 = 1'b1;
  assign _zz_4174 = ($signed(_zz_6463) * $signed(_zz_183));
  assign _zz_2020 = _zz_6464[15 : 0];
  assign _zz_4175 = ($signed(_zz_6465) * $signed(twiddle_factor_table_0_real));
  assign _zz_4176 = ($signed(_zz_6466) * $signed(twiddle_factor_table_0_imag));
  assign _zz_2018 = ($signed(_zz_2020) - $signed(_zz_6467));
  assign _zz_2019 = ($signed(_zz_2020) + $signed(_zz_6469));
  assign _zz_2021 = 1'b1;
  assign _zz_2022 = 1'b1;
  assign _zz_4177 = ($signed(_zz_6487) * $signed(_zz_187));
  assign _zz_2025 = _zz_6488[15 : 0];
  assign _zz_4178 = ($signed(_zz_6489) * $signed(twiddle_factor_table_0_real));
  assign _zz_4179 = ($signed(_zz_6490) * $signed(twiddle_factor_table_0_imag));
  assign _zz_2023 = ($signed(_zz_2025) - $signed(_zz_6491));
  assign _zz_2024 = ($signed(_zz_2025) + $signed(_zz_6493));
  assign _zz_2026 = 1'b1;
  assign _zz_2027 = 1'b1;
  assign _zz_4180 = ($signed(_zz_6511) * $signed(_zz_191));
  assign _zz_2030 = _zz_6512[15 : 0];
  assign _zz_4181 = ($signed(_zz_6513) * $signed(twiddle_factor_table_0_real));
  assign _zz_4182 = ($signed(_zz_6514) * $signed(twiddle_factor_table_0_imag));
  assign _zz_2028 = ($signed(_zz_2030) - $signed(_zz_6515));
  assign _zz_2029 = ($signed(_zz_2030) + $signed(_zz_6517));
  assign _zz_2031 = 1'b1;
  assign _zz_2032 = 1'b1;
  assign _zz_4183 = ($signed(_zz_6535) * $signed(_zz_195));
  assign _zz_2035 = _zz_6536[15 : 0];
  assign _zz_4184 = ($signed(_zz_6537) * $signed(twiddle_factor_table_0_real));
  assign _zz_4185 = ($signed(_zz_6538) * $signed(twiddle_factor_table_0_imag));
  assign _zz_2033 = ($signed(_zz_2035) - $signed(_zz_6539));
  assign _zz_2034 = ($signed(_zz_2035) + $signed(_zz_6541));
  assign _zz_2036 = 1'b1;
  assign _zz_2037 = 1'b1;
  assign _zz_4186 = ($signed(_zz_6559) * $signed(_zz_199));
  assign _zz_2040 = _zz_6560[15 : 0];
  assign _zz_4187 = ($signed(_zz_6561) * $signed(twiddle_factor_table_0_real));
  assign _zz_4188 = ($signed(_zz_6562) * $signed(twiddle_factor_table_0_imag));
  assign _zz_2038 = ($signed(_zz_2040) - $signed(_zz_6563));
  assign _zz_2039 = ($signed(_zz_2040) + $signed(_zz_6565));
  assign _zz_2041 = 1'b1;
  assign _zz_2042 = 1'b1;
  assign _zz_4189 = ($signed(_zz_6583) * $signed(_zz_203));
  assign _zz_2045 = _zz_6584[15 : 0];
  assign _zz_4190 = ($signed(_zz_6585) * $signed(twiddle_factor_table_0_real));
  assign _zz_4191 = ($signed(_zz_6586) * $signed(twiddle_factor_table_0_imag));
  assign _zz_2043 = ($signed(_zz_2045) - $signed(_zz_6587));
  assign _zz_2044 = ($signed(_zz_2045) + $signed(_zz_6589));
  assign _zz_2046 = 1'b1;
  assign _zz_2047 = 1'b1;
  assign _zz_4192 = ($signed(_zz_6607) * $signed(_zz_207));
  assign _zz_2050 = _zz_6608[15 : 0];
  assign _zz_4193 = ($signed(_zz_6609) * $signed(twiddle_factor_table_0_real));
  assign _zz_4194 = ($signed(_zz_6610) * $signed(twiddle_factor_table_0_imag));
  assign _zz_2048 = ($signed(_zz_2050) - $signed(_zz_6611));
  assign _zz_2049 = ($signed(_zz_2050) + $signed(_zz_6613));
  assign _zz_2051 = 1'b1;
  assign _zz_2052 = 1'b1;
  assign _zz_4195 = ($signed(_zz_6631) * $signed(_zz_211));
  assign _zz_2055 = _zz_6632[15 : 0];
  assign _zz_4196 = ($signed(_zz_6633) * $signed(twiddle_factor_table_0_real));
  assign _zz_4197 = ($signed(_zz_6634) * $signed(twiddle_factor_table_0_imag));
  assign _zz_2053 = ($signed(_zz_2055) - $signed(_zz_6635));
  assign _zz_2054 = ($signed(_zz_2055) + $signed(_zz_6637));
  assign _zz_2056 = 1'b1;
  assign _zz_2057 = 1'b1;
  assign _zz_4198 = ($signed(_zz_6655) * $signed(_zz_215));
  assign _zz_2060 = _zz_6656[15 : 0];
  assign _zz_4199 = ($signed(_zz_6657) * $signed(twiddle_factor_table_0_real));
  assign _zz_4200 = ($signed(_zz_6658) * $signed(twiddle_factor_table_0_imag));
  assign _zz_2058 = ($signed(_zz_2060) - $signed(_zz_6659));
  assign _zz_2059 = ($signed(_zz_2060) + $signed(_zz_6661));
  assign _zz_2061 = 1'b1;
  assign _zz_2062 = 1'b1;
  assign _zz_4201 = ($signed(_zz_6679) * $signed(_zz_219));
  assign _zz_2065 = _zz_6680[15 : 0];
  assign _zz_4202 = ($signed(_zz_6681) * $signed(twiddle_factor_table_0_real));
  assign _zz_4203 = ($signed(_zz_6682) * $signed(twiddle_factor_table_0_imag));
  assign _zz_2063 = ($signed(_zz_2065) - $signed(_zz_6683));
  assign _zz_2064 = ($signed(_zz_2065) + $signed(_zz_6685));
  assign _zz_2066 = 1'b1;
  assign _zz_2067 = 1'b1;
  assign _zz_4204 = ($signed(_zz_6703) * $signed(_zz_223));
  assign _zz_2070 = _zz_6704[15 : 0];
  assign _zz_4205 = ($signed(_zz_6705) * $signed(twiddle_factor_table_0_real));
  assign _zz_4206 = ($signed(_zz_6706) * $signed(twiddle_factor_table_0_imag));
  assign _zz_2068 = ($signed(_zz_2070) - $signed(_zz_6707));
  assign _zz_2069 = ($signed(_zz_2070) + $signed(_zz_6709));
  assign _zz_2071 = 1'b1;
  assign _zz_2072 = 1'b1;
  assign _zz_4207 = ($signed(_zz_6727) * $signed(_zz_227));
  assign _zz_2075 = _zz_6728[15 : 0];
  assign _zz_4208 = ($signed(_zz_6729) * $signed(twiddle_factor_table_0_real));
  assign _zz_4209 = ($signed(_zz_6730) * $signed(twiddle_factor_table_0_imag));
  assign _zz_2073 = ($signed(_zz_2075) - $signed(_zz_6731));
  assign _zz_2074 = ($signed(_zz_2075) + $signed(_zz_6733));
  assign _zz_2076 = 1'b1;
  assign _zz_2077 = 1'b1;
  assign _zz_4210 = ($signed(_zz_6751) * $signed(_zz_231));
  assign _zz_2080 = _zz_6752[15 : 0];
  assign _zz_4211 = ($signed(_zz_6753) * $signed(twiddle_factor_table_0_real));
  assign _zz_4212 = ($signed(_zz_6754) * $signed(twiddle_factor_table_0_imag));
  assign _zz_2078 = ($signed(_zz_2080) - $signed(_zz_6755));
  assign _zz_2079 = ($signed(_zz_2080) + $signed(_zz_6757));
  assign _zz_2081 = 1'b1;
  assign _zz_2082 = 1'b1;
  assign _zz_4213 = ($signed(_zz_6775) * $signed(_zz_235));
  assign _zz_2085 = _zz_6776[15 : 0];
  assign _zz_4214 = ($signed(_zz_6777) * $signed(twiddle_factor_table_0_real));
  assign _zz_4215 = ($signed(_zz_6778) * $signed(twiddle_factor_table_0_imag));
  assign _zz_2083 = ($signed(_zz_2085) - $signed(_zz_6779));
  assign _zz_2084 = ($signed(_zz_2085) + $signed(_zz_6781));
  assign _zz_2086 = 1'b1;
  assign _zz_2087 = 1'b1;
  assign _zz_4216 = ($signed(_zz_6799) * $signed(_zz_239));
  assign _zz_2090 = _zz_6800[15 : 0];
  assign _zz_4217 = ($signed(_zz_6801) * $signed(twiddle_factor_table_0_real));
  assign _zz_4218 = ($signed(_zz_6802) * $signed(twiddle_factor_table_0_imag));
  assign _zz_2088 = ($signed(_zz_2090) - $signed(_zz_6803));
  assign _zz_2089 = ($signed(_zz_2090) + $signed(_zz_6805));
  assign _zz_2091 = 1'b1;
  assign _zz_2092 = 1'b1;
  assign _zz_4219 = ($signed(_zz_6823) * $signed(_zz_243));
  assign _zz_2095 = _zz_6824[15 : 0];
  assign _zz_4220 = ($signed(_zz_6825) * $signed(twiddle_factor_table_0_real));
  assign _zz_4221 = ($signed(_zz_6826) * $signed(twiddle_factor_table_0_imag));
  assign _zz_2093 = ($signed(_zz_2095) - $signed(_zz_6827));
  assign _zz_2094 = ($signed(_zz_2095) + $signed(_zz_6829));
  assign _zz_2096 = 1'b1;
  assign _zz_2097 = 1'b1;
  assign _zz_4222 = ($signed(_zz_6847) * $signed(_zz_247));
  assign _zz_2100 = _zz_6848[15 : 0];
  assign _zz_4223 = ($signed(_zz_6849) * $signed(twiddle_factor_table_0_real));
  assign _zz_4224 = ($signed(_zz_6850) * $signed(twiddle_factor_table_0_imag));
  assign _zz_2098 = ($signed(_zz_2100) - $signed(_zz_6851));
  assign _zz_2099 = ($signed(_zz_2100) + $signed(_zz_6853));
  assign _zz_2101 = 1'b1;
  assign _zz_2102 = 1'b1;
  assign _zz_4225 = ($signed(_zz_6871) * $signed(_zz_251));
  assign _zz_2105 = _zz_6872[15 : 0];
  assign _zz_4226 = ($signed(_zz_6873) * $signed(twiddle_factor_table_0_real));
  assign _zz_4227 = ($signed(_zz_6874) * $signed(twiddle_factor_table_0_imag));
  assign _zz_2103 = ($signed(_zz_2105) - $signed(_zz_6875));
  assign _zz_2104 = ($signed(_zz_2105) + $signed(_zz_6877));
  assign _zz_2106 = 1'b1;
  assign _zz_2107 = 1'b1;
  assign _zz_4228 = ($signed(_zz_6895) * $signed(_zz_255));
  assign _zz_2110 = _zz_6896[15 : 0];
  assign _zz_4229 = ($signed(_zz_6897) * $signed(twiddle_factor_table_0_real));
  assign _zz_4230 = ($signed(_zz_6898) * $signed(twiddle_factor_table_0_imag));
  assign _zz_2108 = ($signed(_zz_2110) - $signed(_zz_6899));
  assign _zz_2109 = ($signed(_zz_2110) + $signed(_zz_6901));
  assign _zz_2111 = 1'b1;
  assign _zz_2112 = 1'b1;
  assign _zz_4231 = ($signed(_zz_6919) * $signed(_zz_261));
  assign _zz_2115 = _zz_6920[15 : 0];
  assign _zz_4232 = ($signed(_zz_6921) * $signed(twiddle_factor_table_1_real));
  assign _zz_4233 = ($signed(_zz_6922) * $signed(twiddle_factor_table_1_imag));
  assign _zz_2113 = ($signed(_zz_2115) - $signed(_zz_6923));
  assign _zz_2114 = ($signed(_zz_2115) + $signed(_zz_6925));
  assign _zz_2116 = 1'b1;
  assign _zz_2117 = 1'b1;
  assign _zz_4234 = ($signed(_zz_6943) * $signed(_zz_263));
  assign _zz_2120 = _zz_6944[15 : 0];
  assign _zz_4235 = ($signed(_zz_6945) * $signed(twiddle_factor_table_2_real));
  assign _zz_4236 = ($signed(_zz_6946) * $signed(twiddle_factor_table_2_imag));
  assign _zz_2118 = ($signed(_zz_2120) - $signed(_zz_6947));
  assign _zz_2119 = ($signed(_zz_2120) + $signed(_zz_6949));
  assign _zz_2121 = 1'b1;
  assign _zz_2122 = 1'b1;
  assign _zz_4237 = ($signed(_zz_6967) * $signed(_zz_269));
  assign _zz_2125 = _zz_6968[15 : 0];
  assign _zz_4238 = ($signed(_zz_6969) * $signed(twiddle_factor_table_1_real));
  assign _zz_4239 = ($signed(_zz_6970) * $signed(twiddle_factor_table_1_imag));
  assign _zz_2123 = ($signed(_zz_2125) - $signed(_zz_6971));
  assign _zz_2124 = ($signed(_zz_2125) + $signed(_zz_6973));
  assign _zz_2126 = 1'b1;
  assign _zz_2127 = 1'b1;
  assign _zz_4240 = ($signed(_zz_6991) * $signed(_zz_271));
  assign _zz_2130 = _zz_6992[15 : 0];
  assign _zz_4241 = ($signed(_zz_6993) * $signed(twiddle_factor_table_2_real));
  assign _zz_4242 = ($signed(_zz_6994) * $signed(twiddle_factor_table_2_imag));
  assign _zz_2128 = ($signed(_zz_2130) - $signed(_zz_6995));
  assign _zz_2129 = ($signed(_zz_2130) + $signed(_zz_6997));
  assign _zz_2131 = 1'b1;
  assign _zz_2132 = 1'b1;
  assign _zz_4243 = ($signed(_zz_7015) * $signed(_zz_277));
  assign _zz_2135 = _zz_7016[15 : 0];
  assign _zz_4244 = ($signed(_zz_7017) * $signed(twiddle_factor_table_1_real));
  assign _zz_4245 = ($signed(_zz_7018) * $signed(twiddle_factor_table_1_imag));
  assign _zz_2133 = ($signed(_zz_2135) - $signed(_zz_7019));
  assign _zz_2134 = ($signed(_zz_2135) + $signed(_zz_7021));
  assign _zz_2136 = 1'b1;
  assign _zz_2137 = 1'b1;
  assign _zz_4246 = ($signed(_zz_7039) * $signed(_zz_279));
  assign _zz_2140 = _zz_7040[15 : 0];
  assign _zz_4247 = ($signed(_zz_7041) * $signed(twiddle_factor_table_2_real));
  assign _zz_4248 = ($signed(_zz_7042) * $signed(twiddle_factor_table_2_imag));
  assign _zz_2138 = ($signed(_zz_2140) - $signed(_zz_7043));
  assign _zz_2139 = ($signed(_zz_2140) + $signed(_zz_7045));
  assign _zz_2141 = 1'b1;
  assign _zz_2142 = 1'b1;
  assign _zz_4249 = ($signed(_zz_7063) * $signed(_zz_285));
  assign _zz_2145 = _zz_7064[15 : 0];
  assign _zz_4250 = ($signed(_zz_7065) * $signed(twiddle_factor_table_1_real));
  assign _zz_4251 = ($signed(_zz_7066) * $signed(twiddle_factor_table_1_imag));
  assign _zz_2143 = ($signed(_zz_2145) - $signed(_zz_7067));
  assign _zz_2144 = ($signed(_zz_2145) + $signed(_zz_7069));
  assign _zz_2146 = 1'b1;
  assign _zz_2147 = 1'b1;
  assign _zz_4252 = ($signed(_zz_7087) * $signed(_zz_287));
  assign _zz_2150 = _zz_7088[15 : 0];
  assign _zz_4253 = ($signed(_zz_7089) * $signed(twiddle_factor_table_2_real));
  assign _zz_4254 = ($signed(_zz_7090) * $signed(twiddle_factor_table_2_imag));
  assign _zz_2148 = ($signed(_zz_2150) - $signed(_zz_7091));
  assign _zz_2149 = ($signed(_zz_2150) + $signed(_zz_7093));
  assign _zz_2151 = 1'b1;
  assign _zz_2152 = 1'b1;
  assign _zz_4255 = ($signed(_zz_7111) * $signed(_zz_293));
  assign _zz_2155 = _zz_7112[15 : 0];
  assign _zz_4256 = ($signed(_zz_7113) * $signed(twiddle_factor_table_1_real));
  assign _zz_4257 = ($signed(_zz_7114) * $signed(twiddle_factor_table_1_imag));
  assign _zz_2153 = ($signed(_zz_2155) - $signed(_zz_7115));
  assign _zz_2154 = ($signed(_zz_2155) + $signed(_zz_7117));
  assign _zz_2156 = 1'b1;
  assign _zz_2157 = 1'b1;
  assign _zz_4258 = ($signed(_zz_7135) * $signed(_zz_295));
  assign _zz_2160 = _zz_7136[15 : 0];
  assign _zz_4259 = ($signed(_zz_7137) * $signed(twiddle_factor_table_2_real));
  assign _zz_4260 = ($signed(_zz_7138) * $signed(twiddle_factor_table_2_imag));
  assign _zz_2158 = ($signed(_zz_2160) - $signed(_zz_7139));
  assign _zz_2159 = ($signed(_zz_2160) + $signed(_zz_7141));
  assign _zz_2161 = 1'b1;
  assign _zz_2162 = 1'b1;
  assign _zz_4261 = ($signed(_zz_7159) * $signed(_zz_301));
  assign _zz_2165 = _zz_7160[15 : 0];
  assign _zz_4262 = ($signed(_zz_7161) * $signed(twiddle_factor_table_1_real));
  assign _zz_4263 = ($signed(_zz_7162) * $signed(twiddle_factor_table_1_imag));
  assign _zz_2163 = ($signed(_zz_2165) - $signed(_zz_7163));
  assign _zz_2164 = ($signed(_zz_2165) + $signed(_zz_7165));
  assign _zz_2166 = 1'b1;
  assign _zz_2167 = 1'b1;
  assign _zz_4264 = ($signed(_zz_7183) * $signed(_zz_303));
  assign _zz_2170 = _zz_7184[15 : 0];
  assign _zz_4265 = ($signed(_zz_7185) * $signed(twiddle_factor_table_2_real));
  assign _zz_4266 = ($signed(_zz_7186) * $signed(twiddle_factor_table_2_imag));
  assign _zz_2168 = ($signed(_zz_2170) - $signed(_zz_7187));
  assign _zz_2169 = ($signed(_zz_2170) + $signed(_zz_7189));
  assign _zz_2171 = 1'b1;
  assign _zz_2172 = 1'b1;
  assign _zz_4267 = ($signed(_zz_7207) * $signed(_zz_309));
  assign _zz_2175 = _zz_7208[15 : 0];
  assign _zz_4268 = ($signed(_zz_7209) * $signed(twiddle_factor_table_1_real));
  assign _zz_4269 = ($signed(_zz_7210) * $signed(twiddle_factor_table_1_imag));
  assign _zz_2173 = ($signed(_zz_2175) - $signed(_zz_7211));
  assign _zz_2174 = ($signed(_zz_2175) + $signed(_zz_7213));
  assign _zz_2176 = 1'b1;
  assign _zz_2177 = 1'b1;
  assign _zz_4270 = ($signed(_zz_7231) * $signed(_zz_311));
  assign _zz_2180 = _zz_7232[15 : 0];
  assign _zz_4271 = ($signed(_zz_7233) * $signed(twiddle_factor_table_2_real));
  assign _zz_4272 = ($signed(_zz_7234) * $signed(twiddle_factor_table_2_imag));
  assign _zz_2178 = ($signed(_zz_2180) - $signed(_zz_7235));
  assign _zz_2179 = ($signed(_zz_2180) + $signed(_zz_7237));
  assign _zz_2181 = 1'b1;
  assign _zz_2182 = 1'b1;
  assign _zz_4273 = ($signed(_zz_7255) * $signed(_zz_317));
  assign _zz_2185 = _zz_7256[15 : 0];
  assign _zz_4274 = ($signed(_zz_7257) * $signed(twiddle_factor_table_1_real));
  assign _zz_4275 = ($signed(_zz_7258) * $signed(twiddle_factor_table_1_imag));
  assign _zz_2183 = ($signed(_zz_2185) - $signed(_zz_7259));
  assign _zz_2184 = ($signed(_zz_2185) + $signed(_zz_7261));
  assign _zz_2186 = 1'b1;
  assign _zz_2187 = 1'b1;
  assign _zz_4276 = ($signed(_zz_7279) * $signed(_zz_319));
  assign _zz_2190 = _zz_7280[15 : 0];
  assign _zz_4277 = ($signed(_zz_7281) * $signed(twiddle_factor_table_2_real));
  assign _zz_4278 = ($signed(_zz_7282) * $signed(twiddle_factor_table_2_imag));
  assign _zz_2188 = ($signed(_zz_2190) - $signed(_zz_7283));
  assign _zz_2189 = ($signed(_zz_2190) + $signed(_zz_7285));
  assign _zz_2191 = 1'b1;
  assign _zz_2192 = 1'b1;
  assign _zz_4279 = ($signed(_zz_7303) * $signed(_zz_325));
  assign _zz_2195 = _zz_7304[15 : 0];
  assign _zz_4280 = ($signed(_zz_7305) * $signed(twiddle_factor_table_1_real));
  assign _zz_4281 = ($signed(_zz_7306) * $signed(twiddle_factor_table_1_imag));
  assign _zz_2193 = ($signed(_zz_2195) - $signed(_zz_7307));
  assign _zz_2194 = ($signed(_zz_2195) + $signed(_zz_7309));
  assign _zz_2196 = 1'b1;
  assign _zz_2197 = 1'b1;
  assign _zz_4282 = ($signed(_zz_7327) * $signed(_zz_327));
  assign _zz_2200 = _zz_7328[15 : 0];
  assign _zz_4283 = ($signed(_zz_7329) * $signed(twiddle_factor_table_2_real));
  assign _zz_4284 = ($signed(_zz_7330) * $signed(twiddle_factor_table_2_imag));
  assign _zz_2198 = ($signed(_zz_2200) - $signed(_zz_7331));
  assign _zz_2199 = ($signed(_zz_2200) + $signed(_zz_7333));
  assign _zz_2201 = 1'b1;
  assign _zz_2202 = 1'b1;
  assign _zz_4285 = ($signed(_zz_7351) * $signed(_zz_333));
  assign _zz_2205 = _zz_7352[15 : 0];
  assign _zz_4286 = ($signed(_zz_7353) * $signed(twiddle_factor_table_1_real));
  assign _zz_4287 = ($signed(_zz_7354) * $signed(twiddle_factor_table_1_imag));
  assign _zz_2203 = ($signed(_zz_2205) - $signed(_zz_7355));
  assign _zz_2204 = ($signed(_zz_2205) + $signed(_zz_7357));
  assign _zz_2206 = 1'b1;
  assign _zz_2207 = 1'b1;
  assign _zz_4288 = ($signed(_zz_7375) * $signed(_zz_335));
  assign _zz_2210 = _zz_7376[15 : 0];
  assign _zz_4289 = ($signed(_zz_7377) * $signed(twiddle_factor_table_2_real));
  assign _zz_4290 = ($signed(_zz_7378) * $signed(twiddle_factor_table_2_imag));
  assign _zz_2208 = ($signed(_zz_2210) - $signed(_zz_7379));
  assign _zz_2209 = ($signed(_zz_2210) + $signed(_zz_7381));
  assign _zz_2211 = 1'b1;
  assign _zz_2212 = 1'b1;
  assign _zz_4291 = ($signed(_zz_7399) * $signed(_zz_341));
  assign _zz_2215 = _zz_7400[15 : 0];
  assign _zz_4292 = ($signed(_zz_7401) * $signed(twiddle_factor_table_1_real));
  assign _zz_4293 = ($signed(_zz_7402) * $signed(twiddle_factor_table_1_imag));
  assign _zz_2213 = ($signed(_zz_2215) - $signed(_zz_7403));
  assign _zz_2214 = ($signed(_zz_2215) + $signed(_zz_7405));
  assign _zz_2216 = 1'b1;
  assign _zz_2217 = 1'b1;
  assign _zz_4294 = ($signed(_zz_7423) * $signed(_zz_343));
  assign _zz_2220 = _zz_7424[15 : 0];
  assign _zz_4295 = ($signed(_zz_7425) * $signed(twiddle_factor_table_2_real));
  assign _zz_4296 = ($signed(_zz_7426) * $signed(twiddle_factor_table_2_imag));
  assign _zz_2218 = ($signed(_zz_2220) - $signed(_zz_7427));
  assign _zz_2219 = ($signed(_zz_2220) + $signed(_zz_7429));
  assign _zz_2221 = 1'b1;
  assign _zz_2222 = 1'b1;
  assign _zz_4297 = ($signed(_zz_7447) * $signed(_zz_349));
  assign _zz_2225 = _zz_7448[15 : 0];
  assign _zz_4298 = ($signed(_zz_7449) * $signed(twiddle_factor_table_1_real));
  assign _zz_4299 = ($signed(_zz_7450) * $signed(twiddle_factor_table_1_imag));
  assign _zz_2223 = ($signed(_zz_2225) - $signed(_zz_7451));
  assign _zz_2224 = ($signed(_zz_2225) + $signed(_zz_7453));
  assign _zz_2226 = 1'b1;
  assign _zz_2227 = 1'b1;
  assign _zz_4300 = ($signed(_zz_7471) * $signed(_zz_351));
  assign _zz_2230 = _zz_7472[15 : 0];
  assign _zz_4301 = ($signed(_zz_7473) * $signed(twiddle_factor_table_2_real));
  assign _zz_4302 = ($signed(_zz_7474) * $signed(twiddle_factor_table_2_imag));
  assign _zz_2228 = ($signed(_zz_2230) - $signed(_zz_7475));
  assign _zz_2229 = ($signed(_zz_2230) + $signed(_zz_7477));
  assign _zz_2231 = 1'b1;
  assign _zz_2232 = 1'b1;
  assign _zz_4303 = ($signed(_zz_7495) * $signed(_zz_357));
  assign _zz_2235 = _zz_7496[15 : 0];
  assign _zz_4304 = ($signed(_zz_7497) * $signed(twiddle_factor_table_1_real));
  assign _zz_4305 = ($signed(_zz_7498) * $signed(twiddle_factor_table_1_imag));
  assign _zz_2233 = ($signed(_zz_2235) - $signed(_zz_7499));
  assign _zz_2234 = ($signed(_zz_2235) + $signed(_zz_7501));
  assign _zz_2236 = 1'b1;
  assign _zz_2237 = 1'b1;
  assign _zz_4306 = ($signed(_zz_7519) * $signed(_zz_359));
  assign _zz_2240 = _zz_7520[15 : 0];
  assign _zz_4307 = ($signed(_zz_7521) * $signed(twiddle_factor_table_2_real));
  assign _zz_4308 = ($signed(_zz_7522) * $signed(twiddle_factor_table_2_imag));
  assign _zz_2238 = ($signed(_zz_2240) - $signed(_zz_7523));
  assign _zz_2239 = ($signed(_zz_2240) + $signed(_zz_7525));
  assign _zz_2241 = 1'b1;
  assign _zz_2242 = 1'b1;
  assign _zz_4309 = ($signed(_zz_7543) * $signed(_zz_365));
  assign _zz_2245 = _zz_7544[15 : 0];
  assign _zz_4310 = ($signed(_zz_7545) * $signed(twiddle_factor_table_1_real));
  assign _zz_4311 = ($signed(_zz_7546) * $signed(twiddle_factor_table_1_imag));
  assign _zz_2243 = ($signed(_zz_2245) - $signed(_zz_7547));
  assign _zz_2244 = ($signed(_zz_2245) + $signed(_zz_7549));
  assign _zz_2246 = 1'b1;
  assign _zz_2247 = 1'b1;
  assign _zz_4312 = ($signed(_zz_7567) * $signed(_zz_367));
  assign _zz_2250 = _zz_7568[15 : 0];
  assign _zz_4313 = ($signed(_zz_7569) * $signed(twiddle_factor_table_2_real));
  assign _zz_4314 = ($signed(_zz_7570) * $signed(twiddle_factor_table_2_imag));
  assign _zz_2248 = ($signed(_zz_2250) - $signed(_zz_7571));
  assign _zz_2249 = ($signed(_zz_2250) + $signed(_zz_7573));
  assign _zz_2251 = 1'b1;
  assign _zz_2252 = 1'b1;
  assign _zz_4315 = ($signed(_zz_7591) * $signed(_zz_373));
  assign _zz_2255 = _zz_7592[15 : 0];
  assign _zz_4316 = ($signed(_zz_7593) * $signed(twiddle_factor_table_1_real));
  assign _zz_4317 = ($signed(_zz_7594) * $signed(twiddle_factor_table_1_imag));
  assign _zz_2253 = ($signed(_zz_2255) - $signed(_zz_7595));
  assign _zz_2254 = ($signed(_zz_2255) + $signed(_zz_7597));
  assign _zz_2256 = 1'b1;
  assign _zz_2257 = 1'b1;
  assign _zz_4318 = ($signed(_zz_7615) * $signed(_zz_375));
  assign _zz_2260 = _zz_7616[15 : 0];
  assign _zz_4319 = ($signed(_zz_7617) * $signed(twiddle_factor_table_2_real));
  assign _zz_4320 = ($signed(_zz_7618) * $signed(twiddle_factor_table_2_imag));
  assign _zz_2258 = ($signed(_zz_2260) - $signed(_zz_7619));
  assign _zz_2259 = ($signed(_zz_2260) + $signed(_zz_7621));
  assign _zz_2261 = 1'b1;
  assign _zz_2262 = 1'b1;
  assign _zz_4321 = ($signed(_zz_7639) * $signed(_zz_381));
  assign _zz_2265 = _zz_7640[15 : 0];
  assign _zz_4322 = ($signed(_zz_7641) * $signed(twiddle_factor_table_1_real));
  assign _zz_4323 = ($signed(_zz_7642) * $signed(twiddle_factor_table_1_imag));
  assign _zz_2263 = ($signed(_zz_2265) - $signed(_zz_7643));
  assign _zz_2264 = ($signed(_zz_2265) + $signed(_zz_7645));
  assign _zz_2266 = 1'b1;
  assign _zz_2267 = 1'b1;
  assign _zz_4324 = ($signed(_zz_7663) * $signed(_zz_383));
  assign _zz_2270 = _zz_7664[15 : 0];
  assign _zz_4325 = ($signed(_zz_7665) * $signed(twiddle_factor_table_2_real));
  assign _zz_4326 = ($signed(_zz_7666) * $signed(twiddle_factor_table_2_imag));
  assign _zz_2268 = ($signed(_zz_2270) - $signed(_zz_7667));
  assign _zz_2269 = ($signed(_zz_2270) + $signed(_zz_7669));
  assign _zz_2271 = 1'b1;
  assign _zz_2272 = 1'b1;
  assign _zz_4327 = ($signed(_zz_7687) * $signed(_zz_389));
  assign _zz_2275 = _zz_7688[15 : 0];
  assign _zz_4328 = ($signed(_zz_7689) * $signed(twiddle_factor_table_1_real));
  assign _zz_4329 = ($signed(_zz_7690) * $signed(twiddle_factor_table_1_imag));
  assign _zz_2273 = ($signed(_zz_2275) - $signed(_zz_7691));
  assign _zz_2274 = ($signed(_zz_2275) + $signed(_zz_7693));
  assign _zz_2276 = 1'b1;
  assign _zz_2277 = 1'b1;
  assign _zz_4330 = ($signed(_zz_7711) * $signed(_zz_391));
  assign _zz_2280 = _zz_7712[15 : 0];
  assign _zz_4331 = ($signed(_zz_7713) * $signed(twiddle_factor_table_2_real));
  assign _zz_4332 = ($signed(_zz_7714) * $signed(twiddle_factor_table_2_imag));
  assign _zz_2278 = ($signed(_zz_2280) - $signed(_zz_7715));
  assign _zz_2279 = ($signed(_zz_2280) + $signed(_zz_7717));
  assign _zz_2281 = 1'b1;
  assign _zz_2282 = 1'b1;
  assign _zz_4333 = ($signed(_zz_7735) * $signed(_zz_397));
  assign _zz_2285 = _zz_7736[15 : 0];
  assign _zz_4334 = ($signed(_zz_7737) * $signed(twiddle_factor_table_1_real));
  assign _zz_4335 = ($signed(_zz_7738) * $signed(twiddle_factor_table_1_imag));
  assign _zz_2283 = ($signed(_zz_2285) - $signed(_zz_7739));
  assign _zz_2284 = ($signed(_zz_2285) + $signed(_zz_7741));
  assign _zz_2286 = 1'b1;
  assign _zz_2287 = 1'b1;
  assign _zz_4336 = ($signed(_zz_7759) * $signed(_zz_399));
  assign _zz_2290 = _zz_7760[15 : 0];
  assign _zz_4337 = ($signed(_zz_7761) * $signed(twiddle_factor_table_2_real));
  assign _zz_4338 = ($signed(_zz_7762) * $signed(twiddle_factor_table_2_imag));
  assign _zz_2288 = ($signed(_zz_2290) - $signed(_zz_7763));
  assign _zz_2289 = ($signed(_zz_2290) + $signed(_zz_7765));
  assign _zz_2291 = 1'b1;
  assign _zz_2292 = 1'b1;
  assign _zz_4339 = ($signed(_zz_7783) * $signed(_zz_405));
  assign _zz_2295 = _zz_7784[15 : 0];
  assign _zz_4340 = ($signed(_zz_7785) * $signed(twiddle_factor_table_1_real));
  assign _zz_4341 = ($signed(_zz_7786) * $signed(twiddle_factor_table_1_imag));
  assign _zz_2293 = ($signed(_zz_2295) - $signed(_zz_7787));
  assign _zz_2294 = ($signed(_zz_2295) + $signed(_zz_7789));
  assign _zz_2296 = 1'b1;
  assign _zz_2297 = 1'b1;
  assign _zz_4342 = ($signed(_zz_7807) * $signed(_zz_407));
  assign _zz_2300 = _zz_7808[15 : 0];
  assign _zz_4343 = ($signed(_zz_7809) * $signed(twiddle_factor_table_2_real));
  assign _zz_4344 = ($signed(_zz_7810) * $signed(twiddle_factor_table_2_imag));
  assign _zz_2298 = ($signed(_zz_2300) - $signed(_zz_7811));
  assign _zz_2299 = ($signed(_zz_2300) + $signed(_zz_7813));
  assign _zz_2301 = 1'b1;
  assign _zz_2302 = 1'b1;
  assign _zz_4345 = ($signed(_zz_7831) * $signed(_zz_413));
  assign _zz_2305 = _zz_7832[15 : 0];
  assign _zz_4346 = ($signed(_zz_7833) * $signed(twiddle_factor_table_1_real));
  assign _zz_4347 = ($signed(_zz_7834) * $signed(twiddle_factor_table_1_imag));
  assign _zz_2303 = ($signed(_zz_2305) - $signed(_zz_7835));
  assign _zz_2304 = ($signed(_zz_2305) + $signed(_zz_7837));
  assign _zz_2306 = 1'b1;
  assign _zz_2307 = 1'b1;
  assign _zz_4348 = ($signed(_zz_7855) * $signed(_zz_415));
  assign _zz_2310 = _zz_7856[15 : 0];
  assign _zz_4349 = ($signed(_zz_7857) * $signed(twiddle_factor_table_2_real));
  assign _zz_4350 = ($signed(_zz_7858) * $signed(twiddle_factor_table_2_imag));
  assign _zz_2308 = ($signed(_zz_2310) - $signed(_zz_7859));
  assign _zz_2309 = ($signed(_zz_2310) + $signed(_zz_7861));
  assign _zz_2311 = 1'b1;
  assign _zz_2312 = 1'b1;
  assign _zz_4351 = ($signed(_zz_7879) * $signed(_zz_421));
  assign _zz_2315 = _zz_7880[15 : 0];
  assign _zz_4352 = ($signed(_zz_7881) * $signed(twiddle_factor_table_1_real));
  assign _zz_4353 = ($signed(_zz_7882) * $signed(twiddle_factor_table_1_imag));
  assign _zz_2313 = ($signed(_zz_2315) - $signed(_zz_7883));
  assign _zz_2314 = ($signed(_zz_2315) + $signed(_zz_7885));
  assign _zz_2316 = 1'b1;
  assign _zz_2317 = 1'b1;
  assign _zz_4354 = ($signed(_zz_7903) * $signed(_zz_423));
  assign _zz_2320 = _zz_7904[15 : 0];
  assign _zz_4355 = ($signed(_zz_7905) * $signed(twiddle_factor_table_2_real));
  assign _zz_4356 = ($signed(_zz_7906) * $signed(twiddle_factor_table_2_imag));
  assign _zz_2318 = ($signed(_zz_2320) - $signed(_zz_7907));
  assign _zz_2319 = ($signed(_zz_2320) + $signed(_zz_7909));
  assign _zz_2321 = 1'b1;
  assign _zz_2322 = 1'b1;
  assign _zz_4357 = ($signed(_zz_7927) * $signed(_zz_429));
  assign _zz_2325 = _zz_7928[15 : 0];
  assign _zz_4358 = ($signed(_zz_7929) * $signed(twiddle_factor_table_1_real));
  assign _zz_4359 = ($signed(_zz_7930) * $signed(twiddle_factor_table_1_imag));
  assign _zz_2323 = ($signed(_zz_2325) - $signed(_zz_7931));
  assign _zz_2324 = ($signed(_zz_2325) + $signed(_zz_7933));
  assign _zz_2326 = 1'b1;
  assign _zz_2327 = 1'b1;
  assign _zz_4360 = ($signed(_zz_7951) * $signed(_zz_431));
  assign _zz_2330 = _zz_7952[15 : 0];
  assign _zz_4361 = ($signed(_zz_7953) * $signed(twiddle_factor_table_2_real));
  assign _zz_4362 = ($signed(_zz_7954) * $signed(twiddle_factor_table_2_imag));
  assign _zz_2328 = ($signed(_zz_2330) - $signed(_zz_7955));
  assign _zz_2329 = ($signed(_zz_2330) + $signed(_zz_7957));
  assign _zz_2331 = 1'b1;
  assign _zz_2332 = 1'b1;
  assign _zz_4363 = ($signed(_zz_7975) * $signed(_zz_437));
  assign _zz_2335 = _zz_7976[15 : 0];
  assign _zz_4364 = ($signed(_zz_7977) * $signed(twiddle_factor_table_1_real));
  assign _zz_4365 = ($signed(_zz_7978) * $signed(twiddle_factor_table_1_imag));
  assign _zz_2333 = ($signed(_zz_2335) - $signed(_zz_7979));
  assign _zz_2334 = ($signed(_zz_2335) + $signed(_zz_7981));
  assign _zz_2336 = 1'b1;
  assign _zz_2337 = 1'b1;
  assign _zz_4366 = ($signed(_zz_7999) * $signed(_zz_439));
  assign _zz_2340 = _zz_8000[15 : 0];
  assign _zz_4367 = ($signed(_zz_8001) * $signed(twiddle_factor_table_2_real));
  assign _zz_4368 = ($signed(_zz_8002) * $signed(twiddle_factor_table_2_imag));
  assign _zz_2338 = ($signed(_zz_2340) - $signed(_zz_8003));
  assign _zz_2339 = ($signed(_zz_2340) + $signed(_zz_8005));
  assign _zz_2341 = 1'b1;
  assign _zz_2342 = 1'b1;
  assign _zz_4369 = ($signed(_zz_8023) * $signed(_zz_445));
  assign _zz_2345 = _zz_8024[15 : 0];
  assign _zz_4370 = ($signed(_zz_8025) * $signed(twiddle_factor_table_1_real));
  assign _zz_4371 = ($signed(_zz_8026) * $signed(twiddle_factor_table_1_imag));
  assign _zz_2343 = ($signed(_zz_2345) - $signed(_zz_8027));
  assign _zz_2344 = ($signed(_zz_2345) + $signed(_zz_8029));
  assign _zz_2346 = 1'b1;
  assign _zz_2347 = 1'b1;
  assign _zz_4372 = ($signed(_zz_8047) * $signed(_zz_447));
  assign _zz_2350 = _zz_8048[15 : 0];
  assign _zz_4373 = ($signed(_zz_8049) * $signed(twiddle_factor_table_2_real));
  assign _zz_4374 = ($signed(_zz_8050) * $signed(twiddle_factor_table_2_imag));
  assign _zz_2348 = ($signed(_zz_2350) - $signed(_zz_8051));
  assign _zz_2349 = ($signed(_zz_2350) + $signed(_zz_8053));
  assign _zz_2351 = 1'b1;
  assign _zz_2352 = 1'b1;
  assign _zz_4375 = ($signed(_zz_8071) * $signed(_zz_453));
  assign _zz_2355 = _zz_8072[15 : 0];
  assign _zz_4376 = ($signed(_zz_8073) * $signed(twiddle_factor_table_1_real));
  assign _zz_4377 = ($signed(_zz_8074) * $signed(twiddle_factor_table_1_imag));
  assign _zz_2353 = ($signed(_zz_2355) - $signed(_zz_8075));
  assign _zz_2354 = ($signed(_zz_2355) + $signed(_zz_8077));
  assign _zz_2356 = 1'b1;
  assign _zz_2357 = 1'b1;
  assign _zz_4378 = ($signed(_zz_8095) * $signed(_zz_455));
  assign _zz_2360 = _zz_8096[15 : 0];
  assign _zz_4379 = ($signed(_zz_8097) * $signed(twiddle_factor_table_2_real));
  assign _zz_4380 = ($signed(_zz_8098) * $signed(twiddle_factor_table_2_imag));
  assign _zz_2358 = ($signed(_zz_2360) - $signed(_zz_8099));
  assign _zz_2359 = ($signed(_zz_2360) + $signed(_zz_8101));
  assign _zz_2361 = 1'b1;
  assign _zz_2362 = 1'b1;
  assign _zz_4381 = ($signed(_zz_8119) * $signed(_zz_461));
  assign _zz_2365 = _zz_8120[15 : 0];
  assign _zz_4382 = ($signed(_zz_8121) * $signed(twiddle_factor_table_1_real));
  assign _zz_4383 = ($signed(_zz_8122) * $signed(twiddle_factor_table_1_imag));
  assign _zz_2363 = ($signed(_zz_2365) - $signed(_zz_8123));
  assign _zz_2364 = ($signed(_zz_2365) + $signed(_zz_8125));
  assign _zz_2366 = 1'b1;
  assign _zz_2367 = 1'b1;
  assign _zz_4384 = ($signed(_zz_8143) * $signed(_zz_463));
  assign _zz_2370 = _zz_8144[15 : 0];
  assign _zz_4385 = ($signed(_zz_8145) * $signed(twiddle_factor_table_2_real));
  assign _zz_4386 = ($signed(_zz_8146) * $signed(twiddle_factor_table_2_imag));
  assign _zz_2368 = ($signed(_zz_2370) - $signed(_zz_8147));
  assign _zz_2369 = ($signed(_zz_2370) + $signed(_zz_8149));
  assign _zz_2371 = 1'b1;
  assign _zz_2372 = 1'b1;
  assign _zz_4387 = ($signed(_zz_8167) * $signed(_zz_469));
  assign _zz_2375 = _zz_8168[15 : 0];
  assign _zz_4388 = ($signed(_zz_8169) * $signed(twiddle_factor_table_1_real));
  assign _zz_4389 = ($signed(_zz_8170) * $signed(twiddle_factor_table_1_imag));
  assign _zz_2373 = ($signed(_zz_2375) - $signed(_zz_8171));
  assign _zz_2374 = ($signed(_zz_2375) + $signed(_zz_8173));
  assign _zz_2376 = 1'b1;
  assign _zz_2377 = 1'b1;
  assign _zz_4390 = ($signed(_zz_8191) * $signed(_zz_471));
  assign _zz_2380 = _zz_8192[15 : 0];
  assign _zz_4391 = ($signed(_zz_8193) * $signed(twiddle_factor_table_2_real));
  assign _zz_4392 = ($signed(_zz_8194) * $signed(twiddle_factor_table_2_imag));
  assign _zz_2378 = ($signed(_zz_2380) - $signed(_zz_8195));
  assign _zz_2379 = ($signed(_zz_2380) + $signed(_zz_8197));
  assign _zz_2381 = 1'b1;
  assign _zz_2382 = 1'b1;
  assign _zz_4393 = ($signed(_zz_8215) * $signed(_zz_477));
  assign _zz_2385 = _zz_8216[15 : 0];
  assign _zz_4394 = ($signed(_zz_8217) * $signed(twiddle_factor_table_1_real));
  assign _zz_4395 = ($signed(_zz_8218) * $signed(twiddle_factor_table_1_imag));
  assign _zz_2383 = ($signed(_zz_2385) - $signed(_zz_8219));
  assign _zz_2384 = ($signed(_zz_2385) + $signed(_zz_8221));
  assign _zz_2386 = 1'b1;
  assign _zz_2387 = 1'b1;
  assign _zz_4396 = ($signed(_zz_8239) * $signed(_zz_479));
  assign _zz_2390 = _zz_8240[15 : 0];
  assign _zz_4397 = ($signed(_zz_8241) * $signed(twiddle_factor_table_2_real));
  assign _zz_4398 = ($signed(_zz_8242) * $signed(twiddle_factor_table_2_imag));
  assign _zz_2388 = ($signed(_zz_2390) - $signed(_zz_8243));
  assign _zz_2389 = ($signed(_zz_2390) + $signed(_zz_8245));
  assign _zz_2391 = 1'b1;
  assign _zz_2392 = 1'b1;
  assign _zz_4399 = ($signed(_zz_8263) * $signed(_zz_485));
  assign _zz_2395 = _zz_8264[15 : 0];
  assign _zz_4400 = ($signed(_zz_8265) * $signed(twiddle_factor_table_1_real));
  assign _zz_4401 = ($signed(_zz_8266) * $signed(twiddle_factor_table_1_imag));
  assign _zz_2393 = ($signed(_zz_2395) - $signed(_zz_8267));
  assign _zz_2394 = ($signed(_zz_2395) + $signed(_zz_8269));
  assign _zz_2396 = 1'b1;
  assign _zz_2397 = 1'b1;
  assign _zz_4402 = ($signed(_zz_8287) * $signed(_zz_487));
  assign _zz_2400 = _zz_8288[15 : 0];
  assign _zz_4403 = ($signed(_zz_8289) * $signed(twiddle_factor_table_2_real));
  assign _zz_4404 = ($signed(_zz_8290) * $signed(twiddle_factor_table_2_imag));
  assign _zz_2398 = ($signed(_zz_2400) - $signed(_zz_8291));
  assign _zz_2399 = ($signed(_zz_2400) + $signed(_zz_8293));
  assign _zz_2401 = 1'b1;
  assign _zz_2402 = 1'b1;
  assign _zz_4405 = ($signed(_zz_8311) * $signed(_zz_493));
  assign _zz_2405 = _zz_8312[15 : 0];
  assign _zz_4406 = ($signed(_zz_8313) * $signed(twiddle_factor_table_1_real));
  assign _zz_4407 = ($signed(_zz_8314) * $signed(twiddle_factor_table_1_imag));
  assign _zz_2403 = ($signed(_zz_2405) - $signed(_zz_8315));
  assign _zz_2404 = ($signed(_zz_2405) + $signed(_zz_8317));
  assign _zz_2406 = 1'b1;
  assign _zz_2407 = 1'b1;
  assign _zz_4408 = ($signed(_zz_8335) * $signed(_zz_495));
  assign _zz_2410 = _zz_8336[15 : 0];
  assign _zz_4409 = ($signed(_zz_8337) * $signed(twiddle_factor_table_2_real));
  assign _zz_4410 = ($signed(_zz_8338) * $signed(twiddle_factor_table_2_imag));
  assign _zz_2408 = ($signed(_zz_2410) - $signed(_zz_8339));
  assign _zz_2409 = ($signed(_zz_2410) + $signed(_zz_8341));
  assign _zz_2411 = 1'b1;
  assign _zz_2412 = 1'b1;
  assign _zz_4411 = ($signed(_zz_8359) * $signed(_zz_501));
  assign _zz_2415 = _zz_8360[15 : 0];
  assign _zz_4412 = ($signed(_zz_8361) * $signed(twiddle_factor_table_1_real));
  assign _zz_4413 = ($signed(_zz_8362) * $signed(twiddle_factor_table_1_imag));
  assign _zz_2413 = ($signed(_zz_2415) - $signed(_zz_8363));
  assign _zz_2414 = ($signed(_zz_2415) + $signed(_zz_8365));
  assign _zz_2416 = 1'b1;
  assign _zz_2417 = 1'b1;
  assign _zz_4414 = ($signed(_zz_8383) * $signed(_zz_503));
  assign _zz_2420 = _zz_8384[15 : 0];
  assign _zz_4415 = ($signed(_zz_8385) * $signed(twiddle_factor_table_2_real));
  assign _zz_4416 = ($signed(_zz_8386) * $signed(twiddle_factor_table_2_imag));
  assign _zz_2418 = ($signed(_zz_2420) - $signed(_zz_8387));
  assign _zz_2419 = ($signed(_zz_2420) + $signed(_zz_8389));
  assign _zz_2421 = 1'b1;
  assign _zz_2422 = 1'b1;
  assign _zz_4417 = ($signed(_zz_8407) * $signed(_zz_509));
  assign _zz_2425 = _zz_8408[15 : 0];
  assign _zz_4418 = ($signed(_zz_8409) * $signed(twiddle_factor_table_1_real));
  assign _zz_4419 = ($signed(_zz_8410) * $signed(twiddle_factor_table_1_imag));
  assign _zz_2423 = ($signed(_zz_2425) - $signed(_zz_8411));
  assign _zz_2424 = ($signed(_zz_2425) + $signed(_zz_8413));
  assign _zz_2426 = 1'b1;
  assign _zz_2427 = 1'b1;
  assign _zz_4420 = ($signed(_zz_8431) * $signed(_zz_511));
  assign _zz_2430 = _zz_8432[15 : 0];
  assign _zz_4421 = ($signed(_zz_8433) * $signed(twiddle_factor_table_2_real));
  assign _zz_4422 = ($signed(_zz_8434) * $signed(twiddle_factor_table_2_imag));
  assign _zz_2428 = ($signed(_zz_2430) - $signed(_zz_8435));
  assign _zz_2429 = ($signed(_zz_2430) + $signed(_zz_8437));
  assign _zz_2431 = 1'b1;
  assign _zz_2432 = 1'b1;
  assign _zz_4423 = ($signed(_zz_8455) * $signed(_zz_521));
  assign _zz_2435 = _zz_8456[15 : 0];
  assign _zz_4424 = ($signed(_zz_8457) * $signed(twiddle_factor_table_3_real));
  assign _zz_4425 = ($signed(_zz_8458) * $signed(twiddle_factor_table_3_imag));
  assign _zz_2433 = ($signed(_zz_2435) - $signed(_zz_8459));
  assign _zz_2434 = ($signed(_zz_2435) + $signed(_zz_8461));
  assign _zz_2436 = 1'b1;
  assign _zz_2437 = 1'b1;
  assign _zz_4426 = ($signed(_zz_8479) * $signed(_zz_523));
  assign _zz_2440 = _zz_8480[15 : 0];
  assign _zz_4427 = ($signed(_zz_8481) * $signed(twiddle_factor_table_4_real));
  assign _zz_4428 = ($signed(_zz_8482) * $signed(twiddle_factor_table_4_imag));
  assign _zz_2438 = ($signed(_zz_2440) - $signed(_zz_8483));
  assign _zz_2439 = ($signed(_zz_2440) + $signed(_zz_8485));
  assign _zz_2441 = 1'b1;
  assign _zz_2442 = 1'b1;
  assign _zz_4429 = ($signed(_zz_8503) * $signed(_zz_525));
  assign _zz_2445 = _zz_8504[15 : 0];
  assign _zz_4430 = ($signed(_zz_8505) * $signed(twiddle_factor_table_5_real));
  assign _zz_4431 = ($signed(_zz_8506) * $signed(twiddle_factor_table_5_imag));
  assign _zz_2443 = ($signed(_zz_2445) - $signed(_zz_8507));
  assign _zz_2444 = ($signed(_zz_2445) + $signed(_zz_8509));
  assign _zz_2446 = 1'b1;
  assign _zz_2447 = 1'b1;
  assign _zz_4432 = ($signed(_zz_8527) * $signed(_zz_527));
  assign _zz_2450 = _zz_8528[15 : 0];
  assign _zz_4433 = ($signed(_zz_8529) * $signed(twiddle_factor_table_6_real));
  assign _zz_4434 = ($signed(_zz_8530) * $signed(twiddle_factor_table_6_imag));
  assign _zz_2448 = ($signed(_zz_2450) - $signed(_zz_8531));
  assign _zz_2449 = ($signed(_zz_2450) + $signed(_zz_8533));
  assign _zz_2451 = 1'b1;
  assign _zz_2452 = 1'b1;
  assign _zz_4435 = ($signed(_zz_8551) * $signed(_zz_537));
  assign _zz_2455 = _zz_8552[15 : 0];
  assign _zz_4436 = ($signed(_zz_8553) * $signed(twiddle_factor_table_3_real));
  assign _zz_4437 = ($signed(_zz_8554) * $signed(twiddle_factor_table_3_imag));
  assign _zz_2453 = ($signed(_zz_2455) - $signed(_zz_8555));
  assign _zz_2454 = ($signed(_zz_2455) + $signed(_zz_8557));
  assign _zz_2456 = 1'b1;
  assign _zz_2457 = 1'b1;
  assign _zz_4438 = ($signed(_zz_8575) * $signed(_zz_539));
  assign _zz_2460 = _zz_8576[15 : 0];
  assign _zz_4439 = ($signed(_zz_8577) * $signed(twiddle_factor_table_4_real));
  assign _zz_4440 = ($signed(_zz_8578) * $signed(twiddle_factor_table_4_imag));
  assign _zz_2458 = ($signed(_zz_2460) - $signed(_zz_8579));
  assign _zz_2459 = ($signed(_zz_2460) + $signed(_zz_8581));
  assign _zz_2461 = 1'b1;
  assign _zz_2462 = 1'b1;
  assign _zz_4441 = ($signed(_zz_8599) * $signed(_zz_541));
  assign _zz_2465 = _zz_8600[15 : 0];
  assign _zz_4442 = ($signed(_zz_8601) * $signed(twiddle_factor_table_5_real));
  assign _zz_4443 = ($signed(_zz_8602) * $signed(twiddle_factor_table_5_imag));
  assign _zz_2463 = ($signed(_zz_2465) - $signed(_zz_8603));
  assign _zz_2464 = ($signed(_zz_2465) + $signed(_zz_8605));
  assign _zz_2466 = 1'b1;
  assign _zz_2467 = 1'b1;
  assign _zz_4444 = ($signed(_zz_8623) * $signed(_zz_543));
  assign _zz_2470 = _zz_8624[15 : 0];
  assign _zz_4445 = ($signed(_zz_8625) * $signed(twiddle_factor_table_6_real));
  assign _zz_4446 = ($signed(_zz_8626) * $signed(twiddle_factor_table_6_imag));
  assign _zz_2468 = ($signed(_zz_2470) - $signed(_zz_8627));
  assign _zz_2469 = ($signed(_zz_2470) + $signed(_zz_8629));
  assign _zz_2471 = 1'b1;
  assign _zz_2472 = 1'b1;
  assign _zz_4447 = ($signed(_zz_8647) * $signed(_zz_553));
  assign _zz_2475 = _zz_8648[15 : 0];
  assign _zz_4448 = ($signed(_zz_8649) * $signed(twiddle_factor_table_3_real));
  assign _zz_4449 = ($signed(_zz_8650) * $signed(twiddle_factor_table_3_imag));
  assign _zz_2473 = ($signed(_zz_2475) - $signed(_zz_8651));
  assign _zz_2474 = ($signed(_zz_2475) + $signed(_zz_8653));
  assign _zz_2476 = 1'b1;
  assign _zz_2477 = 1'b1;
  assign _zz_4450 = ($signed(_zz_8671) * $signed(_zz_555));
  assign _zz_2480 = _zz_8672[15 : 0];
  assign _zz_4451 = ($signed(_zz_8673) * $signed(twiddle_factor_table_4_real));
  assign _zz_4452 = ($signed(_zz_8674) * $signed(twiddle_factor_table_4_imag));
  assign _zz_2478 = ($signed(_zz_2480) - $signed(_zz_8675));
  assign _zz_2479 = ($signed(_zz_2480) + $signed(_zz_8677));
  assign _zz_2481 = 1'b1;
  assign _zz_2482 = 1'b1;
  assign _zz_4453 = ($signed(_zz_8695) * $signed(_zz_557));
  assign _zz_2485 = _zz_8696[15 : 0];
  assign _zz_4454 = ($signed(_zz_8697) * $signed(twiddle_factor_table_5_real));
  assign _zz_4455 = ($signed(_zz_8698) * $signed(twiddle_factor_table_5_imag));
  assign _zz_2483 = ($signed(_zz_2485) - $signed(_zz_8699));
  assign _zz_2484 = ($signed(_zz_2485) + $signed(_zz_8701));
  assign _zz_2486 = 1'b1;
  assign _zz_2487 = 1'b1;
  assign _zz_4456 = ($signed(_zz_8719) * $signed(_zz_559));
  assign _zz_2490 = _zz_8720[15 : 0];
  assign _zz_4457 = ($signed(_zz_8721) * $signed(twiddle_factor_table_6_real));
  assign _zz_4458 = ($signed(_zz_8722) * $signed(twiddle_factor_table_6_imag));
  assign _zz_2488 = ($signed(_zz_2490) - $signed(_zz_8723));
  assign _zz_2489 = ($signed(_zz_2490) + $signed(_zz_8725));
  assign _zz_2491 = 1'b1;
  assign _zz_2492 = 1'b1;
  assign _zz_4459 = ($signed(_zz_8743) * $signed(_zz_569));
  assign _zz_2495 = _zz_8744[15 : 0];
  assign _zz_4460 = ($signed(_zz_8745) * $signed(twiddle_factor_table_3_real));
  assign _zz_4461 = ($signed(_zz_8746) * $signed(twiddle_factor_table_3_imag));
  assign _zz_2493 = ($signed(_zz_2495) - $signed(_zz_8747));
  assign _zz_2494 = ($signed(_zz_2495) + $signed(_zz_8749));
  assign _zz_2496 = 1'b1;
  assign _zz_2497 = 1'b1;
  assign _zz_4462 = ($signed(_zz_8767) * $signed(_zz_571));
  assign _zz_2500 = _zz_8768[15 : 0];
  assign _zz_4463 = ($signed(_zz_8769) * $signed(twiddle_factor_table_4_real));
  assign _zz_4464 = ($signed(_zz_8770) * $signed(twiddle_factor_table_4_imag));
  assign _zz_2498 = ($signed(_zz_2500) - $signed(_zz_8771));
  assign _zz_2499 = ($signed(_zz_2500) + $signed(_zz_8773));
  assign _zz_2501 = 1'b1;
  assign _zz_2502 = 1'b1;
  assign _zz_4465 = ($signed(_zz_8791) * $signed(_zz_573));
  assign _zz_2505 = _zz_8792[15 : 0];
  assign _zz_4466 = ($signed(_zz_8793) * $signed(twiddle_factor_table_5_real));
  assign _zz_4467 = ($signed(_zz_8794) * $signed(twiddle_factor_table_5_imag));
  assign _zz_2503 = ($signed(_zz_2505) - $signed(_zz_8795));
  assign _zz_2504 = ($signed(_zz_2505) + $signed(_zz_8797));
  assign _zz_2506 = 1'b1;
  assign _zz_2507 = 1'b1;
  assign _zz_4468 = ($signed(_zz_8815) * $signed(_zz_575));
  assign _zz_2510 = _zz_8816[15 : 0];
  assign _zz_4469 = ($signed(_zz_8817) * $signed(twiddle_factor_table_6_real));
  assign _zz_4470 = ($signed(_zz_8818) * $signed(twiddle_factor_table_6_imag));
  assign _zz_2508 = ($signed(_zz_2510) - $signed(_zz_8819));
  assign _zz_2509 = ($signed(_zz_2510) + $signed(_zz_8821));
  assign _zz_2511 = 1'b1;
  assign _zz_2512 = 1'b1;
  assign _zz_4471 = ($signed(_zz_8839) * $signed(_zz_585));
  assign _zz_2515 = _zz_8840[15 : 0];
  assign _zz_4472 = ($signed(_zz_8841) * $signed(twiddle_factor_table_3_real));
  assign _zz_4473 = ($signed(_zz_8842) * $signed(twiddle_factor_table_3_imag));
  assign _zz_2513 = ($signed(_zz_2515) - $signed(_zz_8843));
  assign _zz_2514 = ($signed(_zz_2515) + $signed(_zz_8845));
  assign _zz_2516 = 1'b1;
  assign _zz_2517 = 1'b1;
  assign _zz_4474 = ($signed(_zz_8863) * $signed(_zz_587));
  assign _zz_2520 = _zz_8864[15 : 0];
  assign _zz_4475 = ($signed(_zz_8865) * $signed(twiddle_factor_table_4_real));
  assign _zz_4476 = ($signed(_zz_8866) * $signed(twiddle_factor_table_4_imag));
  assign _zz_2518 = ($signed(_zz_2520) - $signed(_zz_8867));
  assign _zz_2519 = ($signed(_zz_2520) + $signed(_zz_8869));
  assign _zz_2521 = 1'b1;
  assign _zz_2522 = 1'b1;
  assign _zz_4477 = ($signed(_zz_8887) * $signed(_zz_589));
  assign _zz_2525 = _zz_8888[15 : 0];
  assign _zz_4478 = ($signed(_zz_8889) * $signed(twiddle_factor_table_5_real));
  assign _zz_4479 = ($signed(_zz_8890) * $signed(twiddle_factor_table_5_imag));
  assign _zz_2523 = ($signed(_zz_2525) - $signed(_zz_8891));
  assign _zz_2524 = ($signed(_zz_2525) + $signed(_zz_8893));
  assign _zz_2526 = 1'b1;
  assign _zz_2527 = 1'b1;
  assign _zz_4480 = ($signed(_zz_8911) * $signed(_zz_591));
  assign _zz_2530 = _zz_8912[15 : 0];
  assign _zz_4481 = ($signed(_zz_8913) * $signed(twiddle_factor_table_6_real));
  assign _zz_4482 = ($signed(_zz_8914) * $signed(twiddle_factor_table_6_imag));
  assign _zz_2528 = ($signed(_zz_2530) - $signed(_zz_8915));
  assign _zz_2529 = ($signed(_zz_2530) + $signed(_zz_8917));
  assign _zz_2531 = 1'b1;
  assign _zz_2532 = 1'b1;
  assign _zz_4483 = ($signed(_zz_8935) * $signed(_zz_601));
  assign _zz_2535 = _zz_8936[15 : 0];
  assign _zz_4484 = ($signed(_zz_8937) * $signed(twiddle_factor_table_3_real));
  assign _zz_4485 = ($signed(_zz_8938) * $signed(twiddle_factor_table_3_imag));
  assign _zz_2533 = ($signed(_zz_2535) - $signed(_zz_8939));
  assign _zz_2534 = ($signed(_zz_2535) + $signed(_zz_8941));
  assign _zz_2536 = 1'b1;
  assign _zz_2537 = 1'b1;
  assign _zz_4486 = ($signed(_zz_8959) * $signed(_zz_603));
  assign _zz_2540 = _zz_8960[15 : 0];
  assign _zz_4487 = ($signed(_zz_8961) * $signed(twiddle_factor_table_4_real));
  assign _zz_4488 = ($signed(_zz_8962) * $signed(twiddle_factor_table_4_imag));
  assign _zz_2538 = ($signed(_zz_2540) - $signed(_zz_8963));
  assign _zz_2539 = ($signed(_zz_2540) + $signed(_zz_8965));
  assign _zz_2541 = 1'b1;
  assign _zz_2542 = 1'b1;
  assign _zz_4489 = ($signed(_zz_8983) * $signed(_zz_605));
  assign _zz_2545 = _zz_8984[15 : 0];
  assign _zz_4490 = ($signed(_zz_8985) * $signed(twiddle_factor_table_5_real));
  assign _zz_4491 = ($signed(_zz_8986) * $signed(twiddle_factor_table_5_imag));
  assign _zz_2543 = ($signed(_zz_2545) - $signed(_zz_8987));
  assign _zz_2544 = ($signed(_zz_2545) + $signed(_zz_8989));
  assign _zz_2546 = 1'b1;
  assign _zz_2547 = 1'b1;
  assign _zz_4492 = ($signed(_zz_9007) * $signed(_zz_607));
  assign _zz_2550 = _zz_9008[15 : 0];
  assign _zz_4493 = ($signed(_zz_9009) * $signed(twiddle_factor_table_6_real));
  assign _zz_4494 = ($signed(_zz_9010) * $signed(twiddle_factor_table_6_imag));
  assign _zz_2548 = ($signed(_zz_2550) - $signed(_zz_9011));
  assign _zz_2549 = ($signed(_zz_2550) + $signed(_zz_9013));
  assign _zz_2551 = 1'b1;
  assign _zz_2552 = 1'b1;
  assign _zz_4495 = ($signed(_zz_9031) * $signed(_zz_617));
  assign _zz_2555 = _zz_9032[15 : 0];
  assign _zz_4496 = ($signed(_zz_9033) * $signed(twiddle_factor_table_3_real));
  assign _zz_4497 = ($signed(_zz_9034) * $signed(twiddle_factor_table_3_imag));
  assign _zz_2553 = ($signed(_zz_2555) - $signed(_zz_9035));
  assign _zz_2554 = ($signed(_zz_2555) + $signed(_zz_9037));
  assign _zz_2556 = 1'b1;
  assign _zz_2557 = 1'b1;
  assign _zz_4498 = ($signed(_zz_9055) * $signed(_zz_619));
  assign _zz_2560 = _zz_9056[15 : 0];
  assign _zz_4499 = ($signed(_zz_9057) * $signed(twiddle_factor_table_4_real));
  assign _zz_4500 = ($signed(_zz_9058) * $signed(twiddle_factor_table_4_imag));
  assign _zz_2558 = ($signed(_zz_2560) - $signed(_zz_9059));
  assign _zz_2559 = ($signed(_zz_2560) + $signed(_zz_9061));
  assign _zz_2561 = 1'b1;
  assign _zz_2562 = 1'b1;
  assign _zz_4501 = ($signed(_zz_9079) * $signed(_zz_621));
  assign _zz_2565 = _zz_9080[15 : 0];
  assign _zz_4502 = ($signed(_zz_9081) * $signed(twiddle_factor_table_5_real));
  assign _zz_4503 = ($signed(_zz_9082) * $signed(twiddle_factor_table_5_imag));
  assign _zz_2563 = ($signed(_zz_2565) - $signed(_zz_9083));
  assign _zz_2564 = ($signed(_zz_2565) + $signed(_zz_9085));
  assign _zz_2566 = 1'b1;
  assign _zz_2567 = 1'b1;
  assign _zz_4504 = ($signed(_zz_9103) * $signed(_zz_623));
  assign _zz_2570 = _zz_9104[15 : 0];
  assign _zz_4505 = ($signed(_zz_9105) * $signed(twiddle_factor_table_6_real));
  assign _zz_4506 = ($signed(_zz_9106) * $signed(twiddle_factor_table_6_imag));
  assign _zz_2568 = ($signed(_zz_2570) - $signed(_zz_9107));
  assign _zz_2569 = ($signed(_zz_2570) + $signed(_zz_9109));
  assign _zz_2571 = 1'b1;
  assign _zz_2572 = 1'b1;
  assign _zz_4507 = ($signed(_zz_9127) * $signed(_zz_633));
  assign _zz_2575 = _zz_9128[15 : 0];
  assign _zz_4508 = ($signed(_zz_9129) * $signed(twiddle_factor_table_3_real));
  assign _zz_4509 = ($signed(_zz_9130) * $signed(twiddle_factor_table_3_imag));
  assign _zz_2573 = ($signed(_zz_2575) - $signed(_zz_9131));
  assign _zz_2574 = ($signed(_zz_2575) + $signed(_zz_9133));
  assign _zz_2576 = 1'b1;
  assign _zz_2577 = 1'b1;
  assign _zz_4510 = ($signed(_zz_9151) * $signed(_zz_635));
  assign _zz_2580 = _zz_9152[15 : 0];
  assign _zz_4511 = ($signed(_zz_9153) * $signed(twiddle_factor_table_4_real));
  assign _zz_4512 = ($signed(_zz_9154) * $signed(twiddle_factor_table_4_imag));
  assign _zz_2578 = ($signed(_zz_2580) - $signed(_zz_9155));
  assign _zz_2579 = ($signed(_zz_2580) + $signed(_zz_9157));
  assign _zz_2581 = 1'b1;
  assign _zz_2582 = 1'b1;
  assign _zz_4513 = ($signed(_zz_9175) * $signed(_zz_637));
  assign _zz_2585 = _zz_9176[15 : 0];
  assign _zz_4514 = ($signed(_zz_9177) * $signed(twiddle_factor_table_5_real));
  assign _zz_4515 = ($signed(_zz_9178) * $signed(twiddle_factor_table_5_imag));
  assign _zz_2583 = ($signed(_zz_2585) - $signed(_zz_9179));
  assign _zz_2584 = ($signed(_zz_2585) + $signed(_zz_9181));
  assign _zz_2586 = 1'b1;
  assign _zz_2587 = 1'b1;
  assign _zz_4516 = ($signed(_zz_9199) * $signed(_zz_639));
  assign _zz_2590 = _zz_9200[15 : 0];
  assign _zz_4517 = ($signed(_zz_9201) * $signed(twiddle_factor_table_6_real));
  assign _zz_4518 = ($signed(_zz_9202) * $signed(twiddle_factor_table_6_imag));
  assign _zz_2588 = ($signed(_zz_2590) - $signed(_zz_9203));
  assign _zz_2589 = ($signed(_zz_2590) + $signed(_zz_9205));
  assign _zz_2591 = 1'b1;
  assign _zz_2592 = 1'b1;
  assign _zz_4519 = ($signed(_zz_9223) * $signed(_zz_649));
  assign _zz_2595 = _zz_9224[15 : 0];
  assign _zz_4520 = ($signed(_zz_9225) * $signed(twiddle_factor_table_3_real));
  assign _zz_4521 = ($signed(_zz_9226) * $signed(twiddle_factor_table_3_imag));
  assign _zz_2593 = ($signed(_zz_2595) - $signed(_zz_9227));
  assign _zz_2594 = ($signed(_zz_2595) + $signed(_zz_9229));
  assign _zz_2596 = 1'b1;
  assign _zz_2597 = 1'b1;
  assign _zz_4522 = ($signed(_zz_9247) * $signed(_zz_651));
  assign _zz_2600 = _zz_9248[15 : 0];
  assign _zz_4523 = ($signed(_zz_9249) * $signed(twiddle_factor_table_4_real));
  assign _zz_4524 = ($signed(_zz_9250) * $signed(twiddle_factor_table_4_imag));
  assign _zz_2598 = ($signed(_zz_2600) - $signed(_zz_9251));
  assign _zz_2599 = ($signed(_zz_2600) + $signed(_zz_9253));
  assign _zz_2601 = 1'b1;
  assign _zz_2602 = 1'b1;
  assign _zz_4525 = ($signed(_zz_9271) * $signed(_zz_653));
  assign _zz_2605 = _zz_9272[15 : 0];
  assign _zz_4526 = ($signed(_zz_9273) * $signed(twiddle_factor_table_5_real));
  assign _zz_4527 = ($signed(_zz_9274) * $signed(twiddle_factor_table_5_imag));
  assign _zz_2603 = ($signed(_zz_2605) - $signed(_zz_9275));
  assign _zz_2604 = ($signed(_zz_2605) + $signed(_zz_9277));
  assign _zz_2606 = 1'b1;
  assign _zz_2607 = 1'b1;
  assign _zz_4528 = ($signed(_zz_9295) * $signed(_zz_655));
  assign _zz_2610 = _zz_9296[15 : 0];
  assign _zz_4529 = ($signed(_zz_9297) * $signed(twiddle_factor_table_6_real));
  assign _zz_4530 = ($signed(_zz_9298) * $signed(twiddle_factor_table_6_imag));
  assign _zz_2608 = ($signed(_zz_2610) - $signed(_zz_9299));
  assign _zz_2609 = ($signed(_zz_2610) + $signed(_zz_9301));
  assign _zz_2611 = 1'b1;
  assign _zz_2612 = 1'b1;
  assign _zz_4531 = ($signed(_zz_9319) * $signed(_zz_665));
  assign _zz_2615 = _zz_9320[15 : 0];
  assign _zz_4532 = ($signed(_zz_9321) * $signed(twiddle_factor_table_3_real));
  assign _zz_4533 = ($signed(_zz_9322) * $signed(twiddle_factor_table_3_imag));
  assign _zz_2613 = ($signed(_zz_2615) - $signed(_zz_9323));
  assign _zz_2614 = ($signed(_zz_2615) + $signed(_zz_9325));
  assign _zz_2616 = 1'b1;
  assign _zz_2617 = 1'b1;
  assign _zz_4534 = ($signed(_zz_9343) * $signed(_zz_667));
  assign _zz_2620 = _zz_9344[15 : 0];
  assign _zz_4535 = ($signed(_zz_9345) * $signed(twiddle_factor_table_4_real));
  assign _zz_4536 = ($signed(_zz_9346) * $signed(twiddle_factor_table_4_imag));
  assign _zz_2618 = ($signed(_zz_2620) - $signed(_zz_9347));
  assign _zz_2619 = ($signed(_zz_2620) + $signed(_zz_9349));
  assign _zz_2621 = 1'b1;
  assign _zz_2622 = 1'b1;
  assign _zz_4537 = ($signed(_zz_9367) * $signed(_zz_669));
  assign _zz_2625 = _zz_9368[15 : 0];
  assign _zz_4538 = ($signed(_zz_9369) * $signed(twiddle_factor_table_5_real));
  assign _zz_4539 = ($signed(_zz_9370) * $signed(twiddle_factor_table_5_imag));
  assign _zz_2623 = ($signed(_zz_2625) - $signed(_zz_9371));
  assign _zz_2624 = ($signed(_zz_2625) + $signed(_zz_9373));
  assign _zz_2626 = 1'b1;
  assign _zz_2627 = 1'b1;
  assign _zz_4540 = ($signed(_zz_9391) * $signed(_zz_671));
  assign _zz_2630 = _zz_9392[15 : 0];
  assign _zz_4541 = ($signed(_zz_9393) * $signed(twiddle_factor_table_6_real));
  assign _zz_4542 = ($signed(_zz_9394) * $signed(twiddle_factor_table_6_imag));
  assign _zz_2628 = ($signed(_zz_2630) - $signed(_zz_9395));
  assign _zz_2629 = ($signed(_zz_2630) + $signed(_zz_9397));
  assign _zz_2631 = 1'b1;
  assign _zz_2632 = 1'b1;
  assign _zz_4543 = ($signed(_zz_9415) * $signed(_zz_681));
  assign _zz_2635 = _zz_9416[15 : 0];
  assign _zz_4544 = ($signed(_zz_9417) * $signed(twiddle_factor_table_3_real));
  assign _zz_4545 = ($signed(_zz_9418) * $signed(twiddle_factor_table_3_imag));
  assign _zz_2633 = ($signed(_zz_2635) - $signed(_zz_9419));
  assign _zz_2634 = ($signed(_zz_2635) + $signed(_zz_9421));
  assign _zz_2636 = 1'b1;
  assign _zz_2637 = 1'b1;
  assign _zz_4546 = ($signed(_zz_9439) * $signed(_zz_683));
  assign _zz_2640 = _zz_9440[15 : 0];
  assign _zz_4547 = ($signed(_zz_9441) * $signed(twiddle_factor_table_4_real));
  assign _zz_4548 = ($signed(_zz_9442) * $signed(twiddle_factor_table_4_imag));
  assign _zz_2638 = ($signed(_zz_2640) - $signed(_zz_9443));
  assign _zz_2639 = ($signed(_zz_2640) + $signed(_zz_9445));
  assign _zz_2641 = 1'b1;
  assign _zz_2642 = 1'b1;
  assign _zz_4549 = ($signed(_zz_9463) * $signed(_zz_685));
  assign _zz_2645 = _zz_9464[15 : 0];
  assign _zz_4550 = ($signed(_zz_9465) * $signed(twiddle_factor_table_5_real));
  assign _zz_4551 = ($signed(_zz_9466) * $signed(twiddle_factor_table_5_imag));
  assign _zz_2643 = ($signed(_zz_2645) - $signed(_zz_9467));
  assign _zz_2644 = ($signed(_zz_2645) + $signed(_zz_9469));
  assign _zz_2646 = 1'b1;
  assign _zz_2647 = 1'b1;
  assign _zz_4552 = ($signed(_zz_9487) * $signed(_zz_687));
  assign _zz_2650 = _zz_9488[15 : 0];
  assign _zz_4553 = ($signed(_zz_9489) * $signed(twiddle_factor_table_6_real));
  assign _zz_4554 = ($signed(_zz_9490) * $signed(twiddle_factor_table_6_imag));
  assign _zz_2648 = ($signed(_zz_2650) - $signed(_zz_9491));
  assign _zz_2649 = ($signed(_zz_2650) + $signed(_zz_9493));
  assign _zz_2651 = 1'b1;
  assign _zz_2652 = 1'b1;
  assign _zz_4555 = ($signed(_zz_9511) * $signed(_zz_697));
  assign _zz_2655 = _zz_9512[15 : 0];
  assign _zz_4556 = ($signed(_zz_9513) * $signed(twiddle_factor_table_3_real));
  assign _zz_4557 = ($signed(_zz_9514) * $signed(twiddle_factor_table_3_imag));
  assign _zz_2653 = ($signed(_zz_2655) - $signed(_zz_9515));
  assign _zz_2654 = ($signed(_zz_2655) + $signed(_zz_9517));
  assign _zz_2656 = 1'b1;
  assign _zz_2657 = 1'b1;
  assign _zz_4558 = ($signed(_zz_9535) * $signed(_zz_699));
  assign _zz_2660 = _zz_9536[15 : 0];
  assign _zz_4559 = ($signed(_zz_9537) * $signed(twiddle_factor_table_4_real));
  assign _zz_4560 = ($signed(_zz_9538) * $signed(twiddle_factor_table_4_imag));
  assign _zz_2658 = ($signed(_zz_2660) - $signed(_zz_9539));
  assign _zz_2659 = ($signed(_zz_2660) + $signed(_zz_9541));
  assign _zz_2661 = 1'b1;
  assign _zz_2662 = 1'b1;
  assign _zz_4561 = ($signed(_zz_9559) * $signed(_zz_701));
  assign _zz_2665 = _zz_9560[15 : 0];
  assign _zz_4562 = ($signed(_zz_9561) * $signed(twiddle_factor_table_5_real));
  assign _zz_4563 = ($signed(_zz_9562) * $signed(twiddle_factor_table_5_imag));
  assign _zz_2663 = ($signed(_zz_2665) - $signed(_zz_9563));
  assign _zz_2664 = ($signed(_zz_2665) + $signed(_zz_9565));
  assign _zz_2666 = 1'b1;
  assign _zz_2667 = 1'b1;
  assign _zz_4564 = ($signed(_zz_9583) * $signed(_zz_703));
  assign _zz_2670 = _zz_9584[15 : 0];
  assign _zz_4565 = ($signed(_zz_9585) * $signed(twiddle_factor_table_6_real));
  assign _zz_4566 = ($signed(_zz_9586) * $signed(twiddle_factor_table_6_imag));
  assign _zz_2668 = ($signed(_zz_2670) - $signed(_zz_9587));
  assign _zz_2669 = ($signed(_zz_2670) + $signed(_zz_9589));
  assign _zz_2671 = 1'b1;
  assign _zz_2672 = 1'b1;
  assign _zz_4567 = ($signed(_zz_9607) * $signed(_zz_713));
  assign _zz_2675 = _zz_9608[15 : 0];
  assign _zz_4568 = ($signed(_zz_9609) * $signed(twiddle_factor_table_3_real));
  assign _zz_4569 = ($signed(_zz_9610) * $signed(twiddle_factor_table_3_imag));
  assign _zz_2673 = ($signed(_zz_2675) - $signed(_zz_9611));
  assign _zz_2674 = ($signed(_zz_2675) + $signed(_zz_9613));
  assign _zz_2676 = 1'b1;
  assign _zz_2677 = 1'b1;
  assign _zz_4570 = ($signed(_zz_9631) * $signed(_zz_715));
  assign _zz_2680 = _zz_9632[15 : 0];
  assign _zz_4571 = ($signed(_zz_9633) * $signed(twiddle_factor_table_4_real));
  assign _zz_4572 = ($signed(_zz_9634) * $signed(twiddle_factor_table_4_imag));
  assign _zz_2678 = ($signed(_zz_2680) - $signed(_zz_9635));
  assign _zz_2679 = ($signed(_zz_2680) + $signed(_zz_9637));
  assign _zz_2681 = 1'b1;
  assign _zz_2682 = 1'b1;
  assign _zz_4573 = ($signed(_zz_9655) * $signed(_zz_717));
  assign _zz_2685 = _zz_9656[15 : 0];
  assign _zz_4574 = ($signed(_zz_9657) * $signed(twiddle_factor_table_5_real));
  assign _zz_4575 = ($signed(_zz_9658) * $signed(twiddle_factor_table_5_imag));
  assign _zz_2683 = ($signed(_zz_2685) - $signed(_zz_9659));
  assign _zz_2684 = ($signed(_zz_2685) + $signed(_zz_9661));
  assign _zz_2686 = 1'b1;
  assign _zz_2687 = 1'b1;
  assign _zz_4576 = ($signed(_zz_9679) * $signed(_zz_719));
  assign _zz_2690 = _zz_9680[15 : 0];
  assign _zz_4577 = ($signed(_zz_9681) * $signed(twiddle_factor_table_6_real));
  assign _zz_4578 = ($signed(_zz_9682) * $signed(twiddle_factor_table_6_imag));
  assign _zz_2688 = ($signed(_zz_2690) - $signed(_zz_9683));
  assign _zz_2689 = ($signed(_zz_2690) + $signed(_zz_9685));
  assign _zz_2691 = 1'b1;
  assign _zz_2692 = 1'b1;
  assign _zz_4579 = ($signed(_zz_9703) * $signed(_zz_729));
  assign _zz_2695 = _zz_9704[15 : 0];
  assign _zz_4580 = ($signed(_zz_9705) * $signed(twiddle_factor_table_3_real));
  assign _zz_4581 = ($signed(_zz_9706) * $signed(twiddle_factor_table_3_imag));
  assign _zz_2693 = ($signed(_zz_2695) - $signed(_zz_9707));
  assign _zz_2694 = ($signed(_zz_2695) + $signed(_zz_9709));
  assign _zz_2696 = 1'b1;
  assign _zz_2697 = 1'b1;
  assign _zz_4582 = ($signed(_zz_9727) * $signed(_zz_731));
  assign _zz_2700 = _zz_9728[15 : 0];
  assign _zz_4583 = ($signed(_zz_9729) * $signed(twiddle_factor_table_4_real));
  assign _zz_4584 = ($signed(_zz_9730) * $signed(twiddle_factor_table_4_imag));
  assign _zz_2698 = ($signed(_zz_2700) - $signed(_zz_9731));
  assign _zz_2699 = ($signed(_zz_2700) + $signed(_zz_9733));
  assign _zz_2701 = 1'b1;
  assign _zz_2702 = 1'b1;
  assign _zz_4585 = ($signed(_zz_9751) * $signed(_zz_733));
  assign _zz_2705 = _zz_9752[15 : 0];
  assign _zz_4586 = ($signed(_zz_9753) * $signed(twiddle_factor_table_5_real));
  assign _zz_4587 = ($signed(_zz_9754) * $signed(twiddle_factor_table_5_imag));
  assign _zz_2703 = ($signed(_zz_2705) - $signed(_zz_9755));
  assign _zz_2704 = ($signed(_zz_2705) + $signed(_zz_9757));
  assign _zz_2706 = 1'b1;
  assign _zz_2707 = 1'b1;
  assign _zz_4588 = ($signed(_zz_9775) * $signed(_zz_735));
  assign _zz_2710 = _zz_9776[15 : 0];
  assign _zz_4589 = ($signed(_zz_9777) * $signed(twiddle_factor_table_6_real));
  assign _zz_4590 = ($signed(_zz_9778) * $signed(twiddle_factor_table_6_imag));
  assign _zz_2708 = ($signed(_zz_2710) - $signed(_zz_9779));
  assign _zz_2709 = ($signed(_zz_2710) + $signed(_zz_9781));
  assign _zz_2711 = 1'b1;
  assign _zz_2712 = 1'b1;
  assign _zz_4591 = ($signed(_zz_9799) * $signed(_zz_745));
  assign _zz_2715 = _zz_9800[15 : 0];
  assign _zz_4592 = ($signed(_zz_9801) * $signed(twiddle_factor_table_3_real));
  assign _zz_4593 = ($signed(_zz_9802) * $signed(twiddle_factor_table_3_imag));
  assign _zz_2713 = ($signed(_zz_2715) - $signed(_zz_9803));
  assign _zz_2714 = ($signed(_zz_2715) + $signed(_zz_9805));
  assign _zz_2716 = 1'b1;
  assign _zz_2717 = 1'b1;
  assign _zz_4594 = ($signed(_zz_9823) * $signed(_zz_747));
  assign _zz_2720 = _zz_9824[15 : 0];
  assign _zz_4595 = ($signed(_zz_9825) * $signed(twiddle_factor_table_4_real));
  assign _zz_4596 = ($signed(_zz_9826) * $signed(twiddle_factor_table_4_imag));
  assign _zz_2718 = ($signed(_zz_2720) - $signed(_zz_9827));
  assign _zz_2719 = ($signed(_zz_2720) + $signed(_zz_9829));
  assign _zz_2721 = 1'b1;
  assign _zz_2722 = 1'b1;
  assign _zz_4597 = ($signed(_zz_9847) * $signed(_zz_749));
  assign _zz_2725 = _zz_9848[15 : 0];
  assign _zz_4598 = ($signed(_zz_9849) * $signed(twiddle_factor_table_5_real));
  assign _zz_4599 = ($signed(_zz_9850) * $signed(twiddle_factor_table_5_imag));
  assign _zz_2723 = ($signed(_zz_2725) - $signed(_zz_9851));
  assign _zz_2724 = ($signed(_zz_2725) + $signed(_zz_9853));
  assign _zz_2726 = 1'b1;
  assign _zz_2727 = 1'b1;
  assign _zz_4600 = ($signed(_zz_9871) * $signed(_zz_751));
  assign _zz_2730 = _zz_9872[15 : 0];
  assign _zz_4601 = ($signed(_zz_9873) * $signed(twiddle_factor_table_6_real));
  assign _zz_4602 = ($signed(_zz_9874) * $signed(twiddle_factor_table_6_imag));
  assign _zz_2728 = ($signed(_zz_2730) - $signed(_zz_9875));
  assign _zz_2729 = ($signed(_zz_2730) + $signed(_zz_9877));
  assign _zz_2731 = 1'b1;
  assign _zz_2732 = 1'b1;
  assign _zz_4603 = ($signed(_zz_9895) * $signed(_zz_761));
  assign _zz_2735 = _zz_9896[15 : 0];
  assign _zz_4604 = ($signed(_zz_9897) * $signed(twiddle_factor_table_3_real));
  assign _zz_4605 = ($signed(_zz_9898) * $signed(twiddle_factor_table_3_imag));
  assign _zz_2733 = ($signed(_zz_2735) - $signed(_zz_9899));
  assign _zz_2734 = ($signed(_zz_2735) + $signed(_zz_9901));
  assign _zz_2736 = 1'b1;
  assign _zz_2737 = 1'b1;
  assign _zz_4606 = ($signed(_zz_9919) * $signed(_zz_763));
  assign _zz_2740 = _zz_9920[15 : 0];
  assign _zz_4607 = ($signed(_zz_9921) * $signed(twiddle_factor_table_4_real));
  assign _zz_4608 = ($signed(_zz_9922) * $signed(twiddle_factor_table_4_imag));
  assign _zz_2738 = ($signed(_zz_2740) - $signed(_zz_9923));
  assign _zz_2739 = ($signed(_zz_2740) + $signed(_zz_9925));
  assign _zz_2741 = 1'b1;
  assign _zz_2742 = 1'b1;
  assign _zz_4609 = ($signed(_zz_9943) * $signed(_zz_765));
  assign _zz_2745 = _zz_9944[15 : 0];
  assign _zz_4610 = ($signed(_zz_9945) * $signed(twiddle_factor_table_5_real));
  assign _zz_4611 = ($signed(_zz_9946) * $signed(twiddle_factor_table_5_imag));
  assign _zz_2743 = ($signed(_zz_2745) - $signed(_zz_9947));
  assign _zz_2744 = ($signed(_zz_2745) + $signed(_zz_9949));
  assign _zz_2746 = 1'b1;
  assign _zz_2747 = 1'b1;
  assign _zz_4612 = ($signed(_zz_9967) * $signed(_zz_767));
  assign _zz_2750 = _zz_9968[15 : 0];
  assign _zz_4613 = ($signed(_zz_9969) * $signed(twiddle_factor_table_6_real));
  assign _zz_4614 = ($signed(_zz_9970) * $signed(twiddle_factor_table_6_imag));
  assign _zz_2748 = ($signed(_zz_2750) - $signed(_zz_9971));
  assign _zz_2749 = ($signed(_zz_2750) + $signed(_zz_9973));
  assign _zz_2751 = 1'b1;
  assign _zz_2752 = 1'b1;
  assign _zz_4615 = ($signed(_zz_9991) * $signed(_zz_785));
  assign _zz_2755 = _zz_9992[15 : 0];
  assign _zz_4616 = ($signed(_zz_9993) * $signed(twiddle_factor_table_7_real));
  assign _zz_4617 = ($signed(_zz_9994) * $signed(twiddle_factor_table_7_imag));
  assign _zz_2753 = ($signed(_zz_2755) - $signed(_zz_9995));
  assign _zz_2754 = ($signed(_zz_2755) + $signed(_zz_9997));
  assign _zz_2756 = 1'b1;
  assign _zz_2757 = 1'b1;
  assign _zz_4618 = ($signed(_zz_10015) * $signed(_zz_787));
  assign _zz_2760 = _zz_10016[15 : 0];
  assign _zz_4619 = ($signed(_zz_10017) * $signed(twiddle_factor_table_8_real));
  assign _zz_4620 = ($signed(_zz_10018) * $signed(twiddle_factor_table_8_imag));
  assign _zz_2758 = ($signed(_zz_2760) - $signed(_zz_10019));
  assign _zz_2759 = ($signed(_zz_2760) + $signed(_zz_10021));
  assign _zz_2761 = 1'b1;
  assign _zz_2762 = 1'b1;
  assign _zz_4621 = ($signed(_zz_10039) * $signed(_zz_789));
  assign _zz_2765 = _zz_10040[15 : 0];
  assign _zz_4622 = ($signed(_zz_10041) * $signed(twiddle_factor_table_9_real));
  assign _zz_4623 = ($signed(_zz_10042) * $signed(twiddle_factor_table_9_imag));
  assign _zz_2763 = ($signed(_zz_2765) - $signed(_zz_10043));
  assign _zz_2764 = ($signed(_zz_2765) + $signed(_zz_10045));
  assign _zz_2766 = 1'b1;
  assign _zz_2767 = 1'b1;
  assign _zz_4624 = ($signed(_zz_10063) * $signed(_zz_791));
  assign _zz_2770 = _zz_10064[15 : 0];
  assign _zz_4625 = ($signed(_zz_10065) * $signed(twiddle_factor_table_10_real));
  assign _zz_4626 = ($signed(_zz_10066) * $signed(twiddle_factor_table_10_imag));
  assign _zz_2768 = ($signed(_zz_2770) - $signed(_zz_10067));
  assign _zz_2769 = ($signed(_zz_2770) + $signed(_zz_10069));
  assign _zz_2771 = 1'b1;
  assign _zz_2772 = 1'b1;
  assign _zz_4627 = ($signed(_zz_10087) * $signed(_zz_793));
  assign _zz_2775 = _zz_10088[15 : 0];
  assign _zz_4628 = ($signed(_zz_10089) * $signed(twiddle_factor_table_11_real));
  assign _zz_4629 = ($signed(_zz_10090) * $signed(twiddle_factor_table_11_imag));
  assign _zz_2773 = ($signed(_zz_2775) - $signed(_zz_10091));
  assign _zz_2774 = ($signed(_zz_2775) + $signed(_zz_10093));
  assign _zz_2776 = 1'b1;
  assign _zz_2777 = 1'b1;
  assign _zz_4630 = ($signed(_zz_10111) * $signed(_zz_795));
  assign _zz_2780 = _zz_10112[15 : 0];
  assign _zz_4631 = ($signed(_zz_10113) * $signed(twiddle_factor_table_12_real));
  assign _zz_4632 = ($signed(_zz_10114) * $signed(twiddle_factor_table_12_imag));
  assign _zz_2778 = ($signed(_zz_2780) - $signed(_zz_10115));
  assign _zz_2779 = ($signed(_zz_2780) + $signed(_zz_10117));
  assign _zz_2781 = 1'b1;
  assign _zz_2782 = 1'b1;
  assign _zz_4633 = ($signed(_zz_10135) * $signed(_zz_797));
  assign _zz_2785 = _zz_10136[15 : 0];
  assign _zz_4634 = ($signed(_zz_10137) * $signed(twiddle_factor_table_13_real));
  assign _zz_4635 = ($signed(_zz_10138) * $signed(twiddle_factor_table_13_imag));
  assign _zz_2783 = ($signed(_zz_2785) - $signed(_zz_10139));
  assign _zz_2784 = ($signed(_zz_2785) + $signed(_zz_10141));
  assign _zz_2786 = 1'b1;
  assign _zz_2787 = 1'b1;
  assign _zz_4636 = ($signed(_zz_10159) * $signed(_zz_799));
  assign _zz_2790 = _zz_10160[15 : 0];
  assign _zz_4637 = ($signed(_zz_10161) * $signed(twiddle_factor_table_14_real));
  assign _zz_4638 = ($signed(_zz_10162) * $signed(twiddle_factor_table_14_imag));
  assign _zz_2788 = ($signed(_zz_2790) - $signed(_zz_10163));
  assign _zz_2789 = ($signed(_zz_2790) + $signed(_zz_10165));
  assign _zz_2791 = 1'b1;
  assign _zz_2792 = 1'b1;
  assign _zz_4639 = ($signed(_zz_10183) * $signed(_zz_817));
  assign _zz_2795 = _zz_10184[15 : 0];
  assign _zz_4640 = ($signed(_zz_10185) * $signed(twiddle_factor_table_7_real));
  assign _zz_4641 = ($signed(_zz_10186) * $signed(twiddle_factor_table_7_imag));
  assign _zz_2793 = ($signed(_zz_2795) - $signed(_zz_10187));
  assign _zz_2794 = ($signed(_zz_2795) + $signed(_zz_10189));
  assign _zz_2796 = 1'b1;
  assign _zz_2797 = 1'b1;
  assign _zz_4642 = ($signed(_zz_10207) * $signed(_zz_819));
  assign _zz_2800 = _zz_10208[15 : 0];
  assign _zz_4643 = ($signed(_zz_10209) * $signed(twiddle_factor_table_8_real));
  assign _zz_4644 = ($signed(_zz_10210) * $signed(twiddle_factor_table_8_imag));
  assign _zz_2798 = ($signed(_zz_2800) - $signed(_zz_10211));
  assign _zz_2799 = ($signed(_zz_2800) + $signed(_zz_10213));
  assign _zz_2801 = 1'b1;
  assign _zz_2802 = 1'b1;
  assign _zz_4645 = ($signed(_zz_10231) * $signed(_zz_821));
  assign _zz_2805 = _zz_10232[15 : 0];
  assign _zz_4646 = ($signed(_zz_10233) * $signed(twiddle_factor_table_9_real));
  assign _zz_4647 = ($signed(_zz_10234) * $signed(twiddle_factor_table_9_imag));
  assign _zz_2803 = ($signed(_zz_2805) - $signed(_zz_10235));
  assign _zz_2804 = ($signed(_zz_2805) + $signed(_zz_10237));
  assign _zz_2806 = 1'b1;
  assign _zz_2807 = 1'b1;
  assign _zz_4648 = ($signed(_zz_10255) * $signed(_zz_823));
  assign _zz_2810 = _zz_10256[15 : 0];
  assign _zz_4649 = ($signed(_zz_10257) * $signed(twiddle_factor_table_10_real));
  assign _zz_4650 = ($signed(_zz_10258) * $signed(twiddle_factor_table_10_imag));
  assign _zz_2808 = ($signed(_zz_2810) - $signed(_zz_10259));
  assign _zz_2809 = ($signed(_zz_2810) + $signed(_zz_10261));
  assign _zz_2811 = 1'b1;
  assign _zz_2812 = 1'b1;
  assign _zz_4651 = ($signed(_zz_10279) * $signed(_zz_825));
  assign _zz_2815 = _zz_10280[15 : 0];
  assign _zz_4652 = ($signed(_zz_10281) * $signed(twiddle_factor_table_11_real));
  assign _zz_4653 = ($signed(_zz_10282) * $signed(twiddle_factor_table_11_imag));
  assign _zz_2813 = ($signed(_zz_2815) - $signed(_zz_10283));
  assign _zz_2814 = ($signed(_zz_2815) + $signed(_zz_10285));
  assign _zz_2816 = 1'b1;
  assign _zz_2817 = 1'b1;
  assign _zz_4654 = ($signed(_zz_10303) * $signed(_zz_827));
  assign _zz_2820 = _zz_10304[15 : 0];
  assign _zz_4655 = ($signed(_zz_10305) * $signed(twiddle_factor_table_12_real));
  assign _zz_4656 = ($signed(_zz_10306) * $signed(twiddle_factor_table_12_imag));
  assign _zz_2818 = ($signed(_zz_2820) - $signed(_zz_10307));
  assign _zz_2819 = ($signed(_zz_2820) + $signed(_zz_10309));
  assign _zz_2821 = 1'b1;
  assign _zz_2822 = 1'b1;
  assign _zz_4657 = ($signed(_zz_10327) * $signed(_zz_829));
  assign _zz_2825 = _zz_10328[15 : 0];
  assign _zz_4658 = ($signed(_zz_10329) * $signed(twiddle_factor_table_13_real));
  assign _zz_4659 = ($signed(_zz_10330) * $signed(twiddle_factor_table_13_imag));
  assign _zz_2823 = ($signed(_zz_2825) - $signed(_zz_10331));
  assign _zz_2824 = ($signed(_zz_2825) + $signed(_zz_10333));
  assign _zz_2826 = 1'b1;
  assign _zz_2827 = 1'b1;
  assign _zz_4660 = ($signed(_zz_10351) * $signed(_zz_831));
  assign _zz_2830 = _zz_10352[15 : 0];
  assign _zz_4661 = ($signed(_zz_10353) * $signed(twiddle_factor_table_14_real));
  assign _zz_4662 = ($signed(_zz_10354) * $signed(twiddle_factor_table_14_imag));
  assign _zz_2828 = ($signed(_zz_2830) - $signed(_zz_10355));
  assign _zz_2829 = ($signed(_zz_2830) + $signed(_zz_10357));
  assign _zz_2831 = 1'b1;
  assign _zz_2832 = 1'b1;
  assign _zz_4663 = ($signed(_zz_10375) * $signed(_zz_849));
  assign _zz_2835 = _zz_10376[15 : 0];
  assign _zz_4664 = ($signed(_zz_10377) * $signed(twiddle_factor_table_7_real));
  assign _zz_4665 = ($signed(_zz_10378) * $signed(twiddle_factor_table_7_imag));
  assign _zz_2833 = ($signed(_zz_2835) - $signed(_zz_10379));
  assign _zz_2834 = ($signed(_zz_2835) + $signed(_zz_10381));
  assign _zz_2836 = 1'b1;
  assign _zz_2837 = 1'b1;
  assign _zz_4666 = ($signed(_zz_10399) * $signed(_zz_851));
  assign _zz_2840 = _zz_10400[15 : 0];
  assign _zz_4667 = ($signed(_zz_10401) * $signed(twiddle_factor_table_8_real));
  assign _zz_4668 = ($signed(_zz_10402) * $signed(twiddle_factor_table_8_imag));
  assign _zz_2838 = ($signed(_zz_2840) - $signed(_zz_10403));
  assign _zz_2839 = ($signed(_zz_2840) + $signed(_zz_10405));
  assign _zz_2841 = 1'b1;
  assign _zz_2842 = 1'b1;
  assign _zz_4669 = ($signed(_zz_10423) * $signed(_zz_853));
  assign _zz_2845 = _zz_10424[15 : 0];
  assign _zz_4670 = ($signed(_zz_10425) * $signed(twiddle_factor_table_9_real));
  assign _zz_4671 = ($signed(_zz_10426) * $signed(twiddle_factor_table_9_imag));
  assign _zz_2843 = ($signed(_zz_2845) - $signed(_zz_10427));
  assign _zz_2844 = ($signed(_zz_2845) + $signed(_zz_10429));
  assign _zz_2846 = 1'b1;
  assign _zz_2847 = 1'b1;
  assign _zz_4672 = ($signed(_zz_10447) * $signed(_zz_855));
  assign _zz_2850 = _zz_10448[15 : 0];
  assign _zz_4673 = ($signed(_zz_10449) * $signed(twiddle_factor_table_10_real));
  assign _zz_4674 = ($signed(_zz_10450) * $signed(twiddle_factor_table_10_imag));
  assign _zz_2848 = ($signed(_zz_2850) - $signed(_zz_10451));
  assign _zz_2849 = ($signed(_zz_2850) + $signed(_zz_10453));
  assign _zz_2851 = 1'b1;
  assign _zz_2852 = 1'b1;
  assign _zz_4675 = ($signed(_zz_10471) * $signed(_zz_857));
  assign _zz_2855 = _zz_10472[15 : 0];
  assign _zz_4676 = ($signed(_zz_10473) * $signed(twiddle_factor_table_11_real));
  assign _zz_4677 = ($signed(_zz_10474) * $signed(twiddle_factor_table_11_imag));
  assign _zz_2853 = ($signed(_zz_2855) - $signed(_zz_10475));
  assign _zz_2854 = ($signed(_zz_2855) + $signed(_zz_10477));
  assign _zz_2856 = 1'b1;
  assign _zz_2857 = 1'b1;
  assign _zz_4678 = ($signed(_zz_10495) * $signed(_zz_859));
  assign _zz_2860 = _zz_10496[15 : 0];
  assign _zz_4679 = ($signed(_zz_10497) * $signed(twiddle_factor_table_12_real));
  assign _zz_4680 = ($signed(_zz_10498) * $signed(twiddle_factor_table_12_imag));
  assign _zz_2858 = ($signed(_zz_2860) - $signed(_zz_10499));
  assign _zz_2859 = ($signed(_zz_2860) + $signed(_zz_10501));
  assign _zz_2861 = 1'b1;
  assign _zz_2862 = 1'b1;
  assign _zz_4681 = ($signed(_zz_10519) * $signed(_zz_861));
  assign _zz_2865 = _zz_10520[15 : 0];
  assign _zz_4682 = ($signed(_zz_10521) * $signed(twiddle_factor_table_13_real));
  assign _zz_4683 = ($signed(_zz_10522) * $signed(twiddle_factor_table_13_imag));
  assign _zz_2863 = ($signed(_zz_2865) - $signed(_zz_10523));
  assign _zz_2864 = ($signed(_zz_2865) + $signed(_zz_10525));
  assign _zz_2866 = 1'b1;
  assign _zz_2867 = 1'b1;
  assign _zz_4684 = ($signed(_zz_10543) * $signed(_zz_863));
  assign _zz_2870 = _zz_10544[15 : 0];
  assign _zz_4685 = ($signed(_zz_10545) * $signed(twiddle_factor_table_14_real));
  assign _zz_4686 = ($signed(_zz_10546) * $signed(twiddle_factor_table_14_imag));
  assign _zz_2868 = ($signed(_zz_2870) - $signed(_zz_10547));
  assign _zz_2869 = ($signed(_zz_2870) + $signed(_zz_10549));
  assign _zz_2871 = 1'b1;
  assign _zz_2872 = 1'b1;
  assign _zz_4687 = ($signed(_zz_10567) * $signed(_zz_881));
  assign _zz_2875 = _zz_10568[15 : 0];
  assign _zz_4688 = ($signed(_zz_10569) * $signed(twiddle_factor_table_7_real));
  assign _zz_4689 = ($signed(_zz_10570) * $signed(twiddle_factor_table_7_imag));
  assign _zz_2873 = ($signed(_zz_2875) - $signed(_zz_10571));
  assign _zz_2874 = ($signed(_zz_2875) + $signed(_zz_10573));
  assign _zz_2876 = 1'b1;
  assign _zz_2877 = 1'b1;
  assign _zz_4690 = ($signed(_zz_10591) * $signed(_zz_883));
  assign _zz_2880 = _zz_10592[15 : 0];
  assign _zz_4691 = ($signed(_zz_10593) * $signed(twiddle_factor_table_8_real));
  assign _zz_4692 = ($signed(_zz_10594) * $signed(twiddle_factor_table_8_imag));
  assign _zz_2878 = ($signed(_zz_2880) - $signed(_zz_10595));
  assign _zz_2879 = ($signed(_zz_2880) + $signed(_zz_10597));
  assign _zz_2881 = 1'b1;
  assign _zz_2882 = 1'b1;
  assign _zz_4693 = ($signed(_zz_10615) * $signed(_zz_885));
  assign _zz_2885 = _zz_10616[15 : 0];
  assign _zz_4694 = ($signed(_zz_10617) * $signed(twiddle_factor_table_9_real));
  assign _zz_4695 = ($signed(_zz_10618) * $signed(twiddle_factor_table_9_imag));
  assign _zz_2883 = ($signed(_zz_2885) - $signed(_zz_10619));
  assign _zz_2884 = ($signed(_zz_2885) + $signed(_zz_10621));
  assign _zz_2886 = 1'b1;
  assign _zz_2887 = 1'b1;
  assign _zz_4696 = ($signed(_zz_10639) * $signed(_zz_887));
  assign _zz_2890 = _zz_10640[15 : 0];
  assign _zz_4697 = ($signed(_zz_10641) * $signed(twiddle_factor_table_10_real));
  assign _zz_4698 = ($signed(_zz_10642) * $signed(twiddle_factor_table_10_imag));
  assign _zz_2888 = ($signed(_zz_2890) - $signed(_zz_10643));
  assign _zz_2889 = ($signed(_zz_2890) + $signed(_zz_10645));
  assign _zz_2891 = 1'b1;
  assign _zz_2892 = 1'b1;
  assign _zz_4699 = ($signed(_zz_10663) * $signed(_zz_889));
  assign _zz_2895 = _zz_10664[15 : 0];
  assign _zz_4700 = ($signed(_zz_10665) * $signed(twiddle_factor_table_11_real));
  assign _zz_4701 = ($signed(_zz_10666) * $signed(twiddle_factor_table_11_imag));
  assign _zz_2893 = ($signed(_zz_2895) - $signed(_zz_10667));
  assign _zz_2894 = ($signed(_zz_2895) + $signed(_zz_10669));
  assign _zz_2896 = 1'b1;
  assign _zz_2897 = 1'b1;
  assign _zz_4702 = ($signed(_zz_10687) * $signed(_zz_891));
  assign _zz_2900 = _zz_10688[15 : 0];
  assign _zz_4703 = ($signed(_zz_10689) * $signed(twiddle_factor_table_12_real));
  assign _zz_4704 = ($signed(_zz_10690) * $signed(twiddle_factor_table_12_imag));
  assign _zz_2898 = ($signed(_zz_2900) - $signed(_zz_10691));
  assign _zz_2899 = ($signed(_zz_2900) + $signed(_zz_10693));
  assign _zz_2901 = 1'b1;
  assign _zz_2902 = 1'b1;
  assign _zz_4705 = ($signed(_zz_10711) * $signed(_zz_893));
  assign _zz_2905 = _zz_10712[15 : 0];
  assign _zz_4706 = ($signed(_zz_10713) * $signed(twiddle_factor_table_13_real));
  assign _zz_4707 = ($signed(_zz_10714) * $signed(twiddle_factor_table_13_imag));
  assign _zz_2903 = ($signed(_zz_2905) - $signed(_zz_10715));
  assign _zz_2904 = ($signed(_zz_2905) + $signed(_zz_10717));
  assign _zz_2906 = 1'b1;
  assign _zz_2907 = 1'b1;
  assign _zz_4708 = ($signed(_zz_10735) * $signed(_zz_895));
  assign _zz_2910 = _zz_10736[15 : 0];
  assign _zz_4709 = ($signed(_zz_10737) * $signed(twiddle_factor_table_14_real));
  assign _zz_4710 = ($signed(_zz_10738) * $signed(twiddle_factor_table_14_imag));
  assign _zz_2908 = ($signed(_zz_2910) - $signed(_zz_10739));
  assign _zz_2909 = ($signed(_zz_2910) + $signed(_zz_10741));
  assign _zz_2911 = 1'b1;
  assign _zz_2912 = 1'b1;
  assign _zz_4711 = ($signed(_zz_10759) * $signed(_zz_913));
  assign _zz_2915 = _zz_10760[15 : 0];
  assign _zz_4712 = ($signed(_zz_10761) * $signed(twiddle_factor_table_7_real));
  assign _zz_4713 = ($signed(_zz_10762) * $signed(twiddle_factor_table_7_imag));
  assign _zz_2913 = ($signed(_zz_2915) - $signed(_zz_10763));
  assign _zz_2914 = ($signed(_zz_2915) + $signed(_zz_10765));
  assign _zz_2916 = 1'b1;
  assign _zz_2917 = 1'b1;
  assign _zz_4714 = ($signed(_zz_10783) * $signed(_zz_915));
  assign _zz_2920 = _zz_10784[15 : 0];
  assign _zz_4715 = ($signed(_zz_10785) * $signed(twiddle_factor_table_8_real));
  assign _zz_4716 = ($signed(_zz_10786) * $signed(twiddle_factor_table_8_imag));
  assign _zz_2918 = ($signed(_zz_2920) - $signed(_zz_10787));
  assign _zz_2919 = ($signed(_zz_2920) + $signed(_zz_10789));
  assign _zz_2921 = 1'b1;
  assign _zz_2922 = 1'b1;
  assign _zz_4717 = ($signed(_zz_10807) * $signed(_zz_917));
  assign _zz_2925 = _zz_10808[15 : 0];
  assign _zz_4718 = ($signed(_zz_10809) * $signed(twiddle_factor_table_9_real));
  assign _zz_4719 = ($signed(_zz_10810) * $signed(twiddle_factor_table_9_imag));
  assign _zz_2923 = ($signed(_zz_2925) - $signed(_zz_10811));
  assign _zz_2924 = ($signed(_zz_2925) + $signed(_zz_10813));
  assign _zz_2926 = 1'b1;
  assign _zz_2927 = 1'b1;
  assign _zz_4720 = ($signed(_zz_10831) * $signed(_zz_919));
  assign _zz_2930 = _zz_10832[15 : 0];
  assign _zz_4721 = ($signed(_zz_10833) * $signed(twiddle_factor_table_10_real));
  assign _zz_4722 = ($signed(_zz_10834) * $signed(twiddle_factor_table_10_imag));
  assign _zz_2928 = ($signed(_zz_2930) - $signed(_zz_10835));
  assign _zz_2929 = ($signed(_zz_2930) + $signed(_zz_10837));
  assign _zz_2931 = 1'b1;
  assign _zz_2932 = 1'b1;
  assign _zz_4723 = ($signed(_zz_10855) * $signed(_zz_921));
  assign _zz_2935 = _zz_10856[15 : 0];
  assign _zz_4724 = ($signed(_zz_10857) * $signed(twiddle_factor_table_11_real));
  assign _zz_4725 = ($signed(_zz_10858) * $signed(twiddle_factor_table_11_imag));
  assign _zz_2933 = ($signed(_zz_2935) - $signed(_zz_10859));
  assign _zz_2934 = ($signed(_zz_2935) + $signed(_zz_10861));
  assign _zz_2936 = 1'b1;
  assign _zz_2937 = 1'b1;
  assign _zz_4726 = ($signed(_zz_10879) * $signed(_zz_923));
  assign _zz_2940 = _zz_10880[15 : 0];
  assign _zz_4727 = ($signed(_zz_10881) * $signed(twiddle_factor_table_12_real));
  assign _zz_4728 = ($signed(_zz_10882) * $signed(twiddle_factor_table_12_imag));
  assign _zz_2938 = ($signed(_zz_2940) - $signed(_zz_10883));
  assign _zz_2939 = ($signed(_zz_2940) + $signed(_zz_10885));
  assign _zz_2941 = 1'b1;
  assign _zz_2942 = 1'b1;
  assign _zz_4729 = ($signed(_zz_10903) * $signed(_zz_925));
  assign _zz_2945 = _zz_10904[15 : 0];
  assign _zz_4730 = ($signed(_zz_10905) * $signed(twiddle_factor_table_13_real));
  assign _zz_4731 = ($signed(_zz_10906) * $signed(twiddle_factor_table_13_imag));
  assign _zz_2943 = ($signed(_zz_2945) - $signed(_zz_10907));
  assign _zz_2944 = ($signed(_zz_2945) + $signed(_zz_10909));
  assign _zz_2946 = 1'b1;
  assign _zz_2947 = 1'b1;
  assign _zz_4732 = ($signed(_zz_10927) * $signed(_zz_927));
  assign _zz_2950 = _zz_10928[15 : 0];
  assign _zz_4733 = ($signed(_zz_10929) * $signed(twiddle_factor_table_14_real));
  assign _zz_4734 = ($signed(_zz_10930) * $signed(twiddle_factor_table_14_imag));
  assign _zz_2948 = ($signed(_zz_2950) - $signed(_zz_10931));
  assign _zz_2949 = ($signed(_zz_2950) + $signed(_zz_10933));
  assign _zz_2951 = 1'b1;
  assign _zz_2952 = 1'b1;
  assign _zz_4735 = ($signed(_zz_10951) * $signed(_zz_945));
  assign _zz_2955 = _zz_10952[15 : 0];
  assign _zz_4736 = ($signed(_zz_10953) * $signed(twiddle_factor_table_7_real));
  assign _zz_4737 = ($signed(_zz_10954) * $signed(twiddle_factor_table_7_imag));
  assign _zz_2953 = ($signed(_zz_2955) - $signed(_zz_10955));
  assign _zz_2954 = ($signed(_zz_2955) + $signed(_zz_10957));
  assign _zz_2956 = 1'b1;
  assign _zz_2957 = 1'b1;
  assign _zz_4738 = ($signed(_zz_10975) * $signed(_zz_947));
  assign _zz_2960 = _zz_10976[15 : 0];
  assign _zz_4739 = ($signed(_zz_10977) * $signed(twiddle_factor_table_8_real));
  assign _zz_4740 = ($signed(_zz_10978) * $signed(twiddle_factor_table_8_imag));
  assign _zz_2958 = ($signed(_zz_2960) - $signed(_zz_10979));
  assign _zz_2959 = ($signed(_zz_2960) + $signed(_zz_10981));
  assign _zz_2961 = 1'b1;
  assign _zz_2962 = 1'b1;
  assign _zz_4741 = ($signed(_zz_10999) * $signed(_zz_949));
  assign _zz_2965 = _zz_11000[15 : 0];
  assign _zz_4742 = ($signed(_zz_11001) * $signed(twiddle_factor_table_9_real));
  assign _zz_4743 = ($signed(_zz_11002) * $signed(twiddle_factor_table_9_imag));
  assign _zz_2963 = ($signed(_zz_2965) - $signed(_zz_11003));
  assign _zz_2964 = ($signed(_zz_2965) + $signed(_zz_11005));
  assign _zz_2966 = 1'b1;
  assign _zz_2967 = 1'b1;
  assign _zz_4744 = ($signed(_zz_11023) * $signed(_zz_951));
  assign _zz_2970 = _zz_11024[15 : 0];
  assign _zz_4745 = ($signed(_zz_11025) * $signed(twiddle_factor_table_10_real));
  assign _zz_4746 = ($signed(_zz_11026) * $signed(twiddle_factor_table_10_imag));
  assign _zz_2968 = ($signed(_zz_2970) - $signed(_zz_11027));
  assign _zz_2969 = ($signed(_zz_2970) + $signed(_zz_11029));
  assign _zz_2971 = 1'b1;
  assign _zz_2972 = 1'b1;
  assign _zz_4747 = ($signed(_zz_11047) * $signed(_zz_953));
  assign _zz_2975 = _zz_11048[15 : 0];
  assign _zz_4748 = ($signed(_zz_11049) * $signed(twiddle_factor_table_11_real));
  assign _zz_4749 = ($signed(_zz_11050) * $signed(twiddle_factor_table_11_imag));
  assign _zz_2973 = ($signed(_zz_2975) - $signed(_zz_11051));
  assign _zz_2974 = ($signed(_zz_2975) + $signed(_zz_11053));
  assign _zz_2976 = 1'b1;
  assign _zz_2977 = 1'b1;
  assign _zz_4750 = ($signed(_zz_11071) * $signed(_zz_955));
  assign _zz_2980 = _zz_11072[15 : 0];
  assign _zz_4751 = ($signed(_zz_11073) * $signed(twiddle_factor_table_12_real));
  assign _zz_4752 = ($signed(_zz_11074) * $signed(twiddle_factor_table_12_imag));
  assign _zz_2978 = ($signed(_zz_2980) - $signed(_zz_11075));
  assign _zz_2979 = ($signed(_zz_2980) + $signed(_zz_11077));
  assign _zz_2981 = 1'b1;
  assign _zz_2982 = 1'b1;
  assign _zz_4753 = ($signed(_zz_11095) * $signed(_zz_957));
  assign _zz_2985 = _zz_11096[15 : 0];
  assign _zz_4754 = ($signed(_zz_11097) * $signed(twiddle_factor_table_13_real));
  assign _zz_4755 = ($signed(_zz_11098) * $signed(twiddle_factor_table_13_imag));
  assign _zz_2983 = ($signed(_zz_2985) - $signed(_zz_11099));
  assign _zz_2984 = ($signed(_zz_2985) + $signed(_zz_11101));
  assign _zz_2986 = 1'b1;
  assign _zz_2987 = 1'b1;
  assign _zz_4756 = ($signed(_zz_11119) * $signed(_zz_959));
  assign _zz_2990 = _zz_11120[15 : 0];
  assign _zz_4757 = ($signed(_zz_11121) * $signed(twiddle_factor_table_14_real));
  assign _zz_4758 = ($signed(_zz_11122) * $signed(twiddle_factor_table_14_imag));
  assign _zz_2988 = ($signed(_zz_2990) - $signed(_zz_11123));
  assign _zz_2989 = ($signed(_zz_2990) + $signed(_zz_11125));
  assign _zz_2991 = 1'b1;
  assign _zz_2992 = 1'b1;
  assign _zz_4759 = ($signed(_zz_11143) * $signed(_zz_977));
  assign _zz_2995 = _zz_11144[15 : 0];
  assign _zz_4760 = ($signed(_zz_11145) * $signed(twiddle_factor_table_7_real));
  assign _zz_4761 = ($signed(_zz_11146) * $signed(twiddle_factor_table_7_imag));
  assign _zz_2993 = ($signed(_zz_2995) - $signed(_zz_11147));
  assign _zz_2994 = ($signed(_zz_2995) + $signed(_zz_11149));
  assign _zz_2996 = 1'b1;
  assign _zz_2997 = 1'b1;
  assign _zz_4762 = ($signed(_zz_11167) * $signed(_zz_979));
  assign _zz_3000 = _zz_11168[15 : 0];
  assign _zz_4763 = ($signed(_zz_11169) * $signed(twiddle_factor_table_8_real));
  assign _zz_4764 = ($signed(_zz_11170) * $signed(twiddle_factor_table_8_imag));
  assign _zz_2998 = ($signed(_zz_3000) - $signed(_zz_11171));
  assign _zz_2999 = ($signed(_zz_3000) + $signed(_zz_11173));
  assign _zz_3001 = 1'b1;
  assign _zz_3002 = 1'b1;
  assign _zz_4765 = ($signed(_zz_11191) * $signed(_zz_981));
  assign _zz_3005 = _zz_11192[15 : 0];
  assign _zz_4766 = ($signed(_zz_11193) * $signed(twiddle_factor_table_9_real));
  assign _zz_4767 = ($signed(_zz_11194) * $signed(twiddle_factor_table_9_imag));
  assign _zz_3003 = ($signed(_zz_3005) - $signed(_zz_11195));
  assign _zz_3004 = ($signed(_zz_3005) + $signed(_zz_11197));
  assign _zz_3006 = 1'b1;
  assign _zz_3007 = 1'b1;
  assign _zz_4768 = ($signed(_zz_11215) * $signed(_zz_983));
  assign _zz_3010 = _zz_11216[15 : 0];
  assign _zz_4769 = ($signed(_zz_11217) * $signed(twiddle_factor_table_10_real));
  assign _zz_4770 = ($signed(_zz_11218) * $signed(twiddle_factor_table_10_imag));
  assign _zz_3008 = ($signed(_zz_3010) - $signed(_zz_11219));
  assign _zz_3009 = ($signed(_zz_3010) + $signed(_zz_11221));
  assign _zz_3011 = 1'b1;
  assign _zz_3012 = 1'b1;
  assign _zz_4771 = ($signed(_zz_11239) * $signed(_zz_985));
  assign _zz_3015 = _zz_11240[15 : 0];
  assign _zz_4772 = ($signed(_zz_11241) * $signed(twiddle_factor_table_11_real));
  assign _zz_4773 = ($signed(_zz_11242) * $signed(twiddle_factor_table_11_imag));
  assign _zz_3013 = ($signed(_zz_3015) - $signed(_zz_11243));
  assign _zz_3014 = ($signed(_zz_3015) + $signed(_zz_11245));
  assign _zz_3016 = 1'b1;
  assign _zz_3017 = 1'b1;
  assign _zz_4774 = ($signed(_zz_11263) * $signed(_zz_987));
  assign _zz_3020 = _zz_11264[15 : 0];
  assign _zz_4775 = ($signed(_zz_11265) * $signed(twiddle_factor_table_12_real));
  assign _zz_4776 = ($signed(_zz_11266) * $signed(twiddle_factor_table_12_imag));
  assign _zz_3018 = ($signed(_zz_3020) - $signed(_zz_11267));
  assign _zz_3019 = ($signed(_zz_3020) + $signed(_zz_11269));
  assign _zz_3021 = 1'b1;
  assign _zz_3022 = 1'b1;
  assign _zz_4777 = ($signed(_zz_11287) * $signed(_zz_989));
  assign _zz_3025 = _zz_11288[15 : 0];
  assign _zz_4778 = ($signed(_zz_11289) * $signed(twiddle_factor_table_13_real));
  assign _zz_4779 = ($signed(_zz_11290) * $signed(twiddle_factor_table_13_imag));
  assign _zz_3023 = ($signed(_zz_3025) - $signed(_zz_11291));
  assign _zz_3024 = ($signed(_zz_3025) + $signed(_zz_11293));
  assign _zz_3026 = 1'b1;
  assign _zz_3027 = 1'b1;
  assign _zz_4780 = ($signed(_zz_11311) * $signed(_zz_991));
  assign _zz_3030 = _zz_11312[15 : 0];
  assign _zz_4781 = ($signed(_zz_11313) * $signed(twiddle_factor_table_14_real));
  assign _zz_4782 = ($signed(_zz_11314) * $signed(twiddle_factor_table_14_imag));
  assign _zz_3028 = ($signed(_zz_3030) - $signed(_zz_11315));
  assign _zz_3029 = ($signed(_zz_3030) + $signed(_zz_11317));
  assign _zz_3031 = 1'b1;
  assign _zz_3032 = 1'b1;
  assign _zz_4783 = ($signed(_zz_11335) * $signed(_zz_1009));
  assign _zz_3035 = _zz_11336[15 : 0];
  assign _zz_4784 = ($signed(_zz_11337) * $signed(twiddle_factor_table_7_real));
  assign _zz_4785 = ($signed(_zz_11338) * $signed(twiddle_factor_table_7_imag));
  assign _zz_3033 = ($signed(_zz_3035) - $signed(_zz_11339));
  assign _zz_3034 = ($signed(_zz_3035) + $signed(_zz_11341));
  assign _zz_3036 = 1'b1;
  assign _zz_3037 = 1'b1;
  assign _zz_4786 = ($signed(_zz_11359) * $signed(_zz_1011));
  assign _zz_3040 = _zz_11360[15 : 0];
  assign _zz_4787 = ($signed(_zz_11361) * $signed(twiddle_factor_table_8_real));
  assign _zz_4788 = ($signed(_zz_11362) * $signed(twiddle_factor_table_8_imag));
  assign _zz_3038 = ($signed(_zz_3040) - $signed(_zz_11363));
  assign _zz_3039 = ($signed(_zz_3040) + $signed(_zz_11365));
  assign _zz_3041 = 1'b1;
  assign _zz_3042 = 1'b1;
  assign _zz_4789 = ($signed(_zz_11383) * $signed(_zz_1013));
  assign _zz_3045 = _zz_11384[15 : 0];
  assign _zz_4790 = ($signed(_zz_11385) * $signed(twiddle_factor_table_9_real));
  assign _zz_4791 = ($signed(_zz_11386) * $signed(twiddle_factor_table_9_imag));
  assign _zz_3043 = ($signed(_zz_3045) - $signed(_zz_11387));
  assign _zz_3044 = ($signed(_zz_3045) + $signed(_zz_11389));
  assign _zz_3046 = 1'b1;
  assign _zz_3047 = 1'b1;
  assign _zz_4792 = ($signed(_zz_11407) * $signed(_zz_1015));
  assign _zz_3050 = _zz_11408[15 : 0];
  assign _zz_4793 = ($signed(_zz_11409) * $signed(twiddle_factor_table_10_real));
  assign _zz_4794 = ($signed(_zz_11410) * $signed(twiddle_factor_table_10_imag));
  assign _zz_3048 = ($signed(_zz_3050) - $signed(_zz_11411));
  assign _zz_3049 = ($signed(_zz_3050) + $signed(_zz_11413));
  assign _zz_3051 = 1'b1;
  assign _zz_3052 = 1'b1;
  assign _zz_4795 = ($signed(_zz_11431) * $signed(_zz_1017));
  assign _zz_3055 = _zz_11432[15 : 0];
  assign _zz_4796 = ($signed(_zz_11433) * $signed(twiddle_factor_table_11_real));
  assign _zz_4797 = ($signed(_zz_11434) * $signed(twiddle_factor_table_11_imag));
  assign _zz_3053 = ($signed(_zz_3055) - $signed(_zz_11435));
  assign _zz_3054 = ($signed(_zz_3055) + $signed(_zz_11437));
  assign _zz_3056 = 1'b1;
  assign _zz_3057 = 1'b1;
  assign _zz_4798 = ($signed(_zz_11455) * $signed(_zz_1019));
  assign _zz_3060 = _zz_11456[15 : 0];
  assign _zz_4799 = ($signed(_zz_11457) * $signed(twiddle_factor_table_12_real));
  assign _zz_4800 = ($signed(_zz_11458) * $signed(twiddle_factor_table_12_imag));
  assign _zz_3058 = ($signed(_zz_3060) - $signed(_zz_11459));
  assign _zz_3059 = ($signed(_zz_3060) + $signed(_zz_11461));
  assign _zz_3061 = 1'b1;
  assign _zz_3062 = 1'b1;
  assign _zz_4801 = ($signed(_zz_11479) * $signed(_zz_1021));
  assign _zz_3065 = _zz_11480[15 : 0];
  assign _zz_4802 = ($signed(_zz_11481) * $signed(twiddle_factor_table_13_real));
  assign _zz_4803 = ($signed(_zz_11482) * $signed(twiddle_factor_table_13_imag));
  assign _zz_3063 = ($signed(_zz_3065) - $signed(_zz_11483));
  assign _zz_3064 = ($signed(_zz_3065) + $signed(_zz_11485));
  assign _zz_3066 = 1'b1;
  assign _zz_3067 = 1'b1;
  assign _zz_4804 = ($signed(_zz_11503) * $signed(_zz_1023));
  assign _zz_3070 = _zz_11504[15 : 0];
  assign _zz_4805 = ($signed(_zz_11505) * $signed(twiddle_factor_table_14_real));
  assign _zz_4806 = ($signed(_zz_11506) * $signed(twiddle_factor_table_14_imag));
  assign _zz_3068 = ($signed(_zz_3070) - $signed(_zz_11507));
  assign _zz_3069 = ($signed(_zz_3070) + $signed(_zz_11509));
  assign _zz_3071 = 1'b1;
  assign _zz_3072 = 1'b1;
  assign _zz_4807 = ($signed(_zz_11527) * $signed(_zz_1057));
  assign _zz_3075 = _zz_11528[15 : 0];
  assign _zz_4808 = ($signed(_zz_11529) * $signed(twiddle_factor_table_15_real));
  assign _zz_4809 = ($signed(_zz_11530) * $signed(twiddle_factor_table_15_imag));
  assign _zz_3073 = ($signed(_zz_3075) - $signed(_zz_11531));
  assign _zz_3074 = ($signed(_zz_3075) + $signed(_zz_11533));
  assign _zz_3076 = 1'b1;
  assign _zz_3077 = 1'b1;
  assign _zz_4810 = ($signed(_zz_11551) * $signed(_zz_1059));
  assign _zz_3080 = _zz_11552[15 : 0];
  assign _zz_4811 = ($signed(_zz_11553) * $signed(twiddle_factor_table_16_real));
  assign _zz_4812 = ($signed(_zz_11554) * $signed(twiddle_factor_table_16_imag));
  assign _zz_3078 = ($signed(_zz_3080) - $signed(_zz_11555));
  assign _zz_3079 = ($signed(_zz_3080) + $signed(_zz_11557));
  assign _zz_3081 = 1'b1;
  assign _zz_3082 = 1'b1;
  assign _zz_4813 = ($signed(_zz_11575) * $signed(_zz_1061));
  assign _zz_3085 = _zz_11576[15 : 0];
  assign _zz_4814 = ($signed(_zz_11577) * $signed(twiddle_factor_table_17_real));
  assign _zz_4815 = ($signed(_zz_11578) * $signed(twiddle_factor_table_17_imag));
  assign _zz_3083 = ($signed(_zz_3085) - $signed(_zz_11579));
  assign _zz_3084 = ($signed(_zz_3085) + $signed(_zz_11581));
  assign _zz_3086 = 1'b1;
  assign _zz_3087 = 1'b1;
  assign _zz_4816 = ($signed(_zz_11599) * $signed(_zz_1063));
  assign _zz_3090 = _zz_11600[15 : 0];
  assign _zz_4817 = ($signed(_zz_11601) * $signed(twiddle_factor_table_18_real));
  assign _zz_4818 = ($signed(_zz_11602) * $signed(twiddle_factor_table_18_imag));
  assign _zz_3088 = ($signed(_zz_3090) - $signed(_zz_11603));
  assign _zz_3089 = ($signed(_zz_3090) + $signed(_zz_11605));
  assign _zz_3091 = 1'b1;
  assign _zz_3092 = 1'b1;
  assign _zz_4819 = ($signed(_zz_11623) * $signed(_zz_1065));
  assign _zz_3095 = _zz_11624[15 : 0];
  assign _zz_4820 = ($signed(_zz_11625) * $signed(twiddle_factor_table_19_real));
  assign _zz_4821 = ($signed(_zz_11626) * $signed(twiddle_factor_table_19_imag));
  assign _zz_3093 = ($signed(_zz_3095) - $signed(_zz_11627));
  assign _zz_3094 = ($signed(_zz_3095) + $signed(_zz_11629));
  assign _zz_3096 = 1'b1;
  assign _zz_3097 = 1'b1;
  assign _zz_4822 = ($signed(_zz_11647) * $signed(_zz_1067));
  assign _zz_3100 = _zz_11648[15 : 0];
  assign _zz_4823 = ($signed(_zz_11649) * $signed(twiddle_factor_table_20_real));
  assign _zz_4824 = ($signed(_zz_11650) * $signed(twiddle_factor_table_20_imag));
  assign _zz_3098 = ($signed(_zz_3100) - $signed(_zz_11651));
  assign _zz_3099 = ($signed(_zz_3100) + $signed(_zz_11653));
  assign _zz_3101 = 1'b1;
  assign _zz_3102 = 1'b1;
  assign _zz_4825 = ($signed(_zz_11671) * $signed(_zz_1069));
  assign _zz_3105 = _zz_11672[15 : 0];
  assign _zz_4826 = ($signed(_zz_11673) * $signed(twiddle_factor_table_21_real));
  assign _zz_4827 = ($signed(_zz_11674) * $signed(twiddle_factor_table_21_imag));
  assign _zz_3103 = ($signed(_zz_3105) - $signed(_zz_11675));
  assign _zz_3104 = ($signed(_zz_3105) + $signed(_zz_11677));
  assign _zz_3106 = 1'b1;
  assign _zz_3107 = 1'b1;
  assign _zz_4828 = ($signed(_zz_11695) * $signed(_zz_1071));
  assign _zz_3110 = _zz_11696[15 : 0];
  assign _zz_4829 = ($signed(_zz_11697) * $signed(twiddle_factor_table_22_real));
  assign _zz_4830 = ($signed(_zz_11698) * $signed(twiddle_factor_table_22_imag));
  assign _zz_3108 = ($signed(_zz_3110) - $signed(_zz_11699));
  assign _zz_3109 = ($signed(_zz_3110) + $signed(_zz_11701));
  assign _zz_3111 = 1'b1;
  assign _zz_3112 = 1'b1;
  assign _zz_4831 = ($signed(_zz_11719) * $signed(_zz_1073));
  assign _zz_3115 = _zz_11720[15 : 0];
  assign _zz_4832 = ($signed(_zz_11721) * $signed(twiddle_factor_table_23_real));
  assign _zz_4833 = ($signed(_zz_11722) * $signed(twiddle_factor_table_23_imag));
  assign _zz_3113 = ($signed(_zz_3115) - $signed(_zz_11723));
  assign _zz_3114 = ($signed(_zz_3115) + $signed(_zz_11725));
  assign _zz_3116 = 1'b1;
  assign _zz_3117 = 1'b1;
  assign _zz_4834 = ($signed(_zz_11743) * $signed(_zz_1075));
  assign _zz_3120 = _zz_11744[15 : 0];
  assign _zz_4835 = ($signed(_zz_11745) * $signed(twiddle_factor_table_24_real));
  assign _zz_4836 = ($signed(_zz_11746) * $signed(twiddle_factor_table_24_imag));
  assign _zz_3118 = ($signed(_zz_3120) - $signed(_zz_11747));
  assign _zz_3119 = ($signed(_zz_3120) + $signed(_zz_11749));
  assign _zz_3121 = 1'b1;
  assign _zz_3122 = 1'b1;
  assign _zz_4837 = ($signed(_zz_11767) * $signed(_zz_1077));
  assign _zz_3125 = _zz_11768[15 : 0];
  assign _zz_4838 = ($signed(_zz_11769) * $signed(twiddle_factor_table_25_real));
  assign _zz_4839 = ($signed(_zz_11770) * $signed(twiddle_factor_table_25_imag));
  assign _zz_3123 = ($signed(_zz_3125) - $signed(_zz_11771));
  assign _zz_3124 = ($signed(_zz_3125) + $signed(_zz_11773));
  assign _zz_3126 = 1'b1;
  assign _zz_3127 = 1'b1;
  assign _zz_4840 = ($signed(_zz_11791) * $signed(_zz_1079));
  assign _zz_3130 = _zz_11792[15 : 0];
  assign _zz_4841 = ($signed(_zz_11793) * $signed(twiddle_factor_table_26_real));
  assign _zz_4842 = ($signed(_zz_11794) * $signed(twiddle_factor_table_26_imag));
  assign _zz_3128 = ($signed(_zz_3130) - $signed(_zz_11795));
  assign _zz_3129 = ($signed(_zz_3130) + $signed(_zz_11797));
  assign _zz_3131 = 1'b1;
  assign _zz_3132 = 1'b1;
  assign _zz_4843 = ($signed(_zz_11815) * $signed(_zz_1081));
  assign _zz_3135 = _zz_11816[15 : 0];
  assign _zz_4844 = ($signed(_zz_11817) * $signed(twiddle_factor_table_27_real));
  assign _zz_4845 = ($signed(_zz_11818) * $signed(twiddle_factor_table_27_imag));
  assign _zz_3133 = ($signed(_zz_3135) - $signed(_zz_11819));
  assign _zz_3134 = ($signed(_zz_3135) + $signed(_zz_11821));
  assign _zz_3136 = 1'b1;
  assign _zz_3137 = 1'b1;
  assign _zz_4846 = ($signed(_zz_11839) * $signed(_zz_1083));
  assign _zz_3140 = _zz_11840[15 : 0];
  assign _zz_4847 = ($signed(_zz_11841) * $signed(twiddle_factor_table_28_real));
  assign _zz_4848 = ($signed(_zz_11842) * $signed(twiddle_factor_table_28_imag));
  assign _zz_3138 = ($signed(_zz_3140) - $signed(_zz_11843));
  assign _zz_3139 = ($signed(_zz_3140) + $signed(_zz_11845));
  assign _zz_3141 = 1'b1;
  assign _zz_3142 = 1'b1;
  assign _zz_4849 = ($signed(_zz_11863) * $signed(_zz_1085));
  assign _zz_3145 = _zz_11864[15 : 0];
  assign _zz_4850 = ($signed(_zz_11865) * $signed(twiddle_factor_table_29_real));
  assign _zz_4851 = ($signed(_zz_11866) * $signed(twiddle_factor_table_29_imag));
  assign _zz_3143 = ($signed(_zz_3145) - $signed(_zz_11867));
  assign _zz_3144 = ($signed(_zz_3145) + $signed(_zz_11869));
  assign _zz_3146 = 1'b1;
  assign _zz_3147 = 1'b1;
  assign _zz_4852 = ($signed(_zz_11887) * $signed(_zz_1087));
  assign _zz_3150 = _zz_11888[15 : 0];
  assign _zz_4853 = ($signed(_zz_11889) * $signed(twiddle_factor_table_30_real));
  assign _zz_4854 = ($signed(_zz_11890) * $signed(twiddle_factor_table_30_imag));
  assign _zz_3148 = ($signed(_zz_3150) - $signed(_zz_11891));
  assign _zz_3149 = ($signed(_zz_3150) + $signed(_zz_11893));
  assign _zz_3151 = 1'b1;
  assign _zz_3152 = 1'b1;
  assign _zz_4855 = ($signed(_zz_11911) * $signed(_zz_1121));
  assign _zz_3155 = _zz_11912[15 : 0];
  assign _zz_4856 = ($signed(_zz_11913) * $signed(twiddle_factor_table_15_real));
  assign _zz_4857 = ($signed(_zz_11914) * $signed(twiddle_factor_table_15_imag));
  assign _zz_3153 = ($signed(_zz_3155) - $signed(_zz_11915));
  assign _zz_3154 = ($signed(_zz_3155) + $signed(_zz_11917));
  assign _zz_3156 = 1'b1;
  assign _zz_3157 = 1'b1;
  assign _zz_4858 = ($signed(_zz_11935) * $signed(_zz_1123));
  assign _zz_3160 = _zz_11936[15 : 0];
  assign _zz_4859 = ($signed(_zz_11937) * $signed(twiddle_factor_table_16_real));
  assign _zz_4860 = ($signed(_zz_11938) * $signed(twiddle_factor_table_16_imag));
  assign _zz_3158 = ($signed(_zz_3160) - $signed(_zz_11939));
  assign _zz_3159 = ($signed(_zz_3160) + $signed(_zz_11941));
  assign _zz_3161 = 1'b1;
  assign _zz_3162 = 1'b1;
  assign _zz_4861 = ($signed(_zz_11959) * $signed(_zz_1125));
  assign _zz_3165 = _zz_11960[15 : 0];
  assign _zz_4862 = ($signed(_zz_11961) * $signed(twiddle_factor_table_17_real));
  assign _zz_4863 = ($signed(_zz_11962) * $signed(twiddle_factor_table_17_imag));
  assign _zz_3163 = ($signed(_zz_3165) - $signed(_zz_11963));
  assign _zz_3164 = ($signed(_zz_3165) + $signed(_zz_11965));
  assign _zz_3166 = 1'b1;
  assign _zz_3167 = 1'b1;
  assign _zz_4864 = ($signed(_zz_11983) * $signed(_zz_1127));
  assign _zz_3170 = _zz_11984[15 : 0];
  assign _zz_4865 = ($signed(_zz_11985) * $signed(twiddle_factor_table_18_real));
  assign _zz_4866 = ($signed(_zz_11986) * $signed(twiddle_factor_table_18_imag));
  assign _zz_3168 = ($signed(_zz_3170) - $signed(_zz_11987));
  assign _zz_3169 = ($signed(_zz_3170) + $signed(_zz_11989));
  assign _zz_3171 = 1'b1;
  assign _zz_3172 = 1'b1;
  assign _zz_4867 = ($signed(_zz_12007) * $signed(_zz_1129));
  assign _zz_3175 = _zz_12008[15 : 0];
  assign _zz_4868 = ($signed(_zz_12009) * $signed(twiddle_factor_table_19_real));
  assign _zz_4869 = ($signed(_zz_12010) * $signed(twiddle_factor_table_19_imag));
  assign _zz_3173 = ($signed(_zz_3175) - $signed(_zz_12011));
  assign _zz_3174 = ($signed(_zz_3175) + $signed(_zz_12013));
  assign _zz_3176 = 1'b1;
  assign _zz_3177 = 1'b1;
  assign _zz_4870 = ($signed(_zz_12031) * $signed(_zz_1131));
  assign _zz_3180 = _zz_12032[15 : 0];
  assign _zz_4871 = ($signed(_zz_12033) * $signed(twiddle_factor_table_20_real));
  assign _zz_4872 = ($signed(_zz_12034) * $signed(twiddle_factor_table_20_imag));
  assign _zz_3178 = ($signed(_zz_3180) - $signed(_zz_12035));
  assign _zz_3179 = ($signed(_zz_3180) + $signed(_zz_12037));
  assign _zz_3181 = 1'b1;
  assign _zz_3182 = 1'b1;
  assign _zz_4873 = ($signed(_zz_12055) * $signed(_zz_1133));
  assign _zz_3185 = _zz_12056[15 : 0];
  assign _zz_4874 = ($signed(_zz_12057) * $signed(twiddle_factor_table_21_real));
  assign _zz_4875 = ($signed(_zz_12058) * $signed(twiddle_factor_table_21_imag));
  assign _zz_3183 = ($signed(_zz_3185) - $signed(_zz_12059));
  assign _zz_3184 = ($signed(_zz_3185) + $signed(_zz_12061));
  assign _zz_3186 = 1'b1;
  assign _zz_3187 = 1'b1;
  assign _zz_4876 = ($signed(_zz_12079) * $signed(_zz_1135));
  assign _zz_3190 = _zz_12080[15 : 0];
  assign _zz_4877 = ($signed(_zz_12081) * $signed(twiddle_factor_table_22_real));
  assign _zz_4878 = ($signed(_zz_12082) * $signed(twiddle_factor_table_22_imag));
  assign _zz_3188 = ($signed(_zz_3190) - $signed(_zz_12083));
  assign _zz_3189 = ($signed(_zz_3190) + $signed(_zz_12085));
  assign _zz_3191 = 1'b1;
  assign _zz_3192 = 1'b1;
  assign _zz_4879 = ($signed(_zz_12103) * $signed(_zz_1137));
  assign _zz_3195 = _zz_12104[15 : 0];
  assign _zz_4880 = ($signed(_zz_12105) * $signed(twiddle_factor_table_23_real));
  assign _zz_4881 = ($signed(_zz_12106) * $signed(twiddle_factor_table_23_imag));
  assign _zz_3193 = ($signed(_zz_3195) - $signed(_zz_12107));
  assign _zz_3194 = ($signed(_zz_3195) + $signed(_zz_12109));
  assign _zz_3196 = 1'b1;
  assign _zz_3197 = 1'b1;
  assign _zz_4882 = ($signed(_zz_12127) * $signed(_zz_1139));
  assign _zz_3200 = _zz_12128[15 : 0];
  assign _zz_4883 = ($signed(_zz_12129) * $signed(twiddle_factor_table_24_real));
  assign _zz_4884 = ($signed(_zz_12130) * $signed(twiddle_factor_table_24_imag));
  assign _zz_3198 = ($signed(_zz_3200) - $signed(_zz_12131));
  assign _zz_3199 = ($signed(_zz_3200) + $signed(_zz_12133));
  assign _zz_3201 = 1'b1;
  assign _zz_3202 = 1'b1;
  assign _zz_4885 = ($signed(_zz_12151) * $signed(_zz_1141));
  assign _zz_3205 = _zz_12152[15 : 0];
  assign _zz_4886 = ($signed(_zz_12153) * $signed(twiddle_factor_table_25_real));
  assign _zz_4887 = ($signed(_zz_12154) * $signed(twiddle_factor_table_25_imag));
  assign _zz_3203 = ($signed(_zz_3205) - $signed(_zz_12155));
  assign _zz_3204 = ($signed(_zz_3205) + $signed(_zz_12157));
  assign _zz_3206 = 1'b1;
  assign _zz_3207 = 1'b1;
  assign _zz_4888 = ($signed(_zz_12175) * $signed(_zz_1143));
  assign _zz_3210 = _zz_12176[15 : 0];
  assign _zz_4889 = ($signed(_zz_12177) * $signed(twiddle_factor_table_26_real));
  assign _zz_4890 = ($signed(_zz_12178) * $signed(twiddle_factor_table_26_imag));
  assign _zz_3208 = ($signed(_zz_3210) - $signed(_zz_12179));
  assign _zz_3209 = ($signed(_zz_3210) + $signed(_zz_12181));
  assign _zz_3211 = 1'b1;
  assign _zz_3212 = 1'b1;
  assign _zz_4891 = ($signed(_zz_12199) * $signed(_zz_1145));
  assign _zz_3215 = _zz_12200[15 : 0];
  assign _zz_4892 = ($signed(_zz_12201) * $signed(twiddle_factor_table_27_real));
  assign _zz_4893 = ($signed(_zz_12202) * $signed(twiddle_factor_table_27_imag));
  assign _zz_3213 = ($signed(_zz_3215) - $signed(_zz_12203));
  assign _zz_3214 = ($signed(_zz_3215) + $signed(_zz_12205));
  assign _zz_3216 = 1'b1;
  assign _zz_3217 = 1'b1;
  assign _zz_4894 = ($signed(_zz_12223) * $signed(_zz_1147));
  assign _zz_3220 = _zz_12224[15 : 0];
  assign _zz_4895 = ($signed(_zz_12225) * $signed(twiddle_factor_table_28_real));
  assign _zz_4896 = ($signed(_zz_12226) * $signed(twiddle_factor_table_28_imag));
  assign _zz_3218 = ($signed(_zz_3220) - $signed(_zz_12227));
  assign _zz_3219 = ($signed(_zz_3220) + $signed(_zz_12229));
  assign _zz_3221 = 1'b1;
  assign _zz_3222 = 1'b1;
  assign _zz_4897 = ($signed(_zz_12247) * $signed(_zz_1149));
  assign _zz_3225 = _zz_12248[15 : 0];
  assign _zz_4898 = ($signed(_zz_12249) * $signed(twiddle_factor_table_29_real));
  assign _zz_4899 = ($signed(_zz_12250) * $signed(twiddle_factor_table_29_imag));
  assign _zz_3223 = ($signed(_zz_3225) - $signed(_zz_12251));
  assign _zz_3224 = ($signed(_zz_3225) + $signed(_zz_12253));
  assign _zz_3226 = 1'b1;
  assign _zz_3227 = 1'b1;
  assign _zz_4900 = ($signed(_zz_12271) * $signed(_zz_1151));
  assign _zz_3230 = _zz_12272[15 : 0];
  assign _zz_4901 = ($signed(_zz_12273) * $signed(twiddle_factor_table_30_real));
  assign _zz_4902 = ($signed(_zz_12274) * $signed(twiddle_factor_table_30_imag));
  assign _zz_3228 = ($signed(_zz_3230) - $signed(_zz_12275));
  assign _zz_3229 = ($signed(_zz_3230) + $signed(_zz_12277));
  assign _zz_3231 = 1'b1;
  assign _zz_3232 = 1'b1;
  assign _zz_4903 = ($signed(_zz_12295) * $signed(_zz_1185));
  assign _zz_3235 = _zz_12296[15 : 0];
  assign _zz_4904 = ($signed(_zz_12297) * $signed(twiddle_factor_table_15_real));
  assign _zz_4905 = ($signed(_zz_12298) * $signed(twiddle_factor_table_15_imag));
  assign _zz_3233 = ($signed(_zz_3235) - $signed(_zz_12299));
  assign _zz_3234 = ($signed(_zz_3235) + $signed(_zz_12301));
  assign _zz_3236 = 1'b1;
  assign _zz_3237 = 1'b1;
  assign _zz_4906 = ($signed(_zz_12319) * $signed(_zz_1187));
  assign _zz_3240 = _zz_12320[15 : 0];
  assign _zz_4907 = ($signed(_zz_12321) * $signed(twiddle_factor_table_16_real));
  assign _zz_4908 = ($signed(_zz_12322) * $signed(twiddle_factor_table_16_imag));
  assign _zz_3238 = ($signed(_zz_3240) - $signed(_zz_12323));
  assign _zz_3239 = ($signed(_zz_3240) + $signed(_zz_12325));
  assign _zz_3241 = 1'b1;
  assign _zz_3242 = 1'b1;
  assign _zz_4909 = ($signed(_zz_12343) * $signed(_zz_1189));
  assign _zz_3245 = _zz_12344[15 : 0];
  assign _zz_4910 = ($signed(_zz_12345) * $signed(twiddle_factor_table_17_real));
  assign _zz_4911 = ($signed(_zz_12346) * $signed(twiddle_factor_table_17_imag));
  assign _zz_3243 = ($signed(_zz_3245) - $signed(_zz_12347));
  assign _zz_3244 = ($signed(_zz_3245) + $signed(_zz_12349));
  assign _zz_3246 = 1'b1;
  assign _zz_3247 = 1'b1;
  assign _zz_4912 = ($signed(_zz_12367) * $signed(_zz_1191));
  assign _zz_3250 = _zz_12368[15 : 0];
  assign _zz_4913 = ($signed(_zz_12369) * $signed(twiddle_factor_table_18_real));
  assign _zz_4914 = ($signed(_zz_12370) * $signed(twiddle_factor_table_18_imag));
  assign _zz_3248 = ($signed(_zz_3250) - $signed(_zz_12371));
  assign _zz_3249 = ($signed(_zz_3250) + $signed(_zz_12373));
  assign _zz_3251 = 1'b1;
  assign _zz_3252 = 1'b1;
  assign _zz_4915 = ($signed(_zz_12391) * $signed(_zz_1193));
  assign _zz_3255 = _zz_12392[15 : 0];
  assign _zz_4916 = ($signed(_zz_12393) * $signed(twiddle_factor_table_19_real));
  assign _zz_4917 = ($signed(_zz_12394) * $signed(twiddle_factor_table_19_imag));
  assign _zz_3253 = ($signed(_zz_3255) - $signed(_zz_12395));
  assign _zz_3254 = ($signed(_zz_3255) + $signed(_zz_12397));
  assign _zz_3256 = 1'b1;
  assign _zz_3257 = 1'b1;
  assign _zz_4918 = ($signed(_zz_12415) * $signed(_zz_1195));
  assign _zz_3260 = _zz_12416[15 : 0];
  assign _zz_4919 = ($signed(_zz_12417) * $signed(twiddle_factor_table_20_real));
  assign _zz_4920 = ($signed(_zz_12418) * $signed(twiddle_factor_table_20_imag));
  assign _zz_3258 = ($signed(_zz_3260) - $signed(_zz_12419));
  assign _zz_3259 = ($signed(_zz_3260) + $signed(_zz_12421));
  assign _zz_3261 = 1'b1;
  assign _zz_3262 = 1'b1;
  assign _zz_4921 = ($signed(_zz_12439) * $signed(_zz_1197));
  assign _zz_3265 = _zz_12440[15 : 0];
  assign _zz_4922 = ($signed(_zz_12441) * $signed(twiddle_factor_table_21_real));
  assign _zz_4923 = ($signed(_zz_12442) * $signed(twiddle_factor_table_21_imag));
  assign _zz_3263 = ($signed(_zz_3265) - $signed(_zz_12443));
  assign _zz_3264 = ($signed(_zz_3265) + $signed(_zz_12445));
  assign _zz_3266 = 1'b1;
  assign _zz_3267 = 1'b1;
  assign _zz_4924 = ($signed(_zz_12463) * $signed(_zz_1199));
  assign _zz_3270 = _zz_12464[15 : 0];
  assign _zz_4925 = ($signed(_zz_12465) * $signed(twiddle_factor_table_22_real));
  assign _zz_4926 = ($signed(_zz_12466) * $signed(twiddle_factor_table_22_imag));
  assign _zz_3268 = ($signed(_zz_3270) - $signed(_zz_12467));
  assign _zz_3269 = ($signed(_zz_3270) + $signed(_zz_12469));
  assign _zz_3271 = 1'b1;
  assign _zz_3272 = 1'b1;
  assign _zz_4927 = ($signed(_zz_12487) * $signed(_zz_1201));
  assign _zz_3275 = _zz_12488[15 : 0];
  assign _zz_4928 = ($signed(_zz_12489) * $signed(twiddle_factor_table_23_real));
  assign _zz_4929 = ($signed(_zz_12490) * $signed(twiddle_factor_table_23_imag));
  assign _zz_3273 = ($signed(_zz_3275) - $signed(_zz_12491));
  assign _zz_3274 = ($signed(_zz_3275) + $signed(_zz_12493));
  assign _zz_3276 = 1'b1;
  assign _zz_3277 = 1'b1;
  assign _zz_4930 = ($signed(_zz_12511) * $signed(_zz_1203));
  assign _zz_3280 = _zz_12512[15 : 0];
  assign _zz_4931 = ($signed(_zz_12513) * $signed(twiddle_factor_table_24_real));
  assign _zz_4932 = ($signed(_zz_12514) * $signed(twiddle_factor_table_24_imag));
  assign _zz_3278 = ($signed(_zz_3280) - $signed(_zz_12515));
  assign _zz_3279 = ($signed(_zz_3280) + $signed(_zz_12517));
  assign _zz_3281 = 1'b1;
  assign _zz_3282 = 1'b1;
  assign _zz_4933 = ($signed(_zz_12535) * $signed(_zz_1205));
  assign _zz_3285 = _zz_12536[15 : 0];
  assign _zz_4934 = ($signed(_zz_12537) * $signed(twiddle_factor_table_25_real));
  assign _zz_4935 = ($signed(_zz_12538) * $signed(twiddle_factor_table_25_imag));
  assign _zz_3283 = ($signed(_zz_3285) - $signed(_zz_12539));
  assign _zz_3284 = ($signed(_zz_3285) + $signed(_zz_12541));
  assign _zz_3286 = 1'b1;
  assign _zz_3287 = 1'b1;
  assign _zz_4936 = ($signed(_zz_12559) * $signed(_zz_1207));
  assign _zz_3290 = _zz_12560[15 : 0];
  assign _zz_4937 = ($signed(_zz_12561) * $signed(twiddle_factor_table_26_real));
  assign _zz_4938 = ($signed(_zz_12562) * $signed(twiddle_factor_table_26_imag));
  assign _zz_3288 = ($signed(_zz_3290) - $signed(_zz_12563));
  assign _zz_3289 = ($signed(_zz_3290) + $signed(_zz_12565));
  assign _zz_3291 = 1'b1;
  assign _zz_3292 = 1'b1;
  assign _zz_4939 = ($signed(_zz_12583) * $signed(_zz_1209));
  assign _zz_3295 = _zz_12584[15 : 0];
  assign _zz_4940 = ($signed(_zz_12585) * $signed(twiddle_factor_table_27_real));
  assign _zz_4941 = ($signed(_zz_12586) * $signed(twiddle_factor_table_27_imag));
  assign _zz_3293 = ($signed(_zz_3295) - $signed(_zz_12587));
  assign _zz_3294 = ($signed(_zz_3295) + $signed(_zz_12589));
  assign _zz_3296 = 1'b1;
  assign _zz_3297 = 1'b1;
  assign _zz_4942 = ($signed(_zz_12607) * $signed(_zz_1211));
  assign _zz_3300 = _zz_12608[15 : 0];
  assign _zz_4943 = ($signed(_zz_12609) * $signed(twiddle_factor_table_28_real));
  assign _zz_4944 = ($signed(_zz_12610) * $signed(twiddle_factor_table_28_imag));
  assign _zz_3298 = ($signed(_zz_3300) - $signed(_zz_12611));
  assign _zz_3299 = ($signed(_zz_3300) + $signed(_zz_12613));
  assign _zz_3301 = 1'b1;
  assign _zz_3302 = 1'b1;
  assign _zz_4945 = ($signed(_zz_12631) * $signed(_zz_1213));
  assign _zz_3305 = _zz_12632[15 : 0];
  assign _zz_4946 = ($signed(_zz_12633) * $signed(twiddle_factor_table_29_real));
  assign _zz_4947 = ($signed(_zz_12634) * $signed(twiddle_factor_table_29_imag));
  assign _zz_3303 = ($signed(_zz_3305) - $signed(_zz_12635));
  assign _zz_3304 = ($signed(_zz_3305) + $signed(_zz_12637));
  assign _zz_3306 = 1'b1;
  assign _zz_3307 = 1'b1;
  assign _zz_4948 = ($signed(_zz_12655) * $signed(_zz_1215));
  assign _zz_3310 = _zz_12656[15 : 0];
  assign _zz_4949 = ($signed(_zz_12657) * $signed(twiddle_factor_table_30_real));
  assign _zz_4950 = ($signed(_zz_12658) * $signed(twiddle_factor_table_30_imag));
  assign _zz_3308 = ($signed(_zz_3310) - $signed(_zz_12659));
  assign _zz_3309 = ($signed(_zz_3310) + $signed(_zz_12661));
  assign _zz_3311 = 1'b1;
  assign _zz_3312 = 1'b1;
  assign _zz_4951 = ($signed(_zz_12679) * $signed(_zz_1249));
  assign _zz_3315 = _zz_12680[15 : 0];
  assign _zz_4952 = ($signed(_zz_12681) * $signed(twiddle_factor_table_15_real));
  assign _zz_4953 = ($signed(_zz_12682) * $signed(twiddle_factor_table_15_imag));
  assign _zz_3313 = ($signed(_zz_3315) - $signed(_zz_12683));
  assign _zz_3314 = ($signed(_zz_3315) + $signed(_zz_12685));
  assign _zz_3316 = 1'b1;
  assign _zz_3317 = 1'b1;
  assign _zz_4954 = ($signed(_zz_12703) * $signed(_zz_1251));
  assign _zz_3320 = _zz_12704[15 : 0];
  assign _zz_4955 = ($signed(_zz_12705) * $signed(twiddle_factor_table_16_real));
  assign _zz_4956 = ($signed(_zz_12706) * $signed(twiddle_factor_table_16_imag));
  assign _zz_3318 = ($signed(_zz_3320) - $signed(_zz_12707));
  assign _zz_3319 = ($signed(_zz_3320) + $signed(_zz_12709));
  assign _zz_3321 = 1'b1;
  assign _zz_3322 = 1'b1;
  assign _zz_4957 = ($signed(_zz_12727) * $signed(_zz_1253));
  assign _zz_3325 = _zz_12728[15 : 0];
  assign _zz_4958 = ($signed(_zz_12729) * $signed(twiddle_factor_table_17_real));
  assign _zz_4959 = ($signed(_zz_12730) * $signed(twiddle_factor_table_17_imag));
  assign _zz_3323 = ($signed(_zz_3325) - $signed(_zz_12731));
  assign _zz_3324 = ($signed(_zz_3325) + $signed(_zz_12733));
  assign _zz_3326 = 1'b1;
  assign _zz_3327 = 1'b1;
  assign _zz_4960 = ($signed(_zz_12751) * $signed(_zz_1255));
  assign _zz_3330 = _zz_12752[15 : 0];
  assign _zz_4961 = ($signed(_zz_12753) * $signed(twiddle_factor_table_18_real));
  assign _zz_4962 = ($signed(_zz_12754) * $signed(twiddle_factor_table_18_imag));
  assign _zz_3328 = ($signed(_zz_3330) - $signed(_zz_12755));
  assign _zz_3329 = ($signed(_zz_3330) + $signed(_zz_12757));
  assign _zz_3331 = 1'b1;
  assign _zz_3332 = 1'b1;
  assign _zz_4963 = ($signed(_zz_12775) * $signed(_zz_1257));
  assign _zz_3335 = _zz_12776[15 : 0];
  assign _zz_4964 = ($signed(_zz_12777) * $signed(twiddle_factor_table_19_real));
  assign _zz_4965 = ($signed(_zz_12778) * $signed(twiddle_factor_table_19_imag));
  assign _zz_3333 = ($signed(_zz_3335) - $signed(_zz_12779));
  assign _zz_3334 = ($signed(_zz_3335) + $signed(_zz_12781));
  assign _zz_3336 = 1'b1;
  assign _zz_3337 = 1'b1;
  assign _zz_4966 = ($signed(_zz_12799) * $signed(_zz_1259));
  assign _zz_3340 = _zz_12800[15 : 0];
  assign _zz_4967 = ($signed(_zz_12801) * $signed(twiddle_factor_table_20_real));
  assign _zz_4968 = ($signed(_zz_12802) * $signed(twiddle_factor_table_20_imag));
  assign _zz_3338 = ($signed(_zz_3340) - $signed(_zz_12803));
  assign _zz_3339 = ($signed(_zz_3340) + $signed(_zz_12805));
  assign _zz_3341 = 1'b1;
  assign _zz_3342 = 1'b1;
  assign _zz_4969 = ($signed(_zz_12823) * $signed(_zz_1261));
  assign _zz_3345 = _zz_12824[15 : 0];
  assign _zz_4970 = ($signed(_zz_12825) * $signed(twiddle_factor_table_21_real));
  assign _zz_4971 = ($signed(_zz_12826) * $signed(twiddle_factor_table_21_imag));
  assign _zz_3343 = ($signed(_zz_3345) - $signed(_zz_12827));
  assign _zz_3344 = ($signed(_zz_3345) + $signed(_zz_12829));
  assign _zz_3346 = 1'b1;
  assign _zz_3347 = 1'b1;
  assign _zz_4972 = ($signed(_zz_12847) * $signed(_zz_1263));
  assign _zz_3350 = _zz_12848[15 : 0];
  assign _zz_4973 = ($signed(_zz_12849) * $signed(twiddle_factor_table_22_real));
  assign _zz_4974 = ($signed(_zz_12850) * $signed(twiddle_factor_table_22_imag));
  assign _zz_3348 = ($signed(_zz_3350) - $signed(_zz_12851));
  assign _zz_3349 = ($signed(_zz_3350) + $signed(_zz_12853));
  assign _zz_3351 = 1'b1;
  assign _zz_3352 = 1'b1;
  assign _zz_4975 = ($signed(_zz_12871) * $signed(_zz_1265));
  assign _zz_3355 = _zz_12872[15 : 0];
  assign _zz_4976 = ($signed(_zz_12873) * $signed(twiddle_factor_table_23_real));
  assign _zz_4977 = ($signed(_zz_12874) * $signed(twiddle_factor_table_23_imag));
  assign _zz_3353 = ($signed(_zz_3355) - $signed(_zz_12875));
  assign _zz_3354 = ($signed(_zz_3355) + $signed(_zz_12877));
  assign _zz_3356 = 1'b1;
  assign _zz_3357 = 1'b1;
  assign _zz_4978 = ($signed(_zz_12895) * $signed(_zz_1267));
  assign _zz_3360 = _zz_12896[15 : 0];
  assign _zz_4979 = ($signed(_zz_12897) * $signed(twiddle_factor_table_24_real));
  assign _zz_4980 = ($signed(_zz_12898) * $signed(twiddle_factor_table_24_imag));
  assign _zz_3358 = ($signed(_zz_3360) - $signed(_zz_12899));
  assign _zz_3359 = ($signed(_zz_3360) + $signed(_zz_12901));
  assign _zz_3361 = 1'b1;
  assign _zz_3362 = 1'b1;
  assign _zz_4981 = ($signed(_zz_12919) * $signed(_zz_1269));
  assign _zz_3365 = _zz_12920[15 : 0];
  assign _zz_4982 = ($signed(_zz_12921) * $signed(twiddle_factor_table_25_real));
  assign _zz_4983 = ($signed(_zz_12922) * $signed(twiddle_factor_table_25_imag));
  assign _zz_3363 = ($signed(_zz_3365) - $signed(_zz_12923));
  assign _zz_3364 = ($signed(_zz_3365) + $signed(_zz_12925));
  assign _zz_3366 = 1'b1;
  assign _zz_3367 = 1'b1;
  assign _zz_4984 = ($signed(_zz_12943) * $signed(_zz_1271));
  assign _zz_3370 = _zz_12944[15 : 0];
  assign _zz_4985 = ($signed(_zz_12945) * $signed(twiddle_factor_table_26_real));
  assign _zz_4986 = ($signed(_zz_12946) * $signed(twiddle_factor_table_26_imag));
  assign _zz_3368 = ($signed(_zz_3370) - $signed(_zz_12947));
  assign _zz_3369 = ($signed(_zz_3370) + $signed(_zz_12949));
  assign _zz_3371 = 1'b1;
  assign _zz_3372 = 1'b1;
  assign _zz_4987 = ($signed(_zz_12967) * $signed(_zz_1273));
  assign _zz_3375 = _zz_12968[15 : 0];
  assign _zz_4988 = ($signed(_zz_12969) * $signed(twiddle_factor_table_27_real));
  assign _zz_4989 = ($signed(_zz_12970) * $signed(twiddle_factor_table_27_imag));
  assign _zz_3373 = ($signed(_zz_3375) - $signed(_zz_12971));
  assign _zz_3374 = ($signed(_zz_3375) + $signed(_zz_12973));
  assign _zz_3376 = 1'b1;
  assign _zz_3377 = 1'b1;
  assign _zz_4990 = ($signed(_zz_12991) * $signed(_zz_1275));
  assign _zz_3380 = _zz_12992[15 : 0];
  assign _zz_4991 = ($signed(_zz_12993) * $signed(twiddle_factor_table_28_real));
  assign _zz_4992 = ($signed(_zz_12994) * $signed(twiddle_factor_table_28_imag));
  assign _zz_3378 = ($signed(_zz_3380) - $signed(_zz_12995));
  assign _zz_3379 = ($signed(_zz_3380) + $signed(_zz_12997));
  assign _zz_3381 = 1'b1;
  assign _zz_3382 = 1'b1;
  assign _zz_4993 = ($signed(_zz_13015) * $signed(_zz_1277));
  assign _zz_3385 = _zz_13016[15 : 0];
  assign _zz_4994 = ($signed(_zz_13017) * $signed(twiddle_factor_table_29_real));
  assign _zz_4995 = ($signed(_zz_13018) * $signed(twiddle_factor_table_29_imag));
  assign _zz_3383 = ($signed(_zz_3385) - $signed(_zz_13019));
  assign _zz_3384 = ($signed(_zz_3385) + $signed(_zz_13021));
  assign _zz_3386 = 1'b1;
  assign _zz_3387 = 1'b1;
  assign _zz_4996 = ($signed(_zz_13039) * $signed(_zz_1279));
  assign _zz_3390 = _zz_13040[15 : 0];
  assign _zz_4997 = ($signed(_zz_13041) * $signed(twiddle_factor_table_30_real));
  assign _zz_4998 = ($signed(_zz_13042) * $signed(twiddle_factor_table_30_imag));
  assign _zz_3388 = ($signed(_zz_3390) - $signed(_zz_13043));
  assign _zz_3389 = ($signed(_zz_3390) + $signed(_zz_13045));
  assign _zz_3391 = 1'b1;
  assign _zz_3392 = 1'b1;
  assign _zz_4999 = ($signed(_zz_13063) * $signed(_zz_1345));
  assign _zz_3395 = _zz_13064[15 : 0];
  assign _zz_5000 = ($signed(_zz_13065) * $signed(twiddle_factor_table_31_real));
  assign _zz_5001 = ($signed(_zz_13066) * $signed(twiddle_factor_table_31_imag));
  assign _zz_3393 = ($signed(_zz_3395) - $signed(_zz_13067));
  assign _zz_3394 = ($signed(_zz_3395) + $signed(_zz_13069));
  assign _zz_3396 = 1'b1;
  assign _zz_3397 = 1'b1;
  assign _zz_5002 = ($signed(_zz_13087) * $signed(_zz_1347));
  assign _zz_3400 = _zz_13088[15 : 0];
  assign _zz_5003 = ($signed(_zz_13089) * $signed(twiddle_factor_table_32_real));
  assign _zz_5004 = ($signed(_zz_13090) * $signed(twiddle_factor_table_32_imag));
  assign _zz_3398 = ($signed(_zz_3400) - $signed(_zz_13091));
  assign _zz_3399 = ($signed(_zz_3400) + $signed(_zz_13093));
  assign _zz_3401 = 1'b1;
  assign _zz_3402 = 1'b1;
  assign _zz_5005 = ($signed(_zz_13111) * $signed(_zz_1349));
  assign _zz_3405 = _zz_13112[15 : 0];
  assign _zz_5006 = ($signed(_zz_13113) * $signed(twiddle_factor_table_33_real));
  assign _zz_5007 = ($signed(_zz_13114) * $signed(twiddle_factor_table_33_imag));
  assign _zz_3403 = ($signed(_zz_3405) - $signed(_zz_13115));
  assign _zz_3404 = ($signed(_zz_3405) + $signed(_zz_13117));
  assign _zz_3406 = 1'b1;
  assign _zz_3407 = 1'b1;
  assign _zz_5008 = ($signed(_zz_13135) * $signed(_zz_1351));
  assign _zz_3410 = _zz_13136[15 : 0];
  assign _zz_5009 = ($signed(_zz_13137) * $signed(twiddle_factor_table_34_real));
  assign _zz_5010 = ($signed(_zz_13138) * $signed(twiddle_factor_table_34_imag));
  assign _zz_3408 = ($signed(_zz_3410) - $signed(_zz_13139));
  assign _zz_3409 = ($signed(_zz_3410) + $signed(_zz_13141));
  assign _zz_3411 = 1'b1;
  assign _zz_3412 = 1'b1;
  assign _zz_5011 = ($signed(_zz_13159) * $signed(_zz_1353));
  assign _zz_3415 = _zz_13160[15 : 0];
  assign _zz_5012 = ($signed(_zz_13161) * $signed(twiddle_factor_table_35_real));
  assign _zz_5013 = ($signed(_zz_13162) * $signed(twiddle_factor_table_35_imag));
  assign _zz_3413 = ($signed(_zz_3415) - $signed(_zz_13163));
  assign _zz_3414 = ($signed(_zz_3415) + $signed(_zz_13165));
  assign _zz_3416 = 1'b1;
  assign _zz_3417 = 1'b1;
  assign _zz_5014 = ($signed(_zz_13183) * $signed(_zz_1355));
  assign _zz_3420 = _zz_13184[15 : 0];
  assign _zz_5015 = ($signed(_zz_13185) * $signed(twiddle_factor_table_36_real));
  assign _zz_5016 = ($signed(_zz_13186) * $signed(twiddle_factor_table_36_imag));
  assign _zz_3418 = ($signed(_zz_3420) - $signed(_zz_13187));
  assign _zz_3419 = ($signed(_zz_3420) + $signed(_zz_13189));
  assign _zz_3421 = 1'b1;
  assign _zz_3422 = 1'b1;
  assign _zz_5017 = ($signed(_zz_13207) * $signed(_zz_1357));
  assign _zz_3425 = _zz_13208[15 : 0];
  assign _zz_5018 = ($signed(_zz_13209) * $signed(twiddle_factor_table_37_real));
  assign _zz_5019 = ($signed(_zz_13210) * $signed(twiddle_factor_table_37_imag));
  assign _zz_3423 = ($signed(_zz_3425) - $signed(_zz_13211));
  assign _zz_3424 = ($signed(_zz_3425) + $signed(_zz_13213));
  assign _zz_3426 = 1'b1;
  assign _zz_3427 = 1'b1;
  assign _zz_5020 = ($signed(_zz_13231) * $signed(_zz_1359));
  assign _zz_3430 = _zz_13232[15 : 0];
  assign _zz_5021 = ($signed(_zz_13233) * $signed(twiddle_factor_table_38_real));
  assign _zz_5022 = ($signed(_zz_13234) * $signed(twiddle_factor_table_38_imag));
  assign _zz_3428 = ($signed(_zz_3430) - $signed(_zz_13235));
  assign _zz_3429 = ($signed(_zz_3430) + $signed(_zz_13237));
  assign _zz_3431 = 1'b1;
  assign _zz_3432 = 1'b1;
  assign _zz_5023 = ($signed(_zz_13255) * $signed(_zz_1361));
  assign _zz_3435 = _zz_13256[15 : 0];
  assign _zz_5024 = ($signed(_zz_13257) * $signed(twiddle_factor_table_39_real));
  assign _zz_5025 = ($signed(_zz_13258) * $signed(twiddle_factor_table_39_imag));
  assign _zz_3433 = ($signed(_zz_3435) - $signed(_zz_13259));
  assign _zz_3434 = ($signed(_zz_3435) + $signed(_zz_13261));
  assign _zz_3436 = 1'b1;
  assign _zz_3437 = 1'b1;
  assign _zz_5026 = ($signed(_zz_13279) * $signed(_zz_1363));
  assign _zz_3440 = _zz_13280[15 : 0];
  assign _zz_5027 = ($signed(_zz_13281) * $signed(twiddle_factor_table_40_real));
  assign _zz_5028 = ($signed(_zz_13282) * $signed(twiddle_factor_table_40_imag));
  assign _zz_3438 = ($signed(_zz_3440) - $signed(_zz_13283));
  assign _zz_3439 = ($signed(_zz_3440) + $signed(_zz_13285));
  assign _zz_3441 = 1'b1;
  assign _zz_3442 = 1'b1;
  assign _zz_5029 = ($signed(_zz_13303) * $signed(_zz_1365));
  assign _zz_3445 = _zz_13304[15 : 0];
  assign _zz_5030 = ($signed(_zz_13305) * $signed(twiddle_factor_table_41_real));
  assign _zz_5031 = ($signed(_zz_13306) * $signed(twiddle_factor_table_41_imag));
  assign _zz_3443 = ($signed(_zz_3445) - $signed(_zz_13307));
  assign _zz_3444 = ($signed(_zz_3445) + $signed(_zz_13309));
  assign _zz_3446 = 1'b1;
  assign _zz_3447 = 1'b1;
  assign _zz_5032 = ($signed(_zz_13327) * $signed(_zz_1367));
  assign _zz_3450 = _zz_13328[15 : 0];
  assign _zz_5033 = ($signed(_zz_13329) * $signed(twiddle_factor_table_42_real));
  assign _zz_5034 = ($signed(_zz_13330) * $signed(twiddle_factor_table_42_imag));
  assign _zz_3448 = ($signed(_zz_3450) - $signed(_zz_13331));
  assign _zz_3449 = ($signed(_zz_3450) + $signed(_zz_13333));
  assign _zz_3451 = 1'b1;
  assign _zz_3452 = 1'b1;
  assign _zz_5035 = ($signed(_zz_13351) * $signed(_zz_1369));
  assign _zz_3455 = _zz_13352[15 : 0];
  assign _zz_5036 = ($signed(_zz_13353) * $signed(twiddle_factor_table_43_real));
  assign _zz_5037 = ($signed(_zz_13354) * $signed(twiddle_factor_table_43_imag));
  assign _zz_3453 = ($signed(_zz_3455) - $signed(_zz_13355));
  assign _zz_3454 = ($signed(_zz_3455) + $signed(_zz_13357));
  assign _zz_3456 = 1'b1;
  assign _zz_3457 = 1'b1;
  assign _zz_5038 = ($signed(_zz_13375) * $signed(_zz_1371));
  assign _zz_3460 = _zz_13376[15 : 0];
  assign _zz_5039 = ($signed(_zz_13377) * $signed(twiddle_factor_table_44_real));
  assign _zz_5040 = ($signed(_zz_13378) * $signed(twiddle_factor_table_44_imag));
  assign _zz_3458 = ($signed(_zz_3460) - $signed(_zz_13379));
  assign _zz_3459 = ($signed(_zz_3460) + $signed(_zz_13381));
  assign _zz_3461 = 1'b1;
  assign _zz_3462 = 1'b1;
  assign _zz_5041 = ($signed(_zz_13399) * $signed(_zz_1373));
  assign _zz_3465 = _zz_13400[15 : 0];
  assign _zz_5042 = ($signed(_zz_13401) * $signed(twiddle_factor_table_45_real));
  assign _zz_5043 = ($signed(_zz_13402) * $signed(twiddle_factor_table_45_imag));
  assign _zz_3463 = ($signed(_zz_3465) - $signed(_zz_13403));
  assign _zz_3464 = ($signed(_zz_3465) + $signed(_zz_13405));
  assign _zz_3466 = 1'b1;
  assign _zz_3467 = 1'b1;
  assign _zz_5044 = ($signed(_zz_13423) * $signed(_zz_1375));
  assign _zz_3470 = _zz_13424[15 : 0];
  assign _zz_5045 = ($signed(_zz_13425) * $signed(twiddle_factor_table_46_real));
  assign _zz_5046 = ($signed(_zz_13426) * $signed(twiddle_factor_table_46_imag));
  assign _zz_3468 = ($signed(_zz_3470) - $signed(_zz_13427));
  assign _zz_3469 = ($signed(_zz_3470) + $signed(_zz_13429));
  assign _zz_3471 = 1'b1;
  assign _zz_3472 = 1'b1;
  assign _zz_5047 = ($signed(_zz_13447) * $signed(_zz_1377));
  assign _zz_3475 = _zz_13448[15 : 0];
  assign _zz_5048 = ($signed(_zz_13449) * $signed(twiddle_factor_table_47_real));
  assign _zz_5049 = ($signed(_zz_13450) * $signed(twiddle_factor_table_47_imag));
  assign _zz_3473 = ($signed(_zz_3475) - $signed(_zz_13451));
  assign _zz_3474 = ($signed(_zz_3475) + $signed(_zz_13453));
  assign _zz_3476 = 1'b1;
  assign _zz_3477 = 1'b1;
  assign _zz_5050 = ($signed(_zz_13471) * $signed(_zz_1379));
  assign _zz_3480 = _zz_13472[15 : 0];
  assign _zz_5051 = ($signed(_zz_13473) * $signed(twiddle_factor_table_48_real));
  assign _zz_5052 = ($signed(_zz_13474) * $signed(twiddle_factor_table_48_imag));
  assign _zz_3478 = ($signed(_zz_3480) - $signed(_zz_13475));
  assign _zz_3479 = ($signed(_zz_3480) + $signed(_zz_13477));
  assign _zz_3481 = 1'b1;
  assign _zz_3482 = 1'b1;
  assign _zz_5053 = ($signed(_zz_13495) * $signed(_zz_1381));
  assign _zz_3485 = _zz_13496[15 : 0];
  assign _zz_5054 = ($signed(_zz_13497) * $signed(twiddle_factor_table_49_real));
  assign _zz_5055 = ($signed(_zz_13498) * $signed(twiddle_factor_table_49_imag));
  assign _zz_3483 = ($signed(_zz_3485) - $signed(_zz_13499));
  assign _zz_3484 = ($signed(_zz_3485) + $signed(_zz_13501));
  assign _zz_3486 = 1'b1;
  assign _zz_3487 = 1'b1;
  assign _zz_5056 = ($signed(_zz_13519) * $signed(_zz_1383));
  assign _zz_3490 = _zz_13520[15 : 0];
  assign _zz_5057 = ($signed(_zz_13521) * $signed(twiddle_factor_table_50_real));
  assign _zz_5058 = ($signed(_zz_13522) * $signed(twiddle_factor_table_50_imag));
  assign _zz_3488 = ($signed(_zz_3490) - $signed(_zz_13523));
  assign _zz_3489 = ($signed(_zz_3490) + $signed(_zz_13525));
  assign _zz_3491 = 1'b1;
  assign _zz_3492 = 1'b1;
  assign _zz_5059 = ($signed(_zz_13543) * $signed(_zz_1385));
  assign _zz_3495 = _zz_13544[15 : 0];
  assign _zz_5060 = ($signed(_zz_13545) * $signed(twiddle_factor_table_51_real));
  assign _zz_5061 = ($signed(_zz_13546) * $signed(twiddle_factor_table_51_imag));
  assign _zz_3493 = ($signed(_zz_3495) - $signed(_zz_13547));
  assign _zz_3494 = ($signed(_zz_3495) + $signed(_zz_13549));
  assign _zz_3496 = 1'b1;
  assign _zz_3497 = 1'b1;
  assign _zz_5062 = ($signed(_zz_13567) * $signed(_zz_1387));
  assign _zz_3500 = _zz_13568[15 : 0];
  assign _zz_5063 = ($signed(_zz_13569) * $signed(twiddle_factor_table_52_real));
  assign _zz_5064 = ($signed(_zz_13570) * $signed(twiddle_factor_table_52_imag));
  assign _zz_3498 = ($signed(_zz_3500) - $signed(_zz_13571));
  assign _zz_3499 = ($signed(_zz_3500) + $signed(_zz_13573));
  assign _zz_3501 = 1'b1;
  assign _zz_3502 = 1'b1;
  assign _zz_5065 = ($signed(_zz_13591) * $signed(_zz_1389));
  assign _zz_3505 = _zz_13592[15 : 0];
  assign _zz_5066 = ($signed(_zz_13593) * $signed(twiddle_factor_table_53_real));
  assign _zz_5067 = ($signed(_zz_13594) * $signed(twiddle_factor_table_53_imag));
  assign _zz_3503 = ($signed(_zz_3505) - $signed(_zz_13595));
  assign _zz_3504 = ($signed(_zz_3505) + $signed(_zz_13597));
  assign _zz_3506 = 1'b1;
  assign _zz_3507 = 1'b1;
  assign _zz_5068 = ($signed(_zz_13615) * $signed(_zz_1391));
  assign _zz_3510 = _zz_13616[15 : 0];
  assign _zz_5069 = ($signed(_zz_13617) * $signed(twiddle_factor_table_54_real));
  assign _zz_5070 = ($signed(_zz_13618) * $signed(twiddle_factor_table_54_imag));
  assign _zz_3508 = ($signed(_zz_3510) - $signed(_zz_13619));
  assign _zz_3509 = ($signed(_zz_3510) + $signed(_zz_13621));
  assign _zz_3511 = 1'b1;
  assign _zz_3512 = 1'b1;
  assign _zz_5071 = ($signed(_zz_13639) * $signed(_zz_1393));
  assign _zz_3515 = _zz_13640[15 : 0];
  assign _zz_5072 = ($signed(_zz_13641) * $signed(twiddle_factor_table_55_real));
  assign _zz_5073 = ($signed(_zz_13642) * $signed(twiddle_factor_table_55_imag));
  assign _zz_3513 = ($signed(_zz_3515) - $signed(_zz_13643));
  assign _zz_3514 = ($signed(_zz_3515) + $signed(_zz_13645));
  assign _zz_3516 = 1'b1;
  assign _zz_3517 = 1'b1;
  assign _zz_5074 = ($signed(_zz_13663) * $signed(_zz_1395));
  assign _zz_3520 = _zz_13664[15 : 0];
  assign _zz_5075 = ($signed(_zz_13665) * $signed(twiddle_factor_table_56_real));
  assign _zz_5076 = ($signed(_zz_13666) * $signed(twiddle_factor_table_56_imag));
  assign _zz_3518 = ($signed(_zz_3520) - $signed(_zz_13667));
  assign _zz_3519 = ($signed(_zz_3520) + $signed(_zz_13669));
  assign _zz_3521 = 1'b1;
  assign _zz_3522 = 1'b1;
  assign _zz_5077 = ($signed(_zz_13687) * $signed(_zz_1397));
  assign _zz_3525 = _zz_13688[15 : 0];
  assign _zz_5078 = ($signed(_zz_13689) * $signed(twiddle_factor_table_57_real));
  assign _zz_5079 = ($signed(_zz_13690) * $signed(twiddle_factor_table_57_imag));
  assign _zz_3523 = ($signed(_zz_3525) - $signed(_zz_13691));
  assign _zz_3524 = ($signed(_zz_3525) + $signed(_zz_13693));
  assign _zz_3526 = 1'b1;
  assign _zz_3527 = 1'b1;
  assign _zz_5080 = ($signed(_zz_13711) * $signed(_zz_1399));
  assign _zz_3530 = _zz_13712[15 : 0];
  assign _zz_5081 = ($signed(_zz_13713) * $signed(twiddle_factor_table_58_real));
  assign _zz_5082 = ($signed(_zz_13714) * $signed(twiddle_factor_table_58_imag));
  assign _zz_3528 = ($signed(_zz_3530) - $signed(_zz_13715));
  assign _zz_3529 = ($signed(_zz_3530) + $signed(_zz_13717));
  assign _zz_3531 = 1'b1;
  assign _zz_3532 = 1'b1;
  assign _zz_5083 = ($signed(_zz_13735) * $signed(_zz_1401));
  assign _zz_3535 = _zz_13736[15 : 0];
  assign _zz_5084 = ($signed(_zz_13737) * $signed(twiddle_factor_table_59_real));
  assign _zz_5085 = ($signed(_zz_13738) * $signed(twiddle_factor_table_59_imag));
  assign _zz_3533 = ($signed(_zz_3535) - $signed(_zz_13739));
  assign _zz_3534 = ($signed(_zz_3535) + $signed(_zz_13741));
  assign _zz_3536 = 1'b1;
  assign _zz_3537 = 1'b1;
  assign _zz_5086 = ($signed(_zz_13759) * $signed(_zz_1403));
  assign _zz_3540 = _zz_13760[15 : 0];
  assign _zz_5087 = ($signed(_zz_13761) * $signed(twiddle_factor_table_60_real));
  assign _zz_5088 = ($signed(_zz_13762) * $signed(twiddle_factor_table_60_imag));
  assign _zz_3538 = ($signed(_zz_3540) - $signed(_zz_13763));
  assign _zz_3539 = ($signed(_zz_3540) + $signed(_zz_13765));
  assign _zz_3541 = 1'b1;
  assign _zz_3542 = 1'b1;
  assign _zz_5089 = ($signed(_zz_13783) * $signed(_zz_1405));
  assign _zz_3545 = _zz_13784[15 : 0];
  assign _zz_5090 = ($signed(_zz_13785) * $signed(twiddle_factor_table_61_real));
  assign _zz_5091 = ($signed(_zz_13786) * $signed(twiddle_factor_table_61_imag));
  assign _zz_3543 = ($signed(_zz_3545) - $signed(_zz_13787));
  assign _zz_3544 = ($signed(_zz_3545) + $signed(_zz_13789));
  assign _zz_3546 = 1'b1;
  assign _zz_3547 = 1'b1;
  assign _zz_5092 = ($signed(_zz_13807) * $signed(_zz_1407));
  assign _zz_3550 = _zz_13808[15 : 0];
  assign _zz_5093 = ($signed(_zz_13809) * $signed(twiddle_factor_table_62_real));
  assign _zz_5094 = ($signed(_zz_13810) * $signed(twiddle_factor_table_62_imag));
  assign _zz_3548 = ($signed(_zz_3550) - $signed(_zz_13811));
  assign _zz_3549 = ($signed(_zz_3550) + $signed(_zz_13813));
  assign _zz_3551 = 1'b1;
  assign _zz_3552 = 1'b1;
  assign _zz_5095 = ($signed(_zz_13831) * $signed(_zz_1473));
  assign _zz_3555 = _zz_13832[15 : 0];
  assign _zz_5096 = ($signed(_zz_13833) * $signed(twiddle_factor_table_31_real));
  assign _zz_5097 = ($signed(_zz_13834) * $signed(twiddle_factor_table_31_imag));
  assign _zz_3553 = ($signed(_zz_3555) - $signed(_zz_13835));
  assign _zz_3554 = ($signed(_zz_3555) + $signed(_zz_13837));
  assign _zz_3556 = 1'b1;
  assign _zz_3557 = 1'b1;
  assign _zz_5098 = ($signed(_zz_13855) * $signed(_zz_1475));
  assign _zz_3560 = _zz_13856[15 : 0];
  assign _zz_5099 = ($signed(_zz_13857) * $signed(twiddle_factor_table_32_real));
  assign _zz_5100 = ($signed(_zz_13858) * $signed(twiddle_factor_table_32_imag));
  assign _zz_3558 = ($signed(_zz_3560) - $signed(_zz_13859));
  assign _zz_3559 = ($signed(_zz_3560) + $signed(_zz_13861));
  assign _zz_3561 = 1'b1;
  assign _zz_3562 = 1'b1;
  assign _zz_5101 = ($signed(_zz_13879) * $signed(_zz_1477));
  assign _zz_3565 = _zz_13880[15 : 0];
  assign _zz_5102 = ($signed(_zz_13881) * $signed(twiddle_factor_table_33_real));
  assign _zz_5103 = ($signed(_zz_13882) * $signed(twiddle_factor_table_33_imag));
  assign _zz_3563 = ($signed(_zz_3565) - $signed(_zz_13883));
  assign _zz_3564 = ($signed(_zz_3565) + $signed(_zz_13885));
  assign _zz_3566 = 1'b1;
  assign _zz_3567 = 1'b1;
  assign _zz_5104 = ($signed(_zz_13903) * $signed(_zz_1479));
  assign _zz_3570 = _zz_13904[15 : 0];
  assign _zz_5105 = ($signed(_zz_13905) * $signed(twiddle_factor_table_34_real));
  assign _zz_5106 = ($signed(_zz_13906) * $signed(twiddle_factor_table_34_imag));
  assign _zz_3568 = ($signed(_zz_3570) - $signed(_zz_13907));
  assign _zz_3569 = ($signed(_zz_3570) + $signed(_zz_13909));
  assign _zz_3571 = 1'b1;
  assign _zz_3572 = 1'b1;
  assign _zz_5107 = ($signed(_zz_13927) * $signed(_zz_1481));
  assign _zz_3575 = _zz_13928[15 : 0];
  assign _zz_5108 = ($signed(_zz_13929) * $signed(twiddle_factor_table_35_real));
  assign _zz_5109 = ($signed(_zz_13930) * $signed(twiddle_factor_table_35_imag));
  assign _zz_3573 = ($signed(_zz_3575) - $signed(_zz_13931));
  assign _zz_3574 = ($signed(_zz_3575) + $signed(_zz_13933));
  assign _zz_3576 = 1'b1;
  assign _zz_3577 = 1'b1;
  assign _zz_5110 = ($signed(_zz_13951) * $signed(_zz_1483));
  assign _zz_3580 = _zz_13952[15 : 0];
  assign _zz_5111 = ($signed(_zz_13953) * $signed(twiddle_factor_table_36_real));
  assign _zz_5112 = ($signed(_zz_13954) * $signed(twiddle_factor_table_36_imag));
  assign _zz_3578 = ($signed(_zz_3580) - $signed(_zz_13955));
  assign _zz_3579 = ($signed(_zz_3580) + $signed(_zz_13957));
  assign _zz_3581 = 1'b1;
  assign _zz_3582 = 1'b1;
  assign _zz_5113 = ($signed(_zz_13975) * $signed(_zz_1485));
  assign _zz_3585 = _zz_13976[15 : 0];
  assign _zz_5114 = ($signed(_zz_13977) * $signed(twiddle_factor_table_37_real));
  assign _zz_5115 = ($signed(_zz_13978) * $signed(twiddle_factor_table_37_imag));
  assign _zz_3583 = ($signed(_zz_3585) - $signed(_zz_13979));
  assign _zz_3584 = ($signed(_zz_3585) + $signed(_zz_13981));
  assign _zz_3586 = 1'b1;
  assign _zz_3587 = 1'b1;
  assign _zz_5116 = ($signed(_zz_13999) * $signed(_zz_1487));
  assign _zz_3590 = _zz_14000[15 : 0];
  assign _zz_5117 = ($signed(_zz_14001) * $signed(twiddle_factor_table_38_real));
  assign _zz_5118 = ($signed(_zz_14002) * $signed(twiddle_factor_table_38_imag));
  assign _zz_3588 = ($signed(_zz_3590) - $signed(_zz_14003));
  assign _zz_3589 = ($signed(_zz_3590) + $signed(_zz_14005));
  assign _zz_3591 = 1'b1;
  assign _zz_3592 = 1'b1;
  assign _zz_5119 = ($signed(_zz_14023) * $signed(_zz_1489));
  assign _zz_3595 = _zz_14024[15 : 0];
  assign _zz_5120 = ($signed(_zz_14025) * $signed(twiddle_factor_table_39_real));
  assign _zz_5121 = ($signed(_zz_14026) * $signed(twiddle_factor_table_39_imag));
  assign _zz_3593 = ($signed(_zz_3595) - $signed(_zz_14027));
  assign _zz_3594 = ($signed(_zz_3595) + $signed(_zz_14029));
  assign _zz_3596 = 1'b1;
  assign _zz_3597 = 1'b1;
  assign _zz_5122 = ($signed(_zz_14047) * $signed(_zz_1491));
  assign _zz_3600 = _zz_14048[15 : 0];
  assign _zz_5123 = ($signed(_zz_14049) * $signed(twiddle_factor_table_40_real));
  assign _zz_5124 = ($signed(_zz_14050) * $signed(twiddle_factor_table_40_imag));
  assign _zz_3598 = ($signed(_zz_3600) - $signed(_zz_14051));
  assign _zz_3599 = ($signed(_zz_3600) + $signed(_zz_14053));
  assign _zz_3601 = 1'b1;
  assign _zz_3602 = 1'b1;
  assign _zz_5125 = ($signed(_zz_14071) * $signed(_zz_1493));
  assign _zz_3605 = _zz_14072[15 : 0];
  assign _zz_5126 = ($signed(_zz_14073) * $signed(twiddle_factor_table_41_real));
  assign _zz_5127 = ($signed(_zz_14074) * $signed(twiddle_factor_table_41_imag));
  assign _zz_3603 = ($signed(_zz_3605) - $signed(_zz_14075));
  assign _zz_3604 = ($signed(_zz_3605) + $signed(_zz_14077));
  assign _zz_3606 = 1'b1;
  assign _zz_3607 = 1'b1;
  assign _zz_5128 = ($signed(_zz_14095) * $signed(_zz_1495));
  assign _zz_3610 = _zz_14096[15 : 0];
  assign _zz_5129 = ($signed(_zz_14097) * $signed(twiddle_factor_table_42_real));
  assign _zz_5130 = ($signed(_zz_14098) * $signed(twiddle_factor_table_42_imag));
  assign _zz_3608 = ($signed(_zz_3610) - $signed(_zz_14099));
  assign _zz_3609 = ($signed(_zz_3610) + $signed(_zz_14101));
  assign _zz_3611 = 1'b1;
  assign _zz_3612 = 1'b1;
  assign _zz_5131 = ($signed(_zz_14119) * $signed(_zz_1497));
  assign _zz_3615 = _zz_14120[15 : 0];
  assign _zz_5132 = ($signed(_zz_14121) * $signed(twiddle_factor_table_43_real));
  assign _zz_5133 = ($signed(_zz_14122) * $signed(twiddle_factor_table_43_imag));
  assign _zz_3613 = ($signed(_zz_3615) - $signed(_zz_14123));
  assign _zz_3614 = ($signed(_zz_3615) + $signed(_zz_14125));
  assign _zz_3616 = 1'b1;
  assign _zz_3617 = 1'b1;
  assign _zz_5134 = ($signed(_zz_14143) * $signed(_zz_1499));
  assign _zz_3620 = _zz_14144[15 : 0];
  assign _zz_5135 = ($signed(_zz_14145) * $signed(twiddle_factor_table_44_real));
  assign _zz_5136 = ($signed(_zz_14146) * $signed(twiddle_factor_table_44_imag));
  assign _zz_3618 = ($signed(_zz_3620) - $signed(_zz_14147));
  assign _zz_3619 = ($signed(_zz_3620) + $signed(_zz_14149));
  assign _zz_3621 = 1'b1;
  assign _zz_3622 = 1'b1;
  assign _zz_5137 = ($signed(_zz_14167) * $signed(_zz_1501));
  assign _zz_3625 = _zz_14168[15 : 0];
  assign _zz_5138 = ($signed(_zz_14169) * $signed(twiddle_factor_table_45_real));
  assign _zz_5139 = ($signed(_zz_14170) * $signed(twiddle_factor_table_45_imag));
  assign _zz_3623 = ($signed(_zz_3625) - $signed(_zz_14171));
  assign _zz_3624 = ($signed(_zz_3625) + $signed(_zz_14173));
  assign _zz_3626 = 1'b1;
  assign _zz_3627 = 1'b1;
  assign _zz_5140 = ($signed(_zz_14191) * $signed(_zz_1503));
  assign _zz_3630 = _zz_14192[15 : 0];
  assign _zz_5141 = ($signed(_zz_14193) * $signed(twiddle_factor_table_46_real));
  assign _zz_5142 = ($signed(_zz_14194) * $signed(twiddle_factor_table_46_imag));
  assign _zz_3628 = ($signed(_zz_3630) - $signed(_zz_14195));
  assign _zz_3629 = ($signed(_zz_3630) + $signed(_zz_14197));
  assign _zz_3631 = 1'b1;
  assign _zz_3632 = 1'b1;
  assign _zz_5143 = ($signed(_zz_14215) * $signed(_zz_1505));
  assign _zz_3635 = _zz_14216[15 : 0];
  assign _zz_5144 = ($signed(_zz_14217) * $signed(twiddle_factor_table_47_real));
  assign _zz_5145 = ($signed(_zz_14218) * $signed(twiddle_factor_table_47_imag));
  assign _zz_3633 = ($signed(_zz_3635) - $signed(_zz_14219));
  assign _zz_3634 = ($signed(_zz_3635) + $signed(_zz_14221));
  assign _zz_3636 = 1'b1;
  assign _zz_3637 = 1'b1;
  assign _zz_5146 = ($signed(_zz_14239) * $signed(_zz_1507));
  assign _zz_3640 = _zz_14240[15 : 0];
  assign _zz_5147 = ($signed(_zz_14241) * $signed(twiddle_factor_table_48_real));
  assign _zz_5148 = ($signed(_zz_14242) * $signed(twiddle_factor_table_48_imag));
  assign _zz_3638 = ($signed(_zz_3640) - $signed(_zz_14243));
  assign _zz_3639 = ($signed(_zz_3640) + $signed(_zz_14245));
  assign _zz_3641 = 1'b1;
  assign _zz_3642 = 1'b1;
  assign _zz_5149 = ($signed(_zz_14263) * $signed(_zz_1509));
  assign _zz_3645 = _zz_14264[15 : 0];
  assign _zz_5150 = ($signed(_zz_14265) * $signed(twiddle_factor_table_49_real));
  assign _zz_5151 = ($signed(_zz_14266) * $signed(twiddle_factor_table_49_imag));
  assign _zz_3643 = ($signed(_zz_3645) - $signed(_zz_14267));
  assign _zz_3644 = ($signed(_zz_3645) + $signed(_zz_14269));
  assign _zz_3646 = 1'b1;
  assign _zz_3647 = 1'b1;
  assign _zz_5152 = ($signed(_zz_14287) * $signed(_zz_1511));
  assign _zz_3650 = _zz_14288[15 : 0];
  assign _zz_5153 = ($signed(_zz_14289) * $signed(twiddle_factor_table_50_real));
  assign _zz_5154 = ($signed(_zz_14290) * $signed(twiddle_factor_table_50_imag));
  assign _zz_3648 = ($signed(_zz_3650) - $signed(_zz_14291));
  assign _zz_3649 = ($signed(_zz_3650) + $signed(_zz_14293));
  assign _zz_3651 = 1'b1;
  assign _zz_3652 = 1'b1;
  assign _zz_5155 = ($signed(_zz_14311) * $signed(_zz_1513));
  assign _zz_3655 = _zz_14312[15 : 0];
  assign _zz_5156 = ($signed(_zz_14313) * $signed(twiddle_factor_table_51_real));
  assign _zz_5157 = ($signed(_zz_14314) * $signed(twiddle_factor_table_51_imag));
  assign _zz_3653 = ($signed(_zz_3655) - $signed(_zz_14315));
  assign _zz_3654 = ($signed(_zz_3655) + $signed(_zz_14317));
  assign _zz_3656 = 1'b1;
  assign _zz_3657 = 1'b1;
  assign _zz_5158 = ($signed(_zz_14335) * $signed(_zz_1515));
  assign _zz_3660 = _zz_14336[15 : 0];
  assign _zz_5159 = ($signed(_zz_14337) * $signed(twiddle_factor_table_52_real));
  assign _zz_5160 = ($signed(_zz_14338) * $signed(twiddle_factor_table_52_imag));
  assign _zz_3658 = ($signed(_zz_3660) - $signed(_zz_14339));
  assign _zz_3659 = ($signed(_zz_3660) + $signed(_zz_14341));
  assign _zz_3661 = 1'b1;
  assign _zz_3662 = 1'b1;
  assign _zz_5161 = ($signed(_zz_14359) * $signed(_zz_1517));
  assign _zz_3665 = _zz_14360[15 : 0];
  assign _zz_5162 = ($signed(_zz_14361) * $signed(twiddle_factor_table_53_real));
  assign _zz_5163 = ($signed(_zz_14362) * $signed(twiddle_factor_table_53_imag));
  assign _zz_3663 = ($signed(_zz_3665) - $signed(_zz_14363));
  assign _zz_3664 = ($signed(_zz_3665) + $signed(_zz_14365));
  assign _zz_3666 = 1'b1;
  assign _zz_3667 = 1'b1;
  assign _zz_5164 = ($signed(_zz_14383) * $signed(_zz_1519));
  assign _zz_3670 = _zz_14384[15 : 0];
  assign _zz_5165 = ($signed(_zz_14385) * $signed(twiddle_factor_table_54_real));
  assign _zz_5166 = ($signed(_zz_14386) * $signed(twiddle_factor_table_54_imag));
  assign _zz_3668 = ($signed(_zz_3670) - $signed(_zz_14387));
  assign _zz_3669 = ($signed(_zz_3670) + $signed(_zz_14389));
  assign _zz_3671 = 1'b1;
  assign _zz_3672 = 1'b1;
  assign _zz_5167 = ($signed(_zz_14407) * $signed(_zz_1521));
  assign _zz_3675 = _zz_14408[15 : 0];
  assign _zz_5168 = ($signed(_zz_14409) * $signed(twiddle_factor_table_55_real));
  assign _zz_5169 = ($signed(_zz_14410) * $signed(twiddle_factor_table_55_imag));
  assign _zz_3673 = ($signed(_zz_3675) - $signed(_zz_14411));
  assign _zz_3674 = ($signed(_zz_3675) + $signed(_zz_14413));
  assign _zz_3676 = 1'b1;
  assign _zz_3677 = 1'b1;
  assign _zz_5170 = ($signed(_zz_14431) * $signed(_zz_1523));
  assign _zz_3680 = _zz_14432[15 : 0];
  assign _zz_5171 = ($signed(_zz_14433) * $signed(twiddle_factor_table_56_real));
  assign _zz_5172 = ($signed(_zz_14434) * $signed(twiddle_factor_table_56_imag));
  assign _zz_3678 = ($signed(_zz_3680) - $signed(_zz_14435));
  assign _zz_3679 = ($signed(_zz_3680) + $signed(_zz_14437));
  assign _zz_3681 = 1'b1;
  assign _zz_3682 = 1'b1;
  assign _zz_5173 = ($signed(_zz_14455) * $signed(_zz_1525));
  assign _zz_3685 = _zz_14456[15 : 0];
  assign _zz_5174 = ($signed(_zz_14457) * $signed(twiddle_factor_table_57_real));
  assign _zz_5175 = ($signed(_zz_14458) * $signed(twiddle_factor_table_57_imag));
  assign _zz_3683 = ($signed(_zz_3685) - $signed(_zz_14459));
  assign _zz_3684 = ($signed(_zz_3685) + $signed(_zz_14461));
  assign _zz_3686 = 1'b1;
  assign _zz_3687 = 1'b1;
  assign _zz_5176 = ($signed(_zz_14479) * $signed(_zz_1527));
  assign _zz_3690 = _zz_14480[15 : 0];
  assign _zz_5177 = ($signed(_zz_14481) * $signed(twiddle_factor_table_58_real));
  assign _zz_5178 = ($signed(_zz_14482) * $signed(twiddle_factor_table_58_imag));
  assign _zz_3688 = ($signed(_zz_3690) - $signed(_zz_14483));
  assign _zz_3689 = ($signed(_zz_3690) + $signed(_zz_14485));
  assign _zz_3691 = 1'b1;
  assign _zz_3692 = 1'b1;
  assign _zz_5179 = ($signed(_zz_14503) * $signed(_zz_1529));
  assign _zz_3695 = _zz_14504[15 : 0];
  assign _zz_5180 = ($signed(_zz_14505) * $signed(twiddle_factor_table_59_real));
  assign _zz_5181 = ($signed(_zz_14506) * $signed(twiddle_factor_table_59_imag));
  assign _zz_3693 = ($signed(_zz_3695) - $signed(_zz_14507));
  assign _zz_3694 = ($signed(_zz_3695) + $signed(_zz_14509));
  assign _zz_3696 = 1'b1;
  assign _zz_3697 = 1'b1;
  assign _zz_5182 = ($signed(_zz_14527) * $signed(_zz_1531));
  assign _zz_3700 = _zz_14528[15 : 0];
  assign _zz_5183 = ($signed(_zz_14529) * $signed(twiddle_factor_table_60_real));
  assign _zz_5184 = ($signed(_zz_14530) * $signed(twiddle_factor_table_60_imag));
  assign _zz_3698 = ($signed(_zz_3700) - $signed(_zz_14531));
  assign _zz_3699 = ($signed(_zz_3700) + $signed(_zz_14533));
  assign _zz_3701 = 1'b1;
  assign _zz_3702 = 1'b1;
  assign _zz_5185 = ($signed(_zz_14551) * $signed(_zz_1533));
  assign _zz_3705 = _zz_14552[15 : 0];
  assign _zz_5186 = ($signed(_zz_14553) * $signed(twiddle_factor_table_61_real));
  assign _zz_5187 = ($signed(_zz_14554) * $signed(twiddle_factor_table_61_imag));
  assign _zz_3703 = ($signed(_zz_3705) - $signed(_zz_14555));
  assign _zz_3704 = ($signed(_zz_3705) + $signed(_zz_14557));
  assign _zz_3706 = 1'b1;
  assign _zz_3707 = 1'b1;
  assign _zz_5188 = ($signed(_zz_14575) * $signed(_zz_1535));
  assign _zz_3710 = _zz_14576[15 : 0];
  assign _zz_5189 = ($signed(_zz_14577) * $signed(twiddle_factor_table_62_real));
  assign _zz_5190 = ($signed(_zz_14578) * $signed(twiddle_factor_table_62_imag));
  assign _zz_3708 = ($signed(_zz_3710) - $signed(_zz_14579));
  assign _zz_3709 = ($signed(_zz_3710) + $signed(_zz_14581));
  assign _zz_3711 = 1'b1;
  assign _zz_3712 = 1'b1;
  assign _zz_5191 = ($signed(_zz_14599) * $signed(_zz_1665));
  assign _zz_3715 = _zz_14600[15 : 0];
  assign _zz_5192 = ($signed(_zz_14601) * $signed(twiddle_factor_table_63_real));
  assign _zz_5193 = ($signed(_zz_14602) * $signed(twiddle_factor_table_63_imag));
  assign _zz_3713 = ($signed(_zz_3715) - $signed(_zz_14603));
  assign _zz_3714 = ($signed(_zz_3715) + $signed(_zz_14605));
  assign _zz_3716 = 1'b1;
  assign _zz_3717 = 1'b1;
  assign _zz_5194 = ($signed(_zz_14623) * $signed(_zz_1667));
  assign _zz_3720 = _zz_14624[15 : 0];
  assign _zz_5195 = ($signed(_zz_14625) * $signed(twiddle_factor_table_64_real));
  assign _zz_5196 = ($signed(_zz_14626) * $signed(twiddle_factor_table_64_imag));
  assign _zz_3718 = ($signed(_zz_3720) - $signed(_zz_14627));
  assign _zz_3719 = ($signed(_zz_3720) + $signed(_zz_14629));
  assign _zz_3721 = 1'b1;
  assign _zz_3722 = 1'b1;
  assign _zz_5197 = ($signed(_zz_14647) * $signed(_zz_1669));
  assign _zz_3725 = _zz_14648[15 : 0];
  assign _zz_5198 = ($signed(_zz_14649) * $signed(twiddle_factor_table_65_real));
  assign _zz_5199 = ($signed(_zz_14650) * $signed(twiddle_factor_table_65_imag));
  assign _zz_3723 = ($signed(_zz_3725) - $signed(_zz_14651));
  assign _zz_3724 = ($signed(_zz_3725) + $signed(_zz_14653));
  assign _zz_3726 = 1'b1;
  assign _zz_3727 = 1'b1;
  assign _zz_5200 = ($signed(_zz_14671) * $signed(_zz_1671));
  assign _zz_3730 = _zz_14672[15 : 0];
  assign _zz_5201 = ($signed(_zz_14673) * $signed(twiddle_factor_table_66_real));
  assign _zz_5202 = ($signed(_zz_14674) * $signed(twiddle_factor_table_66_imag));
  assign _zz_3728 = ($signed(_zz_3730) - $signed(_zz_14675));
  assign _zz_3729 = ($signed(_zz_3730) + $signed(_zz_14677));
  assign _zz_3731 = 1'b1;
  assign _zz_3732 = 1'b1;
  assign _zz_5203 = ($signed(_zz_14695) * $signed(_zz_1673));
  assign _zz_3735 = _zz_14696[15 : 0];
  assign _zz_5204 = ($signed(_zz_14697) * $signed(twiddle_factor_table_67_real));
  assign _zz_5205 = ($signed(_zz_14698) * $signed(twiddle_factor_table_67_imag));
  assign _zz_3733 = ($signed(_zz_3735) - $signed(_zz_14699));
  assign _zz_3734 = ($signed(_zz_3735) + $signed(_zz_14701));
  assign _zz_3736 = 1'b1;
  assign _zz_3737 = 1'b1;
  assign _zz_5206 = ($signed(_zz_14719) * $signed(_zz_1675));
  assign _zz_3740 = _zz_14720[15 : 0];
  assign _zz_5207 = ($signed(_zz_14721) * $signed(twiddle_factor_table_68_real));
  assign _zz_5208 = ($signed(_zz_14722) * $signed(twiddle_factor_table_68_imag));
  assign _zz_3738 = ($signed(_zz_3740) - $signed(_zz_14723));
  assign _zz_3739 = ($signed(_zz_3740) + $signed(_zz_14725));
  assign _zz_3741 = 1'b1;
  assign _zz_3742 = 1'b1;
  assign _zz_5209 = ($signed(_zz_14743) * $signed(_zz_1677));
  assign _zz_3745 = _zz_14744[15 : 0];
  assign _zz_5210 = ($signed(_zz_14745) * $signed(twiddle_factor_table_69_real));
  assign _zz_5211 = ($signed(_zz_14746) * $signed(twiddle_factor_table_69_imag));
  assign _zz_3743 = ($signed(_zz_3745) - $signed(_zz_14747));
  assign _zz_3744 = ($signed(_zz_3745) + $signed(_zz_14749));
  assign _zz_3746 = 1'b1;
  assign _zz_3747 = 1'b1;
  assign _zz_5212 = ($signed(_zz_14767) * $signed(_zz_1679));
  assign _zz_3750 = _zz_14768[15 : 0];
  assign _zz_5213 = ($signed(_zz_14769) * $signed(twiddle_factor_table_70_real));
  assign _zz_5214 = ($signed(_zz_14770) * $signed(twiddle_factor_table_70_imag));
  assign _zz_3748 = ($signed(_zz_3750) - $signed(_zz_14771));
  assign _zz_3749 = ($signed(_zz_3750) + $signed(_zz_14773));
  assign _zz_3751 = 1'b1;
  assign _zz_3752 = 1'b1;
  assign _zz_5215 = ($signed(_zz_14791) * $signed(_zz_1681));
  assign _zz_3755 = _zz_14792[15 : 0];
  assign _zz_5216 = ($signed(_zz_14793) * $signed(twiddle_factor_table_71_real));
  assign _zz_5217 = ($signed(_zz_14794) * $signed(twiddle_factor_table_71_imag));
  assign _zz_3753 = ($signed(_zz_3755) - $signed(_zz_14795));
  assign _zz_3754 = ($signed(_zz_3755) + $signed(_zz_14797));
  assign _zz_3756 = 1'b1;
  assign _zz_3757 = 1'b1;
  assign _zz_5218 = ($signed(_zz_14815) * $signed(_zz_1683));
  assign _zz_3760 = _zz_14816[15 : 0];
  assign _zz_5219 = ($signed(_zz_14817) * $signed(twiddle_factor_table_72_real));
  assign _zz_5220 = ($signed(_zz_14818) * $signed(twiddle_factor_table_72_imag));
  assign _zz_3758 = ($signed(_zz_3760) - $signed(_zz_14819));
  assign _zz_3759 = ($signed(_zz_3760) + $signed(_zz_14821));
  assign _zz_3761 = 1'b1;
  assign _zz_3762 = 1'b1;
  assign _zz_5221 = ($signed(_zz_14839) * $signed(_zz_1685));
  assign _zz_3765 = _zz_14840[15 : 0];
  assign _zz_5222 = ($signed(_zz_14841) * $signed(twiddle_factor_table_73_real));
  assign _zz_5223 = ($signed(_zz_14842) * $signed(twiddle_factor_table_73_imag));
  assign _zz_3763 = ($signed(_zz_3765) - $signed(_zz_14843));
  assign _zz_3764 = ($signed(_zz_3765) + $signed(_zz_14845));
  assign _zz_3766 = 1'b1;
  assign _zz_3767 = 1'b1;
  assign _zz_5224 = ($signed(_zz_14863) * $signed(_zz_1687));
  assign _zz_3770 = _zz_14864[15 : 0];
  assign _zz_5225 = ($signed(_zz_14865) * $signed(twiddle_factor_table_74_real));
  assign _zz_5226 = ($signed(_zz_14866) * $signed(twiddle_factor_table_74_imag));
  assign _zz_3768 = ($signed(_zz_3770) - $signed(_zz_14867));
  assign _zz_3769 = ($signed(_zz_3770) + $signed(_zz_14869));
  assign _zz_3771 = 1'b1;
  assign _zz_3772 = 1'b1;
  assign _zz_5227 = ($signed(_zz_14887) * $signed(_zz_1689));
  assign _zz_3775 = _zz_14888[15 : 0];
  assign _zz_5228 = ($signed(_zz_14889) * $signed(twiddle_factor_table_75_real));
  assign _zz_5229 = ($signed(_zz_14890) * $signed(twiddle_factor_table_75_imag));
  assign _zz_3773 = ($signed(_zz_3775) - $signed(_zz_14891));
  assign _zz_3774 = ($signed(_zz_3775) + $signed(_zz_14893));
  assign _zz_3776 = 1'b1;
  assign _zz_3777 = 1'b1;
  assign _zz_5230 = ($signed(_zz_14911) * $signed(_zz_1691));
  assign _zz_3780 = _zz_14912[15 : 0];
  assign _zz_5231 = ($signed(_zz_14913) * $signed(twiddle_factor_table_76_real));
  assign _zz_5232 = ($signed(_zz_14914) * $signed(twiddle_factor_table_76_imag));
  assign _zz_3778 = ($signed(_zz_3780) - $signed(_zz_14915));
  assign _zz_3779 = ($signed(_zz_3780) + $signed(_zz_14917));
  assign _zz_3781 = 1'b1;
  assign _zz_3782 = 1'b1;
  assign _zz_5233 = ($signed(_zz_14935) * $signed(_zz_1693));
  assign _zz_3785 = _zz_14936[15 : 0];
  assign _zz_5234 = ($signed(_zz_14937) * $signed(twiddle_factor_table_77_real));
  assign _zz_5235 = ($signed(_zz_14938) * $signed(twiddle_factor_table_77_imag));
  assign _zz_3783 = ($signed(_zz_3785) - $signed(_zz_14939));
  assign _zz_3784 = ($signed(_zz_3785) + $signed(_zz_14941));
  assign _zz_3786 = 1'b1;
  assign _zz_3787 = 1'b1;
  assign _zz_5236 = ($signed(_zz_14959) * $signed(_zz_1695));
  assign _zz_3790 = _zz_14960[15 : 0];
  assign _zz_5237 = ($signed(_zz_14961) * $signed(twiddle_factor_table_78_real));
  assign _zz_5238 = ($signed(_zz_14962) * $signed(twiddle_factor_table_78_imag));
  assign _zz_3788 = ($signed(_zz_3790) - $signed(_zz_14963));
  assign _zz_3789 = ($signed(_zz_3790) + $signed(_zz_14965));
  assign _zz_3791 = 1'b1;
  assign _zz_3792 = 1'b1;
  assign _zz_5239 = ($signed(_zz_14983) * $signed(_zz_1697));
  assign _zz_3795 = _zz_14984[15 : 0];
  assign _zz_5240 = ($signed(_zz_14985) * $signed(twiddle_factor_table_79_real));
  assign _zz_5241 = ($signed(_zz_14986) * $signed(twiddle_factor_table_79_imag));
  assign _zz_3793 = ($signed(_zz_3795) - $signed(_zz_14987));
  assign _zz_3794 = ($signed(_zz_3795) + $signed(_zz_14989));
  assign _zz_3796 = 1'b1;
  assign _zz_3797 = 1'b1;
  assign _zz_5242 = ($signed(_zz_15007) * $signed(_zz_1699));
  assign _zz_3800 = _zz_15008[15 : 0];
  assign _zz_5243 = ($signed(_zz_15009) * $signed(twiddle_factor_table_80_real));
  assign _zz_5244 = ($signed(_zz_15010) * $signed(twiddle_factor_table_80_imag));
  assign _zz_3798 = ($signed(_zz_3800) - $signed(_zz_15011));
  assign _zz_3799 = ($signed(_zz_3800) + $signed(_zz_15013));
  assign _zz_3801 = 1'b1;
  assign _zz_3802 = 1'b1;
  assign _zz_5245 = ($signed(_zz_15031) * $signed(_zz_1701));
  assign _zz_3805 = _zz_15032[15 : 0];
  assign _zz_5246 = ($signed(_zz_15033) * $signed(twiddle_factor_table_81_real));
  assign _zz_5247 = ($signed(_zz_15034) * $signed(twiddle_factor_table_81_imag));
  assign _zz_3803 = ($signed(_zz_3805) - $signed(_zz_15035));
  assign _zz_3804 = ($signed(_zz_3805) + $signed(_zz_15037));
  assign _zz_3806 = 1'b1;
  assign _zz_3807 = 1'b1;
  assign _zz_5248 = ($signed(_zz_15055) * $signed(_zz_1703));
  assign _zz_3810 = _zz_15056[15 : 0];
  assign _zz_5249 = ($signed(_zz_15057) * $signed(twiddle_factor_table_82_real));
  assign _zz_5250 = ($signed(_zz_15058) * $signed(twiddle_factor_table_82_imag));
  assign _zz_3808 = ($signed(_zz_3810) - $signed(_zz_15059));
  assign _zz_3809 = ($signed(_zz_3810) + $signed(_zz_15061));
  assign _zz_3811 = 1'b1;
  assign _zz_3812 = 1'b1;
  assign _zz_5251 = ($signed(_zz_15079) * $signed(_zz_1705));
  assign _zz_3815 = _zz_15080[15 : 0];
  assign _zz_5252 = ($signed(_zz_15081) * $signed(twiddle_factor_table_83_real));
  assign _zz_5253 = ($signed(_zz_15082) * $signed(twiddle_factor_table_83_imag));
  assign _zz_3813 = ($signed(_zz_3815) - $signed(_zz_15083));
  assign _zz_3814 = ($signed(_zz_3815) + $signed(_zz_15085));
  assign _zz_3816 = 1'b1;
  assign _zz_3817 = 1'b1;
  assign _zz_5254 = ($signed(_zz_15103) * $signed(_zz_1707));
  assign _zz_3820 = _zz_15104[15 : 0];
  assign _zz_5255 = ($signed(_zz_15105) * $signed(twiddle_factor_table_84_real));
  assign _zz_5256 = ($signed(_zz_15106) * $signed(twiddle_factor_table_84_imag));
  assign _zz_3818 = ($signed(_zz_3820) - $signed(_zz_15107));
  assign _zz_3819 = ($signed(_zz_3820) + $signed(_zz_15109));
  assign _zz_3821 = 1'b1;
  assign _zz_3822 = 1'b1;
  assign _zz_5257 = ($signed(_zz_15127) * $signed(_zz_1709));
  assign _zz_3825 = _zz_15128[15 : 0];
  assign _zz_5258 = ($signed(_zz_15129) * $signed(twiddle_factor_table_85_real));
  assign _zz_5259 = ($signed(_zz_15130) * $signed(twiddle_factor_table_85_imag));
  assign _zz_3823 = ($signed(_zz_3825) - $signed(_zz_15131));
  assign _zz_3824 = ($signed(_zz_3825) + $signed(_zz_15133));
  assign _zz_3826 = 1'b1;
  assign _zz_3827 = 1'b1;
  assign _zz_5260 = ($signed(_zz_15151) * $signed(_zz_1711));
  assign _zz_3830 = _zz_15152[15 : 0];
  assign _zz_5261 = ($signed(_zz_15153) * $signed(twiddle_factor_table_86_real));
  assign _zz_5262 = ($signed(_zz_15154) * $signed(twiddle_factor_table_86_imag));
  assign _zz_3828 = ($signed(_zz_3830) - $signed(_zz_15155));
  assign _zz_3829 = ($signed(_zz_3830) + $signed(_zz_15157));
  assign _zz_3831 = 1'b1;
  assign _zz_3832 = 1'b1;
  assign _zz_5263 = ($signed(_zz_15175) * $signed(_zz_1713));
  assign _zz_3835 = _zz_15176[15 : 0];
  assign _zz_5264 = ($signed(_zz_15177) * $signed(twiddle_factor_table_87_real));
  assign _zz_5265 = ($signed(_zz_15178) * $signed(twiddle_factor_table_87_imag));
  assign _zz_3833 = ($signed(_zz_3835) - $signed(_zz_15179));
  assign _zz_3834 = ($signed(_zz_3835) + $signed(_zz_15181));
  assign _zz_3836 = 1'b1;
  assign _zz_3837 = 1'b1;
  assign _zz_5266 = ($signed(_zz_15199) * $signed(_zz_1715));
  assign _zz_3840 = _zz_15200[15 : 0];
  assign _zz_5267 = ($signed(_zz_15201) * $signed(twiddle_factor_table_88_real));
  assign _zz_5268 = ($signed(_zz_15202) * $signed(twiddle_factor_table_88_imag));
  assign _zz_3838 = ($signed(_zz_3840) - $signed(_zz_15203));
  assign _zz_3839 = ($signed(_zz_3840) + $signed(_zz_15205));
  assign _zz_3841 = 1'b1;
  assign _zz_3842 = 1'b1;
  assign _zz_5269 = ($signed(_zz_15223) * $signed(_zz_1717));
  assign _zz_3845 = _zz_15224[15 : 0];
  assign _zz_5270 = ($signed(_zz_15225) * $signed(twiddle_factor_table_89_real));
  assign _zz_5271 = ($signed(_zz_15226) * $signed(twiddle_factor_table_89_imag));
  assign _zz_3843 = ($signed(_zz_3845) - $signed(_zz_15227));
  assign _zz_3844 = ($signed(_zz_3845) + $signed(_zz_15229));
  assign _zz_3846 = 1'b1;
  assign _zz_3847 = 1'b1;
  assign _zz_5272 = ($signed(_zz_15247) * $signed(_zz_1719));
  assign _zz_3850 = _zz_15248[15 : 0];
  assign _zz_5273 = ($signed(_zz_15249) * $signed(twiddle_factor_table_90_real));
  assign _zz_5274 = ($signed(_zz_15250) * $signed(twiddle_factor_table_90_imag));
  assign _zz_3848 = ($signed(_zz_3850) - $signed(_zz_15251));
  assign _zz_3849 = ($signed(_zz_3850) + $signed(_zz_15253));
  assign _zz_3851 = 1'b1;
  assign _zz_3852 = 1'b1;
  assign _zz_5275 = ($signed(_zz_15271) * $signed(_zz_1721));
  assign _zz_3855 = _zz_15272[15 : 0];
  assign _zz_5276 = ($signed(_zz_15273) * $signed(twiddle_factor_table_91_real));
  assign _zz_5277 = ($signed(_zz_15274) * $signed(twiddle_factor_table_91_imag));
  assign _zz_3853 = ($signed(_zz_3855) - $signed(_zz_15275));
  assign _zz_3854 = ($signed(_zz_3855) + $signed(_zz_15277));
  assign _zz_3856 = 1'b1;
  assign _zz_3857 = 1'b1;
  assign _zz_5278 = ($signed(_zz_15295) * $signed(_zz_1723));
  assign _zz_3860 = _zz_15296[15 : 0];
  assign _zz_5279 = ($signed(_zz_15297) * $signed(twiddle_factor_table_92_real));
  assign _zz_5280 = ($signed(_zz_15298) * $signed(twiddle_factor_table_92_imag));
  assign _zz_3858 = ($signed(_zz_3860) - $signed(_zz_15299));
  assign _zz_3859 = ($signed(_zz_3860) + $signed(_zz_15301));
  assign _zz_3861 = 1'b1;
  assign _zz_3862 = 1'b1;
  assign _zz_5281 = ($signed(_zz_15319) * $signed(_zz_1725));
  assign _zz_3865 = _zz_15320[15 : 0];
  assign _zz_5282 = ($signed(_zz_15321) * $signed(twiddle_factor_table_93_real));
  assign _zz_5283 = ($signed(_zz_15322) * $signed(twiddle_factor_table_93_imag));
  assign _zz_3863 = ($signed(_zz_3865) - $signed(_zz_15323));
  assign _zz_3864 = ($signed(_zz_3865) + $signed(_zz_15325));
  assign _zz_3866 = 1'b1;
  assign _zz_3867 = 1'b1;
  assign _zz_5284 = ($signed(_zz_15343) * $signed(_zz_1727));
  assign _zz_3870 = _zz_15344[15 : 0];
  assign _zz_5285 = ($signed(_zz_15345) * $signed(twiddle_factor_table_94_real));
  assign _zz_5286 = ($signed(_zz_15346) * $signed(twiddle_factor_table_94_imag));
  assign _zz_3868 = ($signed(_zz_3870) - $signed(_zz_15347));
  assign _zz_3869 = ($signed(_zz_3870) + $signed(_zz_15349));
  assign _zz_3871 = 1'b1;
  assign _zz_3872 = 1'b1;
  assign _zz_5287 = ($signed(_zz_15367) * $signed(_zz_1729));
  assign _zz_3875 = _zz_15368[15 : 0];
  assign _zz_5288 = ($signed(_zz_15369) * $signed(twiddle_factor_table_95_real));
  assign _zz_5289 = ($signed(_zz_15370) * $signed(twiddle_factor_table_95_imag));
  assign _zz_3873 = ($signed(_zz_3875) - $signed(_zz_15371));
  assign _zz_3874 = ($signed(_zz_3875) + $signed(_zz_15373));
  assign _zz_3876 = 1'b1;
  assign _zz_3877 = 1'b1;
  assign _zz_5290 = ($signed(_zz_15391) * $signed(_zz_1731));
  assign _zz_3880 = _zz_15392[15 : 0];
  assign _zz_5291 = ($signed(_zz_15393) * $signed(twiddle_factor_table_96_real));
  assign _zz_5292 = ($signed(_zz_15394) * $signed(twiddle_factor_table_96_imag));
  assign _zz_3878 = ($signed(_zz_3880) - $signed(_zz_15395));
  assign _zz_3879 = ($signed(_zz_3880) + $signed(_zz_15397));
  assign _zz_3881 = 1'b1;
  assign _zz_3882 = 1'b1;
  assign _zz_5293 = ($signed(_zz_15415) * $signed(_zz_1733));
  assign _zz_3885 = _zz_15416[15 : 0];
  assign _zz_5294 = ($signed(_zz_15417) * $signed(twiddle_factor_table_97_real));
  assign _zz_5295 = ($signed(_zz_15418) * $signed(twiddle_factor_table_97_imag));
  assign _zz_3883 = ($signed(_zz_3885) - $signed(_zz_15419));
  assign _zz_3884 = ($signed(_zz_3885) + $signed(_zz_15421));
  assign _zz_3886 = 1'b1;
  assign _zz_3887 = 1'b1;
  assign _zz_5296 = ($signed(_zz_15439) * $signed(_zz_1735));
  assign _zz_3890 = _zz_15440[15 : 0];
  assign _zz_5297 = ($signed(_zz_15441) * $signed(twiddle_factor_table_98_real));
  assign _zz_5298 = ($signed(_zz_15442) * $signed(twiddle_factor_table_98_imag));
  assign _zz_3888 = ($signed(_zz_3890) - $signed(_zz_15443));
  assign _zz_3889 = ($signed(_zz_3890) + $signed(_zz_15445));
  assign _zz_3891 = 1'b1;
  assign _zz_3892 = 1'b1;
  assign _zz_5299 = ($signed(_zz_15463) * $signed(_zz_1737));
  assign _zz_3895 = _zz_15464[15 : 0];
  assign _zz_5300 = ($signed(_zz_15465) * $signed(twiddle_factor_table_99_real));
  assign _zz_5301 = ($signed(_zz_15466) * $signed(twiddle_factor_table_99_imag));
  assign _zz_3893 = ($signed(_zz_3895) - $signed(_zz_15467));
  assign _zz_3894 = ($signed(_zz_3895) + $signed(_zz_15469));
  assign _zz_3896 = 1'b1;
  assign _zz_3897 = 1'b1;
  assign _zz_5302 = ($signed(_zz_15487) * $signed(_zz_1739));
  assign _zz_3900 = _zz_15488[15 : 0];
  assign _zz_5303 = ($signed(_zz_15489) * $signed(twiddle_factor_table_100_real));
  assign _zz_5304 = ($signed(_zz_15490) * $signed(twiddle_factor_table_100_imag));
  assign _zz_3898 = ($signed(_zz_3900) - $signed(_zz_15491));
  assign _zz_3899 = ($signed(_zz_3900) + $signed(_zz_15493));
  assign _zz_3901 = 1'b1;
  assign _zz_3902 = 1'b1;
  assign _zz_5305 = ($signed(_zz_15511) * $signed(_zz_1741));
  assign _zz_3905 = _zz_15512[15 : 0];
  assign _zz_5306 = ($signed(_zz_15513) * $signed(twiddle_factor_table_101_real));
  assign _zz_5307 = ($signed(_zz_15514) * $signed(twiddle_factor_table_101_imag));
  assign _zz_3903 = ($signed(_zz_3905) - $signed(_zz_15515));
  assign _zz_3904 = ($signed(_zz_3905) + $signed(_zz_15517));
  assign _zz_3906 = 1'b1;
  assign _zz_3907 = 1'b1;
  assign _zz_5308 = ($signed(_zz_15535) * $signed(_zz_1743));
  assign _zz_3910 = _zz_15536[15 : 0];
  assign _zz_5309 = ($signed(_zz_15537) * $signed(twiddle_factor_table_102_real));
  assign _zz_5310 = ($signed(_zz_15538) * $signed(twiddle_factor_table_102_imag));
  assign _zz_3908 = ($signed(_zz_3910) - $signed(_zz_15539));
  assign _zz_3909 = ($signed(_zz_3910) + $signed(_zz_15541));
  assign _zz_3911 = 1'b1;
  assign _zz_3912 = 1'b1;
  assign _zz_5311 = ($signed(_zz_15559) * $signed(_zz_1745));
  assign _zz_3915 = _zz_15560[15 : 0];
  assign _zz_5312 = ($signed(_zz_15561) * $signed(twiddle_factor_table_103_real));
  assign _zz_5313 = ($signed(_zz_15562) * $signed(twiddle_factor_table_103_imag));
  assign _zz_3913 = ($signed(_zz_3915) - $signed(_zz_15563));
  assign _zz_3914 = ($signed(_zz_3915) + $signed(_zz_15565));
  assign _zz_3916 = 1'b1;
  assign _zz_3917 = 1'b1;
  assign _zz_5314 = ($signed(_zz_15583) * $signed(_zz_1747));
  assign _zz_3920 = _zz_15584[15 : 0];
  assign _zz_5315 = ($signed(_zz_15585) * $signed(twiddle_factor_table_104_real));
  assign _zz_5316 = ($signed(_zz_15586) * $signed(twiddle_factor_table_104_imag));
  assign _zz_3918 = ($signed(_zz_3920) - $signed(_zz_15587));
  assign _zz_3919 = ($signed(_zz_3920) + $signed(_zz_15589));
  assign _zz_3921 = 1'b1;
  assign _zz_3922 = 1'b1;
  assign _zz_5317 = ($signed(_zz_15607) * $signed(_zz_1749));
  assign _zz_3925 = _zz_15608[15 : 0];
  assign _zz_5318 = ($signed(_zz_15609) * $signed(twiddle_factor_table_105_real));
  assign _zz_5319 = ($signed(_zz_15610) * $signed(twiddle_factor_table_105_imag));
  assign _zz_3923 = ($signed(_zz_3925) - $signed(_zz_15611));
  assign _zz_3924 = ($signed(_zz_3925) + $signed(_zz_15613));
  assign _zz_3926 = 1'b1;
  assign _zz_3927 = 1'b1;
  assign _zz_5320 = ($signed(_zz_15631) * $signed(_zz_1751));
  assign _zz_3930 = _zz_15632[15 : 0];
  assign _zz_5321 = ($signed(_zz_15633) * $signed(twiddle_factor_table_106_real));
  assign _zz_5322 = ($signed(_zz_15634) * $signed(twiddle_factor_table_106_imag));
  assign _zz_3928 = ($signed(_zz_3930) - $signed(_zz_15635));
  assign _zz_3929 = ($signed(_zz_3930) + $signed(_zz_15637));
  assign _zz_3931 = 1'b1;
  assign _zz_3932 = 1'b1;
  assign _zz_5323 = ($signed(_zz_15655) * $signed(_zz_1753));
  assign _zz_3935 = _zz_15656[15 : 0];
  assign _zz_5324 = ($signed(_zz_15657) * $signed(twiddle_factor_table_107_real));
  assign _zz_5325 = ($signed(_zz_15658) * $signed(twiddle_factor_table_107_imag));
  assign _zz_3933 = ($signed(_zz_3935) - $signed(_zz_15659));
  assign _zz_3934 = ($signed(_zz_3935) + $signed(_zz_15661));
  assign _zz_3936 = 1'b1;
  assign _zz_3937 = 1'b1;
  assign _zz_5326 = ($signed(_zz_15679) * $signed(_zz_1755));
  assign _zz_3940 = _zz_15680[15 : 0];
  assign _zz_5327 = ($signed(_zz_15681) * $signed(twiddle_factor_table_108_real));
  assign _zz_5328 = ($signed(_zz_15682) * $signed(twiddle_factor_table_108_imag));
  assign _zz_3938 = ($signed(_zz_3940) - $signed(_zz_15683));
  assign _zz_3939 = ($signed(_zz_3940) + $signed(_zz_15685));
  assign _zz_3941 = 1'b1;
  assign _zz_3942 = 1'b1;
  assign _zz_5329 = ($signed(_zz_15703) * $signed(_zz_1757));
  assign _zz_3945 = _zz_15704[15 : 0];
  assign _zz_5330 = ($signed(_zz_15705) * $signed(twiddle_factor_table_109_real));
  assign _zz_5331 = ($signed(_zz_15706) * $signed(twiddle_factor_table_109_imag));
  assign _zz_3943 = ($signed(_zz_3945) - $signed(_zz_15707));
  assign _zz_3944 = ($signed(_zz_3945) + $signed(_zz_15709));
  assign _zz_3946 = 1'b1;
  assign _zz_3947 = 1'b1;
  assign _zz_5332 = ($signed(_zz_15727) * $signed(_zz_1759));
  assign _zz_3950 = _zz_15728[15 : 0];
  assign _zz_5333 = ($signed(_zz_15729) * $signed(twiddle_factor_table_110_real));
  assign _zz_5334 = ($signed(_zz_15730) * $signed(twiddle_factor_table_110_imag));
  assign _zz_3948 = ($signed(_zz_3950) - $signed(_zz_15731));
  assign _zz_3949 = ($signed(_zz_3950) + $signed(_zz_15733));
  assign _zz_3951 = 1'b1;
  assign _zz_3952 = 1'b1;
  assign _zz_5335 = ($signed(_zz_15751) * $signed(_zz_1761));
  assign _zz_3955 = _zz_15752[15 : 0];
  assign _zz_5336 = ($signed(_zz_15753) * $signed(twiddle_factor_table_111_real));
  assign _zz_5337 = ($signed(_zz_15754) * $signed(twiddle_factor_table_111_imag));
  assign _zz_3953 = ($signed(_zz_3955) - $signed(_zz_15755));
  assign _zz_3954 = ($signed(_zz_3955) + $signed(_zz_15757));
  assign _zz_3956 = 1'b1;
  assign _zz_3957 = 1'b1;
  assign _zz_5338 = ($signed(_zz_15775) * $signed(_zz_1763));
  assign _zz_3960 = _zz_15776[15 : 0];
  assign _zz_5339 = ($signed(_zz_15777) * $signed(twiddle_factor_table_112_real));
  assign _zz_5340 = ($signed(_zz_15778) * $signed(twiddle_factor_table_112_imag));
  assign _zz_3958 = ($signed(_zz_3960) - $signed(_zz_15779));
  assign _zz_3959 = ($signed(_zz_3960) + $signed(_zz_15781));
  assign _zz_3961 = 1'b1;
  assign _zz_3962 = 1'b1;
  assign _zz_5341 = ($signed(_zz_15799) * $signed(_zz_1765));
  assign _zz_3965 = _zz_15800[15 : 0];
  assign _zz_5342 = ($signed(_zz_15801) * $signed(twiddle_factor_table_113_real));
  assign _zz_5343 = ($signed(_zz_15802) * $signed(twiddle_factor_table_113_imag));
  assign _zz_3963 = ($signed(_zz_3965) - $signed(_zz_15803));
  assign _zz_3964 = ($signed(_zz_3965) + $signed(_zz_15805));
  assign _zz_3966 = 1'b1;
  assign _zz_3967 = 1'b1;
  assign _zz_5344 = ($signed(_zz_15823) * $signed(_zz_1767));
  assign _zz_3970 = _zz_15824[15 : 0];
  assign _zz_5345 = ($signed(_zz_15825) * $signed(twiddle_factor_table_114_real));
  assign _zz_5346 = ($signed(_zz_15826) * $signed(twiddle_factor_table_114_imag));
  assign _zz_3968 = ($signed(_zz_3970) - $signed(_zz_15827));
  assign _zz_3969 = ($signed(_zz_3970) + $signed(_zz_15829));
  assign _zz_3971 = 1'b1;
  assign _zz_3972 = 1'b1;
  assign _zz_5347 = ($signed(_zz_15847) * $signed(_zz_1769));
  assign _zz_3975 = _zz_15848[15 : 0];
  assign _zz_5348 = ($signed(_zz_15849) * $signed(twiddle_factor_table_115_real));
  assign _zz_5349 = ($signed(_zz_15850) * $signed(twiddle_factor_table_115_imag));
  assign _zz_3973 = ($signed(_zz_3975) - $signed(_zz_15851));
  assign _zz_3974 = ($signed(_zz_3975) + $signed(_zz_15853));
  assign _zz_3976 = 1'b1;
  assign _zz_3977 = 1'b1;
  assign _zz_5350 = ($signed(_zz_15871) * $signed(_zz_1771));
  assign _zz_3980 = _zz_15872[15 : 0];
  assign _zz_5351 = ($signed(_zz_15873) * $signed(twiddle_factor_table_116_real));
  assign _zz_5352 = ($signed(_zz_15874) * $signed(twiddle_factor_table_116_imag));
  assign _zz_3978 = ($signed(_zz_3980) - $signed(_zz_15875));
  assign _zz_3979 = ($signed(_zz_3980) + $signed(_zz_15877));
  assign _zz_3981 = 1'b1;
  assign _zz_3982 = 1'b1;
  assign _zz_5353 = ($signed(_zz_15895) * $signed(_zz_1773));
  assign _zz_3985 = _zz_15896[15 : 0];
  assign _zz_5354 = ($signed(_zz_15897) * $signed(twiddle_factor_table_117_real));
  assign _zz_5355 = ($signed(_zz_15898) * $signed(twiddle_factor_table_117_imag));
  assign _zz_3983 = ($signed(_zz_3985) - $signed(_zz_15899));
  assign _zz_3984 = ($signed(_zz_3985) + $signed(_zz_15901));
  assign _zz_3986 = 1'b1;
  assign _zz_3987 = 1'b1;
  assign _zz_5356 = ($signed(_zz_15919) * $signed(_zz_1775));
  assign _zz_3990 = _zz_15920[15 : 0];
  assign _zz_5357 = ($signed(_zz_15921) * $signed(twiddle_factor_table_118_real));
  assign _zz_5358 = ($signed(_zz_15922) * $signed(twiddle_factor_table_118_imag));
  assign _zz_3988 = ($signed(_zz_3990) - $signed(_zz_15923));
  assign _zz_3989 = ($signed(_zz_3990) + $signed(_zz_15925));
  assign _zz_3991 = 1'b1;
  assign _zz_3992 = 1'b1;
  assign _zz_5359 = ($signed(_zz_15943) * $signed(_zz_1777));
  assign _zz_3995 = _zz_15944[15 : 0];
  assign _zz_5360 = ($signed(_zz_15945) * $signed(twiddle_factor_table_119_real));
  assign _zz_5361 = ($signed(_zz_15946) * $signed(twiddle_factor_table_119_imag));
  assign _zz_3993 = ($signed(_zz_3995) - $signed(_zz_15947));
  assign _zz_3994 = ($signed(_zz_3995) + $signed(_zz_15949));
  assign _zz_3996 = 1'b1;
  assign _zz_3997 = 1'b1;
  assign _zz_5362 = ($signed(_zz_15967) * $signed(_zz_1779));
  assign _zz_4000 = _zz_15968[15 : 0];
  assign _zz_5363 = ($signed(_zz_15969) * $signed(twiddle_factor_table_120_real));
  assign _zz_5364 = ($signed(_zz_15970) * $signed(twiddle_factor_table_120_imag));
  assign _zz_3998 = ($signed(_zz_4000) - $signed(_zz_15971));
  assign _zz_3999 = ($signed(_zz_4000) + $signed(_zz_15973));
  assign _zz_4001 = 1'b1;
  assign _zz_4002 = 1'b1;
  assign _zz_5365 = ($signed(_zz_15991) * $signed(_zz_1781));
  assign _zz_4005 = _zz_15992[15 : 0];
  assign _zz_5366 = ($signed(_zz_15993) * $signed(twiddle_factor_table_121_real));
  assign _zz_5367 = ($signed(_zz_15994) * $signed(twiddle_factor_table_121_imag));
  assign _zz_4003 = ($signed(_zz_4005) - $signed(_zz_15995));
  assign _zz_4004 = ($signed(_zz_4005) + $signed(_zz_15997));
  assign _zz_4006 = 1'b1;
  assign _zz_4007 = 1'b1;
  assign _zz_5368 = ($signed(_zz_16015) * $signed(_zz_1783));
  assign _zz_4010 = _zz_16016[15 : 0];
  assign _zz_5369 = ($signed(_zz_16017) * $signed(twiddle_factor_table_122_real));
  assign _zz_5370 = ($signed(_zz_16018) * $signed(twiddle_factor_table_122_imag));
  assign _zz_4008 = ($signed(_zz_4010) - $signed(_zz_16019));
  assign _zz_4009 = ($signed(_zz_4010) + $signed(_zz_16021));
  assign _zz_4011 = 1'b1;
  assign _zz_4012 = 1'b1;
  assign _zz_5371 = ($signed(_zz_16039) * $signed(_zz_1785));
  assign _zz_4015 = _zz_16040[15 : 0];
  assign _zz_5372 = ($signed(_zz_16041) * $signed(twiddle_factor_table_123_real));
  assign _zz_5373 = ($signed(_zz_16042) * $signed(twiddle_factor_table_123_imag));
  assign _zz_4013 = ($signed(_zz_4015) - $signed(_zz_16043));
  assign _zz_4014 = ($signed(_zz_4015) + $signed(_zz_16045));
  assign _zz_4016 = 1'b1;
  assign _zz_4017 = 1'b1;
  assign _zz_5374 = ($signed(_zz_16063) * $signed(_zz_1787));
  assign _zz_4020 = _zz_16064[15 : 0];
  assign _zz_5375 = ($signed(_zz_16065) * $signed(twiddle_factor_table_124_real));
  assign _zz_5376 = ($signed(_zz_16066) * $signed(twiddle_factor_table_124_imag));
  assign _zz_4018 = ($signed(_zz_4020) - $signed(_zz_16067));
  assign _zz_4019 = ($signed(_zz_4020) + $signed(_zz_16069));
  assign _zz_4021 = 1'b1;
  assign _zz_4022 = 1'b1;
  assign _zz_5377 = ($signed(_zz_16087) * $signed(_zz_1789));
  assign _zz_4025 = _zz_16088[15 : 0];
  assign _zz_5378 = ($signed(_zz_16089) * $signed(twiddle_factor_table_125_real));
  assign _zz_5379 = ($signed(_zz_16090) * $signed(twiddle_factor_table_125_imag));
  assign _zz_4023 = ($signed(_zz_4025) - $signed(_zz_16091));
  assign _zz_4024 = ($signed(_zz_4025) + $signed(_zz_16093));
  assign _zz_4026 = 1'b1;
  assign _zz_4027 = 1'b1;
  assign _zz_5380 = ($signed(_zz_16111) * $signed(_zz_1791));
  assign _zz_4030 = _zz_16112[15 : 0];
  assign _zz_5381 = ($signed(_zz_16113) * $signed(twiddle_factor_table_126_real));
  assign _zz_5382 = ($signed(_zz_16114) * $signed(twiddle_factor_table_126_imag));
  assign _zz_4028 = ($signed(_zz_4030) - $signed(_zz_16115));
  assign _zz_4029 = ($signed(_zz_4030) + $signed(_zz_16117));
  assign _zz_4031 = 1'b1;
  assign _zz_4032 = 1'b1;
  always @ (*) begin
    _zz_4033 = 1'b0;
    if((io_data_in_valid_regNext || _zz_4038))begin
      _zz_4033 = 1'b1;
    end
  end

  assign _zz_4036 = (_zz_4035 == 4'b1000);
  assign _zz_4037 = (_zz_4036 && _zz_4033);
  always @ (*) begin
    if(_zz_4037)begin
      _zz_4034 = 4'b0000;
    end else begin
      _zz_4034 = (_zz_4035 + _zz_16136);
    end
    if(1'b0)begin
      _zz_4034 = 4'b0000;
    end
  end

  assign io_data_out_valid = _zz_4037;
  assign io_data_out_payload_0_real = _zz_1537;
  assign io_data_out_payload_0_imag = _zz_1538;
  assign io_data_out_payload_1_real = _zz_1539;
  assign io_data_out_payload_1_imag = _zz_1540;
  assign io_data_out_payload_2_real = _zz_1541;
  assign io_data_out_payload_2_imag = _zz_1542;
  assign io_data_out_payload_3_real = _zz_1543;
  assign io_data_out_payload_3_imag = _zz_1544;
  assign io_data_out_payload_4_real = _zz_1545;
  assign io_data_out_payload_4_imag = _zz_1546;
  assign io_data_out_payload_5_real = _zz_1547;
  assign io_data_out_payload_5_imag = _zz_1548;
  assign io_data_out_payload_6_real = _zz_1549;
  assign io_data_out_payload_6_imag = _zz_1550;
  assign io_data_out_payload_7_real = _zz_1551;
  assign io_data_out_payload_7_imag = _zz_1552;
  assign io_data_out_payload_8_real = _zz_1553;
  assign io_data_out_payload_8_imag = _zz_1554;
  assign io_data_out_payload_9_real = _zz_1555;
  assign io_data_out_payload_9_imag = _zz_1556;
  assign io_data_out_payload_10_real = _zz_1557;
  assign io_data_out_payload_10_imag = _zz_1558;
  assign io_data_out_payload_11_real = _zz_1559;
  assign io_data_out_payload_11_imag = _zz_1560;
  assign io_data_out_payload_12_real = _zz_1561;
  assign io_data_out_payload_12_imag = _zz_1562;
  assign io_data_out_payload_13_real = _zz_1563;
  assign io_data_out_payload_13_imag = _zz_1564;
  assign io_data_out_payload_14_real = _zz_1565;
  assign io_data_out_payload_14_imag = _zz_1566;
  assign io_data_out_payload_15_real = _zz_1567;
  assign io_data_out_payload_15_imag = _zz_1568;
  assign io_data_out_payload_16_real = _zz_1569;
  assign io_data_out_payload_16_imag = _zz_1570;
  assign io_data_out_payload_17_real = _zz_1571;
  assign io_data_out_payload_17_imag = _zz_1572;
  assign io_data_out_payload_18_real = _zz_1573;
  assign io_data_out_payload_18_imag = _zz_1574;
  assign io_data_out_payload_19_real = _zz_1575;
  assign io_data_out_payload_19_imag = _zz_1576;
  assign io_data_out_payload_20_real = _zz_1577;
  assign io_data_out_payload_20_imag = _zz_1578;
  assign io_data_out_payload_21_real = _zz_1579;
  assign io_data_out_payload_21_imag = _zz_1580;
  assign io_data_out_payload_22_real = _zz_1581;
  assign io_data_out_payload_22_imag = _zz_1582;
  assign io_data_out_payload_23_real = _zz_1583;
  assign io_data_out_payload_23_imag = _zz_1584;
  assign io_data_out_payload_24_real = _zz_1585;
  assign io_data_out_payload_24_imag = _zz_1586;
  assign io_data_out_payload_25_real = _zz_1587;
  assign io_data_out_payload_25_imag = _zz_1588;
  assign io_data_out_payload_26_real = _zz_1589;
  assign io_data_out_payload_26_imag = _zz_1590;
  assign io_data_out_payload_27_real = _zz_1591;
  assign io_data_out_payload_27_imag = _zz_1592;
  assign io_data_out_payload_28_real = _zz_1593;
  assign io_data_out_payload_28_imag = _zz_1594;
  assign io_data_out_payload_29_real = _zz_1595;
  assign io_data_out_payload_29_imag = _zz_1596;
  assign io_data_out_payload_30_real = _zz_1597;
  assign io_data_out_payload_30_imag = _zz_1598;
  assign io_data_out_payload_31_real = _zz_1599;
  assign io_data_out_payload_31_imag = _zz_1600;
  assign io_data_out_payload_32_real = _zz_1601;
  assign io_data_out_payload_32_imag = _zz_1602;
  assign io_data_out_payload_33_real = _zz_1603;
  assign io_data_out_payload_33_imag = _zz_1604;
  assign io_data_out_payload_34_real = _zz_1605;
  assign io_data_out_payload_34_imag = _zz_1606;
  assign io_data_out_payload_35_real = _zz_1607;
  assign io_data_out_payload_35_imag = _zz_1608;
  assign io_data_out_payload_36_real = _zz_1609;
  assign io_data_out_payload_36_imag = _zz_1610;
  assign io_data_out_payload_37_real = _zz_1611;
  assign io_data_out_payload_37_imag = _zz_1612;
  assign io_data_out_payload_38_real = _zz_1613;
  assign io_data_out_payload_38_imag = _zz_1614;
  assign io_data_out_payload_39_real = _zz_1615;
  assign io_data_out_payload_39_imag = _zz_1616;
  assign io_data_out_payload_40_real = _zz_1617;
  assign io_data_out_payload_40_imag = _zz_1618;
  assign io_data_out_payload_41_real = _zz_1619;
  assign io_data_out_payload_41_imag = _zz_1620;
  assign io_data_out_payload_42_real = _zz_1621;
  assign io_data_out_payload_42_imag = _zz_1622;
  assign io_data_out_payload_43_real = _zz_1623;
  assign io_data_out_payload_43_imag = _zz_1624;
  assign io_data_out_payload_44_real = _zz_1625;
  assign io_data_out_payload_44_imag = _zz_1626;
  assign io_data_out_payload_45_real = _zz_1627;
  assign io_data_out_payload_45_imag = _zz_1628;
  assign io_data_out_payload_46_real = _zz_1629;
  assign io_data_out_payload_46_imag = _zz_1630;
  assign io_data_out_payload_47_real = _zz_1631;
  assign io_data_out_payload_47_imag = _zz_1632;
  assign io_data_out_payload_48_real = _zz_1633;
  assign io_data_out_payload_48_imag = _zz_1634;
  assign io_data_out_payload_49_real = _zz_1635;
  assign io_data_out_payload_49_imag = _zz_1636;
  assign io_data_out_payload_50_real = _zz_1637;
  assign io_data_out_payload_50_imag = _zz_1638;
  assign io_data_out_payload_51_real = _zz_1639;
  assign io_data_out_payload_51_imag = _zz_1640;
  assign io_data_out_payload_52_real = _zz_1641;
  assign io_data_out_payload_52_imag = _zz_1642;
  assign io_data_out_payload_53_real = _zz_1643;
  assign io_data_out_payload_53_imag = _zz_1644;
  assign io_data_out_payload_54_real = _zz_1645;
  assign io_data_out_payload_54_imag = _zz_1646;
  assign io_data_out_payload_55_real = _zz_1647;
  assign io_data_out_payload_55_imag = _zz_1648;
  assign io_data_out_payload_56_real = _zz_1649;
  assign io_data_out_payload_56_imag = _zz_1650;
  assign io_data_out_payload_57_real = _zz_1651;
  assign io_data_out_payload_57_imag = _zz_1652;
  assign io_data_out_payload_58_real = _zz_1653;
  assign io_data_out_payload_58_imag = _zz_1654;
  assign io_data_out_payload_59_real = _zz_1655;
  assign io_data_out_payload_59_imag = _zz_1656;
  assign io_data_out_payload_60_real = _zz_1657;
  assign io_data_out_payload_60_imag = _zz_1658;
  assign io_data_out_payload_61_real = _zz_1659;
  assign io_data_out_payload_61_imag = _zz_1660;
  assign io_data_out_payload_62_real = _zz_1661;
  assign io_data_out_payload_62_imag = _zz_1662;
  assign io_data_out_payload_63_real = _zz_1663;
  assign io_data_out_payload_63_imag = _zz_1664;
  assign io_data_out_payload_64_real = _zz_1665;
  assign io_data_out_payload_64_imag = _zz_1666;
  assign io_data_out_payload_65_real = _zz_1667;
  assign io_data_out_payload_65_imag = _zz_1668;
  assign io_data_out_payload_66_real = _zz_1669;
  assign io_data_out_payload_66_imag = _zz_1670;
  assign io_data_out_payload_67_real = _zz_1671;
  assign io_data_out_payload_67_imag = _zz_1672;
  assign io_data_out_payload_68_real = _zz_1673;
  assign io_data_out_payload_68_imag = _zz_1674;
  assign io_data_out_payload_69_real = _zz_1675;
  assign io_data_out_payload_69_imag = _zz_1676;
  assign io_data_out_payload_70_real = _zz_1677;
  assign io_data_out_payload_70_imag = _zz_1678;
  assign io_data_out_payload_71_real = _zz_1679;
  assign io_data_out_payload_71_imag = _zz_1680;
  assign io_data_out_payload_72_real = _zz_1681;
  assign io_data_out_payload_72_imag = _zz_1682;
  assign io_data_out_payload_73_real = _zz_1683;
  assign io_data_out_payload_73_imag = _zz_1684;
  assign io_data_out_payload_74_real = _zz_1685;
  assign io_data_out_payload_74_imag = _zz_1686;
  assign io_data_out_payload_75_real = _zz_1687;
  assign io_data_out_payload_75_imag = _zz_1688;
  assign io_data_out_payload_76_real = _zz_1689;
  assign io_data_out_payload_76_imag = _zz_1690;
  assign io_data_out_payload_77_real = _zz_1691;
  assign io_data_out_payload_77_imag = _zz_1692;
  assign io_data_out_payload_78_real = _zz_1693;
  assign io_data_out_payload_78_imag = _zz_1694;
  assign io_data_out_payload_79_real = _zz_1695;
  assign io_data_out_payload_79_imag = _zz_1696;
  assign io_data_out_payload_80_real = _zz_1697;
  assign io_data_out_payload_80_imag = _zz_1698;
  assign io_data_out_payload_81_real = _zz_1699;
  assign io_data_out_payload_81_imag = _zz_1700;
  assign io_data_out_payload_82_real = _zz_1701;
  assign io_data_out_payload_82_imag = _zz_1702;
  assign io_data_out_payload_83_real = _zz_1703;
  assign io_data_out_payload_83_imag = _zz_1704;
  assign io_data_out_payload_84_real = _zz_1705;
  assign io_data_out_payload_84_imag = _zz_1706;
  assign io_data_out_payload_85_real = _zz_1707;
  assign io_data_out_payload_85_imag = _zz_1708;
  assign io_data_out_payload_86_real = _zz_1709;
  assign io_data_out_payload_86_imag = _zz_1710;
  assign io_data_out_payload_87_real = _zz_1711;
  assign io_data_out_payload_87_imag = _zz_1712;
  assign io_data_out_payload_88_real = _zz_1713;
  assign io_data_out_payload_88_imag = _zz_1714;
  assign io_data_out_payload_89_real = _zz_1715;
  assign io_data_out_payload_89_imag = _zz_1716;
  assign io_data_out_payload_90_real = _zz_1717;
  assign io_data_out_payload_90_imag = _zz_1718;
  assign io_data_out_payload_91_real = _zz_1719;
  assign io_data_out_payload_91_imag = _zz_1720;
  assign io_data_out_payload_92_real = _zz_1721;
  assign io_data_out_payload_92_imag = _zz_1722;
  assign io_data_out_payload_93_real = _zz_1723;
  assign io_data_out_payload_93_imag = _zz_1724;
  assign io_data_out_payload_94_real = _zz_1725;
  assign io_data_out_payload_94_imag = _zz_1726;
  assign io_data_out_payload_95_real = _zz_1727;
  assign io_data_out_payload_95_imag = _zz_1728;
  assign io_data_out_payload_96_real = _zz_1729;
  assign io_data_out_payload_96_imag = _zz_1730;
  assign io_data_out_payload_97_real = _zz_1731;
  assign io_data_out_payload_97_imag = _zz_1732;
  assign io_data_out_payload_98_real = _zz_1733;
  assign io_data_out_payload_98_imag = _zz_1734;
  assign io_data_out_payload_99_real = _zz_1735;
  assign io_data_out_payload_99_imag = _zz_1736;
  assign io_data_out_payload_100_real = _zz_1737;
  assign io_data_out_payload_100_imag = _zz_1738;
  assign io_data_out_payload_101_real = _zz_1739;
  assign io_data_out_payload_101_imag = _zz_1740;
  assign io_data_out_payload_102_real = _zz_1741;
  assign io_data_out_payload_102_imag = _zz_1742;
  assign io_data_out_payload_103_real = _zz_1743;
  assign io_data_out_payload_103_imag = _zz_1744;
  assign io_data_out_payload_104_real = _zz_1745;
  assign io_data_out_payload_104_imag = _zz_1746;
  assign io_data_out_payload_105_real = _zz_1747;
  assign io_data_out_payload_105_imag = _zz_1748;
  assign io_data_out_payload_106_real = _zz_1749;
  assign io_data_out_payload_106_imag = _zz_1750;
  assign io_data_out_payload_107_real = _zz_1751;
  assign io_data_out_payload_107_imag = _zz_1752;
  assign io_data_out_payload_108_real = _zz_1753;
  assign io_data_out_payload_108_imag = _zz_1754;
  assign io_data_out_payload_109_real = _zz_1755;
  assign io_data_out_payload_109_imag = _zz_1756;
  assign io_data_out_payload_110_real = _zz_1757;
  assign io_data_out_payload_110_imag = _zz_1758;
  assign io_data_out_payload_111_real = _zz_1759;
  assign io_data_out_payload_111_imag = _zz_1760;
  assign io_data_out_payload_112_real = _zz_1761;
  assign io_data_out_payload_112_imag = _zz_1762;
  assign io_data_out_payload_113_real = _zz_1763;
  assign io_data_out_payload_113_imag = _zz_1764;
  assign io_data_out_payload_114_real = _zz_1765;
  assign io_data_out_payload_114_imag = _zz_1766;
  assign io_data_out_payload_115_real = _zz_1767;
  assign io_data_out_payload_115_imag = _zz_1768;
  assign io_data_out_payload_116_real = _zz_1769;
  assign io_data_out_payload_116_imag = _zz_1770;
  assign io_data_out_payload_117_real = _zz_1771;
  assign io_data_out_payload_117_imag = _zz_1772;
  assign io_data_out_payload_118_real = _zz_1773;
  assign io_data_out_payload_118_imag = _zz_1774;
  assign io_data_out_payload_119_real = _zz_1775;
  assign io_data_out_payload_119_imag = _zz_1776;
  assign io_data_out_payload_120_real = _zz_1777;
  assign io_data_out_payload_120_imag = _zz_1778;
  assign io_data_out_payload_121_real = _zz_1779;
  assign io_data_out_payload_121_imag = _zz_1780;
  assign io_data_out_payload_122_real = _zz_1781;
  assign io_data_out_payload_122_imag = _zz_1782;
  assign io_data_out_payload_123_real = _zz_1783;
  assign io_data_out_payload_123_imag = _zz_1784;
  assign io_data_out_payload_124_real = _zz_1785;
  assign io_data_out_payload_124_imag = _zz_1786;
  assign io_data_out_payload_125_real = _zz_1787;
  assign io_data_out_payload_125_imag = _zz_1788;
  assign io_data_out_payload_126_real = _zz_1789;
  assign io_data_out_payload_126_imag = _zz_1790;
  assign io_data_out_payload_127_real = _zz_1791;
  assign io_data_out_payload_127_imag = _zz_1792;
  always @ (posedge clk) begin
    if(io_data_in_valid)begin
      data_in_0_real <= io_data_in_payload_0_real;
      data_in_0_imag <= io_data_in_payload_0_imag;
      data_in_1_real <= io_data_in_payload_1_real;
      data_in_1_imag <= io_data_in_payload_1_imag;
      data_in_2_real <= io_data_in_payload_2_real;
      data_in_2_imag <= io_data_in_payload_2_imag;
      data_in_3_real <= io_data_in_payload_3_real;
      data_in_3_imag <= io_data_in_payload_3_imag;
      data_in_4_real <= io_data_in_payload_4_real;
      data_in_4_imag <= io_data_in_payload_4_imag;
      data_in_5_real <= io_data_in_payload_5_real;
      data_in_5_imag <= io_data_in_payload_5_imag;
      data_in_6_real <= io_data_in_payload_6_real;
      data_in_6_imag <= io_data_in_payload_6_imag;
      data_in_7_real <= io_data_in_payload_7_real;
      data_in_7_imag <= io_data_in_payload_7_imag;
      data_in_8_real <= io_data_in_payload_8_real;
      data_in_8_imag <= io_data_in_payload_8_imag;
      data_in_9_real <= io_data_in_payload_9_real;
      data_in_9_imag <= io_data_in_payload_9_imag;
      data_in_10_real <= io_data_in_payload_10_real;
      data_in_10_imag <= io_data_in_payload_10_imag;
      data_in_11_real <= io_data_in_payload_11_real;
      data_in_11_imag <= io_data_in_payload_11_imag;
      data_in_12_real <= io_data_in_payload_12_real;
      data_in_12_imag <= io_data_in_payload_12_imag;
      data_in_13_real <= io_data_in_payload_13_real;
      data_in_13_imag <= io_data_in_payload_13_imag;
      data_in_14_real <= io_data_in_payload_14_real;
      data_in_14_imag <= io_data_in_payload_14_imag;
      data_in_15_real <= io_data_in_payload_15_real;
      data_in_15_imag <= io_data_in_payload_15_imag;
      data_in_16_real <= io_data_in_payload_16_real;
      data_in_16_imag <= io_data_in_payload_16_imag;
      data_in_17_real <= io_data_in_payload_17_real;
      data_in_17_imag <= io_data_in_payload_17_imag;
      data_in_18_real <= io_data_in_payload_18_real;
      data_in_18_imag <= io_data_in_payload_18_imag;
      data_in_19_real <= io_data_in_payload_19_real;
      data_in_19_imag <= io_data_in_payload_19_imag;
      data_in_20_real <= io_data_in_payload_20_real;
      data_in_20_imag <= io_data_in_payload_20_imag;
      data_in_21_real <= io_data_in_payload_21_real;
      data_in_21_imag <= io_data_in_payload_21_imag;
      data_in_22_real <= io_data_in_payload_22_real;
      data_in_22_imag <= io_data_in_payload_22_imag;
      data_in_23_real <= io_data_in_payload_23_real;
      data_in_23_imag <= io_data_in_payload_23_imag;
      data_in_24_real <= io_data_in_payload_24_real;
      data_in_24_imag <= io_data_in_payload_24_imag;
      data_in_25_real <= io_data_in_payload_25_real;
      data_in_25_imag <= io_data_in_payload_25_imag;
      data_in_26_real <= io_data_in_payload_26_real;
      data_in_26_imag <= io_data_in_payload_26_imag;
      data_in_27_real <= io_data_in_payload_27_real;
      data_in_27_imag <= io_data_in_payload_27_imag;
      data_in_28_real <= io_data_in_payload_28_real;
      data_in_28_imag <= io_data_in_payload_28_imag;
      data_in_29_real <= io_data_in_payload_29_real;
      data_in_29_imag <= io_data_in_payload_29_imag;
      data_in_30_real <= io_data_in_payload_30_real;
      data_in_30_imag <= io_data_in_payload_30_imag;
      data_in_31_real <= io_data_in_payload_31_real;
      data_in_31_imag <= io_data_in_payload_31_imag;
      data_in_32_real <= io_data_in_payload_32_real;
      data_in_32_imag <= io_data_in_payload_32_imag;
      data_in_33_real <= io_data_in_payload_33_real;
      data_in_33_imag <= io_data_in_payload_33_imag;
      data_in_34_real <= io_data_in_payload_34_real;
      data_in_34_imag <= io_data_in_payload_34_imag;
      data_in_35_real <= io_data_in_payload_35_real;
      data_in_35_imag <= io_data_in_payload_35_imag;
      data_in_36_real <= io_data_in_payload_36_real;
      data_in_36_imag <= io_data_in_payload_36_imag;
      data_in_37_real <= io_data_in_payload_37_real;
      data_in_37_imag <= io_data_in_payload_37_imag;
      data_in_38_real <= io_data_in_payload_38_real;
      data_in_38_imag <= io_data_in_payload_38_imag;
      data_in_39_real <= io_data_in_payload_39_real;
      data_in_39_imag <= io_data_in_payload_39_imag;
      data_in_40_real <= io_data_in_payload_40_real;
      data_in_40_imag <= io_data_in_payload_40_imag;
      data_in_41_real <= io_data_in_payload_41_real;
      data_in_41_imag <= io_data_in_payload_41_imag;
      data_in_42_real <= io_data_in_payload_42_real;
      data_in_42_imag <= io_data_in_payload_42_imag;
      data_in_43_real <= io_data_in_payload_43_real;
      data_in_43_imag <= io_data_in_payload_43_imag;
      data_in_44_real <= io_data_in_payload_44_real;
      data_in_44_imag <= io_data_in_payload_44_imag;
      data_in_45_real <= io_data_in_payload_45_real;
      data_in_45_imag <= io_data_in_payload_45_imag;
      data_in_46_real <= io_data_in_payload_46_real;
      data_in_46_imag <= io_data_in_payload_46_imag;
      data_in_47_real <= io_data_in_payload_47_real;
      data_in_47_imag <= io_data_in_payload_47_imag;
      data_in_48_real <= io_data_in_payload_48_real;
      data_in_48_imag <= io_data_in_payload_48_imag;
      data_in_49_real <= io_data_in_payload_49_real;
      data_in_49_imag <= io_data_in_payload_49_imag;
      data_in_50_real <= io_data_in_payload_50_real;
      data_in_50_imag <= io_data_in_payload_50_imag;
      data_in_51_real <= io_data_in_payload_51_real;
      data_in_51_imag <= io_data_in_payload_51_imag;
      data_in_52_real <= io_data_in_payload_52_real;
      data_in_52_imag <= io_data_in_payload_52_imag;
      data_in_53_real <= io_data_in_payload_53_real;
      data_in_53_imag <= io_data_in_payload_53_imag;
      data_in_54_real <= io_data_in_payload_54_real;
      data_in_54_imag <= io_data_in_payload_54_imag;
      data_in_55_real <= io_data_in_payload_55_real;
      data_in_55_imag <= io_data_in_payload_55_imag;
      data_in_56_real <= io_data_in_payload_56_real;
      data_in_56_imag <= io_data_in_payload_56_imag;
      data_in_57_real <= io_data_in_payload_57_real;
      data_in_57_imag <= io_data_in_payload_57_imag;
      data_in_58_real <= io_data_in_payload_58_real;
      data_in_58_imag <= io_data_in_payload_58_imag;
      data_in_59_real <= io_data_in_payload_59_real;
      data_in_59_imag <= io_data_in_payload_59_imag;
      data_in_60_real <= io_data_in_payload_60_real;
      data_in_60_imag <= io_data_in_payload_60_imag;
      data_in_61_real <= io_data_in_payload_61_real;
      data_in_61_imag <= io_data_in_payload_61_imag;
      data_in_62_real <= io_data_in_payload_62_real;
      data_in_62_imag <= io_data_in_payload_62_imag;
      data_in_63_real <= io_data_in_payload_63_real;
      data_in_63_imag <= io_data_in_payload_63_imag;
      data_in_64_real <= io_data_in_payload_64_real;
      data_in_64_imag <= io_data_in_payload_64_imag;
      data_in_65_real <= io_data_in_payload_65_real;
      data_in_65_imag <= io_data_in_payload_65_imag;
      data_in_66_real <= io_data_in_payload_66_real;
      data_in_66_imag <= io_data_in_payload_66_imag;
      data_in_67_real <= io_data_in_payload_67_real;
      data_in_67_imag <= io_data_in_payload_67_imag;
      data_in_68_real <= io_data_in_payload_68_real;
      data_in_68_imag <= io_data_in_payload_68_imag;
      data_in_69_real <= io_data_in_payload_69_real;
      data_in_69_imag <= io_data_in_payload_69_imag;
      data_in_70_real <= io_data_in_payload_70_real;
      data_in_70_imag <= io_data_in_payload_70_imag;
      data_in_71_real <= io_data_in_payload_71_real;
      data_in_71_imag <= io_data_in_payload_71_imag;
      data_in_72_real <= io_data_in_payload_72_real;
      data_in_72_imag <= io_data_in_payload_72_imag;
      data_in_73_real <= io_data_in_payload_73_real;
      data_in_73_imag <= io_data_in_payload_73_imag;
      data_in_74_real <= io_data_in_payload_74_real;
      data_in_74_imag <= io_data_in_payload_74_imag;
      data_in_75_real <= io_data_in_payload_75_real;
      data_in_75_imag <= io_data_in_payload_75_imag;
      data_in_76_real <= io_data_in_payload_76_real;
      data_in_76_imag <= io_data_in_payload_76_imag;
      data_in_77_real <= io_data_in_payload_77_real;
      data_in_77_imag <= io_data_in_payload_77_imag;
      data_in_78_real <= io_data_in_payload_78_real;
      data_in_78_imag <= io_data_in_payload_78_imag;
      data_in_79_real <= io_data_in_payload_79_real;
      data_in_79_imag <= io_data_in_payload_79_imag;
      data_in_80_real <= io_data_in_payload_80_real;
      data_in_80_imag <= io_data_in_payload_80_imag;
      data_in_81_real <= io_data_in_payload_81_real;
      data_in_81_imag <= io_data_in_payload_81_imag;
      data_in_82_real <= io_data_in_payload_82_real;
      data_in_82_imag <= io_data_in_payload_82_imag;
      data_in_83_real <= io_data_in_payload_83_real;
      data_in_83_imag <= io_data_in_payload_83_imag;
      data_in_84_real <= io_data_in_payload_84_real;
      data_in_84_imag <= io_data_in_payload_84_imag;
      data_in_85_real <= io_data_in_payload_85_real;
      data_in_85_imag <= io_data_in_payload_85_imag;
      data_in_86_real <= io_data_in_payload_86_real;
      data_in_86_imag <= io_data_in_payload_86_imag;
      data_in_87_real <= io_data_in_payload_87_real;
      data_in_87_imag <= io_data_in_payload_87_imag;
      data_in_88_real <= io_data_in_payload_88_real;
      data_in_88_imag <= io_data_in_payload_88_imag;
      data_in_89_real <= io_data_in_payload_89_real;
      data_in_89_imag <= io_data_in_payload_89_imag;
      data_in_90_real <= io_data_in_payload_90_real;
      data_in_90_imag <= io_data_in_payload_90_imag;
      data_in_91_real <= io_data_in_payload_91_real;
      data_in_91_imag <= io_data_in_payload_91_imag;
      data_in_92_real <= io_data_in_payload_92_real;
      data_in_92_imag <= io_data_in_payload_92_imag;
      data_in_93_real <= io_data_in_payload_93_real;
      data_in_93_imag <= io_data_in_payload_93_imag;
      data_in_94_real <= io_data_in_payload_94_real;
      data_in_94_imag <= io_data_in_payload_94_imag;
      data_in_95_real <= io_data_in_payload_95_real;
      data_in_95_imag <= io_data_in_payload_95_imag;
      data_in_96_real <= io_data_in_payload_96_real;
      data_in_96_imag <= io_data_in_payload_96_imag;
      data_in_97_real <= io_data_in_payload_97_real;
      data_in_97_imag <= io_data_in_payload_97_imag;
      data_in_98_real <= io_data_in_payload_98_real;
      data_in_98_imag <= io_data_in_payload_98_imag;
      data_in_99_real <= io_data_in_payload_99_real;
      data_in_99_imag <= io_data_in_payload_99_imag;
      data_in_100_real <= io_data_in_payload_100_real;
      data_in_100_imag <= io_data_in_payload_100_imag;
      data_in_101_real <= io_data_in_payload_101_real;
      data_in_101_imag <= io_data_in_payload_101_imag;
      data_in_102_real <= io_data_in_payload_102_real;
      data_in_102_imag <= io_data_in_payload_102_imag;
      data_in_103_real <= io_data_in_payload_103_real;
      data_in_103_imag <= io_data_in_payload_103_imag;
      data_in_104_real <= io_data_in_payload_104_real;
      data_in_104_imag <= io_data_in_payload_104_imag;
      data_in_105_real <= io_data_in_payload_105_real;
      data_in_105_imag <= io_data_in_payload_105_imag;
      data_in_106_real <= io_data_in_payload_106_real;
      data_in_106_imag <= io_data_in_payload_106_imag;
      data_in_107_real <= io_data_in_payload_107_real;
      data_in_107_imag <= io_data_in_payload_107_imag;
      data_in_108_real <= io_data_in_payload_108_real;
      data_in_108_imag <= io_data_in_payload_108_imag;
      data_in_109_real <= io_data_in_payload_109_real;
      data_in_109_imag <= io_data_in_payload_109_imag;
      data_in_110_real <= io_data_in_payload_110_real;
      data_in_110_imag <= io_data_in_payload_110_imag;
      data_in_111_real <= io_data_in_payload_111_real;
      data_in_111_imag <= io_data_in_payload_111_imag;
      data_in_112_real <= io_data_in_payload_112_real;
      data_in_112_imag <= io_data_in_payload_112_imag;
      data_in_113_real <= io_data_in_payload_113_real;
      data_in_113_imag <= io_data_in_payload_113_imag;
      data_in_114_real <= io_data_in_payload_114_real;
      data_in_114_imag <= io_data_in_payload_114_imag;
      data_in_115_real <= io_data_in_payload_115_real;
      data_in_115_imag <= io_data_in_payload_115_imag;
      data_in_116_real <= io_data_in_payload_116_real;
      data_in_116_imag <= io_data_in_payload_116_imag;
      data_in_117_real <= io_data_in_payload_117_real;
      data_in_117_imag <= io_data_in_payload_117_imag;
      data_in_118_real <= io_data_in_payload_118_real;
      data_in_118_imag <= io_data_in_payload_118_imag;
      data_in_119_real <= io_data_in_payload_119_real;
      data_in_119_imag <= io_data_in_payload_119_imag;
      data_in_120_real <= io_data_in_payload_120_real;
      data_in_120_imag <= io_data_in_payload_120_imag;
      data_in_121_real <= io_data_in_payload_121_real;
      data_in_121_imag <= io_data_in_payload_121_imag;
      data_in_122_real <= io_data_in_payload_122_real;
      data_in_122_imag <= io_data_in_payload_122_imag;
      data_in_123_real <= io_data_in_payload_123_real;
      data_in_123_imag <= io_data_in_payload_123_imag;
      data_in_124_real <= io_data_in_payload_124_real;
      data_in_124_imag <= io_data_in_payload_124_imag;
      data_in_125_real <= io_data_in_payload_125_real;
      data_in_125_imag <= io_data_in_payload_125_imag;
      data_in_126_real <= io_data_in_payload_126_real;
      data_in_126_imag <= io_data_in_payload_126_imag;
      data_in_127_real <= io_data_in_payload_127_real;
      data_in_127_imag <= io_data_in_payload_127_imag;
    end
    _zz_3 <= _zz_5391[15 : 0];
    _zz_4 <= _zz_5395[15 : 0];
    _zz_1 <= _zz_5399[15 : 0];
    _zz_2 <= _zz_5403[15 : 0];
    _zz_7 <= _zz_5415[15 : 0];
    _zz_8 <= _zz_5419[15 : 0];
    _zz_5 <= _zz_5423[15 : 0];
    _zz_6 <= _zz_5427[15 : 0];
    _zz_11 <= _zz_5439[15 : 0];
    _zz_12 <= _zz_5443[15 : 0];
    _zz_9 <= _zz_5447[15 : 0];
    _zz_10 <= _zz_5451[15 : 0];
    _zz_15 <= _zz_5463[15 : 0];
    _zz_16 <= _zz_5467[15 : 0];
    _zz_13 <= _zz_5471[15 : 0];
    _zz_14 <= _zz_5475[15 : 0];
    _zz_19 <= _zz_5487[15 : 0];
    _zz_20 <= _zz_5491[15 : 0];
    _zz_17 <= _zz_5495[15 : 0];
    _zz_18 <= _zz_5499[15 : 0];
    _zz_23 <= _zz_5511[15 : 0];
    _zz_24 <= _zz_5515[15 : 0];
    _zz_21 <= _zz_5519[15 : 0];
    _zz_22 <= _zz_5523[15 : 0];
    _zz_27 <= _zz_5535[15 : 0];
    _zz_28 <= _zz_5539[15 : 0];
    _zz_25 <= _zz_5543[15 : 0];
    _zz_26 <= _zz_5547[15 : 0];
    _zz_31 <= _zz_5559[15 : 0];
    _zz_32 <= _zz_5563[15 : 0];
    _zz_29 <= _zz_5567[15 : 0];
    _zz_30 <= _zz_5571[15 : 0];
    _zz_35 <= _zz_5583[15 : 0];
    _zz_36 <= _zz_5587[15 : 0];
    _zz_33 <= _zz_5591[15 : 0];
    _zz_34 <= _zz_5595[15 : 0];
    _zz_39 <= _zz_5607[15 : 0];
    _zz_40 <= _zz_5611[15 : 0];
    _zz_37 <= _zz_5615[15 : 0];
    _zz_38 <= _zz_5619[15 : 0];
    _zz_43 <= _zz_5631[15 : 0];
    _zz_44 <= _zz_5635[15 : 0];
    _zz_41 <= _zz_5639[15 : 0];
    _zz_42 <= _zz_5643[15 : 0];
    _zz_47 <= _zz_5655[15 : 0];
    _zz_48 <= _zz_5659[15 : 0];
    _zz_45 <= _zz_5663[15 : 0];
    _zz_46 <= _zz_5667[15 : 0];
    _zz_51 <= _zz_5679[15 : 0];
    _zz_52 <= _zz_5683[15 : 0];
    _zz_49 <= _zz_5687[15 : 0];
    _zz_50 <= _zz_5691[15 : 0];
    _zz_55 <= _zz_5703[15 : 0];
    _zz_56 <= _zz_5707[15 : 0];
    _zz_53 <= _zz_5711[15 : 0];
    _zz_54 <= _zz_5715[15 : 0];
    _zz_59 <= _zz_5727[15 : 0];
    _zz_60 <= _zz_5731[15 : 0];
    _zz_57 <= _zz_5735[15 : 0];
    _zz_58 <= _zz_5739[15 : 0];
    _zz_63 <= _zz_5751[15 : 0];
    _zz_64 <= _zz_5755[15 : 0];
    _zz_61 <= _zz_5759[15 : 0];
    _zz_62 <= _zz_5763[15 : 0];
    _zz_67 <= _zz_5775[15 : 0];
    _zz_68 <= _zz_5779[15 : 0];
    _zz_65 <= _zz_5783[15 : 0];
    _zz_66 <= _zz_5787[15 : 0];
    _zz_71 <= _zz_5799[15 : 0];
    _zz_72 <= _zz_5803[15 : 0];
    _zz_69 <= _zz_5807[15 : 0];
    _zz_70 <= _zz_5811[15 : 0];
    _zz_75 <= _zz_5823[15 : 0];
    _zz_76 <= _zz_5827[15 : 0];
    _zz_73 <= _zz_5831[15 : 0];
    _zz_74 <= _zz_5835[15 : 0];
    _zz_79 <= _zz_5847[15 : 0];
    _zz_80 <= _zz_5851[15 : 0];
    _zz_77 <= _zz_5855[15 : 0];
    _zz_78 <= _zz_5859[15 : 0];
    _zz_83 <= _zz_5871[15 : 0];
    _zz_84 <= _zz_5875[15 : 0];
    _zz_81 <= _zz_5879[15 : 0];
    _zz_82 <= _zz_5883[15 : 0];
    _zz_87 <= _zz_5895[15 : 0];
    _zz_88 <= _zz_5899[15 : 0];
    _zz_85 <= _zz_5903[15 : 0];
    _zz_86 <= _zz_5907[15 : 0];
    _zz_91 <= _zz_5919[15 : 0];
    _zz_92 <= _zz_5923[15 : 0];
    _zz_89 <= _zz_5927[15 : 0];
    _zz_90 <= _zz_5931[15 : 0];
    _zz_95 <= _zz_5943[15 : 0];
    _zz_96 <= _zz_5947[15 : 0];
    _zz_93 <= _zz_5951[15 : 0];
    _zz_94 <= _zz_5955[15 : 0];
    _zz_99 <= _zz_5967[15 : 0];
    _zz_100 <= _zz_5971[15 : 0];
    _zz_97 <= _zz_5975[15 : 0];
    _zz_98 <= _zz_5979[15 : 0];
    _zz_103 <= _zz_5991[15 : 0];
    _zz_104 <= _zz_5995[15 : 0];
    _zz_101 <= _zz_5999[15 : 0];
    _zz_102 <= _zz_6003[15 : 0];
    _zz_107 <= _zz_6015[15 : 0];
    _zz_108 <= _zz_6019[15 : 0];
    _zz_105 <= _zz_6023[15 : 0];
    _zz_106 <= _zz_6027[15 : 0];
    _zz_111 <= _zz_6039[15 : 0];
    _zz_112 <= _zz_6043[15 : 0];
    _zz_109 <= _zz_6047[15 : 0];
    _zz_110 <= _zz_6051[15 : 0];
    _zz_115 <= _zz_6063[15 : 0];
    _zz_116 <= _zz_6067[15 : 0];
    _zz_113 <= _zz_6071[15 : 0];
    _zz_114 <= _zz_6075[15 : 0];
    _zz_119 <= _zz_6087[15 : 0];
    _zz_120 <= _zz_6091[15 : 0];
    _zz_117 <= _zz_6095[15 : 0];
    _zz_118 <= _zz_6099[15 : 0];
    _zz_123 <= _zz_6111[15 : 0];
    _zz_124 <= _zz_6115[15 : 0];
    _zz_121 <= _zz_6119[15 : 0];
    _zz_122 <= _zz_6123[15 : 0];
    _zz_127 <= _zz_6135[15 : 0];
    _zz_128 <= _zz_6139[15 : 0];
    _zz_125 <= _zz_6143[15 : 0];
    _zz_126 <= _zz_6147[15 : 0];
    _zz_131 <= _zz_6159[15 : 0];
    _zz_132 <= _zz_6163[15 : 0];
    _zz_129 <= _zz_6167[15 : 0];
    _zz_130 <= _zz_6171[15 : 0];
    _zz_135 <= _zz_6183[15 : 0];
    _zz_136 <= _zz_6187[15 : 0];
    _zz_133 <= _zz_6191[15 : 0];
    _zz_134 <= _zz_6195[15 : 0];
    _zz_139 <= _zz_6207[15 : 0];
    _zz_140 <= _zz_6211[15 : 0];
    _zz_137 <= _zz_6215[15 : 0];
    _zz_138 <= _zz_6219[15 : 0];
    _zz_143 <= _zz_6231[15 : 0];
    _zz_144 <= _zz_6235[15 : 0];
    _zz_141 <= _zz_6239[15 : 0];
    _zz_142 <= _zz_6243[15 : 0];
    _zz_147 <= _zz_6255[15 : 0];
    _zz_148 <= _zz_6259[15 : 0];
    _zz_145 <= _zz_6263[15 : 0];
    _zz_146 <= _zz_6267[15 : 0];
    _zz_151 <= _zz_6279[15 : 0];
    _zz_152 <= _zz_6283[15 : 0];
    _zz_149 <= _zz_6287[15 : 0];
    _zz_150 <= _zz_6291[15 : 0];
    _zz_155 <= _zz_6303[15 : 0];
    _zz_156 <= _zz_6307[15 : 0];
    _zz_153 <= _zz_6311[15 : 0];
    _zz_154 <= _zz_6315[15 : 0];
    _zz_159 <= _zz_6327[15 : 0];
    _zz_160 <= _zz_6331[15 : 0];
    _zz_157 <= _zz_6335[15 : 0];
    _zz_158 <= _zz_6339[15 : 0];
    _zz_163 <= _zz_6351[15 : 0];
    _zz_164 <= _zz_6355[15 : 0];
    _zz_161 <= _zz_6359[15 : 0];
    _zz_162 <= _zz_6363[15 : 0];
    _zz_167 <= _zz_6375[15 : 0];
    _zz_168 <= _zz_6379[15 : 0];
    _zz_165 <= _zz_6383[15 : 0];
    _zz_166 <= _zz_6387[15 : 0];
    _zz_171 <= _zz_6399[15 : 0];
    _zz_172 <= _zz_6403[15 : 0];
    _zz_169 <= _zz_6407[15 : 0];
    _zz_170 <= _zz_6411[15 : 0];
    _zz_175 <= _zz_6423[15 : 0];
    _zz_176 <= _zz_6427[15 : 0];
    _zz_173 <= _zz_6431[15 : 0];
    _zz_174 <= _zz_6435[15 : 0];
    _zz_179 <= _zz_6447[15 : 0];
    _zz_180 <= _zz_6451[15 : 0];
    _zz_177 <= _zz_6455[15 : 0];
    _zz_178 <= _zz_6459[15 : 0];
    _zz_183 <= _zz_6471[15 : 0];
    _zz_184 <= _zz_6475[15 : 0];
    _zz_181 <= _zz_6479[15 : 0];
    _zz_182 <= _zz_6483[15 : 0];
    _zz_187 <= _zz_6495[15 : 0];
    _zz_188 <= _zz_6499[15 : 0];
    _zz_185 <= _zz_6503[15 : 0];
    _zz_186 <= _zz_6507[15 : 0];
    _zz_191 <= _zz_6519[15 : 0];
    _zz_192 <= _zz_6523[15 : 0];
    _zz_189 <= _zz_6527[15 : 0];
    _zz_190 <= _zz_6531[15 : 0];
    _zz_195 <= _zz_6543[15 : 0];
    _zz_196 <= _zz_6547[15 : 0];
    _zz_193 <= _zz_6551[15 : 0];
    _zz_194 <= _zz_6555[15 : 0];
    _zz_199 <= _zz_6567[15 : 0];
    _zz_200 <= _zz_6571[15 : 0];
    _zz_197 <= _zz_6575[15 : 0];
    _zz_198 <= _zz_6579[15 : 0];
    _zz_203 <= _zz_6591[15 : 0];
    _zz_204 <= _zz_6595[15 : 0];
    _zz_201 <= _zz_6599[15 : 0];
    _zz_202 <= _zz_6603[15 : 0];
    _zz_207 <= _zz_6615[15 : 0];
    _zz_208 <= _zz_6619[15 : 0];
    _zz_205 <= _zz_6623[15 : 0];
    _zz_206 <= _zz_6627[15 : 0];
    _zz_211 <= _zz_6639[15 : 0];
    _zz_212 <= _zz_6643[15 : 0];
    _zz_209 <= _zz_6647[15 : 0];
    _zz_210 <= _zz_6651[15 : 0];
    _zz_215 <= _zz_6663[15 : 0];
    _zz_216 <= _zz_6667[15 : 0];
    _zz_213 <= _zz_6671[15 : 0];
    _zz_214 <= _zz_6675[15 : 0];
    _zz_219 <= _zz_6687[15 : 0];
    _zz_220 <= _zz_6691[15 : 0];
    _zz_217 <= _zz_6695[15 : 0];
    _zz_218 <= _zz_6699[15 : 0];
    _zz_223 <= _zz_6711[15 : 0];
    _zz_224 <= _zz_6715[15 : 0];
    _zz_221 <= _zz_6719[15 : 0];
    _zz_222 <= _zz_6723[15 : 0];
    _zz_227 <= _zz_6735[15 : 0];
    _zz_228 <= _zz_6739[15 : 0];
    _zz_225 <= _zz_6743[15 : 0];
    _zz_226 <= _zz_6747[15 : 0];
    _zz_231 <= _zz_6759[15 : 0];
    _zz_232 <= _zz_6763[15 : 0];
    _zz_229 <= _zz_6767[15 : 0];
    _zz_230 <= _zz_6771[15 : 0];
    _zz_235 <= _zz_6783[15 : 0];
    _zz_236 <= _zz_6787[15 : 0];
    _zz_233 <= _zz_6791[15 : 0];
    _zz_234 <= _zz_6795[15 : 0];
    _zz_239 <= _zz_6807[15 : 0];
    _zz_240 <= _zz_6811[15 : 0];
    _zz_237 <= _zz_6815[15 : 0];
    _zz_238 <= _zz_6819[15 : 0];
    _zz_243 <= _zz_6831[15 : 0];
    _zz_244 <= _zz_6835[15 : 0];
    _zz_241 <= _zz_6839[15 : 0];
    _zz_242 <= _zz_6843[15 : 0];
    _zz_247 <= _zz_6855[15 : 0];
    _zz_248 <= _zz_6859[15 : 0];
    _zz_245 <= _zz_6863[15 : 0];
    _zz_246 <= _zz_6867[15 : 0];
    _zz_251 <= _zz_6879[15 : 0];
    _zz_252 <= _zz_6883[15 : 0];
    _zz_249 <= _zz_6887[15 : 0];
    _zz_250 <= _zz_6891[15 : 0];
    _zz_255 <= _zz_6903[15 : 0];
    _zz_256 <= _zz_6907[15 : 0];
    _zz_253 <= _zz_6911[15 : 0];
    _zz_254 <= _zz_6915[15 : 0];
    _zz_261 <= _zz_6927[15 : 0];
    _zz_262 <= _zz_6931[15 : 0];
    _zz_257 <= _zz_6935[15 : 0];
    _zz_258 <= _zz_6939[15 : 0];
    _zz_263 <= _zz_6951[15 : 0];
    _zz_264 <= _zz_6955[15 : 0];
    _zz_259 <= _zz_6959[15 : 0];
    _zz_260 <= _zz_6963[15 : 0];
    _zz_269 <= _zz_6975[15 : 0];
    _zz_270 <= _zz_6979[15 : 0];
    _zz_265 <= _zz_6983[15 : 0];
    _zz_266 <= _zz_6987[15 : 0];
    _zz_271 <= _zz_6999[15 : 0];
    _zz_272 <= _zz_7003[15 : 0];
    _zz_267 <= _zz_7007[15 : 0];
    _zz_268 <= _zz_7011[15 : 0];
    _zz_277 <= _zz_7023[15 : 0];
    _zz_278 <= _zz_7027[15 : 0];
    _zz_273 <= _zz_7031[15 : 0];
    _zz_274 <= _zz_7035[15 : 0];
    _zz_279 <= _zz_7047[15 : 0];
    _zz_280 <= _zz_7051[15 : 0];
    _zz_275 <= _zz_7055[15 : 0];
    _zz_276 <= _zz_7059[15 : 0];
    _zz_285 <= _zz_7071[15 : 0];
    _zz_286 <= _zz_7075[15 : 0];
    _zz_281 <= _zz_7079[15 : 0];
    _zz_282 <= _zz_7083[15 : 0];
    _zz_287 <= _zz_7095[15 : 0];
    _zz_288 <= _zz_7099[15 : 0];
    _zz_283 <= _zz_7103[15 : 0];
    _zz_284 <= _zz_7107[15 : 0];
    _zz_293 <= _zz_7119[15 : 0];
    _zz_294 <= _zz_7123[15 : 0];
    _zz_289 <= _zz_7127[15 : 0];
    _zz_290 <= _zz_7131[15 : 0];
    _zz_295 <= _zz_7143[15 : 0];
    _zz_296 <= _zz_7147[15 : 0];
    _zz_291 <= _zz_7151[15 : 0];
    _zz_292 <= _zz_7155[15 : 0];
    _zz_301 <= _zz_7167[15 : 0];
    _zz_302 <= _zz_7171[15 : 0];
    _zz_297 <= _zz_7175[15 : 0];
    _zz_298 <= _zz_7179[15 : 0];
    _zz_303 <= _zz_7191[15 : 0];
    _zz_304 <= _zz_7195[15 : 0];
    _zz_299 <= _zz_7199[15 : 0];
    _zz_300 <= _zz_7203[15 : 0];
    _zz_309 <= _zz_7215[15 : 0];
    _zz_310 <= _zz_7219[15 : 0];
    _zz_305 <= _zz_7223[15 : 0];
    _zz_306 <= _zz_7227[15 : 0];
    _zz_311 <= _zz_7239[15 : 0];
    _zz_312 <= _zz_7243[15 : 0];
    _zz_307 <= _zz_7247[15 : 0];
    _zz_308 <= _zz_7251[15 : 0];
    _zz_317 <= _zz_7263[15 : 0];
    _zz_318 <= _zz_7267[15 : 0];
    _zz_313 <= _zz_7271[15 : 0];
    _zz_314 <= _zz_7275[15 : 0];
    _zz_319 <= _zz_7287[15 : 0];
    _zz_320 <= _zz_7291[15 : 0];
    _zz_315 <= _zz_7295[15 : 0];
    _zz_316 <= _zz_7299[15 : 0];
    _zz_325 <= _zz_7311[15 : 0];
    _zz_326 <= _zz_7315[15 : 0];
    _zz_321 <= _zz_7319[15 : 0];
    _zz_322 <= _zz_7323[15 : 0];
    _zz_327 <= _zz_7335[15 : 0];
    _zz_328 <= _zz_7339[15 : 0];
    _zz_323 <= _zz_7343[15 : 0];
    _zz_324 <= _zz_7347[15 : 0];
    _zz_333 <= _zz_7359[15 : 0];
    _zz_334 <= _zz_7363[15 : 0];
    _zz_329 <= _zz_7367[15 : 0];
    _zz_330 <= _zz_7371[15 : 0];
    _zz_335 <= _zz_7383[15 : 0];
    _zz_336 <= _zz_7387[15 : 0];
    _zz_331 <= _zz_7391[15 : 0];
    _zz_332 <= _zz_7395[15 : 0];
    _zz_341 <= _zz_7407[15 : 0];
    _zz_342 <= _zz_7411[15 : 0];
    _zz_337 <= _zz_7415[15 : 0];
    _zz_338 <= _zz_7419[15 : 0];
    _zz_343 <= _zz_7431[15 : 0];
    _zz_344 <= _zz_7435[15 : 0];
    _zz_339 <= _zz_7439[15 : 0];
    _zz_340 <= _zz_7443[15 : 0];
    _zz_349 <= _zz_7455[15 : 0];
    _zz_350 <= _zz_7459[15 : 0];
    _zz_345 <= _zz_7463[15 : 0];
    _zz_346 <= _zz_7467[15 : 0];
    _zz_351 <= _zz_7479[15 : 0];
    _zz_352 <= _zz_7483[15 : 0];
    _zz_347 <= _zz_7487[15 : 0];
    _zz_348 <= _zz_7491[15 : 0];
    _zz_357 <= _zz_7503[15 : 0];
    _zz_358 <= _zz_7507[15 : 0];
    _zz_353 <= _zz_7511[15 : 0];
    _zz_354 <= _zz_7515[15 : 0];
    _zz_359 <= _zz_7527[15 : 0];
    _zz_360 <= _zz_7531[15 : 0];
    _zz_355 <= _zz_7535[15 : 0];
    _zz_356 <= _zz_7539[15 : 0];
    _zz_365 <= _zz_7551[15 : 0];
    _zz_366 <= _zz_7555[15 : 0];
    _zz_361 <= _zz_7559[15 : 0];
    _zz_362 <= _zz_7563[15 : 0];
    _zz_367 <= _zz_7575[15 : 0];
    _zz_368 <= _zz_7579[15 : 0];
    _zz_363 <= _zz_7583[15 : 0];
    _zz_364 <= _zz_7587[15 : 0];
    _zz_373 <= _zz_7599[15 : 0];
    _zz_374 <= _zz_7603[15 : 0];
    _zz_369 <= _zz_7607[15 : 0];
    _zz_370 <= _zz_7611[15 : 0];
    _zz_375 <= _zz_7623[15 : 0];
    _zz_376 <= _zz_7627[15 : 0];
    _zz_371 <= _zz_7631[15 : 0];
    _zz_372 <= _zz_7635[15 : 0];
    _zz_381 <= _zz_7647[15 : 0];
    _zz_382 <= _zz_7651[15 : 0];
    _zz_377 <= _zz_7655[15 : 0];
    _zz_378 <= _zz_7659[15 : 0];
    _zz_383 <= _zz_7671[15 : 0];
    _zz_384 <= _zz_7675[15 : 0];
    _zz_379 <= _zz_7679[15 : 0];
    _zz_380 <= _zz_7683[15 : 0];
    _zz_389 <= _zz_7695[15 : 0];
    _zz_390 <= _zz_7699[15 : 0];
    _zz_385 <= _zz_7703[15 : 0];
    _zz_386 <= _zz_7707[15 : 0];
    _zz_391 <= _zz_7719[15 : 0];
    _zz_392 <= _zz_7723[15 : 0];
    _zz_387 <= _zz_7727[15 : 0];
    _zz_388 <= _zz_7731[15 : 0];
    _zz_397 <= _zz_7743[15 : 0];
    _zz_398 <= _zz_7747[15 : 0];
    _zz_393 <= _zz_7751[15 : 0];
    _zz_394 <= _zz_7755[15 : 0];
    _zz_399 <= _zz_7767[15 : 0];
    _zz_400 <= _zz_7771[15 : 0];
    _zz_395 <= _zz_7775[15 : 0];
    _zz_396 <= _zz_7779[15 : 0];
    _zz_405 <= _zz_7791[15 : 0];
    _zz_406 <= _zz_7795[15 : 0];
    _zz_401 <= _zz_7799[15 : 0];
    _zz_402 <= _zz_7803[15 : 0];
    _zz_407 <= _zz_7815[15 : 0];
    _zz_408 <= _zz_7819[15 : 0];
    _zz_403 <= _zz_7823[15 : 0];
    _zz_404 <= _zz_7827[15 : 0];
    _zz_413 <= _zz_7839[15 : 0];
    _zz_414 <= _zz_7843[15 : 0];
    _zz_409 <= _zz_7847[15 : 0];
    _zz_410 <= _zz_7851[15 : 0];
    _zz_415 <= _zz_7863[15 : 0];
    _zz_416 <= _zz_7867[15 : 0];
    _zz_411 <= _zz_7871[15 : 0];
    _zz_412 <= _zz_7875[15 : 0];
    _zz_421 <= _zz_7887[15 : 0];
    _zz_422 <= _zz_7891[15 : 0];
    _zz_417 <= _zz_7895[15 : 0];
    _zz_418 <= _zz_7899[15 : 0];
    _zz_423 <= _zz_7911[15 : 0];
    _zz_424 <= _zz_7915[15 : 0];
    _zz_419 <= _zz_7919[15 : 0];
    _zz_420 <= _zz_7923[15 : 0];
    _zz_429 <= _zz_7935[15 : 0];
    _zz_430 <= _zz_7939[15 : 0];
    _zz_425 <= _zz_7943[15 : 0];
    _zz_426 <= _zz_7947[15 : 0];
    _zz_431 <= _zz_7959[15 : 0];
    _zz_432 <= _zz_7963[15 : 0];
    _zz_427 <= _zz_7967[15 : 0];
    _zz_428 <= _zz_7971[15 : 0];
    _zz_437 <= _zz_7983[15 : 0];
    _zz_438 <= _zz_7987[15 : 0];
    _zz_433 <= _zz_7991[15 : 0];
    _zz_434 <= _zz_7995[15 : 0];
    _zz_439 <= _zz_8007[15 : 0];
    _zz_440 <= _zz_8011[15 : 0];
    _zz_435 <= _zz_8015[15 : 0];
    _zz_436 <= _zz_8019[15 : 0];
    _zz_445 <= _zz_8031[15 : 0];
    _zz_446 <= _zz_8035[15 : 0];
    _zz_441 <= _zz_8039[15 : 0];
    _zz_442 <= _zz_8043[15 : 0];
    _zz_447 <= _zz_8055[15 : 0];
    _zz_448 <= _zz_8059[15 : 0];
    _zz_443 <= _zz_8063[15 : 0];
    _zz_444 <= _zz_8067[15 : 0];
    _zz_453 <= _zz_8079[15 : 0];
    _zz_454 <= _zz_8083[15 : 0];
    _zz_449 <= _zz_8087[15 : 0];
    _zz_450 <= _zz_8091[15 : 0];
    _zz_455 <= _zz_8103[15 : 0];
    _zz_456 <= _zz_8107[15 : 0];
    _zz_451 <= _zz_8111[15 : 0];
    _zz_452 <= _zz_8115[15 : 0];
    _zz_461 <= _zz_8127[15 : 0];
    _zz_462 <= _zz_8131[15 : 0];
    _zz_457 <= _zz_8135[15 : 0];
    _zz_458 <= _zz_8139[15 : 0];
    _zz_463 <= _zz_8151[15 : 0];
    _zz_464 <= _zz_8155[15 : 0];
    _zz_459 <= _zz_8159[15 : 0];
    _zz_460 <= _zz_8163[15 : 0];
    _zz_469 <= _zz_8175[15 : 0];
    _zz_470 <= _zz_8179[15 : 0];
    _zz_465 <= _zz_8183[15 : 0];
    _zz_466 <= _zz_8187[15 : 0];
    _zz_471 <= _zz_8199[15 : 0];
    _zz_472 <= _zz_8203[15 : 0];
    _zz_467 <= _zz_8207[15 : 0];
    _zz_468 <= _zz_8211[15 : 0];
    _zz_477 <= _zz_8223[15 : 0];
    _zz_478 <= _zz_8227[15 : 0];
    _zz_473 <= _zz_8231[15 : 0];
    _zz_474 <= _zz_8235[15 : 0];
    _zz_479 <= _zz_8247[15 : 0];
    _zz_480 <= _zz_8251[15 : 0];
    _zz_475 <= _zz_8255[15 : 0];
    _zz_476 <= _zz_8259[15 : 0];
    _zz_485 <= _zz_8271[15 : 0];
    _zz_486 <= _zz_8275[15 : 0];
    _zz_481 <= _zz_8279[15 : 0];
    _zz_482 <= _zz_8283[15 : 0];
    _zz_487 <= _zz_8295[15 : 0];
    _zz_488 <= _zz_8299[15 : 0];
    _zz_483 <= _zz_8303[15 : 0];
    _zz_484 <= _zz_8307[15 : 0];
    _zz_493 <= _zz_8319[15 : 0];
    _zz_494 <= _zz_8323[15 : 0];
    _zz_489 <= _zz_8327[15 : 0];
    _zz_490 <= _zz_8331[15 : 0];
    _zz_495 <= _zz_8343[15 : 0];
    _zz_496 <= _zz_8347[15 : 0];
    _zz_491 <= _zz_8351[15 : 0];
    _zz_492 <= _zz_8355[15 : 0];
    _zz_501 <= _zz_8367[15 : 0];
    _zz_502 <= _zz_8371[15 : 0];
    _zz_497 <= _zz_8375[15 : 0];
    _zz_498 <= _zz_8379[15 : 0];
    _zz_503 <= _zz_8391[15 : 0];
    _zz_504 <= _zz_8395[15 : 0];
    _zz_499 <= _zz_8399[15 : 0];
    _zz_500 <= _zz_8403[15 : 0];
    _zz_509 <= _zz_8415[15 : 0];
    _zz_510 <= _zz_8419[15 : 0];
    _zz_505 <= _zz_8423[15 : 0];
    _zz_506 <= _zz_8427[15 : 0];
    _zz_511 <= _zz_8439[15 : 0];
    _zz_512 <= _zz_8443[15 : 0];
    _zz_507 <= _zz_8447[15 : 0];
    _zz_508 <= _zz_8451[15 : 0];
    _zz_521 <= _zz_8463[15 : 0];
    _zz_522 <= _zz_8467[15 : 0];
    _zz_513 <= _zz_8471[15 : 0];
    _zz_514 <= _zz_8475[15 : 0];
    _zz_523 <= _zz_8487[15 : 0];
    _zz_524 <= _zz_8491[15 : 0];
    _zz_515 <= _zz_8495[15 : 0];
    _zz_516 <= _zz_8499[15 : 0];
    _zz_525 <= _zz_8511[15 : 0];
    _zz_526 <= _zz_8515[15 : 0];
    _zz_517 <= _zz_8519[15 : 0];
    _zz_518 <= _zz_8523[15 : 0];
    _zz_527 <= _zz_8535[15 : 0];
    _zz_528 <= _zz_8539[15 : 0];
    _zz_519 <= _zz_8543[15 : 0];
    _zz_520 <= _zz_8547[15 : 0];
    _zz_537 <= _zz_8559[15 : 0];
    _zz_538 <= _zz_8563[15 : 0];
    _zz_529 <= _zz_8567[15 : 0];
    _zz_530 <= _zz_8571[15 : 0];
    _zz_539 <= _zz_8583[15 : 0];
    _zz_540 <= _zz_8587[15 : 0];
    _zz_531 <= _zz_8591[15 : 0];
    _zz_532 <= _zz_8595[15 : 0];
    _zz_541 <= _zz_8607[15 : 0];
    _zz_542 <= _zz_8611[15 : 0];
    _zz_533 <= _zz_8615[15 : 0];
    _zz_534 <= _zz_8619[15 : 0];
    _zz_543 <= _zz_8631[15 : 0];
    _zz_544 <= _zz_8635[15 : 0];
    _zz_535 <= _zz_8639[15 : 0];
    _zz_536 <= _zz_8643[15 : 0];
    _zz_553 <= _zz_8655[15 : 0];
    _zz_554 <= _zz_8659[15 : 0];
    _zz_545 <= _zz_8663[15 : 0];
    _zz_546 <= _zz_8667[15 : 0];
    _zz_555 <= _zz_8679[15 : 0];
    _zz_556 <= _zz_8683[15 : 0];
    _zz_547 <= _zz_8687[15 : 0];
    _zz_548 <= _zz_8691[15 : 0];
    _zz_557 <= _zz_8703[15 : 0];
    _zz_558 <= _zz_8707[15 : 0];
    _zz_549 <= _zz_8711[15 : 0];
    _zz_550 <= _zz_8715[15 : 0];
    _zz_559 <= _zz_8727[15 : 0];
    _zz_560 <= _zz_8731[15 : 0];
    _zz_551 <= _zz_8735[15 : 0];
    _zz_552 <= _zz_8739[15 : 0];
    _zz_569 <= _zz_8751[15 : 0];
    _zz_570 <= _zz_8755[15 : 0];
    _zz_561 <= _zz_8759[15 : 0];
    _zz_562 <= _zz_8763[15 : 0];
    _zz_571 <= _zz_8775[15 : 0];
    _zz_572 <= _zz_8779[15 : 0];
    _zz_563 <= _zz_8783[15 : 0];
    _zz_564 <= _zz_8787[15 : 0];
    _zz_573 <= _zz_8799[15 : 0];
    _zz_574 <= _zz_8803[15 : 0];
    _zz_565 <= _zz_8807[15 : 0];
    _zz_566 <= _zz_8811[15 : 0];
    _zz_575 <= _zz_8823[15 : 0];
    _zz_576 <= _zz_8827[15 : 0];
    _zz_567 <= _zz_8831[15 : 0];
    _zz_568 <= _zz_8835[15 : 0];
    _zz_585 <= _zz_8847[15 : 0];
    _zz_586 <= _zz_8851[15 : 0];
    _zz_577 <= _zz_8855[15 : 0];
    _zz_578 <= _zz_8859[15 : 0];
    _zz_587 <= _zz_8871[15 : 0];
    _zz_588 <= _zz_8875[15 : 0];
    _zz_579 <= _zz_8879[15 : 0];
    _zz_580 <= _zz_8883[15 : 0];
    _zz_589 <= _zz_8895[15 : 0];
    _zz_590 <= _zz_8899[15 : 0];
    _zz_581 <= _zz_8903[15 : 0];
    _zz_582 <= _zz_8907[15 : 0];
    _zz_591 <= _zz_8919[15 : 0];
    _zz_592 <= _zz_8923[15 : 0];
    _zz_583 <= _zz_8927[15 : 0];
    _zz_584 <= _zz_8931[15 : 0];
    _zz_601 <= _zz_8943[15 : 0];
    _zz_602 <= _zz_8947[15 : 0];
    _zz_593 <= _zz_8951[15 : 0];
    _zz_594 <= _zz_8955[15 : 0];
    _zz_603 <= _zz_8967[15 : 0];
    _zz_604 <= _zz_8971[15 : 0];
    _zz_595 <= _zz_8975[15 : 0];
    _zz_596 <= _zz_8979[15 : 0];
    _zz_605 <= _zz_8991[15 : 0];
    _zz_606 <= _zz_8995[15 : 0];
    _zz_597 <= _zz_8999[15 : 0];
    _zz_598 <= _zz_9003[15 : 0];
    _zz_607 <= _zz_9015[15 : 0];
    _zz_608 <= _zz_9019[15 : 0];
    _zz_599 <= _zz_9023[15 : 0];
    _zz_600 <= _zz_9027[15 : 0];
    _zz_617 <= _zz_9039[15 : 0];
    _zz_618 <= _zz_9043[15 : 0];
    _zz_609 <= _zz_9047[15 : 0];
    _zz_610 <= _zz_9051[15 : 0];
    _zz_619 <= _zz_9063[15 : 0];
    _zz_620 <= _zz_9067[15 : 0];
    _zz_611 <= _zz_9071[15 : 0];
    _zz_612 <= _zz_9075[15 : 0];
    _zz_621 <= _zz_9087[15 : 0];
    _zz_622 <= _zz_9091[15 : 0];
    _zz_613 <= _zz_9095[15 : 0];
    _zz_614 <= _zz_9099[15 : 0];
    _zz_623 <= _zz_9111[15 : 0];
    _zz_624 <= _zz_9115[15 : 0];
    _zz_615 <= _zz_9119[15 : 0];
    _zz_616 <= _zz_9123[15 : 0];
    _zz_633 <= _zz_9135[15 : 0];
    _zz_634 <= _zz_9139[15 : 0];
    _zz_625 <= _zz_9143[15 : 0];
    _zz_626 <= _zz_9147[15 : 0];
    _zz_635 <= _zz_9159[15 : 0];
    _zz_636 <= _zz_9163[15 : 0];
    _zz_627 <= _zz_9167[15 : 0];
    _zz_628 <= _zz_9171[15 : 0];
    _zz_637 <= _zz_9183[15 : 0];
    _zz_638 <= _zz_9187[15 : 0];
    _zz_629 <= _zz_9191[15 : 0];
    _zz_630 <= _zz_9195[15 : 0];
    _zz_639 <= _zz_9207[15 : 0];
    _zz_640 <= _zz_9211[15 : 0];
    _zz_631 <= _zz_9215[15 : 0];
    _zz_632 <= _zz_9219[15 : 0];
    _zz_649 <= _zz_9231[15 : 0];
    _zz_650 <= _zz_9235[15 : 0];
    _zz_641 <= _zz_9239[15 : 0];
    _zz_642 <= _zz_9243[15 : 0];
    _zz_651 <= _zz_9255[15 : 0];
    _zz_652 <= _zz_9259[15 : 0];
    _zz_643 <= _zz_9263[15 : 0];
    _zz_644 <= _zz_9267[15 : 0];
    _zz_653 <= _zz_9279[15 : 0];
    _zz_654 <= _zz_9283[15 : 0];
    _zz_645 <= _zz_9287[15 : 0];
    _zz_646 <= _zz_9291[15 : 0];
    _zz_655 <= _zz_9303[15 : 0];
    _zz_656 <= _zz_9307[15 : 0];
    _zz_647 <= _zz_9311[15 : 0];
    _zz_648 <= _zz_9315[15 : 0];
    _zz_665 <= _zz_9327[15 : 0];
    _zz_666 <= _zz_9331[15 : 0];
    _zz_657 <= _zz_9335[15 : 0];
    _zz_658 <= _zz_9339[15 : 0];
    _zz_667 <= _zz_9351[15 : 0];
    _zz_668 <= _zz_9355[15 : 0];
    _zz_659 <= _zz_9359[15 : 0];
    _zz_660 <= _zz_9363[15 : 0];
    _zz_669 <= _zz_9375[15 : 0];
    _zz_670 <= _zz_9379[15 : 0];
    _zz_661 <= _zz_9383[15 : 0];
    _zz_662 <= _zz_9387[15 : 0];
    _zz_671 <= _zz_9399[15 : 0];
    _zz_672 <= _zz_9403[15 : 0];
    _zz_663 <= _zz_9407[15 : 0];
    _zz_664 <= _zz_9411[15 : 0];
    _zz_681 <= _zz_9423[15 : 0];
    _zz_682 <= _zz_9427[15 : 0];
    _zz_673 <= _zz_9431[15 : 0];
    _zz_674 <= _zz_9435[15 : 0];
    _zz_683 <= _zz_9447[15 : 0];
    _zz_684 <= _zz_9451[15 : 0];
    _zz_675 <= _zz_9455[15 : 0];
    _zz_676 <= _zz_9459[15 : 0];
    _zz_685 <= _zz_9471[15 : 0];
    _zz_686 <= _zz_9475[15 : 0];
    _zz_677 <= _zz_9479[15 : 0];
    _zz_678 <= _zz_9483[15 : 0];
    _zz_687 <= _zz_9495[15 : 0];
    _zz_688 <= _zz_9499[15 : 0];
    _zz_679 <= _zz_9503[15 : 0];
    _zz_680 <= _zz_9507[15 : 0];
    _zz_697 <= _zz_9519[15 : 0];
    _zz_698 <= _zz_9523[15 : 0];
    _zz_689 <= _zz_9527[15 : 0];
    _zz_690 <= _zz_9531[15 : 0];
    _zz_699 <= _zz_9543[15 : 0];
    _zz_700 <= _zz_9547[15 : 0];
    _zz_691 <= _zz_9551[15 : 0];
    _zz_692 <= _zz_9555[15 : 0];
    _zz_701 <= _zz_9567[15 : 0];
    _zz_702 <= _zz_9571[15 : 0];
    _zz_693 <= _zz_9575[15 : 0];
    _zz_694 <= _zz_9579[15 : 0];
    _zz_703 <= _zz_9591[15 : 0];
    _zz_704 <= _zz_9595[15 : 0];
    _zz_695 <= _zz_9599[15 : 0];
    _zz_696 <= _zz_9603[15 : 0];
    _zz_713 <= _zz_9615[15 : 0];
    _zz_714 <= _zz_9619[15 : 0];
    _zz_705 <= _zz_9623[15 : 0];
    _zz_706 <= _zz_9627[15 : 0];
    _zz_715 <= _zz_9639[15 : 0];
    _zz_716 <= _zz_9643[15 : 0];
    _zz_707 <= _zz_9647[15 : 0];
    _zz_708 <= _zz_9651[15 : 0];
    _zz_717 <= _zz_9663[15 : 0];
    _zz_718 <= _zz_9667[15 : 0];
    _zz_709 <= _zz_9671[15 : 0];
    _zz_710 <= _zz_9675[15 : 0];
    _zz_719 <= _zz_9687[15 : 0];
    _zz_720 <= _zz_9691[15 : 0];
    _zz_711 <= _zz_9695[15 : 0];
    _zz_712 <= _zz_9699[15 : 0];
    _zz_729 <= _zz_9711[15 : 0];
    _zz_730 <= _zz_9715[15 : 0];
    _zz_721 <= _zz_9719[15 : 0];
    _zz_722 <= _zz_9723[15 : 0];
    _zz_731 <= _zz_9735[15 : 0];
    _zz_732 <= _zz_9739[15 : 0];
    _zz_723 <= _zz_9743[15 : 0];
    _zz_724 <= _zz_9747[15 : 0];
    _zz_733 <= _zz_9759[15 : 0];
    _zz_734 <= _zz_9763[15 : 0];
    _zz_725 <= _zz_9767[15 : 0];
    _zz_726 <= _zz_9771[15 : 0];
    _zz_735 <= _zz_9783[15 : 0];
    _zz_736 <= _zz_9787[15 : 0];
    _zz_727 <= _zz_9791[15 : 0];
    _zz_728 <= _zz_9795[15 : 0];
    _zz_745 <= _zz_9807[15 : 0];
    _zz_746 <= _zz_9811[15 : 0];
    _zz_737 <= _zz_9815[15 : 0];
    _zz_738 <= _zz_9819[15 : 0];
    _zz_747 <= _zz_9831[15 : 0];
    _zz_748 <= _zz_9835[15 : 0];
    _zz_739 <= _zz_9839[15 : 0];
    _zz_740 <= _zz_9843[15 : 0];
    _zz_749 <= _zz_9855[15 : 0];
    _zz_750 <= _zz_9859[15 : 0];
    _zz_741 <= _zz_9863[15 : 0];
    _zz_742 <= _zz_9867[15 : 0];
    _zz_751 <= _zz_9879[15 : 0];
    _zz_752 <= _zz_9883[15 : 0];
    _zz_743 <= _zz_9887[15 : 0];
    _zz_744 <= _zz_9891[15 : 0];
    _zz_761 <= _zz_9903[15 : 0];
    _zz_762 <= _zz_9907[15 : 0];
    _zz_753 <= _zz_9911[15 : 0];
    _zz_754 <= _zz_9915[15 : 0];
    _zz_763 <= _zz_9927[15 : 0];
    _zz_764 <= _zz_9931[15 : 0];
    _zz_755 <= _zz_9935[15 : 0];
    _zz_756 <= _zz_9939[15 : 0];
    _zz_765 <= _zz_9951[15 : 0];
    _zz_766 <= _zz_9955[15 : 0];
    _zz_757 <= _zz_9959[15 : 0];
    _zz_758 <= _zz_9963[15 : 0];
    _zz_767 <= _zz_9975[15 : 0];
    _zz_768 <= _zz_9979[15 : 0];
    _zz_759 <= _zz_9983[15 : 0];
    _zz_760 <= _zz_9987[15 : 0];
    _zz_785 <= _zz_9999[15 : 0];
    _zz_786 <= _zz_10003[15 : 0];
    _zz_769 <= _zz_10007[15 : 0];
    _zz_770 <= _zz_10011[15 : 0];
    _zz_787 <= _zz_10023[15 : 0];
    _zz_788 <= _zz_10027[15 : 0];
    _zz_771 <= _zz_10031[15 : 0];
    _zz_772 <= _zz_10035[15 : 0];
    _zz_789 <= _zz_10047[15 : 0];
    _zz_790 <= _zz_10051[15 : 0];
    _zz_773 <= _zz_10055[15 : 0];
    _zz_774 <= _zz_10059[15 : 0];
    _zz_791 <= _zz_10071[15 : 0];
    _zz_792 <= _zz_10075[15 : 0];
    _zz_775 <= _zz_10079[15 : 0];
    _zz_776 <= _zz_10083[15 : 0];
    _zz_793 <= _zz_10095[15 : 0];
    _zz_794 <= _zz_10099[15 : 0];
    _zz_777 <= _zz_10103[15 : 0];
    _zz_778 <= _zz_10107[15 : 0];
    _zz_795 <= _zz_10119[15 : 0];
    _zz_796 <= _zz_10123[15 : 0];
    _zz_779 <= _zz_10127[15 : 0];
    _zz_780 <= _zz_10131[15 : 0];
    _zz_797 <= _zz_10143[15 : 0];
    _zz_798 <= _zz_10147[15 : 0];
    _zz_781 <= _zz_10151[15 : 0];
    _zz_782 <= _zz_10155[15 : 0];
    _zz_799 <= _zz_10167[15 : 0];
    _zz_800 <= _zz_10171[15 : 0];
    _zz_783 <= _zz_10175[15 : 0];
    _zz_784 <= _zz_10179[15 : 0];
    _zz_817 <= _zz_10191[15 : 0];
    _zz_818 <= _zz_10195[15 : 0];
    _zz_801 <= _zz_10199[15 : 0];
    _zz_802 <= _zz_10203[15 : 0];
    _zz_819 <= _zz_10215[15 : 0];
    _zz_820 <= _zz_10219[15 : 0];
    _zz_803 <= _zz_10223[15 : 0];
    _zz_804 <= _zz_10227[15 : 0];
    _zz_821 <= _zz_10239[15 : 0];
    _zz_822 <= _zz_10243[15 : 0];
    _zz_805 <= _zz_10247[15 : 0];
    _zz_806 <= _zz_10251[15 : 0];
    _zz_823 <= _zz_10263[15 : 0];
    _zz_824 <= _zz_10267[15 : 0];
    _zz_807 <= _zz_10271[15 : 0];
    _zz_808 <= _zz_10275[15 : 0];
    _zz_825 <= _zz_10287[15 : 0];
    _zz_826 <= _zz_10291[15 : 0];
    _zz_809 <= _zz_10295[15 : 0];
    _zz_810 <= _zz_10299[15 : 0];
    _zz_827 <= _zz_10311[15 : 0];
    _zz_828 <= _zz_10315[15 : 0];
    _zz_811 <= _zz_10319[15 : 0];
    _zz_812 <= _zz_10323[15 : 0];
    _zz_829 <= _zz_10335[15 : 0];
    _zz_830 <= _zz_10339[15 : 0];
    _zz_813 <= _zz_10343[15 : 0];
    _zz_814 <= _zz_10347[15 : 0];
    _zz_831 <= _zz_10359[15 : 0];
    _zz_832 <= _zz_10363[15 : 0];
    _zz_815 <= _zz_10367[15 : 0];
    _zz_816 <= _zz_10371[15 : 0];
    _zz_849 <= _zz_10383[15 : 0];
    _zz_850 <= _zz_10387[15 : 0];
    _zz_833 <= _zz_10391[15 : 0];
    _zz_834 <= _zz_10395[15 : 0];
    _zz_851 <= _zz_10407[15 : 0];
    _zz_852 <= _zz_10411[15 : 0];
    _zz_835 <= _zz_10415[15 : 0];
    _zz_836 <= _zz_10419[15 : 0];
    _zz_853 <= _zz_10431[15 : 0];
    _zz_854 <= _zz_10435[15 : 0];
    _zz_837 <= _zz_10439[15 : 0];
    _zz_838 <= _zz_10443[15 : 0];
    _zz_855 <= _zz_10455[15 : 0];
    _zz_856 <= _zz_10459[15 : 0];
    _zz_839 <= _zz_10463[15 : 0];
    _zz_840 <= _zz_10467[15 : 0];
    _zz_857 <= _zz_10479[15 : 0];
    _zz_858 <= _zz_10483[15 : 0];
    _zz_841 <= _zz_10487[15 : 0];
    _zz_842 <= _zz_10491[15 : 0];
    _zz_859 <= _zz_10503[15 : 0];
    _zz_860 <= _zz_10507[15 : 0];
    _zz_843 <= _zz_10511[15 : 0];
    _zz_844 <= _zz_10515[15 : 0];
    _zz_861 <= _zz_10527[15 : 0];
    _zz_862 <= _zz_10531[15 : 0];
    _zz_845 <= _zz_10535[15 : 0];
    _zz_846 <= _zz_10539[15 : 0];
    _zz_863 <= _zz_10551[15 : 0];
    _zz_864 <= _zz_10555[15 : 0];
    _zz_847 <= _zz_10559[15 : 0];
    _zz_848 <= _zz_10563[15 : 0];
    _zz_881 <= _zz_10575[15 : 0];
    _zz_882 <= _zz_10579[15 : 0];
    _zz_865 <= _zz_10583[15 : 0];
    _zz_866 <= _zz_10587[15 : 0];
    _zz_883 <= _zz_10599[15 : 0];
    _zz_884 <= _zz_10603[15 : 0];
    _zz_867 <= _zz_10607[15 : 0];
    _zz_868 <= _zz_10611[15 : 0];
    _zz_885 <= _zz_10623[15 : 0];
    _zz_886 <= _zz_10627[15 : 0];
    _zz_869 <= _zz_10631[15 : 0];
    _zz_870 <= _zz_10635[15 : 0];
    _zz_887 <= _zz_10647[15 : 0];
    _zz_888 <= _zz_10651[15 : 0];
    _zz_871 <= _zz_10655[15 : 0];
    _zz_872 <= _zz_10659[15 : 0];
    _zz_889 <= _zz_10671[15 : 0];
    _zz_890 <= _zz_10675[15 : 0];
    _zz_873 <= _zz_10679[15 : 0];
    _zz_874 <= _zz_10683[15 : 0];
    _zz_891 <= _zz_10695[15 : 0];
    _zz_892 <= _zz_10699[15 : 0];
    _zz_875 <= _zz_10703[15 : 0];
    _zz_876 <= _zz_10707[15 : 0];
    _zz_893 <= _zz_10719[15 : 0];
    _zz_894 <= _zz_10723[15 : 0];
    _zz_877 <= _zz_10727[15 : 0];
    _zz_878 <= _zz_10731[15 : 0];
    _zz_895 <= _zz_10743[15 : 0];
    _zz_896 <= _zz_10747[15 : 0];
    _zz_879 <= _zz_10751[15 : 0];
    _zz_880 <= _zz_10755[15 : 0];
    _zz_913 <= _zz_10767[15 : 0];
    _zz_914 <= _zz_10771[15 : 0];
    _zz_897 <= _zz_10775[15 : 0];
    _zz_898 <= _zz_10779[15 : 0];
    _zz_915 <= _zz_10791[15 : 0];
    _zz_916 <= _zz_10795[15 : 0];
    _zz_899 <= _zz_10799[15 : 0];
    _zz_900 <= _zz_10803[15 : 0];
    _zz_917 <= _zz_10815[15 : 0];
    _zz_918 <= _zz_10819[15 : 0];
    _zz_901 <= _zz_10823[15 : 0];
    _zz_902 <= _zz_10827[15 : 0];
    _zz_919 <= _zz_10839[15 : 0];
    _zz_920 <= _zz_10843[15 : 0];
    _zz_903 <= _zz_10847[15 : 0];
    _zz_904 <= _zz_10851[15 : 0];
    _zz_921 <= _zz_10863[15 : 0];
    _zz_922 <= _zz_10867[15 : 0];
    _zz_905 <= _zz_10871[15 : 0];
    _zz_906 <= _zz_10875[15 : 0];
    _zz_923 <= _zz_10887[15 : 0];
    _zz_924 <= _zz_10891[15 : 0];
    _zz_907 <= _zz_10895[15 : 0];
    _zz_908 <= _zz_10899[15 : 0];
    _zz_925 <= _zz_10911[15 : 0];
    _zz_926 <= _zz_10915[15 : 0];
    _zz_909 <= _zz_10919[15 : 0];
    _zz_910 <= _zz_10923[15 : 0];
    _zz_927 <= _zz_10935[15 : 0];
    _zz_928 <= _zz_10939[15 : 0];
    _zz_911 <= _zz_10943[15 : 0];
    _zz_912 <= _zz_10947[15 : 0];
    _zz_945 <= _zz_10959[15 : 0];
    _zz_946 <= _zz_10963[15 : 0];
    _zz_929 <= _zz_10967[15 : 0];
    _zz_930 <= _zz_10971[15 : 0];
    _zz_947 <= _zz_10983[15 : 0];
    _zz_948 <= _zz_10987[15 : 0];
    _zz_931 <= _zz_10991[15 : 0];
    _zz_932 <= _zz_10995[15 : 0];
    _zz_949 <= _zz_11007[15 : 0];
    _zz_950 <= _zz_11011[15 : 0];
    _zz_933 <= _zz_11015[15 : 0];
    _zz_934 <= _zz_11019[15 : 0];
    _zz_951 <= _zz_11031[15 : 0];
    _zz_952 <= _zz_11035[15 : 0];
    _zz_935 <= _zz_11039[15 : 0];
    _zz_936 <= _zz_11043[15 : 0];
    _zz_953 <= _zz_11055[15 : 0];
    _zz_954 <= _zz_11059[15 : 0];
    _zz_937 <= _zz_11063[15 : 0];
    _zz_938 <= _zz_11067[15 : 0];
    _zz_955 <= _zz_11079[15 : 0];
    _zz_956 <= _zz_11083[15 : 0];
    _zz_939 <= _zz_11087[15 : 0];
    _zz_940 <= _zz_11091[15 : 0];
    _zz_957 <= _zz_11103[15 : 0];
    _zz_958 <= _zz_11107[15 : 0];
    _zz_941 <= _zz_11111[15 : 0];
    _zz_942 <= _zz_11115[15 : 0];
    _zz_959 <= _zz_11127[15 : 0];
    _zz_960 <= _zz_11131[15 : 0];
    _zz_943 <= _zz_11135[15 : 0];
    _zz_944 <= _zz_11139[15 : 0];
    _zz_977 <= _zz_11151[15 : 0];
    _zz_978 <= _zz_11155[15 : 0];
    _zz_961 <= _zz_11159[15 : 0];
    _zz_962 <= _zz_11163[15 : 0];
    _zz_979 <= _zz_11175[15 : 0];
    _zz_980 <= _zz_11179[15 : 0];
    _zz_963 <= _zz_11183[15 : 0];
    _zz_964 <= _zz_11187[15 : 0];
    _zz_981 <= _zz_11199[15 : 0];
    _zz_982 <= _zz_11203[15 : 0];
    _zz_965 <= _zz_11207[15 : 0];
    _zz_966 <= _zz_11211[15 : 0];
    _zz_983 <= _zz_11223[15 : 0];
    _zz_984 <= _zz_11227[15 : 0];
    _zz_967 <= _zz_11231[15 : 0];
    _zz_968 <= _zz_11235[15 : 0];
    _zz_985 <= _zz_11247[15 : 0];
    _zz_986 <= _zz_11251[15 : 0];
    _zz_969 <= _zz_11255[15 : 0];
    _zz_970 <= _zz_11259[15 : 0];
    _zz_987 <= _zz_11271[15 : 0];
    _zz_988 <= _zz_11275[15 : 0];
    _zz_971 <= _zz_11279[15 : 0];
    _zz_972 <= _zz_11283[15 : 0];
    _zz_989 <= _zz_11295[15 : 0];
    _zz_990 <= _zz_11299[15 : 0];
    _zz_973 <= _zz_11303[15 : 0];
    _zz_974 <= _zz_11307[15 : 0];
    _zz_991 <= _zz_11319[15 : 0];
    _zz_992 <= _zz_11323[15 : 0];
    _zz_975 <= _zz_11327[15 : 0];
    _zz_976 <= _zz_11331[15 : 0];
    _zz_1009 <= _zz_11343[15 : 0];
    _zz_1010 <= _zz_11347[15 : 0];
    _zz_993 <= _zz_11351[15 : 0];
    _zz_994 <= _zz_11355[15 : 0];
    _zz_1011 <= _zz_11367[15 : 0];
    _zz_1012 <= _zz_11371[15 : 0];
    _zz_995 <= _zz_11375[15 : 0];
    _zz_996 <= _zz_11379[15 : 0];
    _zz_1013 <= _zz_11391[15 : 0];
    _zz_1014 <= _zz_11395[15 : 0];
    _zz_997 <= _zz_11399[15 : 0];
    _zz_998 <= _zz_11403[15 : 0];
    _zz_1015 <= _zz_11415[15 : 0];
    _zz_1016 <= _zz_11419[15 : 0];
    _zz_999 <= _zz_11423[15 : 0];
    _zz_1000 <= _zz_11427[15 : 0];
    _zz_1017 <= _zz_11439[15 : 0];
    _zz_1018 <= _zz_11443[15 : 0];
    _zz_1001 <= _zz_11447[15 : 0];
    _zz_1002 <= _zz_11451[15 : 0];
    _zz_1019 <= _zz_11463[15 : 0];
    _zz_1020 <= _zz_11467[15 : 0];
    _zz_1003 <= _zz_11471[15 : 0];
    _zz_1004 <= _zz_11475[15 : 0];
    _zz_1021 <= _zz_11487[15 : 0];
    _zz_1022 <= _zz_11491[15 : 0];
    _zz_1005 <= _zz_11495[15 : 0];
    _zz_1006 <= _zz_11499[15 : 0];
    _zz_1023 <= _zz_11511[15 : 0];
    _zz_1024 <= _zz_11515[15 : 0];
    _zz_1007 <= _zz_11519[15 : 0];
    _zz_1008 <= _zz_11523[15 : 0];
    _zz_1057 <= _zz_11535[15 : 0];
    _zz_1058 <= _zz_11539[15 : 0];
    _zz_1025 <= _zz_11543[15 : 0];
    _zz_1026 <= _zz_11547[15 : 0];
    _zz_1059 <= _zz_11559[15 : 0];
    _zz_1060 <= _zz_11563[15 : 0];
    _zz_1027 <= _zz_11567[15 : 0];
    _zz_1028 <= _zz_11571[15 : 0];
    _zz_1061 <= _zz_11583[15 : 0];
    _zz_1062 <= _zz_11587[15 : 0];
    _zz_1029 <= _zz_11591[15 : 0];
    _zz_1030 <= _zz_11595[15 : 0];
    _zz_1063 <= _zz_11607[15 : 0];
    _zz_1064 <= _zz_11611[15 : 0];
    _zz_1031 <= _zz_11615[15 : 0];
    _zz_1032 <= _zz_11619[15 : 0];
    _zz_1065 <= _zz_11631[15 : 0];
    _zz_1066 <= _zz_11635[15 : 0];
    _zz_1033 <= _zz_11639[15 : 0];
    _zz_1034 <= _zz_11643[15 : 0];
    _zz_1067 <= _zz_11655[15 : 0];
    _zz_1068 <= _zz_11659[15 : 0];
    _zz_1035 <= _zz_11663[15 : 0];
    _zz_1036 <= _zz_11667[15 : 0];
    _zz_1069 <= _zz_11679[15 : 0];
    _zz_1070 <= _zz_11683[15 : 0];
    _zz_1037 <= _zz_11687[15 : 0];
    _zz_1038 <= _zz_11691[15 : 0];
    _zz_1071 <= _zz_11703[15 : 0];
    _zz_1072 <= _zz_11707[15 : 0];
    _zz_1039 <= _zz_11711[15 : 0];
    _zz_1040 <= _zz_11715[15 : 0];
    _zz_1073 <= _zz_11727[15 : 0];
    _zz_1074 <= _zz_11731[15 : 0];
    _zz_1041 <= _zz_11735[15 : 0];
    _zz_1042 <= _zz_11739[15 : 0];
    _zz_1075 <= _zz_11751[15 : 0];
    _zz_1076 <= _zz_11755[15 : 0];
    _zz_1043 <= _zz_11759[15 : 0];
    _zz_1044 <= _zz_11763[15 : 0];
    _zz_1077 <= _zz_11775[15 : 0];
    _zz_1078 <= _zz_11779[15 : 0];
    _zz_1045 <= _zz_11783[15 : 0];
    _zz_1046 <= _zz_11787[15 : 0];
    _zz_1079 <= _zz_11799[15 : 0];
    _zz_1080 <= _zz_11803[15 : 0];
    _zz_1047 <= _zz_11807[15 : 0];
    _zz_1048 <= _zz_11811[15 : 0];
    _zz_1081 <= _zz_11823[15 : 0];
    _zz_1082 <= _zz_11827[15 : 0];
    _zz_1049 <= _zz_11831[15 : 0];
    _zz_1050 <= _zz_11835[15 : 0];
    _zz_1083 <= _zz_11847[15 : 0];
    _zz_1084 <= _zz_11851[15 : 0];
    _zz_1051 <= _zz_11855[15 : 0];
    _zz_1052 <= _zz_11859[15 : 0];
    _zz_1085 <= _zz_11871[15 : 0];
    _zz_1086 <= _zz_11875[15 : 0];
    _zz_1053 <= _zz_11879[15 : 0];
    _zz_1054 <= _zz_11883[15 : 0];
    _zz_1087 <= _zz_11895[15 : 0];
    _zz_1088 <= _zz_11899[15 : 0];
    _zz_1055 <= _zz_11903[15 : 0];
    _zz_1056 <= _zz_11907[15 : 0];
    _zz_1121 <= _zz_11919[15 : 0];
    _zz_1122 <= _zz_11923[15 : 0];
    _zz_1089 <= _zz_11927[15 : 0];
    _zz_1090 <= _zz_11931[15 : 0];
    _zz_1123 <= _zz_11943[15 : 0];
    _zz_1124 <= _zz_11947[15 : 0];
    _zz_1091 <= _zz_11951[15 : 0];
    _zz_1092 <= _zz_11955[15 : 0];
    _zz_1125 <= _zz_11967[15 : 0];
    _zz_1126 <= _zz_11971[15 : 0];
    _zz_1093 <= _zz_11975[15 : 0];
    _zz_1094 <= _zz_11979[15 : 0];
    _zz_1127 <= _zz_11991[15 : 0];
    _zz_1128 <= _zz_11995[15 : 0];
    _zz_1095 <= _zz_11999[15 : 0];
    _zz_1096 <= _zz_12003[15 : 0];
    _zz_1129 <= _zz_12015[15 : 0];
    _zz_1130 <= _zz_12019[15 : 0];
    _zz_1097 <= _zz_12023[15 : 0];
    _zz_1098 <= _zz_12027[15 : 0];
    _zz_1131 <= _zz_12039[15 : 0];
    _zz_1132 <= _zz_12043[15 : 0];
    _zz_1099 <= _zz_12047[15 : 0];
    _zz_1100 <= _zz_12051[15 : 0];
    _zz_1133 <= _zz_12063[15 : 0];
    _zz_1134 <= _zz_12067[15 : 0];
    _zz_1101 <= _zz_12071[15 : 0];
    _zz_1102 <= _zz_12075[15 : 0];
    _zz_1135 <= _zz_12087[15 : 0];
    _zz_1136 <= _zz_12091[15 : 0];
    _zz_1103 <= _zz_12095[15 : 0];
    _zz_1104 <= _zz_12099[15 : 0];
    _zz_1137 <= _zz_12111[15 : 0];
    _zz_1138 <= _zz_12115[15 : 0];
    _zz_1105 <= _zz_12119[15 : 0];
    _zz_1106 <= _zz_12123[15 : 0];
    _zz_1139 <= _zz_12135[15 : 0];
    _zz_1140 <= _zz_12139[15 : 0];
    _zz_1107 <= _zz_12143[15 : 0];
    _zz_1108 <= _zz_12147[15 : 0];
    _zz_1141 <= _zz_12159[15 : 0];
    _zz_1142 <= _zz_12163[15 : 0];
    _zz_1109 <= _zz_12167[15 : 0];
    _zz_1110 <= _zz_12171[15 : 0];
    _zz_1143 <= _zz_12183[15 : 0];
    _zz_1144 <= _zz_12187[15 : 0];
    _zz_1111 <= _zz_12191[15 : 0];
    _zz_1112 <= _zz_12195[15 : 0];
    _zz_1145 <= _zz_12207[15 : 0];
    _zz_1146 <= _zz_12211[15 : 0];
    _zz_1113 <= _zz_12215[15 : 0];
    _zz_1114 <= _zz_12219[15 : 0];
    _zz_1147 <= _zz_12231[15 : 0];
    _zz_1148 <= _zz_12235[15 : 0];
    _zz_1115 <= _zz_12239[15 : 0];
    _zz_1116 <= _zz_12243[15 : 0];
    _zz_1149 <= _zz_12255[15 : 0];
    _zz_1150 <= _zz_12259[15 : 0];
    _zz_1117 <= _zz_12263[15 : 0];
    _zz_1118 <= _zz_12267[15 : 0];
    _zz_1151 <= _zz_12279[15 : 0];
    _zz_1152 <= _zz_12283[15 : 0];
    _zz_1119 <= _zz_12287[15 : 0];
    _zz_1120 <= _zz_12291[15 : 0];
    _zz_1185 <= _zz_12303[15 : 0];
    _zz_1186 <= _zz_12307[15 : 0];
    _zz_1153 <= _zz_12311[15 : 0];
    _zz_1154 <= _zz_12315[15 : 0];
    _zz_1187 <= _zz_12327[15 : 0];
    _zz_1188 <= _zz_12331[15 : 0];
    _zz_1155 <= _zz_12335[15 : 0];
    _zz_1156 <= _zz_12339[15 : 0];
    _zz_1189 <= _zz_12351[15 : 0];
    _zz_1190 <= _zz_12355[15 : 0];
    _zz_1157 <= _zz_12359[15 : 0];
    _zz_1158 <= _zz_12363[15 : 0];
    _zz_1191 <= _zz_12375[15 : 0];
    _zz_1192 <= _zz_12379[15 : 0];
    _zz_1159 <= _zz_12383[15 : 0];
    _zz_1160 <= _zz_12387[15 : 0];
    _zz_1193 <= _zz_12399[15 : 0];
    _zz_1194 <= _zz_12403[15 : 0];
    _zz_1161 <= _zz_12407[15 : 0];
    _zz_1162 <= _zz_12411[15 : 0];
    _zz_1195 <= _zz_12423[15 : 0];
    _zz_1196 <= _zz_12427[15 : 0];
    _zz_1163 <= _zz_12431[15 : 0];
    _zz_1164 <= _zz_12435[15 : 0];
    _zz_1197 <= _zz_12447[15 : 0];
    _zz_1198 <= _zz_12451[15 : 0];
    _zz_1165 <= _zz_12455[15 : 0];
    _zz_1166 <= _zz_12459[15 : 0];
    _zz_1199 <= _zz_12471[15 : 0];
    _zz_1200 <= _zz_12475[15 : 0];
    _zz_1167 <= _zz_12479[15 : 0];
    _zz_1168 <= _zz_12483[15 : 0];
    _zz_1201 <= _zz_12495[15 : 0];
    _zz_1202 <= _zz_12499[15 : 0];
    _zz_1169 <= _zz_12503[15 : 0];
    _zz_1170 <= _zz_12507[15 : 0];
    _zz_1203 <= _zz_12519[15 : 0];
    _zz_1204 <= _zz_12523[15 : 0];
    _zz_1171 <= _zz_12527[15 : 0];
    _zz_1172 <= _zz_12531[15 : 0];
    _zz_1205 <= _zz_12543[15 : 0];
    _zz_1206 <= _zz_12547[15 : 0];
    _zz_1173 <= _zz_12551[15 : 0];
    _zz_1174 <= _zz_12555[15 : 0];
    _zz_1207 <= _zz_12567[15 : 0];
    _zz_1208 <= _zz_12571[15 : 0];
    _zz_1175 <= _zz_12575[15 : 0];
    _zz_1176 <= _zz_12579[15 : 0];
    _zz_1209 <= _zz_12591[15 : 0];
    _zz_1210 <= _zz_12595[15 : 0];
    _zz_1177 <= _zz_12599[15 : 0];
    _zz_1178 <= _zz_12603[15 : 0];
    _zz_1211 <= _zz_12615[15 : 0];
    _zz_1212 <= _zz_12619[15 : 0];
    _zz_1179 <= _zz_12623[15 : 0];
    _zz_1180 <= _zz_12627[15 : 0];
    _zz_1213 <= _zz_12639[15 : 0];
    _zz_1214 <= _zz_12643[15 : 0];
    _zz_1181 <= _zz_12647[15 : 0];
    _zz_1182 <= _zz_12651[15 : 0];
    _zz_1215 <= _zz_12663[15 : 0];
    _zz_1216 <= _zz_12667[15 : 0];
    _zz_1183 <= _zz_12671[15 : 0];
    _zz_1184 <= _zz_12675[15 : 0];
    _zz_1249 <= _zz_12687[15 : 0];
    _zz_1250 <= _zz_12691[15 : 0];
    _zz_1217 <= _zz_12695[15 : 0];
    _zz_1218 <= _zz_12699[15 : 0];
    _zz_1251 <= _zz_12711[15 : 0];
    _zz_1252 <= _zz_12715[15 : 0];
    _zz_1219 <= _zz_12719[15 : 0];
    _zz_1220 <= _zz_12723[15 : 0];
    _zz_1253 <= _zz_12735[15 : 0];
    _zz_1254 <= _zz_12739[15 : 0];
    _zz_1221 <= _zz_12743[15 : 0];
    _zz_1222 <= _zz_12747[15 : 0];
    _zz_1255 <= _zz_12759[15 : 0];
    _zz_1256 <= _zz_12763[15 : 0];
    _zz_1223 <= _zz_12767[15 : 0];
    _zz_1224 <= _zz_12771[15 : 0];
    _zz_1257 <= _zz_12783[15 : 0];
    _zz_1258 <= _zz_12787[15 : 0];
    _zz_1225 <= _zz_12791[15 : 0];
    _zz_1226 <= _zz_12795[15 : 0];
    _zz_1259 <= _zz_12807[15 : 0];
    _zz_1260 <= _zz_12811[15 : 0];
    _zz_1227 <= _zz_12815[15 : 0];
    _zz_1228 <= _zz_12819[15 : 0];
    _zz_1261 <= _zz_12831[15 : 0];
    _zz_1262 <= _zz_12835[15 : 0];
    _zz_1229 <= _zz_12839[15 : 0];
    _zz_1230 <= _zz_12843[15 : 0];
    _zz_1263 <= _zz_12855[15 : 0];
    _zz_1264 <= _zz_12859[15 : 0];
    _zz_1231 <= _zz_12863[15 : 0];
    _zz_1232 <= _zz_12867[15 : 0];
    _zz_1265 <= _zz_12879[15 : 0];
    _zz_1266 <= _zz_12883[15 : 0];
    _zz_1233 <= _zz_12887[15 : 0];
    _zz_1234 <= _zz_12891[15 : 0];
    _zz_1267 <= _zz_12903[15 : 0];
    _zz_1268 <= _zz_12907[15 : 0];
    _zz_1235 <= _zz_12911[15 : 0];
    _zz_1236 <= _zz_12915[15 : 0];
    _zz_1269 <= _zz_12927[15 : 0];
    _zz_1270 <= _zz_12931[15 : 0];
    _zz_1237 <= _zz_12935[15 : 0];
    _zz_1238 <= _zz_12939[15 : 0];
    _zz_1271 <= _zz_12951[15 : 0];
    _zz_1272 <= _zz_12955[15 : 0];
    _zz_1239 <= _zz_12959[15 : 0];
    _zz_1240 <= _zz_12963[15 : 0];
    _zz_1273 <= _zz_12975[15 : 0];
    _zz_1274 <= _zz_12979[15 : 0];
    _zz_1241 <= _zz_12983[15 : 0];
    _zz_1242 <= _zz_12987[15 : 0];
    _zz_1275 <= _zz_12999[15 : 0];
    _zz_1276 <= _zz_13003[15 : 0];
    _zz_1243 <= _zz_13007[15 : 0];
    _zz_1244 <= _zz_13011[15 : 0];
    _zz_1277 <= _zz_13023[15 : 0];
    _zz_1278 <= _zz_13027[15 : 0];
    _zz_1245 <= _zz_13031[15 : 0];
    _zz_1246 <= _zz_13035[15 : 0];
    _zz_1279 <= _zz_13047[15 : 0];
    _zz_1280 <= _zz_13051[15 : 0];
    _zz_1247 <= _zz_13055[15 : 0];
    _zz_1248 <= _zz_13059[15 : 0];
    _zz_1345 <= _zz_13071[15 : 0];
    _zz_1346 <= _zz_13075[15 : 0];
    _zz_1281 <= _zz_13079[15 : 0];
    _zz_1282 <= _zz_13083[15 : 0];
    _zz_1347 <= _zz_13095[15 : 0];
    _zz_1348 <= _zz_13099[15 : 0];
    _zz_1283 <= _zz_13103[15 : 0];
    _zz_1284 <= _zz_13107[15 : 0];
    _zz_1349 <= _zz_13119[15 : 0];
    _zz_1350 <= _zz_13123[15 : 0];
    _zz_1285 <= _zz_13127[15 : 0];
    _zz_1286 <= _zz_13131[15 : 0];
    _zz_1351 <= _zz_13143[15 : 0];
    _zz_1352 <= _zz_13147[15 : 0];
    _zz_1287 <= _zz_13151[15 : 0];
    _zz_1288 <= _zz_13155[15 : 0];
    _zz_1353 <= _zz_13167[15 : 0];
    _zz_1354 <= _zz_13171[15 : 0];
    _zz_1289 <= _zz_13175[15 : 0];
    _zz_1290 <= _zz_13179[15 : 0];
    _zz_1355 <= _zz_13191[15 : 0];
    _zz_1356 <= _zz_13195[15 : 0];
    _zz_1291 <= _zz_13199[15 : 0];
    _zz_1292 <= _zz_13203[15 : 0];
    _zz_1357 <= _zz_13215[15 : 0];
    _zz_1358 <= _zz_13219[15 : 0];
    _zz_1293 <= _zz_13223[15 : 0];
    _zz_1294 <= _zz_13227[15 : 0];
    _zz_1359 <= _zz_13239[15 : 0];
    _zz_1360 <= _zz_13243[15 : 0];
    _zz_1295 <= _zz_13247[15 : 0];
    _zz_1296 <= _zz_13251[15 : 0];
    _zz_1361 <= _zz_13263[15 : 0];
    _zz_1362 <= _zz_13267[15 : 0];
    _zz_1297 <= _zz_13271[15 : 0];
    _zz_1298 <= _zz_13275[15 : 0];
    _zz_1363 <= _zz_13287[15 : 0];
    _zz_1364 <= _zz_13291[15 : 0];
    _zz_1299 <= _zz_13295[15 : 0];
    _zz_1300 <= _zz_13299[15 : 0];
    _zz_1365 <= _zz_13311[15 : 0];
    _zz_1366 <= _zz_13315[15 : 0];
    _zz_1301 <= _zz_13319[15 : 0];
    _zz_1302 <= _zz_13323[15 : 0];
    _zz_1367 <= _zz_13335[15 : 0];
    _zz_1368 <= _zz_13339[15 : 0];
    _zz_1303 <= _zz_13343[15 : 0];
    _zz_1304 <= _zz_13347[15 : 0];
    _zz_1369 <= _zz_13359[15 : 0];
    _zz_1370 <= _zz_13363[15 : 0];
    _zz_1305 <= _zz_13367[15 : 0];
    _zz_1306 <= _zz_13371[15 : 0];
    _zz_1371 <= _zz_13383[15 : 0];
    _zz_1372 <= _zz_13387[15 : 0];
    _zz_1307 <= _zz_13391[15 : 0];
    _zz_1308 <= _zz_13395[15 : 0];
    _zz_1373 <= _zz_13407[15 : 0];
    _zz_1374 <= _zz_13411[15 : 0];
    _zz_1309 <= _zz_13415[15 : 0];
    _zz_1310 <= _zz_13419[15 : 0];
    _zz_1375 <= _zz_13431[15 : 0];
    _zz_1376 <= _zz_13435[15 : 0];
    _zz_1311 <= _zz_13439[15 : 0];
    _zz_1312 <= _zz_13443[15 : 0];
    _zz_1377 <= _zz_13455[15 : 0];
    _zz_1378 <= _zz_13459[15 : 0];
    _zz_1313 <= _zz_13463[15 : 0];
    _zz_1314 <= _zz_13467[15 : 0];
    _zz_1379 <= _zz_13479[15 : 0];
    _zz_1380 <= _zz_13483[15 : 0];
    _zz_1315 <= _zz_13487[15 : 0];
    _zz_1316 <= _zz_13491[15 : 0];
    _zz_1381 <= _zz_13503[15 : 0];
    _zz_1382 <= _zz_13507[15 : 0];
    _zz_1317 <= _zz_13511[15 : 0];
    _zz_1318 <= _zz_13515[15 : 0];
    _zz_1383 <= _zz_13527[15 : 0];
    _zz_1384 <= _zz_13531[15 : 0];
    _zz_1319 <= _zz_13535[15 : 0];
    _zz_1320 <= _zz_13539[15 : 0];
    _zz_1385 <= _zz_13551[15 : 0];
    _zz_1386 <= _zz_13555[15 : 0];
    _zz_1321 <= _zz_13559[15 : 0];
    _zz_1322 <= _zz_13563[15 : 0];
    _zz_1387 <= _zz_13575[15 : 0];
    _zz_1388 <= _zz_13579[15 : 0];
    _zz_1323 <= _zz_13583[15 : 0];
    _zz_1324 <= _zz_13587[15 : 0];
    _zz_1389 <= _zz_13599[15 : 0];
    _zz_1390 <= _zz_13603[15 : 0];
    _zz_1325 <= _zz_13607[15 : 0];
    _zz_1326 <= _zz_13611[15 : 0];
    _zz_1391 <= _zz_13623[15 : 0];
    _zz_1392 <= _zz_13627[15 : 0];
    _zz_1327 <= _zz_13631[15 : 0];
    _zz_1328 <= _zz_13635[15 : 0];
    _zz_1393 <= _zz_13647[15 : 0];
    _zz_1394 <= _zz_13651[15 : 0];
    _zz_1329 <= _zz_13655[15 : 0];
    _zz_1330 <= _zz_13659[15 : 0];
    _zz_1395 <= _zz_13671[15 : 0];
    _zz_1396 <= _zz_13675[15 : 0];
    _zz_1331 <= _zz_13679[15 : 0];
    _zz_1332 <= _zz_13683[15 : 0];
    _zz_1397 <= _zz_13695[15 : 0];
    _zz_1398 <= _zz_13699[15 : 0];
    _zz_1333 <= _zz_13703[15 : 0];
    _zz_1334 <= _zz_13707[15 : 0];
    _zz_1399 <= _zz_13719[15 : 0];
    _zz_1400 <= _zz_13723[15 : 0];
    _zz_1335 <= _zz_13727[15 : 0];
    _zz_1336 <= _zz_13731[15 : 0];
    _zz_1401 <= _zz_13743[15 : 0];
    _zz_1402 <= _zz_13747[15 : 0];
    _zz_1337 <= _zz_13751[15 : 0];
    _zz_1338 <= _zz_13755[15 : 0];
    _zz_1403 <= _zz_13767[15 : 0];
    _zz_1404 <= _zz_13771[15 : 0];
    _zz_1339 <= _zz_13775[15 : 0];
    _zz_1340 <= _zz_13779[15 : 0];
    _zz_1405 <= _zz_13791[15 : 0];
    _zz_1406 <= _zz_13795[15 : 0];
    _zz_1341 <= _zz_13799[15 : 0];
    _zz_1342 <= _zz_13803[15 : 0];
    _zz_1407 <= _zz_13815[15 : 0];
    _zz_1408 <= _zz_13819[15 : 0];
    _zz_1343 <= _zz_13823[15 : 0];
    _zz_1344 <= _zz_13827[15 : 0];
    _zz_1473 <= _zz_13839[15 : 0];
    _zz_1474 <= _zz_13843[15 : 0];
    _zz_1409 <= _zz_13847[15 : 0];
    _zz_1410 <= _zz_13851[15 : 0];
    _zz_1475 <= _zz_13863[15 : 0];
    _zz_1476 <= _zz_13867[15 : 0];
    _zz_1411 <= _zz_13871[15 : 0];
    _zz_1412 <= _zz_13875[15 : 0];
    _zz_1477 <= _zz_13887[15 : 0];
    _zz_1478 <= _zz_13891[15 : 0];
    _zz_1413 <= _zz_13895[15 : 0];
    _zz_1414 <= _zz_13899[15 : 0];
    _zz_1479 <= _zz_13911[15 : 0];
    _zz_1480 <= _zz_13915[15 : 0];
    _zz_1415 <= _zz_13919[15 : 0];
    _zz_1416 <= _zz_13923[15 : 0];
    _zz_1481 <= _zz_13935[15 : 0];
    _zz_1482 <= _zz_13939[15 : 0];
    _zz_1417 <= _zz_13943[15 : 0];
    _zz_1418 <= _zz_13947[15 : 0];
    _zz_1483 <= _zz_13959[15 : 0];
    _zz_1484 <= _zz_13963[15 : 0];
    _zz_1419 <= _zz_13967[15 : 0];
    _zz_1420 <= _zz_13971[15 : 0];
    _zz_1485 <= _zz_13983[15 : 0];
    _zz_1486 <= _zz_13987[15 : 0];
    _zz_1421 <= _zz_13991[15 : 0];
    _zz_1422 <= _zz_13995[15 : 0];
    _zz_1487 <= _zz_14007[15 : 0];
    _zz_1488 <= _zz_14011[15 : 0];
    _zz_1423 <= _zz_14015[15 : 0];
    _zz_1424 <= _zz_14019[15 : 0];
    _zz_1489 <= _zz_14031[15 : 0];
    _zz_1490 <= _zz_14035[15 : 0];
    _zz_1425 <= _zz_14039[15 : 0];
    _zz_1426 <= _zz_14043[15 : 0];
    _zz_1491 <= _zz_14055[15 : 0];
    _zz_1492 <= _zz_14059[15 : 0];
    _zz_1427 <= _zz_14063[15 : 0];
    _zz_1428 <= _zz_14067[15 : 0];
    _zz_1493 <= _zz_14079[15 : 0];
    _zz_1494 <= _zz_14083[15 : 0];
    _zz_1429 <= _zz_14087[15 : 0];
    _zz_1430 <= _zz_14091[15 : 0];
    _zz_1495 <= _zz_14103[15 : 0];
    _zz_1496 <= _zz_14107[15 : 0];
    _zz_1431 <= _zz_14111[15 : 0];
    _zz_1432 <= _zz_14115[15 : 0];
    _zz_1497 <= _zz_14127[15 : 0];
    _zz_1498 <= _zz_14131[15 : 0];
    _zz_1433 <= _zz_14135[15 : 0];
    _zz_1434 <= _zz_14139[15 : 0];
    _zz_1499 <= _zz_14151[15 : 0];
    _zz_1500 <= _zz_14155[15 : 0];
    _zz_1435 <= _zz_14159[15 : 0];
    _zz_1436 <= _zz_14163[15 : 0];
    _zz_1501 <= _zz_14175[15 : 0];
    _zz_1502 <= _zz_14179[15 : 0];
    _zz_1437 <= _zz_14183[15 : 0];
    _zz_1438 <= _zz_14187[15 : 0];
    _zz_1503 <= _zz_14199[15 : 0];
    _zz_1504 <= _zz_14203[15 : 0];
    _zz_1439 <= _zz_14207[15 : 0];
    _zz_1440 <= _zz_14211[15 : 0];
    _zz_1505 <= _zz_14223[15 : 0];
    _zz_1506 <= _zz_14227[15 : 0];
    _zz_1441 <= _zz_14231[15 : 0];
    _zz_1442 <= _zz_14235[15 : 0];
    _zz_1507 <= _zz_14247[15 : 0];
    _zz_1508 <= _zz_14251[15 : 0];
    _zz_1443 <= _zz_14255[15 : 0];
    _zz_1444 <= _zz_14259[15 : 0];
    _zz_1509 <= _zz_14271[15 : 0];
    _zz_1510 <= _zz_14275[15 : 0];
    _zz_1445 <= _zz_14279[15 : 0];
    _zz_1446 <= _zz_14283[15 : 0];
    _zz_1511 <= _zz_14295[15 : 0];
    _zz_1512 <= _zz_14299[15 : 0];
    _zz_1447 <= _zz_14303[15 : 0];
    _zz_1448 <= _zz_14307[15 : 0];
    _zz_1513 <= _zz_14319[15 : 0];
    _zz_1514 <= _zz_14323[15 : 0];
    _zz_1449 <= _zz_14327[15 : 0];
    _zz_1450 <= _zz_14331[15 : 0];
    _zz_1515 <= _zz_14343[15 : 0];
    _zz_1516 <= _zz_14347[15 : 0];
    _zz_1451 <= _zz_14351[15 : 0];
    _zz_1452 <= _zz_14355[15 : 0];
    _zz_1517 <= _zz_14367[15 : 0];
    _zz_1518 <= _zz_14371[15 : 0];
    _zz_1453 <= _zz_14375[15 : 0];
    _zz_1454 <= _zz_14379[15 : 0];
    _zz_1519 <= _zz_14391[15 : 0];
    _zz_1520 <= _zz_14395[15 : 0];
    _zz_1455 <= _zz_14399[15 : 0];
    _zz_1456 <= _zz_14403[15 : 0];
    _zz_1521 <= _zz_14415[15 : 0];
    _zz_1522 <= _zz_14419[15 : 0];
    _zz_1457 <= _zz_14423[15 : 0];
    _zz_1458 <= _zz_14427[15 : 0];
    _zz_1523 <= _zz_14439[15 : 0];
    _zz_1524 <= _zz_14443[15 : 0];
    _zz_1459 <= _zz_14447[15 : 0];
    _zz_1460 <= _zz_14451[15 : 0];
    _zz_1525 <= _zz_14463[15 : 0];
    _zz_1526 <= _zz_14467[15 : 0];
    _zz_1461 <= _zz_14471[15 : 0];
    _zz_1462 <= _zz_14475[15 : 0];
    _zz_1527 <= _zz_14487[15 : 0];
    _zz_1528 <= _zz_14491[15 : 0];
    _zz_1463 <= _zz_14495[15 : 0];
    _zz_1464 <= _zz_14499[15 : 0];
    _zz_1529 <= _zz_14511[15 : 0];
    _zz_1530 <= _zz_14515[15 : 0];
    _zz_1465 <= _zz_14519[15 : 0];
    _zz_1466 <= _zz_14523[15 : 0];
    _zz_1531 <= _zz_14535[15 : 0];
    _zz_1532 <= _zz_14539[15 : 0];
    _zz_1467 <= _zz_14543[15 : 0];
    _zz_1468 <= _zz_14547[15 : 0];
    _zz_1533 <= _zz_14559[15 : 0];
    _zz_1534 <= _zz_14563[15 : 0];
    _zz_1469 <= _zz_14567[15 : 0];
    _zz_1470 <= _zz_14571[15 : 0];
    _zz_1535 <= _zz_14583[15 : 0];
    _zz_1536 <= _zz_14587[15 : 0];
    _zz_1471 <= _zz_14591[15 : 0];
    _zz_1472 <= _zz_14595[15 : 0];
    _zz_1665 <= _zz_14607[15 : 0];
    _zz_1666 <= _zz_14611[15 : 0];
    _zz_1537 <= _zz_14615[15 : 0];
    _zz_1538 <= _zz_14619[15 : 0];
    _zz_1667 <= _zz_14631[15 : 0];
    _zz_1668 <= _zz_14635[15 : 0];
    _zz_1539 <= _zz_14639[15 : 0];
    _zz_1540 <= _zz_14643[15 : 0];
    _zz_1669 <= _zz_14655[15 : 0];
    _zz_1670 <= _zz_14659[15 : 0];
    _zz_1541 <= _zz_14663[15 : 0];
    _zz_1542 <= _zz_14667[15 : 0];
    _zz_1671 <= _zz_14679[15 : 0];
    _zz_1672 <= _zz_14683[15 : 0];
    _zz_1543 <= _zz_14687[15 : 0];
    _zz_1544 <= _zz_14691[15 : 0];
    _zz_1673 <= _zz_14703[15 : 0];
    _zz_1674 <= _zz_14707[15 : 0];
    _zz_1545 <= _zz_14711[15 : 0];
    _zz_1546 <= _zz_14715[15 : 0];
    _zz_1675 <= _zz_14727[15 : 0];
    _zz_1676 <= _zz_14731[15 : 0];
    _zz_1547 <= _zz_14735[15 : 0];
    _zz_1548 <= _zz_14739[15 : 0];
    _zz_1677 <= _zz_14751[15 : 0];
    _zz_1678 <= _zz_14755[15 : 0];
    _zz_1549 <= _zz_14759[15 : 0];
    _zz_1550 <= _zz_14763[15 : 0];
    _zz_1679 <= _zz_14775[15 : 0];
    _zz_1680 <= _zz_14779[15 : 0];
    _zz_1551 <= _zz_14783[15 : 0];
    _zz_1552 <= _zz_14787[15 : 0];
    _zz_1681 <= _zz_14799[15 : 0];
    _zz_1682 <= _zz_14803[15 : 0];
    _zz_1553 <= _zz_14807[15 : 0];
    _zz_1554 <= _zz_14811[15 : 0];
    _zz_1683 <= _zz_14823[15 : 0];
    _zz_1684 <= _zz_14827[15 : 0];
    _zz_1555 <= _zz_14831[15 : 0];
    _zz_1556 <= _zz_14835[15 : 0];
    _zz_1685 <= _zz_14847[15 : 0];
    _zz_1686 <= _zz_14851[15 : 0];
    _zz_1557 <= _zz_14855[15 : 0];
    _zz_1558 <= _zz_14859[15 : 0];
    _zz_1687 <= _zz_14871[15 : 0];
    _zz_1688 <= _zz_14875[15 : 0];
    _zz_1559 <= _zz_14879[15 : 0];
    _zz_1560 <= _zz_14883[15 : 0];
    _zz_1689 <= _zz_14895[15 : 0];
    _zz_1690 <= _zz_14899[15 : 0];
    _zz_1561 <= _zz_14903[15 : 0];
    _zz_1562 <= _zz_14907[15 : 0];
    _zz_1691 <= _zz_14919[15 : 0];
    _zz_1692 <= _zz_14923[15 : 0];
    _zz_1563 <= _zz_14927[15 : 0];
    _zz_1564 <= _zz_14931[15 : 0];
    _zz_1693 <= _zz_14943[15 : 0];
    _zz_1694 <= _zz_14947[15 : 0];
    _zz_1565 <= _zz_14951[15 : 0];
    _zz_1566 <= _zz_14955[15 : 0];
    _zz_1695 <= _zz_14967[15 : 0];
    _zz_1696 <= _zz_14971[15 : 0];
    _zz_1567 <= _zz_14975[15 : 0];
    _zz_1568 <= _zz_14979[15 : 0];
    _zz_1697 <= _zz_14991[15 : 0];
    _zz_1698 <= _zz_14995[15 : 0];
    _zz_1569 <= _zz_14999[15 : 0];
    _zz_1570 <= _zz_15003[15 : 0];
    _zz_1699 <= _zz_15015[15 : 0];
    _zz_1700 <= _zz_15019[15 : 0];
    _zz_1571 <= _zz_15023[15 : 0];
    _zz_1572 <= _zz_15027[15 : 0];
    _zz_1701 <= _zz_15039[15 : 0];
    _zz_1702 <= _zz_15043[15 : 0];
    _zz_1573 <= _zz_15047[15 : 0];
    _zz_1574 <= _zz_15051[15 : 0];
    _zz_1703 <= _zz_15063[15 : 0];
    _zz_1704 <= _zz_15067[15 : 0];
    _zz_1575 <= _zz_15071[15 : 0];
    _zz_1576 <= _zz_15075[15 : 0];
    _zz_1705 <= _zz_15087[15 : 0];
    _zz_1706 <= _zz_15091[15 : 0];
    _zz_1577 <= _zz_15095[15 : 0];
    _zz_1578 <= _zz_15099[15 : 0];
    _zz_1707 <= _zz_15111[15 : 0];
    _zz_1708 <= _zz_15115[15 : 0];
    _zz_1579 <= _zz_15119[15 : 0];
    _zz_1580 <= _zz_15123[15 : 0];
    _zz_1709 <= _zz_15135[15 : 0];
    _zz_1710 <= _zz_15139[15 : 0];
    _zz_1581 <= _zz_15143[15 : 0];
    _zz_1582 <= _zz_15147[15 : 0];
    _zz_1711 <= _zz_15159[15 : 0];
    _zz_1712 <= _zz_15163[15 : 0];
    _zz_1583 <= _zz_15167[15 : 0];
    _zz_1584 <= _zz_15171[15 : 0];
    _zz_1713 <= _zz_15183[15 : 0];
    _zz_1714 <= _zz_15187[15 : 0];
    _zz_1585 <= _zz_15191[15 : 0];
    _zz_1586 <= _zz_15195[15 : 0];
    _zz_1715 <= _zz_15207[15 : 0];
    _zz_1716 <= _zz_15211[15 : 0];
    _zz_1587 <= _zz_15215[15 : 0];
    _zz_1588 <= _zz_15219[15 : 0];
    _zz_1717 <= _zz_15231[15 : 0];
    _zz_1718 <= _zz_15235[15 : 0];
    _zz_1589 <= _zz_15239[15 : 0];
    _zz_1590 <= _zz_15243[15 : 0];
    _zz_1719 <= _zz_15255[15 : 0];
    _zz_1720 <= _zz_15259[15 : 0];
    _zz_1591 <= _zz_15263[15 : 0];
    _zz_1592 <= _zz_15267[15 : 0];
    _zz_1721 <= _zz_15279[15 : 0];
    _zz_1722 <= _zz_15283[15 : 0];
    _zz_1593 <= _zz_15287[15 : 0];
    _zz_1594 <= _zz_15291[15 : 0];
    _zz_1723 <= _zz_15303[15 : 0];
    _zz_1724 <= _zz_15307[15 : 0];
    _zz_1595 <= _zz_15311[15 : 0];
    _zz_1596 <= _zz_15315[15 : 0];
    _zz_1725 <= _zz_15327[15 : 0];
    _zz_1726 <= _zz_15331[15 : 0];
    _zz_1597 <= _zz_15335[15 : 0];
    _zz_1598 <= _zz_15339[15 : 0];
    _zz_1727 <= _zz_15351[15 : 0];
    _zz_1728 <= _zz_15355[15 : 0];
    _zz_1599 <= _zz_15359[15 : 0];
    _zz_1600 <= _zz_15363[15 : 0];
    _zz_1729 <= _zz_15375[15 : 0];
    _zz_1730 <= _zz_15379[15 : 0];
    _zz_1601 <= _zz_15383[15 : 0];
    _zz_1602 <= _zz_15387[15 : 0];
    _zz_1731 <= _zz_15399[15 : 0];
    _zz_1732 <= _zz_15403[15 : 0];
    _zz_1603 <= _zz_15407[15 : 0];
    _zz_1604 <= _zz_15411[15 : 0];
    _zz_1733 <= _zz_15423[15 : 0];
    _zz_1734 <= _zz_15427[15 : 0];
    _zz_1605 <= _zz_15431[15 : 0];
    _zz_1606 <= _zz_15435[15 : 0];
    _zz_1735 <= _zz_15447[15 : 0];
    _zz_1736 <= _zz_15451[15 : 0];
    _zz_1607 <= _zz_15455[15 : 0];
    _zz_1608 <= _zz_15459[15 : 0];
    _zz_1737 <= _zz_15471[15 : 0];
    _zz_1738 <= _zz_15475[15 : 0];
    _zz_1609 <= _zz_15479[15 : 0];
    _zz_1610 <= _zz_15483[15 : 0];
    _zz_1739 <= _zz_15495[15 : 0];
    _zz_1740 <= _zz_15499[15 : 0];
    _zz_1611 <= _zz_15503[15 : 0];
    _zz_1612 <= _zz_15507[15 : 0];
    _zz_1741 <= _zz_15519[15 : 0];
    _zz_1742 <= _zz_15523[15 : 0];
    _zz_1613 <= _zz_15527[15 : 0];
    _zz_1614 <= _zz_15531[15 : 0];
    _zz_1743 <= _zz_15543[15 : 0];
    _zz_1744 <= _zz_15547[15 : 0];
    _zz_1615 <= _zz_15551[15 : 0];
    _zz_1616 <= _zz_15555[15 : 0];
    _zz_1745 <= _zz_15567[15 : 0];
    _zz_1746 <= _zz_15571[15 : 0];
    _zz_1617 <= _zz_15575[15 : 0];
    _zz_1618 <= _zz_15579[15 : 0];
    _zz_1747 <= _zz_15591[15 : 0];
    _zz_1748 <= _zz_15595[15 : 0];
    _zz_1619 <= _zz_15599[15 : 0];
    _zz_1620 <= _zz_15603[15 : 0];
    _zz_1749 <= _zz_15615[15 : 0];
    _zz_1750 <= _zz_15619[15 : 0];
    _zz_1621 <= _zz_15623[15 : 0];
    _zz_1622 <= _zz_15627[15 : 0];
    _zz_1751 <= _zz_15639[15 : 0];
    _zz_1752 <= _zz_15643[15 : 0];
    _zz_1623 <= _zz_15647[15 : 0];
    _zz_1624 <= _zz_15651[15 : 0];
    _zz_1753 <= _zz_15663[15 : 0];
    _zz_1754 <= _zz_15667[15 : 0];
    _zz_1625 <= _zz_15671[15 : 0];
    _zz_1626 <= _zz_15675[15 : 0];
    _zz_1755 <= _zz_15687[15 : 0];
    _zz_1756 <= _zz_15691[15 : 0];
    _zz_1627 <= _zz_15695[15 : 0];
    _zz_1628 <= _zz_15699[15 : 0];
    _zz_1757 <= _zz_15711[15 : 0];
    _zz_1758 <= _zz_15715[15 : 0];
    _zz_1629 <= _zz_15719[15 : 0];
    _zz_1630 <= _zz_15723[15 : 0];
    _zz_1759 <= _zz_15735[15 : 0];
    _zz_1760 <= _zz_15739[15 : 0];
    _zz_1631 <= _zz_15743[15 : 0];
    _zz_1632 <= _zz_15747[15 : 0];
    _zz_1761 <= _zz_15759[15 : 0];
    _zz_1762 <= _zz_15763[15 : 0];
    _zz_1633 <= _zz_15767[15 : 0];
    _zz_1634 <= _zz_15771[15 : 0];
    _zz_1763 <= _zz_15783[15 : 0];
    _zz_1764 <= _zz_15787[15 : 0];
    _zz_1635 <= _zz_15791[15 : 0];
    _zz_1636 <= _zz_15795[15 : 0];
    _zz_1765 <= _zz_15807[15 : 0];
    _zz_1766 <= _zz_15811[15 : 0];
    _zz_1637 <= _zz_15815[15 : 0];
    _zz_1638 <= _zz_15819[15 : 0];
    _zz_1767 <= _zz_15831[15 : 0];
    _zz_1768 <= _zz_15835[15 : 0];
    _zz_1639 <= _zz_15839[15 : 0];
    _zz_1640 <= _zz_15843[15 : 0];
    _zz_1769 <= _zz_15855[15 : 0];
    _zz_1770 <= _zz_15859[15 : 0];
    _zz_1641 <= _zz_15863[15 : 0];
    _zz_1642 <= _zz_15867[15 : 0];
    _zz_1771 <= _zz_15879[15 : 0];
    _zz_1772 <= _zz_15883[15 : 0];
    _zz_1643 <= _zz_15887[15 : 0];
    _zz_1644 <= _zz_15891[15 : 0];
    _zz_1773 <= _zz_15903[15 : 0];
    _zz_1774 <= _zz_15907[15 : 0];
    _zz_1645 <= _zz_15911[15 : 0];
    _zz_1646 <= _zz_15915[15 : 0];
    _zz_1775 <= _zz_15927[15 : 0];
    _zz_1776 <= _zz_15931[15 : 0];
    _zz_1647 <= _zz_15935[15 : 0];
    _zz_1648 <= _zz_15939[15 : 0];
    _zz_1777 <= _zz_15951[15 : 0];
    _zz_1778 <= _zz_15955[15 : 0];
    _zz_1649 <= _zz_15959[15 : 0];
    _zz_1650 <= _zz_15963[15 : 0];
    _zz_1779 <= _zz_15975[15 : 0];
    _zz_1780 <= _zz_15979[15 : 0];
    _zz_1651 <= _zz_15983[15 : 0];
    _zz_1652 <= _zz_15987[15 : 0];
    _zz_1781 <= _zz_15999[15 : 0];
    _zz_1782 <= _zz_16003[15 : 0];
    _zz_1653 <= _zz_16007[15 : 0];
    _zz_1654 <= _zz_16011[15 : 0];
    _zz_1783 <= _zz_16023[15 : 0];
    _zz_1784 <= _zz_16027[15 : 0];
    _zz_1655 <= _zz_16031[15 : 0];
    _zz_1656 <= _zz_16035[15 : 0];
    _zz_1785 <= _zz_16047[15 : 0];
    _zz_1786 <= _zz_16051[15 : 0];
    _zz_1657 <= _zz_16055[15 : 0];
    _zz_1658 <= _zz_16059[15 : 0];
    _zz_1787 <= _zz_16071[15 : 0];
    _zz_1788 <= _zz_16075[15 : 0];
    _zz_1659 <= _zz_16079[15 : 0];
    _zz_1660 <= _zz_16083[15 : 0];
    _zz_1789 <= _zz_16095[15 : 0];
    _zz_1790 <= _zz_16099[15 : 0];
    _zz_1661 <= _zz_16103[15 : 0];
    _zz_1662 <= _zz_16107[15 : 0];
    _zz_1791 <= _zz_16119[15 : 0];
    _zz_1792 <= _zz_16123[15 : 0];
    _zz_1663 <= _zz_16127[15 : 0];
    _zz_1664 <= _zz_16131[15 : 0];
    io_data_in_valid_regNext <= io_data_in_valid;
  end

  always @ (posedge clk or posedge reset) begin
    if (reset) begin
      _zz_4035 <= 4'b0000;
      _zz_4038 <= 1'b0;
    end else begin
      _zz_4035 <= _zz_4034;
      if(io_data_in_valid_regNext)begin
        _zz_4038 <= 1'b1;
      end else begin
        if(_zz_4037)begin
          _zz_4038 <= 1'b0;
        end
      end
    end
  end


endmodule

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

module SInt32fixTo23_8_ROUNDTOINF (
  input      [31:0]   din,
  output     [15:0]   dout
);
  wire       [32:0]   _zz_9;
  wire       [32:0]   _zz_10;
  wire       [7:0]    _zz_11;
  wire       [24:0]   _zz_12;
  wire       [24:0]   _zz_13;
  wire       [32:0]   _zz_14;
  wire       [32:0]   _zz_15;
  wire       [32:0]   _zz_16;
  wire       [9:0]    _zz_17;
  wire       [8:0]    _zz_18;
  reg        [24:0]   _zz_1;
  wire       [31:0]   _zz_2;
  wire       [31:0]   _zz_3;
  wire       [31:0]   _zz_4;
  wire       [32:0]   _zz_5;
  wire       [31:0]   _zz_6;
  reg        [24:0]   _zz_7;
  reg        [15:0]   _zz_8;

  assign _zz_9 = {_zz_4[31],_zz_4};
  assign _zz_10 = {_zz_3[31],_zz_3};
  assign _zz_11 = _zz_5[7 : 0];
  assign _zz_12 = _zz_5[32 : 8];
  assign _zz_13 = 25'h0000001;
  assign _zz_14 = ($signed(_zz_15) + $signed(_zz_16));
  assign _zz_15 = {_zz_6[31],_zz_6};
  assign _zz_16 = {_zz_2[31],_zz_2};
  assign _zz_17 = _zz_1[24 : 15];
  assign _zz_18 = _zz_1[23 : 15];
  assign _zz_2 = {{24'h0,1'b1},7'h0};
  assign _zz_3 = {25'h1ffffff,7'h0};
  assign _zz_4 = din[31 : 0];
  assign _zz_5 = ($signed(_zz_9) + $signed(_zz_10));
  assign _zz_6 = din[31 : 0];
  always @ (*) begin
    if((_zz_11 != 8'h0))begin
      _zz_7 = ($signed(_zz_12) + $signed(_zz_13));
    end else begin
      _zz_7 = _zz_5[32 : 8];
    end
  end

  always @ (*) begin
    if(_zz_5[32])begin
      _zz_1 = _zz_7;
    end else begin
      _zz_1 = (_zz_14 >>> 8);
    end
  end

  always @ (*) begin
    if(_zz_1[24])begin
      if((! (_zz_17 == 10'h3ff)))begin
        _zz_8 = 16'h8000;
      end else begin
        _zz_8 = _zz_1[15 : 0];
      end
    end else begin
      if((_zz_18 != 9'h0))begin
        _zz_8 = 16'h7fff;
      end else begin
        _zz_8 = _zz_1[15 : 0];
      end
    end
  end

  assign dout = _zz_8;

endmodule
