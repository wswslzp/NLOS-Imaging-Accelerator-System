// Generator : SpinalHDL v1.4.1    git head : d1b4746673438bc5f242515335278fa39a666c38
// Component : SFFT
// Git hash  : ef30208e6bb081eaf187cc4ad996c905dde29f11



module SFFT (
  input               data_in_valid,
  input      [15:0]   data_in_payload_real,
  input      [15:0]   data_in_payload_imag,
  output              data_out_valid,
  output     [15:0]   data_out_payload_real,
  output     [15:0]   data_out_payload_imag,
  input               clk,
  input               reset
);
  reg        [15:0]   _zz_65;
  reg        [15:0]   _zz_66;
  wire                myFFT_1_sdata_out_valid;
  wire       [15:0]   myFFT_1_sdata_out_payload_0_real;
  wire       [15:0]   myFFT_1_sdata_out_payload_0_imag;
  wire       [15:0]   myFFT_1_sdata_out_payload_1_real;
  wire       [15:0]   myFFT_1_sdata_out_payload_1_imag;
  wire       [15:0]   myFFT_1_sdata_out_payload_2_real;
  wire       [15:0]   myFFT_1_sdata_out_payload_2_imag;
  wire       [15:0]   myFFT_1_sdata_out_payload_3_real;
  wire       [15:0]   myFFT_1_sdata_out_payload_3_imag;
  wire       [15:0]   myFFT_1_sdata_out_payload_4_real;
  wire       [15:0]   myFFT_1_sdata_out_payload_4_imag;
  wire       [15:0]   myFFT_1_sdata_out_payload_5_real;
  wire       [15:0]   myFFT_1_sdata_out_payload_5_imag;
  wire       [15:0]   myFFT_1_sdata_out_payload_6_real;
  wire       [15:0]   myFFT_1_sdata_out_payload_6_imag;
  wire       [15:0]   myFFT_1_sdata_out_payload_7_real;
  wire       [15:0]   myFFT_1_sdata_out_payload_7_imag;
  wire       [15:0]   myFFT_1_sdata_out_payload_8_real;
  wire       [15:0]   myFFT_1_sdata_out_payload_8_imag;
  wire       [15:0]   myFFT_1_sdata_out_payload_9_real;
  wire       [15:0]   myFFT_1_sdata_out_payload_9_imag;
  wire       [15:0]   myFFT_1_sdata_out_payload_10_real;
  wire       [15:0]   myFFT_1_sdata_out_payload_10_imag;
  wire       [15:0]   myFFT_1_sdata_out_payload_11_real;
  wire       [15:0]   myFFT_1_sdata_out_payload_11_imag;
  wire       [15:0]   myFFT_1_sdata_out_payload_12_real;
  wire       [15:0]   myFFT_1_sdata_out_payload_12_imag;
  wire       [15:0]   myFFT_1_sdata_out_payload_13_real;
  wire       [15:0]   myFFT_1_sdata_out_payload_13_imag;
  wire       [15:0]   myFFT_1_sdata_out_payload_14_real;
  wire       [15:0]   myFFT_1_sdata_out_payload_14_imag;
  wire       [15:0]   myFFT_1_sdata_out_payload_15_real;
  wire       [15:0]   myFFT_1_sdata_out_payload_15_imag;
  wire       [15:0]   myFFT_1_sdata_out_payload_16_real;
  wire       [15:0]   myFFT_1_sdata_out_payload_16_imag;
  wire       [15:0]   myFFT_1_sdata_out_payload_17_real;
  wire       [15:0]   myFFT_1_sdata_out_payload_17_imag;
  wire       [15:0]   myFFT_1_sdata_out_payload_18_real;
  wire       [15:0]   myFFT_1_sdata_out_payload_18_imag;
  wire       [15:0]   myFFT_1_sdata_out_payload_19_real;
  wire       [15:0]   myFFT_1_sdata_out_payload_19_imag;
  wire       [15:0]   myFFT_1_sdata_out_payload_20_real;
  wire       [15:0]   myFFT_1_sdata_out_payload_20_imag;
  wire       [15:0]   myFFT_1_sdata_out_payload_21_real;
  wire       [15:0]   myFFT_1_sdata_out_payload_21_imag;
  wire       [15:0]   myFFT_1_sdata_out_payload_22_real;
  wire       [15:0]   myFFT_1_sdata_out_payload_22_imag;
  wire       [15:0]   myFFT_1_sdata_out_payload_23_real;
  wire       [15:0]   myFFT_1_sdata_out_payload_23_imag;
  wire       [15:0]   myFFT_1_sdata_out_payload_24_real;
  wire       [15:0]   myFFT_1_sdata_out_payload_24_imag;
  wire       [15:0]   myFFT_1_sdata_out_payload_25_real;
  wire       [15:0]   myFFT_1_sdata_out_payload_25_imag;
  wire       [15:0]   myFFT_1_sdata_out_payload_26_real;
  wire       [15:0]   myFFT_1_sdata_out_payload_26_imag;
  wire       [15:0]   myFFT_1_sdata_out_payload_27_real;
  wire       [15:0]   myFFT_1_sdata_out_payload_27_imag;
  wire       [15:0]   myFFT_1_sdata_out_payload_28_real;
  wire       [15:0]   myFFT_1_sdata_out_payload_28_imag;
  wire       [15:0]   myFFT_1_sdata_out_payload_29_real;
  wire       [15:0]   myFFT_1_sdata_out_payload_29_imag;
  wire       [15:0]   myFFT_1_sdata_out_payload_30_real;
  wire       [15:0]   myFFT_1_sdata_out_payload_30_imag;
  wire       [15:0]   myFFT_1_sdata_out_payload_31_real;
  wire       [15:0]   myFFT_1_sdata_out_payload_31_imag;
  wire       [0:0]    _zz_67;
  wire       [4:0]    _zz_68;
  wire       [0:0]    _zz_69;
  wire       [4:0]    _zz_70;
  wire       [15:0]   _zz_1;
  wire       [15:0]   _zz_2;
  reg        [15:0]   _zz_3;
  reg        [15:0]   _zz_4;
  reg        [15:0]   _zz_5;
  reg        [15:0]   _zz_6;
  reg        [15:0]   _zz_7;
  reg        [15:0]   _zz_8;
  reg        [15:0]   _zz_9;
  reg        [15:0]   _zz_10;
  reg        [15:0]   _zz_11;
  reg        [15:0]   _zz_12;
  reg        [15:0]   _zz_13;
  reg        [15:0]   _zz_14;
  reg        [15:0]   _zz_15;
  reg        [15:0]   _zz_16;
  reg        [15:0]   _zz_17;
  reg        [15:0]   _zz_18;
  reg        [15:0]   _zz_19;
  reg        [15:0]   _zz_20;
  reg        [15:0]   _zz_21;
  reg        [15:0]   _zz_22;
  reg        [15:0]   _zz_23;
  reg        [15:0]   _zz_24;
  reg        [15:0]   _zz_25;
  reg        [15:0]   _zz_26;
  reg        [15:0]   _zz_27;
  reg        [15:0]   _zz_28;
  reg        [15:0]   _zz_29;
  reg        [15:0]   _zz_30;
  reg        [15:0]   _zz_31;
  reg        [15:0]   _zz_32;
  reg        [15:0]   _zz_33;
  reg        [15:0]   _zz_34;
  reg        [15:0]   _zz_35;
  reg        [15:0]   _zz_36;
  reg        [15:0]   _zz_37;
  reg        [15:0]   _zz_38;
  reg        [15:0]   _zz_39;
  reg        [15:0]   _zz_40;
  reg        [15:0]   _zz_41;
  reg        [15:0]   _zz_42;
  reg        [15:0]   _zz_43;
  reg        [15:0]   _zz_44;
  reg        [15:0]   _zz_45;
  reg        [15:0]   _zz_46;
  reg        [15:0]   _zz_47;
  reg        [15:0]   _zz_48;
  reg        [15:0]   _zz_49;
  reg        [15:0]   _zz_50;
  reg        [15:0]   _zz_51;
  reg        [15:0]   _zz_52;
  reg        [15:0]   _zz_53;
  reg        [15:0]   _zz_54;
  reg        [15:0]   _zz_55;
  reg        [15:0]   _zz_56;
  reg        [15:0]   _zz_57;
  reg        [15:0]   _zz_58;
  reg        [15:0]   _zz_59;
  reg        [15:0]   _zz_60;
  reg        [15:0]   _zz_61;
  reg        [15:0]   _zz_62;
  reg        [15:0]   _zz_63;
  reg        [15:0]   _zz_64;
  wire                fft_input_flow_valid;
  wire       [15:0]   fft_input_flow_payload_0_real;
  wire       [15:0]   fft_input_flow_payload_0_imag;
  wire       [15:0]   fft_input_flow_payload_1_real;
  wire       [15:0]   fft_input_flow_payload_1_imag;
  wire       [15:0]   fft_input_flow_payload_2_real;
  wire       [15:0]   fft_input_flow_payload_2_imag;
  wire       [15:0]   fft_input_flow_payload_3_real;
  wire       [15:0]   fft_input_flow_payload_3_imag;
  wire       [15:0]   fft_input_flow_payload_4_real;
  wire       [15:0]   fft_input_flow_payload_4_imag;
  wire       [15:0]   fft_input_flow_payload_5_real;
  wire       [15:0]   fft_input_flow_payload_5_imag;
  wire       [15:0]   fft_input_flow_payload_6_real;
  wire       [15:0]   fft_input_flow_payload_6_imag;
  wire       [15:0]   fft_input_flow_payload_7_real;
  wire       [15:0]   fft_input_flow_payload_7_imag;
  wire       [15:0]   fft_input_flow_payload_8_real;
  wire       [15:0]   fft_input_flow_payload_8_imag;
  wire       [15:0]   fft_input_flow_payload_9_real;
  wire       [15:0]   fft_input_flow_payload_9_imag;
  wire       [15:0]   fft_input_flow_payload_10_real;
  wire       [15:0]   fft_input_flow_payload_10_imag;
  wire       [15:0]   fft_input_flow_payload_11_real;
  wire       [15:0]   fft_input_flow_payload_11_imag;
  wire       [15:0]   fft_input_flow_payload_12_real;
  wire       [15:0]   fft_input_flow_payload_12_imag;
  wire       [15:0]   fft_input_flow_payload_13_real;
  wire       [15:0]   fft_input_flow_payload_13_imag;
  wire       [15:0]   fft_input_flow_payload_14_real;
  wire       [15:0]   fft_input_flow_payload_14_imag;
  wire       [15:0]   fft_input_flow_payload_15_real;
  wire       [15:0]   fft_input_flow_payload_15_imag;
  wire       [15:0]   fft_input_flow_payload_16_real;
  wire       [15:0]   fft_input_flow_payload_16_imag;
  wire       [15:0]   fft_input_flow_payload_17_real;
  wire       [15:0]   fft_input_flow_payload_17_imag;
  wire       [15:0]   fft_input_flow_payload_18_real;
  wire       [15:0]   fft_input_flow_payload_18_imag;
  wire       [15:0]   fft_input_flow_payload_19_real;
  wire       [15:0]   fft_input_flow_payload_19_imag;
  wire       [15:0]   fft_input_flow_payload_20_real;
  wire       [15:0]   fft_input_flow_payload_20_imag;
  wire       [15:0]   fft_input_flow_payload_21_real;
  wire       [15:0]   fft_input_flow_payload_21_imag;
  wire       [15:0]   fft_input_flow_payload_22_real;
  wire       [15:0]   fft_input_flow_payload_22_imag;
  wire       [15:0]   fft_input_flow_payload_23_real;
  wire       [15:0]   fft_input_flow_payload_23_imag;
  wire       [15:0]   fft_input_flow_payload_24_real;
  wire       [15:0]   fft_input_flow_payload_24_imag;
  wire       [15:0]   fft_input_flow_payload_25_real;
  wire       [15:0]   fft_input_flow_payload_25_imag;
  wire       [15:0]   fft_input_flow_payload_26_real;
  wire       [15:0]   fft_input_flow_payload_26_imag;
  wire       [15:0]   fft_input_flow_payload_27_real;
  wire       [15:0]   fft_input_flow_payload_27_imag;
  wire       [15:0]   fft_input_flow_payload_28_real;
  wire       [15:0]   fft_input_flow_payload_28_imag;
  wire       [15:0]   fft_input_flow_payload_29_real;
  wire       [15:0]   fft_input_flow_payload_29_imag;
  wire       [15:0]   fft_input_flow_payload_30_real;
  wire       [15:0]   fft_input_flow_payload_30_imag;
  wire       [15:0]   fft_input_flow_payload_31_real;
  wire       [15:0]   fft_input_flow_payload_31_imag;
  reg                 count_up_inside_cnt_willIncrement;
  wire                count_up_inside_cnt_willClear;
  reg        [4:0]    count_up_inside_cnt_valueNext;
  reg        [4:0]    count_up_inside_cnt_value;
  wire                count_up_inside_cnt_willOverflowIfInc;
  wire                count_up_inside_cnt_willOverflow;
  reg                 myFFT_1_sdata_out_valid_regNext;
  reg                 null_cnt_willIncrement;
  wire                null_cnt_willClear;
  reg        [4:0]    null_cnt_valueNext;
  reg        [4:0]    null_cnt_value;
  wire                null_cnt_willOverflowIfInc;
  wire                null_cnt_willOverflow;
  reg                 null_cond_period_minus_1;
  wire                null_cond_period;
  reg        [15:0]   sdata_out_regs_0_real;
  reg        [15:0]   sdata_out_regs_0_imag;
  reg        [15:0]   sdata_out_regs_1_real;
  reg        [15:0]   sdata_out_regs_1_imag;
  reg        [15:0]   sdata_out_regs_2_real;
  reg        [15:0]   sdata_out_regs_2_imag;
  reg        [15:0]   sdata_out_regs_3_real;
  reg        [15:0]   sdata_out_regs_3_imag;
  reg        [15:0]   sdata_out_regs_4_real;
  reg        [15:0]   sdata_out_regs_4_imag;
  reg        [15:0]   sdata_out_regs_5_real;
  reg        [15:0]   sdata_out_regs_5_imag;
  reg        [15:0]   sdata_out_regs_6_real;
  reg        [15:0]   sdata_out_regs_6_imag;
  reg        [15:0]   sdata_out_regs_7_real;
  reg        [15:0]   sdata_out_regs_7_imag;
  reg        [15:0]   sdata_out_regs_8_real;
  reg        [15:0]   sdata_out_regs_8_imag;
  reg        [15:0]   sdata_out_regs_9_real;
  reg        [15:0]   sdata_out_regs_9_imag;
  reg        [15:0]   sdata_out_regs_10_real;
  reg        [15:0]   sdata_out_regs_10_imag;
  reg        [15:0]   sdata_out_regs_11_real;
  reg        [15:0]   sdata_out_regs_11_imag;
  reg        [15:0]   sdata_out_regs_12_real;
  reg        [15:0]   sdata_out_regs_12_imag;
  reg        [15:0]   sdata_out_regs_13_real;
  reg        [15:0]   sdata_out_regs_13_imag;
  reg        [15:0]   sdata_out_regs_14_real;
  reg        [15:0]   sdata_out_regs_14_imag;
  reg        [15:0]   sdata_out_regs_15_real;
  reg        [15:0]   sdata_out_regs_15_imag;
  reg        [15:0]   sdata_out_regs_16_real;
  reg        [15:0]   sdata_out_regs_16_imag;
  reg        [15:0]   sdata_out_regs_17_real;
  reg        [15:0]   sdata_out_regs_17_imag;
  reg        [15:0]   sdata_out_regs_18_real;
  reg        [15:0]   sdata_out_regs_18_imag;
  reg        [15:0]   sdata_out_regs_19_real;
  reg        [15:0]   sdata_out_regs_19_imag;
  reg        [15:0]   sdata_out_regs_20_real;
  reg        [15:0]   sdata_out_regs_20_imag;
  reg        [15:0]   sdata_out_regs_21_real;
  reg        [15:0]   sdata_out_regs_21_imag;
  reg        [15:0]   sdata_out_regs_22_real;
  reg        [15:0]   sdata_out_regs_22_imag;
  reg        [15:0]   sdata_out_regs_23_real;
  reg        [15:0]   sdata_out_regs_23_imag;
  reg        [15:0]   sdata_out_regs_24_real;
  reg        [15:0]   sdata_out_regs_24_imag;
  reg        [15:0]   sdata_out_regs_25_real;
  reg        [15:0]   sdata_out_regs_25_imag;
  reg        [15:0]   sdata_out_regs_26_real;
  reg        [15:0]   sdata_out_regs_26_imag;
  reg        [15:0]   sdata_out_regs_27_real;
  reg        [15:0]   sdata_out_regs_27_imag;
  reg        [15:0]   sdata_out_regs_28_real;
  reg        [15:0]   sdata_out_regs_28_imag;
  reg        [15:0]   sdata_out_regs_29_real;
  reg        [15:0]   sdata_out_regs_29_imag;
  reg        [15:0]   sdata_out_regs_30_real;
  reg        [15:0]   sdata_out_regs_30_imag;
  reg        [15:0]   sdata_out_regs_31_real;
  reg        [15:0]   sdata_out_regs_31_imag;
  wire                output_valid;
  wire       [15:0]   output_payload_real;
  wire       [15:0]   output_payload_imag;

  assign _zz_67 = count_up_inside_cnt_willIncrement;
  assign _zz_68 = {4'd0, _zz_67};
  assign _zz_69 = null_cnt_willIncrement;
  assign _zz_70 = {4'd0, _zz_69};
  MyFFT myFFT_1 (
    .io_data_in_valid              (fft_input_flow_valid                     ), //i
    .io_data_in_payload_0_real     (fft_input_flow_payload_0_real[15:0]      ), //i
    .io_data_in_payload_0_imag     (fft_input_flow_payload_0_imag[15:0]      ), //i
    .io_data_in_payload_1_real     (fft_input_flow_payload_1_real[15:0]      ), //i
    .io_data_in_payload_1_imag     (fft_input_flow_payload_1_imag[15:0]      ), //i
    .io_data_in_payload_2_real     (fft_input_flow_payload_2_real[15:0]      ), //i
    .io_data_in_payload_2_imag     (fft_input_flow_payload_2_imag[15:0]      ), //i
    .io_data_in_payload_3_real     (fft_input_flow_payload_3_real[15:0]      ), //i
    .io_data_in_payload_3_imag     (fft_input_flow_payload_3_imag[15:0]      ), //i
    .io_data_in_payload_4_real     (fft_input_flow_payload_4_real[15:0]      ), //i
    .io_data_in_payload_4_imag     (fft_input_flow_payload_4_imag[15:0]      ), //i
    .io_data_in_payload_5_real     (fft_input_flow_payload_5_real[15:0]      ), //i
    .io_data_in_payload_5_imag     (fft_input_flow_payload_5_imag[15:0]      ), //i
    .io_data_in_payload_6_real     (fft_input_flow_payload_6_real[15:0]      ), //i
    .io_data_in_payload_6_imag     (fft_input_flow_payload_6_imag[15:0]      ), //i
    .io_data_in_payload_7_real     (fft_input_flow_payload_7_real[15:0]      ), //i
    .io_data_in_payload_7_imag     (fft_input_flow_payload_7_imag[15:0]      ), //i
    .io_data_in_payload_8_real     (fft_input_flow_payload_8_real[15:0]      ), //i
    .io_data_in_payload_8_imag     (fft_input_flow_payload_8_imag[15:0]      ), //i
    .io_data_in_payload_9_real     (fft_input_flow_payload_9_real[15:0]      ), //i
    .io_data_in_payload_9_imag     (fft_input_flow_payload_9_imag[15:0]      ), //i
    .io_data_in_payload_10_real    (fft_input_flow_payload_10_real[15:0]     ), //i
    .io_data_in_payload_10_imag    (fft_input_flow_payload_10_imag[15:0]     ), //i
    .io_data_in_payload_11_real    (fft_input_flow_payload_11_real[15:0]     ), //i
    .io_data_in_payload_11_imag    (fft_input_flow_payload_11_imag[15:0]     ), //i
    .io_data_in_payload_12_real    (fft_input_flow_payload_12_real[15:0]     ), //i
    .io_data_in_payload_12_imag    (fft_input_flow_payload_12_imag[15:0]     ), //i
    .io_data_in_payload_13_real    (fft_input_flow_payload_13_real[15:0]     ), //i
    .io_data_in_payload_13_imag    (fft_input_flow_payload_13_imag[15:0]     ), //i
    .io_data_in_payload_14_real    (fft_input_flow_payload_14_real[15:0]     ), //i
    .io_data_in_payload_14_imag    (fft_input_flow_payload_14_imag[15:0]     ), //i
    .io_data_in_payload_15_real    (fft_input_flow_payload_15_real[15:0]     ), //i
    .io_data_in_payload_15_imag    (fft_input_flow_payload_15_imag[15:0]     ), //i
    .io_data_in_payload_16_real    (fft_input_flow_payload_16_real[15:0]     ), //i
    .io_data_in_payload_16_imag    (fft_input_flow_payload_16_imag[15:0]     ), //i
    .io_data_in_payload_17_real    (fft_input_flow_payload_17_real[15:0]     ), //i
    .io_data_in_payload_17_imag    (fft_input_flow_payload_17_imag[15:0]     ), //i
    .io_data_in_payload_18_real    (fft_input_flow_payload_18_real[15:0]     ), //i
    .io_data_in_payload_18_imag    (fft_input_flow_payload_18_imag[15:0]     ), //i
    .io_data_in_payload_19_real    (fft_input_flow_payload_19_real[15:0]     ), //i
    .io_data_in_payload_19_imag    (fft_input_flow_payload_19_imag[15:0]     ), //i
    .io_data_in_payload_20_real    (fft_input_flow_payload_20_real[15:0]     ), //i
    .io_data_in_payload_20_imag    (fft_input_flow_payload_20_imag[15:0]     ), //i
    .io_data_in_payload_21_real    (fft_input_flow_payload_21_real[15:0]     ), //i
    .io_data_in_payload_21_imag    (fft_input_flow_payload_21_imag[15:0]     ), //i
    .io_data_in_payload_22_real    (fft_input_flow_payload_22_real[15:0]     ), //i
    .io_data_in_payload_22_imag    (fft_input_flow_payload_22_imag[15:0]     ), //i
    .io_data_in_payload_23_real    (fft_input_flow_payload_23_real[15:0]     ), //i
    .io_data_in_payload_23_imag    (fft_input_flow_payload_23_imag[15:0]     ), //i
    .io_data_in_payload_24_real    (fft_input_flow_payload_24_real[15:0]     ), //i
    .io_data_in_payload_24_imag    (fft_input_flow_payload_24_imag[15:0]     ), //i
    .io_data_in_payload_25_real    (fft_input_flow_payload_25_real[15:0]     ), //i
    .io_data_in_payload_25_imag    (fft_input_flow_payload_25_imag[15:0]     ), //i
    .io_data_in_payload_26_real    (fft_input_flow_payload_26_real[15:0]     ), //i
    .io_data_in_payload_26_imag    (fft_input_flow_payload_26_imag[15:0]     ), //i
    .io_data_in_payload_27_real    (fft_input_flow_payload_27_real[15:0]     ), //i
    .io_data_in_payload_27_imag    (fft_input_flow_payload_27_imag[15:0]     ), //i
    .io_data_in_payload_28_real    (fft_input_flow_payload_28_real[15:0]     ), //i
    .io_data_in_payload_28_imag    (fft_input_flow_payload_28_imag[15:0]     ), //i
    .io_data_in_payload_29_real    (fft_input_flow_payload_29_real[15:0]     ), //i
    .io_data_in_payload_29_imag    (fft_input_flow_payload_29_imag[15:0]     ), //i
    .io_data_in_payload_30_real    (fft_input_flow_payload_30_real[15:0]     ), //i
    .io_data_in_payload_30_imag    (fft_input_flow_payload_30_imag[15:0]     ), //i
    .io_data_in_payload_31_real    (fft_input_flow_payload_31_real[15:0]     ), //i
    .io_data_in_payload_31_imag    (fft_input_flow_payload_31_imag[15:0]     ), //i
    .sdata_out_valid               (myFFT_1_sdata_out_valid                  ), //o
    .sdata_out_payload_0_real      (myFFT_1_sdata_out_payload_0_real[15:0]   ), //o
    .sdata_out_payload_0_imag      (myFFT_1_sdata_out_payload_0_imag[15:0]   ), //o
    .sdata_out_payload_1_real      (myFFT_1_sdata_out_payload_1_real[15:0]   ), //o
    .sdata_out_payload_1_imag      (myFFT_1_sdata_out_payload_1_imag[15:0]   ), //o
    .sdata_out_payload_2_real      (myFFT_1_sdata_out_payload_2_real[15:0]   ), //o
    .sdata_out_payload_2_imag      (myFFT_1_sdata_out_payload_2_imag[15:0]   ), //o
    .sdata_out_payload_3_real      (myFFT_1_sdata_out_payload_3_real[15:0]   ), //o
    .sdata_out_payload_3_imag      (myFFT_1_sdata_out_payload_3_imag[15:0]   ), //o
    .sdata_out_payload_4_real      (myFFT_1_sdata_out_payload_4_real[15:0]   ), //o
    .sdata_out_payload_4_imag      (myFFT_1_sdata_out_payload_4_imag[15:0]   ), //o
    .sdata_out_payload_5_real      (myFFT_1_sdata_out_payload_5_real[15:0]   ), //o
    .sdata_out_payload_5_imag      (myFFT_1_sdata_out_payload_5_imag[15:0]   ), //o
    .sdata_out_payload_6_real      (myFFT_1_sdata_out_payload_6_real[15:0]   ), //o
    .sdata_out_payload_6_imag      (myFFT_1_sdata_out_payload_6_imag[15:0]   ), //o
    .sdata_out_payload_7_real      (myFFT_1_sdata_out_payload_7_real[15:0]   ), //o
    .sdata_out_payload_7_imag      (myFFT_1_sdata_out_payload_7_imag[15:0]   ), //o
    .sdata_out_payload_8_real      (myFFT_1_sdata_out_payload_8_real[15:0]   ), //o
    .sdata_out_payload_8_imag      (myFFT_1_sdata_out_payload_8_imag[15:0]   ), //o
    .sdata_out_payload_9_real      (myFFT_1_sdata_out_payload_9_real[15:0]   ), //o
    .sdata_out_payload_9_imag      (myFFT_1_sdata_out_payload_9_imag[15:0]   ), //o
    .sdata_out_payload_10_real     (myFFT_1_sdata_out_payload_10_real[15:0]  ), //o
    .sdata_out_payload_10_imag     (myFFT_1_sdata_out_payload_10_imag[15:0]  ), //o
    .sdata_out_payload_11_real     (myFFT_1_sdata_out_payload_11_real[15:0]  ), //o
    .sdata_out_payload_11_imag     (myFFT_1_sdata_out_payload_11_imag[15:0]  ), //o
    .sdata_out_payload_12_real     (myFFT_1_sdata_out_payload_12_real[15:0]  ), //o
    .sdata_out_payload_12_imag     (myFFT_1_sdata_out_payload_12_imag[15:0]  ), //o
    .sdata_out_payload_13_real     (myFFT_1_sdata_out_payload_13_real[15:0]  ), //o
    .sdata_out_payload_13_imag     (myFFT_1_sdata_out_payload_13_imag[15:0]  ), //o
    .sdata_out_payload_14_real     (myFFT_1_sdata_out_payload_14_real[15:0]  ), //o
    .sdata_out_payload_14_imag     (myFFT_1_sdata_out_payload_14_imag[15:0]  ), //o
    .sdata_out_payload_15_real     (myFFT_1_sdata_out_payload_15_real[15:0]  ), //o
    .sdata_out_payload_15_imag     (myFFT_1_sdata_out_payload_15_imag[15:0]  ), //o
    .sdata_out_payload_16_real     (myFFT_1_sdata_out_payload_16_real[15:0]  ), //o
    .sdata_out_payload_16_imag     (myFFT_1_sdata_out_payload_16_imag[15:0]  ), //o
    .sdata_out_payload_17_real     (myFFT_1_sdata_out_payload_17_real[15:0]  ), //o
    .sdata_out_payload_17_imag     (myFFT_1_sdata_out_payload_17_imag[15:0]  ), //o
    .sdata_out_payload_18_real     (myFFT_1_sdata_out_payload_18_real[15:0]  ), //o
    .sdata_out_payload_18_imag     (myFFT_1_sdata_out_payload_18_imag[15:0]  ), //o
    .sdata_out_payload_19_real     (myFFT_1_sdata_out_payload_19_real[15:0]  ), //o
    .sdata_out_payload_19_imag     (myFFT_1_sdata_out_payload_19_imag[15:0]  ), //o
    .sdata_out_payload_20_real     (myFFT_1_sdata_out_payload_20_real[15:0]  ), //o
    .sdata_out_payload_20_imag     (myFFT_1_sdata_out_payload_20_imag[15:0]  ), //o
    .sdata_out_payload_21_real     (myFFT_1_sdata_out_payload_21_real[15:0]  ), //o
    .sdata_out_payload_21_imag     (myFFT_1_sdata_out_payload_21_imag[15:0]  ), //o
    .sdata_out_payload_22_real     (myFFT_1_sdata_out_payload_22_real[15:0]  ), //o
    .sdata_out_payload_22_imag     (myFFT_1_sdata_out_payload_22_imag[15:0]  ), //o
    .sdata_out_payload_23_real     (myFFT_1_sdata_out_payload_23_real[15:0]  ), //o
    .sdata_out_payload_23_imag     (myFFT_1_sdata_out_payload_23_imag[15:0]  ), //o
    .sdata_out_payload_24_real     (myFFT_1_sdata_out_payload_24_real[15:0]  ), //o
    .sdata_out_payload_24_imag     (myFFT_1_sdata_out_payload_24_imag[15:0]  ), //o
    .sdata_out_payload_25_real     (myFFT_1_sdata_out_payload_25_real[15:0]  ), //o
    .sdata_out_payload_25_imag     (myFFT_1_sdata_out_payload_25_imag[15:0]  ), //o
    .sdata_out_payload_26_real     (myFFT_1_sdata_out_payload_26_real[15:0]  ), //o
    .sdata_out_payload_26_imag     (myFFT_1_sdata_out_payload_26_imag[15:0]  ), //o
    .sdata_out_payload_27_real     (myFFT_1_sdata_out_payload_27_real[15:0]  ), //o
    .sdata_out_payload_27_imag     (myFFT_1_sdata_out_payload_27_imag[15:0]  ), //o
    .sdata_out_payload_28_real     (myFFT_1_sdata_out_payload_28_real[15:0]  ), //o
    .sdata_out_payload_28_imag     (myFFT_1_sdata_out_payload_28_imag[15:0]  ), //o
    .sdata_out_payload_29_real     (myFFT_1_sdata_out_payload_29_real[15:0]  ), //o
    .sdata_out_payload_29_imag     (myFFT_1_sdata_out_payload_29_imag[15:0]  ), //o
    .sdata_out_payload_30_real     (myFFT_1_sdata_out_payload_30_real[15:0]  ), //o
    .sdata_out_payload_30_imag     (myFFT_1_sdata_out_payload_30_imag[15:0]  ), //o
    .sdata_out_payload_31_real     (myFFT_1_sdata_out_payload_31_real[15:0]  ), //o
    .sdata_out_payload_31_imag     (myFFT_1_sdata_out_payload_31_imag[15:0]  ), //o
    .clk                           (clk                                      ), //i
    .reset                         (reset                                    )  //i
  );
  always @(*) begin
    case(null_cnt_value)
      5'b00000 : begin
        _zz_65 = sdata_out_regs_0_real;
        _zz_66 = sdata_out_regs_0_imag;
      end
      5'b00001 : begin
        _zz_65 = sdata_out_regs_1_real;
        _zz_66 = sdata_out_regs_1_imag;
      end
      5'b00010 : begin
        _zz_65 = sdata_out_regs_2_real;
        _zz_66 = sdata_out_regs_2_imag;
      end
      5'b00011 : begin
        _zz_65 = sdata_out_regs_3_real;
        _zz_66 = sdata_out_regs_3_imag;
      end
      5'b00100 : begin
        _zz_65 = sdata_out_regs_4_real;
        _zz_66 = sdata_out_regs_4_imag;
      end
      5'b00101 : begin
        _zz_65 = sdata_out_regs_5_real;
        _zz_66 = sdata_out_regs_5_imag;
      end
      5'b00110 : begin
        _zz_65 = sdata_out_regs_6_real;
        _zz_66 = sdata_out_regs_6_imag;
      end
      5'b00111 : begin
        _zz_65 = sdata_out_regs_7_real;
        _zz_66 = sdata_out_regs_7_imag;
      end
      5'b01000 : begin
        _zz_65 = sdata_out_regs_8_real;
        _zz_66 = sdata_out_regs_8_imag;
      end
      5'b01001 : begin
        _zz_65 = sdata_out_regs_9_real;
        _zz_66 = sdata_out_regs_9_imag;
      end
      5'b01010 : begin
        _zz_65 = sdata_out_regs_10_real;
        _zz_66 = sdata_out_regs_10_imag;
      end
      5'b01011 : begin
        _zz_65 = sdata_out_regs_11_real;
        _zz_66 = sdata_out_regs_11_imag;
      end
      5'b01100 : begin
        _zz_65 = sdata_out_regs_12_real;
        _zz_66 = sdata_out_regs_12_imag;
      end
      5'b01101 : begin
        _zz_65 = sdata_out_regs_13_real;
        _zz_66 = sdata_out_regs_13_imag;
      end
      5'b01110 : begin
        _zz_65 = sdata_out_regs_14_real;
        _zz_66 = sdata_out_regs_14_imag;
      end
      5'b01111 : begin
        _zz_65 = sdata_out_regs_15_real;
        _zz_66 = sdata_out_regs_15_imag;
      end
      5'b10000 : begin
        _zz_65 = sdata_out_regs_16_real;
        _zz_66 = sdata_out_regs_16_imag;
      end
      5'b10001 : begin
        _zz_65 = sdata_out_regs_17_real;
        _zz_66 = sdata_out_regs_17_imag;
      end
      5'b10010 : begin
        _zz_65 = sdata_out_regs_18_real;
        _zz_66 = sdata_out_regs_18_imag;
      end
      5'b10011 : begin
        _zz_65 = sdata_out_regs_19_real;
        _zz_66 = sdata_out_regs_19_imag;
      end
      5'b10100 : begin
        _zz_65 = sdata_out_regs_20_real;
        _zz_66 = sdata_out_regs_20_imag;
      end
      5'b10101 : begin
        _zz_65 = sdata_out_regs_21_real;
        _zz_66 = sdata_out_regs_21_imag;
      end
      5'b10110 : begin
        _zz_65 = sdata_out_regs_22_real;
        _zz_66 = sdata_out_regs_22_imag;
      end
      5'b10111 : begin
        _zz_65 = sdata_out_regs_23_real;
        _zz_66 = sdata_out_regs_23_imag;
      end
      5'b11000 : begin
        _zz_65 = sdata_out_regs_24_real;
        _zz_66 = sdata_out_regs_24_imag;
      end
      5'b11001 : begin
        _zz_65 = sdata_out_regs_25_real;
        _zz_66 = sdata_out_regs_25_imag;
      end
      5'b11010 : begin
        _zz_65 = sdata_out_regs_26_real;
        _zz_66 = sdata_out_regs_26_imag;
      end
      5'b11011 : begin
        _zz_65 = sdata_out_regs_27_real;
        _zz_66 = sdata_out_regs_27_imag;
      end
      5'b11100 : begin
        _zz_65 = sdata_out_regs_28_real;
        _zz_66 = sdata_out_regs_28_imag;
      end
      5'b11101 : begin
        _zz_65 = sdata_out_regs_29_real;
        _zz_66 = sdata_out_regs_29_imag;
      end
      5'b11110 : begin
        _zz_65 = sdata_out_regs_30_real;
        _zz_66 = sdata_out_regs_30_imag;
      end
      default : begin
        _zz_65 = sdata_out_regs_31_real;
        _zz_66 = sdata_out_regs_31_imag;
      end
    endcase
  end

  assign _zz_1 = data_in_payload_real;
  assign _zz_2 = data_in_payload_imag;
  assign fft_input_flow_payload_0_real = _zz_63;
  assign fft_input_flow_payload_0_imag = _zz_64;
  assign fft_input_flow_payload_1_real = _zz_61;
  assign fft_input_flow_payload_1_imag = _zz_62;
  assign fft_input_flow_payload_2_real = _zz_59;
  assign fft_input_flow_payload_2_imag = _zz_60;
  assign fft_input_flow_payload_3_real = _zz_57;
  assign fft_input_flow_payload_3_imag = _zz_58;
  assign fft_input_flow_payload_4_real = _zz_55;
  assign fft_input_flow_payload_4_imag = _zz_56;
  assign fft_input_flow_payload_5_real = _zz_53;
  assign fft_input_flow_payload_5_imag = _zz_54;
  assign fft_input_flow_payload_6_real = _zz_51;
  assign fft_input_flow_payload_6_imag = _zz_52;
  assign fft_input_flow_payload_7_real = _zz_49;
  assign fft_input_flow_payload_7_imag = _zz_50;
  assign fft_input_flow_payload_8_real = _zz_47;
  assign fft_input_flow_payload_8_imag = _zz_48;
  assign fft_input_flow_payload_9_real = _zz_45;
  assign fft_input_flow_payload_9_imag = _zz_46;
  assign fft_input_flow_payload_10_real = _zz_43;
  assign fft_input_flow_payload_10_imag = _zz_44;
  assign fft_input_flow_payload_11_real = _zz_41;
  assign fft_input_flow_payload_11_imag = _zz_42;
  assign fft_input_flow_payload_12_real = _zz_39;
  assign fft_input_flow_payload_12_imag = _zz_40;
  assign fft_input_flow_payload_13_real = _zz_37;
  assign fft_input_flow_payload_13_imag = _zz_38;
  assign fft_input_flow_payload_14_real = _zz_35;
  assign fft_input_flow_payload_14_imag = _zz_36;
  assign fft_input_flow_payload_15_real = _zz_33;
  assign fft_input_flow_payload_15_imag = _zz_34;
  assign fft_input_flow_payload_16_real = _zz_31;
  assign fft_input_flow_payload_16_imag = _zz_32;
  assign fft_input_flow_payload_17_real = _zz_29;
  assign fft_input_flow_payload_17_imag = _zz_30;
  assign fft_input_flow_payload_18_real = _zz_27;
  assign fft_input_flow_payload_18_imag = _zz_28;
  assign fft_input_flow_payload_19_real = _zz_25;
  assign fft_input_flow_payload_19_imag = _zz_26;
  assign fft_input_flow_payload_20_real = _zz_23;
  assign fft_input_flow_payload_20_imag = _zz_24;
  assign fft_input_flow_payload_21_real = _zz_21;
  assign fft_input_flow_payload_21_imag = _zz_22;
  assign fft_input_flow_payload_22_real = _zz_19;
  assign fft_input_flow_payload_22_imag = _zz_20;
  assign fft_input_flow_payload_23_real = _zz_17;
  assign fft_input_flow_payload_23_imag = _zz_18;
  assign fft_input_flow_payload_24_real = _zz_15;
  assign fft_input_flow_payload_24_imag = _zz_16;
  assign fft_input_flow_payload_25_real = _zz_13;
  assign fft_input_flow_payload_25_imag = _zz_14;
  assign fft_input_flow_payload_26_real = _zz_11;
  assign fft_input_flow_payload_26_imag = _zz_12;
  assign fft_input_flow_payload_27_real = _zz_9;
  assign fft_input_flow_payload_27_imag = _zz_10;
  assign fft_input_flow_payload_28_real = _zz_7;
  assign fft_input_flow_payload_28_imag = _zz_8;
  assign fft_input_flow_payload_29_real = _zz_5;
  assign fft_input_flow_payload_29_imag = _zz_6;
  assign fft_input_flow_payload_30_real = _zz_3;
  assign fft_input_flow_payload_30_imag = _zz_4;
  assign fft_input_flow_payload_31_real = _zz_1;
  assign fft_input_flow_payload_31_imag = _zz_2;
  always @ (*) begin
    count_up_inside_cnt_willIncrement = 1'b0;
    if(data_in_valid)begin
      count_up_inside_cnt_willIncrement = 1'b1;
    end
  end

  assign count_up_inside_cnt_willClear = 1'b0;
  assign count_up_inside_cnt_willOverflowIfInc = (count_up_inside_cnt_value == 5'h1f);
  assign count_up_inside_cnt_willOverflow = (count_up_inside_cnt_willOverflowIfInc && count_up_inside_cnt_willIncrement);
  always @ (*) begin
    count_up_inside_cnt_valueNext = (count_up_inside_cnt_value + _zz_68);
    if(count_up_inside_cnt_willClear)begin
      count_up_inside_cnt_valueNext = 5'h0;
    end
  end

  assign fft_input_flow_valid = count_up_inside_cnt_willOverflow;
  always @ (*) begin
    null_cnt_willIncrement = 1'b0;
    if(null_cond_period)begin
      null_cnt_willIncrement = 1'b1;
    end
  end

  assign null_cnt_willClear = 1'b0;
  assign null_cnt_willOverflowIfInc = (null_cnt_value == 5'h1f);
  assign null_cnt_willOverflow = (null_cnt_willOverflowIfInc && null_cnt_willIncrement);
  always @ (*) begin
    null_cnt_valueNext = (null_cnt_value + _zz_70);
    if(null_cnt_willClear)begin
      null_cnt_valueNext = 5'h0;
    end
  end

  assign null_cond_period = (myFFT_1_sdata_out_valid_regNext || null_cond_period_minus_1);
  assign output_payload_real = _zz_65;
  assign output_payload_imag = _zz_66;
  assign output_valid = null_cond_period;
  assign data_out_valid = output_valid;
  assign data_out_payload_real = output_payload_real;
  assign data_out_payload_imag = output_payload_imag;
  always @ (posedge clk) begin
    if(data_in_valid)begin
      _zz_3 <= _zz_1;
      _zz_4 <= _zz_2;
    end
    if(data_in_valid)begin
      _zz_5 <= _zz_3;
      _zz_6 <= _zz_4;
    end
    if(data_in_valid)begin
      _zz_7 <= _zz_5;
      _zz_8 <= _zz_6;
    end
    if(data_in_valid)begin
      _zz_9 <= _zz_7;
      _zz_10 <= _zz_8;
    end
    if(data_in_valid)begin
      _zz_11 <= _zz_9;
      _zz_12 <= _zz_10;
    end
    if(data_in_valid)begin
      _zz_13 <= _zz_11;
      _zz_14 <= _zz_12;
    end
    if(data_in_valid)begin
      _zz_15 <= _zz_13;
      _zz_16 <= _zz_14;
    end
    if(data_in_valid)begin
      _zz_17 <= _zz_15;
      _zz_18 <= _zz_16;
    end
    if(data_in_valid)begin
      _zz_19 <= _zz_17;
      _zz_20 <= _zz_18;
    end
    if(data_in_valid)begin
      _zz_21 <= _zz_19;
      _zz_22 <= _zz_20;
    end
    if(data_in_valid)begin
      _zz_23 <= _zz_21;
      _zz_24 <= _zz_22;
    end
    if(data_in_valid)begin
      _zz_25 <= _zz_23;
      _zz_26 <= _zz_24;
    end
    if(data_in_valid)begin
      _zz_27 <= _zz_25;
      _zz_28 <= _zz_26;
    end
    if(data_in_valid)begin
      _zz_29 <= _zz_27;
      _zz_30 <= _zz_28;
    end
    if(data_in_valid)begin
      _zz_31 <= _zz_29;
      _zz_32 <= _zz_30;
    end
    if(data_in_valid)begin
      _zz_33 <= _zz_31;
      _zz_34 <= _zz_32;
    end
    if(data_in_valid)begin
      _zz_35 <= _zz_33;
      _zz_36 <= _zz_34;
    end
    if(data_in_valid)begin
      _zz_37 <= _zz_35;
      _zz_38 <= _zz_36;
    end
    if(data_in_valid)begin
      _zz_39 <= _zz_37;
      _zz_40 <= _zz_38;
    end
    if(data_in_valid)begin
      _zz_41 <= _zz_39;
      _zz_42 <= _zz_40;
    end
    if(data_in_valid)begin
      _zz_43 <= _zz_41;
      _zz_44 <= _zz_42;
    end
    if(data_in_valid)begin
      _zz_45 <= _zz_43;
      _zz_46 <= _zz_44;
    end
    if(data_in_valid)begin
      _zz_47 <= _zz_45;
      _zz_48 <= _zz_46;
    end
    if(data_in_valid)begin
      _zz_49 <= _zz_47;
      _zz_50 <= _zz_48;
    end
    if(data_in_valid)begin
      _zz_51 <= _zz_49;
      _zz_52 <= _zz_50;
    end
    if(data_in_valid)begin
      _zz_53 <= _zz_51;
      _zz_54 <= _zz_52;
    end
    if(data_in_valid)begin
      _zz_55 <= _zz_53;
      _zz_56 <= _zz_54;
    end
    if(data_in_valid)begin
      _zz_57 <= _zz_55;
      _zz_58 <= _zz_56;
    end
    if(data_in_valid)begin
      _zz_59 <= _zz_57;
      _zz_60 <= _zz_58;
    end
    if(data_in_valid)begin
      _zz_61 <= _zz_59;
      _zz_62 <= _zz_60;
    end
    if(data_in_valid)begin
      _zz_63 <= _zz_61;
      _zz_64 <= _zz_62;
    end
    if(myFFT_1_sdata_out_valid)begin
      sdata_out_regs_0_real <= myFFT_1_sdata_out_payload_0_real;
      sdata_out_regs_0_imag <= myFFT_1_sdata_out_payload_0_imag;
      sdata_out_regs_1_real <= myFFT_1_sdata_out_payload_1_real;
      sdata_out_regs_1_imag <= myFFT_1_sdata_out_payload_1_imag;
      sdata_out_regs_2_real <= myFFT_1_sdata_out_payload_2_real;
      sdata_out_regs_2_imag <= myFFT_1_sdata_out_payload_2_imag;
      sdata_out_regs_3_real <= myFFT_1_sdata_out_payload_3_real;
      sdata_out_regs_3_imag <= myFFT_1_sdata_out_payload_3_imag;
      sdata_out_regs_4_real <= myFFT_1_sdata_out_payload_4_real;
      sdata_out_regs_4_imag <= myFFT_1_sdata_out_payload_4_imag;
      sdata_out_regs_5_real <= myFFT_1_sdata_out_payload_5_real;
      sdata_out_regs_5_imag <= myFFT_1_sdata_out_payload_5_imag;
      sdata_out_regs_6_real <= myFFT_1_sdata_out_payload_6_real;
      sdata_out_regs_6_imag <= myFFT_1_sdata_out_payload_6_imag;
      sdata_out_regs_7_real <= myFFT_1_sdata_out_payload_7_real;
      sdata_out_regs_7_imag <= myFFT_1_sdata_out_payload_7_imag;
      sdata_out_regs_8_real <= myFFT_1_sdata_out_payload_8_real;
      sdata_out_regs_8_imag <= myFFT_1_sdata_out_payload_8_imag;
      sdata_out_regs_9_real <= myFFT_1_sdata_out_payload_9_real;
      sdata_out_regs_9_imag <= myFFT_1_sdata_out_payload_9_imag;
      sdata_out_regs_10_real <= myFFT_1_sdata_out_payload_10_real;
      sdata_out_regs_10_imag <= myFFT_1_sdata_out_payload_10_imag;
      sdata_out_regs_11_real <= myFFT_1_sdata_out_payload_11_real;
      sdata_out_regs_11_imag <= myFFT_1_sdata_out_payload_11_imag;
      sdata_out_regs_12_real <= myFFT_1_sdata_out_payload_12_real;
      sdata_out_regs_12_imag <= myFFT_1_sdata_out_payload_12_imag;
      sdata_out_regs_13_real <= myFFT_1_sdata_out_payload_13_real;
      sdata_out_regs_13_imag <= myFFT_1_sdata_out_payload_13_imag;
      sdata_out_regs_14_real <= myFFT_1_sdata_out_payload_14_real;
      sdata_out_regs_14_imag <= myFFT_1_sdata_out_payload_14_imag;
      sdata_out_regs_15_real <= myFFT_1_sdata_out_payload_15_real;
      sdata_out_regs_15_imag <= myFFT_1_sdata_out_payload_15_imag;
      sdata_out_regs_16_real <= myFFT_1_sdata_out_payload_16_real;
      sdata_out_regs_16_imag <= myFFT_1_sdata_out_payload_16_imag;
      sdata_out_regs_17_real <= myFFT_1_sdata_out_payload_17_real;
      sdata_out_regs_17_imag <= myFFT_1_sdata_out_payload_17_imag;
      sdata_out_regs_18_real <= myFFT_1_sdata_out_payload_18_real;
      sdata_out_regs_18_imag <= myFFT_1_sdata_out_payload_18_imag;
      sdata_out_regs_19_real <= myFFT_1_sdata_out_payload_19_real;
      sdata_out_regs_19_imag <= myFFT_1_sdata_out_payload_19_imag;
      sdata_out_regs_20_real <= myFFT_1_sdata_out_payload_20_real;
      sdata_out_regs_20_imag <= myFFT_1_sdata_out_payload_20_imag;
      sdata_out_regs_21_real <= myFFT_1_sdata_out_payload_21_real;
      sdata_out_regs_21_imag <= myFFT_1_sdata_out_payload_21_imag;
      sdata_out_regs_22_real <= myFFT_1_sdata_out_payload_22_real;
      sdata_out_regs_22_imag <= myFFT_1_sdata_out_payload_22_imag;
      sdata_out_regs_23_real <= myFFT_1_sdata_out_payload_23_real;
      sdata_out_regs_23_imag <= myFFT_1_sdata_out_payload_23_imag;
      sdata_out_regs_24_real <= myFFT_1_sdata_out_payload_24_real;
      sdata_out_regs_24_imag <= myFFT_1_sdata_out_payload_24_imag;
      sdata_out_regs_25_real <= myFFT_1_sdata_out_payload_25_real;
      sdata_out_regs_25_imag <= myFFT_1_sdata_out_payload_25_imag;
      sdata_out_regs_26_real <= myFFT_1_sdata_out_payload_26_real;
      sdata_out_regs_26_imag <= myFFT_1_sdata_out_payload_26_imag;
      sdata_out_regs_27_real <= myFFT_1_sdata_out_payload_27_real;
      sdata_out_regs_27_imag <= myFFT_1_sdata_out_payload_27_imag;
      sdata_out_regs_28_real <= myFFT_1_sdata_out_payload_28_real;
      sdata_out_regs_28_imag <= myFFT_1_sdata_out_payload_28_imag;
      sdata_out_regs_29_real <= myFFT_1_sdata_out_payload_29_real;
      sdata_out_regs_29_imag <= myFFT_1_sdata_out_payload_29_imag;
      sdata_out_regs_30_real <= myFFT_1_sdata_out_payload_30_real;
      sdata_out_regs_30_imag <= myFFT_1_sdata_out_payload_30_imag;
      sdata_out_regs_31_real <= myFFT_1_sdata_out_payload_31_real;
      sdata_out_regs_31_imag <= myFFT_1_sdata_out_payload_31_imag;
    end
  end

  always @ (posedge clk or posedge reset) begin
    if (reset) begin
      count_up_inside_cnt_value <= 5'h0;
      myFFT_1_sdata_out_valid_regNext <= 1'b0;
      null_cnt_value <= 5'h0;
      null_cond_period_minus_1 <= 1'b0;
    end else begin
      count_up_inside_cnt_value <= count_up_inside_cnt_valueNext;
      myFFT_1_sdata_out_valid_regNext <= myFFT_1_sdata_out_valid;
      null_cnt_value <= null_cnt_valueNext;
      if(myFFT_1_sdata_out_valid_regNext)begin
        null_cond_period_minus_1 <= 1'b1;
      end else begin
        if(null_cnt_willOverflow)begin
          null_cond_period_minus_1 <= 1'b0;
        end
      end
    end
  end


endmodule

module MyFFT (
  input               io_data_in_valid,
  input      [15:0]   io_data_in_payload_0_real,
  input      [15:0]   io_data_in_payload_0_imag,
  input      [15:0]   io_data_in_payload_1_real,
  input      [15:0]   io_data_in_payload_1_imag,
  input      [15:0]   io_data_in_payload_2_real,
  input      [15:0]   io_data_in_payload_2_imag,
  input      [15:0]   io_data_in_payload_3_real,
  input      [15:0]   io_data_in_payload_3_imag,
  input      [15:0]   io_data_in_payload_4_real,
  input      [15:0]   io_data_in_payload_4_imag,
  input      [15:0]   io_data_in_payload_5_real,
  input      [15:0]   io_data_in_payload_5_imag,
  input      [15:0]   io_data_in_payload_6_real,
  input      [15:0]   io_data_in_payload_6_imag,
  input      [15:0]   io_data_in_payload_7_real,
  input      [15:0]   io_data_in_payload_7_imag,
  input      [15:0]   io_data_in_payload_8_real,
  input      [15:0]   io_data_in_payload_8_imag,
  input      [15:0]   io_data_in_payload_9_real,
  input      [15:0]   io_data_in_payload_9_imag,
  input      [15:0]   io_data_in_payload_10_real,
  input      [15:0]   io_data_in_payload_10_imag,
  input      [15:0]   io_data_in_payload_11_real,
  input      [15:0]   io_data_in_payload_11_imag,
  input      [15:0]   io_data_in_payload_12_real,
  input      [15:0]   io_data_in_payload_12_imag,
  input      [15:0]   io_data_in_payload_13_real,
  input      [15:0]   io_data_in_payload_13_imag,
  input      [15:0]   io_data_in_payload_14_real,
  input      [15:0]   io_data_in_payload_14_imag,
  input      [15:0]   io_data_in_payload_15_real,
  input      [15:0]   io_data_in_payload_15_imag,
  input      [15:0]   io_data_in_payload_16_real,
  input      [15:0]   io_data_in_payload_16_imag,
  input      [15:0]   io_data_in_payload_17_real,
  input      [15:0]   io_data_in_payload_17_imag,
  input      [15:0]   io_data_in_payload_18_real,
  input      [15:0]   io_data_in_payload_18_imag,
  input      [15:0]   io_data_in_payload_19_real,
  input      [15:0]   io_data_in_payload_19_imag,
  input      [15:0]   io_data_in_payload_20_real,
  input      [15:0]   io_data_in_payload_20_imag,
  input      [15:0]   io_data_in_payload_21_real,
  input      [15:0]   io_data_in_payload_21_imag,
  input      [15:0]   io_data_in_payload_22_real,
  input      [15:0]   io_data_in_payload_22_imag,
  input      [15:0]   io_data_in_payload_23_real,
  input      [15:0]   io_data_in_payload_23_imag,
  input      [15:0]   io_data_in_payload_24_real,
  input      [15:0]   io_data_in_payload_24_imag,
  input      [15:0]   io_data_in_payload_25_real,
  input      [15:0]   io_data_in_payload_25_imag,
  input      [15:0]   io_data_in_payload_26_real,
  input      [15:0]   io_data_in_payload_26_imag,
  input      [15:0]   io_data_in_payload_27_real,
  input      [15:0]   io_data_in_payload_27_imag,
  input      [15:0]   io_data_in_payload_28_real,
  input      [15:0]   io_data_in_payload_28_imag,
  input      [15:0]   io_data_in_payload_29_real,
  input      [15:0]   io_data_in_payload_29_imag,
  input      [15:0]   io_data_in_payload_30_real,
  input      [15:0]   io_data_in_payload_30_imag,
  input      [15:0]   io_data_in_payload_31_real,
  input      [15:0]   io_data_in_payload_31_imag,
  output              sdata_out_valid,
  output     [15:0]   sdata_out_payload_0_real,
  output     [15:0]   sdata_out_payload_0_imag,
  output     [15:0]   sdata_out_payload_1_real,
  output     [15:0]   sdata_out_payload_1_imag,
  output     [15:0]   sdata_out_payload_2_real,
  output     [15:0]   sdata_out_payload_2_imag,
  output     [15:0]   sdata_out_payload_3_real,
  output     [15:0]   sdata_out_payload_3_imag,
  output     [15:0]   sdata_out_payload_4_real,
  output     [15:0]   sdata_out_payload_4_imag,
  output     [15:0]   sdata_out_payload_5_real,
  output     [15:0]   sdata_out_payload_5_imag,
  output     [15:0]   sdata_out_payload_6_real,
  output     [15:0]   sdata_out_payload_6_imag,
  output     [15:0]   sdata_out_payload_7_real,
  output     [15:0]   sdata_out_payload_7_imag,
  output     [15:0]   sdata_out_payload_8_real,
  output     [15:0]   sdata_out_payload_8_imag,
  output     [15:0]   sdata_out_payload_9_real,
  output     [15:0]   sdata_out_payload_9_imag,
  output     [15:0]   sdata_out_payload_10_real,
  output     [15:0]   sdata_out_payload_10_imag,
  output     [15:0]   sdata_out_payload_11_real,
  output     [15:0]   sdata_out_payload_11_imag,
  output     [15:0]   sdata_out_payload_12_real,
  output     [15:0]   sdata_out_payload_12_imag,
  output     [15:0]   sdata_out_payload_13_real,
  output     [15:0]   sdata_out_payload_13_imag,
  output     [15:0]   sdata_out_payload_14_real,
  output     [15:0]   sdata_out_payload_14_imag,
  output     [15:0]   sdata_out_payload_15_real,
  output     [15:0]   sdata_out_payload_15_imag,
  output     [15:0]   sdata_out_payload_16_real,
  output     [15:0]   sdata_out_payload_16_imag,
  output     [15:0]   sdata_out_payload_17_real,
  output     [15:0]   sdata_out_payload_17_imag,
  output     [15:0]   sdata_out_payload_18_real,
  output     [15:0]   sdata_out_payload_18_imag,
  output     [15:0]   sdata_out_payload_19_real,
  output     [15:0]   sdata_out_payload_19_imag,
  output     [15:0]   sdata_out_payload_20_real,
  output     [15:0]   sdata_out_payload_20_imag,
  output     [15:0]   sdata_out_payload_21_real,
  output     [15:0]   sdata_out_payload_21_imag,
  output     [15:0]   sdata_out_payload_22_real,
  output     [15:0]   sdata_out_payload_22_imag,
  output     [15:0]   sdata_out_payload_23_real,
  output     [15:0]   sdata_out_payload_23_imag,
  output     [15:0]   sdata_out_payload_24_real,
  output     [15:0]   sdata_out_payload_24_imag,
  output     [15:0]   sdata_out_payload_25_real,
  output     [15:0]   sdata_out_payload_25_imag,
  output     [15:0]   sdata_out_payload_26_real,
  output     [15:0]   sdata_out_payload_26_imag,
  output     [15:0]   sdata_out_payload_27_real,
  output     [15:0]   sdata_out_payload_27_imag,
  output     [15:0]   sdata_out_payload_28_real,
  output     [15:0]   sdata_out_payload_28_imag,
  output     [15:0]   sdata_out_payload_29_real,
  output     [15:0]   sdata_out_payload_29_imag,
  output     [15:0]   sdata_out_payload_30_real,
  output     [15:0]   sdata_out_payload_30_imag,
  output     [15:0]   sdata_out_payload_31_real,
  output     [15:0]   sdata_out_payload_31_imag,
  input               clk,
  input               reset
);
  wire       [31:0]   _zz_401;
  wire       [31:0]   _zz_402;
  wire       [31:0]   _zz_403;
  wire       [31:0]   _zz_404;
  wire       [31:0]   _zz_405;
  wire       [31:0]   _zz_406;
  wire       [31:0]   _zz_407;
  wire       [31:0]   _zz_408;
  wire       [31:0]   _zz_409;
  wire       [31:0]   _zz_410;
  wire       [31:0]   _zz_411;
  wire       [31:0]   _zz_412;
  wire       [31:0]   _zz_413;
  wire       [31:0]   _zz_414;
  wire       [31:0]   _zz_415;
  wire       [31:0]   _zz_416;
  wire       [31:0]   _zz_417;
  wire       [31:0]   _zz_418;
  wire       [31:0]   _zz_419;
  wire       [31:0]   _zz_420;
  wire       [31:0]   _zz_421;
  wire       [31:0]   _zz_422;
  wire       [31:0]   _zz_423;
  wire       [31:0]   _zz_424;
  wire       [31:0]   _zz_425;
  wire       [31:0]   _zz_426;
  wire       [31:0]   _zz_427;
  wire       [31:0]   _zz_428;
  wire       [31:0]   _zz_429;
  wire       [31:0]   _zz_430;
  wire       [31:0]   _zz_431;
  wire       [31:0]   _zz_432;
  wire       [31:0]   _zz_433;
  wire       [31:0]   _zz_434;
  wire       [31:0]   _zz_435;
  wire       [31:0]   _zz_436;
  wire       [31:0]   _zz_437;
  wire       [31:0]   _zz_438;
  wire       [31:0]   _zz_439;
  wire       [31:0]   _zz_440;
  wire       [31:0]   _zz_441;
  wire       [31:0]   _zz_442;
  wire       [31:0]   _zz_443;
  wire       [31:0]   _zz_444;
  wire       [31:0]   _zz_445;
  wire       [31:0]   _zz_446;
  wire       [31:0]   _zz_447;
  wire       [31:0]   _zz_448;
  wire       [31:0]   _zz_449;
  wire       [31:0]   _zz_450;
  wire       [31:0]   _zz_451;
  wire       [31:0]   _zz_452;
  wire       [31:0]   _zz_453;
  wire       [31:0]   _zz_454;
  wire       [31:0]   _zz_455;
  wire       [31:0]   _zz_456;
  wire       [31:0]   _zz_457;
  wire       [31:0]   _zz_458;
  wire       [31:0]   _zz_459;
  wire       [31:0]   _zz_460;
  wire       [31:0]   _zz_461;
  wire       [31:0]   _zz_462;
  wire       [31:0]   _zz_463;
  wire       [31:0]   _zz_464;
  wire       [31:0]   _zz_465;
  wire       [31:0]   _zz_466;
  wire       [31:0]   _zz_467;
  wire       [31:0]   _zz_468;
  wire       [31:0]   _zz_469;
  wire       [31:0]   _zz_470;
  wire       [31:0]   _zz_471;
  wire       [31:0]   _zz_472;
  wire       [31:0]   _zz_473;
  wire       [31:0]   _zz_474;
  wire       [31:0]   _zz_475;
  wire       [31:0]   _zz_476;
  wire       [31:0]   _zz_477;
  wire       [31:0]   _zz_478;
  wire       [31:0]   _zz_479;
  wire       [31:0]   _zz_480;
  wire       [31:0]   _zz_481;
  wire       [31:0]   _zz_482;
  wire       [31:0]   _zz_483;
  wire       [31:0]   _zz_484;
  wire       [31:0]   _zz_485;
  wire       [31:0]   _zz_486;
  wire       [31:0]   _zz_487;
  wire       [31:0]   _zz_488;
  wire       [31:0]   _zz_489;
  wire       [31:0]   _zz_490;
  wire       [31:0]   _zz_491;
  wire       [31:0]   _zz_492;
  wire       [31:0]   _zz_493;
  wire       [31:0]   _zz_494;
  wire       [31:0]   _zz_495;
  wire       [31:0]   _zz_496;
  wire       [31:0]   _zz_497;
  wire       [31:0]   _zz_498;
  wire       [31:0]   _zz_499;
  wire       [31:0]   _zz_500;
  wire       [31:0]   _zz_501;
  wire       [31:0]   _zz_502;
  wire       [31:0]   _zz_503;
  wire       [31:0]   _zz_504;
  wire       [31:0]   _zz_505;
  wire       [31:0]   _zz_506;
  wire       [31:0]   _zz_507;
  wire       [31:0]   _zz_508;
  wire       [31:0]   _zz_509;
  wire       [31:0]   _zz_510;
  wire       [31:0]   _zz_511;
  wire       [31:0]   _zz_512;
  wire       [31:0]   _zz_513;
  wire       [31:0]   _zz_514;
  wire       [31:0]   _zz_515;
  wire       [31:0]   _zz_516;
  wire       [31:0]   _zz_517;
  wire       [31:0]   _zz_518;
  wire       [31:0]   _zz_519;
  wire       [31:0]   _zz_520;
  wire       [31:0]   _zz_521;
  wire       [31:0]   _zz_522;
  wire       [31:0]   _zz_523;
  wire       [31:0]   _zz_524;
  wire       [31:0]   _zz_525;
  wire       [31:0]   _zz_526;
  wire       [31:0]   _zz_527;
  wire       [31:0]   _zz_528;
  wire       [31:0]   _zz_529;
  wire       [31:0]   _zz_530;
  wire       [31:0]   _zz_531;
  wire       [31:0]   _zz_532;
  wire       [31:0]   _zz_533;
  wire       [31:0]   _zz_534;
  wire       [31:0]   _zz_535;
  wire       [31:0]   _zz_536;
  wire       [31:0]   _zz_537;
  wire       [31:0]   _zz_538;
  wire       [31:0]   _zz_539;
  wire       [31:0]   _zz_540;
  wire       [31:0]   _zz_541;
  wire       [31:0]   _zz_542;
  wire       [31:0]   _zz_543;
  wire       [31:0]   _zz_544;
  wire       [31:0]   _zz_545;
  wire       [31:0]   _zz_546;
  wire       [31:0]   _zz_547;
  wire       [31:0]   _zz_548;
  wire       [31:0]   _zz_549;
  wire       [31:0]   _zz_550;
  wire       [31:0]   _zz_551;
  wire       [31:0]   _zz_552;
  wire       [31:0]   _zz_553;
  wire       [31:0]   _zz_554;
  wire       [31:0]   _zz_555;
  wire       [31:0]   _zz_556;
  wire       [31:0]   _zz_557;
  wire       [31:0]   _zz_558;
  wire       [31:0]   _zz_559;
  wire       [31:0]   _zz_560;
  wire       [31:0]   _zz_561;
  wire       [31:0]   _zz_562;
  wire       [31:0]   _zz_563;
  wire       [31:0]   _zz_564;
  wire       [31:0]   _zz_565;
  wire       [31:0]   _zz_566;
  wire       [31:0]   _zz_567;
  wire       [31:0]   _zz_568;
  wire       [31:0]   _zz_569;
  wire       [31:0]   _zz_570;
  wire       [31:0]   _zz_571;
  wire       [31:0]   _zz_572;
  wire       [31:0]   _zz_573;
  wire       [31:0]   _zz_574;
  wire       [31:0]   _zz_575;
  wire       [31:0]   _zz_576;
  wire       [31:0]   _zz_577;
  wire       [31:0]   _zz_578;
  wire       [31:0]   _zz_579;
  wire       [31:0]   _zz_580;
  wire       [31:0]   _zz_581;
  wire       [31:0]   _zz_582;
  wire       [31:0]   _zz_583;
  wire       [31:0]   _zz_584;
  wire       [31:0]   _zz_585;
  wire       [31:0]   _zz_586;
  wire       [31:0]   _zz_587;
  wire       [31:0]   _zz_588;
  wire       [31:0]   _zz_589;
  wire       [31:0]   _zz_590;
  wire       [31:0]   _zz_591;
  wire       [31:0]   _zz_592;
  wire       [31:0]   _zz_593;
  wire       [31:0]   _zz_594;
  wire       [31:0]   _zz_595;
  wire       [31:0]   _zz_596;
  wire       [31:0]   _zz_597;
  wire       [31:0]   _zz_598;
  wire       [31:0]   _zz_599;
  wire       [31:0]   _zz_600;
  wire       [31:0]   _zz_601;
  wire       [31:0]   _zz_602;
  wire       [31:0]   _zz_603;
  wire       [31:0]   _zz_604;
  wire       [31:0]   _zz_605;
  wire       [31:0]   _zz_606;
  wire       [31:0]   _zz_607;
  wire       [31:0]   _zz_608;
  wire       [31:0]   _zz_609;
  wire       [31:0]   _zz_610;
  wire       [31:0]   _zz_611;
  wire       [31:0]   _zz_612;
  wire       [31:0]   _zz_613;
  wire       [31:0]   _zz_614;
  wire       [31:0]   _zz_615;
  wire       [31:0]   _zz_616;
  wire       [31:0]   _zz_617;
  wire       [31:0]   _zz_618;
  wire       [31:0]   _zz_619;
  wire       [31:0]   _zz_620;
  wire       [31:0]   _zz_621;
  wire       [31:0]   _zz_622;
  wire       [31:0]   _zz_623;
  wire       [31:0]   _zz_624;
  wire       [31:0]   _zz_625;
  wire       [31:0]   _zz_626;
  wire       [31:0]   _zz_627;
  wire       [31:0]   _zz_628;
  wire       [31:0]   _zz_629;
  wire       [31:0]   _zz_630;
  wire       [31:0]   _zz_631;
  wire       [31:0]   _zz_632;
  wire       [31:0]   _zz_633;
  wire       [31:0]   _zz_634;
  wire       [31:0]   _zz_635;
  wire       [31:0]   _zz_636;
  wire       [31:0]   _zz_637;
  wire       [31:0]   _zz_638;
  wire       [31:0]   _zz_639;
  wire       [31:0]   _zz_640;
  wire       [31:0]   _zz_641;
  wire       [31:0]   _zz_642;
  wire       [31:0]   _zz_643;
  wire       [31:0]   _zz_644;
  wire       [31:0]   _zz_645;
  wire       [31:0]   _zz_646;
  wire       [31:0]   _zz_647;
  wire       [31:0]   _zz_648;
  wire       [31:0]   _zz_649;
  wire       [31:0]   _zz_650;
  wire       [31:0]   _zz_651;
  wire       [31:0]   _zz_652;
  wire       [31:0]   _zz_653;
  wire       [31:0]   _zz_654;
  wire       [31:0]   _zz_655;
  wire       [31:0]   _zz_656;
  wire       [31:0]   _zz_657;
  wire       [31:0]   _zz_658;
  wire       [31:0]   _zz_659;
  wire       [31:0]   _zz_660;
  wire       [31:0]   _zz_661;
  wire       [31:0]   _zz_662;
  wire       [31:0]   _zz_663;
  wire       [31:0]   _zz_664;
  wire       [31:0]   _zz_665;
  wire       [31:0]   _zz_666;
  wire       [31:0]   _zz_667;
  wire       [31:0]   _zz_668;
  wire       [31:0]   _zz_669;
  wire       [31:0]   _zz_670;
  wire       [31:0]   _zz_671;
  wire       [31:0]   _zz_672;
  wire       [31:0]   _zz_673;
  wire       [31:0]   _zz_674;
  wire       [31:0]   _zz_675;
  wire       [31:0]   _zz_676;
  wire       [31:0]   _zz_677;
  wire       [31:0]   _zz_678;
  wire       [31:0]   _zz_679;
  wire       [31:0]   _zz_680;
  wire       [31:0]   _zz_681;
  wire       [31:0]   _zz_682;
  wire       [31:0]   _zz_683;
  wire       [31:0]   _zz_684;
  wire       [31:0]   _zz_685;
  wire       [31:0]   _zz_686;
  wire       [31:0]   _zz_687;
  wire       [31:0]   _zz_688;
  wire       [31:0]   _zz_689;
  wire       [31:0]   _zz_690;
  wire       [31:0]   _zz_691;
  wire       [31:0]   _zz_692;
  wire       [31:0]   _zz_693;
  wire       [31:0]   _zz_694;
  wire       [31:0]   _zz_695;
  wire       [31:0]   _zz_696;
  wire       [31:0]   _zz_697;
  wire       [31:0]   _zz_698;
  wire       [31:0]   _zz_699;
  wire       [31:0]   _zz_700;
  wire       [31:0]   _zz_701;
  wire       [31:0]   _zz_702;
  wire       [31:0]   _zz_703;
  wire       [31:0]   _zz_704;
  wire       [31:0]   _zz_705;
  wire       [31:0]   _zz_706;
  wire       [31:0]   _zz_707;
  wire       [31:0]   _zz_708;
  wire       [31:0]   _zz_709;
  wire       [31:0]   _zz_710;
  wire       [31:0]   _zz_711;
  wire       [31:0]   _zz_712;
  wire       [31:0]   _zz_713;
  wire       [31:0]   _zz_714;
  wire       [31:0]   _zz_715;
  wire       [31:0]   _zz_716;
  wire       [31:0]   _zz_717;
  wire       [31:0]   _zz_718;
  wire       [31:0]   _zz_719;
  wire       [31:0]   _zz_720;
  wire       [31:0]   _zz_721;
  wire       [31:0]   _zz_722;
  wire       [31:0]   _zz_723;
  wire       [31:0]   _zz_724;
  wire       [31:0]   _zz_725;
  wire       [31:0]   _zz_726;
  wire       [31:0]   _zz_727;
  wire       [31:0]   _zz_728;
  wire       [31:0]   _zz_729;
  wire       [31:0]   _zz_730;
  wire       [31:0]   _zz_731;
  wire       [31:0]   _zz_732;
  wire       [31:0]   _zz_733;
  wire       [31:0]   _zz_734;
  wire       [31:0]   _zz_735;
  wire       [31:0]   _zz_736;
  wire       [31:0]   _zz_737;
  wire       [31:0]   _zz_738;
  wire       [31:0]   _zz_739;
  wire       [31:0]   _zz_740;
  wire       [31:0]   _zz_741;
  wire       [31:0]   _zz_742;
  wire       [31:0]   _zz_743;
  wire       [31:0]   _zz_744;
  wire       [31:0]   _zz_745;
  wire       [31:0]   _zz_746;
  wire       [31:0]   _zz_747;
  wire       [31:0]   _zz_748;
  wire       [31:0]   _zz_749;
  wire       [31:0]   _zz_750;
  wire       [31:0]   _zz_751;
  wire       [31:0]   _zz_752;
  wire       [31:0]   _zz_753;
  wire       [31:0]   _zz_754;
  wire       [31:0]   _zz_755;
  wire       [31:0]   _zz_756;
  wire       [31:0]   _zz_757;
  wire       [31:0]   _zz_758;
  wire       [31:0]   _zz_759;
  wire       [31:0]   _zz_760;
  wire       [31:0]   _zz_761;
  wire       [31:0]   _zz_762;
  wire       [31:0]   _zz_763;
  wire       [31:0]   _zz_764;
  wire       [31:0]   _zz_765;
  wire       [31:0]   _zz_766;
  wire       [31:0]   _zz_767;
  wire       [31:0]   _zz_768;
  wire       [31:0]   _zz_769;
  wire       [31:0]   _zz_770;
  wire       [31:0]   _zz_771;
  wire       [31:0]   _zz_772;
  wire       [31:0]   _zz_773;
  wire       [31:0]   _zz_774;
  wire       [31:0]   _zz_775;
  wire       [31:0]   _zz_776;
  wire       [31:0]   _zz_777;
  wire       [31:0]   _zz_778;
  wire       [31:0]   _zz_779;
  wire       [31:0]   _zz_780;
  wire       [31:0]   _zz_781;
  wire       [31:0]   _zz_782;
  wire       [31:0]   _zz_783;
  wire       [31:0]   _zz_784;
  wire       [31:0]   _zz_785;
  wire       [31:0]   _zz_786;
  wire       [31:0]   _zz_787;
  wire       [31:0]   _zz_788;
  wire       [31:0]   _zz_789;
  wire       [31:0]   _zz_790;
  wire       [31:0]   _zz_791;
  wire       [31:0]   _zz_792;
  wire       [31:0]   _zz_793;
  wire       [31:0]   _zz_794;
  wire       [31:0]   _zz_795;
  wire       [31:0]   _zz_796;
  wire       [31:0]   _zz_797;
  wire       [31:0]   _zz_798;
  wire       [31:0]   _zz_799;
  wire       [31:0]   _zz_800;
  wire       [31:0]   _zz_801;
  wire       [31:0]   _zz_802;
  wire       [31:0]   _zz_803;
  wire       [31:0]   _zz_804;
  wire       [31:0]   _zz_805;
  wire       [31:0]   _zz_806;
  wire       [31:0]   _zz_807;
  wire       [31:0]   _zz_808;
  wire       [31:0]   _zz_809;
  wire       [31:0]   _zz_810;
  wire       [31:0]   _zz_811;
  wire       [31:0]   _zz_812;
  wire       [31:0]   _zz_813;
  wire       [31:0]   _zz_814;
  wire       [31:0]   _zz_815;
  wire       [31:0]   _zz_816;
  wire       [31:0]   _zz_817;
  wire       [31:0]   _zz_818;
  wire       [31:0]   _zz_819;
  wire       [31:0]   _zz_820;
  wire       [31:0]   _zz_821;
  wire       [31:0]   _zz_822;
  wire       [31:0]   _zz_823;
  wire       [31:0]   _zz_824;
  wire       [31:0]   _zz_825;
  wire       [31:0]   _zz_826;
  wire       [31:0]   _zz_827;
  wire       [31:0]   _zz_828;
  wire       [31:0]   _zz_829;
  wire       [31:0]   _zz_830;
  wire       [31:0]   _zz_831;
  wire       [31:0]   _zz_832;
  wire       [31:0]   _zz_833;
  wire       [31:0]   _zz_834;
  wire       [31:0]   _zz_835;
  wire       [31:0]   _zz_836;
  wire       [31:0]   _zz_837;
  wire       [31:0]   _zz_838;
  wire       [31:0]   _zz_839;
  wire       [31:0]   _zz_840;
  wire       [31:0]   _zz_841;
  wire       [31:0]   _zz_842;
  wire       [31:0]   _zz_843;
  wire       [31:0]   _zz_844;
  wire       [31:0]   _zz_845;
  wire       [31:0]   _zz_846;
  wire       [31:0]   _zz_847;
  wire       [31:0]   _zz_848;
  wire       [31:0]   _zz_849;
  wire       [31:0]   _zz_850;
  wire       [31:0]   _zz_851;
  wire       [31:0]   _zz_852;
  wire       [31:0]   _zz_853;
  wire       [31:0]   _zz_854;
  wire       [31:0]   _zz_855;
  wire       [31:0]   _zz_856;
  wire       [31:0]   _zz_857;
  wire       [31:0]   _zz_858;
  wire       [31:0]   _zz_859;
  wire       [31:0]   _zz_860;
  wire       [31:0]   _zz_861;
  wire       [31:0]   _zz_862;
  wire       [31:0]   _zz_863;
  wire       [31:0]   _zz_864;
  wire       [31:0]   _zz_865;
  wire       [31:0]   _zz_866;
  wire       [31:0]   _zz_867;
  wire       [31:0]   _zz_868;
  wire       [31:0]   _zz_869;
  wire       [31:0]   _zz_870;
  wire       [31:0]   _zz_871;
  wire       [31:0]   _zz_872;
  wire       [31:0]   _zz_873;
  wire       [31:0]   _zz_874;
  wire       [31:0]   _zz_875;
  wire       [31:0]   _zz_876;
  wire       [31:0]   _zz_877;
  wire       [31:0]   _zz_878;
  wire       [31:0]   _zz_879;
  wire       [31:0]   _zz_880;
  wire       [31:0]   fixTo_dout;
  wire       [31:0]   fixTo_1_dout;
  wire       [15:0]   fixTo_2_dout;
  wire       [15:0]   fixTo_3_dout;
  wire       [15:0]   fixTo_4_dout;
  wire       [15:0]   fixTo_5_dout;
  wire       [31:0]   fixTo_6_dout;
  wire       [31:0]   fixTo_7_dout;
  wire       [15:0]   fixTo_8_dout;
  wire       [15:0]   fixTo_9_dout;
  wire       [15:0]   fixTo_10_dout;
  wire       [15:0]   fixTo_11_dout;
  wire       [31:0]   fixTo_12_dout;
  wire       [31:0]   fixTo_13_dout;
  wire       [15:0]   fixTo_14_dout;
  wire       [15:0]   fixTo_15_dout;
  wire       [15:0]   fixTo_16_dout;
  wire       [15:0]   fixTo_17_dout;
  wire       [31:0]   fixTo_18_dout;
  wire       [31:0]   fixTo_19_dout;
  wire       [15:0]   fixTo_20_dout;
  wire       [15:0]   fixTo_21_dout;
  wire       [15:0]   fixTo_22_dout;
  wire       [15:0]   fixTo_23_dout;
  wire       [31:0]   fixTo_24_dout;
  wire       [31:0]   fixTo_25_dout;
  wire       [15:0]   fixTo_26_dout;
  wire       [15:0]   fixTo_27_dout;
  wire       [15:0]   fixTo_28_dout;
  wire       [15:0]   fixTo_29_dout;
  wire       [31:0]   fixTo_30_dout;
  wire       [31:0]   fixTo_31_dout;
  wire       [15:0]   fixTo_32_dout;
  wire       [15:0]   fixTo_33_dout;
  wire       [15:0]   fixTo_34_dout;
  wire       [15:0]   fixTo_35_dout;
  wire       [31:0]   fixTo_36_dout;
  wire       [31:0]   fixTo_37_dout;
  wire       [15:0]   fixTo_38_dout;
  wire       [15:0]   fixTo_39_dout;
  wire       [15:0]   fixTo_40_dout;
  wire       [15:0]   fixTo_41_dout;
  wire       [31:0]   fixTo_42_dout;
  wire       [31:0]   fixTo_43_dout;
  wire       [15:0]   fixTo_44_dout;
  wire       [15:0]   fixTo_45_dout;
  wire       [15:0]   fixTo_46_dout;
  wire       [15:0]   fixTo_47_dout;
  wire       [31:0]   fixTo_48_dout;
  wire       [31:0]   fixTo_49_dout;
  wire       [15:0]   fixTo_50_dout;
  wire       [15:0]   fixTo_51_dout;
  wire       [15:0]   fixTo_52_dout;
  wire       [15:0]   fixTo_53_dout;
  wire       [31:0]   fixTo_54_dout;
  wire       [31:0]   fixTo_55_dout;
  wire       [15:0]   fixTo_56_dout;
  wire       [15:0]   fixTo_57_dout;
  wire       [15:0]   fixTo_58_dout;
  wire       [15:0]   fixTo_59_dout;
  wire       [31:0]   fixTo_60_dout;
  wire       [31:0]   fixTo_61_dout;
  wire       [15:0]   fixTo_62_dout;
  wire       [15:0]   fixTo_63_dout;
  wire       [15:0]   fixTo_64_dout;
  wire       [15:0]   fixTo_65_dout;
  wire       [31:0]   fixTo_66_dout;
  wire       [31:0]   fixTo_67_dout;
  wire       [15:0]   fixTo_68_dout;
  wire       [15:0]   fixTo_69_dout;
  wire       [15:0]   fixTo_70_dout;
  wire       [15:0]   fixTo_71_dout;
  wire       [31:0]   fixTo_72_dout;
  wire       [31:0]   fixTo_73_dout;
  wire       [15:0]   fixTo_74_dout;
  wire       [15:0]   fixTo_75_dout;
  wire       [15:0]   fixTo_76_dout;
  wire       [15:0]   fixTo_77_dout;
  wire       [31:0]   fixTo_78_dout;
  wire       [31:0]   fixTo_79_dout;
  wire       [15:0]   fixTo_80_dout;
  wire       [15:0]   fixTo_81_dout;
  wire       [15:0]   fixTo_82_dout;
  wire       [15:0]   fixTo_83_dout;
  wire       [31:0]   fixTo_84_dout;
  wire       [31:0]   fixTo_85_dout;
  wire       [15:0]   fixTo_86_dout;
  wire       [15:0]   fixTo_87_dout;
  wire       [15:0]   fixTo_88_dout;
  wire       [15:0]   fixTo_89_dout;
  wire       [31:0]   fixTo_90_dout;
  wire       [31:0]   fixTo_91_dout;
  wire       [15:0]   fixTo_92_dout;
  wire       [15:0]   fixTo_93_dout;
  wire       [15:0]   fixTo_94_dout;
  wire       [15:0]   fixTo_95_dout;
  wire       [31:0]   fixTo_96_dout;
  wire       [31:0]   fixTo_97_dout;
  wire       [15:0]   fixTo_98_dout;
  wire       [15:0]   fixTo_99_dout;
  wire       [15:0]   fixTo_100_dout;
  wire       [15:0]   fixTo_101_dout;
  wire       [31:0]   fixTo_102_dout;
  wire       [31:0]   fixTo_103_dout;
  wire       [15:0]   fixTo_104_dout;
  wire       [15:0]   fixTo_105_dout;
  wire       [15:0]   fixTo_106_dout;
  wire       [15:0]   fixTo_107_dout;
  wire       [31:0]   fixTo_108_dout;
  wire       [31:0]   fixTo_109_dout;
  wire       [15:0]   fixTo_110_dout;
  wire       [15:0]   fixTo_111_dout;
  wire       [15:0]   fixTo_112_dout;
  wire       [15:0]   fixTo_113_dout;
  wire       [31:0]   fixTo_114_dout;
  wire       [31:0]   fixTo_115_dout;
  wire       [15:0]   fixTo_116_dout;
  wire       [15:0]   fixTo_117_dout;
  wire       [15:0]   fixTo_118_dout;
  wire       [15:0]   fixTo_119_dout;
  wire       [31:0]   fixTo_120_dout;
  wire       [31:0]   fixTo_121_dout;
  wire       [15:0]   fixTo_122_dout;
  wire       [15:0]   fixTo_123_dout;
  wire       [15:0]   fixTo_124_dout;
  wire       [15:0]   fixTo_125_dout;
  wire       [31:0]   fixTo_126_dout;
  wire       [31:0]   fixTo_127_dout;
  wire       [15:0]   fixTo_128_dout;
  wire       [15:0]   fixTo_129_dout;
  wire       [15:0]   fixTo_130_dout;
  wire       [15:0]   fixTo_131_dout;
  wire       [31:0]   fixTo_132_dout;
  wire       [31:0]   fixTo_133_dout;
  wire       [15:0]   fixTo_134_dout;
  wire       [15:0]   fixTo_135_dout;
  wire       [15:0]   fixTo_136_dout;
  wire       [15:0]   fixTo_137_dout;
  wire       [31:0]   fixTo_138_dout;
  wire       [31:0]   fixTo_139_dout;
  wire       [15:0]   fixTo_140_dout;
  wire       [15:0]   fixTo_141_dout;
  wire       [15:0]   fixTo_142_dout;
  wire       [15:0]   fixTo_143_dout;
  wire       [31:0]   fixTo_144_dout;
  wire       [31:0]   fixTo_145_dout;
  wire       [15:0]   fixTo_146_dout;
  wire       [15:0]   fixTo_147_dout;
  wire       [15:0]   fixTo_148_dout;
  wire       [15:0]   fixTo_149_dout;
  wire       [31:0]   fixTo_150_dout;
  wire       [31:0]   fixTo_151_dout;
  wire       [15:0]   fixTo_152_dout;
  wire       [15:0]   fixTo_153_dout;
  wire       [15:0]   fixTo_154_dout;
  wire       [15:0]   fixTo_155_dout;
  wire       [31:0]   fixTo_156_dout;
  wire       [31:0]   fixTo_157_dout;
  wire       [15:0]   fixTo_158_dout;
  wire       [15:0]   fixTo_159_dout;
  wire       [15:0]   fixTo_160_dout;
  wire       [15:0]   fixTo_161_dout;
  wire       [31:0]   fixTo_162_dout;
  wire       [31:0]   fixTo_163_dout;
  wire       [15:0]   fixTo_164_dout;
  wire       [15:0]   fixTo_165_dout;
  wire       [15:0]   fixTo_166_dout;
  wire       [15:0]   fixTo_167_dout;
  wire       [31:0]   fixTo_168_dout;
  wire       [31:0]   fixTo_169_dout;
  wire       [15:0]   fixTo_170_dout;
  wire       [15:0]   fixTo_171_dout;
  wire       [15:0]   fixTo_172_dout;
  wire       [15:0]   fixTo_173_dout;
  wire       [31:0]   fixTo_174_dout;
  wire       [31:0]   fixTo_175_dout;
  wire       [15:0]   fixTo_176_dout;
  wire       [15:0]   fixTo_177_dout;
  wire       [15:0]   fixTo_178_dout;
  wire       [15:0]   fixTo_179_dout;
  wire       [31:0]   fixTo_180_dout;
  wire       [31:0]   fixTo_181_dout;
  wire       [15:0]   fixTo_182_dout;
  wire       [15:0]   fixTo_183_dout;
  wire       [15:0]   fixTo_184_dout;
  wire       [15:0]   fixTo_185_dout;
  wire       [31:0]   fixTo_186_dout;
  wire       [31:0]   fixTo_187_dout;
  wire       [15:0]   fixTo_188_dout;
  wire       [15:0]   fixTo_189_dout;
  wire       [15:0]   fixTo_190_dout;
  wire       [15:0]   fixTo_191_dout;
  wire       [31:0]   fixTo_192_dout;
  wire       [31:0]   fixTo_193_dout;
  wire       [15:0]   fixTo_194_dout;
  wire       [15:0]   fixTo_195_dout;
  wire       [15:0]   fixTo_196_dout;
  wire       [15:0]   fixTo_197_dout;
  wire       [31:0]   fixTo_198_dout;
  wire       [31:0]   fixTo_199_dout;
  wire       [15:0]   fixTo_200_dout;
  wire       [15:0]   fixTo_201_dout;
  wire       [15:0]   fixTo_202_dout;
  wire       [15:0]   fixTo_203_dout;
  wire       [31:0]   fixTo_204_dout;
  wire       [31:0]   fixTo_205_dout;
  wire       [15:0]   fixTo_206_dout;
  wire       [15:0]   fixTo_207_dout;
  wire       [15:0]   fixTo_208_dout;
  wire       [15:0]   fixTo_209_dout;
  wire       [31:0]   fixTo_210_dout;
  wire       [31:0]   fixTo_211_dout;
  wire       [15:0]   fixTo_212_dout;
  wire       [15:0]   fixTo_213_dout;
  wire       [15:0]   fixTo_214_dout;
  wire       [15:0]   fixTo_215_dout;
  wire       [31:0]   fixTo_216_dout;
  wire       [31:0]   fixTo_217_dout;
  wire       [15:0]   fixTo_218_dout;
  wire       [15:0]   fixTo_219_dout;
  wire       [15:0]   fixTo_220_dout;
  wire       [15:0]   fixTo_221_dout;
  wire       [31:0]   fixTo_222_dout;
  wire       [31:0]   fixTo_223_dout;
  wire       [15:0]   fixTo_224_dout;
  wire       [15:0]   fixTo_225_dout;
  wire       [15:0]   fixTo_226_dout;
  wire       [15:0]   fixTo_227_dout;
  wire       [31:0]   fixTo_228_dout;
  wire       [31:0]   fixTo_229_dout;
  wire       [15:0]   fixTo_230_dout;
  wire       [15:0]   fixTo_231_dout;
  wire       [15:0]   fixTo_232_dout;
  wire       [15:0]   fixTo_233_dout;
  wire       [31:0]   fixTo_234_dout;
  wire       [31:0]   fixTo_235_dout;
  wire       [15:0]   fixTo_236_dout;
  wire       [15:0]   fixTo_237_dout;
  wire       [15:0]   fixTo_238_dout;
  wire       [15:0]   fixTo_239_dout;
  wire       [31:0]   fixTo_240_dout;
  wire       [31:0]   fixTo_241_dout;
  wire       [15:0]   fixTo_242_dout;
  wire       [15:0]   fixTo_243_dout;
  wire       [15:0]   fixTo_244_dout;
  wire       [15:0]   fixTo_245_dout;
  wire       [31:0]   fixTo_246_dout;
  wire       [31:0]   fixTo_247_dout;
  wire       [15:0]   fixTo_248_dout;
  wire       [15:0]   fixTo_249_dout;
  wire       [15:0]   fixTo_250_dout;
  wire       [15:0]   fixTo_251_dout;
  wire       [31:0]   fixTo_252_dout;
  wire       [31:0]   fixTo_253_dout;
  wire       [15:0]   fixTo_254_dout;
  wire       [15:0]   fixTo_255_dout;
  wire       [15:0]   fixTo_256_dout;
  wire       [15:0]   fixTo_257_dout;
  wire       [31:0]   fixTo_258_dout;
  wire       [31:0]   fixTo_259_dout;
  wire       [15:0]   fixTo_260_dout;
  wire       [15:0]   fixTo_261_dout;
  wire       [15:0]   fixTo_262_dout;
  wire       [15:0]   fixTo_263_dout;
  wire       [31:0]   fixTo_264_dout;
  wire       [31:0]   fixTo_265_dout;
  wire       [15:0]   fixTo_266_dout;
  wire       [15:0]   fixTo_267_dout;
  wire       [15:0]   fixTo_268_dout;
  wire       [15:0]   fixTo_269_dout;
  wire       [31:0]   fixTo_270_dout;
  wire       [31:0]   fixTo_271_dout;
  wire       [15:0]   fixTo_272_dout;
  wire       [15:0]   fixTo_273_dout;
  wire       [15:0]   fixTo_274_dout;
  wire       [15:0]   fixTo_275_dout;
  wire       [31:0]   fixTo_276_dout;
  wire       [31:0]   fixTo_277_dout;
  wire       [15:0]   fixTo_278_dout;
  wire       [15:0]   fixTo_279_dout;
  wire       [15:0]   fixTo_280_dout;
  wire       [15:0]   fixTo_281_dout;
  wire       [31:0]   fixTo_282_dout;
  wire       [31:0]   fixTo_283_dout;
  wire       [15:0]   fixTo_284_dout;
  wire       [15:0]   fixTo_285_dout;
  wire       [15:0]   fixTo_286_dout;
  wire       [15:0]   fixTo_287_dout;
  wire       [31:0]   fixTo_288_dout;
  wire       [31:0]   fixTo_289_dout;
  wire       [15:0]   fixTo_290_dout;
  wire       [15:0]   fixTo_291_dout;
  wire       [15:0]   fixTo_292_dout;
  wire       [15:0]   fixTo_293_dout;
  wire       [31:0]   fixTo_294_dout;
  wire       [31:0]   fixTo_295_dout;
  wire       [15:0]   fixTo_296_dout;
  wire       [15:0]   fixTo_297_dout;
  wire       [15:0]   fixTo_298_dout;
  wire       [15:0]   fixTo_299_dout;
  wire       [31:0]   fixTo_300_dout;
  wire       [31:0]   fixTo_301_dout;
  wire       [15:0]   fixTo_302_dout;
  wire       [15:0]   fixTo_303_dout;
  wire       [15:0]   fixTo_304_dout;
  wire       [15:0]   fixTo_305_dout;
  wire       [31:0]   fixTo_306_dout;
  wire       [31:0]   fixTo_307_dout;
  wire       [15:0]   fixTo_308_dout;
  wire       [15:0]   fixTo_309_dout;
  wire       [15:0]   fixTo_310_dout;
  wire       [15:0]   fixTo_311_dout;
  wire       [31:0]   fixTo_312_dout;
  wire       [31:0]   fixTo_313_dout;
  wire       [15:0]   fixTo_314_dout;
  wire       [15:0]   fixTo_315_dout;
  wire       [15:0]   fixTo_316_dout;
  wire       [15:0]   fixTo_317_dout;
  wire       [31:0]   fixTo_318_dout;
  wire       [31:0]   fixTo_319_dout;
  wire       [15:0]   fixTo_320_dout;
  wire       [15:0]   fixTo_321_dout;
  wire       [15:0]   fixTo_322_dout;
  wire       [15:0]   fixTo_323_dout;
  wire       [31:0]   fixTo_324_dout;
  wire       [31:0]   fixTo_325_dout;
  wire       [15:0]   fixTo_326_dout;
  wire       [15:0]   fixTo_327_dout;
  wire       [15:0]   fixTo_328_dout;
  wire       [15:0]   fixTo_329_dout;
  wire       [31:0]   fixTo_330_dout;
  wire       [31:0]   fixTo_331_dout;
  wire       [15:0]   fixTo_332_dout;
  wire       [15:0]   fixTo_333_dout;
  wire       [15:0]   fixTo_334_dout;
  wire       [15:0]   fixTo_335_dout;
  wire       [31:0]   fixTo_336_dout;
  wire       [31:0]   fixTo_337_dout;
  wire       [15:0]   fixTo_338_dout;
  wire       [15:0]   fixTo_339_dout;
  wire       [15:0]   fixTo_340_dout;
  wire       [15:0]   fixTo_341_dout;
  wire       [31:0]   fixTo_342_dout;
  wire       [31:0]   fixTo_343_dout;
  wire       [15:0]   fixTo_344_dout;
  wire       [15:0]   fixTo_345_dout;
  wire       [15:0]   fixTo_346_dout;
  wire       [15:0]   fixTo_347_dout;
  wire       [31:0]   fixTo_348_dout;
  wire       [31:0]   fixTo_349_dout;
  wire       [15:0]   fixTo_350_dout;
  wire       [15:0]   fixTo_351_dout;
  wire       [15:0]   fixTo_352_dout;
  wire       [15:0]   fixTo_353_dout;
  wire       [31:0]   fixTo_354_dout;
  wire       [31:0]   fixTo_355_dout;
  wire       [15:0]   fixTo_356_dout;
  wire       [15:0]   fixTo_357_dout;
  wire       [15:0]   fixTo_358_dout;
  wire       [15:0]   fixTo_359_dout;
  wire       [31:0]   fixTo_360_dout;
  wire       [31:0]   fixTo_361_dout;
  wire       [15:0]   fixTo_362_dout;
  wire       [15:0]   fixTo_363_dout;
  wire       [15:0]   fixTo_364_dout;
  wire       [15:0]   fixTo_365_dout;
  wire       [31:0]   fixTo_366_dout;
  wire       [31:0]   fixTo_367_dout;
  wire       [15:0]   fixTo_368_dout;
  wire       [15:0]   fixTo_369_dout;
  wire       [15:0]   fixTo_370_dout;
  wire       [15:0]   fixTo_371_dout;
  wire       [31:0]   fixTo_372_dout;
  wire       [31:0]   fixTo_373_dout;
  wire       [15:0]   fixTo_374_dout;
  wire       [15:0]   fixTo_375_dout;
  wire       [15:0]   fixTo_376_dout;
  wire       [15:0]   fixTo_377_dout;
  wire       [31:0]   fixTo_378_dout;
  wire       [31:0]   fixTo_379_dout;
  wire       [15:0]   fixTo_380_dout;
  wire       [15:0]   fixTo_381_dout;
  wire       [15:0]   fixTo_382_dout;
  wire       [15:0]   fixTo_383_dout;
  wire       [31:0]   fixTo_384_dout;
  wire       [31:0]   fixTo_385_dout;
  wire       [15:0]   fixTo_386_dout;
  wire       [15:0]   fixTo_387_dout;
  wire       [15:0]   fixTo_388_dout;
  wire       [15:0]   fixTo_389_dout;
  wire       [31:0]   fixTo_390_dout;
  wire       [31:0]   fixTo_391_dout;
  wire       [15:0]   fixTo_392_dout;
  wire       [15:0]   fixTo_393_dout;
  wire       [15:0]   fixTo_394_dout;
  wire       [15:0]   fixTo_395_dout;
  wire       [31:0]   fixTo_396_dout;
  wire       [31:0]   fixTo_397_dout;
  wire       [15:0]   fixTo_398_dout;
  wire       [15:0]   fixTo_399_dout;
  wire       [15:0]   fixTo_400_dout;
  wire       [15:0]   fixTo_401_dout;
  wire       [31:0]   fixTo_402_dout;
  wire       [31:0]   fixTo_403_dout;
  wire       [15:0]   fixTo_404_dout;
  wire       [15:0]   fixTo_405_dout;
  wire       [15:0]   fixTo_406_dout;
  wire       [15:0]   fixTo_407_dout;
  wire       [31:0]   fixTo_408_dout;
  wire       [31:0]   fixTo_409_dout;
  wire       [15:0]   fixTo_410_dout;
  wire       [15:0]   fixTo_411_dout;
  wire       [15:0]   fixTo_412_dout;
  wire       [15:0]   fixTo_413_dout;
  wire       [31:0]   fixTo_414_dout;
  wire       [31:0]   fixTo_415_dout;
  wire       [15:0]   fixTo_416_dout;
  wire       [15:0]   fixTo_417_dout;
  wire       [15:0]   fixTo_418_dout;
  wire       [15:0]   fixTo_419_dout;
  wire       [31:0]   fixTo_420_dout;
  wire       [31:0]   fixTo_421_dout;
  wire       [15:0]   fixTo_422_dout;
  wire       [15:0]   fixTo_423_dout;
  wire       [15:0]   fixTo_424_dout;
  wire       [15:0]   fixTo_425_dout;
  wire       [31:0]   fixTo_426_dout;
  wire       [31:0]   fixTo_427_dout;
  wire       [15:0]   fixTo_428_dout;
  wire       [15:0]   fixTo_429_dout;
  wire       [15:0]   fixTo_430_dout;
  wire       [15:0]   fixTo_431_dout;
  wire       [31:0]   fixTo_432_dout;
  wire       [31:0]   fixTo_433_dout;
  wire       [15:0]   fixTo_434_dout;
  wire       [15:0]   fixTo_435_dout;
  wire       [15:0]   fixTo_436_dout;
  wire       [15:0]   fixTo_437_dout;
  wire       [31:0]   fixTo_438_dout;
  wire       [31:0]   fixTo_439_dout;
  wire       [15:0]   fixTo_440_dout;
  wire       [15:0]   fixTo_441_dout;
  wire       [15:0]   fixTo_442_dout;
  wire       [15:0]   fixTo_443_dout;
  wire       [31:0]   fixTo_444_dout;
  wire       [31:0]   fixTo_445_dout;
  wire       [15:0]   fixTo_446_dout;
  wire       [15:0]   fixTo_447_dout;
  wire       [15:0]   fixTo_448_dout;
  wire       [15:0]   fixTo_449_dout;
  wire       [31:0]   fixTo_450_dout;
  wire       [31:0]   fixTo_451_dout;
  wire       [15:0]   fixTo_452_dout;
  wire       [15:0]   fixTo_453_dout;
  wire       [15:0]   fixTo_454_dout;
  wire       [15:0]   fixTo_455_dout;
  wire       [31:0]   fixTo_456_dout;
  wire       [31:0]   fixTo_457_dout;
  wire       [15:0]   fixTo_458_dout;
  wire       [15:0]   fixTo_459_dout;
  wire       [15:0]   fixTo_460_dout;
  wire       [15:0]   fixTo_461_dout;
  wire       [31:0]   fixTo_462_dout;
  wire       [31:0]   fixTo_463_dout;
  wire       [15:0]   fixTo_464_dout;
  wire       [15:0]   fixTo_465_dout;
  wire       [15:0]   fixTo_466_dout;
  wire       [15:0]   fixTo_467_dout;
  wire       [31:0]   fixTo_468_dout;
  wire       [31:0]   fixTo_469_dout;
  wire       [15:0]   fixTo_470_dout;
  wire       [15:0]   fixTo_471_dout;
  wire       [15:0]   fixTo_472_dout;
  wire       [15:0]   fixTo_473_dout;
  wire       [31:0]   fixTo_474_dout;
  wire       [31:0]   fixTo_475_dout;
  wire       [15:0]   fixTo_476_dout;
  wire       [15:0]   fixTo_477_dout;
  wire       [15:0]   fixTo_478_dout;
  wire       [15:0]   fixTo_479_dout;
  wire       [0:0]    _zz_881;
  wire       [2:0]    _zz_882;
  wire       [15:0]   _zz_883;
  wire       [31:0]   _zz_884;
  wire       [31:0]   _zz_885;
  wire       [15:0]   _zz_886;
  wire       [31:0]   _zz_887;
  wire       [31:0]   _zz_888;
  wire       [31:0]   _zz_889;
  wire       [15:0]   _zz_890;
  wire       [31:0]   _zz_891;
  wire       [31:0]   _zz_892;
  wire       [31:0]   _zz_893;
  wire       [31:0]   _zz_894;
  wire       [31:0]   _zz_895;
  wire       [31:0]   _zz_896;
  wire       [23:0]   _zz_897;
  wire       [31:0]   _zz_898;
  wire       [15:0]   _zz_899;
  wire       [31:0]   _zz_900;
  wire       [31:0]   _zz_901;
  wire       [31:0]   _zz_902;
  wire       [31:0]   _zz_903;
  wire       [31:0]   _zz_904;
  wire       [23:0]   _zz_905;
  wire       [31:0]   _zz_906;
  wire       [15:0]   _zz_907;
  wire       [31:0]   _zz_908;
  wire       [31:0]   _zz_909;
  wire       [31:0]   _zz_910;
  wire       [31:0]   _zz_911;
  wire       [31:0]   _zz_912;
  wire       [23:0]   _zz_913;
  wire       [31:0]   _zz_914;
  wire       [15:0]   _zz_915;
  wire       [31:0]   _zz_916;
  wire       [31:0]   _zz_917;
  wire       [31:0]   _zz_918;
  wire       [31:0]   _zz_919;
  wire       [31:0]   _zz_920;
  wire       [23:0]   _zz_921;
  wire       [31:0]   _zz_922;
  wire       [15:0]   _zz_923;
  wire       [15:0]   _zz_924;
  wire       [31:0]   _zz_925;
  wire       [31:0]   _zz_926;
  wire       [15:0]   _zz_927;
  wire       [31:0]   _zz_928;
  wire       [31:0]   _zz_929;
  wire       [31:0]   _zz_930;
  wire       [15:0]   _zz_931;
  wire       [31:0]   _zz_932;
  wire       [31:0]   _zz_933;
  wire       [31:0]   _zz_934;
  wire       [31:0]   _zz_935;
  wire       [31:0]   _zz_936;
  wire       [31:0]   _zz_937;
  wire       [23:0]   _zz_938;
  wire       [31:0]   _zz_939;
  wire       [15:0]   _zz_940;
  wire       [31:0]   _zz_941;
  wire       [31:0]   _zz_942;
  wire       [31:0]   _zz_943;
  wire       [31:0]   _zz_944;
  wire       [31:0]   _zz_945;
  wire       [23:0]   _zz_946;
  wire       [31:0]   _zz_947;
  wire       [15:0]   _zz_948;
  wire       [31:0]   _zz_949;
  wire       [31:0]   _zz_950;
  wire       [31:0]   _zz_951;
  wire       [31:0]   _zz_952;
  wire       [31:0]   _zz_953;
  wire       [23:0]   _zz_954;
  wire       [31:0]   _zz_955;
  wire       [15:0]   _zz_956;
  wire       [31:0]   _zz_957;
  wire       [31:0]   _zz_958;
  wire       [31:0]   _zz_959;
  wire       [31:0]   _zz_960;
  wire       [31:0]   _zz_961;
  wire       [23:0]   _zz_962;
  wire       [31:0]   _zz_963;
  wire       [15:0]   _zz_964;
  wire       [15:0]   _zz_965;
  wire       [31:0]   _zz_966;
  wire       [31:0]   _zz_967;
  wire       [15:0]   _zz_968;
  wire       [31:0]   _zz_969;
  wire       [31:0]   _zz_970;
  wire       [31:0]   _zz_971;
  wire       [15:0]   _zz_972;
  wire       [31:0]   _zz_973;
  wire       [31:0]   _zz_974;
  wire       [31:0]   _zz_975;
  wire       [31:0]   _zz_976;
  wire       [31:0]   _zz_977;
  wire       [31:0]   _zz_978;
  wire       [23:0]   _zz_979;
  wire       [31:0]   _zz_980;
  wire       [15:0]   _zz_981;
  wire       [31:0]   _zz_982;
  wire       [31:0]   _zz_983;
  wire       [31:0]   _zz_984;
  wire       [31:0]   _zz_985;
  wire       [31:0]   _zz_986;
  wire       [23:0]   _zz_987;
  wire       [31:0]   _zz_988;
  wire       [15:0]   _zz_989;
  wire       [31:0]   _zz_990;
  wire       [31:0]   _zz_991;
  wire       [31:0]   _zz_992;
  wire       [31:0]   _zz_993;
  wire       [31:0]   _zz_994;
  wire       [23:0]   _zz_995;
  wire       [31:0]   _zz_996;
  wire       [15:0]   _zz_997;
  wire       [31:0]   _zz_998;
  wire       [31:0]   _zz_999;
  wire       [31:0]   _zz_1000;
  wire       [31:0]   _zz_1001;
  wire       [31:0]   _zz_1002;
  wire       [23:0]   _zz_1003;
  wire       [31:0]   _zz_1004;
  wire       [15:0]   _zz_1005;
  wire       [15:0]   _zz_1006;
  wire       [31:0]   _zz_1007;
  wire       [31:0]   _zz_1008;
  wire       [15:0]   _zz_1009;
  wire       [31:0]   _zz_1010;
  wire       [31:0]   _zz_1011;
  wire       [31:0]   _zz_1012;
  wire       [15:0]   _zz_1013;
  wire       [31:0]   _zz_1014;
  wire       [31:0]   _zz_1015;
  wire       [31:0]   _zz_1016;
  wire       [31:0]   _zz_1017;
  wire       [31:0]   _zz_1018;
  wire       [31:0]   _zz_1019;
  wire       [23:0]   _zz_1020;
  wire       [31:0]   _zz_1021;
  wire       [15:0]   _zz_1022;
  wire       [31:0]   _zz_1023;
  wire       [31:0]   _zz_1024;
  wire       [31:0]   _zz_1025;
  wire       [31:0]   _zz_1026;
  wire       [31:0]   _zz_1027;
  wire       [23:0]   _zz_1028;
  wire       [31:0]   _zz_1029;
  wire       [15:0]   _zz_1030;
  wire       [31:0]   _zz_1031;
  wire       [31:0]   _zz_1032;
  wire       [31:0]   _zz_1033;
  wire       [31:0]   _zz_1034;
  wire       [31:0]   _zz_1035;
  wire       [23:0]   _zz_1036;
  wire       [31:0]   _zz_1037;
  wire       [15:0]   _zz_1038;
  wire       [31:0]   _zz_1039;
  wire       [31:0]   _zz_1040;
  wire       [31:0]   _zz_1041;
  wire       [31:0]   _zz_1042;
  wire       [31:0]   _zz_1043;
  wire       [23:0]   _zz_1044;
  wire       [31:0]   _zz_1045;
  wire       [15:0]   _zz_1046;
  wire       [15:0]   _zz_1047;
  wire       [31:0]   _zz_1048;
  wire       [31:0]   _zz_1049;
  wire       [15:0]   _zz_1050;
  wire       [31:0]   _zz_1051;
  wire       [31:0]   _zz_1052;
  wire       [31:0]   _zz_1053;
  wire       [15:0]   _zz_1054;
  wire       [31:0]   _zz_1055;
  wire       [31:0]   _zz_1056;
  wire       [31:0]   _zz_1057;
  wire       [31:0]   _zz_1058;
  wire       [31:0]   _zz_1059;
  wire       [31:0]   _zz_1060;
  wire       [23:0]   _zz_1061;
  wire       [31:0]   _zz_1062;
  wire       [15:0]   _zz_1063;
  wire       [31:0]   _zz_1064;
  wire       [31:0]   _zz_1065;
  wire       [31:0]   _zz_1066;
  wire       [31:0]   _zz_1067;
  wire       [31:0]   _zz_1068;
  wire       [23:0]   _zz_1069;
  wire       [31:0]   _zz_1070;
  wire       [15:0]   _zz_1071;
  wire       [31:0]   _zz_1072;
  wire       [31:0]   _zz_1073;
  wire       [31:0]   _zz_1074;
  wire       [31:0]   _zz_1075;
  wire       [31:0]   _zz_1076;
  wire       [23:0]   _zz_1077;
  wire       [31:0]   _zz_1078;
  wire       [15:0]   _zz_1079;
  wire       [31:0]   _zz_1080;
  wire       [31:0]   _zz_1081;
  wire       [31:0]   _zz_1082;
  wire       [31:0]   _zz_1083;
  wire       [31:0]   _zz_1084;
  wire       [23:0]   _zz_1085;
  wire       [31:0]   _zz_1086;
  wire       [15:0]   _zz_1087;
  wire       [15:0]   _zz_1088;
  wire       [31:0]   _zz_1089;
  wire       [31:0]   _zz_1090;
  wire       [15:0]   _zz_1091;
  wire       [31:0]   _zz_1092;
  wire       [31:0]   _zz_1093;
  wire       [31:0]   _zz_1094;
  wire       [15:0]   _zz_1095;
  wire       [31:0]   _zz_1096;
  wire       [31:0]   _zz_1097;
  wire       [31:0]   _zz_1098;
  wire       [31:0]   _zz_1099;
  wire       [31:0]   _zz_1100;
  wire       [31:0]   _zz_1101;
  wire       [23:0]   _zz_1102;
  wire       [31:0]   _zz_1103;
  wire       [15:0]   _zz_1104;
  wire       [31:0]   _zz_1105;
  wire       [31:0]   _zz_1106;
  wire       [31:0]   _zz_1107;
  wire       [31:0]   _zz_1108;
  wire       [31:0]   _zz_1109;
  wire       [23:0]   _zz_1110;
  wire       [31:0]   _zz_1111;
  wire       [15:0]   _zz_1112;
  wire       [31:0]   _zz_1113;
  wire       [31:0]   _zz_1114;
  wire       [31:0]   _zz_1115;
  wire       [31:0]   _zz_1116;
  wire       [31:0]   _zz_1117;
  wire       [23:0]   _zz_1118;
  wire       [31:0]   _zz_1119;
  wire       [15:0]   _zz_1120;
  wire       [31:0]   _zz_1121;
  wire       [31:0]   _zz_1122;
  wire       [31:0]   _zz_1123;
  wire       [31:0]   _zz_1124;
  wire       [31:0]   _zz_1125;
  wire       [23:0]   _zz_1126;
  wire       [31:0]   _zz_1127;
  wire       [15:0]   _zz_1128;
  wire       [15:0]   _zz_1129;
  wire       [31:0]   _zz_1130;
  wire       [31:0]   _zz_1131;
  wire       [15:0]   _zz_1132;
  wire       [31:0]   _zz_1133;
  wire       [31:0]   _zz_1134;
  wire       [31:0]   _zz_1135;
  wire       [15:0]   _zz_1136;
  wire       [31:0]   _zz_1137;
  wire       [31:0]   _zz_1138;
  wire       [31:0]   _zz_1139;
  wire       [31:0]   _zz_1140;
  wire       [31:0]   _zz_1141;
  wire       [31:0]   _zz_1142;
  wire       [23:0]   _zz_1143;
  wire       [31:0]   _zz_1144;
  wire       [15:0]   _zz_1145;
  wire       [31:0]   _zz_1146;
  wire       [31:0]   _zz_1147;
  wire       [31:0]   _zz_1148;
  wire       [31:0]   _zz_1149;
  wire       [31:0]   _zz_1150;
  wire       [23:0]   _zz_1151;
  wire       [31:0]   _zz_1152;
  wire       [15:0]   _zz_1153;
  wire       [31:0]   _zz_1154;
  wire       [31:0]   _zz_1155;
  wire       [31:0]   _zz_1156;
  wire       [31:0]   _zz_1157;
  wire       [31:0]   _zz_1158;
  wire       [23:0]   _zz_1159;
  wire       [31:0]   _zz_1160;
  wire       [15:0]   _zz_1161;
  wire       [31:0]   _zz_1162;
  wire       [31:0]   _zz_1163;
  wire       [31:0]   _zz_1164;
  wire       [31:0]   _zz_1165;
  wire       [31:0]   _zz_1166;
  wire       [23:0]   _zz_1167;
  wire       [31:0]   _zz_1168;
  wire       [15:0]   _zz_1169;
  wire       [15:0]   _zz_1170;
  wire       [31:0]   _zz_1171;
  wire       [31:0]   _zz_1172;
  wire       [15:0]   _zz_1173;
  wire       [31:0]   _zz_1174;
  wire       [31:0]   _zz_1175;
  wire       [31:0]   _zz_1176;
  wire       [15:0]   _zz_1177;
  wire       [31:0]   _zz_1178;
  wire       [31:0]   _zz_1179;
  wire       [31:0]   _zz_1180;
  wire       [31:0]   _zz_1181;
  wire       [31:0]   _zz_1182;
  wire       [31:0]   _zz_1183;
  wire       [23:0]   _zz_1184;
  wire       [31:0]   _zz_1185;
  wire       [15:0]   _zz_1186;
  wire       [31:0]   _zz_1187;
  wire       [31:0]   _zz_1188;
  wire       [31:0]   _zz_1189;
  wire       [31:0]   _zz_1190;
  wire       [31:0]   _zz_1191;
  wire       [23:0]   _zz_1192;
  wire       [31:0]   _zz_1193;
  wire       [15:0]   _zz_1194;
  wire       [31:0]   _zz_1195;
  wire       [31:0]   _zz_1196;
  wire       [31:0]   _zz_1197;
  wire       [31:0]   _zz_1198;
  wire       [31:0]   _zz_1199;
  wire       [23:0]   _zz_1200;
  wire       [31:0]   _zz_1201;
  wire       [15:0]   _zz_1202;
  wire       [31:0]   _zz_1203;
  wire       [31:0]   _zz_1204;
  wire       [31:0]   _zz_1205;
  wire       [31:0]   _zz_1206;
  wire       [31:0]   _zz_1207;
  wire       [23:0]   _zz_1208;
  wire       [31:0]   _zz_1209;
  wire       [15:0]   _zz_1210;
  wire       [15:0]   _zz_1211;
  wire       [31:0]   _zz_1212;
  wire       [31:0]   _zz_1213;
  wire       [15:0]   _zz_1214;
  wire       [31:0]   _zz_1215;
  wire       [31:0]   _zz_1216;
  wire       [31:0]   _zz_1217;
  wire       [15:0]   _zz_1218;
  wire       [31:0]   _zz_1219;
  wire       [31:0]   _zz_1220;
  wire       [31:0]   _zz_1221;
  wire       [31:0]   _zz_1222;
  wire       [31:0]   _zz_1223;
  wire       [31:0]   _zz_1224;
  wire       [23:0]   _zz_1225;
  wire       [31:0]   _zz_1226;
  wire       [15:0]   _zz_1227;
  wire       [31:0]   _zz_1228;
  wire       [31:0]   _zz_1229;
  wire       [31:0]   _zz_1230;
  wire       [31:0]   _zz_1231;
  wire       [31:0]   _zz_1232;
  wire       [23:0]   _zz_1233;
  wire       [31:0]   _zz_1234;
  wire       [15:0]   _zz_1235;
  wire       [31:0]   _zz_1236;
  wire       [31:0]   _zz_1237;
  wire       [31:0]   _zz_1238;
  wire       [31:0]   _zz_1239;
  wire       [31:0]   _zz_1240;
  wire       [23:0]   _zz_1241;
  wire       [31:0]   _zz_1242;
  wire       [15:0]   _zz_1243;
  wire       [31:0]   _zz_1244;
  wire       [31:0]   _zz_1245;
  wire       [31:0]   _zz_1246;
  wire       [31:0]   _zz_1247;
  wire       [31:0]   _zz_1248;
  wire       [23:0]   _zz_1249;
  wire       [31:0]   _zz_1250;
  wire       [15:0]   _zz_1251;
  wire       [15:0]   _zz_1252;
  wire       [31:0]   _zz_1253;
  wire       [31:0]   _zz_1254;
  wire       [15:0]   _zz_1255;
  wire       [31:0]   _zz_1256;
  wire       [31:0]   _zz_1257;
  wire       [31:0]   _zz_1258;
  wire       [15:0]   _zz_1259;
  wire       [31:0]   _zz_1260;
  wire       [31:0]   _zz_1261;
  wire       [31:0]   _zz_1262;
  wire       [31:0]   _zz_1263;
  wire       [31:0]   _zz_1264;
  wire       [31:0]   _zz_1265;
  wire       [23:0]   _zz_1266;
  wire       [31:0]   _zz_1267;
  wire       [15:0]   _zz_1268;
  wire       [31:0]   _zz_1269;
  wire       [31:0]   _zz_1270;
  wire       [31:0]   _zz_1271;
  wire       [31:0]   _zz_1272;
  wire       [31:0]   _zz_1273;
  wire       [23:0]   _zz_1274;
  wire       [31:0]   _zz_1275;
  wire       [15:0]   _zz_1276;
  wire       [31:0]   _zz_1277;
  wire       [31:0]   _zz_1278;
  wire       [31:0]   _zz_1279;
  wire       [31:0]   _zz_1280;
  wire       [31:0]   _zz_1281;
  wire       [23:0]   _zz_1282;
  wire       [31:0]   _zz_1283;
  wire       [15:0]   _zz_1284;
  wire       [31:0]   _zz_1285;
  wire       [31:0]   _zz_1286;
  wire       [31:0]   _zz_1287;
  wire       [31:0]   _zz_1288;
  wire       [31:0]   _zz_1289;
  wire       [23:0]   _zz_1290;
  wire       [31:0]   _zz_1291;
  wire       [15:0]   _zz_1292;
  wire       [15:0]   _zz_1293;
  wire       [31:0]   _zz_1294;
  wire       [31:0]   _zz_1295;
  wire       [15:0]   _zz_1296;
  wire       [31:0]   _zz_1297;
  wire       [31:0]   _zz_1298;
  wire       [31:0]   _zz_1299;
  wire       [15:0]   _zz_1300;
  wire       [31:0]   _zz_1301;
  wire       [31:0]   _zz_1302;
  wire       [31:0]   _zz_1303;
  wire       [31:0]   _zz_1304;
  wire       [31:0]   _zz_1305;
  wire       [31:0]   _zz_1306;
  wire       [23:0]   _zz_1307;
  wire       [31:0]   _zz_1308;
  wire       [15:0]   _zz_1309;
  wire       [31:0]   _zz_1310;
  wire       [31:0]   _zz_1311;
  wire       [31:0]   _zz_1312;
  wire       [31:0]   _zz_1313;
  wire       [31:0]   _zz_1314;
  wire       [23:0]   _zz_1315;
  wire       [31:0]   _zz_1316;
  wire       [15:0]   _zz_1317;
  wire       [31:0]   _zz_1318;
  wire       [31:0]   _zz_1319;
  wire       [31:0]   _zz_1320;
  wire       [31:0]   _zz_1321;
  wire       [31:0]   _zz_1322;
  wire       [23:0]   _zz_1323;
  wire       [31:0]   _zz_1324;
  wire       [15:0]   _zz_1325;
  wire       [31:0]   _zz_1326;
  wire       [31:0]   _zz_1327;
  wire       [31:0]   _zz_1328;
  wire       [31:0]   _zz_1329;
  wire       [31:0]   _zz_1330;
  wire       [23:0]   _zz_1331;
  wire       [31:0]   _zz_1332;
  wire       [15:0]   _zz_1333;
  wire       [15:0]   _zz_1334;
  wire       [31:0]   _zz_1335;
  wire       [31:0]   _zz_1336;
  wire       [15:0]   _zz_1337;
  wire       [31:0]   _zz_1338;
  wire       [31:0]   _zz_1339;
  wire       [31:0]   _zz_1340;
  wire       [15:0]   _zz_1341;
  wire       [31:0]   _zz_1342;
  wire       [31:0]   _zz_1343;
  wire       [31:0]   _zz_1344;
  wire       [31:0]   _zz_1345;
  wire       [31:0]   _zz_1346;
  wire       [31:0]   _zz_1347;
  wire       [23:0]   _zz_1348;
  wire       [31:0]   _zz_1349;
  wire       [15:0]   _zz_1350;
  wire       [31:0]   _zz_1351;
  wire       [31:0]   _zz_1352;
  wire       [31:0]   _zz_1353;
  wire       [31:0]   _zz_1354;
  wire       [31:0]   _zz_1355;
  wire       [23:0]   _zz_1356;
  wire       [31:0]   _zz_1357;
  wire       [15:0]   _zz_1358;
  wire       [31:0]   _zz_1359;
  wire       [31:0]   _zz_1360;
  wire       [31:0]   _zz_1361;
  wire       [31:0]   _zz_1362;
  wire       [31:0]   _zz_1363;
  wire       [23:0]   _zz_1364;
  wire       [31:0]   _zz_1365;
  wire       [15:0]   _zz_1366;
  wire       [31:0]   _zz_1367;
  wire       [31:0]   _zz_1368;
  wire       [31:0]   _zz_1369;
  wire       [31:0]   _zz_1370;
  wire       [31:0]   _zz_1371;
  wire       [23:0]   _zz_1372;
  wire       [31:0]   _zz_1373;
  wire       [15:0]   _zz_1374;
  wire       [15:0]   _zz_1375;
  wire       [31:0]   _zz_1376;
  wire       [31:0]   _zz_1377;
  wire       [15:0]   _zz_1378;
  wire       [31:0]   _zz_1379;
  wire       [31:0]   _zz_1380;
  wire       [31:0]   _zz_1381;
  wire       [15:0]   _zz_1382;
  wire       [31:0]   _zz_1383;
  wire       [31:0]   _zz_1384;
  wire       [31:0]   _zz_1385;
  wire       [31:0]   _zz_1386;
  wire       [31:0]   _zz_1387;
  wire       [31:0]   _zz_1388;
  wire       [23:0]   _zz_1389;
  wire       [31:0]   _zz_1390;
  wire       [15:0]   _zz_1391;
  wire       [31:0]   _zz_1392;
  wire       [31:0]   _zz_1393;
  wire       [31:0]   _zz_1394;
  wire       [31:0]   _zz_1395;
  wire       [31:0]   _zz_1396;
  wire       [23:0]   _zz_1397;
  wire       [31:0]   _zz_1398;
  wire       [15:0]   _zz_1399;
  wire       [31:0]   _zz_1400;
  wire       [31:0]   _zz_1401;
  wire       [31:0]   _zz_1402;
  wire       [31:0]   _zz_1403;
  wire       [31:0]   _zz_1404;
  wire       [23:0]   _zz_1405;
  wire       [31:0]   _zz_1406;
  wire       [15:0]   _zz_1407;
  wire       [31:0]   _zz_1408;
  wire       [31:0]   _zz_1409;
  wire       [31:0]   _zz_1410;
  wire       [31:0]   _zz_1411;
  wire       [31:0]   _zz_1412;
  wire       [23:0]   _zz_1413;
  wire       [31:0]   _zz_1414;
  wire       [15:0]   _zz_1415;
  wire       [15:0]   _zz_1416;
  wire       [31:0]   _zz_1417;
  wire       [31:0]   _zz_1418;
  wire       [15:0]   _zz_1419;
  wire       [31:0]   _zz_1420;
  wire       [31:0]   _zz_1421;
  wire       [31:0]   _zz_1422;
  wire       [15:0]   _zz_1423;
  wire       [31:0]   _zz_1424;
  wire       [31:0]   _zz_1425;
  wire       [31:0]   _zz_1426;
  wire       [31:0]   _zz_1427;
  wire       [31:0]   _zz_1428;
  wire       [31:0]   _zz_1429;
  wire       [23:0]   _zz_1430;
  wire       [31:0]   _zz_1431;
  wire       [15:0]   _zz_1432;
  wire       [31:0]   _zz_1433;
  wire       [31:0]   _zz_1434;
  wire       [31:0]   _zz_1435;
  wire       [31:0]   _zz_1436;
  wire       [31:0]   _zz_1437;
  wire       [23:0]   _zz_1438;
  wire       [31:0]   _zz_1439;
  wire       [15:0]   _zz_1440;
  wire       [31:0]   _zz_1441;
  wire       [31:0]   _zz_1442;
  wire       [31:0]   _zz_1443;
  wire       [31:0]   _zz_1444;
  wire       [31:0]   _zz_1445;
  wire       [23:0]   _zz_1446;
  wire       [31:0]   _zz_1447;
  wire       [15:0]   _zz_1448;
  wire       [31:0]   _zz_1449;
  wire       [31:0]   _zz_1450;
  wire       [31:0]   _zz_1451;
  wire       [31:0]   _zz_1452;
  wire       [31:0]   _zz_1453;
  wire       [23:0]   _zz_1454;
  wire       [31:0]   _zz_1455;
  wire       [15:0]   _zz_1456;
  wire       [15:0]   _zz_1457;
  wire       [31:0]   _zz_1458;
  wire       [31:0]   _zz_1459;
  wire       [15:0]   _zz_1460;
  wire       [31:0]   _zz_1461;
  wire       [31:0]   _zz_1462;
  wire       [31:0]   _zz_1463;
  wire       [15:0]   _zz_1464;
  wire       [31:0]   _zz_1465;
  wire       [31:0]   _zz_1466;
  wire       [31:0]   _zz_1467;
  wire       [31:0]   _zz_1468;
  wire       [31:0]   _zz_1469;
  wire       [31:0]   _zz_1470;
  wire       [23:0]   _zz_1471;
  wire       [31:0]   _zz_1472;
  wire       [15:0]   _zz_1473;
  wire       [31:0]   _zz_1474;
  wire       [31:0]   _zz_1475;
  wire       [31:0]   _zz_1476;
  wire       [31:0]   _zz_1477;
  wire       [31:0]   _zz_1478;
  wire       [23:0]   _zz_1479;
  wire       [31:0]   _zz_1480;
  wire       [15:0]   _zz_1481;
  wire       [31:0]   _zz_1482;
  wire       [31:0]   _zz_1483;
  wire       [31:0]   _zz_1484;
  wire       [31:0]   _zz_1485;
  wire       [31:0]   _zz_1486;
  wire       [23:0]   _zz_1487;
  wire       [31:0]   _zz_1488;
  wire       [15:0]   _zz_1489;
  wire       [31:0]   _zz_1490;
  wire       [31:0]   _zz_1491;
  wire       [31:0]   _zz_1492;
  wire       [31:0]   _zz_1493;
  wire       [31:0]   _zz_1494;
  wire       [23:0]   _zz_1495;
  wire       [31:0]   _zz_1496;
  wire       [15:0]   _zz_1497;
  wire       [15:0]   _zz_1498;
  wire       [31:0]   _zz_1499;
  wire       [31:0]   _zz_1500;
  wire       [15:0]   _zz_1501;
  wire       [31:0]   _zz_1502;
  wire       [31:0]   _zz_1503;
  wire       [31:0]   _zz_1504;
  wire       [15:0]   _zz_1505;
  wire       [31:0]   _zz_1506;
  wire       [31:0]   _zz_1507;
  wire       [31:0]   _zz_1508;
  wire       [31:0]   _zz_1509;
  wire       [31:0]   _zz_1510;
  wire       [31:0]   _zz_1511;
  wire       [23:0]   _zz_1512;
  wire       [31:0]   _zz_1513;
  wire       [15:0]   _zz_1514;
  wire       [31:0]   _zz_1515;
  wire       [31:0]   _zz_1516;
  wire       [31:0]   _zz_1517;
  wire       [31:0]   _zz_1518;
  wire       [31:0]   _zz_1519;
  wire       [23:0]   _zz_1520;
  wire       [31:0]   _zz_1521;
  wire       [15:0]   _zz_1522;
  wire       [31:0]   _zz_1523;
  wire       [31:0]   _zz_1524;
  wire       [31:0]   _zz_1525;
  wire       [31:0]   _zz_1526;
  wire       [31:0]   _zz_1527;
  wire       [23:0]   _zz_1528;
  wire       [31:0]   _zz_1529;
  wire       [15:0]   _zz_1530;
  wire       [31:0]   _zz_1531;
  wire       [31:0]   _zz_1532;
  wire       [31:0]   _zz_1533;
  wire       [31:0]   _zz_1534;
  wire       [31:0]   _zz_1535;
  wire       [23:0]   _zz_1536;
  wire       [31:0]   _zz_1537;
  wire       [15:0]   _zz_1538;
  wire       [15:0]   _zz_1539;
  wire       [31:0]   _zz_1540;
  wire       [31:0]   _zz_1541;
  wire       [15:0]   _zz_1542;
  wire       [31:0]   _zz_1543;
  wire       [31:0]   _zz_1544;
  wire       [31:0]   _zz_1545;
  wire       [15:0]   _zz_1546;
  wire       [31:0]   _zz_1547;
  wire       [31:0]   _zz_1548;
  wire       [31:0]   _zz_1549;
  wire       [31:0]   _zz_1550;
  wire       [31:0]   _zz_1551;
  wire       [31:0]   _zz_1552;
  wire       [23:0]   _zz_1553;
  wire       [31:0]   _zz_1554;
  wire       [15:0]   _zz_1555;
  wire       [31:0]   _zz_1556;
  wire       [31:0]   _zz_1557;
  wire       [31:0]   _zz_1558;
  wire       [31:0]   _zz_1559;
  wire       [31:0]   _zz_1560;
  wire       [23:0]   _zz_1561;
  wire       [31:0]   _zz_1562;
  wire       [15:0]   _zz_1563;
  wire       [31:0]   _zz_1564;
  wire       [31:0]   _zz_1565;
  wire       [31:0]   _zz_1566;
  wire       [31:0]   _zz_1567;
  wire       [31:0]   _zz_1568;
  wire       [23:0]   _zz_1569;
  wire       [31:0]   _zz_1570;
  wire       [15:0]   _zz_1571;
  wire       [31:0]   _zz_1572;
  wire       [31:0]   _zz_1573;
  wire       [31:0]   _zz_1574;
  wire       [31:0]   _zz_1575;
  wire       [31:0]   _zz_1576;
  wire       [23:0]   _zz_1577;
  wire       [31:0]   _zz_1578;
  wire       [15:0]   _zz_1579;
  wire       [15:0]   _zz_1580;
  wire       [31:0]   _zz_1581;
  wire       [31:0]   _zz_1582;
  wire       [15:0]   _zz_1583;
  wire       [31:0]   _zz_1584;
  wire       [31:0]   _zz_1585;
  wire       [31:0]   _zz_1586;
  wire       [15:0]   _zz_1587;
  wire       [31:0]   _zz_1588;
  wire       [31:0]   _zz_1589;
  wire       [31:0]   _zz_1590;
  wire       [31:0]   _zz_1591;
  wire       [31:0]   _zz_1592;
  wire       [31:0]   _zz_1593;
  wire       [23:0]   _zz_1594;
  wire       [31:0]   _zz_1595;
  wire       [15:0]   _zz_1596;
  wire       [31:0]   _zz_1597;
  wire       [31:0]   _zz_1598;
  wire       [31:0]   _zz_1599;
  wire       [31:0]   _zz_1600;
  wire       [31:0]   _zz_1601;
  wire       [23:0]   _zz_1602;
  wire       [31:0]   _zz_1603;
  wire       [15:0]   _zz_1604;
  wire       [31:0]   _zz_1605;
  wire       [31:0]   _zz_1606;
  wire       [31:0]   _zz_1607;
  wire       [31:0]   _zz_1608;
  wire       [31:0]   _zz_1609;
  wire       [23:0]   _zz_1610;
  wire       [31:0]   _zz_1611;
  wire       [15:0]   _zz_1612;
  wire       [31:0]   _zz_1613;
  wire       [31:0]   _zz_1614;
  wire       [31:0]   _zz_1615;
  wire       [31:0]   _zz_1616;
  wire       [31:0]   _zz_1617;
  wire       [23:0]   _zz_1618;
  wire       [31:0]   _zz_1619;
  wire       [15:0]   _zz_1620;
  wire       [15:0]   _zz_1621;
  wire       [31:0]   _zz_1622;
  wire       [31:0]   _zz_1623;
  wire       [15:0]   _zz_1624;
  wire       [31:0]   _zz_1625;
  wire       [31:0]   _zz_1626;
  wire       [31:0]   _zz_1627;
  wire       [15:0]   _zz_1628;
  wire       [31:0]   _zz_1629;
  wire       [31:0]   _zz_1630;
  wire       [31:0]   _zz_1631;
  wire       [31:0]   _zz_1632;
  wire       [31:0]   _zz_1633;
  wire       [31:0]   _zz_1634;
  wire       [23:0]   _zz_1635;
  wire       [31:0]   _zz_1636;
  wire       [15:0]   _zz_1637;
  wire       [31:0]   _zz_1638;
  wire       [31:0]   _zz_1639;
  wire       [31:0]   _zz_1640;
  wire       [31:0]   _zz_1641;
  wire       [31:0]   _zz_1642;
  wire       [23:0]   _zz_1643;
  wire       [31:0]   _zz_1644;
  wire       [15:0]   _zz_1645;
  wire       [31:0]   _zz_1646;
  wire       [31:0]   _zz_1647;
  wire       [31:0]   _zz_1648;
  wire       [31:0]   _zz_1649;
  wire       [31:0]   _zz_1650;
  wire       [23:0]   _zz_1651;
  wire       [31:0]   _zz_1652;
  wire       [15:0]   _zz_1653;
  wire       [31:0]   _zz_1654;
  wire       [31:0]   _zz_1655;
  wire       [31:0]   _zz_1656;
  wire       [31:0]   _zz_1657;
  wire       [31:0]   _zz_1658;
  wire       [23:0]   _zz_1659;
  wire       [31:0]   _zz_1660;
  wire       [15:0]   _zz_1661;
  wire       [15:0]   _zz_1662;
  wire       [31:0]   _zz_1663;
  wire       [31:0]   _zz_1664;
  wire       [15:0]   _zz_1665;
  wire       [31:0]   _zz_1666;
  wire       [31:0]   _zz_1667;
  wire       [31:0]   _zz_1668;
  wire       [15:0]   _zz_1669;
  wire       [31:0]   _zz_1670;
  wire       [31:0]   _zz_1671;
  wire       [31:0]   _zz_1672;
  wire       [31:0]   _zz_1673;
  wire       [31:0]   _zz_1674;
  wire       [31:0]   _zz_1675;
  wire       [23:0]   _zz_1676;
  wire       [31:0]   _zz_1677;
  wire       [15:0]   _zz_1678;
  wire       [31:0]   _zz_1679;
  wire       [31:0]   _zz_1680;
  wire       [31:0]   _zz_1681;
  wire       [31:0]   _zz_1682;
  wire       [31:0]   _zz_1683;
  wire       [23:0]   _zz_1684;
  wire       [31:0]   _zz_1685;
  wire       [15:0]   _zz_1686;
  wire       [31:0]   _zz_1687;
  wire       [31:0]   _zz_1688;
  wire       [31:0]   _zz_1689;
  wire       [31:0]   _zz_1690;
  wire       [31:0]   _zz_1691;
  wire       [23:0]   _zz_1692;
  wire       [31:0]   _zz_1693;
  wire       [15:0]   _zz_1694;
  wire       [31:0]   _zz_1695;
  wire       [31:0]   _zz_1696;
  wire       [31:0]   _zz_1697;
  wire       [31:0]   _zz_1698;
  wire       [31:0]   _zz_1699;
  wire       [23:0]   _zz_1700;
  wire       [31:0]   _zz_1701;
  wire       [15:0]   _zz_1702;
  wire       [15:0]   _zz_1703;
  wire       [31:0]   _zz_1704;
  wire       [31:0]   _zz_1705;
  wire       [15:0]   _zz_1706;
  wire       [31:0]   _zz_1707;
  wire       [31:0]   _zz_1708;
  wire       [31:0]   _zz_1709;
  wire       [15:0]   _zz_1710;
  wire       [31:0]   _zz_1711;
  wire       [31:0]   _zz_1712;
  wire       [31:0]   _zz_1713;
  wire       [31:0]   _zz_1714;
  wire       [31:0]   _zz_1715;
  wire       [31:0]   _zz_1716;
  wire       [23:0]   _zz_1717;
  wire       [31:0]   _zz_1718;
  wire       [15:0]   _zz_1719;
  wire       [31:0]   _zz_1720;
  wire       [31:0]   _zz_1721;
  wire       [31:0]   _zz_1722;
  wire       [31:0]   _zz_1723;
  wire       [31:0]   _zz_1724;
  wire       [23:0]   _zz_1725;
  wire       [31:0]   _zz_1726;
  wire       [15:0]   _zz_1727;
  wire       [31:0]   _zz_1728;
  wire       [31:0]   _zz_1729;
  wire       [31:0]   _zz_1730;
  wire       [31:0]   _zz_1731;
  wire       [31:0]   _zz_1732;
  wire       [23:0]   _zz_1733;
  wire       [31:0]   _zz_1734;
  wire       [15:0]   _zz_1735;
  wire       [31:0]   _zz_1736;
  wire       [31:0]   _zz_1737;
  wire       [31:0]   _zz_1738;
  wire       [31:0]   _zz_1739;
  wire       [31:0]   _zz_1740;
  wire       [23:0]   _zz_1741;
  wire       [31:0]   _zz_1742;
  wire       [15:0]   _zz_1743;
  wire       [15:0]   _zz_1744;
  wire       [31:0]   _zz_1745;
  wire       [31:0]   _zz_1746;
  wire       [15:0]   _zz_1747;
  wire       [31:0]   _zz_1748;
  wire       [31:0]   _zz_1749;
  wire       [31:0]   _zz_1750;
  wire       [15:0]   _zz_1751;
  wire       [31:0]   _zz_1752;
  wire       [31:0]   _zz_1753;
  wire       [31:0]   _zz_1754;
  wire       [31:0]   _zz_1755;
  wire       [31:0]   _zz_1756;
  wire       [31:0]   _zz_1757;
  wire       [23:0]   _zz_1758;
  wire       [31:0]   _zz_1759;
  wire       [15:0]   _zz_1760;
  wire       [31:0]   _zz_1761;
  wire       [31:0]   _zz_1762;
  wire       [31:0]   _zz_1763;
  wire       [31:0]   _zz_1764;
  wire       [31:0]   _zz_1765;
  wire       [23:0]   _zz_1766;
  wire       [31:0]   _zz_1767;
  wire       [15:0]   _zz_1768;
  wire       [31:0]   _zz_1769;
  wire       [31:0]   _zz_1770;
  wire       [31:0]   _zz_1771;
  wire       [31:0]   _zz_1772;
  wire       [31:0]   _zz_1773;
  wire       [23:0]   _zz_1774;
  wire       [31:0]   _zz_1775;
  wire       [15:0]   _zz_1776;
  wire       [31:0]   _zz_1777;
  wire       [31:0]   _zz_1778;
  wire       [31:0]   _zz_1779;
  wire       [31:0]   _zz_1780;
  wire       [31:0]   _zz_1781;
  wire       [23:0]   _zz_1782;
  wire       [31:0]   _zz_1783;
  wire       [15:0]   _zz_1784;
  wire       [15:0]   _zz_1785;
  wire       [31:0]   _zz_1786;
  wire       [31:0]   _zz_1787;
  wire       [15:0]   _zz_1788;
  wire       [31:0]   _zz_1789;
  wire       [31:0]   _zz_1790;
  wire       [31:0]   _zz_1791;
  wire       [15:0]   _zz_1792;
  wire       [31:0]   _zz_1793;
  wire       [31:0]   _zz_1794;
  wire       [31:0]   _zz_1795;
  wire       [31:0]   _zz_1796;
  wire       [31:0]   _zz_1797;
  wire       [31:0]   _zz_1798;
  wire       [23:0]   _zz_1799;
  wire       [31:0]   _zz_1800;
  wire       [15:0]   _zz_1801;
  wire       [31:0]   _zz_1802;
  wire       [31:0]   _zz_1803;
  wire       [31:0]   _zz_1804;
  wire       [31:0]   _zz_1805;
  wire       [31:0]   _zz_1806;
  wire       [23:0]   _zz_1807;
  wire       [31:0]   _zz_1808;
  wire       [15:0]   _zz_1809;
  wire       [31:0]   _zz_1810;
  wire       [31:0]   _zz_1811;
  wire       [31:0]   _zz_1812;
  wire       [31:0]   _zz_1813;
  wire       [31:0]   _zz_1814;
  wire       [23:0]   _zz_1815;
  wire       [31:0]   _zz_1816;
  wire       [15:0]   _zz_1817;
  wire       [31:0]   _zz_1818;
  wire       [31:0]   _zz_1819;
  wire       [31:0]   _zz_1820;
  wire       [31:0]   _zz_1821;
  wire       [31:0]   _zz_1822;
  wire       [23:0]   _zz_1823;
  wire       [31:0]   _zz_1824;
  wire       [15:0]   _zz_1825;
  wire       [15:0]   _zz_1826;
  wire       [31:0]   _zz_1827;
  wire       [31:0]   _zz_1828;
  wire       [15:0]   _zz_1829;
  wire       [31:0]   _zz_1830;
  wire       [31:0]   _zz_1831;
  wire       [31:0]   _zz_1832;
  wire       [15:0]   _zz_1833;
  wire       [31:0]   _zz_1834;
  wire       [31:0]   _zz_1835;
  wire       [31:0]   _zz_1836;
  wire       [31:0]   _zz_1837;
  wire       [31:0]   _zz_1838;
  wire       [31:0]   _zz_1839;
  wire       [23:0]   _zz_1840;
  wire       [31:0]   _zz_1841;
  wire       [15:0]   _zz_1842;
  wire       [31:0]   _zz_1843;
  wire       [31:0]   _zz_1844;
  wire       [31:0]   _zz_1845;
  wire       [31:0]   _zz_1846;
  wire       [31:0]   _zz_1847;
  wire       [23:0]   _zz_1848;
  wire       [31:0]   _zz_1849;
  wire       [15:0]   _zz_1850;
  wire       [31:0]   _zz_1851;
  wire       [31:0]   _zz_1852;
  wire       [31:0]   _zz_1853;
  wire       [31:0]   _zz_1854;
  wire       [31:0]   _zz_1855;
  wire       [23:0]   _zz_1856;
  wire       [31:0]   _zz_1857;
  wire       [15:0]   _zz_1858;
  wire       [31:0]   _zz_1859;
  wire       [31:0]   _zz_1860;
  wire       [31:0]   _zz_1861;
  wire       [31:0]   _zz_1862;
  wire       [31:0]   _zz_1863;
  wire       [23:0]   _zz_1864;
  wire       [31:0]   _zz_1865;
  wire       [15:0]   _zz_1866;
  wire       [15:0]   _zz_1867;
  wire       [31:0]   _zz_1868;
  wire       [31:0]   _zz_1869;
  wire       [15:0]   _zz_1870;
  wire       [31:0]   _zz_1871;
  wire       [31:0]   _zz_1872;
  wire       [31:0]   _zz_1873;
  wire       [15:0]   _zz_1874;
  wire       [31:0]   _zz_1875;
  wire       [31:0]   _zz_1876;
  wire       [31:0]   _zz_1877;
  wire       [31:0]   _zz_1878;
  wire       [31:0]   _zz_1879;
  wire       [31:0]   _zz_1880;
  wire       [23:0]   _zz_1881;
  wire       [31:0]   _zz_1882;
  wire       [15:0]   _zz_1883;
  wire       [31:0]   _zz_1884;
  wire       [31:0]   _zz_1885;
  wire       [31:0]   _zz_1886;
  wire       [31:0]   _zz_1887;
  wire       [31:0]   _zz_1888;
  wire       [23:0]   _zz_1889;
  wire       [31:0]   _zz_1890;
  wire       [15:0]   _zz_1891;
  wire       [31:0]   _zz_1892;
  wire       [31:0]   _zz_1893;
  wire       [31:0]   _zz_1894;
  wire       [31:0]   _zz_1895;
  wire       [31:0]   _zz_1896;
  wire       [23:0]   _zz_1897;
  wire       [31:0]   _zz_1898;
  wire       [15:0]   _zz_1899;
  wire       [31:0]   _zz_1900;
  wire       [31:0]   _zz_1901;
  wire       [31:0]   _zz_1902;
  wire       [31:0]   _zz_1903;
  wire       [31:0]   _zz_1904;
  wire       [23:0]   _zz_1905;
  wire       [31:0]   _zz_1906;
  wire       [15:0]   _zz_1907;
  wire       [15:0]   _zz_1908;
  wire       [31:0]   _zz_1909;
  wire       [31:0]   _zz_1910;
  wire       [15:0]   _zz_1911;
  wire       [31:0]   _zz_1912;
  wire       [31:0]   _zz_1913;
  wire       [31:0]   _zz_1914;
  wire       [15:0]   _zz_1915;
  wire       [31:0]   _zz_1916;
  wire       [31:0]   _zz_1917;
  wire       [31:0]   _zz_1918;
  wire       [31:0]   _zz_1919;
  wire       [31:0]   _zz_1920;
  wire       [31:0]   _zz_1921;
  wire       [23:0]   _zz_1922;
  wire       [31:0]   _zz_1923;
  wire       [15:0]   _zz_1924;
  wire       [31:0]   _zz_1925;
  wire       [31:0]   _zz_1926;
  wire       [31:0]   _zz_1927;
  wire       [31:0]   _zz_1928;
  wire       [31:0]   _zz_1929;
  wire       [23:0]   _zz_1930;
  wire       [31:0]   _zz_1931;
  wire       [15:0]   _zz_1932;
  wire       [31:0]   _zz_1933;
  wire       [31:0]   _zz_1934;
  wire       [31:0]   _zz_1935;
  wire       [31:0]   _zz_1936;
  wire       [31:0]   _zz_1937;
  wire       [23:0]   _zz_1938;
  wire       [31:0]   _zz_1939;
  wire       [15:0]   _zz_1940;
  wire       [31:0]   _zz_1941;
  wire       [31:0]   _zz_1942;
  wire       [31:0]   _zz_1943;
  wire       [31:0]   _zz_1944;
  wire       [31:0]   _zz_1945;
  wire       [23:0]   _zz_1946;
  wire       [31:0]   _zz_1947;
  wire       [15:0]   _zz_1948;
  wire       [15:0]   _zz_1949;
  wire       [31:0]   _zz_1950;
  wire       [31:0]   _zz_1951;
  wire       [15:0]   _zz_1952;
  wire       [31:0]   _zz_1953;
  wire       [31:0]   _zz_1954;
  wire       [31:0]   _zz_1955;
  wire       [15:0]   _zz_1956;
  wire       [31:0]   _zz_1957;
  wire       [31:0]   _zz_1958;
  wire       [31:0]   _zz_1959;
  wire       [31:0]   _zz_1960;
  wire       [31:0]   _zz_1961;
  wire       [31:0]   _zz_1962;
  wire       [23:0]   _zz_1963;
  wire       [31:0]   _zz_1964;
  wire       [15:0]   _zz_1965;
  wire       [31:0]   _zz_1966;
  wire       [31:0]   _zz_1967;
  wire       [31:0]   _zz_1968;
  wire       [31:0]   _zz_1969;
  wire       [31:0]   _zz_1970;
  wire       [23:0]   _zz_1971;
  wire       [31:0]   _zz_1972;
  wire       [15:0]   _zz_1973;
  wire       [31:0]   _zz_1974;
  wire       [31:0]   _zz_1975;
  wire       [31:0]   _zz_1976;
  wire       [31:0]   _zz_1977;
  wire       [31:0]   _zz_1978;
  wire       [23:0]   _zz_1979;
  wire       [31:0]   _zz_1980;
  wire       [15:0]   _zz_1981;
  wire       [31:0]   _zz_1982;
  wire       [31:0]   _zz_1983;
  wire       [31:0]   _zz_1984;
  wire       [31:0]   _zz_1985;
  wire       [31:0]   _zz_1986;
  wire       [23:0]   _zz_1987;
  wire       [31:0]   _zz_1988;
  wire       [15:0]   _zz_1989;
  wire       [15:0]   _zz_1990;
  wire       [31:0]   _zz_1991;
  wire       [31:0]   _zz_1992;
  wire       [15:0]   _zz_1993;
  wire       [31:0]   _zz_1994;
  wire       [31:0]   _zz_1995;
  wire       [31:0]   _zz_1996;
  wire       [15:0]   _zz_1997;
  wire       [31:0]   _zz_1998;
  wire       [31:0]   _zz_1999;
  wire       [31:0]   _zz_2000;
  wire       [31:0]   _zz_2001;
  wire       [31:0]   _zz_2002;
  wire       [31:0]   _zz_2003;
  wire       [23:0]   _zz_2004;
  wire       [31:0]   _zz_2005;
  wire       [15:0]   _zz_2006;
  wire       [31:0]   _zz_2007;
  wire       [31:0]   _zz_2008;
  wire       [31:0]   _zz_2009;
  wire       [31:0]   _zz_2010;
  wire       [31:0]   _zz_2011;
  wire       [23:0]   _zz_2012;
  wire       [31:0]   _zz_2013;
  wire       [15:0]   _zz_2014;
  wire       [31:0]   _zz_2015;
  wire       [31:0]   _zz_2016;
  wire       [31:0]   _zz_2017;
  wire       [31:0]   _zz_2018;
  wire       [31:0]   _zz_2019;
  wire       [23:0]   _zz_2020;
  wire       [31:0]   _zz_2021;
  wire       [15:0]   _zz_2022;
  wire       [31:0]   _zz_2023;
  wire       [31:0]   _zz_2024;
  wire       [31:0]   _zz_2025;
  wire       [31:0]   _zz_2026;
  wire       [31:0]   _zz_2027;
  wire       [23:0]   _zz_2028;
  wire       [31:0]   _zz_2029;
  wire       [15:0]   _zz_2030;
  wire       [15:0]   _zz_2031;
  wire       [31:0]   _zz_2032;
  wire       [31:0]   _zz_2033;
  wire       [15:0]   _zz_2034;
  wire       [31:0]   _zz_2035;
  wire       [31:0]   _zz_2036;
  wire       [31:0]   _zz_2037;
  wire       [15:0]   _zz_2038;
  wire       [31:0]   _zz_2039;
  wire       [31:0]   _zz_2040;
  wire       [31:0]   _zz_2041;
  wire       [31:0]   _zz_2042;
  wire       [31:0]   _zz_2043;
  wire       [31:0]   _zz_2044;
  wire       [23:0]   _zz_2045;
  wire       [31:0]   _zz_2046;
  wire       [15:0]   _zz_2047;
  wire       [31:0]   _zz_2048;
  wire       [31:0]   _zz_2049;
  wire       [31:0]   _zz_2050;
  wire       [31:0]   _zz_2051;
  wire       [31:0]   _zz_2052;
  wire       [23:0]   _zz_2053;
  wire       [31:0]   _zz_2054;
  wire       [15:0]   _zz_2055;
  wire       [31:0]   _zz_2056;
  wire       [31:0]   _zz_2057;
  wire       [31:0]   _zz_2058;
  wire       [31:0]   _zz_2059;
  wire       [31:0]   _zz_2060;
  wire       [23:0]   _zz_2061;
  wire       [31:0]   _zz_2062;
  wire       [15:0]   _zz_2063;
  wire       [31:0]   _zz_2064;
  wire       [31:0]   _zz_2065;
  wire       [31:0]   _zz_2066;
  wire       [31:0]   _zz_2067;
  wire       [31:0]   _zz_2068;
  wire       [23:0]   _zz_2069;
  wire       [31:0]   _zz_2070;
  wire       [15:0]   _zz_2071;
  wire       [15:0]   _zz_2072;
  wire       [31:0]   _zz_2073;
  wire       [31:0]   _zz_2074;
  wire       [15:0]   _zz_2075;
  wire       [31:0]   _zz_2076;
  wire       [31:0]   _zz_2077;
  wire       [31:0]   _zz_2078;
  wire       [15:0]   _zz_2079;
  wire       [31:0]   _zz_2080;
  wire       [31:0]   _zz_2081;
  wire       [31:0]   _zz_2082;
  wire       [31:0]   _zz_2083;
  wire       [31:0]   _zz_2084;
  wire       [31:0]   _zz_2085;
  wire       [23:0]   _zz_2086;
  wire       [31:0]   _zz_2087;
  wire       [15:0]   _zz_2088;
  wire       [31:0]   _zz_2089;
  wire       [31:0]   _zz_2090;
  wire       [31:0]   _zz_2091;
  wire       [31:0]   _zz_2092;
  wire       [31:0]   _zz_2093;
  wire       [23:0]   _zz_2094;
  wire       [31:0]   _zz_2095;
  wire       [15:0]   _zz_2096;
  wire       [31:0]   _zz_2097;
  wire       [31:0]   _zz_2098;
  wire       [31:0]   _zz_2099;
  wire       [31:0]   _zz_2100;
  wire       [31:0]   _zz_2101;
  wire       [23:0]   _zz_2102;
  wire       [31:0]   _zz_2103;
  wire       [15:0]   _zz_2104;
  wire       [31:0]   _zz_2105;
  wire       [31:0]   _zz_2106;
  wire       [31:0]   _zz_2107;
  wire       [31:0]   _zz_2108;
  wire       [31:0]   _zz_2109;
  wire       [23:0]   _zz_2110;
  wire       [31:0]   _zz_2111;
  wire       [15:0]   _zz_2112;
  wire       [15:0]   _zz_2113;
  wire       [31:0]   _zz_2114;
  wire       [31:0]   _zz_2115;
  wire       [15:0]   _zz_2116;
  wire       [31:0]   _zz_2117;
  wire       [31:0]   _zz_2118;
  wire       [31:0]   _zz_2119;
  wire       [15:0]   _zz_2120;
  wire       [31:0]   _zz_2121;
  wire       [31:0]   _zz_2122;
  wire       [31:0]   _zz_2123;
  wire       [31:0]   _zz_2124;
  wire       [31:0]   _zz_2125;
  wire       [31:0]   _zz_2126;
  wire       [23:0]   _zz_2127;
  wire       [31:0]   _zz_2128;
  wire       [15:0]   _zz_2129;
  wire       [31:0]   _zz_2130;
  wire       [31:0]   _zz_2131;
  wire       [31:0]   _zz_2132;
  wire       [31:0]   _zz_2133;
  wire       [31:0]   _zz_2134;
  wire       [23:0]   _zz_2135;
  wire       [31:0]   _zz_2136;
  wire       [15:0]   _zz_2137;
  wire       [31:0]   _zz_2138;
  wire       [31:0]   _zz_2139;
  wire       [31:0]   _zz_2140;
  wire       [31:0]   _zz_2141;
  wire       [31:0]   _zz_2142;
  wire       [23:0]   _zz_2143;
  wire       [31:0]   _zz_2144;
  wire       [15:0]   _zz_2145;
  wire       [31:0]   _zz_2146;
  wire       [31:0]   _zz_2147;
  wire       [31:0]   _zz_2148;
  wire       [31:0]   _zz_2149;
  wire       [31:0]   _zz_2150;
  wire       [23:0]   _zz_2151;
  wire       [31:0]   _zz_2152;
  wire       [15:0]   _zz_2153;
  wire       [15:0]   _zz_2154;
  wire       [31:0]   _zz_2155;
  wire       [31:0]   _zz_2156;
  wire       [15:0]   _zz_2157;
  wire       [31:0]   _zz_2158;
  wire       [31:0]   _zz_2159;
  wire       [31:0]   _zz_2160;
  wire       [15:0]   _zz_2161;
  wire       [31:0]   _zz_2162;
  wire       [31:0]   _zz_2163;
  wire       [31:0]   _zz_2164;
  wire       [31:0]   _zz_2165;
  wire       [31:0]   _zz_2166;
  wire       [31:0]   _zz_2167;
  wire       [23:0]   _zz_2168;
  wire       [31:0]   _zz_2169;
  wire       [15:0]   _zz_2170;
  wire       [31:0]   _zz_2171;
  wire       [31:0]   _zz_2172;
  wire       [31:0]   _zz_2173;
  wire       [31:0]   _zz_2174;
  wire       [31:0]   _zz_2175;
  wire       [23:0]   _zz_2176;
  wire       [31:0]   _zz_2177;
  wire       [15:0]   _zz_2178;
  wire       [31:0]   _zz_2179;
  wire       [31:0]   _zz_2180;
  wire       [31:0]   _zz_2181;
  wire       [31:0]   _zz_2182;
  wire       [31:0]   _zz_2183;
  wire       [23:0]   _zz_2184;
  wire       [31:0]   _zz_2185;
  wire       [15:0]   _zz_2186;
  wire       [31:0]   _zz_2187;
  wire       [31:0]   _zz_2188;
  wire       [31:0]   _zz_2189;
  wire       [31:0]   _zz_2190;
  wire       [31:0]   _zz_2191;
  wire       [23:0]   _zz_2192;
  wire       [31:0]   _zz_2193;
  wire       [15:0]   _zz_2194;
  wire       [15:0]   _zz_2195;
  wire       [31:0]   _zz_2196;
  wire       [31:0]   _zz_2197;
  wire       [15:0]   _zz_2198;
  wire       [31:0]   _zz_2199;
  wire       [31:0]   _zz_2200;
  wire       [31:0]   _zz_2201;
  wire       [15:0]   _zz_2202;
  wire       [31:0]   _zz_2203;
  wire       [31:0]   _zz_2204;
  wire       [31:0]   _zz_2205;
  wire       [31:0]   _zz_2206;
  wire       [31:0]   _zz_2207;
  wire       [31:0]   _zz_2208;
  wire       [23:0]   _zz_2209;
  wire       [31:0]   _zz_2210;
  wire       [15:0]   _zz_2211;
  wire       [31:0]   _zz_2212;
  wire       [31:0]   _zz_2213;
  wire       [31:0]   _zz_2214;
  wire       [31:0]   _zz_2215;
  wire       [31:0]   _zz_2216;
  wire       [23:0]   _zz_2217;
  wire       [31:0]   _zz_2218;
  wire       [15:0]   _zz_2219;
  wire       [31:0]   _zz_2220;
  wire       [31:0]   _zz_2221;
  wire       [31:0]   _zz_2222;
  wire       [31:0]   _zz_2223;
  wire       [31:0]   _zz_2224;
  wire       [23:0]   _zz_2225;
  wire       [31:0]   _zz_2226;
  wire       [15:0]   _zz_2227;
  wire       [31:0]   _zz_2228;
  wire       [31:0]   _zz_2229;
  wire       [31:0]   _zz_2230;
  wire       [31:0]   _zz_2231;
  wire       [31:0]   _zz_2232;
  wire       [23:0]   _zz_2233;
  wire       [31:0]   _zz_2234;
  wire       [15:0]   _zz_2235;
  wire       [15:0]   _zz_2236;
  wire       [31:0]   _zz_2237;
  wire       [31:0]   _zz_2238;
  wire       [15:0]   _zz_2239;
  wire       [31:0]   _zz_2240;
  wire       [31:0]   _zz_2241;
  wire       [31:0]   _zz_2242;
  wire       [15:0]   _zz_2243;
  wire       [31:0]   _zz_2244;
  wire       [31:0]   _zz_2245;
  wire       [31:0]   _zz_2246;
  wire       [31:0]   _zz_2247;
  wire       [31:0]   _zz_2248;
  wire       [31:0]   _zz_2249;
  wire       [23:0]   _zz_2250;
  wire       [31:0]   _zz_2251;
  wire       [15:0]   _zz_2252;
  wire       [31:0]   _zz_2253;
  wire       [31:0]   _zz_2254;
  wire       [31:0]   _zz_2255;
  wire       [31:0]   _zz_2256;
  wire       [31:0]   _zz_2257;
  wire       [23:0]   _zz_2258;
  wire       [31:0]   _zz_2259;
  wire       [15:0]   _zz_2260;
  wire       [31:0]   _zz_2261;
  wire       [31:0]   _zz_2262;
  wire       [31:0]   _zz_2263;
  wire       [31:0]   _zz_2264;
  wire       [31:0]   _zz_2265;
  wire       [23:0]   _zz_2266;
  wire       [31:0]   _zz_2267;
  wire       [15:0]   _zz_2268;
  wire       [31:0]   _zz_2269;
  wire       [31:0]   _zz_2270;
  wire       [31:0]   _zz_2271;
  wire       [31:0]   _zz_2272;
  wire       [31:0]   _zz_2273;
  wire       [23:0]   _zz_2274;
  wire       [31:0]   _zz_2275;
  wire       [15:0]   _zz_2276;
  wire       [15:0]   _zz_2277;
  wire       [31:0]   _zz_2278;
  wire       [31:0]   _zz_2279;
  wire       [15:0]   _zz_2280;
  wire       [31:0]   _zz_2281;
  wire       [31:0]   _zz_2282;
  wire       [31:0]   _zz_2283;
  wire       [15:0]   _zz_2284;
  wire       [31:0]   _zz_2285;
  wire       [31:0]   _zz_2286;
  wire       [31:0]   _zz_2287;
  wire       [31:0]   _zz_2288;
  wire       [31:0]   _zz_2289;
  wire       [31:0]   _zz_2290;
  wire       [23:0]   _zz_2291;
  wire       [31:0]   _zz_2292;
  wire       [15:0]   _zz_2293;
  wire       [31:0]   _zz_2294;
  wire       [31:0]   _zz_2295;
  wire       [31:0]   _zz_2296;
  wire       [31:0]   _zz_2297;
  wire       [31:0]   _zz_2298;
  wire       [23:0]   _zz_2299;
  wire       [31:0]   _zz_2300;
  wire       [15:0]   _zz_2301;
  wire       [31:0]   _zz_2302;
  wire       [31:0]   _zz_2303;
  wire       [31:0]   _zz_2304;
  wire       [31:0]   _zz_2305;
  wire       [31:0]   _zz_2306;
  wire       [23:0]   _zz_2307;
  wire       [31:0]   _zz_2308;
  wire       [15:0]   _zz_2309;
  wire       [31:0]   _zz_2310;
  wire       [31:0]   _zz_2311;
  wire       [31:0]   _zz_2312;
  wire       [31:0]   _zz_2313;
  wire       [31:0]   _zz_2314;
  wire       [23:0]   _zz_2315;
  wire       [31:0]   _zz_2316;
  wire       [15:0]   _zz_2317;
  wire       [15:0]   _zz_2318;
  wire       [31:0]   _zz_2319;
  wire       [31:0]   _zz_2320;
  wire       [15:0]   _zz_2321;
  wire       [31:0]   _zz_2322;
  wire       [31:0]   _zz_2323;
  wire       [31:0]   _zz_2324;
  wire       [15:0]   _zz_2325;
  wire       [31:0]   _zz_2326;
  wire       [31:0]   _zz_2327;
  wire       [31:0]   _zz_2328;
  wire       [31:0]   _zz_2329;
  wire       [31:0]   _zz_2330;
  wire       [31:0]   _zz_2331;
  wire       [23:0]   _zz_2332;
  wire       [31:0]   _zz_2333;
  wire       [15:0]   _zz_2334;
  wire       [31:0]   _zz_2335;
  wire       [31:0]   _zz_2336;
  wire       [31:0]   _zz_2337;
  wire       [31:0]   _zz_2338;
  wire       [31:0]   _zz_2339;
  wire       [23:0]   _zz_2340;
  wire       [31:0]   _zz_2341;
  wire       [15:0]   _zz_2342;
  wire       [31:0]   _zz_2343;
  wire       [31:0]   _zz_2344;
  wire       [31:0]   _zz_2345;
  wire       [31:0]   _zz_2346;
  wire       [31:0]   _zz_2347;
  wire       [23:0]   _zz_2348;
  wire       [31:0]   _zz_2349;
  wire       [15:0]   _zz_2350;
  wire       [31:0]   _zz_2351;
  wire       [31:0]   _zz_2352;
  wire       [31:0]   _zz_2353;
  wire       [31:0]   _zz_2354;
  wire       [31:0]   _zz_2355;
  wire       [23:0]   _zz_2356;
  wire       [31:0]   _zz_2357;
  wire       [15:0]   _zz_2358;
  wire       [15:0]   _zz_2359;
  wire       [31:0]   _zz_2360;
  wire       [31:0]   _zz_2361;
  wire       [15:0]   _zz_2362;
  wire       [31:0]   _zz_2363;
  wire       [31:0]   _zz_2364;
  wire       [31:0]   _zz_2365;
  wire       [15:0]   _zz_2366;
  wire       [31:0]   _zz_2367;
  wire       [31:0]   _zz_2368;
  wire       [31:0]   _zz_2369;
  wire       [31:0]   _zz_2370;
  wire       [31:0]   _zz_2371;
  wire       [31:0]   _zz_2372;
  wire       [23:0]   _zz_2373;
  wire       [31:0]   _zz_2374;
  wire       [15:0]   _zz_2375;
  wire       [31:0]   _zz_2376;
  wire       [31:0]   _zz_2377;
  wire       [31:0]   _zz_2378;
  wire       [31:0]   _zz_2379;
  wire       [31:0]   _zz_2380;
  wire       [23:0]   _zz_2381;
  wire       [31:0]   _zz_2382;
  wire       [15:0]   _zz_2383;
  wire       [31:0]   _zz_2384;
  wire       [31:0]   _zz_2385;
  wire       [31:0]   _zz_2386;
  wire       [31:0]   _zz_2387;
  wire       [31:0]   _zz_2388;
  wire       [23:0]   _zz_2389;
  wire       [31:0]   _zz_2390;
  wire       [15:0]   _zz_2391;
  wire       [31:0]   _zz_2392;
  wire       [31:0]   _zz_2393;
  wire       [31:0]   _zz_2394;
  wire       [31:0]   _zz_2395;
  wire       [31:0]   _zz_2396;
  wire       [23:0]   _zz_2397;
  wire       [31:0]   _zz_2398;
  wire       [15:0]   _zz_2399;
  wire       [15:0]   _zz_2400;
  wire       [31:0]   _zz_2401;
  wire       [31:0]   _zz_2402;
  wire       [15:0]   _zz_2403;
  wire       [31:0]   _zz_2404;
  wire       [31:0]   _zz_2405;
  wire       [31:0]   _zz_2406;
  wire       [15:0]   _zz_2407;
  wire       [31:0]   _zz_2408;
  wire       [31:0]   _zz_2409;
  wire       [31:0]   _zz_2410;
  wire       [31:0]   _zz_2411;
  wire       [31:0]   _zz_2412;
  wire       [31:0]   _zz_2413;
  wire       [23:0]   _zz_2414;
  wire       [31:0]   _zz_2415;
  wire       [15:0]   _zz_2416;
  wire       [31:0]   _zz_2417;
  wire       [31:0]   _zz_2418;
  wire       [31:0]   _zz_2419;
  wire       [31:0]   _zz_2420;
  wire       [31:0]   _zz_2421;
  wire       [23:0]   _zz_2422;
  wire       [31:0]   _zz_2423;
  wire       [15:0]   _zz_2424;
  wire       [31:0]   _zz_2425;
  wire       [31:0]   _zz_2426;
  wire       [31:0]   _zz_2427;
  wire       [31:0]   _zz_2428;
  wire       [31:0]   _zz_2429;
  wire       [23:0]   _zz_2430;
  wire       [31:0]   _zz_2431;
  wire       [15:0]   _zz_2432;
  wire       [31:0]   _zz_2433;
  wire       [31:0]   _zz_2434;
  wire       [31:0]   _zz_2435;
  wire       [31:0]   _zz_2436;
  wire       [31:0]   _zz_2437;
  wire       [23:0]   _zz_2438;
  wire       [31:0]   _zz_2439;
  wire       [15:0]   _zz_2440;
  wire       [15:0]   _zz_2441;
  wire       [31:0]   _zz_2442;
  wire       [31:0]   _zz_2443;
  wire       [15:0]   _zz_2444;
  wire       [31:0]   _zz_2445;
  wire       [31:0]   _zz_2446;
  wire       [31:0]   _zz_2447;
  wire       [15:0]   _zz_2448;
  wire       [31:0]   _zz_2449;
  wire       [31:0]   _zz_2450;
  wire       [31:0]   _zz_2451;
  wire       [31:0]   _zz_2452;
  wire       [31:0]   _zz_2453;
  wire       [31:0]   _zz_2454;
  wire       [23:0]   _zz_2455;
  wire       [31:0]   _zz_2456;
  wire       [15:0]   _zz_2457;
  wire       [31:0]   _zz_2458;
  wire       [31:0]   _zz_2459;
  wire       [31:0]   _zz_2460;
  wire       [31:0]   _zz_2461;
  wire       [31:0]   _zz_2462;
  wire       [23:0]   _zz_2463;
  wire       [31:0]   _zz_2464;
  wire       [15:0]   _zz_2465;
  wire       [31:0]   _zz_2466;
  wire       [31:0]   _zz_2467;
  wire       [31:0]   _zz_2468;
  wire       [31:0]   _zz_2469;
  wire       [31:0]   _zz_2470;
  wire       [23:0]   _zz_2471;
  wire       [31:0]   _zz_2472;
  wire       [15:0]   _zz_2473;
  wire       [31:0]   _zz_2474;
  wire       [31:0]   _zz_2475;
  wire       [31:0]   _zz_2476;
  wire       [31:0]   _zz_2477;
  wire       [31:0]   _zz_2478;
  wire       [23:0]   _zz_2479;
  wire       [31:0]   _zz_2480;
  wire       [15:0]   _zz_2481;
  wire       [15:0]   _zz_2482;
  wire       [31:0]   _zz_2483;
  wire       [31:0]   _zz_2484;
  wire       [15:0]   _zz_2485;
  wire       [31:0]   _zz_2486;
  wire       [31:0]   _zz_2487;
  wire       [31:0]   _zz_2488;
  wire       [15:0]   _zz_2489;
  wire       [31:0]   _zz_2490;
  wire       [31:0]   _zz_2491;
  wire       [31:0]   _zz_2492;
  wire       [31:0]   _zz_2493;
  wire       [31:0]   _zz_2494;
  wire       [31:0]   _zz_2495;
  wire       [23:0]   _zz_2496;
  wire       [31:0]   _zz_2497;
  wire       [15:0]   _zz_2498;
  wire       [31:0]   _zz_2499;
  wire       [31:0]   _zz_2500;
  wire       [31:0]   _zz_2501;
  wire       [31:0]   _zz_2502;
  wire       [31:0]   _zz_2503;
  wire       [23:0]   _zz_2504;
  wire       [31:0]   _zz_2505;
  wire       [15:0]   _zz_2506;
  wire       [31:0]   _zz_2507;
  wire       [31:0]   _zz_2508;
  wire       [31:0]   _zz_2509;
  wire       [31:0]   _zz_2510;
  wire       [31:0]   _zz_2511;
  wire       [23:0]   _zz_2512;
  wire       [31:0]   _zz_2513;
  wire       [15:0]   _zz_2514;
  wire       [31:0]   _zz_2515;
  wire       [31:0]   _zz_2516;
  wire       [31:0]   _zz_2517;
  wire       [31:0]   _zz_2518;
  wire       [31:0]   _zz_2519;
  wire       [23:0]   _zz_2520;
  wire       [31:0]   _zz_2521;
  wire       [15:0]   _zz_2522;
  wire       [15:0]   _zz_2523;
  wire       [31:0]   _zz_2524;
  wire       [31:0]   _zz_2525;
  wire       [15:0]   _zz_2526;
  wire       [31:0]   _zz_2527;
  wire       [31:0]   _zz_2528;
  wire       [31:0]   _zz_2529;
  wire       [15:0]   _zz_2530;
  wire       [31:0]   _zz_2531;
  wire       [31:0]   _zz_2532;
  wire       [31:0]   _zz_2533;
  wire       [31:0]   _zz_2534;
  wire       [31:0]   _zz_2535;
  wire       [31:0]   _zz_2536;
  wire       [23:0]   _zz_2537;
  wire       [31:0]   _zz_2538;
  wire       [15:0]   _zz_2539;
  wire       [31:0]   _zz_2540;
  wire       [31:0]   _zz_2541;
  wire       [31:0]   _zz_2542;
  wire       [31:0]   _zz_2543;
  wire       [31:0]   _zz_2544;
  wire       [23:0]   _zz_2545;
  wire       [31:0]   _zz_2546;
  wire       [15:0]   _zz_2547;
  wire       [31:0]   _zz_2548;
  wire       [31:0]   _zz_2549;
  wire       [31:0]   _zz_2550;
  wire       [31:0]   _zz_2551;
  wire       [31:0]   _zz_2552;
  wire       [23:0]   _zz_2553;
  wire       [31:0]   _zz_2554;
  wire       [15:0]   _zz_2555;
  wire       [31:0]   _zz_2556;
  wire       [31:0]   _zz_2557;
  wire       [31:0]   _zz_2558;
  wire       [31:0]   _zz_2559;
  wire       [31:0]   _zz_2560;
  wire       [23:0]   _zz_2561;
  wire       [31:0]   _zz_2562;
  wire       [15:0]   _zz_2563;
  wire       [15:0]   _zz_2564;
  wire       [31:0]   _zz_2565;
  wire       [31:0]   _zz_2566;
  wire       [15:0]   _zz_2567;
  wire       [31:0]   _zz_2568;
  wire       [31:0]   _zz_2569;
  wire       [31:0]   _zz_2570;
  wire       [15:0]   _zz_2571;
  wire       [31:0]   _zz_2572;
  wire       [31:0]   _zz_2573;
  wire       [31:0]   _zz_2574;
  wire       [31:0]   _zz_2575;
  wire       [31:0]   _zz_2576;
  wire       [31:0]   _zz_2577;
  wire       [23:0]   _zz_2578;
  wire       [31:0]   _zz_2579;
  wire       [15:0]   _zz_2580;
  wire       [31:0]   _zz_2581;
  wire       [31:0]   _zz_2582;
  wire       [31:0]   _zz_2583;
  wire       [31:0]   _zz_2584;
  wire       [31:0]   _zz_2585;
  wire       [23:0]   _zz_2586;
  wire       [31:0]   _zz_2587;
  wire       [15:0]   _zz_2588;
  wire       [31:0]   _zz_2589;
  wire       [31:0]   _zz_2590;
  wire       [31:0]   _zz_2591;
  wire       [31:0]   _zz_2592;
  wire       [31:0]   _zz_2593;
  wire       [23:0]   _zz_2594;
  wire       [31:0]   _zz_2595;
  wire       [15:0]   _zz_2596;
  wire       [31:0]   _zz_2597;
  wire       [31:0]   _zz_2598;
  wire       [31:0]   _zz_2599;
  wire       [31:0]   _zz_2600;
  wire       [31:0]   _zz_2601;
  wire       [23:0]   _zz_2602;
  wire       [31:0]   _zz_2603;
  wire       [15:0]   _zz_2604;
  wire       [15:0]   _zz_2605;
  wire       [31:0]   _zz_2606;
  wire       [31:0]   _zz_2607;
  wire       [15:0]   _zz_2608;
  wire       [31:0]   _zz_2609;
  wire       [31:0]   _zz_2610;
  wire       [31:0]   _zz_2611;
  wire       [15:0]   _zz_2612;
  wire       [31:0]   _zz_2613;
  wire       [31:0]   _zz_2614;
  wire       [31:0]   _zz_2615;
  wire       [31:0]   _zz_2616;
  wire       [31:0]   _zz_2617;
  wire       [31:0]   _zz_2618;
  wire       [23:0]   _zz_2619;
  wire       [31:0]   _zz_2620;
  wire       [15:0]   _zz_2621;
  wire       [31:0]   _zz_2622;
  wire       [31:0]   _zz_2623;
  wire       [31:0]   _zz_2624;
  wire       [31:0]   _zz_2625;
  wire       [31:0]   _zz_2626;
  wire       [23:0]   _zz_2627;
  wire       [31:0]   _zz_2628;
  wire       [15:0]   _zz_2629;
  wire       [31:0]   _zz_2630;
  wire       [31:0]   _zz_2631;
  wire       [31:0]   _zz_2632;
  wire       [31:0]   _zz_2633;
  wire       [31:0]   _zz_2634;
  wire       [23:0]   _zz_2635;
  wire       [31:0]   _zz_2636;
  wire       [15:0]   _zz_2637;
  wire       [31:0]   _zz_2638;
  wire       [31:0]   _zz_2639;
  wire       [31:0]   _zz_2640;
  wire       [31:0]   _zz_2641;
  wire       [31:0]   _zz_2642;
  wire       [23:0]   _zz_2643;
  wire       [31:0]   _zz_2644;
  wire       [15:0]   _zz_2645;
  wire       [15:0]   _zz_2646;
  wire       [31:0]   _zz_2647;
  wire       [31:0]   _zz_2648;
  wire       [15:0]   _zz_2649;
  wire       [31:0]   _zz_2650;
  wire       [31:0]   _zz_2651;
  wire       [31:0]   _zz_2652;
  wire       [15:0]   _zz_2653;
  wire       [31:0]   _zz_2654;
  wire       [31:0]   _zz_2655;
  wire       [31:0]   _zz_2656;
  wire       [31:0]   _zz_2657;
  wire       [31:0]   _zz_2658;
  wire       [31:0]   _zz_2659;
  wire       [23:0]   _zz_2660;
  wire       [31:0]   _zz_2661;
  wire       [15:0]   _zz_2662;
  wire       [31:0]   _zz_2663;
  wire       [31:0]   _zz_2664;
  wire       [31:0]   _zz_2665;
  wire       [31:0]   _zz_2666;
  wire       [31:0]   _zz_2667;
  wire       [23:0]   _zz_2668;
  wire       [31:0]   _zz_2669;
  wire       [15:0]   _zz_2670;
  wire       [31:0]   _zz_2671;
  wire       [31:0]   _zz_2672;
  wire       [31:0]   _zz_2673;
  wire       [31:0]   _zz_2674;
  wire       [31:0]   _zz_2675;
  wire       [23:0]   _zz_2676;
  wire       [31:0]   _zz_2677;
  wire       [15:0]   _zz_2678;
  wire       [31:0]   _zz_2679;
  wire       [31:0]   _zz_2680;
  wire       [31:0]   _zz_2681;
  wire       [31:0]   _zz_2682;
  wire       [31:0]   _zz_2683;
  wire       [23:0]   _zz_2684;
  wire       [31:0]   _zz_2685;
  wire       [15:0]   _zz_2686;
  wire       [15:0]   _zz_2687;
  wire       [31:0]   _zz_2688;
  wire       [31:0]   _zz_2689;
  wire       [15:0]   _zz_2690;
  wire       [31:0]   _zz_2691;
  wire       [31:0]   _zz_2692;
  wire       [31:0]   _zz_2693;
  wire       [15:0]   _zz_2694;
  wire       [31:0]   _zz_2695;
  wire       [31:0]   _zz_2696;
  wire       [31:0]   _zz_2697;
  wire       [31:0]   _zz_2698;
  wire       [31:0]   _zz_2699;
  wire       [31:0]   _zz_2700;
  wire       [23:0]   _zz_2701;
  wire       [31:0]   _zz_2702;
  wire       [15:0]   _zz_2703;
  wire       [31:0]   _zz_2704;
  wire       [31:0]   _zz_2705;
  wire       [31:0]   _zz_2706;
  wire       [31:0]   _zz_2707;
  wire       [31:0]   _zz_2708;
  wire       [23:0]   _zz_2709;
  wire       [31:0]   _zz_2710;
  wire       [15:0]   _zz_2711;
  wire       [31:0]   _zz_2712;
  wire       [31:0]   _zz_2713;
  wire       [31:0]   _zz_2714;
  wire       [31:0]   _zz_2715;
  wire       [31:0]   _zz_2716;
  wire       [23:0]   _zz_2717;
  wire       [31:0]   _zz_2718;
  wire       [15:0]   _zz_2719;
  wire       [31:0]   _zz_2720;
  wire       [31:0]   _zz_2721;
  wire       [31:0]   _zz_2722;
  wire       [31:0]   _zz_2723;
  wire       [31:0]   _zz_2724;
  wire       [23:0]   _zz_2725;
  wire       [31:0]   _zz_2726;
  wire       [15:0]   _zz_2727;
  wire       [15:0]   _zz_2728;
  wire       [31:0]   _zz_2729;
  wire       [31:0]   _zz_2730;
  wire       [15:0]   _zz_2731;
  wire       [31:0]   _zz_2732;
  wire       [31:0]   _zz_2733;
  wire       [31:0]   _zz_2734;
  wire       [15:0]   _zz_2735;
  wire       [31:0]   _zz_2736;
  wire       [31:0]   _zz_2737;
  wire       [31:0]   _zz_2738;
  wire       [31:0]   _zz_2739;
  wire       [31:0]   _zz_2740;
  wire       [31:0]   _zz_2741;
  wire       [23:0]   _zz_2742;
  wire       [31:0]   _zz_2743;
  wire       [15:0]   _zz_2744;
  wire       [31:0]   _zz_2745;
  wire       [31:0]   _zz_2746;
  wire       [31:0]   _zz_2747;
  wire       [31:0]   _zz_2748;
  wire       [31:0]   _zz_2749;
  wire       [23:0]   _zz_2750;
  wire       [31:0]   _zz_2751;
  wire       [15:0]   _zz_2752;
  wire       [31:0]   _zz_2753;
  wire       [31:0]   _zz_2754;
  wire       [31:0]   _zz_2755;
  wire       [31:0]   _zz_2756;
  wire       [31:0]   _zz_2757;
  wire       [23:0]   _zz_2758;
  wire       [31:0]   _zz_2759;
  wire       [15:0]   _zz_2760;
  wire       [31:0]   _zz_2761;
  wire       [31:0]   _zz_2762;
  wire       [31:0]   _zz_2763;
  wire       [31:0]   _zz_2764;
  wire       [31:0]   _zz_2765;
  wire       [23:0]   _zz_2766;
  wire       [31:0]   _zz_2767;
  wire       [15:0]   _zz_2768;
  wire       [15:0]   _zz_2769;
  wire       [31:0]   _zz_2770;
  wire       [31:0]   _zz_2771;
  wire       [15:0]   _zz_2772;
  wire       [31:0]   _zz_2773;
  wire       [31:0]   _zz_2774;
  wire       [31:0]   _zz_2775;
  wire       [15:0]   _zz_2776;
  wire       [31:0]   _zz_2777;
  wire       [31:0]   _zz_2778;
  wire       [31:0]   _zz_2779;
  wire       [31:0]   _zz_2780;
  wire       [31:0]   _zz_2781;
  wire       [31:0]   _zz_2782;
  wire       [23:0]   _zz_2783;
  wire       [31:0]   _zz_2784;
  wire       [15:0]   _zz_2785;
  wire       [31:0]   _zz_2786;
  wire       [31:0]   _zz_2787;
  wire       [31:0]   _zz_2788;
  wire       [31:0]   _zz_2789;
  wire       [31:0]   _zz_2790;
  wire       [23:0]   _zz_2791;
  wire       [31:0]   _zz_2792;
  wire       [15:0]   _zz_2793;
  wire       [31:0]   _zz_2794;
  wire       [31:0]   _zz_2795;
  wire       [31:0]   _zz_2796;
  wire       [31:0]   _zz_2797;
  wire       [31:0]   _zz_2798;
  wire       [23:0]   _zz_2799;
  wire       [31:0]   _zz_2800;
  wire       [15:0]   _zz_2801;
  wire       [31:0]   _zz_2802;
  wire       [31:0]   _zz_2803;
  wire       [31:0]   _zz_2804;
  wire       [31:0]   _zz_2805;
  wire       [31:0]   _zz_2806;
  wire       [23:0]   _zz_2807;
  wire       [31:0]   _zz_2808;
  wire       [15:0]   _zz_2809;
  wire       [15:0]   _zz_2810;
  wire       [31:0]   _zz_2811;
  wire       [31:0]   _zz_2812;
  wire       [15:0]   _zz_2813;
  wire       [31:0]   _zz_2814;
  wire       [31:0]   _zz_2815;
  wire       [31:0]   _zz_2816;
  wire       [15:0]   _zz_2817;
  wire       [31:0]   _zz_2818;
  wire       [31:0]   _zz_2819;
  wire       [31:0]   _zz_2820;
  wire       [31:0]   _zz_2821;
  wire       [31:0]   _zz_2822;
  wire       [31:0]   _zz_2823;
  wire       [23:0]   _zz_2824;
  wire       [31:0]   _zz_2825;
  wire       [15:0]   _zz_2826;
  wire       [31:0]   _zz_2827;
  wire       [31:0]   _zz_2828;
  wire       [31:0]   _zz_2829;
  wire       [31:0]   _zz_2830;
  wire       [31:0]   _zz_2831;
  wire       [23:0]   _zz_2832;
  wire       [31:0]   _zz_2833;
  wire       [15:0]   _zz_2834;
  wire       [31:0]   _zz_2835;
  wire       [31:0]   _zz_2836;
  wire       [31:0]   _zz_2837;
  wire       [31:0]   _zz_2838;
  wire       [31:0]   _zz_2839;
  wire       [23:0]   _zz_2840;
  wire       [31:0]   _zz_2841;
  wire       [15:0]   _zz_2842;
  wire       [31:0]   _zz_2843;
  wire       [31:0]   _zz_2844;
  wire       [31:0]   _zz_2845;
  wire       [31:0]   _zz_2846;
  wire       [31:0]   _zz_2847;
  wire       [23:0]   _zz_2848;
  wire       [31:0]   _zz_2849;
  wire       [15:0]   _zz_2850;
  wire       [15:0]   _zz_2851;
  wire       [31:0]   _zz_2852;
  wire       [31:0]   _zz_2853;
  wire       [15:0]   _zz_2854;
  wire       [31:0]   _zz_2855;
  wire       [31:0]   _zz_2856;
  wire       [31:0]   _zz_2857;
  wire       [15:0]   _zz_2858;
  wire       [31:0]   _zz_2859;
  wire       [31:0]   _zz_2860;
  wire       [31:0]   _zz_2861;
  wire       [31:0]   _zz_2862;
  wire       [31:0]   _zz_2863;
  wire       [31:0]   _zz_2864;
  wire       [23:0]   _zz_2865;
  wire       [31:0]   _zz_2866;
  wire       [15:0]   _zz_2867;
  wire       [31:0]   _zz_2868;
  wire       [31:0]   _zz_2869;
  wire       [31:0]   _zz_2870;
  wire       [31:0]   _zz_2871;
  wire       [31:0]   _zz_2872;
  wire       [23:0]   _zz_2873;
  wire       [31:0]   _zz_2874;
  wire       [15:0]   _zz_2875;
  wire       [31:0]   _zz_2876;
  wire       [31:0]   _zz_2877;
  wire       [31:0]   _zz_2878;
  wire       [31:0]   _zz_2879;
  wire       [31:0]   _zz_2880;
  wire       [23:0]   _zz_2881;
  wire       [31:0]   _zz_2882;
  wire       [15:0]   _zz_2883;
  wire       [31:0]   _zz_2884;
  wire       [31:0]   _zz_2885;
  wire       [31:0]   _zz_2886;
  wire       [31:0]   _zz_2887;
  wire       [31:0]   _zz_2888;
  wire       [23:0]   _zz_2889;
  wire       [31:0]   _zz_2890;
  wire       [15:0]   _zz_2891;
  wire       [15:0]   _zz_2892;
  wire       [31:0]   _zz_2893;
  wire       [31:0]   _zz_2894;
  wire       [15:0]   _zz_2895;
  wire       [31:0]   _zz_2896;
  wire       [31:0]   _zz_2897;
  wire       [31:0]   _zz_2898;
  wire       [15:0]   _zz_2899;
  wire       [31:0]   _zz_2900;
  wire       [31:0]   _zz_2901;
  wire       [31:0]   _zz_2902;
  wire       [31:0]   _zz_2903;
  wire       [31:0]   _zz_2904;
  wire       [31:0]   _zz_2905;
  wire       [23:0]   _zz_2906;
  wire       [31:0]   _zz_2907;
  wire       [15:0]   _zz_2908;
  wire       [31:0]   _zz_2909;
  wire       [31:0]   _zz_2910;
  wire       [31:0]   _zz_2911;
  wire       [31:0]   _zz_2912;
  wire       [31:0]   _zz_2913;
  wire       [23:0]   _zz_2914;
  wire       [31:0]   _zz_2915;
  wire       [15:0]   _zz_2916;
  wire       [31:0]   _zz_2917;
  wire       [31:0]   _zz_2918;
  wire       [31:0]   _zz_2919;
  wire       [31:0]   _zz_2920;
  wire       [31:0]   _zz_2921;
  wire       [23:0]   _zz_2922;
  wire       [31:0]   _zz_2923;
  wire       [15:0]   _zz_2924;
  wire       [31:0]   _zz_2925;
  wire       [31:0]   _zz_2926;
  wire       [31:0]   _zz_2927;
  wire       [31:0]   _zz_2928;
  wire       [31:0]   _zz_2929;
  wire       [23:0]   _zz_2930;
  wire       [31:0]   _zz_2931;
  wire       [15:0]   _zz_2932;
  wire       [15:0]   _zz_2933;
  wire       [31:0]   _zz_2934;
  wire       [31:0]   _zz_2935;
  wire       [15:0]   _zz_2936;
  wire       [31:0]   _zz_2937;
  wire       [31:0]   _zz_2938;
  wire       [31:0]   _zz_2939;
  wire       [15:0]   _zz_2940;
  wire       [31:0]   _zz_2941;
  wire       [31:0]   _zz_2942;
  wire       [31:0]   _zz_2943;
  wire       [31:0]   _zz_2944;
  wire       [31:0]   _zz_2945;
  wire       [31:0]   _zz_2946;
  wire       [23:0]   _zz_2947;
  wire       [31:0]   _zz_2948;
  wire       [15:0]   _zz_2949;
  wire       [31:0]   _zz_2950;
  wire       [31:0]   _zz_2951;
  wire       [31:0]   _zz_2952;
  wire       [31:0]   _zz_2953;
  wire       [31:0]   _zz_2954;
  wire       [23:0]   _zz_2955;
  wire       [31:0]   _zz_2956;
  wire       [15:0]   _zz_2957;
  wire       [31:0]   _zz_2958;
  wire       [31:0]   _zz_2959;
  wire       [31:0]   _zz_2960;
  wire       [31:0]   _zz_2961;
  wire       [31:0]   _zz_2962;
  wire       [23:0]   _zz_2963;
  wire       [31:0]   _zz_2964;
  wire       [15:0]   _zz_2965;
  wire       [31:0]   _zz_2966;
  wire       [31:0]   _zz_2967;
  wire       [31:0]   _zz_2968;
  wire       [31:0]   _zz_2969;
  wire       [31:0]   _zz_2970;
  wire       [23:0]   _zz_2971;
  wire       [31:0]   _zz_2972;
  wire       [15:0]   _zz_2973;
  wire       [15:0]   _zz_2974;
  wire       [31:0]   _zz_2975;
  wire       [31:0]   _zz_2976;
  wire       [15:0]   _zz_2977;
  wire       [31:0]   _zz_2978;
  wire       [31:0]   _zz_2979;
  wire       [31:0]   _zz_2980;
  wire       [15:0]   _zz_2981;
  wire       [31:0]   _zz_2982;
  wire       [31:0]   _zz_2983;
  wire       [31:0]   _zz_2984;
  wire       [31:0]   _zz_2985;
  wire       [31:0]   _zz_2986;
  wire       [31:0]   _zz_2987;
  wire       [23:0]   _zz_2988;
  wire       [31:0]   _zz_2989;
  wire       [15:0]   _zz_2990;
  wire       [31:0]   _zz_2991;
  wire       [31:0]   _zz_2992;
  wire       [31:0]   _zz_2993;
  wire       [31:0]   _zz_2994;
  wire       [31:0]   _zz_2995;
  wire       [23:0]   _zz_2996;
  wire       [31:0]   _zz_2997;
  wire       [15:0]   _zz_2998;
  wire       [31:0]   _zz_2999;
  wire       [31:0]   _zz_3000;
  wire       [31:0]   _zz_3001;
  wire       [31:0]   _zz_3002;
  wire       [31:0]   _zz_3003;
  wire       [23:0]   _zz_3004;
  wire       [31:0]   _zz_3005;
  wire       [15:0]   _zz_3006;
  wire       [31:0]   _zz_3007;
  wire       [31:0]   _zz_3008;
  wire       [31:0]   _zz_3009;
  wire       [31:0]   _zz_3010;
  wire       [31:0]   _zz_3011;
  wire       [23:0]   _zz_3012;
  wire       [31:0]   _zz_3013;
  wire       [15:0]   _zz_3014;
  wire       [15:0]   _zz_3015;
  wire       [31:0]   _zz_3016;
  wire       [31:0]   _zz_3017;
  wire       [15:0]   _zz_3018;
  wire       [31:0]   _zz_3019;
  wire       [31:0]   _zz_3020;
  wire       [31:0]   _zz_3021;
  wire       [15:0]   _zz_3022;
  wire       [31:0]   _zz_3023;
  wire       [31:0]   _zz_3024;
  wire       [31:0]   _zz_3025;
  wire       [31:0]   _zz_3026;
  wire       [31:0]   _zz_3027;
  wire       [31:0]   _zz_3028;
  wire       [23:0]   _zz_3029;
  wire       [31:0]   _zz_3030;
  wire       [15:0]   _zz_3031;
  wire       [31:0]   _zz_3032;
  wire       [31:0]   _zz_3033;
  wire       [31:0]   _zz_3034;
  wire       [31:0]   _zz_3035;
  wire       [31:0]   _zz_3036;
  wire       [23:0]   _zz_3037;
  wire       [31:0]   _zz_3038;
  wire       [15:0]   _zz_3039;
  wire       [31:0]   _zz_3040;
  wire       [31:0]   _zz_3041;
  wire       [31:0]   _zz_3042;
  wire       [31:0]   _zz_3043;
  wire       [31:0]   _zz_3044;
  wire       [23:0]   _zz_3045;
  wire       [31:0]   _zz_3046;
  wire       [15:0]   _zz_3047;
  wire       [31:0]   _zz_3048;
  wire       [31:0]   _zz_3049;
  wire       [31:0]   _zz_3050;
  wire       [31:0]   _zz_3051;
  wire       [31:0]   _zz_3052;
  wire       [23:0]   _zz_3053;
  wire       [31:0]   _zz_3054;
  wire       [15:0]   _zz_3055;
  wire       [15:0]   _zz_3056;
  wire       [31:0]   _zz_3057;
  wire       [31:0]   _zz_3058;
  wire       [15:0]   _zz_3059;
  wire       [31:0]   _zz_3060;
  wire       [31:0]   _zz_3061;
  wire       [31:0]   _zz_3062;
  wire       [15:0]   _zz_3063;
  wire       [31:0]   _zz_3064;
  wire       [31:0]   _zz_3065;
  wire       [31:0]   _zz_3066;
  wire       [31:0]   _zz_3067;
  wire       [31:0]   _zz_3068;
  wire       [31:0]   _zz_3069;
  wire       [23:0]   _zz_3070;
  wire       [31:0]   _zz_3071;
  wire       [15:0]   _zz_3072;
  wire       [31:0]   _zz_3073;
  wire       [31:0]   _zz_3074;
  wire       [31:0]   _zz_3075;
  wire       [31:0]   _zz_3076;
  wire       [31:0]   _zz_3077;
  wire       [23:0]   _zz_3078;
  wire       [31:0]   _zz_3079;
  wire       [15:0]   _zz_3080;
  wire       [31:0]   _zz_3081;
  wire       [31:0]   _zz_3082;
  wire       [31:0]   _zz_3083;
  wire       [31:0]   _zz_3084;
  wire       [31:0]   _zz_3085;
  wire       [23:0]   _zz_3086;
  wire       [31:0]   _zz_3087;
  wire       [15:0]   _zz_3088;
  wire       [31:0]   _zz_3089;
  wire       [31:0]   _zz_3090;
  wire       [31:0]   _zz_3091;
  wire       [31:0]   _zz_3092;
  wire       [31:0]   _zz_3093;
  wire       [23:0]   _zz_3094;
  wire       [31:0]   _zz_3095;
  wire       [15:0]   _zz_3096;
  wire       [15:0]   _zz_3097;
  wire       [31:0]   _zz_3098;
  wire       [31:0]   _zz_3099;
  wire       [15:0]   _zz_3100;
  wire       [31:0]   _zz_3101;
  wire       [31:0]   _zz_3102;
  wire       [31:0]   _zz_3103;
  wire       [15:0]   _zz_3104;
  wire       [31:0]   _zz_3105;
  wire       [31:0]   _zz_3106;
  wire       [31:0]   _zz_3107;
  wire       [31:0]   _zz_3108;
  wire       [31:0]   _zz_3109;
  wire       [31:0]   _zz_3110;
  wire       [23:0]   _zz_3111;
  wire       [31:0]   _zz_3112;
  wire       [15:0]   _zz_3113;
  wire       [31:0]   _zz_3114;
  wire       [31:0]   _zz_3115;
  wire       [31:0]   _zz_3116;
  wire       [31:0]   _zz_3117;
  wire       [31:0]   _zz_3118;
  wire       [23:0]   _zz_3119;
  wire       [31:0]   _zz_3120;
  wire       [15:0]   _zz_3121;
  wire       [31:0]   _zz_3122;
  wire       [31:0]   _zz_3123;
  wire       [31:0]   _zz_3124;
  wire       [31:0]   _zz_3125;
  wire       [31:0]   _zz_3126;
  wire       [23:0]   _zz_3127;
  wire       [31:0]   _zz_3128;
  wire       [15:0]   _zz_3129;
  wire       [31:0]   _zz_3130;
  wire       [31:0]   _zz_3131;
  wire       [31:0]   _zz_3132;
  wire       [31:0]   _zz_3133;
  wire       [31:0]   _zz_3134;
  wire       [23:0]   _zz_3135;
  wire       [31:0]   _zz_3136;
  wire       [15:0]   _zz_3137;
  wire       [15:0]   _zz_3138;
  wire       [31:0]   _zz_3139;
  wire       [31:0]   _zz_3140;
  wire       [15:0]   _zz_3141;
  wire       [31:0]   _zz_3142;
  wire       [31:0]   _zz_3143;
  wire       [31:0]   _zz_3144;
  wire       [15:0]   _zz_3145;
  wire       [31:0]   _zz_3146;
  wire       [31:0]   _zz_3147;
  wire       [31:0]   _zz_3148;
  wire       [31:0]   _zz_3149;
  wire       [31:0]   _zz_3150;
  wire       [31:0]   _zz_3151;
  wire       [23:0]   _zz_3152;
  wire       [31:0]   _zz_3153;
  wire       [15:0]   _zz_3154;
  wire       [31:0]   _zz_3155;
  wire       [31:0]   _zz_3156;
  wire       [31:0]   _zz_3157;
  wire       [31:0]   _zz_3158;
  wire       [31:0]   _zz_3159;
  wire       [23:0]   _zz_3160;
  wire       [31:0]   _zz_3161;
  wire       [15:0]   _zz_3162;
  wire       [31:0]   _zz_3163;
  wire       [31:0]   _zz_3164;
  wire       [31:0]   _zz_3165;
  wire       [31:0]   _zz_3166;
  wire       [31:0]   _zz_3167;
  wire       [23:0]   _zz_3168;
  wire       [31:0]   _zz_3169;
  wire       [15:0]   _zz_3170;
  wire       [31:0]   _zz_3171;
  wire       [31:0]   _zz_3172;
  wire       [31:0]   _zz_3173;
  wire       [31:0]   _zz_3174;
  wire       [31:0]   _zz_3175;
  wire       [23:0]   _zz_3176;
  wire       [31:0]   _zz_3177;
  wire       [15:0]   _zz_3178;
  wire       [15:0]   _zz_3179;
  wire       [31:0]   _zz_3180;
  wire       [31:0]   _zz_3181;
  wire       [15:0]   _zz_3182;
  wire       [31:0]   _zz_3183;
  wire       [31:0]   _zz_3184;
  wire       [31:0]   _zz_3185;
  wire       [15:0]   _zz_3186;
  wire       [31:0]   _zz_3187;
  wire       [31:0]   _zz_3188;
  wire       [31:0]   _zz_3189;
  wire       [31:0]   _zz_3190;
  wire       [31:0]   _zz_3191;
  wire       [31:0]   _zz_3192;
  wire       [23:0]   _zz_3193;
  wire       [31:0]   _zz_3194;
  wire       [15:0]   _zz_3195;
  wire       [31:0]   _zz_3196;
  wire       [31:0]   _zz_3197;
  wire       [31:0]   _zz_3198;
  wire       [31:0]   _zz_3199;
  wire       [31:0]   _zz_3200;
  wire       [23:0]   _zz_3201;
  wire       [31:0]   _zz_3202;
  wire       [15:0]   _zz_3203;
  wire       [31:0]   _zz_3204;
  wire       [31:0]   _zz_3205;
  wire       [31:0]   _zz_3206;
  wire       [31:0]   _zz_3207;
  wire       [31:0]   _zz_3208;
  wire       [23:0]   _zz_3209;
  wire       [31:0]   _zz_3210;
  wire       [15:0]   _zz_3211;
  wire       [31:0]   _zz_3212;
  wire       [31:0]   _zz_3213;
  wire       [31:0]   _zz_3214;
  wire       [31:0]   _zz_3215;
  wire       [31:0]   _zz_3216;
  wire       [23:0]   _zz_3217;
  wire       [31:0]   _zz_3218;
  wire       [15:0]   _zz_3219;
  wire       [15:0]   _zz_3220;
  wire       [31:0]   _zz_3221;
  wire       [31:0]   _zz_3222;
  wire       [15:0]   _zz_3223;
  wire       [31:0]   _zz_3224;
  wire       [31:0]   _zz_3225;
  wire       [31:0]   _zz_3226;
  wire       [15:0]   _zz_3227;
  wire       [31:0]   _zz_3228;
  wire       [31:0]   _zz_3229;
  wire       [31:0]   _zz_3230;
  wire       [31:0]   _zz_3231;
  wire       [31:0]   _zz_3232;
  wire       [31:0]   _zz_3233;
  wire       [23:0]   _zz_3234;
  wire       [31:0]   _zz_3235;
  wire       [15:0]   _zz_3236;
  wire       [31:0]   _zz_3237;
  wire       [31:0]   _zz_3238;
  wire       [31:0]   _zz_3239;
  wire       [31:0]   _zz_3240;
  wire       [31:0]   _zz_3241;
  wire       [23:0]   _zz_3242;
  wire       [31:0]   _zz_3243;
  wire       [15:0]   _zz_3244;
  wire       [31:0]   _zz_3245;
  wire       [31:0]   _zz_3246;
  wire       [31:0]   _zz_3247;
  wire       [31:0]   _zz_3248;
  wire       [31:0]   _zz_3249;
  wire       [23:0]   _zz_3250;
  wire       [31:0]   _zz_3251;
  wire       [15:0]   _zz_3252;
  wire       [31:0]   _zz_3253;
  wire       [31:0]   _zz_3254;
  wire       [31:0]   _zz_3255;
  wire       [31:0]   _zz_3256;
  wire       [31:0]   _zz_3257;
  wire       [23:0]   _zz_3258;
  wire       [31:0]   _zz_3259;
  wire       [15:0]   _zz_3260;
  wire       [15:0]   _zz_3261;
  wire       [31:0]   _zz_3262;
  wire       [31:0]   _zz_3263;
  wire       [15:0]   _zz_3264;
  wire       [31:0]   _zz_3265;
  wire       [31:0]   _zz_3266;
  wire       [31:0]   _zz_3267;
  wire       [15:0]   _zz_3268;
  wire       [31:0]   _zz_3269;
  wire       [31:0]   _zz_3270;
  wire       [31:0]   _zz_3271;
  wire       [31:0]   _zz_3272;
  wire       [31:0]   _zz_3273;
  wire       [31:0]   _zz_3274;
  wire       [23:0]   _zz_3275;
  wire       [31:0]   _zz_3276;
  wire       [15:0]   _zz_3277;
  wire       [31:0]   _zz_3278;
  wire       [31:0]   _zz_3279;
  wire       [31:0]   _zz_3280;
  wire       [31:0]   _zz_3281;
  wire       [31:0]   _zz_3282;
  wire       [23:0]   _zz_3283;
  wire       [31:0]   _zz_3284;
  wire       [15:0]   _zz_3285;
  wire       [31:0]   _zz_3286;
  wire       [31:0]   _zz_3287;
  wire       [31:0]   _zz_3288;
  wire       [31:0]   _zz_3289;
  wire       [31:0]   _zz_3290;
  wire       [23:0]   _zz_3291;
  wire       [31:0]   _zz_3292;
  wire       [15:0]   _zz_3293;
  wire       [31:0]   _zz_3294;
  wire       [31:0]   _zz_3295;
  wire       [31:0]   _zz_3296;
  wire       [31:0]   _zz_3297;
  wire       [31:0]   _zz_3298;
  wire       [23:0]   _zz_3299;
  wire       [31:0]   _zz_3300;
  wire       [15:0]   _zz_3301;
  wire       [15:0]   _zz_3302;
  wire       [31:0]   _zz_3303;
  wire       [31:0]   _zz_3304;
  wire       [15:0]   _zz_3305;
  wire       [31:0]   _zz_3306;
  wire       [31:0]   _zz_3307;
  wire       [31:0]   _zz_3308;
  wire       [15:0]   _zz_3309;
  wire       [31:0]   _zz_3310;
  wire       [31:0]   _zz_3311;
  wire       [31:0]   _zz_3312;
  wire       [31:0]   _zz_3313;
  wire       [31:0]   _zz_3314;
  wire       [31:0]   _zz_3315;
  wire       [23:0]   _zz_3316;
  wire       [31:0]   _zz_3317;
  wire       [15:0]   _zz_3318;
  wire       [31:0]   _zz_3319;
  wire       [31:0]   _zz_3320;
  wire       [31:0]   _zz_3321;
  wire       [31:0]   _zz_3322;
  wire       [31:0]   _zz_3323;
  wire       [23:0]   _zz_3324;
  wire       [31:0]   _zz_3325;
  wire       [15:0]   _zz_3326;
  wire       [31:0]   _zz_3327;
  wire       [31:0]   _zz_3328;
  wire       [31:0]   _zz_3329;
  wire       [31:0]   _zz_3330;
  wire       [31:0]   _zz_3331;
  wire       [23:0]   _zz_3332;
  wire       [31:0]   _zz_3333;
  wire       [15:0]   _zz_3334;
  wire       [31:0]   _zz_3335;
  wire       [31:0]   _zz_3336;
  wire       [31:0]   _zz_3337;
  wire       [31:0]   _zz_3338;
  wire       [31:0]   _zz_3339;
  wire       [23:0]   _zz_3340;
  wire       [31:0]   _zz_3341;
  wire       [15:0]   _zz_3342;
  wire       [15:0]   _zz_3343;
  wire       [31:0]   _zz_3344;
  wire       [31:0]   _zz_3345;
  wire       [15:0]   _zz_3346;
  wire       [31:0]   _zz_3347;
  wire       [31:0]   _zz_3348;
  wire       [31:0]   _zz_3349;
  wire       [15:0]   _zz_3350;
  wire       [31:0]   _zz_3351;
  wire       [31:0]   _zz_3352;
  wire       [31:0]   _zz_3353;
  wire       [31:0]   _zz_3354;
  wire       [31:0]   _zz_3355;
  wire       [31:0]   _zz_3356;
  wire       [23:0]   _zz_3357;
  wire       [31:0]   _zz_3358;
  wire       [15:0]   _zz_3359;
  wire       [31:0]   _zz_3360;
  wire       [31:0]   _zz_3361;
  wire       [31:0]   _zz_3362;
  wire       [31:0]   _zz_3363;
  wire       [31:0]   _zz_3364;
  wire       [23:0]   _zz_3365;
  wire       [31:0]   _zz_3366;
  wire       [15:0]   _zz_3367;
  wire       [31:0]   _zz_3368;
  wire       [31:0]   _zz_3369;
  wire       [31:0]   _zz_3370;
  wire       [31:0]   _zz_3371;
  wire       [31:0]   _zz_3372;
  wire       [23:0]   _zz_3373;
  wire       [31:0]   _zz_3374;
  wire       [15:0]   _zz_3375;
  wire       [31:0]   _zz_3376;
  wire       [31:0]   _zz_3377;
  wire       [31:0]   _zz_3378;
  wire       [31:0]   _zz_3379;
  wire       [31:0]   _zz_3380;
  wire       [23:0]   _zz_3381;
  wire       [31:0]   _zz_3382;
  wire       [15:0]   _zz_3383;
  wire       [15:0]   _zz_3384;
  wire       [31:0]   _zz_3385;
  wire       [31:0]   _zz_3386;
  wire       [15:0]   _zz_3387;
  wire       [31:0]   _zz_3388;
  wire       [31:0]   _zz_3389;
  wire       [31:0]   _zz_3390;
  wire       [15:0]   _zz_3391;
  wire       [31:0]   _zz_3392;
  wire       [31:0]   _zz_3393;
  wire       [31:0]   _zz_3394;
  wire       [31:0]   _zz_3395;
  wire       [31:0]   _zz_3396;
  wire       [31:0]   _zz_3397;
  wire       [23:0]   _zz_3398;
  wire       [31:0]   _zz_3399;
  wire       [15:0]   _zz_3400;
  wire       [31:0]   _zz_3401;
  wire       [31:0]   _zz_3402;
  wire       [31:0]   _zz_3403;
  wire       [31:0]   _zz_3404;
  wire       [31:0]   _zz_3405;
  wire       [23:0]   _zz_3406;
  wire       [31:0]   _zz_3407;
  wire       [15:0]   _zz_3408;
  wire       [31:0]   _zz_3409;
  wire       [31:0]   _zz_3410;
  wire       [31:0]   _zz_3411;
  wire       [31:0]   _zz_3412;
  wire       [31:0]   _zz_3413;
  wire       [23:0]   _zz_3414;
  wire       [31:0]   _zz_3415;
  wire       [15:0]   _zz_3416;
  wire       [31:0]   _zz_3417;
  wire       [31:0]   _zz_3418;
  wire       [31:0]   _zz_3419;
  wire       [31:0]   _zz_3420;
  wire       [31:0]   _zz_3421;
  wire       [23:0]   _zz_3422;
  wire       [31:0]   _zz_3423;
  wire       [15:0]   _zz_3424;
  wire       [15:0]   _zz_3425;
  wire       [31:0]   _zz_3426;
  wire       [31:0]   _zz_3427;
  wire       [15:0]   _zz_3428;
  wire       [31:0]   _zz_3429;
  wire       [31:0]   _zz_3430;
  wire       [31:0]   _zz_3431;
  wire       [15:0]   _zz_3432;
  wire       [31:0]   _zz_3433;
  wire       [31:0]   _zz_3434;
  wire       [31:0]   _zz_3435;
  wire       [31:0]   _zz_3436;
  wire       [31:0]   _zz_3437;
  wire       [31:0]   _zz_3438;
  wire       [23:0]   _zz_3439;
  wire       [31:0]   _zz_3440;
  wire       [15:0]   _zz_3441;
  wire       [31:0]   _zz_3442;
  wire       [31:0]   _zz_3443;
  wire       [31:0]   _zz_3444;
  wire       [31:0]   _zz_3445;
  wire       [31:0]   _zz_3446;
  wire       [23:0]   _zz_3447;
  wire       [31:0]   _zz_3448;
  wire       [15:0]   _zz_3449;
  wire       [31:0]   _zz_3450;
  wire       [31:0]   _zz_3451;
  wire       [31:0]   _zz_3452;
  wire       [31:0]   _zz_3453;
  wire       [31:0]   _zz_3454;
  wire       [23:0]   _zz_3455;
  wire       [31:0]   _zz_3456;
  wire       [15:0]   _zz_3457;
  wire       [31:0]   _zz_3458;
  wire       [31:0]   _zz_3459;
  wire       [31:0]   _zz_3460;
  wire       [31:0]   _zz_3461;
  wire       [31:0]   _zz_3462;
  wire       [23:0]   _zz_3463;
  wire       [31:0]   _zz_3464;
  wire       [15:0]   _zz_3465;
  wire       [15:0]   _zz_3466;
  wire       [31:0]   _zz_3467;
  wire       [31:0]   _zz_3468;
  wire       [15:0]   _zz_3469;
  wire       [31:0]   _zz_3470;
  wire       [31:0]   _zz_3471;
  wire       [31:0]   _zz_3472;
  wire       [15:0]   _zz_3473;
  wire       [31:0]   _zz_3474;
  wire       [31:0]   _zz_3475;
  wire       [31:0]   _zz_3476;
  wire       [31:0]   _zz_3477;
  wire       [31:0]   _zz_3478;
  wire       [31:0]   _zz_3479;
  wire       [23:0]   _zz_3480;
  wire       [31:0]   _zz_3481;
  wire       [15:0]   _zz_3482;
  wire       [31:0]   _zz_3483;
  wire       [31:0]   _zz_3484;
  wire       [31:0]   _zz_3485;
  wire       [31:0]   _zz_3486;
  wire       [31:0]   _zz_3487;
  wire       [23:0]   _zz_3488;
  wire       [31:0]   _zz_3489;
  wire       [15:0]   _zz_3490;
  wire       [31:0]   _zz_3491;
  wire       [31:0]   _zz_3492;
  wire       [31:0]   _zz_3493;
  wire       [31:0]   _zz_3494;
  wire       [31:0]   _zz_3495;
  wire       [23:0]   _zz_3496;
  wire       [31:0]   _zz_3497;
  wire       [15:0]   _zz_3498;
  wire       [31:0]   _zz_3499;
  wire       [31:0]   _zz_3500;
  wire       [31:0]   _zz_3501;
  wire       [31:0]   _zz_3502;
  wire       [31:0]   _zz_3503;
  wire       [23:0]   _zz_3504;
  wire       [31:0]   _zz_3505;
  wire       [15:0]   _zz_3506;
  wire       [15:0]   _zz_3507;
  wire       [31:0]   _zz_3508;
  wire       [31:0]   _zz_3509;
  wire       [15:0]   _zz_3510;
  wire       [31:0]   _zz_3511;
  wire       [31:0]   _zz_3512;
  wire       [31:0]   _zz_3513;
  wire       [15:0]   _zz_3514;
  wire       [31:0]   _zz_3515;
  wire       [31:0]   _zz_3516;
  wire       [31:0]   _zz_3517;
  wire       [31:0]   _zz_3518;
  wire       [31:0]   _zz_3519;
  wire       [31:0]   _zz_3520;
  wire       [23:0]   _zz_3521;
  wire       [31:0]   _zz_3522;
  wire       [15:0]   _zz_3523;
  wire       [31:0]   _zz_3524;
  wire       [31:0]   _zz_3525;
  wire       [31:0]   _zz_3526;
  wire       [31:0]   _zz_3527;
  wire       [31:0]   _zz_3528;
  wire       [23:0]   _zz_3529;
  wire       [31:0]   _zz_3530;
  wire       [15:0]   _zz_3531;
  wire       [31:0]   _zz_3532;
  wire       [31:0]   _zz_3533;
  wire       [31:0]   _zz_3534;
  wire       [31:0]   _zz_3535;
  wire       [31:0]   _zz_3536;
  wire       [23:0]   _zz_3537;
  wire       [31:0]   _zz_3538;
  wire       [15:0]   _zz_3539;
  wire       [31:0]   _zz_3540;
  wire       [31:0]   _zz_3541;
  wire       [31:0]   _zz_3542;
  wire       [31:0]   _zz_3543;
  wire       [31:0]   _zz_3544;
  wire       [23:0]   _zz_3545;
  wire       [31:0]   _zz_3546;
  wire       [15:0]   _zz_3547;
  wire       [15:0]   _zz_3548;
  wire       [31:0]   _zz_3549;
  wire       [31:0]   _zz_3550;
  wire       [15:0]   _zz_3551;
  wire       [31:0]   _zz_3552;
  wire       [31:0]   _zz_3553;
  wire       [31:0]   _zz_3554;
  wire       [15:0]   _zz_3555;
  wire       [31:0]   _zz_3556;
  wire       [31:0]   _zz_3557;
  wire       [31:0]   _zz_3558;
  wire       [31:0]   _zz_3559;
  wire       [31:0]   _zz_3560;
  wire       [31:0]   _zz_3561;
  wire       [23:0]   _zz_3562;
  wire       [31:0]   _zz_3563;
  wire       [15:0]   _zz_3564;
  wire       [31:0]   _zz_3565;
  wire       [31:0]   _zz_3566;
  wire       [31:0]   _zz_3567;
  wire       [31:0]   _zz_3568;
  wire       [31:0]   _zz_3569;
  wire       [23:0]   _zz_3570;
  wire       [31:0]   _zz_3571;
  wire       [15:0]   _zz_3572;
  wire       [31:0]   _zz_3573;
  wire       [31:0]   _zz_3574;
  wire       [31:0]   _zz_3575;
  wire       [31:0]   _zz_3576;
  wire       [31:0]   _zz_3577;
  wire       [23:0]   _zz_3578;
  wire       [31:0]   _zz_3579;
  wire       [15:0]   _zz_3580;
  wire       [31:0]   _zz_3581;
  wire       [31:0]   _zz_3582;
  wire       [31:0]   _zz_3583;
  wire       [31:0]   _zz_3584;
  wire       [31:0]   _zz_3585;
  wire       [23:0]   _zz_3586;
  wire       [31:0]   _zz_3587;
  wire       [15:0]   _zz_3588;
  wire       [15:0]   _zz_3589;
  wire       [31:0]   _zz_3590;
  wire       [31:0]   _zz_3591;
  wire       [15:0]   _zz_3592;
  wire       [31:0]   _zz_3593;
  wire       [31:0]   _zz_3594;
  wire       [31:0]   _zz_3595;
  wire       [15:0]   _zz_3596;
  wire       [31:0]   _zz_3597;
  wire       [31:0]   _zz_3598;
  wire       [31:0]   _zz_3599;
  wire       [31:0]   _zz_3600;
  wire       [31:0]   _zz_3601;
  wire       [31:0]   _zz_3602;
  wire       [23:0]   _zz_3603;
  wire       [31:0]   _zz_3604;
  wire       [15:0]   _zz_3605;
  wire       [31:0]   _zz_3606;
  wire       [31:0]   _zz_3607;
  wire       [31:0]   _zz_3608;
  wire       [31:0]   _zz_3609;
  wire       [31:0]   _zz_3610;
  wire       [23:0]   _zz_3611;
  wire       [31:0]   _zz_3612;
  wire       [15:0]   _zz_3613;
  wire       [31:0]   _zz_3614;
  wire       [31:0]   _zz_3615;
  wire       [31:0]   _zz_3616;
  wire       [31:0]   _zz_3617;
  wire       [31:0]   _zz_3618;
  wire       [23:0]   _zz_3619;
  wire       [31:0]   _zz_3620;
  wire       [15:0]   _zz_3621;
  wire       [31:0]   _zz_3622;
  wire       [31:0]   _zz_3623;
  wire       [31:0]   _zz_3624;
  wire       [31:0]   _zz_3625;
  wire       [31:0]   _zz_3626;
  wire       [23:0]   _zz_3627;
  wire       [31:0]   _zz_3628;
  wire       [15:0]   _zz_3629;
  wire       [15:0]   _zz_3630;
  wire       [31:0]   _zz_3631;
  wire       [31:0]   _zz_3632;
  wire       [15:0]   _zz_3633;
  wire       [31:0]   _zz_3634;
  wire       [31:0]   _zz_3635;
  wire       [31:0]   _zz_3636;
  wire       [15:0]   _zz_3637;
  wire       [31:0]   _zz_3638;
  wire       [31:0]   _zz_3639;
  wire       [31:0]   _zz_3640;
  wire       [31:0]   _zz_3641;
  wire       [31:0]   _zz_3642;
  wire       [31:0]   _zz_3643;
  wire       [23:0]   _zz_3644;
  wire       [31:0]   _zz_3645;
  wire       [15:0]   _zz_3646;
  wire       [31:0]   _zz_3647;
  wire       [31:0]   _zz_3648;
  wire       [31:0]   _zz_3649;
  wire       [31:0]   _zz_3650;
  wire       [31:0]   _zz_3651;
  wire       [23:0]   _zz_3652;
  wire       [31:0]   _zz_3653;
  wire       [15:0]   _zz_3654;
  wire       [31:0]   _zz_3655;
  wire       [31:0]   _zz_3656;
  wire       [31:0]   _zz_3657;
  wire       [31:0]   _zz_3658;
  wire       [31:0]   _zz_3659;
  wire       [23:0]   _zz_3660;
  wire       [31:0]   _zz_3661;
  wire       [15:0]   _zz_3662;
  wire       [31:0]   _zz_3663;
  wire       [31:0]   _zz_3664;
  wire       [31:0]   _zz_3665;
  wire       [31:0]   _zz_3666;
  wire       [31:0]   _zz_3667;
  wire       [23:0]   _zz_3668;
  wire       [31:0]   _zz_3669;
  wire       [15:0]   _zz_3670;
  wire       [15:0]   _zz_3671;
  wire       [31:0]   _zz_3672;
  wire       [31:0]   _zz_3673;
  wire       [15:0]   _zz_3674;
  wire       [31:0]   _zz_3675;
  wire       [31:0]   _zz_3676;
  wire       [31:0]   _zz_3677;
  wire       [15:0]   _zz_3678;
  wire       [31:0]   _zz_3679;
  wire       [31:0]   _zz_3680;
  wire       [31:0]   _zz_3681;
  wire       [31:0]   _zz_3682;
  wire       [31:0]   _zz_3683;
  wire       [31:0]   _zz_3684;
  wire       [23:0]   _zz_3685;
  wire       [31:0]   _zz_3686;
  wire       [15:0]   _zz_3687;
  wire       [31:0]   _zz_3688;
  wire       [31:0]   _zz_3689;
  wire       [31:0]   _zz_3690;
  wire       [31:0]   _zz_3691;
  wire       [31:0]   _zz_3692;
  wire       [23:0]   _zz_3693;
  wire       [31:0]   _zz_3694;
  wire       [15:0]   _zz_3695;
  wire       [31:0]   _zz_3696;
  wire       [31:0]   _zz_3697;
  wire       [31:0]   _zz_3698;
  wire       [31:0]   _zz_3699;
  wire       [31:0]   _zz_3700;
  wire       [23:0]   _zz_3701;
  wire       [31:0]   _zz_3702;
  wire       [15:0]   _zz_3703;
  wire       [31:0]   _zz_3704;
  wire       [31:0]   _zz_3705;
  wire       [31:0]   _zz_3706;
  wire       [31:0]   _zz_3707;
  wire       [31:0]   _zz_3708;
  wire       [23:0]   _zz_3709;
  wire       [31:0]   _zz_3710;
  wire       [15:0]   _zz_3711;
  wire       [15:0]   _zz_3712;
  wire       [31:0]   _zz_3713;
  wire       [31:0]   _zz_3714;
  wire       [15:0]   _zz_3715;
  wire       [31:0]   _zz_3716;
  wire       [31:0]   _zz_3717;
  wire       [31:0]   _zz_3718;
  wire       [15:0]   _zz_3719;
  wire       [31:0]   _zz_3720;
  wire       [31:0]   _zz_3721;
  wire       [31:0]   _zz_3722;
  wire       [31:0]   _zz_3723;
  wire       [31:0]   _zz_3724;
  wire       [31:0]   _zz_3725;
  wire       [23:0]   _zz_3726;
  wire       [31:0]   _zz_3727;
  wire       [15:0]   _zz_3728;
  wire       [31:0]   _zz_3729;
  wire       [31:0]   _zz_3730;
  wire       [31:0]   _zz_3731;
  wire       [31:0]   _zz_3732;
  wire       [31:0]   _zz_3733;
  wire       [23:0]   _zz_3734;
  wire       [31:0]   _zz_3735;
  wire       [15:0]   _zz_3736;
  wire       [31:0]   _zz_3737;
  wire       [31:0]   _zz_3738;
  wire       [31:0]   _zz_3739;
  wire       [31:0]   _zz_3740;
  wire       [31:0]   _zz_3741;
  wire       [23:0]   _zz_3742;
  wire       [31:0]   _zz_3743;
  wire       [15:0]   _zz_3744;
  wire       [31:0]   _zz_3745;
  wire       [31:0]   _zz_3746;
  wire       [31:0]   _zz_3747;
  wire       [31:0]   _zz_3748;
  wire       [31:0]   _zz_3749;
  wire       [23:0]   _zz_3750;
  wire       [31:0]   _zz_3751;
  wire       [15:0]   _zz_3752;
  wire       [15:0]   _zz_3753;
  wire       [31:0]   _zz_3754;
  wire       [31:0]   _zz_3755;
  wire       [15:0]   _zz_3756;
  wire       [31:0]   _zz_3757;
  wire       [31:0]   _zz_3758;
  wire       [31:0]   _zz_3759;
  wire       [15:0]   _zz_3760;
  wire       [31:0]   _zz_3761;
  wire       [31:0]   _zz_3762;
  wire       [31:0]   _zz_3763;
  wire       [31:0]   _zz_3764;
  wire       [31:0]   _zz_3765;
  wire       [31:0]   _zz_3766;
  wire       [23:0]   _zz_3767;
  wire       [31:0]   _zz_3768;
  wire       [15:0]   _zz_3769;
  wire       [31:0]   _zz_3770;
  wire       [31:0]   _zz_3771;
  wire       [31:0]   _zz_3772;
  wire       [31:0]   _zz_3773;
  wire       [31:0]   _zz_3774;
  wire       [23:0]   _zz_3775;
  wire       [31:0]   _zz_3776;
  wire       [15:0]   _zz_3777;
  wire       [31:0]   _zz_3778;
  wire       [31:0]   _zz_3779;
  wire       [31:0]   _zz_3780;
  wire       [31:0]   _zz_3781;
  wire       [31:0]   _zz_3782;
  wire       [23:0]   _zz_3783;
  wire       [31:0]   _zz_3784;
  wire       [15:0]   _zz_3785;
  wire       [31:0]   _zz_3786;
  wire       [31:0]   _zz_3787;
  wire       [31:0]   _zz_3788;
  wire       [31:0]   _zz_3789;
  wire       [31:0]   _zz_3790;
  wire       [23:0]   _zz_3791;
  wire       [31:0]   _zz_3792;
  wire       [15:0]   _zz_3793;
  wire       [15:0]   _zz_3794;
  wire       [31:0]   _zz_3795;
  wire       [31:0]   _zz_3796;
  wire       [15:0]   _zz_3797;
  wire       [31:0]   _zz_3798;
  wire       [31:0]   _zz_3799;
  wire       [31:0]   _zz_3800;
  wire       [15:0]   _zz_3801;
  wire       [31:0]   _zz_3802;
  wire       [31:0]   _zz_3803;
  wire       [31:0]   _zz_3804;
  wire       [31:0]   _zz_3805;
  wire       [31:0]   _zz_3806;
  wire       [31:0]   _zz_3807;
  wire       [23:0]   _zz_3808;
  wire       [31:0]   _zz_3809;
  wire       [15:0]   _zz_3810;
  wire       [31:0]   _zz_3811;
  wire       [31:0]   _zz_3812;
  wire       [31:0]   _zz_3813;
  wire       [31:0]   _zz_3814;
  wire       [31:0]   _zz_3815;
  wire       [23:0]   _zz_3816;
  wire       [31:0]   _zz_3817;
  wire       [15:0]   _zz_3818;
  wire       [31:0]   _zz_3819;
  wire       [31:0]   _zz_3820;
  wire       [31:0]   _zz_3821;
  wire       [31:0]   _zz_3822;
  wire       [31:0]   _zz_3823;
  wire       [23:0]   _zz_3824;
  wire       [31:0]   _zz_3825;
  wire       [15:0]   _zz_3826;
  wire       [31:0]   _zz_3827;
  wire       [31:0]   _zz_3828;
  wire       [31:0]   _zz_3829;
  wire       [31:0]   _zz_3830;
  wire       [31:0]   _zz_3831;
  wire       [23:0]   _zz_3832;
  wire       [31:0]   _zz_3833;
  wire       [15:0]   _zz_3834;
  wire       [15:0]   _zz_3835;
  wire       [31:0]   _zz_3836;
  wire       [31:0]   _zz_3837;
  wire       [15:0]   _zz_3838;
  wire       [31:0]   _zz_3839;
  wire       [31:0]   _zz_3840;
  wire       [31:0]   _zz_3841;
  wire       [15:0]   _zz_3842;
  wire       [31:0]   _zz_3843;
  wire       [31:0]   _zz_3844;
  wire       [31:0]   _zz_3845;
  wire       [31:0]   _zz_3846;
  wire       [31:0]   _zz_3847;
  wire       [31:0]   _zz_3848;
  wire       [23:0]   _zz_3849;
  wire       [31:0]   _zz_3850;
  wire       [15:0]   _zz_3851;
  wire       [31:0]   _zz_3852;
  wire       [31:0]   _zz_3853;
  wire       [31:0]   _zz_3854;
  wire       [31:0]   _zz_3855;
  wire       [31:0]   _zz_3856;
  wire       [23:0]   _zz_3857;
  wire       [31:0]   _zz_3858;
  wire       [15:0]   _zz_3859;
  wire       [31:0]   _zz_3860;
  wire       [31:0]   _zz_3861;
  wire       [31:0]   _zz_3862;
  wire       [31:0]   _zz_3863;
  wire       [31:0]   _zz_3864;
  wire       [23:0]   _zz_3865;
  wire       [31:0]   _zz_3866;
  wire       [15:0]   _zz_3867;
  wire       [31:0]   _zz_3868;
  wire       [31:0]   _zz_3869;
  wire       [31:0]   _zz_3870;
  wire       [31:0]   _zz_3871;
  wire       [31:0]   _zz_3872;
  wire       [23:0]   _zz_3873;
  wire       [31:0]   _zz_3874;
  wire       [15:0]   _zz_3875;
  wire       [15:0]   _zz_3876;
  wire       [31:0]   _zz_3877;
  wire       [31:0]   _zz_3878;
  wire       [15:0]   _zz_3879;
  wire       [31:0]   _zz_3880;
  wire       [31:0]   _zz_3881;
  wire       [31:0]   _zz_3882;
  wire       [15:0]   _zz_3883;
  wire       [31:0]   _zz_3884;
  wire       [31:0]   _zz_3885;
  wire       [31:0]   _zz_3886;
  wire       [31:0]   _zz_3887;
  wire       [31:0]   _zz_3888;
  wire       [31:0]   _zz_3889;
  wire       [23:0]   _zz_3890;
  wire       [31:0]   _zz_3891;
  wire       [15:0]   _zz_3892;
  wire       [31:0]   _zz_3893;
  wire       [31:0]   _zz_3894;
  wire       [31:0]   _zz_3895;
  wire       [31:0]   _zz_3896;
  wire       [31:0]   _zz_3897;
  wire       [23:0]   _zz_3898;
  wire       [31:0]   _zz_3899;
  wire       [15:0]   _zz_3900;
  wire       [31:0]   _zz_3901;
  wire       [31:0]   _zz_3902;
  wire       [31:0]   _zz_3903;
  wire       [31:0]   _zz_3904;
  wire       [31:0]   _zz_3905;
  wire       [23:0]   _zz_3906;
  wire       [31:0]   _zz_3907;
  wire       [15:0]   _zz_3908;
  wire       [31:0]   _zz_3909;
  wire       [31:0]   _zz_3910;
  wire       [31:0]   _zz_3911;
  wire       [31:0]   _zz_3912;
  wire       [31:0]   _zz_3913;
  wire       [23:0]   _zz_3914;
  wire       [31:0]   _zz_3915;
  wire       [15:0]   _zz_3916;
  wire       [15:0]   _zz_3917;
  wire       [31:0]   _zz_3918;
  wire       [31:0]   _zz_3919;
  wire       [15:0]   _zz_3920;
  wire       [31:0]   _zz_3921;
  wire       [31:0]   _zz_3922;
  wire       [31:0]   _zz_3923;
  wire       [15:0]   _zz_3924;
  wire       [31:0]   _zz_3925;
  wire       [31:0]   _zz_3926;
  wire       [31:0]   _zz_3927;
  wire       [31:0]   _zz_3928;
  wire       [31:0]   _zz_3929;
  wire       [31:0]   _zz_3930;
  wire       [23:0]   _zz_3931;
  wire       [31:0]   _zz_3932;
  wire       [15:0]   _zz_3933;
  wire       [31:0]   _zz_3934;
  wire       [31:0]   _zz_3935;
  wire       [31:0]   _zz_3936;
  wire       [31:0]   _zz_3937;
  wire       [31:0]   _zz_3938;
  wire       [23:0]   _zz_3939;
  wire       [31:0]   _zz_3940;
  wire       [15:0]   _zz_3941;
  wire       [31:0]   _zz_3942;
  wire       [31:0]   _zz_3943;
  wire       [31:0]   _zz_3944;
  wire       [31:0]   _zz_3945;
  wire       [31:0]   _zz_3946;
  wire       [23:0]   _zz_3947;
  wire       [31:0]   _zz_3948;
  wire       [15:0]   _zz_3949;
  wire       [31:0]   _zz_3950;
  wire       [31:0]   _zz_3951;
  wire       [31:0]   _zz_3952;
  wire       [31:0]   _zz_3953;
  wire       [31:0]   _zz_3954;
  wire       [23:0]   _zz_3955;
  wire       [31:0]   _zz_3956;
  wire       [15:0]   _zz_3957;
  wire       [15:0]   _zz_3958;
  wire       [31:0]   _zz_3959;
  wire       [31:0]   _zz_3960;
  wire       [15:0]   _zz_3961;
  wire       [31:0]   _zz_3962;
  wire       [31:0]   _zz_3963;
  wire       [31:0]   _zz_3964;
  wire       [15:0]   _zz_3965;
  wire       [31:0]   _zz_3966;
  wire       [31:0]   _zz_3967;
  wire       [31:0]   _zz_3968;
  wire       [31:0]   _zz_3969;
  wire       [31:0]   _zz_3970;
  wire       [31:0]   _zz_3971;
  wire       [23:0]   _zz_3972;
  wire       [31:0]   _zz_3973;
  wire       [15:0]   _zz_3974;
  wire       [31:0]   _zz_3975;
  wire       [31:0]   _zz_3976;
  wire       [31:0]   _zz_3977;
  wire       [31:0]   _zz_3978;
  wire       [31:0]   _zz_3979;
  wire       [23:0]   _zz_3980;
  wire       [31:0]   _zz_3981;
  wire       [15:0]   _zz_3982;
  wire       [31:0]   _zz_3983;
  wire       [31:0]   _zz_3984;
  wire       [31:0]   _zz_3985;
  wire       [31:0]   _zz_3986;
  wire       [31:0]   _zz_3987;
  wire       [23:0]   _zz_3988;
  wire       [31:0]   _zz_3989;
  wire       [15:0]   _zz_3990;
  wire       [31:0]   _zz_3991;
  wire       [31:0]   _zz_3992;
  wire       [31:0]   _zz_3993;
  wire       [31:0]   _zz_3994;
  wire       [31:0]   _zz_3995;
  wire       [23:0]   _zz_3996;
  wire       [31:0]   _zz_3997;
  wire       [15:0]   _zz_3998;
  wire       [15:0]   _zz_3999;
  wire       [31:0]   _zz_4000;
  wire       [31:0]   _zz_4001;
  wire       [15:0]   _zz_4002;
  wire       [31:0]   _zz_4003;
  wire       [31:0]   _zz_4004;
  wire       [31:0]   _zz_4005;
  wire       [15:0]   _zz_4006;
  wire       [31:0]   _zz_4007;
  wire       [31:0]   _zz_4008;
  wire       [31:0]   _zz_4009;
  wire       [31:0]   _zz_4010;
  wire       [31:0]   _zz_4011;
  wire       [31:0]   _zz_4012;
  wire       [23:0]   _zz_4013;
  wire       [31:0]   _zz_4014;
  wire       [15:0]   _zz_4015;
  wire       [31:0]   _zz_4016;
  wire       [31:0]   _zz_4017;
  wire       [31:0]   _zz_4018;
  wire       [31:0]   _zz_4019;
  wire       [31:0]   _zz_4020;
  wire       [23:0]   _zz_4021;
  wire       [31:0]   _zz_4022;
  wire       [15:0]   _zz_4023;
  wire       [31:0]   _zz_4024;
  wire       [31:0]   _zz_4025;
  wire       [31:0]   _zz_4026;
  wire       [31:0]   _zz_4027;
  wire       [31:0]   _zz_4028;
  wire       [23:0]   _zz_4029;
  wire       [31:0]   _zz_4030;
  wire       [15:0]   _zz_4031;
  wire       [31:0]   _zz_4032;
  wire       [31:0]   _zz_4033;
  wire       [31:0]   _zz_4034;
  wire       [31:0]   _zz_4035;
  wire       [31:0]   _zz_4036;
  wire       [23:0]   _zz_4037;
  wire       [31:0]   _zz_4038;
  wire       [15:0]   _zz_4039;
  wire       [15:0]   _zz_4040;
  wire       [31:0]   _zz_4041;
  wire       [31:0]   _zz_4042;
  wire       [15:0]   _zz_4043;
  wire       [31:0]   _zz_4044;
  wire       [31:0]   _zz_4045;
  wire       [31:0]   _zz_4046;
  wire       [15:0]   _zz_4047;
  wire       [31:0]   _zz_4048;
  wire       [31:0]   _zz_4049;
  wire       [31:0]   _zz_4050;
  wire       [31:0]   _zz_4051;
  wire       [31:0]   _zz_4052;
  wire       [31:0]   _zz_4053;
  wire       [23:0]   _zz_4054;
  wire       [31:0]   _zz_4055;
  wire       [15:0]   _zz_4056;
  wire       [31:0]   _zz_4057;
  wire       [31:0]   _zz_4058;
  wire       [31:0]   _zz_4059;
  wire       [31:0]   _zz_4060;
  wire       [31:0]   _zz_4061;
  wire       [23:0]   _zz_4062;
  wire       [31:0]   _zz_4063;
  wire       [15:0]   _zz_4064;
  wire       [31:0]   _zz_4065;
  wire       [31:0]   _zz_4066;
  wire       [31:0]   _zz_4067;
  wire       [31:0]   _zz_4068;
  wire       [31:0]   _zz_4069;
  wire       [23:0]   _zz_4070;
  wire       [31:0]   _zz_4071;
  wire       [15:0]   _zz_4072;
  wire       [31:0]   _zz_4073;
  wire       [31:0]   _zz_4074;
  wire       [31:0]   _zz_4075;
  wire       [31:0]   _zz_4076;
  wire       [31:0]   _zz_4077;
  wire       [23:0]   _zz_4078;
  wire       [31:0]   _zz_4079;
  wire       [15:0]   _zz_4080;
  wire       [15:0]   _zz_4081;
  wire       [31:0]   _zz_4082;
  wire       [31:0]   _zz_4083;
  wire       [15:0]   _zz_4084;
  wire       [31:0]   _zz_4085;
  wire       [31:0]   _zz_4086;
  wire       [31:0]   _zz_4087;
  wire       [15:0]   _zz_4088;
  wire       [31:0]   _zz_4089;
  wire       [31:0]   _zz_4090;
  wire       [31:0]   _zz_4091;
  wire       [31:0]   _zz_4092;
  wire       [31:0]   _zz_4093;
  wire       [31:0]   _zz_4094;
  wire       [23:0]   _zz_4095;
  wire       [31:0]   _zz_4096;
  wire       [15:0]   _zz_4097;
  wire       [31:0]   _zz_4098;
  wire       [31:0]   _zz_4099;
  wire       [31:0]   _zz_4100;
  wire       [31:0]   _zz_4101;
  wire       [31:0]   _zz_4102;
  wire       [23:0]   _zz_4103;
  wire       [31:0]   _zz_4104;
  wire       [15:0]   _zz_4105;
  wire       [31:0]   _zz_4106;
  wire       [31:0]   _zz_4107;
  wire       [31:0]   _zz_4108;
  wire       [31:0]   _zz_4109;
  wire       [31:0]   _zz_4110;
  wire       [23:0]   _zz_4111;
  wire       [31:0]   _zz_4112;
  wire       [15:0]   _zz_4113;
  wire       [31:0]   _zz_4114;
  wire       [31:0]   _zz_4115;
  wire       [31:0]   _zz_4116;
  wire       [31:0]   _zz_4117;
  wire       [31:0]   _zz_4118;
  wire       [23:0]   _zz_4119;
  wire       [31:0]   _zz_4120;
  wire       [15:0]   _zz_4121;
  wire       [15:0]   _zz_4122;
  wire       [31:0]   _zz_4123;
  wire       [31:0]   _zz_4124;
  wire       [15:0]   _zz_4125;
  wire       [31:0]   _zz_4126;
  wire       [31:0]   _zz_4127;
  wire       [31:0]   _zz_4128;
  wire       [15:0]   _zz_4129;
  wire       [31:0]   _zz_4130;
  wire       [31:0]   _zz_4131;
  wire       [31:0]   _zz_4132;
  wire       [31:0]   _zz_4133;
  wire       [31:0]   _zz_4134;
  wire       [31:0]   _zz_4135;
  wire       [23:0]   _zz_4136;
  wire       [31:0]   _zz_4137;
  wire       [15:0]   _zz_4138;
  wire       [31:0]   _zz_4139;
  wire       [31:0]   _zz_4140;
  wire       [31:0]   _zz_4141;
  wire       [31:0]   _zz_4142;
  wire       [31:0]   _zz_4143;
  wire       [23:0]   _zz_4144;
  wire       [31:0]   _zz_4145;
  wire       [15:0]   _zz_4146;
  wire       [31:0]   _zz_4147;
  wire       [31:0]   _zz_4148;
  wire       [31:0]   _zz_4149;
  wire       [31:0]   _zz_4150;
  wire       [31:0]   _zz_4151;
  wire       [23:0]   _zz_4152;
  wire       [31:0]   _zz_4153;
  wire       [15:0]   _zz_4154;
  wire       [31:0]   _zz_4155;
  wire       [31:0]   _zz_4156;
  wire       [31:0]   _zz_4157;
  wire       [31:0]   _zz_4158;
  wire       [31:0]   _zz_4159;
  wire       [23:0]   _zz_4160;
  wire       [31:0]   _zz_4161;
  wire       [15:0]   _zz_4162;
  reg        [15:0]   data_in_0_real;
  reg        [15:0]   data_in_0_imag;
  reg        [15:0]   data_in_1_real;
  reg        [15:0]   data_in_1_imag;
  reg        [15:0]   data_in_2_real;
  reg        [15:0]   data_in_2_imag;
  reg        [15:0]   data_in_3_real;
  reg        [15:0]   data_in_3_imag;
  reg        [15:0]   data_in_4_real;
  reg        [15:0]   data_in_4_imag;
  reg        [15:0]   data_in_5_real;
  reg        [15:0]   data_in_5_imag;
  reg        [15:0]   data_in_6_real;
  reg        [15:0]   data_in_6_imag;
  reg        [15:0]   data_in_7_real;
  reg        [15:0]   data_in_7_imag;
  reg        [15:0]   data_in_8_real;
  reg        [15:0]   data_in_8_imag;
  reg        [15:0]   data_in_9_real;
  reg        [15:0]   data_in_9_imag;
  reg        [15:0]   data_in_10_real;
  reg        [15:0]   data_in_10_imag;
  reg        [15:0]   data_in_11_real;
  reg        [15:0]   data_in_11_imag;
  reg        [15:0]   data_in_12_real;
  reg        [15:0]   data_in_12_imag;
  reg        [15:0]   data_in_13_real;
  reg        [15:0]   data_in_13_imag;
  reg        [15:0]   data_in_14_real;
  reg        [15:0]   data_in_14_imag;
  reg        [15:0]   data_in_15_real;
  reg        [15:0]   data_in_15_imag;
  reg        [15:0]   data_in_16_real;
  reg        [15:0]   data_in_16_imag;
  reg        [15:0]   data_in_17_real;
  reg        [15:0]   data_in_17_imag;
  reg        [15:0]   data_in_18_real;
  reg        [15:0]   data_in_18_imag;
  reg        [15:0]   data_in_19_real;
  reg        [15:0]   data_in_19_imag;
  reg        [15:0]   data_in_20_real;
  reg        [15:0]   data_in_20_imag;
  reg        [15:0]   data_in_21_real;
  reg        [15:0]   data_in_21_imag;
  reg        [15:0]   data_in_22_real;
  reg        [15:0]   data_in_22_imag;
  reg        [15:0]   data_in_23_real;
  reg        [15:0]   data_in_23_imag;
  reg        [15:0]   data_in_24_real;
  reg        [15:0]   data_in_24_imag;
  reg        [15:0]   data_in_25_real;
  reg        [15:0]   data_in_25_imag;
  reg        [15:0]   data_in_26_real;
  reg        [15:0]   data_in_26_imag;
  reg        [15:0]   data_in_27_real;
  reg        [15:0]   data_in_27_imag;
  reg        [15:0]   data_in_28_real;
  reg        [15:0]   data_in_28_imag;
  reg        [15:0]   data_in_29_real;
  reg        [15:0]   data_in_29_imag;
  reg        [15:0]   data_in_30_real;
  reg        [15:0]   data_in_30_imag;
  reg        [15:0]   data_in_31_real;
  reg        [15:0]   data_in_31_imag;
  wire       [15:0]   twiddle_factor_table_0_real;
  wire       [15:0]   twiddle_factor_table_0_imag;
  wire       [15:0]   twiddle_factor_table_1_real;
  wire       [15:0]   twiddle_factor_table_1_imag;
  wire       [15:0]   twiddle_factor_table_2_real;
  wire       [15:0]   twiddle_factor_table_2_imag;
  wire       [15:0]   twiddle_factor_table_3_real;
  wire       [15:0]   twiddle_factor_table_3_imag;
  wire       [15:0]   twiddle_factor_table_4_real;
  wire       [15:0]   twiddle_factor_table_4_imag;
  wire       [15:0]   twiddle_factor_table_5_real;
  wire       [15:0]   twiddle_factor_table_5_imag;
  wire       [15:0]   twiddle_factor_table_6_real;
  wire       [15:0]   twiddle_factor_table_6_imag;
  wire       [15:0]   twiddle_factor_table_7_real;
  wire       [15:0]   twiddle_factor_table_7_imag;
  wire       [15:0]   twiddle_factor_table_8_real;
  wire       [15:0]   twiddle_factor_table_8_imag;
  wire       [15:0]   twiddle_factor_table_9_real;
  wire       [15:0]   twiddle_factor_table_9_imag;
  wire       [15:0]   twiddle_factor_table_10_real;
  wire       [15:0]   twiddle_factor_table_10_imag;
  wire       [15:0]   twiddle_factor_table_11_real;
  wire       [15:0]   twiddle_factor_table_11_imag;
  wire       [15:0]   twiddle_factor_table_12_real;
  wire       [15:0]   twiddle_factor_table_12_imag;
  wire       [15:0]   twiddle_factor_table_13_real;
  wire       [15:0]   twiddle_factor_table_13_imag;
  wire       [15:0]   twiddle_factor_table_14_real;
  wire       [15:0]   twiddle_factor_table_14_imag;
  wire       [15:0]   twiddle_factor_table_15_real;
  wire       [15:0]   twiddle_factor_table_15_imag;
  wire       [15:0]   twiddle_factor_table_16_real;
  wire       [15:0]   twiddle_factor_table_16_imag;
  wire       [15:0]   twiddle_factor_table_17_real;
  wire       [15:0]   twiddle_factor_table_17_imag;
  wire       [15:0]   twiddle_factor_table_18_real;
  wire       [15:0]   twiddle_factor_table_18_imag;
  wire       [15:0]   twiddle_factor_table_19_real;
  wire       [15:0]   twiddle_factor_table_19_imag;
  wire       [15:0]   twiddle_factor_table_20_real;
  wire       [15:0]   twiddle_factor_table_20_imag;
  wire       [15:0]   twiddle_factor_table_21_real;
  wire       [15:0]   twiddle_factor_table_21_imag;
  wire       [15:0]   twiddle_factor_table_22_real;
  wire       [15:0]   twiddle_factor_table_22_imag;
  wire       [15:0]   twiddle_factor_table_23_real;
  wire       [15:0]   twiddle_factor_table_23_imag;
  wire       [15:0]   twiddle_factor_table_24_real;
  wire       [15:0]   twiddle_factor_table_24_imag;
  wire       [15:0]   twiddle_factor_table_25_real;
  wire       [15:0]   twiddle_factor_table_25_imag;
  wire       [15:0]   twiddle_factor_table_26_real;
  wire       [15:0]   twiddle_factor_table_26_imag;
  wire       [15:0]   twiddle_factor_table_27_real;
  wire       [15:0]   twiddle_factor_table_27_imag;
  wire       [15:0]   twiddle_factor_table_28_real;
  wire       [15:0]   twiddle_factor_table_28_imag;
  wire       [15:0]   twiddle_factor_table_29_real;
  wire       [15:0]   twiddle_factor_table_29_imag;
  wire       [15:0]   twiddle_factor_table_30_real;
  wire       [15:0]   twiddle_factor_table_30_imag;
  wire       [15:0]   data_reorder_0_real;
  wire       [15:0]   data_reorder_0_imag;
  wire       [15:0]   data_reorder_1_real;
  wire       [15:0]   data_reorder_1_imag;
  wire       [15:0]   data_reorder_2_real;
  wire       [15:0]   data_reorder_2_imag;
  wire       [15:0]   data_reorder_3_real;
  wire       [15:0]   data_reorder_3_imag;
  wire       [15:0]   data_reorder_4_real;
  wire       [15:0]   data_reorder_4_imag;
  wire       [15:0]   data_reorder_5_real;
  wire       [15:0]   data_reorder_5_imag;
  wire       [15:0]   data_reorder_6_real;
  wire       [15:0]   data_reorder_6_imag;
  wire       [15:0]   data_reorder_7_real;
  wire       [15:0]   data_reorder_7_imag;
  wire       [15:0]   data_reorder_8_real;
  wire       [15:0]   data_reorder_8_imag;
  wire       [15:0]   data_reorder_9_real;
  wire       [15:0]   data_reorder_9_imag;
  wire       [15:0]   data_reorder_10_real;
  wire       [15:0]   data_reorder_10_imag;
  wire       [15:0]   data_reorder_11_real;
  wire       [15:0]   data_reorder_11_imag;
  wire       [15:0]   data_reorder_12_real;
  wire       [15:0]   data_reorder_12_imag;
  wire       [15:0]   data_reorder_13_real;
  wire       [15:0]   data_reorder_13_imag;
  wire       [15:0]   data_reorder_14_real;
  wire       [15:0]   data_reorder_14_imag;
  wire       [15:0]   data_reorder_15_real;
  wire       [15:0]   data_reorder_15_imag;
  wire       [15:0]   data_reorder_16_real;
  wire       [15:0]   data_reorder_16_imag;
  wire       [15:0]   data_reorder_17_real;
  wire       [15:0]   data_reorder_17_imag;
  wire       [15:0]   data_reorder_18_real;
  wire       [15:0]   data_reorder_18_imag;
  wire       [15:0]   data_reorder_19_real;
  wire       [15:0]   data_reorder_19_imag;
  wire       [15:0]   data_reorder_20_real;
  wire       [15:0]   data_reorder_20_imag;
  wire       [15:0]   data_reorder_21_real;
  wire       [15:0]   data_reorder_21_imag;
  wire       [15:0]   data_reorder_22_real;
  wire       [15:0]   data_reorder_22_imag;
  wire       [15:0]   data_reorder_23_real;
  wire       [15:0]   data_reorder_23_imag;
  wire       [15:0]   data_reorder_24_real;
  wire       [15:0]   data_reorder_24_imag;
  wire       [15:0]   data_reorder_25_real;
  wire       [15:0]   data_reorder_25_imag;
  wire       [15:0]   data_reorder_26_real;
  wire       [15:0]   data_reorder_26_imag;
  wire       [15:0]   data_reorder_27_real;
  wire       [15:0]   data_reorder_27_imag;
  wire       [15:0]   data_reorder_28_real;
  wire       [15:0]   data_reorder_28_imag;
  wire       [15:0]   data_reorder_29_real;
  wire       [15:0]   data_reorder_29_imag;
  wire       [15:0]   data_reorder_30_real;
  wire       [15:0]   data_reorder_30_imag;
  wire       [15:0]   data_reorder_31_real;
  wire       [15:0]   data_reorder_31_imag;
  reg                 io_data_in_valid_regNext;
  reg                 current_level_willIncrement;
  wire                current_level_willClear;
  reg        [2:0]    current_level_valueNext;
  reg        [2:0]    current_level_value;
  wire                current_level_willOverflowIfInc;
  wire                current_level_willOverflow;
  reg                 null_cond_period_minus_1;
  wire                null_cond_period;
  reg        [15:0]   data_mid_0_real;
  reg        [15:0]   data_mid_0_imag;
  reg        [15:0]   data_mid_1_real;
  reg        [15:0]   data_mid_1_imag;
  reg        [15:0]   data_mid_2_real;
  reg        [15:0]   data_mid_2_imag;
  reg        [15:0]   data_mid_3_real;
  reg        [15:0]   data_mid_3_imag;
  reg        [15:0]   data_mid_4_real;
  reg        [15:0]   data_mid_4_imag;
  reg        [15:0]   data_mid_5_real;
  reg        [15:0]   data_mid_5_imag;
  reg        [15:0]   data_mid_6_real;
  reg        [15:0]   data_mid_6_imag;
  reg        [15:0]   data_mid_7_real;
  reg        [15:0]   data_mid_7_imag;
  reg        [15:0]   data_mid_8_real;
  reg        [15:0]   data_mid_8_imag;
  reg        [15:0]   data_mid_9_real;
  reg        [15:0]   data_mid_9_imag;
  reg        [15:0]   data_mid_10_real;
  reg        [15:0]   data_mid_10_imag;
  reg        [15:0]   data_mid_11_real;
  reg        [15:0]   data_mid_11_imag;
  reg        [15:0]   data_mid_12_real;
  reg        [15:0]   data_mid_12_imag;
  reg        [15:0]   data_mid_13_real;
  reg        [15:0]   data_mid_13_imag;
  reg        [15:0]   data_mid_14_real;
  reg        [15:0]   data_mid_14_imag;
  reg        [15:0]   data_mid_15_real;
  reg        [15:0]   data_mid_15_imag;
  reg        [15:0]   data_mid_16_real;
  reg        [15:0]   data_mid_16_imag;
  reg        [15:0]   data_mid_17_real;
  reg        [15:0]   data_mid_17_imag;
  reg        [15:0]   data_mid_18_real;
  reg        [15:0]   data_mid_18_imag;
  reg        [15:0]   data_mid_19_real;
  reg        [15:0]   data_mid_19_imag;
  reg        [15:0]   data_mid_20_real;
  reg        [15:0]   data_mid_20_imag;
  reg        [15:0]   data_mid_21_real;
  reg        [15:0]   data_mid_21_imag;
  reg        [15:0]   data_mid_22_real;
  reg        [15:0]   data_mid_22_imag;
  reg        [15:0]   data_mid_23_real;
  reg        [15:0]   data_mid_23_imag;
  reg        [15:0]   data_mid_24_real;
  reg        [15:0]   data_mid_24_imag;
  reg        [15:0]   data_mid_25_real;
  reg        [15:0]   data_mid_25_imag;
  reg        [15:0]   data_mid_26_real;
  reg        [15:0]   data_mid_26_imag;
  reg        [15:0]   data_mid_27_real;
  reg        [15:0]   data_mid_27_imag;
  reg        [15:0]   data_mid_28_real;
  reg        [15:0]   data_mid_28_imag;
  reg        [15:0]   data_mid_29_real;
  reg        [15:0]   data_mid_29_imag;
  reg        [15:0]   data_mid_30_real;
  reg        [15:0]   data_mid_30_imag;
  reg        [15:0]   data_mid_31_real;
  reg        [15:0]   data_mid_31_imag;
  wire       [31:0]   _zz_1;
  wire       [31:0]   _zz_2;
  wire       [31:0]   _zz_3;
  wire       [0:0]    _zz_4;
  wire       [0:0]    _zz_5;
  wire       [31:0]   _zz_6;
  wire       [31:0]   _zz_7;
  wire       [31:0]   _zz_8;
  wire       [0:0]    _zz_9;
  wire       [0:0]    _zz_10;
  wire       [31:0]   _zz_11;
  wire       [31:0]   _zz_12;
  wire       [31:0]   _zz_13;
  wire       [0:0]    _zz_14;
  wire       [0:0]    _zz_15;
  wire       [31:0]   _zz_16;
  wire       [31:0]   _zz_17;
  wire       [31:0]   _zz_18;
  wire       [0:0]    _zz_19;
  wire       [0:0]    _zz_20;
  wire       [31:0]   _zz_21;
  wire       [31:0]   _zz_22;
  wire       [31:0]   _zz_23;
  wire       [0:0]    _zz_24;
  wire       [0:0]    _zz_25;
  wire       [31:0]   _zz_26;
  wire       [31:0]   _zz_27;
  wire       [31:0]   _zz_28;
  wire       [0:0]    _zz_29;
  wire       [0:0]    _zz_30;
  wire       [31:0]   _zz_31;
  wire       [31:0]   _zz_32;
  wire       [31:0]   _zz_33;
  wire       [0:0]    _zz_34;
  wire       [0:0]    _zz_35;
  wire       [31:0]   _zz_36;
  wire       [31:0]   _zz_37;
  wire       [31:0]   _zz_38;
  wire       [0:0]    _zz_39;
  wire       [0:0]    _zz_40;
  wire       [31:0]   _zz_41;
  wire       [31:0]   _zz_42;
  wire       [31:0]   _zz_43;
  wire       [0:0]    _zz_44;
  wire       [0:0]    _zz_45;
  wire       [31:0]   _zz_46;
  wire       [31:0]   _zz_47;
  wire       [31:0]   _zz_48;
  wire       [0:0]    _zz_49;
  wire       [0:0]    _zz_50;
  wire       [31:0]   _zz_51;
  wire       [31:0]   _zz_52;
  wire       [31:0]   _zz_53;
  wire       [0:0]    _zz_54;
  wire       [0:0]    _zz_55;
  wire       [31:0]   _zz_56;
  wire       [31:0]   _zz_57;
  wire       [31:0]   _zz_58;
  wire       [0:0]    _zz_59;
  wire       [0:0]    _zz_60;
  wire       [31:0]   _zz_61;
  wire       [31:0]   _zz_62;
  wire       [31:0]   _zz_63;
  wire       [0:0]    _zz_64;
  wire       [0:0]    _zz_65;
  wire       [31:0]   _zz_66;
  wire       [31:0]   _zz_67;
  wire       [31:0]   _zz_68;
  wire       [0:0]    _zz_69;
  wire       [0:0]    _zz_70;
  wire       [31:0]   _zz_71;
  wire       [31:0]   _zz_72;
  wire       [31:0]   _zz_73;
  wire       [0:0]    _zz_74;
  wire       [0:0]    _zz_75;
  wire       [31:0]   _zz_76;
  wire       [31:0]   _zz_77;
  wire       [31:0]   _zz_78;
  wire       [0:0]    _zz_79;
  wire       [0:0]    _zz_80;
  wire       [31:0]   _zz_81;
  wire       [31:0]   _zz_82;
  wire       [31:0]   _zz_83;
  wire       [0:0]    _zz_84;
  wire       [0:0]    _zz_85;
  wire       [31:0]   _zz_86;
  wire       [31:0]   _zz_87;
  wire       [31:0]   _zz_88;
  wire       [0:0]    _zz_89;
  wire       [0:0]    _zz_90;
  wire       [31:0]   _zz_91;
  wire       [31:0]   _zz_92;
  wire       [31:0]   _zz_93;
  wire       [0:0]    _zz_94;
  wire       [0:0]    _zz_95;
  wire       [31:0]   _zz_96;
  wire       [31:0]   _zz_97;
  wire       [31:0]   _zz_98;
  wire       [0:0]    _zz_99;
  wire       [0:0]    _zz_100;
  wire       [31:0]   _zz_101;
  wire       [31:0]   _zz_102;
  wire       [31:0]   _zz_103;
  wire       [0:0]    _zz_104;
  wire       [0:0]    _zz_105;
  wire       [31:0]   _zz_106;
  wire       [31:0]   _zz_107;
  wire       [31:0]   _zz_108;
  wire       [0:0]    _zz_109;
  wire       [0:0]    _zz_110;
  wire       [31:0]   _zz_111;
  wire       [31:0]   _zz_112;
  wire       [31:0]   _zz_113;
  wire       [0:0]    _zz_114;
  wire       [0:0]    _zz_115;
  wire       [31:0]   _zz_116;
  wire       [31:0]   _zz_117;
  wire       [31:0]   _zz_118;
  wire       [0:0]    _zz_119;
  wire       [0:0]    _zz_120;
  wire       [31:0]   _zz_121;
  wire       [31:0]   _zz_122;
  wire       [31:0]   _zz_123;
  wire       [0:0]    _zz_124;
  wire       [0:0]    _zz_125;
  wire       [31:0]   _zz_126;
  wire       [31:0]   _zz_127;
  wire       [31:0]   _zz_128;
  wire       [0:0]    _zz_129;
  wire       [0:0]    _zz_130;
  wire       [31:0]   _zz_131;
  wire       [31:0]   _zz_132;
  wire       [31:0]   _zz_133;
  wire       [0:0]    _zz_134;
  wire       [0:0]    _zz_135;
  wire       [31:0]   _zz_136;
  wire       [31:0]   _zz_137;
  wire       [31:0]   _zz_138;
  wire       [0:0]    _zz_139;
  wire       [0:0]    _zz_140;
  wire       [31:0]   _zz_141;
  wire       [31:0]   _zz_142;
  wire       [31:0]   _zz_143;
  wire       [0:0]    _zz_144;
  wire       [0:0]    _zz_145;
  wire       [31:0]   _zz_146;
  wire       [31:0]   _zz_147;
  wire       [31:0]   _zz_148;
  wire       [0:0]    _zz_149;
  wire       [0:0]    _zz_150;
  wire       [31:0]   _zz_151;
  wire       [31:0]   _zz_152;
  wire       [31:0]   _zz_153;
  wire       [0:0]    _zz_154;
  wire       [0:0]    _zz_155;
  wire       [31:0]   _zz_156;
  wire       [31:0]   _zz_157;
  wire       [31:0]   _zz_158;
  wire       [0:0]    _zz_159;
  wire       [0:0]    _zz_160;
  wire       [31:0]   _zz_161;
  wire       [31:0]   _zz_162;
  wire       [31:0]   _zz_163;
  wire       [0:0]    _zz_164;
  wire       [0:0]    _zz_165;
  wire       [31:0]   _zz_166;
  wire       [31:0]   _zz_167;
  wire       [31:0]   _zz_168;
  wire       [0:0]    _zz_169;
  wire       [0:0]    _zz_170;
  wire       [31:0]   _zz_171;
  wire       [31:0]   _zz_172;
  wire       [31:0]   _zz_173;
  wire       [0:0]    _zz_174;
  wire       [0:0]    _zz_175;
  wire       [31:0]   _zz_176;
  wire       [31:0]   _zz_177;
  wire       [31:0]   _zz_178;
  wire       [0:0]    _zz_179;
  wire       [0:0]    _zz_180;
  wire       [31:0]   _zz_181;
  wire       [31:0]   _zz_182;
  wire       [31:0]   _zz_183;
  wire       [0:0]    _zz_184;
  wire       [0:0]    _zz_185;
  wire       [31:0]   _zz_186;
  wire       [31:0]   _zz_187;
  wire       [31:0]   _zz_188;
  wire       [0:0]    _zz_189;
  wire       [0:0]    _zz_190;
  wire       [31:0]   _zz_191;
  wire       [31:0]   _zz_192;
  wire       [31:0]   _zz_193;
  wire       [0:0]    _zz_194;
  wire       [0:0]    _zz_195;
  wire       [31:0]   _zz_196;
  wire       [31:0]   _zz_197;
  wire       [31:0]   _zz_198;
  wire       [0:0]    _zz_199;
  wire       [0:0]    _zz_200;
  wire       [31:0]   _zz_201;
  wire       [31:0]   _zz_202;
  wire       [31:0]   _zz_203;
  wire       [0:0]    _zz_204;
  wire       [0:0]    _zz_205;
  wire       [31:0]   _zz_206;
  wire       [31:0]   _zz_207;
  wire       [31:0]   _zz_208;
  wire       [0:0]    _zz_209;
  wire       [0:0]    _zz_210;
  wire       [31:0]   _zz_211;
  wire       [31:0]   _zz_212;
  wire       [31:0]   _zz_213;
  wire       [0:0]    _zz_214;
  wire       [0:0]    _zz_215;
  wire       [31:0]   _zz_216;
  wire       [31:0]   _zz_217;
  wire       [31:0]   _zz_218;
  wire       [0:0]    _zz_219;
  wire       [0:0]    _zz_220;
  wire       [31:0]   _zz_221;
  wire       [31:0]   _zz_222;
  wire       [31:0]   _zz_223;
  wire       [0:0]    _zz_224;
  wire       [0:0]    _zz_225;
  wire       [31:0]   _zz_226;
  wire       [31:0]   _zz_227;
  wire       [31:0]   _zz_228;
  wire       [0:0]    _zz_229;
  wire       [0:0]    _zz_230;
  wire       [31:0]   _zz_231;
  wire       [31:0]   _zz_232;
  wire       [31:0]   _zz_233;
  wire       [0:0]    _zz_234;
  wire       [0:0]    _zz_235;
  wire       [31:0]   _zz_236;
  wire       [31:0]   _zz_237;
  wire       [31:0]   _zz_238;
  wire       [0:0]    _zz_239;
  wire       [0:0]    _zz_240;
  wire       [31:0]   _zz_241;
  wire       [31:0]   _zz_242;
  wire       [31:0]   _zz_243;
  wire       [0:0]    _zz_244;
  wire       [0:0]    _zz_245;
  wire       [31:0]   _zz_246;
  wire       [31:0]   _zz_247;
  wire       [31:0]   _zz_248;
  wire       [0:0]    _zz_249;
  wire       [0:0]    _zz_250;
  wire       [31:0]   _zz_251;
  wire       [31:0]   _zz_252;
  wire       [31:0]   _zz_253;
  wire       [0:0]    _zz_254;
  wire       [0:0]    _zz_255;
  wire       [31:0]   _zz_256;
  wire       [31:0]   _zz_257;
  wire       [31:0]   _zz_258;
  wire       [0:0]    _zz_259;
  wire       [0:0]    _zz_260;
  wire       [31:0]   _zz_261;
  wire       [31:0]   _zz_262;
  wire       [31:0]   _zz_263;
  wire       [0:0]    _zz_264;
  wire       [0:0]    _zz_265;
  wire       [31:0]   _zz_266;
  wire       [31:0]   _zz_267;
  wire       [31:0]   _zz_268;
  wire       [0:0]    _zz_269;
  wire       [0:0]    _zz_270;
  wire       [31:0]   _zz_271;
  wire       [31:0]   _zz_272;
  wire       [31:0]   _zz_273;
  wire       [0:0]    _zz_274;
  wire       [0:0]    _zz_275;
  wire       [31:0]   _zz_276;
  wire       [31:0]   _zz_277;
  wire       [31:0]   _zz_278;
  wire       [0:0]    _zz_279;
  wire       [0:0]    _zz_280;
  wire       [31:0]   _zz_281;
  wire       [31:0]   _zz_282;
  wire       [31:0]   _zz_283;
  wire       [0:0]    _zz_284;
  wire       [0:0]    _zz_285;
  wire       [31:0]   _zz_286;
  wire       [31:0]   _zz_287;
  wire       [31:0]   _zz_288;
  wire       [0:0]    _zz_289;
  wire       [0:0]    _zz_290;
  wire       [31:0]   _zz_291;
  wire       [31:0]   _zz_292;
  wire       [31:0]   _zz_293;
  wire       [0:0]    _zz_294;
  wire       [0:0]    _zz_295;
  wire       [31:0]   _zz_296;
  wire       [31:0]   _zz_297;
  wire       [31:0]   _zz_298;
  wire       [0:0]    _zz_299;
  wire       [0:0]    _zz_300;
  wire       [31:0]   _zz_301;
  wire       [31:0]   _zz_302;
  wire       [31:0]   _zz_303;
  wire       [0:0]    _zz_304;
  wire       [0:0]    _zz_305;
  wire       [31:0]   _zz_306;
  wire       [31:0]   _zz_307;
  wire       [31:0]   _zz_308;
  wire       [0:0]    _zz_309;
  wire       [0:0]    _zz_310;
  wire       [31:0]   _zz_311;
  wire       [31:0]   _zz_312;
  wire       [31:0]   _zz_313;
  wire       [0:0]    _zz_314;
  wire       [0:0]    _zz_315;
  wire       [31:0]   _zz_316;
  wire       [31:0]   _zz_317;
  wire       [31:0]   _zz_318;
  wire       [0:0]    _zz_319;
  wire       [0:0]    _zz_320;
  wire       [31:0]   _zz_321;
  wire       [31:0]   _zz_322;
  wire       [31:0]   _zz_323;
  wire       [0:0]    _zz_324;
  wire       [0:0]    _zz_325;
  wire       [31:0]   _zz_326;
  wire       [31:0]   _zz_327;
  wire       [31:0]   _zz_328;
  wire       [0:0]    _zz_329;
  wire       [0:0]    _zz_330;
  wire       [31:0]   _zz_331;
  wire       [31:0]   _zz_332;
  wire       [31:0]   _zz_333;
  wire       [0:0]    _zz_334;
  wire       [0:0]    _zz_335;
  wire       [31:0]   _zz_336;
  wire       [31:0]   _zz_337;
  wire       [31:0]   _zz_338;
  wire       [0:0]    _zz_339;
  wire       [0:0]    _zz_340;
  wire       [31:0]   _zz_341;
  wire       [31:0]   _zz_342;
  wire       [31:0]   _zz_343;
  wire       [0:0]    _zz_344;
  wire       [0:0]    _zz_345;
  wire       [31:0]   _zz_346;
  wire       [31:0]   _zz_347;
  wire       [31:0]   _zz_348;
  wire       [0:0]    _zz_349;
  wire       [0:0]    _zz_350;
  wire       [31:0]   _zz_351;
  wire       [31:0]   _zz_352;
  wire       [31:0]   _zz_353;
  wire       [0:0]    _zz_354;
  wire       [0:0]    _zz_355;
  wire       [31:0]   _zz_356;
  wire       [31:0]   _zz_357;
  wire       [31:0]   _zz_358;
  wire       [0:0]    _zz_359;
  wire       [0:0]    _zz_360;
  wire       [31:0]   _zz_361;
  wire       [31:0]   _zz_362;
  wire       [31:0]   _zz_363;
  wire       [0:0]    _zz_364;
  wire       [0:0]    _zz_365;
  wire       [31:0]   _zz_366;
  wire       [31:0]   _zz_367;
  wire       [31:0]   _zz_368;
  wire       [0:0]    _zz_369;
  wire       [0:0]    _zz_370;
  wire       [31:0]   _zz_371;
  wire       [31:0]   _zz_372;
  wire       [31:0]   _zz_373;
  wire       [0:0]    _zz_374;
  wire       [0:0]    _zz_375;
  wire       [31:0]   _zz_376;
  wire       [31:0]   _zz_377;
  wire       [31:0]   _zz_378;
  wire       [0:0]    _zz_379;
  wire       [0:0]    _zz_380;
  wire       [31:0]   _zz_381;
  wire       [31:0]   _zz_382;
  wire       [31:0]   _zz_383;
  wire       [0:0]    _zz_384;
  wire       [0:0]    _zz_385;
  wire       [31:0]   _zz_386;
  wire       [31:0]   _zz_387;
  wire       [31:0]   _zz_388;
  wire       [0:0]    _zz_389;
  wire       [0:0]    _zz_390;
  wire       [31:0]   _zz_391;
  wire       [31:0]   _zz_392;
  wire       [31:0]   _zz_393;
  wire       [0:0]    _zz_394;
  wire       [0:0]    _zz_395;
  wire       [31:0]   _zz_396;
  wire       [31:0]   _zz_397;
  wire       [31:0]   _zz_398;
  wire       [0:0]    _zz_399;
  wire       [0:0]    _zz_400;
  reg                 current_level_willOverflow_regNext;

  assign _zz_881 = current_level_willIncrement;
  assign _zz_882 = {2'd0, _zz_881};
  assign _zz_883 = ($signed(twiddle_factor_table_0_real) + $signed(twiddle_factor_table_0_imag));
  assign _zz_884 = ($signed(_zz_3) - $signed(_zz_885));
  assign _zz_885 = ($signed(_zz_886) * $signed(twiddle_factor_table_0_imag));
  assign _zz_886 = ($signed(data_mid_1_real) + $signed(data_mid_1_imag));
  assign _zz_887 = fixTo_dout;
  assign _zz_888 = ($signed(_zz_3) + $signed(_zz_889));
  assign _zz_889 = ($signed(_zz_890) * $signed(twiddle_factor_table_0_real));
  assign _zz_890 = ($signed(data_mid_1_imag) - $signed(data_mid_1_real));
  assign _zz_891 = fixTo_1_dout;
  assign _zz_892 = _zz_893[31 : 0];
  assign _zz_893 = _zz_894;
  assign _zz_894 = ($signed(_zz_895) >>> _zz_4);
  assign _zz_895 = _zz_896;
  assign _zz_896 = ($signed(_zz_898) - $signed(_zz_1));
  assign _zz_897 = ({8'd0,data_mid_0_real} <<< 8);
  assign _zz_898 = {{8{_zz_897[23]}}, _zz_897};
  assign _zz_899 = fixTo_2_dout;
  assign _zz_900 = _zz_901[31 : 0];
  assign _zz_901 = _zz_902;
  assign _zz_902 = ($signed(_zz_903) >>> _zz_4);
  assign _zz_903 = _zz_904;
  assign _zz_904 = ($signed(_zz_906) - $signed(_zz_2));
  assign _zz_905 = ({8'd0,data_mid_0_imag} <<< 8);
  assign _zz_906 = {{8{_zz_905[23]}}, _zz_905};
  assign _zz_907 = fixTo_3_dout;
  assign _zz_908 = _zz_909[31 : 0];
  assign _zz_909 = _zz_910;
  assign _zz_910 = ($signed(_zz_911) >>> _zz_5);
  assign _zz_911 = _zz_912;
  assign _zz_912 = ($signed(_zz_914) + $signed(_zz_1));
  assign _zz_913 = ({8'd0,data_mid_0_real} <<< 8);
  assign _zz_914 = {{8{_zz_913[23]}}, _zz_913};
  assign _zz_915 = fixTo_4_dout;
  assign _zz_916 = _zz_917[31 : 0];
  assign _zz_917 = _zz_918;
  assign _zz_918 = ($signed(_zz_919) >>> _zz_5);
  assign _zz_919 = _zz_920;
  assign _zz_920 = ($signed(_zz_922) + $signed(_zz_2));
  assign _zz_921 = ({8'd0,data_mid_0_imag} <<< 8);
  assign _zz_922 = {{8{_zz_921[23]}}, _zz_921};
  assign _zz_923 = fixTo_5_dout;
  assign _zz_924 = ($signed(twiddle_factor_table_0_real) + $signed(twiddle_factor_table_0_imag));
  assign _zz_925 = ($signed(_zz_8) - $signed(_zz_926));
  assign _zz_926 = ($signed(_zz_927) * $signed(twiddle_factor_table_0_imag));
  assign _zz_927 = ($signed(data_mid_3_real) + $signed(data_mid_3_imag));
  assign _zz_928 = fixTo_6_dout;
  assign _zz_929 = ($signed(_zz_8) + $signed(_zz_930));
  assign _zz_930 = ($signed(_zz_931) * $signed(twiddle_factor_table_0_real));
  assign _zz_931 = ($signed(data_mid_3_imag) - $signed(data_mid_3_real));
  assign _zz_932 = fixTo_7_dout;
  assign _zz_933 = _zz_934[31 : 0];
  assign _zz_934 = _zz_935;
  assign _zz_935 = ($signed(_zz_936) >>> _zz_9);
  assign _zz_936 = _zz_937;
  assign _zz_937 = ($signed(_zz_939) - $signed(_zz_6));
  assign _zz_938 = ({8'd0,data_mid_2_real} <<< 8);
  assign _zz_939 = {{8{_zz_938[23]}}, _zz_938};
  assign _zz_940 = fixTo_8_dout;
  assign _zz_941 = _zz_942[31 : 0];
  assign _zz_942 = _zz_943;
  assign _zz_943 = ($signed(_zz_944) >>> _zz_9);
  assign _zz_944 = _zz_945;
  assign _zz_945 = ($signed(_zz_947) - $signed(_zz_7));
  assign _zz_946 = ({8'd0,data_mid_2_imag} <<< 8);
  assign _zz_947 = {{8{_zz_946[23]}}, _zz_946};
  assign _zz_948 = fixTo_9_dout;
  assign _zz_949 = _zz_950[31 : 0];
  assign _zz_950 = _zz_951;
  assign _zz_951 = ($signed(_zz_952) >>> _zz_10);
  assign _zz_952 = _zz_953;
  assign _zz_953 = ($signed(_zz_955) + $signed(_zz_6));
  assign _zz_954 = ({8'd0,data_mid_2_real} <<< 8);
  assign _zz_955 = {{8{_zz_954[23]}}, _zz_954};
  assign _zz_956 = fixTo_10_dout;
  assign _zz_957 = _zz_958[31 : 0];
  assign _zz_958 = _zz_959;
  assign _zz_959 = ($signed(_zz_960) >>> _zz_10);
  assign _zz_960 = _zz_961;
  assign _zz_961 = ($signed(_zz_963) + $signed(_zz_7));
  assign _zz_962 = ({8'd0,data_mid_2_imag} <<< 8);
  assign _zz_963 = {{8{_zz_962[23]}}, _zz_962};
  assign _zz_964 = fixTo_11_dout;
  assign _zz_965 = ($signed(twiddle_factor_table_0_real) + $signed(twiddle_factor_table_0_imag));
  assign _zz_966 = ($signed(_zz_13) - $signed(_zz_967));
  assign _zz_967 = ($signed(_zz_968) * $signed(twiddle_factor_table_0_imag));
  assign _zz_968 = ($signed(data_mid_5_real) + $signed(data_mid_5_imag));
  assign _zz_969 = fixTo_12_dout;
  assign _zz_970 = ($signed(_zz_13) + $signed(_zz_971));
  assign _zz_971 = ($signed(_zz_972) * $signed(twiddle_factor_table_0_real));
  assign _zz_972 = ($signed(data_mid_5_imag) - $signed(data_mid_5_real));
  assign _zz_973 = fixTo_13_dout;
  assign _zz_974 = _zz_975[31 : 0];
  assign _zz_975 = _zz_976;
  assign _zz_976 = ($signed(_zz_977) >>> _zz_14);
  assign _zz_977 = _zz_978;
  assign _zz_978 = ($signed(_zz_980) - $signed(_zz_11));
  assign _zz_979 = ({8'd0,data_mid_4_real} <<< 8);
  assign _zz_980 = {{8{_zz_979[23]}}, _zz_979};
  assign _zz_981 = fixTo_14_dout;
  assign _zz_982 = _zz_983[31 : 0];
  assign _zz_983 = _zz_984;
  assign _zz_984 = ($signed(_zz_985) >>> _zz_14);
  assign _zz_985 = _zz_986;
  assign _zz_986 = ($signed(_zz_988) - $signed(_zz_12));
  assign _zz_987 = ({8'd0,data_mid_4_imag} <<< 8);
  assign _zz_988 = {{8{_zz_987[23]}}, _zz_987};
  assign _zz_989 = fixTo_15_dout;
  assign _zz_990 = _zz_991[31 : 0];
  assign _zz_991 = _zz_992;
  assign _zz_992 = ($signed(_zz_993) >>> _zz_15);
  assign _zz_993 = _zz_994;
  assign _zz_994 = ($signed(_zz_996) + $signed(_zz_11));
  assign _zz_995 = ({8'd0,data_mid_4_real} <<< 8);
  assign _zz_996 = {{8{_zz_995[23]}}, _zz_995};
  assign _zz_997 = fixTo_16_dout;
  assign _zz_998 = _zz_999[31 : 0];
  assign _zz_999 = _zz_1000;
  assign _zz_1000 = ($signed(_zz_1001) >>> _zz_15);
  assign _zz_1001 = _zz_1002;
  assign _zz_1002 = ($signed(_zz_1004) + $signed(_zz_12));
  assign _zz_1003 = ({8'd0,data_mid_4_imag} <<< 8);
  assign _zz_1004 = {{8{_zz_1003[23]}}, _zz_1003};
  assign _zz_1005 = fixTo_17_dout;
  assign _zz_1006 = ($signed(twiddle_factor_table_0_real) + $signed(twiddle_factor_table_0_imag));
  assign _zz_1007 = ($signed(_zz_18) - $signed(_zz_1008));
  assign _zz_1008 = ($signed(_zz_1009) * $signed(twiddle_factor_table_0_imag));
  assign _zz_1009 = ($signed(data_mid_7_real) + $signed(data_mid_7_imag));
  assign _zz_1010 = fixTo_18_dout;
  assign _zz_1011 = ($signed(_zz_18) + $signed(_zz_1012));
  assign _zz_1012 = ($signed(_zz_1013) * $signed(twiddle_factor_table_0_real));
  assign _zz_1013 = ($signed(data_mid_7_imag) - $signed(data_mid_7_real));
  assign _zz_1014 = fixTo_19_dout;
  assign _zz_1015 = _zz_1016[31 : 0];
  assign _zz_1016 = _zz_1017;
  assign _zz_1017 = ($signed(_zz_1018) >>> _zz_19);
  assign _zz_1018 = _zz_1019;
  assign _zz_1019 = ($signed(_zz_1021) - $signed(_zz_16));
  assign _zz_1020 = ({8'd0,data_mid_6_real} <<< 8);
  assign _zz_1021 = {{8{_zz_1020[23]}}, _zz_1020};
  assign _zz_1022 = fixTo_20_dout;
  assign _zz_1023 = _zz_1024[31 : 0];
  assign _zz_1024 = _zz_1025;
  assign _zz_1025 = ($signed(_zz_1026) >>> _zz_19);
  assign _zz_1026 = _zz_1027;
  assign _zz_1027 = ($signed(_zz_1029) - $signed(_zz_17));
  assign _zz_1028 = ({8'd0,data_mid_6_imag} <<< 8);
  assign _zz_1029 = {{8{_zz_1028[23]}}, _zz_1028};
  assign _zz_1030 = fixTo_21_dout;
  assign _zz_1031 = _zz_1032[31 : 0];
  assign _zz_1032 = _zz_1033;
  assign _zz_1033 = ($signed(_zz_1034) >>> _zz_20);
  assign _zz_1034 = _zz_1035;
  assign _zz_1035 = ($signed(_zz_1037) + $signed(_zz_16));
  assign _zz_1036 = ({8'd0,data_mid_6_real} <<< 8);
  assign _zz_1037 = {{8{_zz_1036[23]}}, _zz_1036};
  assign _zz_1038 = fixTo_22_dout;
  assign _zz_1039 = _zz_1040[31 : 0];
  assign _zz_1040 = _zz_1041;
  assign _zz_1041 = ($signed(_zz_1042) >>> _zz_20);
  assign _zz_1042 = _zz_1043;
  assign _zz_1043 = ($signed(_zz_1045) + $signed(_zz_17));
  assign _zz_1044 = ({8'd0,data_mid_6_imag} <<< 8);
  assign _zz_1045 = {{8{_zz_1044[23]}}, _zz_1044};
  assign _zz_1046 = fixTo_23_dout;
  assign _zz_1047 = ($signed(twiddle_factor_table_0_real) + $signed(twiddle_factor_table_0_imag));
  assign _zz_1048 = ($signed(_zz_23) - $signed(_zz_1049));
  assign _zz_1049 = ($signed(_zz_1050) * $signed(twiddle_factor_table_0_imag));
  assign _zz_1050 = ($signed(data_mid_9_real) + $signed(data_mid_9_imag));
  assign _zz_1051 = fixTo_24_dout;
  assign _zz_1052 = ($signed(_zz_23) + $signed(_zz_1053));
  assign _zz_1053 = ($signed(_zz_1054) * $signed(twiddle_factor_table_0_real));
  assign _zz_1054 = ($signed(data_mid_9_imag) - $signed(data_mid_9_real));
  assign _zz_1055 = fixTo_25_dout;
  assign _zz_1056 = _zz_1057[31 : 0];
  assign _zz_1057 = _zz_1058;
  assign _zz_1058 = ($signed(_zz_1059) >>> _zz_24);
  assign _zz_1059 = _zz_1060;
  assign _zz_1060 = ($signed(_zz_1062) - $signed(_zz_21));
  assign _zz_1061 = ({8'd0,data_mid_8_real} <<< 8);
  assign _zz_1062 = {{8{_zz_1061[23]}}, _zz_1061};
  assign _zz_1063 = fixTo_26_dout;
  assign _zz_1064 = _zz_1065[31 : 0];
  assign _zz_1065 = _zz_1066;
  assign _zz_1066 = ($signed(_zz_1067) >>> _zz_24);
  assign _zz_1067 = _zz_1068;
  assign _zz_1068 = ($signed(_zz_1070) - $signed(_zz_22));
  assign _zz_1069 = ({8'd0,data_mid_8_imag} <<< 8);
  assign _zz_1070 = {{8{_zz_1069[23]}}, _zz_1069};
  assign _zz_1071 = fixTo_27_dout;
  assign _zz_1072 = _zz_1073[31 : 0];
  assign _zz_1073 = _zz_1074;
  assign _zz_1074 = ($signed(_zz_1075) >>> _zz_25);
  assign _zz_1075 = _zz_1076;
  assign _zz_1076 = ($signed(_zz_1078) + $signed(_zz_21));
  assign _zz_1077 = ({8'd0,data_mid_8_real} <<< 8);
  assign _zz_1078 = {{8{_zz_1077[23]}}, _zz_1077};
  assign _zz_1079 = fixTo_28_dout;
  assign _zz_1080 = _zz_1081[31 : 0];
  assign _zz_1081 = _zz_1082;
  assign _zz_1082 = ($signed(_zz_1083) >>> _zz_25);
  assign _zz_1083 = _zz_1084;
  assign _zz_1084 = ($signed(_zz_1086) + $signed(_zz_22));
  assign _zz_1085 = ({8'd0,data_mid_8_imag} <<< 8);
  assign _zz_1086 = {{8{_zz_1085[23]}}, _zz_1085};
  assign _zz_1087 = fixTo_29_dout;
  assign _zz_1088 = ($signed(twiddle_factor_table_0_real) + $signed(twiddle_factor_table_0_imag));
  assign _zz_1089 = ($signed(_zz_28) - $signed(_zz_1090));
  assign _zz_1090 = ($signed(_zz_1091) * $signed(twiddle_factor_table_0_imag));
  assign _zz_1091 = ($signed(data_mid_11_real) + $signed(data_mid_11_imag));
  assign _zz_1092 = fixTo_30_dout;
  assign _zz_1093 = ($signed(_zz_28) + $signed(_zz_1094));
  assign _zz_1094 = ($signed(_zz_1095) * $signed(twiddle_factor_table_0_real));
  assign _zz_1095 = ($signed(data_mid_11_imag) - $signed(data_mid_11_real));
  assign _zz_1096 = fixTo_31_dout;
  assign _zz_1097 = _zz_1098[31 : 0];
  assign _zz_1098 = _zz_1099;
  assign _zz_1099 = ($signed(_zz_1100) >>> _zz_29);
  assign _zz_1100 = _zz_1101;
  assign _zz_1101 = ($signed(_zz_1103) - $signed(_zz_26));
  assign _zz_1102 = ({8'd0,data_mid_10_real} <<< 8);
  assign _zz_1103 = {{8{_zz_1102[23]}}, _zz_1102};
  assign _zz_1104 = fixTo_32_dout;
  assign _zz_1105 = _zz_1106[31 : 0];
  assign _zz_1106 = _zz_1107;
  assign _zz_1107 = ($signed(_zz_1108) >>> _zz_29);
  assign _zz_1108 = _zz_1109;
  assign _zz_1109 = ($signed(_zz_1111) - $signed(_zz_27));
  assign _zz_1110 = ({8'd0,data_mid_10_imag} <<< 8);
  assign _zz_1111 = {{8{_zz_1110[23]}}, _zz_1110};
  assign _zz_1112 = fixTo_33_dout;
  assign _zz_1113 = _zz_1114[31 : 0];
  assign _zz_1114 = _zz_1115;
  assign _zz_1115 = ($signed(_zz_1116) >>> _zz_30);
  assign _zz_1116 = _zz_1117;
  assign _zz_1117 = ($signed(_zz_1119) + $signed(_zz_26));
  assign _zz_1118 = ({8'd0,data_mid_10_real} <<< 8);
  assign _zz_1119 = {{8{_zz_1118[23]}}, _zz_1118};
  assign _zz_1120 = fixTo_34_dout;
  assign _zz_1121 = _zz_1122[31 : 0];
  assign _zz_1122 = _zz_1123;
  assign _zz_1123 = ($signed(_zz_1124) >>> _zz_30);
  assign _zz_1124 = _zz_1125;
  assign _zz_1125 = ($signed(_zz_1127) + $signed(_zz_27));
  assign _zz_1126 = ({8'd0,data_mid_10_imag} <<< 8);
  assign _zz_1127 = {{8{_zz_1126[23]}}, _zz_1126};
  assign _zz_1128 = fixTo_35_dout;
  assign _zz_1129 = ($signed(twiddle_factor_table_0_real) + $signed(twiddle_factor_table_0_imag));
  assign _zz_1130 = ($signed(_zz_33) - $signed(_zz_1131));
  assign _zz_1131 = ($signed(_zz_1132) * $signed(twiddle_factor_table_0_imag));
  assign _zz_1132 = ($signed(data_mid_13_real) + $signed(data_mid_13_imag));
  assign _zz_1133 = fixTo_36_dout;
  assign _zz_1134 = ($signed(_zz_33) + $signed(_zz_1135));
  assign _zz_1135 = ($signed(_zz_1136) * $signed(twiddle_factor_table_0_real));
  assign _zz_1136 = ($signed(data_mid_13_imag) - $signed(data_mid_13_real));
  assign _zz_1137 = fixTo_37_dout;
  assign _zz_1138 = _zz_1139[31 : 0];
  assign _zz_1139 = _zz_1140;
  assign _zz_1140 = ($signed(_zz_1141) >>> _zz_34);
  assign _zz_1141 = _zz_1142;
  assign _zz_1142 = ($signed(_zz_1144) - $signed(_zz_31));
  assign _zz_1143 = ({8'd0,data_mid_12_real} <<< 8);
  assign _zz_1144 = {{8{_zz_1143[23]}}, _zz_1143};
  assign _zz_1145 = fixTo_38_dout;
  assign _zz_1146 = _zz_1147[31 : 0];
  assign _zz_1147 = _zz_1148;
  assign _zz_1148 = ($signed(_zz_1149) >>> _zz_34);
  assign _zz_1149 = _zz_1150;
  assign _zz_1150 = ($signed(_zz_1152) - $signed(_zz_32));
  assign _zz_1151 = ({8'd0,data_mid_12_imag} <<< 8);
  assign _zz_1152 = {{8{_zz_1151[23]}}, _zz_1151};
  assign _zz_1153 = fixTo_39_dout;
  assign _zz_1154 = _zz_1155[31 : 0];
  assign _zz_1155 = _zz_1156;
  assign _zz_1156 = ($signed(_zz_1157) >>> _zz_35);
  assign _zz_1157 = _zz_1158;
  assign _zz_1158 = ($signed(_zz_1160) + $signed(_zz_31));
  assign _zz_1159 = ({8'd0,data_mid_12_real} <<< 8);
  assign _zz_1160 = {{8{_zz_1159[23]}}, _zz_1159};
  assign _zz_1161 = fixTo_40_dout;
  assign _zz_1162 = _zz_1163[31 : 0];
  assign _zz_1163 = _zz_1164;
  assign _zz_1164 = ($signed(_zz_1165) >>> _zz_35);
  assign _zz_1165 = _zz_1166;
  assign _zz_1166 = ($signed(_zz_1168) + $signed(_zz_32));
  assign _zz_1167 = ({8'd0,data_mid_12_imag} <<< 8);
  assign _zz_1168 = {{8{_zz_1167[23]}}, _zz_1167};
  assign _zz_1169 = fixTo_41_dout;
  assign _zz_1170 = ($signed(twiddle_factor_table_0_real) + $signed(twiddle_factor_table_0_imag));
  assign _zz_1171 = ($signed(_zz_38) - $signed(_zz_1172));
  assign _zz_1172 = ($signed(_zz_1173) * $signed(twiddle_factor_table_0_imag));
  assign _zz_1173 = ($signed(data_mid_15_real) + $signed(data_mid_15_imag));
  assign _zz_1174 = fixTo_42_dout;
  assign _zz_1175 = ($signed(_zz_38) + $signed(_zz_1176));
  assign _zz_1176 = ($signed(_zz_1177) * $signed(twiddle_factor_table_0_real));
  assign _zz_1177 = ($signed(data_mid_15_imag) - $signed(data_mid_15_real));
  assign _zz_1178 = fixTo_43_dout;
  assign _zz_1179 = _zz_1180[31 : 0];
  assign _zz_1180 = _zz_1181;
  assign _zz_1181 = ($signed(_zz_1182) >>> _zz_39);
  assign _zz_1182 = _zz_1183;
  assign _zz_1183 = ($signed(_zz_1185) - $signed(_zz_36));
  assign _zz_1184 = ({8'd0,data_mid_14_real} <<< 8);
  assign _zz_1185 = {{8{_zz_1184[23]}}, _zz_1184};
  assign _zz_1186 = fixTo_44_dout;
  assign _zz_1187 = _zz_1188[31 : 0];
  assign _zz_1188 = _zz_1189;
  assign _zz_1189 = ($signed(_zz_1190) >>> _zz_39);
  assign _zz_1190 = _zz_1191;
  assign _zz_1191 = ($signed(_zz_1193) - $signed(_zz_37));
  assign _zz_1192 = ({8'd0,data_mid_14_imag} <<< 8);
  assign _zz_1193 = {{8{_zz_1192[23]}}, _zz_1192};
  assign _zz_1194 = fixTo_45_dout;
  assign _zz_1195 = _zz_1196[31 : 0];
  assign _zz_1196 = _zz_1197;
  assign _zz_1197 = ($signed(_zz_1198) >>> _zz_40);
  assign _zz_1198 = _zz_1199;
  assign _zz_1199 = ($signed(_zz_1201) + $signed(_zz_36));
  assign _zz_1200 = ({8'd0,data_mid_14_real} <<< 8);
  assign _zz_1201 = {{8{_zz_1200[23]}}, _zz_1200};
  assign _zz_1202 = fixTo_46_dout;
  assign _zz_1203 = _zz_1204[31 : 0];
  assign _zz_1204 = _zz_1205;
  assign _zz_1205 = ($signed(_zz_1206) >>> _zz_40);
  assign _zz_1206 = _zz_1207;
  assign _zz_1207 = ($signed(_zz_1209) + $signed(_zz_37));
  assign _zz_1208 = ({8'd0,data_mid_14_imag} <<< 8);
  assign _zz_1209 = {{8{_zz_1208[23]}}, _zz_1208};
  assign _zz_1210 = fixTo_47_dout;
  assign _zz_1211 = ($signed(twiddle_factor_table_0_real) + $signed(twiddle_factor_table_0_imag));
  assign _zz_1212 = ($signed(_zz_43) - $signed(_zz_1213));
  assign _zz_1213 = ($signed(_zz_1214) * $signed(twiddle_factor_table_0_imag));
  assign _zz_1214 = ($signed(data_mid_17_real) + $signed(data_mid_17_imag));
  assign _zz_1215 = fixTo_48_dout;
  assign _zz_1216 = ($signed(_zz_43) + $signed(_zz_1217));
  assign _zz_1217 = ($signed(_zz_1218) * $signed(twiddle_factor_table_0_real));
  assign _zz_1218 = ($signed(data_mid_17_imag) - $signed(data_mid_17_real));
  assign _zz_1219 = fixTo_49_dout;
  assign _zz_1220 = _zz_1221[31 : 0];
  assign _zz_1221 = _zz_1222;
  assign _zz_1222 = ($signed(_zz_1223) >>> _zz_44);
  assign _zz_1223 = _zz_1224;
  assign _zz_1224 = ($signed(_zz_1226) - $signed(_zz_41));
  assign _zz_1225 = ({8'd0,data_mid_16_real} <<< 8);
  assign _zz_1226 = {{8{_zz_1225[23]}}, _zz_1225};
  assign _zz_1227 = fixTo_50_dout;
  assign _zz_1228 = _zz_1229[31 : 0];
  assign _zz_1229 = _zz_1230;
  assign _zz_1230 = ($signed(_zz_1231) >>> _zz_44);
  assign _zz_1231 = _zz_1232;
  assign _zz_1232 = ($signed(_zz_1234) - $signed(_zz_42));
  assign _zz_1233 = ({8'd0,data_mid_16_imag} <<< 8);
  assign _zz_1234 = {{8{_zz_1233[23]}}, _zz_1233};
  assign _zz_1235 = fixTo_51_dout;
  assign _zz_1236 = _zz_1237[31 : 0];
  assign _zz_1237 = _zz_1238;
  assign _zz_1238 = ($signed(_zz_1239) >>> _zz_45);
  assign _zz_1239 = _zz_1240;
  assign _zz_1240 = ($signed(_zz_1242) + $signed(_zz_41));
  assign _zz_1241 = ({8'd0,data_mid_16_real} <<< 8);
  assign _zz_1242 = {{8{_zz_1241[23]}}, _zz_1241};
  assign _zz_1243 = fixTo_52_dout;
  assign _zz_1244 = _zz_1245[31 : 0];
  assign _zz_1245 = _zz_1246;
  assign _zz_1246 = ($signed(_zz_1247) >>> _zz_45);
  assign _zz_1247 = _zz_1248;
  assign _zz_1248 = ($signed(_zz_1250) + $signed(_zz_42));
  assign _zz_1249 = ({8'd0,data_mid_16_imag} <<< 8);
  assign _zz_1250 = {{8{_zz_1249[23]}}, _zz_1249};
  assign _zz_1251 = fixTo_53_dout;
  assign _zz_1252 = ($signed(twiddle_factor_table_0_real) + $signed(twiddle_factor_table_0_imag));
  assign _zz_1253 = ($signed(_zz_48) - $signed(_zz_1254));
  assign _zz_1254 = ($signed(_zz_1255) * $signed(twiddle_factor_table_0_imag));
  assign _zz_1255 = ($signed(data_mid_19_real) + $signed(data_mid_19_imag));
  assign _zz_1256 = fixTo_54_dout;
  assign _zz_1257 = ($signed(_zz_48) + $signed(_zz_1258));
  assign _zz_1258 = ($signed(_zz_1259) * $signed(twiddle_factor_table_0_real));
  assign _zz_1259 = ($signed(data_mid_19_imag) - $signed(data_mid_19_real));
  assign _zz_1260 = fixTo_55_dout;
  assign _zz_1261 = _zz_1262[31 : 0];
  assign _zz_1262 = _zz_1263;
  assign _zz_1263 = ($signed(_zz_1264) >>> _zz_49);
  assign _zz_1264 = _zz_1265;
  assign _zz_1265 = ($signed(_zz_1267) - $signed(_zz_46));
  assign _zz_1266 = ({8'd0,data_mid_18_real} <<< 8);
  assign _zz_1267 = {{8{_zz_1266[23]}}, _zz_1266};
  assign _zz_1268 = fixTo_56_dout;
  assign _zz_1269 = _zz_1270[31 : 0];
  assign _zz_1270 = _zz_1271;
  assign _zz_1271 = ($signed(_zz_1272) >>> _zz_49);
  assign _zz_1272 = _zz_1273;
  assign _zz_1273 = ($signed(_zz_1275) - $signed(_zz_47));
  assign _zz_1274 = ({8'd0,data_mid_18_imag} <<< 8);
  assign _zz_1275 = {{8{_zz_1274[23]}}, _zz_1274};
  assign _zz_1276 = fixTo_57_dout;
  assign _zz_1277 = _zz_1278[31 : 0];
  assign _zz_1278 = _zz_1279;
  assign _zz_1279 = ($signed(_zz_1280) >>> _zz_50);
  assign _zz_1280 = _zz_1281;
  assign _zz_1281 = ($signed(_zz_1283) + $signed(_zz_46));
  assign _zz_1282 = ({8'd0,data_mid_18_real} <<< 8);
  assign _zz_1283 = {{8{_zz_1282[23]}}, _zz_1282};
  assign _zz_1284 = fixTo_58_dout;
  assign _zz_1285 = _zz_1286[31 : 0];
  assign _zz_1286 = _zz_1287;
  assign _zz_1287 = ($signed(_zz_1288) >>> _zz_50);
  assign _zz_1288 = _zz_1289;
  assign _zz_1289 = ($signed(_zz_1291) + $signed(_zz_47));
  assign _zz_1290 = ({8'd0,data_mid_18_imag} <<< 8);
  assign _zz_1291 = {{8{_zz_1290[23]}}, _zz_1290};
  assign _zz_1292 = fixTo_59_dout;
  assign _zz_1293 = ($signed(twiddle_factor_table_0_real) + $signed(twiddle_factor_table_0_imag));
  assign _zz_1294 = ($signed(_zz_53) - $signed(_zz_1295));
  assign _zz_1295 = ($signed(_zz_1296) * $signed(twiddle_factor_table_0_imag));
  assign _zz_1296 = ($signed(data_mid_21_real) + $signed(data_mid_21_imag));
  assign _zz_1297 = fixTo_60_dout;
  assign _zz_1298 = ($signed(_zz_53) + $signed(_zz_1299));
  assign _zz_1299 = ($signed(_zz_1300) * $signed(twiddle_factor_table_0_real));
  assign _zz_1300 = ($signed(data_mid_21_imag) - $signed(data_mid_21_real));
  assign _zz_1301 = fixTo_61_dout;
  assign _zz_1302 = _zz_1303[31 : 0];
  assign _zz_1303 = _zz_1304;
  assign _zz_1304 = ($signed(_zz_1305) >>> _zz_54);
  assign _zz_1305 = _zz_1306;
  assign _zz_1306 = ($signed(_zz_1308) - $signed(_zz_51));
  assign _zz_1307 = ({8'd0,data_mid_20_real} <<< 8);
  assign _zz_1308 = {{8{_zz_1307[23]}}, _zz_1307};
  assign _zz_1309 = fixTo_62_dout;
  assign _zz_1310 = _zz_1311[31 : 0];
  assign _zz_1311 = _zz_1312;
  assign _zz_1312 = ($signed(_zz_1313) >>> _zz_54);
  assign _zz_1313 = _zz_1314;
  assign _zz_1314 = ($signed(_zz_1316) - $signed(_zz_52));
  assign _zz_1315 = ({8'd0,data_mid_20_imag} <<< 8);
  assign _zz_1316 = {{8{_zz_1315[23]}}, _zz_1315};
  assign _zz_1317 = fixTo_63_dout;
  assign _zz_1318 = _zz_1319[31 : 0];
  assign _zz_1319 = _zz_1320;
  assign _zz_1320 = ($signed(_zz_1321) >>> _zz_55);
  assign _zz_1321 = _zz_1322;
  assign _zz_1322 = ($signed(_zz_1324) + $signed(_zz_51));
  assign _zz_1323 = ({8'd0,data_mid_20_real} <<< 8);
  assign _zz_1324 = {{8{_zz_1323[23]}}, _zz_1323};
  assign _zz_1325 = fixTo_64_dout;
  assign _zz_1326 = _zz_1327[31 : 0];
  assign _zz_1327 = _zz_1328;
  assign _zz_1328 = ($signed(_zz_1329) >>> _zz_55);
  assign _zz_1329 = _zz_1330;
  assign _zz_1330 = ($signed(_zz_1332) + $signed(_zz_52));
  assign _zz_1331 = ({8'd0,data_mid_20_imag} <<< 8);
  assign _zz_1332 = {{8{_zz_1331[23]}}, _zz_1331};
  assign _zz_1333 = fixTo_65_dout;
  assign _zz_1334 = ($signed(twiddle_factor_table_0_real) + $signed(twiddle_factor_table_0_imag));
  assign _zz_1335 = ($signed(_zz_58) - $signed(_zz_1336));
  assign _zz_1336 = ($signed(_zz_1337) * $signed(twiddle_factor_table_0_imag));
  assign _zz_1337 = ($signed(data_mid_23_real) + $signed(data_mid_23_imag));
  assign _zz_1338 = fixTo_66_dout;
  assign _zz_1339 = ($signed(_zz_58) + $signed(_zz_1340));
  assign _zz_1340 = ($signed(_zz_1341) * $signed(twiddle_factor_table_0_real));
  assign _zz_1341 = ($signed(data_mid_23_imag) - $signed(data_mid_23_real));
  assign _zz_1342 = fixTo_67_dout;
  assign _zz_1343 = _zz_1344[31 : 0];
  assign _zz_1344 = _zz_1345;
  assign _zz_1345 = ($signed(_zz_1346) >>> _zz_59);
  assign _zz_1346 = _zz_1347;
  assign _zz_1347 = ($signed(_zz_1349) - $signed(_zz_56));
  assign _zz_1348 = ({8'd0,data_mid_22_real} <<< 8);
  assign _zz_1349 = {{8{_zz_1348[23]}}, _zz_1348};
  assign _zz_1350 = fixTo_68_dout;
  assign _zz_1351 = _zz_1352[31 : 0];
  assign _zz_1352 = _zz_1353;
  assign _zz_1353 = ($signed(_zz_1354) >>> _zz_59);
  assign _zz_1354 = _zz_1355;
  assign _zz_1355 = ($signed(_zz_1357) - $signed(_zz_57));
  assign _zz_1356 = ({8'd0,data_mid_22_imag} <<< 8);
  assign _zz_1357 = {{8{_zz_1356[23]}}, _zz_1356};
  assign _zz_1358 = fixTo_69_dout;
  assign _zz_1359 = _zz_1360[31 : 0];
  assign _zz_1360 = _zz_1361;
  assign _zz_1361 = ($signed(_zz_1362) >>> _zz_60);
  assign _zz_1362 = _zz_1363;
  assign _zz_1363 = ($signed(_zz_1365) + $signed(_zz_56));
  assign _zz_1364 = ({8'd0,data_mid_22_real} <<< 8);
  assign _zz_1365 = {{8{_zz_1364[23]}}, _zz_1364};
  assign _zz_1366 = fixTo_70_dout;
  assign _zz_1367 = _zz_1368[31 : 0];
  assign _zz_1368 = _zz_1369;
  assign _zz_1369 = ($signed(_zz_1370) >>> _zz_60);
  assign _zz_1370 = _zz_1371;
  assign _zz_1371 = ($signed(_zz_1373) + $signed(_zz_57));
  assign _zz_1372 = ({8'd0,data_mid_22_imag} <<< 8);
  assign _zz_1373 = {{8{_zz_1372[23]}}, _zz_1372};
  assign _zz_1374 = fixTo_71_dout;
  assign _zz_1375 = ($signed(twiddle_factor_table_0_real) + $signed(twiddle_factor_table_0_imag));
  assign _zz_1376 = ($signed(_zz_63) - $signed(_zz_1377));
  assign _zz_1377 = ($signed(_zz_1378) * $signed(twiddle_factor_table_0_imag));
  assign _zz_1378 = ($signed(data_mid_25_real) + $signed(data_mid_25_imag));
  assign _zz_1379 = fixTo_72_dout;
  assign _zz_1380 = ($signed(_zz_63) + $signed(_zz_1381));
  assign _zz_1381 = ($signed(_zz_1382) * $signed(twiddle_factor_table_0_real));
  assign _zz_1382 = ($signed(data_mid_25_imag) - $signed(data_mid_25_real));
  assign _zz_1383 = fixTo_73_dout;
  assign _zz_1384 = _zz_1385[31 : 0];
  assign _zz_1385 = _zz_1386;
  assign _zz_1386 = ($signed(_zz_1387) >>> _zz_64);
  assign _zz_1387 = _zz_1388;
  assign _zz_1388 = ($signed(_zz_1390) - $signed(_zz_61));
  assign _zz_1389 = ({8'd0,data_mid_24_real} <<< 8);
  assign _zz_1390 = {{8{_zz_1389[23]}}, _zz_1389};
  assign _zz_1391 = fixTo_74_dout;
  assign _zz_1392 = _zz_1393[31 : 0];
  assign _zz_1393 = _zz_1394;
  assign _zz_1394 = ($signed(_zz_1395) >>> _zz_64);
  assign _zz_1395 = _zz_1396;
  assign _zz_1396 = ($signed(_zz_1398) - $signed(_zz_62));
  assign _zz_1397 = ({8'd0,data_mid_24_imag} <<< 8);
  assign _zz_1398 = {{8{_zz_1397[23]}}, _zz_1397};
  assign _zz_1399 = fixTo_75_dout;
  assign _zz_1400 = _zz_1401[31 : 0];
  assign _zz_1401 = _zz_1402;
  assign _zz_1402 = ($signed(_zz_1403) >>> _zz_65);
  assign _zz_1403 = _zz_1404;
  assign _zz_1404 = ($signed(_zz_1406) + $signed(_zz_61));
  assign _zz_1405 = ({8'd0,data_mid_24_real} <<< 8);
  assign _zz_1406 = {{8{_zz_1405[23]}}, _zz_1405};
  assign _zz_1407 = fixTo_76_dout;
  assign _zz_1408 = _zz_1409[31 : 0];
  assign _zz_1409 = _zz_1410;
  assign _zz_1410 = ($signed(_zz_1411) >>> _zz_65);
  assign _zz_1411 = _zz_1412;
  assign _zz_1412 = ($signed(_zz_1414) + $signed(_zz_62));
  assign _zz_1413 = ({8'd0,data_mid_24_imag} <<< 8);
  assign _zz_1414 = {{8{_zz_1413[23]}}, _zz_1413};
  assign _zz_1415 = fixTo_77_dout;
  assign _zz_1416 = ($signed(twiddle_factor_table_0_real) + $signed(twiddle_factor_table_0_imag));
  assign _zz_1417 = ($signed(_zz_68) - $signed(_zz_1418));
  assign _zz_1418 = ($signed(_zz_1419) * $signed(twiddle_factor_table_0_imag));
  assign _zz_1419 = ($signed(data_mid_27_real) + $signed(data_mid_27_imag));
  assign _zz_1420 = fixTo_78_dout;
  assign _zz_1421 = ($signed(_zz_68) + $signed(_zz_1422));
  assign _zz_1422 = ($signed(_zz_1423) * $signed(twiddle_factor_table_0_real));
  assign _zz_1423 = ($signed(data_mid_27_imag) - $signed(data_mid_27_real));
  assign _zz_1424 = fixTo_79_dout;
  assign _zz_1425 = _zz_1426[31 : 0];
  assign _zz_1426 = _zz_1427;
  assign _zz_1427 = ($signed(_zz_1428) >>> _zz_69);
  assign _zz_1428 = _zz_1429;
  assign _zz_1429 = ($signed(_zz_1431) - $signed(_zz_66));
  assign _zz_1430 = ({8'd0,data_mid_26_real} <<< 8);
  assign _zz_1431 = {{8{_zz_1430[23]}}, _zz_1430};
  assign _zz_1432 = fixTo_80_dout;
  assign _zz_1433 = _zz_1434[31 : 0];
  assign _zz_1434 = _zz_1435;
  assign _zz_1435 = ($signed(_zz_1436) >>> _zz_69);
  assign _zz_1436 = _zz_1437;
  assign _zz_1437 = ($signed(_zz_1439) - $signed(_zz_67));
  assign _zz_1438 = ({8'd0,data_mid_26_imag} <<< 8);
  assign _zz_1439 = {{8{_zz_1438[23]}}, _zz_1438};
  assign _zz_1440 = fixTo_81_dout;
  assign _zz_1441 = _zz_1442[31 : 0];
  assign _zz_1442 = _zz_1443;
  assign _zz_1443 = ($signed(_zz_1444) >>> _zz_70);
  assign _zz_1444 = _zz_1445;
  assign _zz_1445 = ($signed(_zz_1447) + $signed(_zz_66));
  assign _zz_1446 = ({8'd0,data_mid_26_real} <<< 8);
  assign _zz_1447 = {{8{_zz_1446[23]}}, _zz_1446};
  assign _zz_1448 = fixTo_82_dout;
  assign _zz_1449 = _zz_1450[31 : 0];
  assign _zz_1450 = _zz_1451;
  assign _zz_1451 = ($signed(_zz_1452) >>> _zz_70);
  assign _zz_1452 = _zz_1453;
  assign _zz_1453 = ($signed(_zz_1455) + $signed(_zz_67));
  assign _zz_1454 = ({8'd0,data_mid_26_imag} <<< 8);
  assign _zz_1455 = {{8{_zz_1454[23]}}, _zz_1454};
  assign _zz_1456 = fixTo_83_dout;
  assign _zz_1457 = ($signed(twiddle_factor_table_0_real) + $signed(twiddle_factor_table_0_imag));
  assign _zz_1458 = ($signed(_zz_73) - $signed(_zz_1459));
  assign _zz_1459 = ($signed(_zz_1460) * $signed(twiddle_factor_table_0_imag));
  assign _zz_1460 = ($signed(data_mid_29_real) + $signed(data_mid_29_imag));
  assign _zz_1461 = fixTo_84_dout;
  assign _zz_1462 = ($signed(_zz_73) + $signed(_zz_1463));
  assign _zz_1463 = ($signed(_zz_1464) * $signed(twiddle_factor_table_0_real));
  assign _zz_1464 = ($signed(data_mid_29_imag) - $signed(data_mid_29_real));
  assign _zz_1465 = fixTo_85_dout;
  assign _zz_1466 = _zz_1467[31 : 0];
  assign _zz_1467 = _zz_1468;
  assign _zz_1468 = ($signed(_zz_1469) >>> _zz_74);
  assign _zz_1469 = _zz_1470;
  assign _zz_1470 = ($signed(_zz_1472) - $signed(_zz_71));
  assign _zz_1471 = ({8'd0,data_mid_28_real} <<< 8);
  assign _zz_1472 = {{8{_zz_1471[23]}}, _zz_1471};
  assign _zz_1473 = fixTo_86_dout;
  assign _zz_1474 = _zz_1475[31 : 0];
  assign _zz_1475 = _zz_1476;
  assign _zz_1476 = ($signed(_zz_1477) >>> _zz_74);
  assign _zz_1477 = _zz_1478;
  assign _zz_1478 = ($signed(_zz_1480) - $signed(_zz_72));
  assign _zz_1479 = ({8'd0,data_mid_28_imag} <<< 8);
  assign _zz_1480 = {{8{_zz_1479[23]}}, _zz_1479};
  assign _zz_1481 = fixTo_87_dout;
  assign _zz_1482 = _zz_1483[31 : 0];
  assign _zz_1483 = _zz_1484;
  assign _zz_1484 = ($signed(_zz_1485) >>> _zz_75);
  assign _zz_1485 = _zz_1486;
  assign _zz_1486 = ($signed(_zz_1488) + $signed(_zz_71));
  assign _zz_1487 = ({8'd0,data_mid_28_real} <<< 8);
  assign _zz_1488 = {{8{_zz_1487[23]}}, _zz_1487};
  assign _zz_1489 = fixTo_88_dout;
  assign _zz_1490 = _zz_1491[31 : 0];
  assign _zz_1491 = _zz_1492;
  assign _zz_1492 = ($signed(_zz_1493) >>> _zz_75);
  assign _zz_1493 = _zz_1494;
  assign _zz_1494 = ($signed(_zz_1496) + $signed(_zz_72));
  assign _zz_1495 = ({8'd0,data_mid_28_imag} <<< 8);
  assign _zz_1496 = {{8{_zz_1495[23]}}, _zz_1495};
  assign _zz_1497 = fixTo_89_dout;
  assign _zz_1498 = ($signed(twiddle_factor_table_0_real) + $signed(twiddle_factor_table_0_imag));
  assign _zz_1499 = ($signed(_zz_78) - $signed(_zz_1500));
  assign _zz_1500 = ($signed(_zz_1501) * $signed(twiddle_factor_table_0_imag));
  assign _zz_1501 = ($signed(data_mid_31_real) + $signed(data_mid_31_imag));
  assign _zz_1502 = fixTo_90_dout;
  assign _zz_1503 = ($signed(_zz_78) + $signed(_zz_1504));
  assign _zz_1504 = ($signed(_zz_1505) * $signed(twiddle_factor_table_0_real));
  assign _zz_1505 = ($signed(data_mid_31_imag) - $signed(data_mid_31_real));
  assign _zz_1506 = fixTo_91_dout;
  assign _zz_1507 = _zz_1508[31 : 0];
  assign _zz_1508 = _zz_1509;
  assign _zz_1509 = ($signed(_zz_1510) >>> _zz_79);
  assign _zz_1510 = _zz_1511;
  assign _zz_1511 = ($signed(_zz_1513) - $signed(_zz_76));
  assign _zz_1512 = ({8'd0,data_mid_30_real} <<< 8);
  assign _zz_1513 = {{8{_zz_1512[23]}}, _zz_1512};
  assign _zz_1514 = fixTo_92_dout;
  assign _zz_1515 = _zz_1516[31 : 0];
  assign _zz_1516 = _zz_1517;
  assign _zz_1517 = ($signed(_zz_1518) >>> _zz_79);
  assign _zz_1518 = _zz_1519;
  assign _zz_1519 = ($signed(_zz_1521) - $signed(_zz_77));
  assign _zz_1520 = ({8'd0,data_mid_30_imag} <<< 8);
  assign _zz_1521 = {{8{_zz_1520[23]}}, _zz_1520};
  assign _zz_1522 = fixTo_93_dout;
  assign _zz_1523 = _zz_1524[31 : 0];
  assign _zz_1524 = _zz_1525;
  assign _zz_1525 = ($signed(_zz_1526) >>> _zz_80);
  assign _zz_1526 = _zz_1527;
  assign _zz_1527 = ($signed(_zz_1529) + $signed(_zz_76));
  assign _zz_1528 = ({8'd0,data_mid_30_real} <<< 8);
  assign _zz_1529 = {{8{_zz_1528[23]}}, _zz_1528};
  assign _zz_1530 = fixTo_94_dout;
  assign _zz_1531 = _zz_1532[31 : 0];
  assign _zz_1532 = _zz_1533;
  assign _zz_1533 = ($signed(_zz_1534) >>> _zz_80);
  assign _zz_1534 = _zz_1535;
  assign _zz_1535 = ($signed(_zz_1537) + $signed(_zz_77));
  assign _zz_1536 = ({8'd0,data_mid_30_imag} <<< 8);
  assign _zz_1537 = {{8{_zz_1536[23]}}, _zz_1536};
  assign _zz_1538 = fixTo_95_dout;
  assign _zz_1539 = ($signed(twiddle_factor_table_1_real) + $signed(twiddle_factor_table_1_imag));
  assign _zz_1540 = ($signed(_zz_83) - $signed(_zz_1541));
  assign _zz_1541 = ($signed(_zz_1542) * $signed(twiddle_factor_table_1_imag));
  assign _zz_1542 = ($signed(data_mid_2_real) + $signed(data_mid_2_imag));
  assign _zz_1543 = fixTo_96_dout;
  assign _zz_1544 = ($signed(_zz_83) + $signed(_zz_1545));
  assign _zz_1545 = ($signed(_zz_1546) * $signed(twiddle_factor_table_1_real));
  assign _zz_1546 = ($signed(data_mid_2_imag) - $signed(data_mid_2_real));
  assign _zz_1547 = fixTo_97_dout;
  assign _zz_1548 = _zz_1549[31 : 0];
  assign _zz_1549 = _zz_1550;
  assign _zz_1550 = ($signed(_zz_1551) >>> _zz_84);
  assign _zz_1551 = _zz_1552;
  assign _zz_1552 = ($signed(_zz_1554) - $signed(_zz_81));
  assign _zz_1553 = ({8'd0,data_mid_0_real} <<< 8);
  assign _zz_1554 = {{8{_zz_1553[23]}}, _zz_1553};
  assign _zz_1555 = fixTo_98_dout;
  assign _zz_1556 = _zz_1557[31 : 0];
  assign _zz_1557 = _zz_1558;
  assign _zz_1558 = ($signed(_zz_1559) >>> _zz_84);
  assign _zz_1559 = _zz_1560;
  assign _zz_1560 = ($signed(_zz_1562) - $signed(_zz_82));
  assign _zz_1561 = ({8'd0,data_mid_0_imag} <<< 8);
  assign _zz_1562 = {{8{_zz_1561[23]}}, _zz_1561};
  assign _zz_1563 = fixTo_99_dout;
  assign _zz_1564 = _zz_1565[31 : 0];
  assign _zz_1565 = _zz_1566;
  assign _zz_1566 = ($signed(_zz_1567) >>> _zz_85);
  assign _zz_1567 = _zz_1568;
  assign _zz_1568 = ($signed(_zz_1570) + $signed(_zz_81));
  assign _zz_1569 = ({8'd0,data_mid_0_real} <<< 8);
  assign _zz_1570 = {{8{_zz_1569[23]}}, _zz_1569};
  assign _zz_1571 = fixTo_100_dout;
  assign _zz_1572 = _zz_1573[31 : 0];
  assign _zz_1573 = _zz_1574;
  assign _zz_1574 = ($signed(_zz_1575) >>> _zz_85);
  assign _zz_1575 = _zz_1576;
  assign _zz_1576 = ($signed(_zz_1578) + $signed(_zz_82));
  assign _zz_1577 = ({8'd0,data_mid_0_imag} <<< 8);
  assign _zz_1578 = {{8{_zz_1577[23]}}, _zz_1577};
  assign _zz_1579 = fixTo_101_dout;
  assign _zz_1580 = ($signed(twiddle_factor_table_2_real) + $signed(twiddle_factor_table_2_imag));
  assign _zz_1581 = ($signed(_zz_88) - $signed(_zz_1582));
  assign _zz_1582 = ($signed(_zz_1583) * $signed(twiddle_factor_table_2_imag));
  assign _zz_1583 = ($signed(data_mid_3_real) + $signed(data_mid_3_imag));
  assign _zz_1584 = fixTo_102_dout;
  assign _zz_1585 = ($signed(_zz_88) + $signed(_zz_1586));
  assign _zz_1586 = ($signed(_zz_1587) * $signed(twiddle_factor_table_2_real));
  assign _zz_1587 = ($signed(data_mid_3_imag) - $signed(data_mid_3_real));
  assign _zz_1588 = fixTo_103_dout;
  assign _zz_1589 = _zz_1590[31 : 0];
  assign _zz_1590 = _zz_1591;
  assign _zz_1591 = ($signed(_zz_1592) >>> _zz_89);
  assign _zz_1592 = _zz_1593;
  assign _zz_1593 = ($signed(_zz_1595) - $signed(_zz_86));
  assign _zz_1594 = ({8'd0,data_mid_1_real} <<< 8);
  assign _zz_1595 = {{8{_zz_1594[23]}}, _zz_1594};
  assign _zz_1596 = fixTo_104_dout;
  assign _zz_1597 = _zz_1598[31 : 0];
  assign _zz_1598 = _zz_1599;
  assign _zz_1599 = ($signed(_zz_1600) >>> _zz_89);
  assign _zz_1600 = _zz_1601;
  assign _zz_1601 = ($signed(_zz_1603) - $signed(_zz_87));
  assign _zz_1602 = ({8'd0,data_mid_1_imag} <<< 8);
  assign _zz_1603 = {{8{_zz_1602[23]}}, _zz_1602};
  assign _zz_1604 = fixTo_105_dout;
  assign _zz_1605 = _zz_1606[31 : 0];
  assign _zz_1606 = _zz_1607;
  assign _zz_1607 = ($signed(_zz_1608) >>> _zz_90);
  assign _zz_1608 = _zz_1609;
  assign _zz_1609 = ($signed(_zz_1611) + $signed(_zz_86));
  assign _zz_1610 = ({8'd0,data_mid_1_real} <<< 8);
  assign _zz_1611 = {{8{_zz_1610[23]}}, _zz_1610};
  assign _zz_1612 = fixTo_106_dout;
  assign _zz_1613 = _zz_1614[31 : 0];
  assign _zz_1614 = _zz_1615;
  assign _zz_1615 = ($signed(_zz_1616) >>> _zz_90);
  assign _zz_1616 = _zz_1617;
  assign _zz_1617 = ($signed(_zz_1619) + $signed(_zz_87));
  assign _zz_1618 = ({8'd0,data_mid_1_imag} <<< 8);
  assign _zz_1619 = {{8{_zz_1618[23]}}, _zz_1618};
  assign _zz_1620 = fixTo_107_dout;
  assign _zz_1621 = ($signed(twiddle_factor_table_1_real) + $signed(twiddle_factor_table_1_imag));
  assign _zz_1622 = ($signed(_zz_93) - $signed(_zz_1623));
  assign _zz_1623 = ($signed(_zz_1624) * $signed(twiddle_factor_table_1_imag));
  assign _zz_1624 = ($signed(data_mid_6_real) + $signed(data_mid_6_imag));
  assign _zz_1625 = fixTo_108_dout;
  assign _zz_1626 = ($signed(_zz_93) + $signed(_zz_1627));
  assign _zz_1627 = ($signed(_zz_1628) * $signed(twiddle_factor_table_1_real));
  assign _zz_1628 = ($signed(data_mid_6_imag) - $signed(data_mid_6_real));
  assign _zz_1629 = fixTo_109_dout;
  assign _zz_1630 = _zz_1631[31 : 0];
  assign _zz_1631 = _zz_1632;
  assign _zz_1632 = ($signed(_zz_1633) >>> _zz_94);
  assign _zz_1633 = _zz_1634;
  assign _zz_1634 = ($signed(_zz_1636) - $signed(_zz_91));
  assign _zz_1635 = ({8'd0,data_mid_4_real} <<< 8);
  assign _zz_1636 = {{8{_zz_1635[23]}}, _zz_1635};
  assign _zz_1637 = fixTo_110_dout;
  assign _zz_1638 = _zz_1639[31 : 0];
  assign _zz_1639 = _zz_1640;
  assign _zz_1640 = ($signed(_zz_1641) >>> _zz_94);
  assign _zz_1641 = _zz_1642;
  assign _zz_1642 = ($signed(_zz_1644) - $signed(_zz_92));
  assign _zz_1643 = ({8'd0,data_mid_4_imag} <<< 8);
  assign _zz_1644 = {{8{_zz_1643[23]}}, _zz_1643};
  assign _zz_1645 = fixTo_111_dout;
  assign _zz_1646 = _zz_1647[31 : 0];
  assign _zz_1647 = _zz_1648;
  assign _zz_1648 = ($signed(_zz_1649) >>> _zz_95);
  assign _zz_1649 = _zz_1650;
  assign _zz_1650 = ($signed(_zz_1652) + $signed(_zz_91));
  assign _zz_1651 = ({8'd0,data_mid_4_real} <<< 8);
  assign _zz_1652 = {{8{_zz_1651[23]}}, _zz_1651};
  assign _zz_1653 = fixTo_112_dout;
  assign _zz_1654 = _zz_1655[31 : 0];
  assign _zz_1655 = _zz_1656;
  assign _zz_1656 = ($signed(_zz_1657) >>> _zz_95);
  assign _zz_1657 = _zz_1658;
  assign _zz_1658 = ($signed(_zz_1660) + $signed(_zz_92));
  assign _zz_1659 = ({8'd0,data_mid_4_imag} <<< 8);
  assign _zz_1660 = {{8{_zz_1659[23]}}, _zz_1659};
  assign _zz_1661 = fixTo_113_dout;
  assign _zz_1662 = ($signed(twiddle_factor_table_2_real) + $signed(twiddle_factor_table_2_imag));
  assign _zz_1663 = ($signed(_zz_98) - $signed(_zz_1664));
  assign _zz_1664 = ($signed(_zz_1665) * $signed(twiddle_factor_table_2_imag));
  assign _zz_1665 = ($signed(data_mid_7_real) + $signed(data_mid_7_imag));
  assign _zz_1666 = fixTo_114_dout;
  assign _zz_1667 = ($signed(_zz_98) + $signed(_zz_1668));
  assign _zz_1668 = ($signed(_zz_1669) * $signed(twiddle_factor_table_2_real));
  assign _zz_1669 = ($signed(data_mid_7_imag) - $signed(data_mid_7_real));
  assign _zz_1670 = fixTo_115_dout;
  assign _zz_1671 = _zz_1672[31 : 0];
  assign _zz_1672 = _zz_1673;
  assign _zz_1673 = ($signed(_zz_1674) >>> _zz_99);
  assign _zz_1674 = _zz_1675;
  assign _zz_1675 = ($signed(_zz_1677) - $signed(_zz_96));
  assign _zz_1676 = ({8'd0,data_mid_5_real} <<< 8);
  assign _zz_1677 = {{8{_zz_1676[23]}}, _zz_1676};
  assign _zz_1678 = fixTo_116_dout;
  assign _zz_1679 = _zz_1680[31 : 0];
  assign _zz_1680 = _zz_1681;
  assign _zz_1681 = ($signed(_zz_1682) >>> _zz_99);
  assign _zz_1682 = _zz_1683;
  assign _zz_1683 = ($signed(_zz_1685) - $signed(_zz_97));
  assign _zz_1684 = ({8'd0,data_mid_5_imag} <<< 8);
  assign _zz_1685 = {{8{_zz_1684[23]}}, _zz_1684};
  assign _zz_1686 = fixTo_117_dout;
  assign _zz_1687 = _zz_1688[31 : 0];
  assign _zz_1688 = _zz_1689;
  assign _zz_1689 = ($signed(_zz_1690) >>> _zz_100);
  assign _zz_1690 = _zz_1691;
  assign _zz_1691 = ($signed(_zz_1693) + $signed(_zz_96));
  assign _zz_1692 = ({8'd0,data_mid_5_real} <<< 8);
  assign _zz_1693 = {{8{_zz_1692[23]}}, _zz_1692};
  assign _zz_1694 = fixTo_118_dout;
  assign _zz_1695 = _zz_1696[31 : 0];
  assign _zz_1696 = _zz_1697;
  assign _zz_1697 = ($signed(_zz_1698) >>> _zz_100);
  assign _zz_1698 = _zz_1699;
  assign _zz_1699 = ($signed(_zz_1701) + $signed(_zz_97));
  assign _zz_1700 = ({8'd0,data_mid_5_imag} <<< 8);
  assign _zz_1701 = {{8{_zz_1700[23]}}, _zz_1700};
  assign _zz_1702 = fixTo_119_dout;
  assign _zz_1703 = ($signed(twiddle_factor_table_1_real) + $signed(twiddle_factor_table_1_imag));
  assign _zz_1704 = ($signed(_zz_103) - $signed(_zz_1705));
  assign _zz_1705 = ($signed(_zz_1706) * $signed(twiddle_factor_table_1_imag));
  assign _zz_1706 = ($signed(data_mid_10_real) + $signed(data_mid_10_imag));
  assign _zz_1707 = fixTo_120_dout;
  assign _zz_1708 = ($signed(_zz_103) + $signed(_zz_1709));
  assign _zz_1709 = ($signed(_zz_1710) * $signed(twiddle_factor_table_1_real));
  assign _zz_1710 = ($signed(data_mid_10_imag) - $signed(data_mid_10_real));
  assign _zz_1711 = fixTo_121_dout;
  assign _zz_1712 = _zz_1713[31 : 0];
  assign _zz_1713 = _zz_1714;
  assign _zz_1714 = ($signed(_zz_1715) >>> _zz_104);
  assign _zz_1715 = _zz_1716;
  assign _zz_1716 = ($signed(_zz_1718) - $signed(_zz_101));
  assign _zz_1717 = ({8'd0,data_mid_8_real} <<< 8);
  assign _zz_1718 = {{8{_zz_1717[23]}}, _zz_1717};
  assign _zz_1719 = fixTo_122_dout;
  assign _zz_1720 = _zz_1721[31 : 0];
  assign _zz_1721 = _zz_1722;
  assign _zz_1722 = ($signed(_zz_1723) >>> _zz_104);
  assign _zz_1723 = _zz_1724;
  assign _zz_1724 = ($signed(_zz_1726) - $signed(_zz_102));
  assign _zz_1725 = ({8'd0,data_mid_8_imag} <<< 8);
  assign _zz_1726 = {{8{_zz_1725[23]}}, _zz_1725};
  assign _zz_1727 = fixTo_123_dout;
  assign _zz_1728 = _zz_1729[31 : 0];
  assign _zz_1729 = _zz_1730;
  assign _zz_1730 = ($signed(_zz_1731) >>> _zz_105);
  assign _zz_1731 = _zz_1732;
  assign _zz_1732 = ($signed(_zz_1734) + $signed(_zz_101));
  assign _zz_1733 = ({8'd0,data_mid_8_real} <<< 8);
  assign _zz_1734 = {{8{_zz_1733[23]}}, _zz_1733};
  assign _zz_1735 = fixTo_124_dout;
  assign _zz_1736 = _zz_1737[31 : 0];
  assign _zz_1737 = _zz_1738;
  assign _zz_1738 = ($signed(_zz_1739) >>> _zz_105);
  assign _zz_1739 = _zz_1740;
  assign _zz_1740 = ($signed(_zz_1742) + $signed(_zz_102));
  assign _zz_1741 = ({8'd0,data_mid_8_imag} <<< 8);
  assign _zz_1742 = {{8{_zz_1741[23]}}, _zz_1741};
  assign _zz_1743 = fixTo_125_dout;
  assign _zz_1744 = ($signed(twiddle_factor_table_2_real) + $signed(twiddle_factor_table_2_imag));
  assign _zz_1745 = ($signed(_zz_108) - $signed(_zz_1746));
  assign _zz_1746 = ($signed(_zz_1747) * $signed(twiddle_factor_table_2_imag));
  assign _zz_1747 = ($signed(data_mid_11_real) + $signed(data_mid_11_imag));
  assign _zz_1748 = fixTo_126_dout;
  assign _zz_1749 = ($signed(_zz_108) + $signed(_zz_1750));
  assign _zz_1750 = ($signed(_zz_1751) * $signed(twiddle_factor_table_2_real));
  assign _zz_1751 = ($signed(data_mid_11_imag) - $signed(data_mid_11_real));
  assign _zz_1752 = fixTo_127_dout;
  assign _zz_1753 = _zz_1754[31 : 0];
  assign _zz_1754 = _zz_1755;
  assign _zz_1755 = ($signed(_zz_1756) >>> _zz_109);
  assign _zz_1756 = _zz_1757;
  assign _zz_1757 = ($signed(_zz_1759) - $signed(_zz_106));
  assign _zz_1758 = ({8'd0,data_mid_9_real} <<< 8);
  assign _zz_1759 = {{8{_zz_1758[23]}}, _zz_1758};
  assign _zz_1760 = fixTo_128_dout;
  assign _zz_1761 = _zz_1762[31 : 0];
  assign _zz_1762 = _zz_1763;
  assign _zz_1763 = ($signed(_zz_1764) >>> _zz_109);
  assign _zz_1764 = _zz_1765;
  assign _zz_1765 = ($signed(_zz_1767) - $signed(_zz_107));
  assign _zz_1766 = ({8'd0,data_mid_9_imag} <<< 8);
  assign _zz_1767 = {{8{_zz_1766[23]}}, _zz_1766};
  assign _zz_1768 = fixTo_129_dout;
  assign _zz_1769 = _zz_1770[31 : 0];
  assign _zz_1770 = _zz_1771;
  assign _zz_1771 = ($signed(_zz_1772) >>> _zz_110);
  assign _zz_1772 = _zz_1773;
  assign _zz_1773 = ($signed(_zz_1775) + $signed(_zz_106));
  assign _zz_1774 = ({8'd0,data_mid_9_real} <<< 8);
  assign _zz_1775 = {{8{_zz_1774[23]}}, _zz_1774};
  assign _zz_1776 = fixTo_130_dout;
  assign _zz_1777 = _zz_1778[31 : 0];
  assign _zz_1778 = _zz_1779;
  assign _zz_1779 = ($signed(_zz_1780) >>> _zz_110);
  assign _zz_1780 = _zz_1781;
  assign _zz_1781 = ($signed(_zz_1783) + $signed(_zz_107));
  assign _zz_1782 = ({8'd0,data_mid_9_imag} <<< 8);
  assign _zz_1783 = {{8{_zz_1782[23]}}, _zz_1782};
  assign _zz_1784 = fixTo_131_dout;
  assign _zz_1785 = ($signed(twiddle_factor_table_1_real) + $signed(twiddle_factor_table_1_imag));
  assign _zz_1786 = ($signed(_zz_113) - $signed(_zz_1787));
  assign _zz_1787 = ($signed(_zz_1788) * $signed(twiddle_factor_table_1_imag));
  assign _zz_1788 = ($signed(data_mid_14_real) + $signed(data_mid_14_imag));
  assign _zz_1789 = fixTo_132_dout;
  assign _zz_1790 = ($signed(_zz_113) + $signed(_zz_1791));
  assign _zz_1791 = ($signed(_zz_1792) * $signed(twiddle_factor_table_1_real));
  assign _zz_1792 = ($signed(data_mid_14_imag) - $signed(data_mid_14_real));
  assign _zz_1793 = fixTo_133_dout;
  assign _zz_1794 = _zz_1795[31 : 0];
  assign _zz_1795 = _zz_1796;
  assign _zz_1796 = ($signed(_zz_1797) >>> _zz_114);
  assign _zz_1797 = _zz_1798;
  assign _zz_1798 = ($signed(_zz_1800) - $signed(_zz_111));
  assign _zz_1799 = ({8'd0,data_mid_12_real} <<< 8);
  assign _zz_1800 = {{8{_zz_1799[23]}}, _zz_1799};
  assign _zz_1801 = fixTo_134_dout;
  assign _zz_1802 = _zz_1803[31 : 0];
  assign _zz_1803 = _zz_1804;
  assign _zz_1804 = ($signed(_zz_1805) >>> _zz_114);
  assign _zz_1805 = _zz_1806;
  assign _zz_1806 = ($signed(_zz_1808) - $signed(_zz_112));
  assign _zz_1807 = ({8'd0,data_mid_12_imag} <<< 8);
  assign _zz_1808 = {{8{_zz_1807[23]}}, _zz_1807};
  assign _zz_1809 = fixTo_135_dout;
  assign _zz_1810 = _zz_1811[31 : 0];
  assign _zz_1811 = _zz_1812;
  assign _zz_1812 = ($signed(_zz_1813) >>> _zz_115);
  assign _zz_1813 = _zz_1814;
  assign _zz_1814 = ($signed(_zz_1816) + $signed(_zz_111));
  assign _zz_1815 = ({8'd0,data_mid_12_real} <<< 8);
  assign _zz_1816 = {{8{_zz_1815[23]}}, _zz_1815};
  assign _zz_1817 = fixTo_136_dout;
  assign _zz_1818 = _zz_1819[31 : 0];
  assign _zz_1819 = _zz_1820;
  assign _zz_1820 = ($signed(_zz_1821) >>> _zz_115);
  assign _zz_1821 = _zz_1822;
  assign _zz_1822 = ($signed(_zz_1824) + $signed(_zz_112));
  assign _zz_1823 = ({8'd0,data_mid_12_imag} <<< 8);
  assign _zz_1824 = {{8{_zz_1823[23]}}, _zz_1823};
  assign _zz_1825 = fixTo_137_dout;
  assign _zz_1826 = ($signed(twiddle_factor_table_2_real) + $signed(twiddle_factor_table_2_imag));
  assign _zz_1827 = ($signed(_zz_118) - $signed(_zz_1828));
  assign _zz_1828 = ($signed(_zz_1829) * $signed(twiddle_factor_table_2_imag));
  assign _zz_1829 = ($signed(data_mid_15_real) + $signed(data_mid_15_imag));
  assign _zz_1830 = fixTo_138_dout;
  assign _zz_1831 = ($signed(_zz_118) + $signed(_zz_1832));
  assign _zz_1832 = ($signed(_zz_1833) * $signed(twiddle_factor_table_2_real));
  assign _zz_1833 = ($signed(data_mid_15_imag) - $signed(data_mid_15_real));
  assign _zz_1834 = fixTo_139_dout;
  assign _zz_1835 = _zz_1836[31 : 0];
  assign _zz_1836 = _zz_1837;
  assign _zz_1837 = ($signed(_zz_1838) >>> _zz_119);
  assign _zz_1838 = _zz_1839;
  assign _zz_1839 = ($signed(_zz_1841) - $signed(_zz_116));
  assign _zz_1840 = ({8'd0,data_mid_13_real} <<< 8);
  assign _zz_1841 = {{8{_zz_1840[23]}}, _zz_1840};
  assign _zz_1842 = fixTo_140_dout;
  assign _zz_1843 = _zz_1844[31 : 0];
  assign _zz_1844 = _zz_1845;
  assign _zz_1845 = ($signed(_zz_1846) >>> _zz_119);
  assign _zz_1846 = _zz_1847;
  assign _zz_1847 = ($signed(_zz_1849) - $signed(_zz_117));
  assign _zz_1848 = ({8'd0,data_mid_13_imag} <<< 8);
  assign _zz_1849 = {{8{_zz_1848[23]}}, _zz_1848};
  assign _zz_1850 = fixTo_141_dout;
  assign _zz_1851 = _zz_1852[31 : 0];
  assign _zz_1852 = _zz_1853;
  assign _zz_1853 = ($signed(_zz_1854) >>> _zz_120);
  assign _zz_1854 = _zz_1855;
  assign _zz_1855 = ($signed(_zz_1857) + $signed(_zz_116));
  assign _zz_1856 = ({8'd0,data_mid_13_real} <<< 8);
  assign _zz_1857 = {{8{_zz_1856[23]}}, _zz_1856};
  assign _zz_1858 = fixTo_142_dout;
  assign _zz_1859 = _zz_1860[31 : 0];
  assign _zz_1860 = _zz_1861;
  assign _zz_1861 = ($signed(_zz_1862) >>> _zz_120);
  assign _zz_1862 = _zz_1863;
  assign _zz_1863 = ($signed(_zz_1865) + $signed(_zz_117));
  assign _zz_1864 = ({8'd0,data_mid_13_imag} <<< 8);
  assign _zz_1865 = {{8{_zz_1864[23]}}, _zz_1864};
  assign _zz_1866 = fixTo_143_dout;
  assign _zz_1867 = ($signed(twiddle_factor_table_1_real) + $signed(twiddle_factor_table_1_imag));
  assign _zz_1868 = ($signed(_zz_123) - $signed(_zz_1869));
  assign _zz_1869 = ($signed(_zz_1870) * $signed(twiddle_factor_table_1_imag));
  assign _zz_1870 = ($signed(data_mid_18_real) + $signed(data_mid_18_imag));
  assign _zz_1871 = fixTo_144_dout;
  assign _zz_1872 = ($signed(_zz_123) + $signed(_zz_1873));
  assign _zz_1873 = ($signed(_zz_1874) * $signed(twiddle_factor_table_1_real));
  assign _zz_1874 = ($signed(data_mid_18_imag) - $signed(data_mid_18_real));
  assign _zz_1875 = fixTo_145_dout;
  assign _zz_1876 = _zz_1877[31 : 0];
  assign _zz_1877 = _zz_1878;
  assign _zz_1878 = ($signed(_zz_1879) >>> _zz_124);
  assign _zz_1879 = _zz_1880;
  assign _zz_1880 = ($signed(_zz_1882) - $signed(_zz_121));
  assign _zz_1881 = ({8'd0,data_mid_16_real} <<< 8);
  assign _zz_1882 = {{8{_zz_1881[23]}}, _zz_1881};
  assign _zz_1883 = fixTo_146_dout;
  assign _zz_1884 = _zz_1885[31 : 0];
  assign _zz_1885 = _zz_1886;
  assign _zz_1886 = ($signed(_zz_1887) >>> _zz_124);
  assign _zz_1887 = _zz_1888;
  assign _zz_1888 = ($signed(_zz_1890) - $signed(_zz_122));
  assign _zz_1889 = ({8'd0,data_mid_16_imag} <<< 8);
  assign _zz_1890 = {{8{_zz_1889[23]}}, _zz_1889};
  assign _zz_1891 = fixTo_147_dout;
  assign _zz_1892 = _zz_1893[31 : 0];
  assign _zz_1893 = _zz_1894;
  assign _zz_1894 = ($signed(_zz_1895) >>> _zz_125);
  assign _zz_1895 = _zz_1896;
  assign _zz_1896 = ($signed(_zz_1898) + $signed(_zz_121));
  assign _zz_1897 = ({8'd0,data_mid_16_real} <<< 8);
  assign _zz_1898 = {{8{_zz_1897[23]}}, _zz_1897};
  assign _zz_1899 = fixTo_148_dout;
  assign _zz_1900 = _zz_1901[31 : 0];
  assign _zz_1901 = _zz_1902;
  assign _zz_1902 = ($signed(_zz_1903) >>> _zz_125);
  assign _zz_1903 = _zz_1904;
  assign _zz_1904 = ($signed(_zz_1906) + $signed(_zz_122));
  assign _zz_1905 = ({8'd0,data_mid_16_imag} <<< 8);
  assign _zz_1906 = {{8{_zz_1905[23]}}, _zz_1905};
  assign _zz_1907 = fixTo_149_dout;
  assign _zz_1908 = ($signed(twiddle_factor_table_2_real) + $signed(twiddle_factor_table_2_imag));
  assign _zz_1909 = ($signed(_zz_128) - $signed(_zz_1910));
  assign _zz_1910 = ($signed(_zz_1911) * $signed(twiddle_factor_table_2_imag));
  assign _zz_1911 = ($signed(data_mid_19_real) + $signed(data_mid_19_imag));
  assign _zz_1912 = fixTo_150_dout;
  assign _zz_1913 = ($signed(_zz_128) + $signed(_zz_1914));
  assign _zz_1914 = ($signed(_zz_1915) * $signed(twiddle_factor_table_2_real));
  assign _zz_1915 = ($signed(data_mid_19_imag) - $signed(data_mid_19_real));
  assign _zz_1916 = fixTo_151_dout;
  assign _zz_1917 = _zz_1918[31 : 0];
  assign _zz_1918 = _zz_1919;
  assign _zz_1919 = ($signed(_zz_1920) >>> _zz_129);
  assign _zz_1920 = _zz_1921;
  assign _zz_1921 = ($signed(_zz_1923) - $signed(_zz_126));
  assign _zz_1922 = ({8'd0,data_mid_17_real} <<< 8);
  assign _zz_1923 = {{8{_zz_1922[23]}}, _zz_1922};
  assign _zz_1924 = fixTo_152_dout;
  assign _zz_1925 = _zz_1926[31 : 0];
  assign _zz_1926 = _zz_1927;
  assign _zz_1927 = ($signed(_zz_1928) >>> _zz_129);
  assign _zz_1928 = _zz_1929;
  assign _zz_1929 = ($signed(_zz_1931) - $signed(_zz_127));
  assign _zz_1930 = ({8'd0,data_mid_17_imag} <<< 8);
  assign _zz_1931 = {{8{_zz_1930[23]}}, _zz_1930};
  assign _zz_1932 = fixTo_153_dout;
  assign _zz_1933 = _zz_1934[31 : 0];
  assign _zz_1934 = _zz_1935;
  assign _zz_1935 = ($signed(_zz_1936) >>> _zz_130);
  assign _zz_1936 = _zz_1937;
  assign _zz_1937 = ($signed(_zz_1939) + $signed(_zz_126));
  assign _zz_1938 = ({8'd0,data_mid_17_real} <<< 8);
  assign _zz_1939 = {{8{_zz_1938[23]}}, _zz_1938};
  assign _zz_1940 = fixTo_154_dout;
  assign _zz_1941 = _zz_1942[31 : 0];
  assign _zz_1942 = _zz_1943;
  assign _zz_1943 = ($signed(_zz_1944) >>> _zz_130);
  assign _zz_1944 = _zz_1945;
  assign _zz_1945 = ($signed(_zz_1947) + $signed(_zz_127));
  assign _zz_1946 = ({8'd0,data_mid_17_imag} <<< 8);
  assign _zz_1947 = {{8{_zz_1946[23]}}, _zz_1946};
  assign _zz_1948 = fixTo_155_dout;
  assign _zz_1949 = ($signed(twiddle_factor_table_1_real) + $signed(twiddle_factor_table_1_imag));
  assign _zz_1950 = ($signed(_zz_133) - $signed(_zz_1951));
  assign _zz_1951 = ($signed(_zz_1952) * $signed(twiddle_factor_table_1_imag));
  assign _zz_1952 = ($signed(data_mid_22_real) + $signed(data_mid_22_imag));
  assign _zz_1953 = fixTo_156_dout;
  assign _zz_1954 = ($signed(_zz_133) + $signed(_zz_1955));
  assign _zz_1955 = ($signed(_zz_1956) * $signed(twiddle_factor_table_1_real));
  assign _zz_1956 = ($signed(data_mid_22_imag) - $signed(data_mid_22_real));
  assign _zz_1957 = fixTo_157_dout;
  assign _zz_1958 = _zz_1959[31 : 0];
  assign _zz_1959 = _zz_1960;
  assign _zz_1960 = ($signed(_zz_1961) >>> _zz_134);
  assign _zz_1961 = _zz_1962;
  assign _zz_1962 = ($signed(_zz_1964) - $signed(_zz_131));
  assign _zz_1963 = ({8'd0,data_mid_20_real} <<< 8);
  assign _zz_1964 = {{8{_zz_1963[23]}}, _zz_1963};
  assign _zz_1965 = fixTo_158_dout;
  assign _zz_1966 = _zz_1967[31 : 0];
  assign _zz_1967 = _zz_1968;
  assign _zz_1968 = ($signed(_zz_1969) >>> _zz_134);
  assign _zz_1969 = _zz_1970;
  assign _zz_1970 = ($signed(_zz_1972) - $signed(_zz_132));
  assign _zz_1971 = ({8'd0,data_mid_20_imag} <<< 8);
  assign _zz_1972 = {{8{_zz_1971[23]}}, _zz_1971};
  assign _zz_1973 = fixTo_159_dout;
  assign _zz_1974 = _zz_1975[31 : 0];
  assign _zz_1975 = _zz_1976;
  assign _zz_1976 = ($signed(_zz_1977) >>> _zz_135);
  assign _zz_1977 = _zz_1978;
  assign _zz_1978 = ($signed(_zz_1980) + $signed(_zz_131));
  assign _zz_1979 = ({8'd0,data_mid_20_real} <<< 8);
  assign _zz_1980 = {{8{_zz_1979[23]}}, _zz_1979};
  assign _zz_1981 = fixTo_160_dout;
  assign _zz_1982 = _zz_1983[31 : 0];
  assign _zz_1983 = _zz_1984;
  assign _zz_1984 = ($signed(_zz_1985) >>> _zz_135);
  assign _zz_1985 = _zz_1986;
  assign _zz_1986 = ($signed(_zz_1988) + $signed(_zz_132));
  assign _zz_1987 = ({8'd0,data_mid_20_imag} <<< 8);
  assign _zz_1988 = {{8{_zz_1987[23]}}, _zz_1987};
  assign _zz_1989 = fixTo_161_dout;
  assign _zz_1990 = ($signed(twiddle_factor_table_2_real) + $signed(twiddle_factor_table_2_imag));
  assign _zz_1991 = ($signed(_zz_138) - $signed(_zz_1992));
  assign _zz_1992 = ($signed(_zz_1993) * $signed(twiddle_factor_table_2_imag));
  assign _zz_1993 = ($signed(data_mid_23_real) + $signed(data_mid_23_imag));
  assign _zz_1994 = fixTo_162_dout;
  assign _zz_1995 = ($signed(_zz_138) + $signed(_zz_1996));
  assign _zz_1996 = ($signed(_zz_1997) * $signed(twiddle_factor_table_2_real));
  assign _zz_1997 = ($signed(data_mid_23_imag) - $signed(data_mid_23_real));
  assign _zz_1998 = fixTo_163_dout;
  assign _zz_1999 = _zz_2000[31 : 0];
  assign _zz_2000 = _zz_2001;
  assign _zz_2001 = ($signed(_zz_2002) >>> _zz_139);
  assign _zz_2002 = _zz_2003;
  assign _zz_2003 = ($signed(_zz_2005) - $signed(_zz_136));
  assign _zz_2004 = ({8'd0,data_mid_21_real} <<< 8);
  assign _zz_2005 = {{8{_zz_2004[23]}}, _zz_2004};
  assign _zz_2006 = fixTo_164_dout;
  assign _zz_2007 = _zz_2008[31 : 0];
  assign _zz_2008 = _zz_2009;
  assign _zz_2009 = ($signed(_zz_2010) >>> _zz_139);
  assign _zz_2010 = _zz_2011;
  assign _zz_2011 = ($signed(_zz_2013) - $signed(_zz_137));
  assign _zz_2012 = ({8'd0,data_mid_21_imag} <<< 8);
  assign _zz_2013 = {{8{_zz_2012[23]}}, _zz_2012};
  assign _zz_2014 = fixTo_165_dout;
  assign _zz_2015 = _zz_2016[31 : 0];
  assign _zz_2016 = _zz_2017;
  assign _zz_2017 = ($signed(_zz_2018) >>> _zz_140);
  assign _zz_2018 = _zz_2019;
  assign _zz_2019 = ($signed(_zz_2021) + $signed(_zz_136));
  assign _zz_2020 = ({8'd0,data_mid_21_real} <<< 8);
  assign _zz_2021 = {{8{_zz_2020[23]}}, _zz_2020};
  assign _zz_2022 = fixTo_166_dout;
  assign _zz_2023 = _zz_2024[31 : 0];
  assign _zz_2024 = _zz_2025;
  assign _zz_2025 = ($signed(_zz_2026) >>> _zz_140);
  assign _zz_2026 = _zz_2027;
  assign _zz_2027 = ($signed(_zz_2029) + $signed(_zz_137));
  assign _zz_2028 = ({8'd0,data_mid_21_imag} <<< 8);
  assign _zz_2029 = {{8{_zz_2028[23]}}, _zz_2028};
  assign _zz_2030 = fixTo_167_dout;
  assign _zz_2031 = ($signed(twiddle_factor_table_1_real) + $signed(twiddle_factor_table_1_imag));
  assign _zz_2032 = ($signed(_zz_143) - $signed(_zz_2033));
  assign _zz_2033 = ($signed(_zz_2034) * $signed(twiddle_factor_table_1_imag));
  assign _zz_2034 = ($signed(data_mid_26_real) + $signed(data_mid_26_imag));
  assign _zz_2035 = fixTo_168_dout;
  assign _zz_2036 = ($signed(_zz_143) + $signed(_zz_2037));
  assign _zz_2037 = ($signed(_zz_2038) * $signed(twiddle_factor_table_1_real));
  assign _zz_2038 = ($signed(data_mid_26_imag) - $signed(data_mid_26_real));
  assign _zz_2039 = fixTo_169_dout;
  assign _zz_2040 = _zz_2041[31 : 0];
  assign _zz_2041 = _zz_2042;
  assign _zz_2042 = ($signed(_zz_2043) >>> _zz_144);
  assign _zz_2043 = _zz_2044;
  assign _zz_2044 = ($signed(_zz_2046) - $signed(_zz_141));
  assign _zz_2045 = ({8'd0,data_mid_24_real} <<< 8);
  assign _zz_2046 = {{8{_zz_2045[23]}}, _zz_2045};
  assign _zz_2047 = fixTo_170_dout;
  assign _zz_2048 = _zz_2049[31 : 0];
  assign _zz_2049 = _zz_2050;
  assign _zz_2050 = ($signed(_zz_2051) >>> _zz_144);
  assign _zz_2051 = _zz_2052;
  assign _zz_2052 = ($signed(_zz_2054) - $signed(_zz_142));
  assign _zz_2053 = ({8'd0,data_mid_24_imag} <<< 8);
  assign _zz_2054 = {{8{_zz_2053[23]}}, _zz_2053};
  assign _zz_2055 = fixTo_171_dout;
  assign _zz_2056 = _zz_2057[31 : 0];
  assign _zz_2057 = _zz_2058;
  assign _zz_2058 = ($signed(_zz_2059) >>> _zz_145);
  assign _zz_2059 = _zz_2060;
  assign _zz_2060 = ($signed(_zz_2062) + $signed(_zz_141));
  assign _zz_2061 = ({8'd0,data_mid_24_real} <<< 8);
  assign _zz_2062 = {{8{_zz_2061[23]}}, _zz_2061};
  assign _zz_2063 = fixTo_172_dout;
  assign _zz_2064 = _zz_2065[31 : 0];
  assign _zz_2065 = _zz_2066;
  assign _zz_2066 = ($signed(_zz_2067) >>> _zz_145);
  assign _zz_2067 = _zz_2068;
  assign _zz_2068 = ($signed(_zz_2070) + $signed(_zz_142));
  assign _zz_2069 = ({8'd0,data_mid_24_imag} <<< 8);
  assign _zz_2070 = {{8{_zz_2069[23]}}, _zz_2069};
  assign _zz_2071 = fixTo_173_dout;
  assign _zz_2072 = ($signed(twiddle_factor_table_2_real) + $signed(twiddle_factor_table_2_imag));
  assign _zz_2073 = ($signed(_zz_148) - $signed(_zz_2074));
  assign _zz_2074 = ($signed(_zz_2075) * $signed(twiddle_factor_table_2_imag));
  assign _zz_2075 = ($signed(data_mid_27_real) + $signed(data_mid_27_imag));
  assign _zz_2076 = fixTo_174_dout;
  assign _zz_2077 = ($signed(_zz_148) + $signed(_zz_2078));
  assign _zz_2078 = ($signed(_zz_2079) * $signed(twiddle_factor_table_2_real));
  assign _zz_2079 = ($signed(data_mid_27_imag) - $signed(data_mid_27_real));
  assign _zz_2080 = fixTo_175_dout;
  assign _zz_2081 = _zz_2082[31 : 0];
  assign _zz_2082 = _zz_2083;
  assign _zz_2083 = ($signed(_zz_2084) >>> _zz_149);
  assign _zz_2084 = _zz_2085;
  assign _zz_2085 = ($signed(_zz_2087) - $signed(_zz_146));
  assign _zz_2086 = ({8'd0,data_mid_25_real} <<< 8);
  assign _zz_2087 = {{8{_zz_2086[23]}}, _zz_2086};
  assign _zz_2088 = fixTo_176_dout;
  assign _zz_2089 = _zz_2090[31 : 0];
  assign _zz_2090 = _zz_2091;
  assign _zz_2091 = ($signed(_zz_2092) >>> _zz_149);
  assign _zz_2092 = _zz_2093;
  assign _zz_2093 = ($signed(_zz_2095) - $signed(_zz_147));
  assign _zz_2094 = ({8'd0,data_mid_25_imag} <<< 8);
  assign _zz_2095 = {{8{_zz_2094[23]}}, _zz_2094};
  assign _zz_2096 = fixTo_177_dout;
  assign _zz_2097 = _zz_2098[31 : 0];
  assign _zz_2098 = _zz_2099;
  assign _zz_2099 = ($signed(_zz_2100) >>> _zz_150);
  assign _zz_2100 = _zz_2101;
  assign _zz_2101 = ($signed(_zz_2103) + $signed(_zz_146));
  assign _zz_2102 = ({8'd0,data_mid_25_real} <<< 8);
  assign _zz_2103 = {{8{_zz_2102[23]}}, _zz_2102};
  assign _zz_2104 = fixTo_178_dout;
  assign _zz_2105 = _zz_2106[31 : 0];
  assign _zz_2106 = _zz_2107;
  assign _zz_2107 = ($signed(_zz_2108) >>> _zz_150);
  assign _zz_2108 = _zz_2109;
  assign _zz_2109 = ($signed(_zz_2111) + $signed(_zz_147));
  assign _zz_2110 = ({8'd0,data_mid_25_imag} <<< 8);
  assign _zz_2111 = {{8{_zz_2110[23]}}, _zz_2110};
  assign _zz_2112 = fixTo_179_dout;
  assign _zz_2113 = ($signed(twiddle_factor_table_1_real) + $signed(twiddle_factor_table_1_imag));
  assign _zz_2114 = ($signed(_zz_153) - $signed(_zz_2115));
  assign _zz_2115 = ($signed(_zz_2116) * $signed(twiddle_factor_table_1_imag));
  assign _zz_2116 = ($signed(data_mid_30_real) + $signed(data_mid_30_imag));
  assign _zz_2117 = fixTo_180_dout;
  assign _zz_2118 = ($signed(_zz_153) + $signed(_zz_2119));
  assign _zz_2119 = ($signed(_zz_2120) * $signed(twiddle_factor_table_1_real));
  assign _zz_2120 = ($signed(data_mid_30_imag) - $signed(data_mid_30_real));
  assign _zz_2121 = fixTo_181_dout;
  assign _zz_2122 = _zz_2123[31 : 0];
  assign _zz_2123 = _zz_2124;
  assign _zz_2124 = ($signed(_zz_2125) >>> _zz_154);
  assign _zz_2125 = _zz_2126;
  assign _zz_2126 = ($signed(_zz_2128) - $signed(_zz_151));
  assign _zz_2127 = ({8'd0,data_mid_28_real} <<< 8);
  assign _zz_2128 = {{8{_zz_2127[23]}}, _zz_2127};
  assign _zz_2129 = fixTo_182_dout;
  assign _zz_2130 = _zz_2131[31 : 0];
  assign _zz_2131 = _zz_2132;
  assign _zz_2132 = ($signed(_zz_2133) >>> _zz_154);
  assign _zz_2133 = _zz_2134;
  assign _zz_2134 = ($signed(_zz_2136) - $signed(_zz_152));
  assign _zz_2135 = ({8'd0,data_mid_28_imag} <<< 8);
  assign _zz_2136 = {{8{_zz_2135[23]}}, _zz_2135};
  assign _zz_2137 = fixTo_183_dout;
  assign _zz_2138 = _zz_2139[31 : 0];
  assign _zz_2139 = _zz_2140;
  assign _zz_2140 = ($signed(_zz_2141) >>> _zz_155);
  assign _zz_2141 = _zz_2142;
  assign _zz_2142 = ($signed(_zz_2144) + $signed(_zz_151));
  assign _zz_2143 = ({8'd0,data_mid_28_real} <<< 8);
  assign _zz_2144 = {{8{_zz_2143[23]}}, _zz_2143};
  assign _zz_2145 = fixTo_184_dout;
  assign _zz_2146 = _zz_2147[31 : 0];
  assign _zz_2147 = _zz_2148;
  assign _zz_2148 = ($signed(_zz_2149) >>> _zz_155);
  assign _zz_2149 = _zz_2150;
  assign _zz_2150 = ($signed(_zz_2152) + $signed(_zz_152));
  assign _zz_2151 = ({8'd0,data_mid_28_imag} <<< 8);
  assign _zz_2152 = {{8{_zz_2151[23]}}, _zz_2151};
  assign _zz_2153 = fixTo_185_dout;
  assign _zz_2154 = ($signed(twiddle_factor_table_2_real) + $signed(twiddle_factor_table_2_imag));
  assign _zz_2155 = ($signed(_zz_158) - $signed(_zz_2156));
  assign _zz_2156 = ($signed(_zz_2157) * $signed(twiddle_factor_table_2_imag));
  assign _zz_2157 = ($signed(data_mid_31_real) + $signed(data_mid_31_imag));
  assign _zz_2158 = fixTo_186_dout;
  assign _zz_2159 = ($signed(_zz_158) + $signed(_zz_2160));
  assign _zz_2160 = ($signed(_zz_2161) * $signed(twiddle_factor_table_2_real));
  assign _zz_2161 = ($signed(data_mid_31_imag) - $signed(data_mid_31_real));
  assign _zz_2162 = fixTo_187_dout;
  assign _zz_2163 = _zz_2164[31 : 0];
  assign _zz_2164 = _zz_2165;
  assign _zz_2165 = ($signed(_zz_2166) >>> _zz_159);
  assign _zz_2166 = _zz_2167;
  assign _zz_2167 = ($signed(_zz_2169) - $signed(_zz_156));
  assign _zz_2168 = ({8'd0,data_mid_29_real} <<< 8);
  assign _zz_2169 = {{8{_zz_2168[23]}}, _zz_2168};
  assign _zz_2170 = fixTo_188_dout;
  assign _zz_2171 = _zz_2172[31 : 0];
  assign _zz_2172 = _zz_2173;
  assign _zz_2173 = ($signed(_zz_2174) >>> _zz_159);
  assign _zz_2174 = _zz_2175;
  assign _zz_2175 = ($signed(_zz_2177) - $signed(_zz_157));
  assign _zz_2176 = ({8'd0,data_mid_29_imag} <<< 8);
  assign _zz_2177 = {{8{_zz_2176[23]}}, _zz_2176};
  assign _zz_2178 = fixTo_189_dout;
  assign _zz_2179 = _zz_2180[31 : 0];
  assign _zz_2180 = _zz_2181;
  assign _zz_2181 = ($signed(_zz_2182) >>> _zz_160);
  assign _zz_2182 = _zz_2183;
  assign _zz_2183 = ($signed(_zz_2185) + $signed(_zz_156));
  assign _zz_2184 = ({8'd0,data_mid_29_real} <<< 8);
  assign _zz_2185 = {{8{_zz_2184[23]}}, _zz_2184};
  assign _zz_2186 = fixTo_190_dout;
  assign _zz_2187 = _zz_2188[31 : 0];
  assign _zz_2188 = _zz_2189;
  assign _zz_2189 = ($signed(_zz_2190) >>> _zz_160);
  assign _zz_2190 = _zz_2191;
  assign _zz_2191 = ($signed(_zz_2193) + $signed(_zz_157));
  assign _zz_2192 = ({8'd0,data_mid_29_imag} <<< 8);
  assign _zz_2193 = {{8{_zz_2192[23]}}, _zz_2192};
  assign _zz_2194 = fixTo_191_dout;
  assign _zz_2195 = ($signed(twiddle_factor_table_3_real) + $signed(twiddle_factor_table_3_imag));
  assign _zz_2196 = ($signed(_zz_163) - $signed(_zz_2197));
  assign _zz_2197 = ($signed(_zz_2198) * $signed(twiddle_factor_table_3_imag));
  assign _zz_2198 = ($signed(data_mid_4_real) + $signed(data_mid_4_imag));
  assign _zz_2199 = fixTo_192_dout;
  assign _zz_2200 = ($signed(_zz_163) + $signed(_zz_2201));
  assign _zz_2201 = ($signed(_zz_2202) * $signed(twiddle_factor_table_3_real));
  assign _zz_2202 = ($signed(data_mid_4_imag) - $signed(data_mid_4_real));
  assign _zz_2203 = fixTo_193_dout;
  assign _zz_2204 = _zz_2205[31 : 0];
  assign _zz_2205 = _zz_2206;
  assign _zz_2206 = ($signed(_zz_2207) >>> _zz_164);
  assign _zz_2207 = _zz_2208;
  assign _zz_2208 = ($signed(_zz_2210) - $signed(_zz_161));
  assign _zz_2209 = ({8'd0,data_mid_0_real} <<< 8);
  assign _zz_2210 = {{8{_zz_2209[23]}}, _zz_2209};
  assign _zz_2211 = fixTo_194_dout;
  assign _zz_2212 = _zz_2213[31 : 0];
  assign _zz_2213 = _zz_2214;
  assign _zz_2214 = ($signed(_zz_2215) >>> _zz_164);
  assign _zz_2215 = _zz_2216;
  assign _zz_2216 = ($signed(_zz_2218) - $signed(_zz_162));
  assign _zz_2217 = ({8'd0,data_mid_0_imag} <<< 8);
  assign _zz_2218 = {{8{_zz_2217[23]}}, _zz_2217};
  assign _zz_2219 = fixTo_195_dout;
  assign _zz_2220 = _zz_2221[31 : 0];
  assign _zz_2221 = _zz_2222;
  assign _zz_2222 = ($signed(_zz_2223) >>> _zz_165);
  assign _zz_2223 = _zz_2224;
  assign _zz_2224 = ($signed(_zz_2226) + $signed(_zz_161));
  assign _zz_2225 = ({8'd0,data_mid_0_real} <<< 8);
  assign _zz_2226 = {{8{_zz_2225[23]}}, _zz_2225};
  assign _zz_2227 = fixTo_196_dout;
  assign _zz_2228 = _zz_2229[31 : 0];
  assign _zz_2229 = _zz_2230;
  assign _zz_2230 = ($signed(_zz_2231) >>> _zz_165);
  assign _zz_2231 = _zz_2232;
  assign _zz_2232 = ($signed(_zz_2234) + $signed(_zz_162));
  assign _zz_2233 = ({8'd0,data_mid_0_imag} <<< 8);
  assign _zz_2234 = {{8{_zz_2233[23]}}, _zz_2233};
  assign _zz_2235 = fixTo_197_dout;
  assign _zz_2236 = ($signed(twiddle_factor_table_4_real) + $signed(twiddle_factor_table_4_imag));
  assign _zz_2237 = ($signed(_zz_168) - $signed(_zz_2238));
  assign _zz_2238 = ($signed(_zz_2239) * $signed(twiddle_factor_table_4_imag));
  assign _zz_2239 = ($signed(data_mid_5_real) + $signed(data_mid_5_imag));
  assign _zz_2240 = fixTo_198_dout;
  assign _zz_2241 = ($signed(_zz_168) + $signed(_zz_2242));
  assign _zz_2242 = ($signed(_zz_2243) * $signed(twiddle_factor_table_4_real));
  assign _zz_2243 = ($signed(data_mid_5_imag) - $signed(data_mid_5_real));
  assign _zz_2244 = fixTo_199_dout;
  assign _zz_2245 = _zz_2246[31 : 0];
  assign _zz_2246 = _zz_2247;
  assign _zz_2247 = ($signed(_zz_2248) >>> _zz_169);
  assign _zz_2248 = _zz_2249;
  assign _zz_2249 = ($signed(_zz_2251) - $signed(_zz_166));
  assign _zz_2250 = ({8'd0,data_mid_1_real} <<< 8);
  assign _zz_2251 = {{8{_zz_2250[23]}}, _zz_2250};
  assign _zz_2252 = fixTo_200_dout;
  assign _zz_2253 = _zz_2254[31 : 0];
  assign _zz_2254 = _zz_2255;
  assign _zz_2255 = ($signed(_zz_2256) >>> _zz_169);
  assign _zz_2256 = _zz_2257;
  assign _zz_2257 = ($signed(_zz_2259) - $signed(_zz_167));
  assign _zz_2258 = ({8'd0,data_mid_1_imag} <<< 8);
  assign _zz_2259 = {{8{_zz_2258[23]}}, _zz_2258};
  assign _zz_2260 = fixTo_201_dout;
  assign _zz_2261 = _zz_2262[31 : 0];
  assign _zz_2262 = _zz_2263;
  assign _zz_2263 = ($signed(_zz_2264) >>> _zz_170);
  assign _zz_2264 = _zz_2265;
  assign _zz_2265 = ($signed(_zz_2267) + $signed(_zz_166));
  assign _zz_2266 = ({8'd0,data_mid_1_real} <<< 8);
  assign _zz_2267 = {{8{_zz_2266[23]}}, _zz_2266};
  assign _zz_2268 = fixTo_202_dout;
  assign _zz_2269 = _zz_2270[31 : 0];
  assign _zz_2270 = _zz_2271;
  assign _zz_2271 = ($signed(_zz_2272) >>> _zz_170);
  assign _zz_2272 = _zz_2273;
  assign _zz_2273 = ($signed(_zz_2275) + $signed(_zz_167));
  assign _zz_2274 = ({8'd0,data_mid_1_imag} <<< 8);
  assign _zz_2275 = {{8{_zz_2274[23]}}, _zz_2274};
  assign _zz_2276 = fixTo_203_dout;
  assign _zz_2277 = ($signed(twiddle_factor_table_5_real) + $signed(twiddle_factor_table_5_imag));
  assign _zz_2278 = ($signed(_zz_173) - $signed(_zz_2279));
  assign _zz_2279 = ($signed(_zz_2280) * $signed(twiddle_factor_table_5_imag));
  assign _zz_2280 = ($signed(data_mid_6_real) + $signed(data_mid_6_imag));
  assign _zz_2281 = fixTo_204_dout;
  assign _zz_2282 = ($signed(_zz_173) + $signed(_zz_2283));
  assign _zz_2283 = ($signed(_zz_2284) * $signed(twiddle_factor_table_5_real));
  assign _zz_2284 = ($signed(data_mid_6_imag) - $signed(data_mid_6_real));
  assign _zz_2285 = fixTo_205_dout;
  assign _zz_2286 = _zz_2287[31 : 0];
  assign _zz_2287 = _zz_2288;
  assign _zz_2288 = ($signed(_zz_2289) >>> _zz_174);
  assign _zz_2289 = _zz_2290;
  assign _zz_2290 = ($signed(_zz_2292) - $signed(_zz_171));
  assign _zz_2291 = ({8'd0,data_mid_2_real} <<< 8);
  assign _zz_2292 = {{8{_zz_2291[23]}}, _zz_2291};
  assign _zz_2293 = fixTo_206_dout;
  assign _zz_2294 = _zz_2295[31 : 0];
  assign _zz_2295 = _zz_2296;
  assign _zz_2296 = ($signed(_zz_2297) >>> _zz_174);
  assign _zz_2297 = _zz_2298;
  assign _zz_2298 = ($signed(_zz_2300) - $signed(_zz_172));
  assign _zz_2299 = ({8'd0,data_mid_2_imag} <<< 8);
  assign _zz_2300 = {{8{_zz_2299[23]}}, _zz_2299};
  assign _zz_2301 = fixTo_207_dout;
  assign _zz_2302 = _zz_2303[31 : 0];
  assign _zz_2303 = _zz_2304;
  assign _zz_2304 = ($signed(_zz_2305) >>> _zz_175);
  assign _zz_2305 = _zz_2306;
  assign _zz_2306 = ($signed(_zz_2308) + $signed(_zz_171));
  assign _zz_2307 = ({8'd0,data_mid_2_real} <<< 8);
  assign _zz_2308 = {{8{_zz_2307[23]}}, _zz_2307};
  assign _zz_2309 = fixTo_208_dout;
  assign _zz_2310 = _zz_2311[31 : 0];
  assign _zz_2311 = _zz_2312;
  assign _zz_2312 = ($signed(_zz_2313) >>> _zz_175);
  assign _zz_2313 = _zz_2314;
  assign _zz_2314 = ($signed(_zz_2316) + $signed(_zz_172));
  assign _zz_2315 = ({8'd0,data_mid_2_imag} <<< 8);
  assign _zz_2316 = {{8{_zz_2315[23]}}, _zz_2315};
  assign _zz_2317 = fixTo_209_dout;
  assign _zz_2318 = ($signed(twiddle_factor_table_6_real) + $signed(twiddle_factor_table_6_imag));
  assign _zz_2319 = ($signed(_zz_178) - $signed(_zz_2320));
  assign _zz_2320 = ($signed(_zz_2321) * $signed(twiddle_factor_table_6_imag));
  assign _zz_2321 = ($signed(data_mid_7_real) + $signed(data_mid_7_imag));
  assign _zz_2322 = fixTo_210_dout;
  assign _zz_2323 = ($signed(_zz_178) + $signed(_zz_2324));
  assign _zz_2324 = ($signed(_zz_2325) * $signed(twiddle_factor_table_6_real));
  assign _zz_2325 = ($signed(data_mid_7_imag) - $signed(data_mid_7_real));
  assign _zz_2326 = fixTo_211_dout;
  assign _zz_2327 = _zz_2328[31 : 0];
  assign _zz_2328 = _zz_2329;
  assign _zz_2329 = ($signed(_zz_2330) >>> _zz_179);
  assign _zz_2330 = _zz_2331;
  assign _zz_2331 = ($signed(_zz_2333) - $signed(_zz_176));
  assign _zz_2332 = ({8'd0,data_mid_3_real} <<< 8);
  assign _zz_2333 = {{8{_zz_2332[23]}}, _zz_2332};
  assign _zz_2334 = fixTo_212_dout;
  assign _zz_2335 = _zz_2336[31 : 0];
  assign _zz_2336 = _zz_2337;
  assign _zz_2337 = ($signed(_zz_2338) >>> _zz_179);
  assign _zz_2338 = _zz_2339;
  assign _zz_2339 = ($signed(_zz_2341) - $signed(_zz_177));
  assign _zz_2340 = ({8'd0,data_mid_3_imag} <<< 8);
  assign _zz_2341 = {{8{_zz_2340[23]}}, _zz_2340};
  assign _zz_2342 = fixTo_213_dout;
  assign _zz_2343 = _zz_2344[31 : 0];
  assign _zz_2344 = _zz_2345;
  assign _zz_2345 = ($signed(_zz_2346) >>> _zz_180);
  assign _zz_2346 = _zz_2347;
  assign _zz_2347 = ($signed(_zz_2349) + $signed(_zz_176));
  assign _zz_2348 = ({8'd0,data_mid_3_real} <<< 8);
  assign _zz_2349 = {{8{_zz_2348[23]}}, _zz_2348};
  assign _zz_2350 = fixTo_214_dout;
  assign _zz_2351 = _zz_2352[31 : 0];
  assign _zz_2352 = _zz_2353;
  assign _zz_2353 = ($signed(_zz_2354) >>> _zz_180);
  assign _zz_2354 = _zz_2355;
  assign _zz_2355 = ($signed(_zz_2357) + $signed(_zz_177));
  assign _zz_2356 = ({8'd0,data_mid_3_imag} <<< 8);
  assign _zz_2357 = {{8{_zz_2356[23]}}, _zz_2356};
  assign _zz_2358 = fixTo_215_dout;
  assign _zz_2359 = ($signed(twiddle_factor_table_3_real) + $signed(twiddle_factor_table_3_imag));
  assign _zz_2360 = ($signed(_zz_183) - $signed(_zz_2361));
  assign _zz_2361 = ($signed(_zz_2362) * $signed(twiddle_factor_table_3_imag));
  assign _zz_2362 = ($signed(data_mid_12_real) + $signed(data_mid_12_imag));
  assign _zz_2363 = fixTo_216_dout;
  assign _zz_2364 = ($signed(_zz_183) + $signed(_zz_2365));
  assign _zz_2365 = ($signed(_zz_2366) * $signed(twiddle_factor_table_3_real));
  assign _zz_2366 = ($signed(data_mid_12_imag) - $signed(data_mid_12_real));
  assign _zz_2367 = fixTo_217_dout;
  assign _zz_2368 = _zz_2369[31 : 0];
  assign _zz_2369 = _zz_2370;
  assign _zz_2370 = ($signed(_zz_2371) >>> _zz_184);
  assign _zz_2371 = _zz_2372;
  assign _zz_2372 = ($signed(_zz_2374) - $signed(_zz_181));
  assign _zz_2373 = ({8'd0,data_mid_8_real} <<< 8);
  assign _zz_2374 = {{8{_zz_2373[23]}}, _zz_2373};
  assign _zz_2375 = fixTo_218_dout;
  assign _zz_2376 = _zz_2377[31 : 0];
  assign _zz_2377 = _zz_2378;
  assign _zz_2378 = ($signed(_zz_2379) >>> _zz_184);
  assign _zz_2379 = _zz_2380;
  assign _zz_2380 = ($signed(_zz_2382) - $signed(_zz_182));
  assign _zz_2381 = ({8'd0,data_mid_8_imag} <<< 8);
  assign _zz_2382 = {{8{_zz_2381[23]}}, _zz_2381};
  assign _zz_2383 = fixTo_219_dout;
  assign _zz_2384 = _zz_2385[31 : 0];
  assign _zz_2385 = _zz_2386;
  assign _zz_2386 = ($signed(_zz_2387) >>> _zz_185);
  assign _zz_2387 = _zz_2388;
  assign _zz_2388 = ($signed(_zz_2390) + $signed(_zz_181));
  assign _zz_2389 = ({8'd0,data_mid_8_real} <<< 8);
  assign _zz_2390 = {{8{_zz_2389[23]}}, _zz_2389};
  assign _zz_2391 = fixTo_220_dout;
  assign _zz_2392 = _zz_2393[31 : 0];
  assign _zz_2393 = _zz_2394;
  assign _zz_2394 = ($signed(_zz_2395) >>> _zz_185);
  assign _zz_2395 = _zz_2396;
  assign _zz_2396 = ($signed(_zz_2398) + $signed(_zz_182));
  assign _zz_2397 = ({8'd0,data_mid_8_imag} <<< 8);
  assign _zz_2398 = {{8{_zz_2397[23]}}, _zz_2397};
  assign _zz_2399 = fixTo_221_dout;
  assign _zz_2400 = ($signed(twiddle_factor_table_4_real) + $signed(twiddle_factor_table_4_imag));
  assign _zz_2401 = ($signed(_zz_188) - $signed(_zz_2402));
  assign _zz_2402 = ($signed(_zz_2403) * $signed(twiddle_factor_table_4_imag));
  assign _zz_2403 = ($signed(data_mid_13_real) + $signed(data_mid_13_imag));
  assign _zz_2404 = fixTo_222_dout;
  assign _zz_2405 = ($signed(_zz_188) + $signed(_zz_2406));
  assign _zz_2406 = ($signed(_zz_2407) * $signed(twiddle_factor_table_4_real));
  assign _zz_2407 = ($signed(data_mid_13_imag) - $signed(data_mid_13_real));
  assign _zz_2408 = fixTo_223_dout;
  assign _zz_2409 = _zz_2410[31 : 0];
  assign _zz_2410 = _zz_2411;
  assign _zz_2411 = ($signed(_zz_2412) >>> _zz_189);
  assign _zz_2412 = _zz_2413;
  assign _zz_2413 = ($signed(_zz_2415) - $signed(_zz_186));
  assign _zz_2414 = ({8'd0,data_mid_9_real} <<< 8);
  assign _zz_2415 = {{8{_zz_2414[23]}}, _zz_2414};
  assign _zz_2416 = fixTo_224_dout;
  assign _zz_2417 = _zz_2418[31 : 0];
  assign _zz_2418 = _zz_2419;
  assign _zz_2419 = ($signed(_zz_2420) >>> _zz_189);
  assign _zz_2420 = _zz_2421;
  assign _zz_2421 = ($signed(_zz_2423) - $signed(_zz_187));
  assign _zz_2422 = ({8'd0,data_mid_9_imag} <<< 8);
  assign _zz_2423 = {{8{_zz_2422[23]}}, _zz_2422};
  assign _zz_2424 = fixTo_225_dout;
  assign _zz_2425 = _zz_2426[31 : 0];
  assign _zz_2426 = _zz_2427;
  assign _zz_2427 = ($signed(_zz_2428) >>> _zz_190);
  assign _zz_2428 = _zz_2429;
  assign _zz_2429 = ($signed(_zz_2431) + $signed(_zz_186));
  assign _zz_2430 = ({8'd0,data_mid_9_real} <<< 8);
  assign _zz_2431 = {{8{_zz_2430[23]}}, _zz_2430};
  assign _zz_2432 = fixTo_226_dout;
  assign _zz_2433 = _zz_2434[31 : 0];
  assign _zz_2434 = _zz_2435;
  assign _zz_2435 = ($signed(_zz_2436) >>> _zz_190);
  assign _zz_2436 = _zz_2437;
  assign _zz_2437 = ($signed(_zz_2439) + $signed(_zz_187));
  assign _zz_2438 = ({8'd0,data_mid_9_imag} <<< 8);
  assign _zz_2439 = {{8{_zz_2438[23]}}, _zz_2438};
  assign _zz_2440 = fixTo_227_dout;
  assign _zz_2441 = ($signed(twiddle_factor_table_5_real) + $signed(twiddle_factor_table_5_imag));
  assign _zz_2442 = ($signed(_zz_193) - $signed(_zz_2443));
  assign _zz_2443 = ($signed(_zz_2444) * $signed(twiddle_factor_table_5_imag));
  assign _zz_2444 = ($signed(data_mid_14_real) + $signed(data_mid_14_imag));
  assign _zz_2445 = fixTo_228_dout;
  assign _zz_2446 = ($signed(_zz_193) + $signed(_zz_2447));
  assign _zz_2447 = ($signed(_zz_2448) * $signed(twiddle_factor_table_5_real));
  assign _zz_2448 = ($signed(data_mid_14_imag) - $signed(data_mid_14_real));
  assign _zz_2449 = fixTo_229_dout;
  assign _zz_2450 = _zz_2451[31 : 0];
  assign _zz_2451 = _zz_2452;
  assign _zz_2452 = ($signed(_zz_2453) >>> _zz_194);
  assign _zz_2453 = _zz_2454;
  assign _zz_2454 = ($signed(_zz_2456) - $signed(_zz_191));
  assign _zz_2455 = ({8'd0,data_mid_10_real} <<< 8);
  assign _zz_2456 = {{8{_zz_2455[23]}}, _zz_2455};
  assign _zz_2457 = fixTo_230_dout;
  assign _zz_2458 = _zz_2459[31 : 0];
  assign _zz_2459 = _zz_2460;
  assign _zz_2460 = ($signed(_zz_2461) >>> _zz_194);
  assign _zz_2461 = _zz_2462;
  assign _zz_2462 = ($signed(_zz_2464) - $signed(_zz_192));
  assign _zz_2463 = ({8'd0,data_mid_10_imag} <<< 8);
  assign _zz_2464 = {{8{_zz_2463[23]}}, _zz_2463};
  assign _zz_2465 = fixTo_231_dout;
  assign _zz_2466 = _zz_2467[31 : 0];
  assign _zz_2467 = _zz_2468;
  assign _zz_2468 = ($signed(_zz_2469) >>> _zz_195);
  assign _zz_2469 = _zz_2470;
  assign _zz_2470 = ($signed(_zz_2472) + $signed(_zz_191));
  assign _zz_2471 = ({8'd0,data_mid_10_real} <<< 8);
  assign _zz_2472 = {{8{_zz_2471[23]}}, _zz_2471};
  assign _zz_2473 = fixTo_232_dout;
  assign _zz_2474 = _zz_2475[31 : 0];
  assign _zz_2475 = _zz_2476;
  assign _zz_2476 = ($signed(_zz_2477) >>> _zz_195);
  assign _zz_2477 = _zz_2478;
  assign _zz_2478 = ($signed(_zz_2480) + $signed(_zz_192));
  assign _zz_2479 = ({8'd0,data_mid_10_imag} <<< 8);
  assign _zz_2480 = {{8{_zz_2479[23]}}, _zz_2479};
  assign _zz_2481 = fixTo_233_dout;
  assign _zz_2482 = ($signed(twiddle_factor_table_6_real) + $signed(twiddle_factor_table_6_imag));
  assign _zz_2483 = ($signed(_zz_198) - $signed(_zz_2484));
  assign _zz_2484 = ($signed(_zz_2485) * $signed(twiddle_factor_table_6_imag));
  assign _zz_2485 = ($signed(data_mid_15_real) + $signed(data_mid_15_imag));
  assign _zz_2486 = fixTo_234_dout;
  assign _zz_2487 = ($signed(_zz_198) + $signed(_zz_2488));
  assign _zz_2488 = ($signed(_zz_2489) * $signed(twiddle_factor_table_6_real));
  assign _zz_2489 = ($signed(data_mid_15_imag) - $signed(data_mid_15_real));
  assign _zz_2490 = fixTo_235_dout;
  assign _zz_2491 = _zz_2492[31 : 0];
  assign _zz_2492 = _zz_2493;
  assign _zz_2493 = ($signed(_zz_2494) >>> _zz_199);
  assign _zz_2494 = _zz_2495;
  assign _zz_2495 = ($signed(_zz_2497) - $signed(_zz_196));
  assign _zz_2496 = ({8'd0,data_mid_11_real} <<< 8);
  assign _zz_2497 = {{8{_zz_2496[23]}}, _zz_2496};
  assign _zz_2498 = fixTo_236_dout;
  assign _zz_2499 = _zz_2500[31 : 0];
  assign _zz_2500 = _zz_2501;
  assign _zz_2501 = ($signed(_zz_2502) >>> _zz_199);
  assign _zz_2502 = _zz_2503;
  assign _zz_2503 = ($signed(_zz_2505) - $signed(_zz_197));
  assign _zz_2504 = ({8'd0,data_mid_11_imag} <<< 8);
  assign _zz_2505 = {{8{_zz_2504[23]}}, _zz_2504};
  assign _zz_2506 = fixTo_237_dout;
  assign _zz_2507 = _zz_2508[31 : 0];
  assign _zz_2508 = _zz_2509;
  assign _zz_2509 = ($signed(_zz_2510) >>> _zz_200);
  assign _zz_2510 = _zz_2511;
  assign _zz_2511 = ($signed(_zz_2513) + $signed(_zz_196));
  assign _zz_2512 = ({8'd0,data_mid_11_real} <<< 8);
  assign _zz_2513 = {{8{_zz_2512[23]}}, _zz_2512};
  assign _zz_2514 = fixTo_238_dout;
  assign _zz_2515 = _zz_2516[31 : 0];
  assign _zz_2516 = _zz_2517;
  assign _zz_2517 = ($signed(_zz_2518) >>> _zz_200);
  assign _zz_2518 = _zz_2519;
  assign _zz_2519 = ($signed(_zz_2521) + $signed(_zz_197));
  assign _zz_2520 = ({8'd0,data_mid_11_imag} <<< 8);
  assign _zz_2521 = {{8{_zz_2520[23]}}, _zz_2520};
  assign _zz_2522 = fixTo_239_dout;
  assign _zz_2523 = ($signed(twiddle_factor_table_3_real) + $signed(twiddle_factor_table_3_imag));
  assign _zz_2524 = ($signed(_zz_203) - $signed(_zz_2525));
  assign _zz_2525 = ($signed(_zz_2526) * $signed(twiddle_factor_table_3_imag));
  assign _zz_2526 = ($signed(data_mid_20_real) + $signed(data_mid_20_imag));
  assign _zz_2527 = fixTo_240_dout;
  assign _zz_2528 = ($signed(_zz_203) + $signed(_zz_2529));
  assign _zz_2529 = ($signed(_zz_2530) * $signed(twiddle_factor_table_3_real));
  assign _zz_2530 = ($signed(data_mid_20_imag) - $signed(data_mid_20_real));
  assign _zz_2531 = fixTo_241_dout;
  assign _zz_2532 = _zz_2533[31 : 0];
  assign _zz_2533 = _zz_2534;
  assign _zz_2534 = ($signed(_zz_2535) >>> _zz_204);
  assign _zz_2535 = _zz_2536;
  assign _zz_2536 = ($signed(_zz_2538) - $signed(_zz_201));
  assign _zz_2537 = ({8'd0,data_mid_16_real} <<< 8);
  assign _zz_2538 = {{8{_zz_2537[23]}}, _zz_2537};
  assign _zz_2539 = fixTo_242_dout;
  assign _zz_2540 = _zz_2541[31 : 0];
  assign _zz_2541 = _zz_2542;
  assign _zz_2542 = ($signed(_zz_2543) >>> _zz_204);
  assign _zz_2543 = _zz_2544;
  assign _zz_2544 = ($signed(_zz_2546) - $signed(_zz_202));
  assign _zz_2545 = ({8'd0,data_mid_16_imag} <<< 8);
  assign _zz_2546 = {{8{_zz_2545[23]}}, _zz_2545};
  assign _zz_2547 = fixTo_243_dout;
  assign _zz_2548 = _zz_2549[31 : 0];
  assign _zz_2549 = _zz_2550;
  assign _zz_2550 = ($signed(_zz_2551) >>> _zz_205);
  assign _zz_2551 = _zz_2552;
  assign _zz_2552 = ($signed(_zz_2554) + $signed(_zz_201));
  assign _zz_2553 = ({8'd0,data_mid_16_real} <<< 8);
  assign _zz_2554 = {{8{_zz_2553[23]}}, _zz_2553};
  assign _zz_2555 = fixTo_244_dout;
  assign _zz_2556 = _zz_2557[31 : 0];
  assign _zz_2557 = _zz_2558;
  assign _zz_2558 = ($signed(_zz_2559) >>> _zz_205);
  assign _zz_2559 = _zz_2560;
  assign _zz_2560 = ($signed(_zz_2562) + $signed(_zz_202));
  assign _zz_2561 = ({8'd0,data_mid_16_imag} <<< 8);
  assign _zz_2562 = {{8{_zz_2561[23]}}, _zz_2561};
  assign _zz_2563 = fixTo_245_dout;
  assign _zz_2564 = ($signed(twiddle_factor_table_4_real) + $signed(twiddle_factor_table_4_imag));
  assign _zz_2565 = ($signed(_zz_208) - $signed(_zz_2566));
  assign _zz_2566 = ($signed(_zz_2567) * $signed(twiddle_factor_table_4_imag));
  assign _zz_2567 = ($signed(data_mid_21_real) + $signed(data_mid_21_imag));
  assign _zz_2568 = fixTo_246_dout;
  assign _zz_2569 = ($signed(_zz_208) + $signed(_zz_2570));
  assign _zz_2570 = ($signed(_zz_2571) * $signed(twiddle_factor_table_4_real));
  assign _zz_2571 = ($signed(data_mid_21_imag) - $signed(data_mid_21_real));
  assign _zz_2572 = fixTo_247_dout;
  assign _zz_2573 = _zz_2574[31 : 0];
  assign _zz_2574 = _zz_2575;
  assign _zz_2575 = ($signed(_zz_2576) >>> _zz_209);
  assign _zz_2576 = _zz_2577;
  assign _zz_2577 = ($signed(_zz_2579) - $signed(_zz_206));
  assign _zz_2578 = ({8'd0,data_mid_17_real} <<< 8);
  assign _zz_2579 = {{8{_zz_2578[23]}}, _zz_2578};
  assign _zz_2580 = fixTo_248_dout;
  assign _zz_2581 = _zz_2582[31 : 0];
  assign _zz_2582 = _zz_2583;
  assign _zz_2583 = ($signed(_zz_2584) >>> _zz_209);
  assign _zz_2584 = _zz_2585;
  assign _zz_2585 = ($signed(_zz_2587) - $signed(_zz_207));
  assign _zz_2586 = ({8'd0,data_mid_17_imag} <<< 8);
  assign _zz_2587 = {{8{_zz_2586[23]}}, _zz_2586};
  assign _zz_2588 = fixTo_249_dout;
  assign _zz_2589 = _zz_2590[31 : 0];
  assign _zz_2590 = _zz_2591;
  assign _zz_2591 = ($signed(_zz_2592) >>> _zz_210);
  assign _zz_2592 = _zz_2593;
  assign _zz_2593 = ($signed(_zz_2595) + $signed(_zz_206));
  assign _zz_2594 = ({8'd0,data_mid_17_real} <<< 8);
  assign _zz_2595 = {{8{_zz_2594[23]}}, _zz_2594};
  assign _zz_2596 = fixTo_250_dout;
  assign _zz_2597 = _zz_2598[31 : 0];
  assign _zz_2598 = _zz_2599;
  assign _zz_2599 = ($signed(_zz_2600) >>> _zz_210);
  assign _zz_2600 = _zz_2601;
  assign _zz_2601 = ($signed(_zz_2603) + $signed(_zz_207));
  assign _zz_2602 = ({8'd0,data_mid_17_imag} <<< 8);
  assign _zz_2603 = {{8{_zz_2602[23]}}, _zz_2602};
  assign _zz_2604 = fixTo_251_dout;
  assign _zz_2605 = ($signed(twiddle_factor_table_5_real) + $signed(twiddle_factor_table_5_imag));
  assign _zz_2606 = ($signed(_zz_213) - $signed(_zz_2607));
  assign _zz_2607 = ($signed(_zz_2608) * $signed(twiddle_factor_table_5_imag));
  assign _zz_2608 = ($signed(data_mid_22_real) + $signed(data_mid_22_imag));
  assign _zz_2609 = fixTo_252_dout;
  assign _zz_2610 = ($signed(_zz_213) + $signed(_zz_2611));
  assign _zz_2611 = ($signed(_zz_2612) * $signed(twiddle_factor_table_5_real));
  assign _zz_2612 = ($signed(data_mid_22_imag) - $signed(data_mid_22_real));
  assign _zz_2613 = fixTo_253_dout;
  assign _zz_2614 = _zz_2615[31 : 0];
  assign _zz_2615 = _zz_2616;
  assign _zz_2616 = ($signed(_zz_2617) >>> _zz_214);
  assign _zz_2617 = _zz_2618;
  assign _zz_2618 = ($signed(_zz_2620) - $signed(_zz_211));
  assign _zz_2619 = ({8'd0,data_mid_18_real} <<< 8);
  assign _zz_2620 = {{8{_zz_2619[23]}}, _zz_2619};
  assign _zz_2621 = fixTo_254_dout;
  assign _zz_2622 = _zz_2623[31 : 0];
  assign _zz_2623 = _zz_2624;
  assign _zz_2624 = ($signed(_zz_2625) >>> _zz_214);
  assign _zz_2625 = _zz_2626;
  assign _zz_2626 = ($signed(_zz_2628) - $signed(_zz_212));
  assign _zz_2627 = ({8'd0,data_mid_18_imag} <<< 8);
  assign _zz_2628 = {{8{_zz_2627[23]}}, _zz_2627};
  assign _zz_2629 = fixTo_255_dout;
  assign _zz_2630 = _zz_2631[31 : 0];
  assign _zz_2631 = _zz_2632;
  assign _zz_2632 = ($signed(_zz_2633) >>> _zz_215);
  assign _zz_2633 = _zz_2634;
  assign _zz_2634 = ($signed(_zz_2636) + $signed(_zz_211));
  assign _zz_2635 = ({8'd0,data_mid_18_real} <<< 8);
  assign _zz_2636 = {{8{_zz_2635[23]}}, _zz_2635};
  assign _zz_2637 = fixTo_256_dout;
  assign _zz_2638 = _zz_2639[31 : 0];
  assign _zz_2639 = _zz_2640;
  assign _zz_2640 = ($signed(_zz_2641) >>> _zz_215);
  assign _zz_2641 = _zz_2642;
  assign _zz_2642 = ($signed(_zz_2644) + $signed(_zz_212));
  assign _zz_2643 = ({8'd0,data_mid_18_imag} <<< 8);
  assign _zz_2644 = {{8{_zz_2643[23]}}, _zz_2643};
  assign _zz_2645 = fixTo_257_dout;
  assign _zz_2646 = ($signed(twiddle_factor_table_6_real) + $signed(twiddle_factor_table_6_imag));
  assign _zz_2647 = ($signed(_zz_218) - $signed(_zz_2648));
  assign _zz_2648 = ($signed(_zz_2649) * $signed(twiddle_factor_table_6_imag));
  assign _zz_2649 = ($signed(data_mid_23_real) + $signed(data_mid_23_imag));
  assign _zz_2650 = fixTo_258_dout;
  assign _zz_2651 = ($signed(_zz_218) + $signed(_zz_2652));
  assign _zz_2652 = ($signed(_zz_2653) * $signed(twiddle_factor_table_6_real));
  assign _zz_2653 = ($signed(data_mid_23_imag) - $signed(data_mid_23_real));
  assign _zz_2654 = fixTo_259_dout;
  assign _zz_2655 = _zz_2656[31 : 0];
  assign _zz_2656 = _zz_2657;
  assign _zz_2657 = ($signed(_zz_2658) >>> _zz_219);
  assign _zz_2658 = _zz_2659;
  assign _zz_2659 = ($signed(_zz_2661) - $signed(_zz_216));
  assign _zz_2660 = ({8'd0,data_mid_19_real} <<< 8);
  assign _zz_2661 = {{8{_zz_2660[23]}}, _zz_2660};
  assign _zz_2662 = fixTo_260_dout;
  assign _zz_2663 = _zz_2664[31 : 0];
  assign _zz_2664 = _zz_2665;
  assign _zz_2665 = ($signed(_zz_2666) >>> _zz_219);
  assign _zz_2666 = _zz_2667;
  assign _zz_2667 = ($signed(_zz_2669) - $signed(_zz_217));
  assign _zz_2668 = ({8'd0,data_mid_19_imag} <<< 8);
  assign _zz_2669 = {{8{_zz_2668[23]}}, _zz_2668};
  assign _zz_2670 = fixTo_261_dout;
  assign _zz_2671 = _zz_2672[31 : 0];
  assign _zz_2672 = _zz_2673;
  assign _zz_2673 = ($signed(_zz_2674) >>> _zz_220);
  assign _zz_2674 = _zz_2675;
  assign _zz_2675 = ($signed(_zz_2677) + $signed(_zz_216));
  assign _zz_2676 = ({8'd0,data_mid_19_real} <<< 8);
  assign _zz_2677 = {{8{_zz_2676[23]}}, _zz_2676};
  assign _zz_2678 = fixTo_262_dout;
  assign _zz_2679 = _zz_2680[31 : 0];
  assign _zz_2680 = _zz_2681;
  assign _zz_2681 = ($signed(_zz_2682) >>> _zz_220);
  assign _zz_2682 = _zz_2683;
  assign _zz_2683 = ($signed(_zz_2685) + $signed(_zz_217));
  assign _zz_2684 = ({8'd0,data_mid_19_imag} <<< 8);
  assign _zz_2685 = {{8{_zz_2684[23]}}, _zz_2684};
  assign _zz_2686 = fixTo_263_dout;
  assign _zz_2687 = ($signed(twiddle_factor_table_3_real) + $signed(twiddle_factor_table_3_imag));
  assign _zz_2688 = ($signed(_zz_223) - $signed(_zz_2689));
  assign _zz_2689 = ($signed(_zz_2690) * $signed(twiddle_factor_table_3_imag));
  assign _zz_2690 = ($signed(data_mid_28_real) + $signed(data_mid_28_imag));
  assign _zz_2691 = fixTo_264_dout;
  assign _zz_2692 = ($signed(_zz_223) + $signed(_zz_2693));
  assign _zz_2693 = ($signed(_zz_2694) * $signed(twiddle_factor_table_3_real));
  assign _zz_2694 = ($signed(data_mid_28_imag) - $signed(data_mid_28_real));
  assign _zz_2695 = fixTo_265_dout;
  assign _zz_2696 = _zz_2697[31 : 0];
  assign _zz_2697 = _zz_2698;
  assign _zz_2698 = ($signed(_zz_2699) >>> _zz_224);
  assign _zz_2699 = _zz_2700;
  assign _zz_2700 = ($signed(_zz_2702) - $signed(_zz_221));
  assign _zz_2701 = ({8'd0,data_mid_24_real} <<< 8);
  assign _zz_2702 = {{8{_zz_2701[23]}}, _zz_2701};
  assign _zz_2703 = fixTo_266_dout;
  assign _zz_2704 = _zz_2705[31 : 0];
  assign _zz_2705 = _zz_2706;
  assign _zz_2706 = ($signed(_zz_2707) >>> _zz_224);
  assign _zz_2707 = _zz_2708;
  assign _zz_2708 = ($signed(_zz_2710) - $signed(_zz_222));
  assign _zz_2709 = ({8'd0,data_mid_24_imag} <<< 8);
  assign _zz_2710 = {{8{_zz_2709[23]}}, _zz_2709};
  assign _zz_2711 = fixTo_267_dout;
  assign _zz_2712 = _zz_2713[31 : 0];
  assign _zz_2713 = _zz_2714;
  assign _zz_2714 = ($signed(_zz_2715) >>> _zz_225);
  assign _zz_2715 = _zz_2716;
  assign _zz_2716 = ($signed(_zz_2718) + $signed(_zz_221));
  assign _zz_2717 = ({8'd0,data_mid_24_real} <<< 8);
  assign _zz_2718 = {{8{_zz_2717[23]}}, _zz_2717};
  assign _zz_2719 = fixTo_268_dout;
  assign _zz_2720 = _zz_2721[31 : 0];
  assign _zz_2721 = _zz_2722;
  assign _zz_2722 = ($signed(_zz_2723) >>> _zz_225);
  assign _zz_2723 = _zz_2724;
  assign _zz_2724 = ($signed(_zz_2726) + $signed(_zz_222));
  assign _zz_2725 = ({8'd0,data_mid_24_imag} <<< 8);
  assign _zz_2726 = {{8{_zz_2725[23]}}, _zz_2725};
  assign _zz_2727 = fixTo_269_dout;
  assign _zz_2728 = ($signed(twiddle_factor_table_4_real) + $signed(twiddle_factor_table_4_imag));
  assign _zz_2729 = ($signed(_zz_228) - $signed(_zz_2730));
  assign _zz_2730 = ($signed(_zz_2731) * $signed(twiddle_factor_table_4_imag));
  assign _zz_2731 = ($signed(data_mid_29_real) + $signed(data_mid_29_imag));
  assign _zz_2732 = fixTo_270_dout;
  assign _zz_2733 = ($signed(_zz_228) + $signed(_zz_2734));
  assign _zz_2734 = ($signed(_zz_2735) * $signed(twiddle_factor_table_4_real));
  assign _zz_2735 = ($signed(data_mid_29_imag) - $signed(data_mid_29_real));
  assign _zz_2736 = fixTo_271_dout;
  assign _zz_2737 = _zz_2738[31 : 0];
  assign _zz_2738 = _zz_2739;
  assign _zz_2739 = ($signed(_zz_2740) >>> _zz_229);
  assign _zz_2740 = _zz_2741;
  assign _zz_2741 = ($signed(_zz_2743) - $signed(_zz_226));
  assign _zz_2742 = ({8'd0,data_mid_25_real} <<< 8);
  assign _zz_2743 = {{8{_zz_2742[23]}}, _zz_2742};
  assign _zz_2744 = fixTo_272_dout;
  assign _zz_2745 = _zz_2746[31 : 0];
  assign _zz_2746 = _zz_2747;
  assign _zz_2747 = ($signed(_zz_2748) >>> _zz_229);
  assign _zz_2748 = _zz_2749;
  assign _zz_2749 = ($signed(_zz_2751) - $signed(_zz_227));
  assign _zz_2750 = ({8'd0,data_mid_25_imag} <<< 8);
  assign _zz_2751 = {{8{_zz_2750[23]}}, _zz_2750};
  assign _zz_2752 = fixTo_273_dout;
  assign _zz_2753 = _zz_2754[31 : 0];
  assign _zz_2754 = _zz_2755;
  assign _zz_2755 = ($signed(_zz_2756) >>> _zz_230);
  assign _zz_2756 = _zz_2757;
  assign _zz_2757 = ($signed(_zz_2759) + $signed(_zz_226));
  assign _zz_2758 = ({8'd0,data_mid_25_real} <<< 8);
  assign _zz_2759 = {{8{_zz_2758[23]}}, _zz_2758};
  assign _zz_2760 = fixTo_274_dout;
  assign _zz_2761 = _zz_2762[31 : 0];
  assign _zz_2762 = _zz_2763;
  assign _zz_2763 = ($signed(_zz_2764) >>> _zz_230);
  assign _zz_2764 = _zz_2765;
  assign _zz_2765 = ($signed(_zz_2767) + $signed(_zz_227));
  assign _zz_2766 = ({8'd0,data_mid_25_imag} <<< 8);
  assign _zz_2767 = {{8{_zz_2766[23]}}, _zz_2766};
  assign _zz_2768 = fixTo_275_dout;
  assign _zz_2769 = ($signed(twiddle_factor_table_5_real) + $signed(twiddle_factor_table_5_imag));
  assign _zz_2770 = ($signed(_zz_233) - $signed(_zz_2771));
  assign _zz_2771 = ($signed(_zz_2772) * $signed(twiddle_factor_table_5_imag));
  assign _zz_2772 = ($signed(data_mid_30_real) + $signed(data_mid_30_imag));
  assign _zz_2773 = fixTo_276_dout;
  assign _zz_2774 = ($signed(_zz_233) + $signed(_zz_2775));
  assign _zz_2775 = ($signed(_zz_2776) * $signed(twiddle_factor_table_5_real));
  assign _zz_2776 = ($signed(data_mid_30_imag) - $signed(data_mid_30_real));
  assign _zz_2777 = fixTo_277_dout;
  assign _zz_2778 = _zz_2779[31 : 0];
  assign _zz_2779 = _zz_2780;
  assign _zz_2780 = ($signed(_zz_2781) >>> _zz_234);
  assign _zz_2781 = _zz_2782;
  assign _zz_2782 = ($signed(_zz_2784) - $signed(_zz_231));
  assign _zz_2783 = ({8'd0,data_mid_26_real} <<< 8);
  assign _zz_2784 = {{8{_zz_2783[23]}}, _zz_2783};
  assign _zz_2785 = fixTo_278_dout;
  assign _zz_2786 = _zz_2787[31 : 0];
  assign _zz_2787 = _zz_2788;
  assign _zz_2788 = ($signed(_zz_2789) >>> _zz_234);
  assign _zz_2789 = _zz_2790;
  assign _zz_2790 = ($signed(_zz_2792) - $signed(_zz_232));
  assign _zz_2791 = ({8'd0,data_mid_26_imag} <<< 8);
  assign _zz_2792 = {{8{_zz_2791[23]}}, _zz_2791};
  assign _zz_2793 = fixTo_279_dout;
  assign _zz_2794 = _zz_2795[31 : 0];
  assign _zz_2795 = _zz_2796;
  assign _zz_2796 = ($signed(_zz_2797) >>> _zz_235);
  assign _zz_2797 = _zz_2798;
  assign _zz_2798 = ($signed(_zz_2800) + $signed(_zz_231));
  assign _zz_2799 = ({8'd0,data_mid_26_real} <<< 8);
  assign _zz_2800 = {{8{_zz_2799[23]}}, _zz_2799};
  assign _zz_2801 = fixTo_280_dout;
  assign _zz_2802 = _zz_2803[31 : 0];
  assign _zz_2803 = _zz_2804;
  assign _zz_2804 = ($signed(_zz_2805) >>> _zz_235);
  assign _zz_2805 = _zz_2806;
  assign _zz_2806 = ($signed(_zz_2808) + $signed(_zz_232));
  assign _zz_2807 = ({8'd0,data_mid_26_imag} <<< 8);
  assign _zz_2808 = {{8{_zz_2807[23]}}, _zz_2807};
  assign _zz_2809 = fixTo_281_dout;
  assign _zz_2810 = ($signed(twiddle_factor_table_6_real) + $signed(twiddle_factor_table_6_imag));
  assign _zz_2811 = ($signed(_zz_238) - $signed(_zz_2812));
  assign _zz_2812 = ($signed(_zz_2813) * $signed(twiddle_factor_table_6_imag));
  assign _zz_2813 = ($signed(data_mid_31_real) + $signed(data_mid_31_imag));
  assign _zz_2814 = fixTo_282_dout;
  assign _zz_2815 = ($signed(_zz_238) + $signed(_zz_2816));
  assign _zz_2816 = ($signed(_zz_2817) * $signed(twiddle_factor_table_6_real));
  assign _zz_2817 = ($signed(data_mid_31_imag) - $signed(data_mid_31_real));
  assign _zz_2818 = fixTo_283_dout;
  assign _zz_2819 = _zz_2820[31 : 0];
  assign _zz_2820 = _zz_2821;
  assign _zz_2821 = ($signed(_zz_2822) >>> _zz_239);
  assign _zz_2822 = _zz_2823;
  assign _zz_2823 = ($signed(_zz_2825) - $signed(_zz_236));
  assign _zz_2824 = ({8'd0,data_mid_27_real} <<< 8);
  assign _zz_2825 = {{8{_zz_2824[23]}}, _zz_2824};
  assign _zz_2826 = fixTo_284_dout;
  assign _zz_2827 = _zz_2828[31 : 0];
  assign _zz_2828 = _zz_2829;
  assign _zz_2829 = ($signed(_zz_2830) >>> _zz_239);
  assign _zz_2830 = _zz_2831;
  assign _zz_2831 = ($signed(_zz_2833) - $signed(_zz_237));
  assign _zz_2832 = ({8'd0,data_mid_27_imag} <<< 8);
  assign _zz_2833 = {{8{_zz_2832[23]}}, _zz_2832};
  assign _zz_2834 = fixTo_285_dout;
  assign _zz_2835 = _zz_2836[31 : 0];
  assign _zz_2836 = _zz_2837;
  assign _zz_2837 = ($signed(_zz_2838) >>> _zz_240);
  assign _zz_2838 = _zz_2839;
  assign _zz_2839 = ($signed(_zz_2841) + $signed(_zz_236));
  assign _zz_2840 = ({8'd0,data_mid_27_real} <<< 8);
  assign _zz_2841 = {{8{_zz_2840[23]}}, _zz_2840};
  assign _zz_2842 = fixTo_286_dout;
  assign _zz_2843 = _zz_2844[31 : 0];
  assign _zz_2844 = _zz_2845;
  assign _zz_2845 = ($signed(_zz_2846) >>> _zz_240);
  assign _zz_2846 = _zz_2847;
  assign _zz_2847 = ($signed(_zz_2849) + $signed(_zz_237));
  assign _zz_2848 = ({8'd0,data_mid_27_imag} <<< 8);
  assign _zz_2849 = {{8{_zz_2848[23]}}, _zz_2848};
  assign _zz_2850 = fixTo_287_dout;
  assign _zz_2851 = ($signed(twiddle_factor_table_7_real) + $signed(twiddle_factor_table_7_imag));
  assign _zz_2852 = ($signed(_zz_243) - $signed(_zz_2853));
  assign _zz_2853 = ($signed(_zz_2854) * $signed(twiddle_factor_table_7_imag));
  assign _zz_2854 = ($signed(data_mid_8_real) + $signed(data_mid_8_imag));
  assign _zz_2855 = fixTo_288_dout;
  assign _zz_2856 = ($signed(_zz_243) + $signed(_zz_2857));
  assign _zz_2857 = ($signed(_zz_2858) * $signed(twiddle_factor_table_7_real));
  assign _zz_2858 = ($signed(data_mid_8_imag) - $signed(data_mid_8_real));
  assign _zz_2859 = fixTo_289_dout;
  assign _zz_2860 = _zz_2861[31 : 0];
  assign _zz_2861 = _zz_2862;
  assign _zz_2862 = ($signed(_zz_2863) >>> _zz_244);
  assign _zz_2863 = _zz_2864;
  assign _zz_2864 = ($signed(_zz_2866) - $signed(_zz_241));
  assign _zz_2865 = ({8'd0,data_mid_0_real} <<< 8);
  assign _zz_2866 = {{8{_zz_2865[23]}}, _zz_2865};
  assign _zz_2867 = fixTo_290_dout;
  assign _zz_2868 = _zz_2869[31 : 0];
  assign _zz_2869 = _zz_2870;
  assign _zz_2870 = ($signed(_zz_2871) >>> _zz_244);
  assign _zz_2871 = _zz_2872;
  assign _zz_2872 = ($signed(_zz_2874) - $signed(_zz_242));
  assign _zz_2873 = ({8'd0,data_mid_0_imag} <<< 8);
  assign _zz_2874 = {{8{_zz_2873[23]}}, _zz_2873};
  assign _zz_2875 = fixTo_291_dout;
  assign _zz_2876 = _zz_2877[31 : 0];
  assign _zz_2877 = _zz_2878;
  assign _zz_2878 = ($signed(_zz_2879) >>> _zz_245);
  assign _zz_2879 = _zz_2880;
  assign _zz_2880 = ($signed(_zz_2882) + $signed(_zz_241));
  assign _zz_2881 = ({8'd0,data_mid_0_real} <<< 8);
  assign _zz_2882 = {{8{_zz_2881[23]}}, _zz_2881};
  assign _zz_2883 = fixTo_292_dout;
  assign _zz_2884 = _zz_2885[31 : 0];
  assign _zz_2885 = _zz_2886;
  assign _zz_2886 = ($signed(_zz_2887) >>> _zz_245);
  assign _zz_2887 = _zz_2888;
  assign _zz_2888 = ($signed(_zz_2890) + $signed(_zz_242));
  assign _zz_2889 = ({8'd0,data_mid_0_imag} <<< 8);
  assign _zz_2890 = {{8{_zz_2889[23]}}, _zz_2889};
  assign _zz_2891 = fixTo_293_dout;
  assign _zz_2892 = ($signed(twiddle_factor_table_8_real) + $signed(twiddle_factor_table_8_imag));
  assign _zz_2893 = ($signed(_zz_248) - $signed(_zz_2894));
  assign _zz_2894 = ($signed(_zz_2895) * $signed(twiddle_factor_table_8_imag));
  assign _zz_2895 = ($signed(data_mid_9_real) + $signed(data_mid_9_imag));
  assign _zz_2896 = fixTo_294_dout;
  assign _zz_2897 = ($signed(_zz_248) + $signed(_zz_2898));
  assign _zz_2898 = ($signed(_zz_2899) * $signed(twiddle_factor_table_8_real));
  assign _zz_2899 = ($signed(data_mid_9_imag) - $signed(data_mid_9_real));
  assign _zz_2900 = fixTo_295_dout;
  assign _zz_2901 = _zz_2902[31 : 0];
  assign _zz_2902 = _zz_2903;
  assign _zz_2903 = ($signed(_zz_2904) >>> _zz_249);
  assign _zz_2904 = _zz_2905;
  assign _zz_2905 = ($signed(_zz_2907) - $signed(_zz_246));
  assign _zz_2906 = ({8'd0,data_mid_1_real} <<< 8);
  assign _zz_2907 = {{8{_zz_2906[23]}}, _zz_2906};
  assign _zz_2908 = fixTo_296_dout;
  assign _zz_2909 = _zz_2910[31 : 0];
  assign _zz_2910 = _zz_2911;
  assign _zz_2911 = ($signed(_zz_2912) >>> _zz_249);
  assign _zz_2912 = _zz_2913;
  assign _zz_2913 = ($signed(_zz_2915) - $signed(_zz_247));
  assign _zz_2914 = ({8'd0,data_mid_1_imag} <<< 8);
  assign _zz_2915 = {{8{_zz_2914[23]}}, _zz_2914};
  assign _zz_2916 = fixTo_297_dout;
  assign _zz_2917 = _zz_2918[31 : 0];
  assign _zz_2918 = _zz_2919;
  assign _zz_2919 = ($signed(_zz_2920) >>> _zz_250);
  assign _zz_2920 = _zz_2921;
  assign _zz_2921 = ($signed(_zz_2923) + $signed(_zz_246));
  assign _zz_2922 = ({8'd0,data_mid_1_real} <<< 8);
  assign _zz_2923 = {{8{_zz_2922[23]}}, _zz_2922};
  assign _zz_2924 = fixTo_298_dout;
  assign _zz_2925 = _zz_2926[31 : 0];
  assign _zz_2926 = _zz_2927;
  assign _zz_2927 = ($signed(_zz_2928) >>> _zz_250);
  assign _zz_2928 = _zz_2929;
  assign _zz_2929 = ($signed(_zz_2931) + $signed(_zz_247));
  assign _zz_2930 = ({8'd0,data_mid_1_imag} <<< 8);
  assign _zz_2931 = {{8{_zz_2930[23]}}, _zz_2930};
  assign _zz_2932 = fixTo_299_dout;
  assign _zz_2933 = ($signed(twiddle_factor_table_9_real) + $signed(twiddle_factor_table_9_imag));
  assign _zz_2934 = ($signed(_zz_253) - $signed(_zz_2935));
  assign _zz_2935 = ($signed(_zz_2936) * $signed(twiddle_factor_table_9_imag));
  assign _zz_2936 = ($signed(data_mid_10_real) + $signed(data_mid_10_imag));
  assign _zz_2937 = fixTo_300_dout;
  assign _zz_2938 = ($signed(_zz_253) + $signed(_zz_2939));
  assign _zz_2939 = ($signed(_zz_2940) * $signed(twiddle_factor_table_9_real));
  assign _zz_2940 = ($signed(data_mid_10_imag) - $signed(data_mid_10_real));
  assign _zz_2941 = fixTo_301_dout;
  assign _zz_2942 = _zz_2943[31 : 0];
  assign _zz_2943 = _zz_2944;
  assign _zz_2944 = ($signed(_zz_2945) >>> _zz_254);
  assign _zz_2945 = _zz_2946;
  assign _zz_2946 = ($signed(_zz_2948) - $signed(_zz_251));
  assign _zz_2947 = ({8'd0,data_mid_2_real} <<< 8);
  assign _zz_2948 = {{8{_zz_2947[23]}}, _zz_2947};
  assign _zz_2949 = fixTo_302_dout;
  assign _zz_2950 = _zz_2951[31 : 0];
  assign _zz_2951 = _zz_2952;
  assign _zz_2952 = ($signed(_zz_2953) >>> _zz_254);
  assign _zz_2953 = _zz_2954;
  assign _zz_2954 = ($signed(_zz_2956) - $signed(_zz_252));
  assign _zz_2955 = ({8'd0,data_mid_2_imag} <<< 8);
  assign _zz_2956 = {{8{_zz_2955[23]}}, _zz_2955};
  assign _zz_2957 = fixTo_303_dout;
  assign _zz_2958 = _zz_2959[31 : 0];
  assign _zz_2959 = _zz_2960;
  assign _zz_2960 = ($signed(_zz_2961) >>> _zz_255);
  assign _zz_2961 = _zz_2962;
  assign _zz_2962 = ($signed(_zz_2964) + $signed(_zz_251));
  assign _zz_2963 = ({8'd0,data_mid_2_real} <<< 8);
  assign _zz_2964 = {{8{_zz_2963[23]}}, _zz_2963};
  assign _zz_2965 = fixTo_304_dout;
  assign _zz_2966 = _zz_2967[31 : 0];
  assign _zz_2967 = _zz_2968;
  assign _zz_2968 = ($signed(_zz_2969) >>> _zz_255);
  assign _zz_2969 = _zz_2970;
  assign _zz_2970 = ($signed(_zz_2972) + $signed(_zz_252));
  assign _zz_2971 = ({8'd0,data_mid_2_imag} <<< 8);
  assign _zz_2972 = {{8{_zz_2971[23]}}, _zz_2971};
  assign _zz_2973 = fixTo_305_dout;
  assign _zz_2974 = ($signed(twiddle_factor_table_10_real) + $signed(twiddle_factor_table_10_imag));
  assign _zz_2975 = ($signed(_zz_258) - $signed(_zz_2976));
  assign _zz_2976 = ($signed(_zz_2977) * $signed(twiddle_factor_table_10_imag));
  assign _zz_2977 = ($signed(data_mid_11_real) + $signed(data_mid_11_imag));
  assign _zz_2978 = fixTo_306_dout;
  assign _zz_2979 = ($signed(_zz_258) + $signed(_zz_2980));
  assign _zz_2980 = ($signed(_zz_2981) * $signed(twiddle_factor_table_10_real));
  assign _zz_2981 = ($signed(data_mid_11_imag) - $signed(data_mid_11_real));
  assign _zz_2982 = fixTo_307_dout;
  assign _zz_2983 = _zz_2984[31 : 0];
  assign _zz_2984 = _zz_2985;
  assign _zz_2985 = ($signed(_zz_2986) >>> _zz_259);
  assign _zz_2986 = _zz_2987;
  assign _zz_2987 = ($signed(_zz_2989) - $signed(_zz_256));
  assign _zz_2988 = ({8'd0,data_mid_3_real} <<< 8);
  assign _zz_2989 = {{8{_zz_2988[23]}}, _zz_2988};
  assign _zz_2990 = fixTo_308_dout;
  assign _zz_2991 = _zz_2992[31 : 0];
  assign _zz_2992 = _zz_2993;
  assign _zz_2993 = ($signed(_zz_2994) >>> _zz_259);
  assign _zz_2994 = _zz_2995;
  assign _zz_2995 = ($signed(_zz_2997) - $signed(_zz_257));
  assign _zz_2996 = ({8'd0,data_mid_3_imag} <<< 8);
  assign _zz_2997 = {{8{_zz_2996[23]}}, _zz_2996};
  assign _zz_2998 = fixTo_309_dout;
  assign _zz_2999 = _zz_3000[31 : 0];
  assign _zz_3000 = _zz_3001;
  assign _zz_3001 = ($signed(_zz_3002) >>> _zz_260);
  assign _zz_3002 = _zz_3003;
  assign _zz_3003 = ($signed(_zz_3005) + $signed(_zz_256));
  assign _zz_3004 = ({8'd0,data_mid_3_real} <<< 8);
  assign _zz_3005 = {{8{_zz_3004[23]}}, _zz_3004};
  assign _zz_3006 = fixTo_310_dout;
  assign _zz_3007 = _zz_3008[31 : 0];
  assign _zz_3008 = _zz_3009;
  assign _zz_3009 = ($signed(_zz_3010) >>> _zz_260);
  assign _zz_3010 = _zz_3011;
  assign _zz_3011 = ($signed(_zz_3013) + $signed(_zz_257));
  assign _zz_3012 = ({8'd0,data_mid_3_imag} <<< 8);
  assign _zz_3013 = {{8{_zz_3012[23]}}, _zz_3012};
  assign _zz_3014 = fixTo_311_dout;
  assign _zz_3015 = ($signed(twiddle_factor_table_11_real) + $signed(twiddle_factor_table_11_imag));
  assign _zz_3016 = ($signed(_zz_263) - $signed(_zz_3017));
  assign _zz_3017 = ($signed(_zz_3018) * $signed(twiddle_factor_table_11_imag));
  assign _zz_3018 = ($signed(data_mid_12_real) + $signed(data_mid_12_imag));
  assign _zz_3019 = fixTo_312_dout;
  assign _zz_3020 = ($signed(_zz_263) + $signed(_zz_3021));
  assign _zz_3021 = ($signed(_zz_3022) * $signed(twiddle_factor_table_11_real));
  assign _zz_3022 = ($signed(data_mid_12_imag) - $signed(data_mid_12_real));
  assign _zz_3023 = fixTo_313_dout;
  assign _zz_3024 = _zz_3025[31 : 0];
  assign _zz_3025 = _zz_3026;
  assign _zz_3026 = ($signed(_zz_3027) >>> _zz_264);
  assign _zz_3027 = _zz_3028;
  assign _zz_3028 = ($signed(_zz_3030) - $signed(_zz_261));
  assign _zz_3029 = ({8'd0,data_mid_4_real} <<< 8);
  assign _zz_3030 = {{8{_zz_3029[23]}}, _zz_3029};
  assign _zz_3031 = fixTo_314_dout;
  assign _zz_3032 = _zz_3033[31 : 0];
  assign _zz_3033 = _zz_3034;
  assign _zz_3034 = ($signed(_zz_3035) >>> _zz_264);
  assign _zz_3035 = _zz_3036;
  assign _zz_3036 = ($signed(_zz_3038) - $signed(_zz_262));
  assign _zz_3037 = ({8'd0,data_mid_4_imag} <<< 8);
  assign _zz_3038 = {{8{_zz_3037[23]}}, _zz_3037};
  assign _zz_3039 = fixTo_315_dout;
  assign _zz_3040 = _zz_3041[31 : 0];
  assign _zz_3041 = _zz_3042;
  assign _zz_3042 = ($signed(_zz_3043) >>> _zz_265);
  assign _zz_3043 = _zz_3044;
  assign _zz_3044 = ($signed(_zz_3046) + $signed(_zz_261));
  assign _zz_3045 = ({8'd0,data_mid_4_real} <<< 8);
  assign _zz_3046 = {{8{_zz_3045[23]}}, _zz_3045};
  assign _zz_3047 = fixTo_316_dout;
  assign _zz_3048 = _zz_3049[31 : 0];
  assign _zz_3049 = _zz_3050;
  assign _zz_3050 = ($signed(_zz_3051) >>> _zz_265);
  assign _zz_3051 = _zz_3052;
  assign _zz_3052 = ($signed(_zz_3054) + $signed(_zz_262));
  assign _zz_3053 = ({8'd0,data_mid_4_imag} <<< 8);
  assign _zz_3054 = {{8{_zz_3053[23]}}, _zz_3053};
  assign _zz_3055 = fixTo_317_dout;
  assign _zz_3056 = ($signed(twiddle_factor_table_12_real) + $signed(twiddle_factor_table_12_imag));
  assign _zz_3057 = ($signed(_zz_268) - $signed(_zz_3058));
  assign _zz_3058 = ($signed(_zz_3059) * $signed(twiddle_factor_table_12_imag));
  assign _zz_3059 = ($signed(data_mid_13_real) + $signed(data_mid_13_imag));
  assign _zz_3060 = fixTo_318_dout;
  assign _zz_3061 = ($signed(_zz_268) + $signed(_zz_3062));
  assign _zz_3062 = ($signed(_zz_3063) * $signed(twiddle_factor_table_12_real));
  assign _zz_3063 = ($signed(data_mid_13_imag) - $signed(data_mid_13_real));
  assign _zz_3064 = fixTo_319_dout;
  assign _zz_3065 = _zz_3066[31 : 0];
  assign _zz_3066 = _zz_3067;
  assign _zz_3067 = ($signed(_zz_3068) >>> _zz_269);
  assign _zz_3068 = _zz_3069;
  assign _zz_3069 = ($signed(_zz_3071) - $signed(_zz_266));
  assign _zz_3070 = ({8'd0,data_mid_5_real} <<< 8);
  assign _zz_3071 = {{8{_zz_3070[23]}}, _zz_3070};
  assign _zz_3072 = fixTo_320_dout;
  assign _zz_3073 = _zz_3074[31 : 0];
  assign _zz_3074 = _zz_3075;
  assign _zz_3075 = ($signed(_zz_3076) >>> _zz_269);
  assign _zz_3076 = _zz_3077;
  assign _zz_3077 = ($signed(_zz_3079) - $signed(_zz_267));
  assign _zz_3078 = ({8'd0,data_mid_5_imag} <<< 8);
  assign _zz_3079 = {{8{_zz_3078[23]}}, _zz_3078};
  assign _zz_3080 = fixTo_321_dout;
  assign _zz_3081 = _zz_3082[31 : 0];
  assign _zz_3082 = _zz_3083;
  assign _zz_3083 = ($signed(_zz_3084) >>> _zz_270);
  assign _zz_3084 = _zz_3085;
  assign _zz_3085 = ($signed(_zz_3087) + $signed(_zz_266));
  assign _zz_3086 = ({8'd0,data_mid_5_real} <<< 8);
  assign _zz_3087 = {{8{_zz_3086[23]}}, _zz_3086};
  assign _zz_3088 = fixTo_322_dout;
  assign _zz_3089 = _zz_3090[31 : 0];
  assign _zz_3090 = _zz_3091;
  assign _zz_3091 = ($signed(_zz_3092) >>> _zz_270);
  assign _zz_3092 = _zz_3093;
  assign _zz_3093 = ($signed(_zz_3095) + $signed(_zz_267));
  assign _zz_3094 = ({8'd0,data_mid_5_imag} <<< 8);
  assign _zz_3095 = {{8{_zz_3094[23]}}, _zz_3094};
  assign _zz_3096 = fixTo_323_dout;
  assign _zz_3097 = ($signed(twiddle_factor_table_13_real) + $signed(twiddle_factor_table_13_imag));
  assign _zz_3098 = ($signed(_zz_273) - $signed(_zz_3099));
  assign _zz_3099 = ($signed(_zz_3100) * $signed(twiddle_factor_table_13_imag));
  assign _zz_3100 = ($signed(data_mid_14_real) + $signed(data_mid_14_imag));
  assign _zz_3101 = fixTo_324_dout;
  assign _zz_3102 = ($signed(_zz_273) + $signed(_zz_3103));
  assign _zz_3103 = ($signed(_zz_3104) * $signed(twiddle_factor_table_13_real));
  assign _zz_3104 = ($signed(data_mid_14_imag) - $signed(data_mid_14_real));
  assign _zz_3105 = fixTo_325_dout;
  assign _zz_3106 = _zz_3107[31 : 0];
  assign _zz_3107 = _zz_3108;
  assign _zz_3108 = ($signed(_zz_3109) >>> _zz_274);
  assign _zz_3109 = _zz_3110;
  assign _zz_3110 = ($signed(_zz_3112) - $signed(_zz_271));
  assign _zz_3111 = ({8'd0,data_mid_6_real} <<< 8);
  assign _zz_3112 = {{8{_zz_3111[23]}}, _zz_3111};
  assign _zz_3113 = fixTo_326_dout;
  assign _zz_3114 = _zz_3115[31 : 0];
  assign _zz_3115 = _zz_3116;
  assign _zz_3116 = ($signed(_zz_3117) >>> _zz_274);
  assign _zz_3117 = _zz_3118;
  assign _zz_3118 = ($signed(_zz_3120) - $signed(_zz_272));
  assign _zz_3119 = ({8'd0,data_mid_6_imag} <<< 8);
  assign _zz_3120 = {{8{_zz_3119[23]}}, _zz_3119};
  assign _zz_3121 = fixTo_327_dout;
  assign _zz_3122 = _zz_3123[31 : 0];
  assign _zz_3123 = _zz_3124;
  assign _zz_3124 = ($signed(_zz_3125) >>> _zz_275);
  assign _zz_3125 = _zz_3126;
  assign _zz_3126 = ($signed(_zz_3128) + $signed(_zz_271));
  assign _zz_3127 = ({8'd0,data_mid_6_real} <<< 8);
  assign _zz_3128 = {{8{_zz_3127[23]}}, _zz_3127};
  assign _zz_3129 = fixTo_328_dout;
  assign _zz_3130 = _zz_3131[31 : 0];
  assign _zz_3131 = _zz_3132;
  assign _zz_3132 = ($signed(_zz_3133) >>> _zz_275);
  assign _zz_3133 = _zz_3134;
  assign _zz_3134 = ($signed(_zz_3136) + $signed(_zz_272));
  assign _zz_3135 = ({8'd0,data_mid_6_imag} <<< 8);
  assign _zz_3136 = {{8{_zz_3135[23]}}, _zz_3135};
  assign _zz_3137 = fixTo_329_dout;
  assign _zz_3138 = ($signed(twiddle_factor_table_14_real) + $signed(twiddle_factor_table_14_imag));
  assign _zz_3139 = ($signed(_zz_278) - $signed(_zz_3140));
  assign _zz_3140 = ($signed(_zz_3141) * $signed(twiddle_factor_table_14_imag));
  assign _zz_3141 = ($signed(data_mid_15_real) + $signed(data_mid_15_imag));
  assign _zz_3142 = fixTo_330_dout;
  assign _zz_3143 = ($signed(_zz_278) + $signed(_zz_3144));
  assign _zz_3144 = ($signed(_zz_3145) * $signed(twiddle_factor_table_14_real));
  assign _zz_3145 = ($signed(data_mid_15_imag) - $signed(data_mid_15_real));
  assign _zz_3146 = fixTo_331_dout;
  assign _zz_3147 = _zz_3148[31 : 0];
  assign _zz_3148 = _zz_3149;
  assign _zz_3149 = ($signed(_zz_3150) >>> _zz_279);
  assign _zz_3150 = _zz_3151;
  assign _zz_3151 = ($signed(_zz_3153) - $signed(_zz_276));
  assign _zz_3152 = ({8'd0,data_mid_7_real} <<< 8);
  assign _zz_3153 = {{8{_zz_3152[23]}}, _zz_3152};
  assign _zz_3154 = fixTo_332_dout;
  assign _zz_3155 = _zz_3156[31 : 0];
  assign _zz_3156 = _zz_3157;
  assign _zz_3157 = ($signed(_zz_3158) >>> _zz_279);
  assign _zz_3158 = _zz_3159;
  assign _zz_3159 = ($signed(_zz_3161) - $signed(_zz_277));
  assign _zz_3160 = ({8'd0,data_mid_7_imag} <<< 8);
  assign _zz_3161 = {{8{_zz_3160[23]}}, _zz_3160};
  assign _zz_3162 = fixTo_333_dout;
  assign _zz_3163 = _zz_3164[31 : 0];
  assign _zz_3164 = _zz_3165;
  assign _zz_3165 = ($signed(_zz_3166) >>> _zz_280);
  assign _zz_3166 = _zz_3167;
  assign _zz_3167 = ($signed(_zz_3169) + $signed(_zz_276));
  assign _zz_3168 = ({8'd0,data_mid_7_real} <<< 8);
  assign _zz_3169 = {{8{_zz_3168[23]}}, _zz_3168};
  assign _zz_3170 = fixTo_334_dout;
  assign _zz_3171 = _zz_3172[31 : 0];
  assign _zz_3172 = _zz_3173;
  assign _zz_3173 = ($signed(_zz_3174) >>> _zz_280);
  assign _zz_3174 = _zz_3175;
  assign _zz_3175 = ($signed(_zz_3177) + $signed(_zz_277));
  assign _zz_3176 = ({8'd0,data_mid_7_imag} <<< 8);
  assign _zz_3177 = {{8{_zz_3176[23]}}, _zz_3176};
  assign _zz_3178 = fixTo_335_dout;
  assign _zz_3179 = ($signed(twiddle_factor_table_7_real) + $signed(twiddle_factor_table_7_imag));
  assign _zz_3180 = ($signed(_zz_283) - $signed(_zz_3181));
  assign _zz_3181 = ($signed(_zz_3182) * $signed(twiddle_factor_table_7_imag));
  assign _zz_3182 = ($signed(data_mid_24_real) + $signed(data_mid_24_imag));
  assign _zz_3183 = fixTo_336_dout;
  assign _zz_3184 = ($signed(_zz_283) + $signed(_zz_3185));
  assign _zz_3185 = ($signed(_zz_3186) * $signed(twiddle_factor_table_7_real));
  assign _zz_3186 = ($signed(data_mid_24_imag) - $signed(data_mid_24_real));
  assign _zz_3187 = fixTo_337_dout;
  assign _zz_3188 = _zz_3189[31 : 0];
  assign _zz_3189 = _zz_3190;
  assign _zz_3190 = ($signed(_zz_3191) >>> _zz_284);
  assign _zz_3191 = _zz_3192;
  assign _zz_3192 = ($signed(_zz_3194) - $signed(_zz_281));
  assign _zz_3193 = ({8'd0,data_mid_16_real} <<< 8);
  assign _zz_3194 = {{8{_zz_3193[23]}}, _zz_3193};
  assign _zz_3195 = fixTo_338_dout;
  assign _zz_3196 = _zz_3197[31 : 0];
  assign _zz_3197 = _zz_3198;
  assign _zz_3198 = ($signed(_zz_3199) >>> _zz_284);
  assign _zz_3199 = _zz_3200;
  assign _zz_3200 = ($signed(_zz_3202) - $signed(_zz_282));
  assign _zz_3201 = ({8'd0,data_mid_16_imag} <<< 8);
  assign _zz_3202 = {{8{_zz_3201[23]}}, _zz_3201};
  assign _zz_3203 = fixTo_339_dout;
  assign _zz_3204 = _zz_3205[31 : 0];
  assign _zz_3205 = _zz_3206;
  assign _zz_3206 = ($signed(_zz_3207) >>> _zz_285);
  assign _zz_3207 = _zz_3208;
  assign _zz_3208 = ($signed(_zz_3210) + $signed(_zz_281));
  assign _zz_3209 = ({8'd0,data_mid_16_real} <<< 8);
  assign _zz_3210 = {{8{_zz_3209[23]}}, _zz_3209};
  assign _zz_3211 = fixTo_340_dout;
  assign _zz_3212 = _zz_3213[31 : 0];
  assign _zz_3213 = _zz_3214;
  assign _zz_3214 = ($signed(_zz_3215) >>> _zz_285);
  assign _zz_3215 = _zz_3216;
  assign _zz_3216 = ($signed(_zz_3218) + $signed(_zz_282));
  assign _zz_3217 = ({8'd0,data_mid_16_imag} <<< 8);
  assign _zz_3218 = {{8{_zz_3217[23]}}, _zz_3217};
  assign _zz_3219 = fixTo_341_dout;
  assign _zz_3220 = ($signed(twiddle_factor_table_8_real) + $signed(twiddle_factor_table_8_imag));
  assign _zz_3221 = ($signed(_zz_288) - $signed(_zz_3222));
  assign _zz_3222 = ($signed(_zz_3223) * $signed(twiddle_factor_table_8_imag));
  assign _zz_3223 = ($signed(data_mid_25_real) + $signed(data_mid_25_imag));
  assign _zz_3224 = fixTo_342_dout;
  assign _zz_3225 = ($signed(_zz_288) + $signed(_zz_3226));
  assign _zz_3226 = ($signed(_zz_3227) * $signed(twiddle_factor_table_8_real));
  assign _zz_3227 = ($signed(data_mid_25_imag) - $signed(data_mid_25_real));
  assign _zz_3228 = fixTo_343_dout;
  assign _zz_3229 = _zz_3230[31 : 0];
  assign _zz_3230 = _zz_3231;
  assign _zz_3231 = ($signed(_zz_3232) >>> _zz_289);
  assign _zz_3232 = _zz_3233;
  assign _zz_3233 = ($signed(_zz_3235) - $signed(_zz_286));
  assign _zz_3234 = ({8'd0,data_mid_17_real} <<< 8);
  assign _zz_3235 = {{8{_zz_3234[23]}}, _zz_3234};
  assign _zz_3236 = fixTo_344_dout;
  assign _zz_3237 = _zz_3238[31 : 0];
  assign _zz_3238 = _zz_3239;
  assign _zz_3239 = ($signed(_zz_3240) >>> _zz_289);
  assign _zz_3240 = _zz_3241;
  assign _zz_3241 = ($signed(_zz_3243) - $signed(_zz_287));
  assign _zz_3242 = ({8'd0,data_mid_17_imag} <<< 8);
  assign _zz_3243 = {{8{_zz_3242[23]}}, _zz_3242};
  assign _zz_3244 = fixTo_345_dout;
  assign _zz_3245 = _zz_3246[31 : 0];
  assign _zz_3246 = _zz_3247;
  assign _zz_3247 = ($signed(_zz_3248) >>> _zz_290);
  assign _zz_3248 = _zz_3249;
  assign _zz_3249 = ($signed(_zz_3251) + $signed(_zz_286));
  assign _zz_3250 = ({8'd0,data_mid_17_real} <<< 8);
  assign _zz_3251 = {{8{_zz_3250[23]}}, _zz_3250};
  assign _zz_3252 = fixTo_346_dout;
  assign _zz_3253 = _zz_3254[31 : 0];
  assign _zz_3254 = _zz_3255;
  assign _zz_3255 = ($signed(_zz_3256) >>> _zz_290);
  assign _zz_3256 = _zz_3257;
  assign _zz_3257 = ($signed(_zz_3259) + $signed(_zz_287));
  assign _zz_3258 = ({8'd0,data_mid_17_imag} <<< 8);
  assign _zz_3259 = {{8{_zz_3258[23]}}, _zz_3258};
  assign _zz_3260 = fixTo_347_dout;
  assign _zz_3261 = ($signed(twiddle_factor_table_9_real) + $signed(twiddle_factor_table_9_imag));
  assign _zz_3262 = ($signed(_zz_293) - $signed(_zz_3263));
  assign _zz_3263 = ($signed(_zz_3264) * $signed(twiddle_factor_table_9_imag));
  assign _zz_3264 = ($signed(data_mid_26_real) + $signed(data_mid_26_imag));
  assign _zz_3265 = fixTo_348_dout;
  assign _zz_3266 = ($signed(_zz_293) + $signed(_zz_3267));
  assign _zz_3267 = ($signed(_zz_3268) * $signed(twiddle_factor_table_9_real));
  assign _zz_3268 = ($signed(data_mid_26_imag) - $signed(data_mid_26_real));
  assign _zz_3269 = fixTo_349_dout;
  assign _zz_3270 = _zz_3271[31 : 0];
  assign _zz_3271 = _zz_3272;
  assign _zz_3272 = ($signed(_zz_3273) >>> _zz_294);
  assign _zz_3273 = _zz_3274;
  assign _zz_3274 = ($signed(_zz_3276) - $signed(_zz_291));
  assign _zz_3275 = ({8'd0,data_mid_18_real} <<< 8);
  assign _zz_3276 = {{8{_zz_3275[23]}}, _zz_3275};
  assign _zz_3277 = fixTo_350_dout;
  assign _zz_3278 = _zz_3279[31 : 0];
  assign _zz_3279 = _zz_3280;
  assign _zz_3280 = ($signed(_zz_3281) >>> _zz_294);
  assign _zz_3281 = _zz_3282;
  assign _zz_3282 = ($signed(_zz_3284) - $signed(_zz_292));
  assign _zz_3283 = ({8'd0,data_mid_18_imag} <<< 8);
  assign _zz_3284 = {{8{_zz_3283[23]}}, _zz_3283};
  assign _zz_3285 = fixTo_351_dout;
  assign _zz_3286 = _zz_3287[31 : 0];
  assign _zz_3287 = _zz_3288;
  assign _zz_3288 = ($signed(_zz_3289) >>> _zz_295);
  assign _zz_3289 = _zz_3290;
  assign _zz_3290 = ($signed(_zz_3292) + $signed(_zz_291));
  assign _zz_3291 = ({8'd0,data_mid_18_real} <<< 8);
  assign _zz_3292 = {{8{_zz_3291[23]}}, _zz_3291};
  assign _zz_3293 = fixTo_352_dout;
  assign _zz_3294 = _zz_3295[31 : 0];
  assign _zz_3295 = _zz_3296;
  assign _zz_3296 = ($signed(_zz_3297) >>> _zz_295);
  assign _zz_3297 = _zz_3298;
  assign _zz_3298 = ($signed(_zz_3300) + $signed(_zz_292));
  assign _zz_3299 = ({8'd0,data_mid_18_imag} <<< 8);
  assign _zz_3300 = {{8{_zz_3299[23]}}, _zz_3299};
  assign _zz_3301 = fixTo_353_dout;
  assign _zz_3302 = ($signed(twiddle_factor_table_10_real) + $signed(twiddle_factor_table_10_imag));
  assign _zz_3303 = ($signed(_zz_298) - $signed(_zz_3304));
  assign _zz_3304 = ($signed(_zz_3305) * $signed(twiddle_factor_table_10_imag));
  assign _zz_3305 = ($signed(data_mid_27_real) + $signed(data_mid_27_imag));
  assign _zz_3306 = fixTo_354_dout;
  assign _zz_3307 = ($signed(_zz_298) + $signed(_zz_3308));
  assign _zz_3308 = ($signed(_zz_3309) * $signed(twiddle_factor_table_10_real));
  assign _zz_3309 = ($signed(data_mid_27_imag) - $signed(data_mid_27_real));
  assign _zz_3310 = fixTo_355_dout;
  assign _zz_3311 = _zz_3312[31 : 0];
  assign _zz_3312 = _zz_3313;
  assign _zz_3313 = ($signed(_zz_3314) >>> _zz_299);
  assign _zz_3314 = _zz_3315;
  assign _zz_3315 = ($signed(_zz_3317) - $signed(_zz_296));
  assign _zz_3316 = ({8'd0,data_mid_19_real} <<< 8);
  assign _zz_3317 = {{8{_zz_3316[23]}}, _zz_3316};
  assign _zz_3318 = fixTo_356_dout;
  assign _zz_3319 = _zz_3320[31 : 0];
  assign _zz_3320 = _zz_3321;
  assign _zz_3321 = ($signed(_zz_3322) >>> _zz_299);
  assign _zz_3322 = _zz_3323;
  assign _zz_3323 = ($signed(_zz_3325) - $signed(_zz_297));
  assign _zz_3324 = ({8'd0,data_mid_19_imag} <<< 8);
  assign _zz_3325 = {{8{_zz_3324[23]}}, _zz_3324};
  assign _zz_3326 = fixTo_357_dout;
  assign _zz_3327 = _zz_3328[31 : 0];
  assign _zz_3328 = _zz_3329;
  assign _zz_3329 = ($signed(_zz_3330) >>> _zz_300);
  assign _zz_3330 = _zz_3331;
  assign _zz_3331 = ($signed(_zz_3333) + $signed(_zz_296));
  assign _zz_3332 = ({8'd0,data_mid_19_real} <<< 8);
  assign _zz_3333 = {{8{_zz_3332[23]}}, _zz_3332};
  assign _zz_3334 = fixTo_358_dout;
  assign _zz_3335 = _zz_3336[31 : 0];
  assign _zz_3336 = _zz_3337;
  assign _zz_3337 = ($signed(_zz_3338) >>> _zz_300);
  assign _zz_3338 = _zz_3339;
  assign _zz_3339 = ($signed(_zz_3341) + $signed(_zz_297));
  assign _zz_3340 = ({8'd0,data_mid_19_imag} <<< 8);
  assign _zz_3341 = {{8{_zz_3340[23]}}, _zz_3340};
  assign _zz_3342 = fixTo_359_dout;
  assign _zz_3343 = ($signed(twiddle_factor_table_11_real) + $signed(twiddle_factor_table_11_imag));
  assign _zz_3344 = ($signed(_zz_303) - $signed(_zz_3345));
  assign _zz_3345 = ($signed(_zz_3346) * $signed(twiddle_factor_table_11_imag));
  assign _zz_3346 = ($signed(data_mid_28_real) + $signed(data_mid_28_imag));
  assign _zz_3347 = fixTo_360_dout;
  assign _zz_3348 = ($signed(_zz_303) + $signed(_zz_3349));
  assign _zz_3349 = ($signed(_zz_3350) * $signed(twiddle_factor_table_11_real));
  assign _zz_3350 = ($signed(data_mid_28_imag) - $signed(data_mid_28_real));
  assign _zz_3351 = fixTo_361_dout;
  assign _zz_3352 = _zz_3353[31 : 0];
  assign _zz_3353 = _zz_3354;
  assign _zz_3354 = ($signed(_zz_3355) >>> _zz_304);
  assign _zz_3355 = _zz_3356;
  assign _zz_3356 = ($signed(_zz_3358) - $signed(_zz_301));
  assign _zz_3357 = ({8'd0,data_mid_20_real} <<< 8);
  assign _zz_3358 = {{8{_zz_3357[23]}}, _zz_3357};
  assign _zz_3359 = fixTo_362_dout;
  assign _zz_3360 = _zz_3361[31 : 0];
  assign _zz_3361 = _zz_3362;
  assign _zz_3362 = ($signed(_zz_3363) >>> _zz_304);
  assign _zz_3363 = _zz_3364;
  assign _zz_3364 = ($signed(_zz_3366) - $signed(_zz_302));
  assign _zz_3365 = ({8'd0,data_mid_20_imag} <<< 8);
  assign _zz_3366 = {{8{_zz_3365[23]}}, _zz_3365};
  assign _zz_3367 = fixTo_363_dout;
  assign _zz_3368 = _zz_3369[31 : 0];
  assign _zz_3369 = _zz_3370;
  assign _zz_3370 = ($signed(_zz_3371) >>> _zz_305);
  assign _zz_3371 = _zz_3372;
  assign _zz_3372 = ($signed(_zz_3374) + $signed(_zz_301));
  assign _zz_3373 = ({8'd0,data_mid_20_real} <<< 8);
  assign _zz_3374 = {{8{_zz_3373[23]}}, _zz_3373};
  assign _zz_3375 = fixTo_364_dout;
  assign _zz_3376 = _zz_3377[31 : 0];
  assign _zz_3377 = _zz_3378;
  assign _zz_3378 = ($signed(_zz_3379) >>> _zz_305);
  assign _zz_3379 = _zz_3380;
  assign _zz_3380 = ($signed(_zz_3382) + $signed(_zz_302));
  assign _zz_3381 = ({8'd0,data_mid_20_imag} <<< 8);
  assign _zz_3382 = {{8{_zz_3381[23]}}, _zz_3381};
  assign _zz_3383 = fixTo_365_dout;
  assign _zz_3384 = ($signed(twiddle_factor_table_12_real) + $signed(twiddle_factor_table_12_imag));
  assign _zz_3385 = ($signed(_zz_308) - $signed(_zz_3386));
  assign _zz_3386 = ($signed(_zz_3387) * $signed(twiddle_factor_table_12_imag));
  assign _zz_3387 = ($signed(data_mid_29_real) + $signed(data_mid_29_imag));
  assign _zz_3388 = fixTo_366_dout;
  assign _zz_3389 = ($signed(_zz_308) + $signed(_zz_3390));
  assign _zz_3390 = ($signed(_zz_3391) * $signed(twiddle_factor_table_12_real));
  assign _zz_3391 = ($signed(data_mid_29_imag) - $signed(data_mid_29_real));
  assign _zz_3392 = fixTo_367_dout;
  assign _zz_3393 = _zz_3394[31 : 0];
  assign _zz_3394 = _zz_3395;
  assign _zz_3395 = ($signed(_zz_3396) >>> _zz_309);
  assign _zz_3396 = _zz_3397;
  assign _zz_3397 = ($signed(_zz_3399) - $signed(_zz_306));
  assign _zz_3398 = ({8'd0,data_mid_21_real} <<< 8);
  assign _zz_3399 = {{8{_zz_3398[23]}}, _zz_3398};
  assign _zz_3400 = fixTo_368_dout;
  assign _zz_3401 = _zz_3402[31 : 0];
  assign _zz_3402 = _zz_3403;
  assign _zz_3403 = ($signed(_zz_3404) >>> _zz_309);
  assign _zz_3404 = _zz_3405;
  assign _zz_3405 = ($signed(_zz_3407) - $signed(_zz_307));
  assign _zz_3406 = ({8'd0,data_mid_21_imag} <<< 8);
  assign _zz_3407 = {{8{_zz_3406[23]}}, _zz_3406};
  assign _zz_3408 = fixTo_369_dout;
  assign _zz_3409 = _zz_3410[31 : 0];
  assign _zz_3410 = _zz_3411;
  assign _zz_3411 = ($signed(_zz_3412) >>> _zz_310);
  assign _zz_3412 = _zz_3413;
  assign _zz_3413 = ($signed(_zz_3415) + $signed(_zz_306));
  assign _zz_3414 = ({8'd0,data_mid_21_real} <<< 8);
  assign _zz_3415 = {{8{_zz_3414[23]}}, _zz_3414};
  assign _zz_3416 = fixTo_370_dout;
  assign _zz_3417 = _zz_3418[31 : 0];
  assign _zz_3418 = _zz_3419;
  assign _zz_3419 = ($signed(_zz_3420) >>> _zz_310);
  assign _zz_3420 = _zz_3421;
  assign _zz_3421 = ($signed(_zz_3423) + $signed(_zz_307));
  assign _zz_3422 = ({8'd0,data_mid_21_imag} <<< 8);
  assign _zz_3423 = {{8{_zz_3422[23]}}, _zz_3422};
  assign _zz_3424 = fixTo_371_dout;
  assign _zz_3425 = ($signed(twiddle_factor_table_13_real) + $signed(twiddle_factor_table_13_imag));
  assign _zz_3426 = ($signed(_zz_313) - $signed(_zz_3427));
  assign _zz_3427 = ($signed(_zz_3428) * $signed(twiddle_factor_table_13_imag));
  assign _zz_3428 = ($signed(data_mid_30_real) + $signed(data_mid_30_imag));
  assign _zz_3429 = fixTo_372_dout;
  assign _zz_3430 = ($signed(_zz_313) + $signed(_zz_3431));
  assign _zz_3431 = ($signed(_zz_3432) * $signed(twiddle_factor_table_13_real));
  assign _zz_3432 = ($signed(data_mid_30_imag) - $signed(data_mid_30_real));
  assign _zz_3433 = fixTo_373_dout;
  assign _zz_3434 = _zz_3435[31 : 0];
  assign _zz_3435 = _zz_3436;
  assign _zz_3436 = ($signed(_zz_3437) >>> _zz_314);
  assign _zz_3437 = _zz_3438;
  assign _zz_3438 = ($signed(_zz_3440) - $signed(_zz_311));
  assign _zz_3439 = ({8'd0,data_mid_22_real} <<< 8);
  assign _zz_3440 = {{8{_zz_3439[23]}}, _zz_3439};
  assign _zz_3441 = fixTo_374_dout;
  assign _zz_3442 = _zz_3443[31 : 0];
  assign _zz_3443 = _zz_3444;
  assign _zz_3444 = ($signed(_zz_3445) >>> _zz_314);
  assign _zz_3445 = _zz_3446;
  assign _zz_3446 = ($signed(_zz_3448) - $signed(_zz_312));
  assign _zz_3447 = ({8'd0,data_mid_22_imag} <<< 8);
  assign _zz_3448 = {{8{_zz_3447[23]}}, _zz_3447};
  assign _zz_3449 = fixTo_375_dout;
  assign _zz_3450 = _zz_3451[31 : 0];
  assign _zz_3451 = _zz_3452;
  assign _zz_3452 = ($signed(_zz_3453) >>> _zz_315);
  assign _zz_3453 = _zz_3454;
  assign _zz_3454 = ($signed(_zz_3456) + $signed(_zz_311));
  assign _zz_3455 = ({8'd0,data_mid_22_real} <<< 8);
  assign _zz_3456 = {{8{_zz_3455[23]}}, _zz_3455};
  assign _zz_3457 = fixTo_376_dout;
  assign _zz_3458 = _zz_3459[31 : 0];
  assign _zz_3459 = _zz_3460;
  assign _zz_3460 = ($signed(_zz_3461) >>> _zz_315);
  assign _zz_3461 = _zz_3462;
  assign _zz_3462 = ($signed(_zz_3464) + $signed(_zz_312));
  assign _zz_3463 = ({8'd0,data_mid_22_imag} <<< 8);
  assign _zz_3464 = {{8{_zz_3463[23]}}, _zz_3463};
  assign _zz_3465 = fixTo_377_dout;
  assign _zz_3466 = ($signed(twiddle_factor_table_14_real) + $signed(twiddle_factor_table_14_imag));
  assign _zz_3467 = ($signed(_zz_318) - $signed(_zz_3468));
  assign _zz_3468 = ($signed(_zz_3469) * $signed(twiddle_factor_table_14_imag));
  assign _zz_3469 = ($signed(data_mid_31_real) + $signed(data_mid_31_imag));
  assign _zz_3470 = fixTo_378_dout;
  assign _zz_3471 = ($signed(_zz_318) + $signed(_zz_3472));
  assign _zz_3472 = ($signed(_zz_3473) * $signed(twiddle_factor_table_14_real));
  assign _zz_3473 = ($signed(data_mid_31_imag) - $signed(data_mid_31_real));
  assign _zz_3474 = fixTo_379_dout;
  assign _zz_3475 = _zz_3476[31 : 0];
  assign _zz_3476 = _zz_3477;
  assign _zz_3477 = ($signed(_zz_3478) >>> _zz_319);
  assign _zz_3478 = _zz_3479;
  assign _zz_3479 = ($signed(_zz_3481) - $signed(_zz_316));
  assign _zz_3480 = ({8'd0,data_mid_23_real} <<< 8);
  assign _zz_3481 = {{8{_zz_3480[23]}}, _zz_3480};
  assign _zz_3482 = fixTo_380_dout;
  assign _zz_3483 = _zz_3484[31 : 0];
  assign _zz_3484 = _zz_3485;
  assign _zz_3485 = ($signed(_zz_3486) >>> _zz_319);
  assign _zz_3486 = _zz_3487;
  assign _zz_3487 = ($signed(_zz_3489) - $signed(_zz_317));
  assign _zz_3488 = ({8'd0,data_mid_23_imag} <<< 8);
  assign _zz_3489 = {{8{_zz_3488[23]}}, _zz_3488};
  assign _zz_3490 = fixTo_381_dout;
  assign _zz_3491 = _zz_3492[31 : 0];
  assign _zz_3492 = _zz_3493;
  assign _zz_3493 = ($signed(_zz_3494) >>> _zz_320);
  assign _zz_3494 = _zz_3495;
  assign _zz_3495 = ($signed(_zz_3497) + $signed(_zz_316));
  assign _zz_3496 = ({8'd0,data_mid_23_real} <<< 8);
  assign _zz_3497 = {{8{_zz_3496[23]}}, _zz_3496};
  assign _zz_3498 = fixTo_382_dout;
  assign _zz_3499 = _zz_3500[31 : 0];
  assign _zz_3500 = _zz_3501;
  assign _zz_3501 = ($signed(_zz_3502) >>> _zz_320);
  assign _zz_3502 = _zz_3503;
  assign _zz_3503 = ($signed(_zz_3505) + $signed(_zz_317));
  assign _zz_3504 = ({8'd0,data_mid_23_imag} <<< 8);
  assign _zz_3505 = {{8{_zz_3504[23]}}, _zz_3504};
  assign _zz_3506 = fixTo_383_dout;
  assign _zz_3507 = ($signed(twiddle_factor_table_15_real) + $signed(twiddle_factor_table_15_imag));
  assign _zz_3508 = ($signed(_zz_323) - $signed(_zz_3509));
  assign _zz_3509 = ($signed(_zz_3510) * $signed(twiddle_factor_table_15_imag));
  assign _zz_3510 = ($signed(data_mid_16_real) + $signed(data_mid_16_imag));
  assign _zz_3511 = fixTo_384_dout;
  assign _zz_3512 = ($signed(_zz_323) + $signed(_zz_3513));
  assign _zz_3513 = ($signed(_zz_3514) * $signed(twiddle_factor_table_15_real));
  assign _zz_3514 = ($signed(data_mid_16_imag) - $signed(data_mid_16_real));
  assign _zz_3515 = fixTo_385_dout;
  assign _zz_3516 = _zz_3517[31 : 0];
  assign _zz_3517 = _zz_3518;
  assign _zz_3518 = ($signed(_zz_3519) >>> _zz_324);
  assign _zz_3519 = _zz_3520;
  assign _zz_3520 = ($signed(_zz_3522) - $signed(_zz_321));
  assign _zz_3521 = ({8'd0,data_mid_0_real} <<< 8);
  assign _zz_3522 = {{8{_zz_3521[23]}}, _zz_3521};
  assign _zz_3523 = fixTo_386_dout;
  assign _zz_3524 = _zz_3525[31 : 0];
  assign _zz_3525 = _zz_3526;
  assign _zz_3526 = ($signed(_zz_3527) >>> _zz_324);
  assign _zz_3527 = _zz_3528;
  assign _zz_3528 = ($signed(_zz_3530) - $signed(_zz_322));
  assign _zz_3529 = ({8'd0,data_mid_0_imag} <<< 8);
  assign _zz_3530 = {{8{_zz_3529[23]}}, _zz_3529};
  assign _zz_3531 = fixTo_387_dout;
  assign _zz_3532 = _zz_3533[31 : 0];
  assign _zz_3533 = _zz_3534;
  assign _zz_3534 = ($signed(_zz_3535) >>> _zz_325);
  assign _zz_3535 = _zz_3536;
  assign _zz_3536 = ($signed(_zz_3538) + $signed(_zz_321));
  assign _zz_3537 = ({8'd0,data_mid_0_real} <<< 8);
  assign _zz_3538 = {{8{_zz_3537[23]}}, _zz_3537};
  assign _zz_3539 = fixTo_388_dout;
  assign _zz_3540 = _zz_3541[31 : 0];
  assign _zz_3541 = _zz_3542;
  assign _zz_3542 = ($signed(_zz_3543) >>> _zz_325);
  assign _zz_3543 = _zz_3544;
  assign _zz_3544 = ($signed(_zz_3546) + $signed(_zz_322));
  assign _zz_3545 = ({8'd0,data_mid_0_imag} <<< 8);
  assign _zz_3546 = {{8{_zz_3545[23]}}, _zz_3545};
  assign _zz_3547 = fixTo_389_dout;
  assign _zz_3548 = ($signed(twiddle_factor_table_16_real) + $signed(twiddle_factor_table_16_imag));
  assign _zz_3549 = ($signed(_zz_328) - $signed(_zz_3550));
  assign _zz_3550 = ($signed(_zz_3551) * $signed(twiddle_factor_table_16_imag));
  assign _zz_3551 = ($signed(data_mid_17_real) + $signed(data_mid_17_imag));
  assign _zz_3552 = fixTo_390_dout;
  assign _zz_3553 = ($signed(_zz_328) + $signed(_zz_3554));
  assign _zz_3554 = ($signed(_zz_3555) * $signed(twiddle_factor_table_16_real));
  assign _zz_3555 = ($signed(data_mid_17_imag) - $signed(data_mid_17_real));
  assign _zz_3556 = fixTo_391_dout;
  assign _zz_3557 = _zz_3558[31 : 0];
  assign _zz_3558 = _zz_3559;
  assign _zz_3559 = ($signed(_zz_3560) >>> _zz_329);
  assign _zz_3560 = _zz_3561;
  assign _zz_3561 = ($signed(_zz_3563) - $signed(_zz_326));
  assign _zz_3562 = ({8'd0,data_mid_1_real} <<< 8);
  assign _zz_3563 = {{8{_zz_3562[23]}}, _zz_3562};
  assign _zz_3564 = fixTo_392_dout;
  assign _zz_3565 = _zz_3566[31 : 0];
  assign _zz_3566 = _zz_3567;
  assign _zz_3567 = ($signed(_zz_3568) >>> _zz_329);
  assign _zz_3568 = _zz_3569;
  assign _zz_3569 = ($signed(_zz_3571) - $signed(_zz_327));
  assign _zz_3570 = ({8'd0,data_mid_1_imag} <<< 8);
  assign _zz_3571 = {{8{_zz_3570[23]}}, _zz_3570};
  assign _zz_3572 = fixTo_393_dout;
  assign _zz_3573 = _zz_3574[31 : 0];
  assign _zz_3574 = _zz_3575;
  assign _zz_3575 = ($signed(_zz_3576) >>> _zz_330);
  assign _zz_3576 = _zz_3577;
  assign _zz_3577 = ($signed(_zz_3579) + $signed(_zz_326));
  assign _zz_3578 = ({8'd0,data_mid_1_real} <<< 8);
  assign _zz_3579 = {{8{_zz_3578[23]}}, _zz_3578};
  assign _zz_3580 = fixTo_394_dout;
  assign _zz_3581 = _zz_3582[31 : 0];
  assign _zz_3582 = _zz_3583;
  assign _zz_3583 = ($signed(_zz_3584) >>> _zz_330);
  assign _zz_3584 = _zz_3585;
  assign _zz_3585 = ($signed(_zz_3587) + $signed(_zz_327));
  assign _zz_3586 = ({8'd0,data_mid_1_imag} <<< 8);
  assign _zz_3587 = {{8{_zz_3586[23]}}, _zz_3586};
  assign _zz_3588 = fixTo_395_dout;
  assign _zz_3589 = ($signed(twiddle_factor_table_17_real) + $signed(twiddle_factor_table_17_imag));
  assign _zz_3590 = ($signed(_zz_333) - $signed(_zz_3591));
  assign _zz_3591 = ($signed(_zz_3592) * $signed(twiddle_factor_table_17_imag));
  assign _zz_3592 = ($signed(data_mid_18_real) + $signed(data_mid_18_imag));
  assign _zz_3593 = fixTo_396_dout;
  assign _zz_3594 = ($signed(_zz_333) + $signed(_zz_3595));
  assign _zz_3595 = ($signed(_zz_3596) * $signed(twiddle_factor_table_17_real));
  assign _zz_3596 = ($signed(data_mid_18_imag) - $signed(data_mid_18_real));
  assign _zz_3597 = fixTo_397_dout;
  assign _zz_3598 = _zz_3599[31 : 0];
  assign _zz_3599 = _zz_3600;
  assign _zz_3600 = ($signed(_zz_3601) >>> _zz_334);
  assign _zz_3601 = _zz_3602;
  assign _zz_3602 = ($signed(_zz_3604) - $signed(_zz_331));
  assign _zz_3603 = ({8'd0,data_mid_2_real} <<< 8);
  assign _zz_3604 = {{8{_zz_3603[23]}}, _zz_3603};
  assign _zz_3605 = fixTo_398_dout;
  assign _zz_3606 = _zz_3607[31 : 0];
  assign _zz_3607 = _zz_3608;
  assign _zz_3608 = ($signed(_zz_3609) >>> _zz_334);
  assign _zz_3609 = _zz_3610;
  assign _zz_3610 = ($signed(_zz_3612) - $signed(_zz_332));
  assign _zz_3611 = ({8'd0,data_mid_2_imag} <<< 8);
  assign _zz_3612 = {{8{_zz_3611[23]}}, _zz_3611};
  assign _zz_3613 = fixTo_399_dout;
  assign _zz_3614 = _zz_3615[31 : 0];
  assign _zz_3615 = _zz_3616;
  assign _zz_3616 = ($signed(_zz_3617) >>> _zz_335);
  assign _zz_3617 = _zz_3618;
  assign _zz_3618 = ($signed(_zz_3620) + $signed(_zz_331));
  assign _zz_3619 = ({8'd0,data_mid_2_real} <<< 8);
  assign _zz_3620 = {{8{_zz_3619[23]}}, _zz_3619};
  assign _zz_3621 = fixTo_400_dout;
  assign _zz_3622 = _zz_3623[31 : 0];
  assign _zz_3623 = _zz_3624;
  assign _zz_3624 = ($signed(_zz_3625) >>> _zz_335);
  assign _zz_3625 = _zz_3626;
  assign _zz_3626 = ($signed(_zz_3628) + $signed(_zz_332));
  assign _zz_3627 = ({8'd0,data_mid_2_imag} <<< 8);
  assign _zz_3628 = {{8{_zz_3627[23]}}, _zz_3627};
  assign _zz_3629 = fixTo_401_dout;
  assign _zz_3630 = ($signed(twiddle_factor_table_18_real) + $signed(twiddle_factor_table_18_imag));
  assign _zz_3631 = ($signed(_zz_338) - $signed(_zz_3632));
  assign _zz_3632 = ($signed(_zz_3633) * $signed(twiddle_factor_table_18_imag));
  assign _zz_3633 = ($signed(data_mid_19_real) + $signed(data_mid_19_imag));
  assign _zz_3634 = fixTo_402_dout;
  assign _zz_3635 = ($signed(_zz_338) + $signed(_zz_3636));
  assign _zz_3636 = ($signed(_zz_3637) * $signed(twiddle_factor_table_18_real));
  assign _zz_3637 = ($signed(data_mid_19_imag) - $signed(data_mid_19_real));
  assign _zz_3638 = fixTo_403_dout;
  assign _zz_3639 = _zz_3640[31 : 0];
  assign _zz_3640 = _zz_3641;
  assign _zz_3641 = ($signed(_zz_3642) >>> _zz_339);
  assign _zz_3642 = _zz_3643;
  assign _zz_3643 = ($signed(_zz_3645) - $signed(_zz_336));
  assign _zz_3644 = ({8'd0,data_mid_3_real} <<< 8);
  assign _zz_3645 = {{8{_zz_3644[23]}}, _zz_3644};
  assign _zz_3646 = fixTo_404_dout;
  assign _zz_3647 = _zz_3648[31 : 0];
  assign _zz_3648 = _zz_3649;
  assign _zz_3649 = ($signed(_zz_3650) >>> _zz_339);
  assign _zz_3650 = _zz_3651;
  assign _zz_3651 = ($signed(_zz_3653) - $signed(_zz_337));
  assign _zz_3652 = ({8'd0,data_mid_3_imag} <<< 8);
  assign _zz_3653 = {{8{_zz_3652[23]}}, _zz_3652};
  assign _zz_3654 = fixTo_405_dout;
  assign _zz_3655 = _zz_3656[31 : 0];
  assign _zz_3656 = _zz_3657;
  assign _zz_3657 = ($signed(_zz_3658) >>> _zz_340);
  assign _zz_3658 = _zz_3659;
  assign _zz_3659 = ($signed(_zz_3661) + $signed(_zz_336));
  assign _zz_3660 = ({8'd0,data_mid_3_real} <<< 8);
  assign _zz_3661 = {{8{_zz_3660[23]}}, _zz_3660};
  assign _zz_3662 = fixTo_406_dout;
  assign _zz_3663 = _zz_3664[31 : 0];
  assign _zz_3664 = _zz_3665;
  assign _zz_3665 = ($signed(_zz_3666) >>> _zz_340);
  assign _zz_3666 = _zz_3667;
  assign _zz_3667 = ($signed(_zz_3669) + $signed(_zz_337));
  assign _zz_3668 = ({8'd0,data_mid_3_imag} <<< 8);
  assign _zz_3669 = {{8{_zz_3668[23]}}, _zz_3668};
  assign _zz_3670 = fixTo_407_dout;
  assign _zz_3671 = ($signed(twiddle_factor_table_19_real) + $signed(twiddle_factor_table_19_imag));
  assign _zz_3672 = ($signed(_zz_343) - $signed(_zz_3673));
  assign _zz_3673 = ($signed(_zz_3674) * $signed(twiddle_factor_table_19_imag));
  assign _zz_3674 = ($signed(data_mid_20_real) + $signed(data_mid_20_imag));
  assign _zz_3675 = fixTo_408_dout;
  assign _zz_3676 = ($signed(_zz_343) + $signed(_zz_3677));
  assign _zz_3677 = ($signed(_zz_3678) * $signed(twiddle_factor_table_19_real));
  assign _zz_3678 = ($signed(data_mid_20_imag) - $signed(data_mid_20_real));
  assign _zz_3679 = fixTo_409_dout;
  assign _zz_3680 = _zz_3681[31 : 0];
  assign _zz_3681 = _zz_3682;
  assign _zz_3682 = ($signed(_zz_3683) >>> _zz_344);
  assign _zz_3683 = _zz_3684;
  assign _zz_3684 = ($signed(_zz_3686) - $signed(_zz_341));
  assign _zz_3685 = ({8'd0,data_mid_4_real} <<< 8);
  assign _zz_3686 = {{8{_zz_3685[23]}}, _zz_3685};
  assign _zz_3687 = fixTo_410_dout;
  assign _zz_3688 = _zz_3689[31 : 0];
  assign _zz_3689 = _zz_3690;
  assign _zz_3690 = ($signed(_zz_3691) >>> _zz_344);
  assign _zz_3691 = _zz_3692;
  assign _zz_3692 = ($signed(_zz_3694) - $signed(_zz_342));
  assign _zz_3693 = ({8'd0,data_mid_4_imag} <<< 8);
  assign _zz_3694 = {{8{_zz_3693[23]}}, _zz_3693};
  assign _zz_3695 = fixTo_411_dout;
  assign _zz_3696 = _zz_3697[31 : 0];
  assign _zz_3697 = _zz_3698;
  assign _zz_3698 = ($signed(_zz_3699) >>> _zz_345);
  assign _zz_3699 = _zz_3700;
  assign _zz_3700 = ($signed(_zz_3702) + $signed(_zz_341));
  assign _zz_3701 = ({8'd0,data_mid_4_real} <<< 8);
  assign _zz_3702 = {{8{_zz_3701[23]}}, _zz_3701};
  assign _zz_3703 = fixTo_412_dout;
  assign _zz_3704 = _zz_3705[31 : 0];
  assign _zz_3705 = _zz_3706;
  assign _zz_3706 = ($signed(_zz_3707) >>> _zz_345);
  assign _zz_3707 = _zz_3708;
  assign _zz_3708 = ($signed(_zz_3710) + $signed(_zz_342));
  assign _zz_3709 = ({8'd0,data_mid_4_imag} <<< 8);
  assign _zz_3710 = {{8{_zz_3709[23]}}, _zz_3709};
  assign _zz_3711 = fixTo_413_dout;
  assign _zz_3712 = ($signed(twiddle_factor_table_20_real) + $signed(twiddle_factor_table_20_imag));
  assign _zz_3713 = ($signed(_zz_348) - $signed(_zz_3714));
  assign _zz_3714 = ($signed(_zz_3715) * $signed(twiddle_factor_table_20_imag));
  assign _zz_3715 = ($signed(data_mid_21_real) + $signed(data_mid_21_imag));
  assign _zz_3716 = fixTo_414_dout;
  assign _zz_3717 = ($signed(_zz_348) + $signed(_zz_3718));
  assign _zz_3718 = ($signed(_zz_3719) * $signed(twiddle_factor_table_20_real));
  assign _zz_3719 = ($signed(data_mid_21_imag) - $signed(data_mid_21_real));
  assign _zz_3720 = fixTo_415_dout;
  assign _zz_3721 = _zz_3722[31 : 0];
  assign _zz_3722 = _zz_3723;
  assign _zz_3723 = ($signed(_zz_3724) >>> _zz_349);
  assign _zz_3724 = _zz_3725;
  assign _zz_3725 = ($signed(_zz_3727) - $signed(_zz_346));
  assign _zz_3726 = ({8'd0,data_mid_5_real} <<< 8);
  assign _zz_3727 = {{8{_zz_3726[23]}}, _zz_3726};
  assign _zz_3728 = fixTo_416_dout;
  assign _zz_3729 = _zz_3730[31 : 0];
  assign _zz_3730 = _zz_3731;
  assign _zz_3731 = ($signed(_zz_3732) >>> _zz_349);
  assign _zz_3732 = _zz_3733;
  assign _zz_3733 = ($signed(_zz_3735) - $signed(_zz_347));
  assign _zz_3734 = ({8'd0,data_mid_5_imag} <<< 8);
  assign _zz_3735 = {{8{_zz_3734[23]}}, _zz_3734};
  assign _zz_3736 = fixTo_417_dout;
  assign _zz_3737 = _zz_3738[31 : 0];
  assign _zz_3738 = _zz_3739;
  assign _zz_3739 = ($signed(_zz_3740) >>> _zz_350);
  assign _zz_3740 = _zz_3741;
  assign _zz_3741 = ($signed(_zz_3743) + $signed(_zz_346));
  assign _zz_3742 = ({8'd0,data_mid_5_real} <<< 8);
  assign _zz_3743 = {{8{_zz_3742[23]}}, _zz_3742};
  assign _zz_3744 = fixTo_418_dout;
  assign _zz_3745 = _zz_3746[31 : 0];
  assign _zz_3746 = _zz_3747;
  assign _zz_3747 = ($signed(_zz_3748) >>> _zz_350);
  assign _zz_3748 = _zz_3749;
  assign _zz_3749 = ($signed(_zz_3751) + $signed(_zz_347));
  assign _zz_3750 = ({8'd0,data_mid_5_imag} <<< 8);
  assign _zz_3751 = {{8{_zz_3750[23]}}, _zz_3750};
  assign _zz_3752 = fixTo_419_dout;
  assign _zz_3753 = ($signed(twiddle_factor_table_21_real) + $signed(twiddle_factor_table_21_imag));
  assign _zz_3754 = ($signed(_zz_353) - $signed(_zz_3755));
  assign _zz_3755 = ($signed(_zz_3756) * $signed(twiddle_factor_table_21_imag));
  assign _zz_3756 = ($signed(data_mid_22_real) + $signed(data_mid_22_imag));
  assign _zz_3757 = fixTo_420_dout;
  assign _zz_3758 = ($signed(_zz_353) + $signed(_zz_3759));
  assign _zz_3759 = ($signed(_zz_3760) * $signed(twiddle_factor_table_21_real));
  assign _zz_3760 = ($signed(data_mid_22_imag) - $signed(data_mid_22_real));
  assign _zz_3761 = fixTo_421_dout;
  assign _zz_3762 = _zz_3763[31 : 0];
  assign _zz_3763 = _zz_3764;
  assign _zz_3764 = ($signed(_zz_3765) >>> _zz_354);
  assign _zz_3765 = _zz_3766;
  assign _zz_3766 = ($signed(_zz_3768) - $signed(_zz_351));
  assign _zz_3767 = ({8'd0,data_mid_6_real} <<< 8);
  assign _zz_3768 = {{8{_zz_3767[23]}}, _zz_3767};
  assign _zz_3769 = fixTo_422_dout;
  assign _zz_3770 = _zz_3771[31 : 0];
  assign _zz_3771 = _zz_3772;
  assign _zz_3772 = ($signed(_zz_3773) >>> _zz_354);
  assign _zz_3773 = _zz_3774;
  assign _zz_3774 = ($signed(_zz_3776) - $signed(_zz_352));
  assign _zz_3775 = ({8'd0,data_mid_6_imag} <<< 8);
  assign _zz_3776 = {{8{_zz_3775[23]}}, _zz_3775};
  assign _zz_3777 = fixTo_423_dout;
  assign _zz_3778 = _zz_3779[31 : 0];
  assign _zz_3779 = _zz_3780;
  assign _zz_3780 = ($signed(_zz_3781) >>> _zz_355);
  assign _zz_3781 = _zz_3782;
  assign _zz_3782 = ($signed(_zz_3784) + $signed(_zz_351));
  assign _zz_3783 = ({8'd0,data_mid_6_real} <<< 8);
  assign _zz_3784 = {{8{_zz_3783[23]}}, _zz_3783};
  assign _zz_3785 = fixTo_424_dout;
  assign _zz_3786 = _zz_3787[31 : 0];
  assign _zz_3787 = _zz_3788;
  assign _zz_3788 = ($signed(_zz_3789) >>> _zz_355);
  assign _zz_3789 = _zz_3790;
  assign _zz_3790 = ($signed(_zz_3792) + $signed(_zz_352));
  assign _zz_3791 = ({8'd0,data_mid_6_imag} <<< 8);
  assign _zz_3792 = {{8{_zz_3791[23]}}, _zz_3791};
  assign _zz_3793 = fixTo_425_dout;
  assign _zz_3794 = ($signed(twiddle_factor_table_22_real) + $signed(twiddle_factor_table_22_imag));
  assign _zz_3795 = ($signed(_zz_358) - $signed(_zz_3796));
  assign _zz_3796 = ($signed(_zz_3797) * $signed(twiddle_factor_table_22_imag));
  assign _zz_3797 = ($signed(data_mid_23_real) + $signed(data_mid_23_imag));
  assign _zz_3798 = fixTo_426_dout;
  assign _zz_3799 = ($signed(_zz_358) + $signed(_zz_3800));
  assign _zz_3800 = ($signed(_zz_3801) * $signed(twiddle_factor_table_22_real));
  assign _zz_3801 = ($signed(data_mid_23_imag) - $signed(data_mid_23_real));
  assign _zz_3802 = fixTo_427_dout;
  assign _zz_3803 = _zz_3804[31 : 0];
  assign _zz_3804 = _zz_3805;
  assign _zz_3805 = ($signed(_zz_3806) >>> _zz_359);
  assign _zz_3806 = _zz_3807;
  assign _zz_3807 = ($signed(_zz_3809) - $signed(_zz_356));
  assign _zz_3808 = ({8'd0,data_mid_7_real} <<< 8);
  assign _zz_3809 = {{8{_zz_3808[23]}}, _zz_3808};
  assign _zz_3810 = fixTo_428_dout;
  assign _zz_3811 = _zz_3812[31 : 0];
  assign _zz_3812 = _zz_3813;
  assign _zz_3813 = ($signed(_zz_3814) >>> _zz_359);
  assign _zz_3814 = _zz_3815;
  assign _zz_3815 = ($signed(_zz_3817) - $signed(_zz_357));
  assign _zz_3816 = ({8'd0,data_mid_7_imag} <<< 8);
  assign _zz_3817 = {{8{_zz_3816[23]}}, _zz_3816};
  assign _zz_3818 = fixTo_429_dout;
  assign _zz_3819 = _zz_3820[31 : 0];
  assign _zz_3820 = _zz_3821;
  assign _zz_3821 = ($signed(_zz_3822) >>> _zz_360);
  assign _zz_3822 = _zz_3823;
  assign _zz_3823 = ($signed(_zz_3825) + $signed(_zz_356));
  assign _zz_3824 = ({8'd0,data_mid_7_real} <<< 8);
  assign _zz_3825 = {{8{_zz_3824[23]}}, _zz_3824};
  assign _zz_3826 = fixTo_430_dout;
  assign _zz_3827 = _zz_3828[31 : 0];
  assign _zz_3828 = _zz_3829;
  assign _zz_3829 = ($signed(_zz_3830) >>> _zz_360);
  assign _zz_3830 = _zz_3831;
  assign _zz_3831 = ($signed(_zz_3833) + $signed(_zz_357));
  assign _zz_3832 = ({8'd0,data_mid_7_imag} <<< 8);
  assign _zz_3833 = {{8{_zz_3832[23]}}, _zz_3832};
  assign _zz_3834 = fixTo_431_dout;
  assign _zz_3835 = ($signed(twiddle_factor_table_23_real) + $signed(twiddle_factor_table_23_imag));
  assign _zz_3836 = ($signed(_zz_363) - $signed(_zz_3837));
  assign _zz_3837 = ($signed(_zz_3838) * $signed(twiddle_factor_table_23_imag));
  assign _zz_3838 = ($signed(data_mid_24_real) + $signed(data_mid_24_imag));
  assign _zz_3839 = fixTo_432_dout;
  assign _zz_3840 = ($signed(_zz_363) + $signed(_zz_3841));
  assign _zz_3841 = ($signed(_zz_3842) * $signed(twiddle_factor_table_23_real));
  assign _zz_3842 = ($signed(data_mid_24_imag) - $signed(data_mid_24_real));
  assign _zz_3843 = fixTo_433_dout;
  assign _zz_3844 = _zz_3845[31 : 0];
  assign _zz_3845 = _zz_3846;
  assign _zz_3846 = ($signed(_zz_3847) >>> _zz_364);
  assign _zz_3847 = _zz_3848;
  assign _zz_3848 = ($signed(_zz_3850) - $signed(_zz_361));
  assign _zz_3849 = ({8'd0,data_mid_8_real} <<< 8);
  assign _zz_3850 = {{8{_zz_3849[23]}}, _zz_3849};
  assign _zz_3851 = fixTo_434_dout;
  assign _zz_3852 = _zz_3853[31 : 0];
  assign _zz_3853 = _zz_3854;
  assign _zz_3854 = ($signed(_zz_3855) >>> _zz_364);
  assign _zz_3855 = _zz_3856;
  assign _zz_3856 = ($signed(_zz_3858) - $signed(_zz_362));
  assign _zz_3857 = ({8'd0,data_mid_8_imag} <<< 8);
  assign _zz_3858 = {{8{_zz_3857[23]}}, _zz_3857};
  assign _zz_3859 = fixTo_435_dout;
  assign _zz_3860 = _zz_3861[31 : 0];
  assign _zz_3861 = _zz_3862;
  assign _zz_3862 = ($signed(_zz_3863) >>> _zz_365);
  assign _zz_3863 = _zz_3864;
  assign _zz_3864 = ($signed(_zz_3866) + $signed(_zz_361));
  assign _zz_3865 = ({8'd0,data_mid_8_real} <<< 8);
  assign _zz_3866 = {{8{_zz_3865[23]}}, _zz_3865};
  assign _zz_3867 = fixTo_436_dout;
  assign _zz_3868 = _zz_3869[31 : 0];
  assign _zz_3869 = _zz_3870;
  assign _zz_3870 = ($signed(_zz_3871) >>> _zz_365);
  assign _zz_3871 = _zz_3872;
  assign _zz_3872 = ($signed(_zz_3874) + $signed(_zz_362));
  assign _zz_3873 = ({8'd0,data_mid_8_imag} <<< 8);
  assign _zz_3874 = {{8{_zz_3873[23]}}, _zz_3873};
  assign _zz_3875 = fixTo_437_dout;
  assign _zz_3876 = ($signed(twiddle_factor_table_24_real) + $signed(twiddle_factor_table_24_imag));
  assign _zz_3877 = ($signed(_zz_368) - $signed(_zz_3878));
  assign _zz_3878 = ($signed(_zz_3879) * $signed(twiddle_factor_table_24_imag));
  assign _zz_3879 = ($signed(data_mid_25_real) + $signed(data_mid_25_imag));
  assign _zz_3880 = fixTo_438_dout;
  assign _zz_3881 = ($signed(_zz_368) + $signed(_zz_3882));
  assign _zz_3882 = ($signed(_zz_3883) * $signed(twiddle_factor_table_24_real));
  assign _zz_3883 = ($signed(data_mid_25_imag) - $signed(data_mid_25_real));
  assign _zz_3884 = fixTo_439_dout;
  assign _zz_3885 = _zz_3886[31 : 0];
  assign _zz_3886 = _zz_3887;
  assign _zz_3887 = ($signed(_zz_3888) >>> _zz_369);
  assign _zz_3888 = _zz_3889;
  assign _zz_3889 = ($signed(_zz_3891) - $signed(_zz_366));
  assign _zz_3890 = ({8'd0,data_mid_9_real} <<< 8);
  assign _zz_3891 = {{8{_zz_3890[23]}}, _zz_3890};
  assign _zz_3892 = fixTo_440_dout;
  assign _zz_3893 = _zz_3894[31 : 0];
  assign _zz_3894 = _zz_3895;
  assign _zz_3895 = ($signed(_zz_3896) >>> _zz_369);
  assign _zz_3896 = _zz_3897;
  assign _zz_3897 = ($signed(_zz_3899) - $signed(_zz_367));
  assign _zz_3898 = ({8'd0,data_mid_9_imag} <<< 8);
  assign _zz_3899 = {{8{_zz_3898[23]}}, _zz_3898};
  assign _zz_3900 = fixTo_441_dout;
  assign _zz_3901 = _zz_3902[31 : 0];
  assign _zz_3902 = _zz_3903;
  assign _zz_3903 = ($signed(_zz_3904) >>> _zz_370);
  assign _zz_3904 = _zz_3905;
  assign _zz_3905 = ($signed(_zz_3907) + $signed(_zz_366));
  assign _zz_3906 = ({8'd0,data_mid_9_real} <<< 8);
  assign _zz_3907 = {{8{_zz_3906[23]}}, _zz_3906};
  assign _zz_3908 = fixTo_442_dout;
  assign _zz_3909 = _zz_3910[31 : 0];
  assign _zz_3910 = _zz_3911;
  assign _zz_3911 = ($signed(_zz_3912) >>> _zz_370);
  assign _zz_3912 = _zz_3913;
  assign _zz_3913 = ($signed(_zz_3915) + $signed(_zz_367));
  assign _zz_3914 = ({8'd0,data_mid_9_imag} <<< 8);
  assign _zz_3915 = {{8{_zz_3914[23]}}, _zz_3914};
  assign _zz_3916 = fixTo_443_dout;
  assign _zz_3917 = ($signed(twiddle_factor_table_25_real) + $signed(twiddle_factor_table_25_imag));
  assign _zz_3918 = ($signed(_zz_373) - $signed(_zz_3919));
  assign _zz_3919 = ($signed(_zz_3920) * $signed(twiddle_factor_table_25_imag));
  assign _zz_3920 = ($signed(data_mid_26_real) + $signed(data_mid_26_imag));
  assign _zz_3921 = fixTo_444_dout;
  assign _zz_3922 = ($signed(_zz_373) + $signed(_zz_3923));
  assign _zz_3923 = ($signed(_zz_3924) * $signed(twiddle_factor_table_25_real));
  assign _zz_3924 = ($signed(data_mid_26_imag) - $signed(data_mid_26_real));
  assign _zz_3925 = fixTo_445_dout;
  assign _zz_3926 = _zz_3927[31 : 0];
  assign _zz_3927 = _zz_3928;
  assign _zz_3928 = ($signed(_zz_3929) >>> _zz_374);
  assign _zz_3929 = _zz_3930;
  assign _zz_3930 = ($signed(_zz_3932) - $signed(_zz_371));
  assign _zz_3931 = ({8'd0,data_mid_10_real} <<< 8);
  assign _zz_3932 = {{8{_zz_3931[23]}}, _zz_3931};
  assign _zz_3933 = fixTo_446_dout;
  assign _zz_3934 = _zz_3935[31 : 0];
  assign _zz_3935 = _zz_3936;
  assign _zz_3936 = ($signed(_zz_3937) >>> _zz_374);
  assign _zz_3937 = _zz_3938;
  assign _zz_3938 = ($signed(_zz_3940) - $signed(_zz_372));
  assign _zz_3939 = ({8'd0,data_mid_10_imag} <<< 8);
  assign _zz_3940 = {{8{_zz_3939[23]}}, _zz_3939};
  assign _zz_3941 = fixTo_447_dout;
  assign _zz_3942 = _zz_3943[31 : 0];
  assign _zz_3943 = _zz_3944;
  assign _zz_3944 = ($signed(_zz_3945) >>> _zz_375);
  assign _zz_3945 = _zz_3946;
  assign _zz_3946 = ($signed(_zz_3948) + $signed(_zz_371));
  assign _zz_3947 = ({8'd0,data_mid_10_real} <<< 8);
  assign _zz_3948 = {{8{_zz_3947[23]}}, _zz_3947};
  assign _zz_3949 = fixTo_448_dout;
  assign _zz_3950 = _zz_3951[31 : 0];
  assign _zz_3951 = _zz_3952;
  assign _zz_3952 = ($signed(_zz_3953) >>> _zz_375);
  assign _zz_3953 = _zz_3954;
  assign _zz_3954 = ($signed(_zz_3956) + $signed(_zz_372));
  assign _zz_3955 = ({8'd0,data_mid_10_imag} <<< 8);
  assign _zz_3956 = {{8{_zz_3955[23]}}, _zz_3955};
  assign _zz_3957 = fixTo_449_dout;
  assign _zz_3958 = ($signed(twiddle_factor_table_26_real) + $signed(twiddle_factor_table_26_imag));
  assign _zz_3959 = ($signed(_zz_378) - $signed(_zz_3960));
  assign _zz_3960 = ($signed(_zz_3961) * $signed(twiddle_factor_table_26_imag));
  assign _zz_3961 = ($signed(data_mid_27_real) + $signed(data_mid_27_imag));
  assign _zz_3962 = fixTo_450_dout;
  assign _zz_3963 = ($signed(_zz_378) + $signed(_zz_3964));
  assign _zz_3964 = ($signed(_zz_3965) * $signed(twiddle_factor_table_26_real));
  assign _zz_3965 = ($signed(data_mid_27_imag) - $signed(data_mid_27_real));
  assign _zz_3966 = fixTo_451_dout;
  assign _zz_3967 = _zz_3968[31 : 0];
  assign _zz_3968 = _zz_3969;
  assign _zz_3969 = ($signed(_zz_3970) >>> _zz_379);
  assign _zz_3970 = _zz_3971;
  assign _zz_3971 = ($signed(_zz_3973) - $signed(_zz_376));
  assign _zz_3972 = ({8'd0,data_mid_11_real} <<< 8);
  assign _zz_3973 = {{8{_zz_3972[23]}}, _zz_3972};
  assign _zz_3974 = fixTo_452_dout;
  assign _zz_3975 = _zz_3976[31 : 0];
  assign _zz_3976 = _zz_3977;
  assign _zz_3977 = ($signed(_zz_3978) >>> _zz_379);
  assign _zz_3978 = _zz_3979;
  assign _zz_3979 = ($signed(_zz_3981) - $signed(_zz_377));
  assign _zz_3980 = ({8'd0,data_mid_11_imag} <<< 8);
  assign _zz_3981 = {{8{_zz_3980[23]}}, _zz_3980};
  assign _zz_3982 = fixTo_453_dout;
  assign _zz_3983 = _zz_3984[31 : 0];
  assign _zz_3984 = _zz_3985;
  assign _zz_3985 = ($signed(_zz_3986) >>> _zz_380);
  assign _zz_3986 = _zz_3987;
  assign _zz_3987 = ($signed(_zz_3989) + $signed(_zz_376));
  assign _zz_3988 = ({8'd0,data_mid_11_real} <<< 8);
  assign _zz_3989 = {{8{_zz_3988[23]}}, _zz_3988};
  assign _zz_3990 = fixTo_454_dout;
  assign _zz_3991 = _zz_3992[31 : 0];
  assign _zz_3992 = _zz_3993;
  assign _zz_3993 = ($signed(_zz_3994) >>> _zz_380);
  assign _zz_3994 = _zz_3995;
  assign _zz_3995 = ($signed(_zz_3997) + $signed(_zz_377));
  assign _zz_3996 = ({8'd0,data_mid_11_imag} <<< 8);
  assign _zz_3997 = {{8{_zz_3996[23]}}, _zz_3996};
  assign _zz_3998 = fixTo_455_dout;
  assign _zz_3999 = ($signed(twiddle_factor_table_27_real) + $signed(twiddle_factor_table_27_imag));
  assign _zz_4000 = ($signed(_zz_383) - $signed(_zz_4001));
  assign _zz_4001 = ($signed(_zz_4002) * $signed(twiddle_factor_table_27_imag));
  assign _zz_4002 = ($signed(data_mid_28_real) + $signed(data_mid_28_imag));
  assign _zz_4003 = fixTo_456_dout;
  assign _zz_4004 = ($signed(_zz_383) + $signed(_zz_4005));
  assign _zz_4005 = ($signed(_zz_4006) * $signed(twiddle_factor_table_27_real));
  assign _zz_4006 = ($signed(data_mid_28_imag) - $signed(data_mid_28_real));
  assign _zz_4007 = fixTo_457_dout;
  assign _zz_4008 = _zz_4009[31 : 0];
  assign _zz_4009 = _zz_4010;
  assign _zz_4010 = ($signed(_zz_4011) >>> _zz_384);
  assign _zz_4011 = _zz_4012;
  assign _zz_4012 = ($signed(_zz_4014) - $signed(_zz_381));
  assign _zz_4013 = ({8'd0,data_mid_12_real} <<< 8);
  assign _zz_4014 = {{8{_zz_4013[23]}}, _zz_4013};
  assign _zz_4015 = fixTo_458_dout;
  assign _zz_4016 = _zz_4017[31 : 0];
  assign _zz_4017 = _zz_4018;
  assign _zz_4018 = ($signed(_zz_4019) >>> _zz_384);
  assign _zz_4019 = _zz_4020;
  assign _zz_4020 = ($signed(_zz_4022) - $signed(_zz_382));
  assign _zz_4021 = ({8'd0,data_mid_12_imag} <<< 8);
  assign _zz_4022 = {{8{_zz_4021[23]}}, _zz_4021};
  assign _zz_4023 = fixTo_459_dout;
  assign _zz_4024 = _zz_4025[31 : 0];
  assign _zz_4025 = _zz_4026;
  assign _zz_4026 = ($signed(_zz_4027) >>> _zz_385);
  assign _zz_4027 = _zz_4028;
  assign _zz_4028 = ($signed(_zz_4030) + $signed(_zz_381));
  assign _zz_4029 = ({8'd0,data_mid_12_real} <<< 8);
  assign _zz_4030 = {{8{_zz_4029[23]}}, _zz_4029};
  assign _zz_4031 = fixTo_460_dout;
  assign _zz_4032 = _zz_4033[31 : 0];
  assign _zz_4033 = _zz_4034;
  assign _zz_4034 = ($signed(_zz_4035) >>> _zz_385);
  assign _zz_4035 = _zz_4036;
  assign _zz_4036 = ($signed(_zz_4038) + $signed(_zz_382));
  assign _zz_4037 = ({8'd0,data_mid_12_imag} <<< 8);
  assign _zz_4038 = {{8{_zz_4037[23]}}, _zz_4037};
  assign _zz_4039 = fixTo_461_dout;
  assign _zz_4040 = ($signed(twiddle_factor_table_28_real) + $signed(twiddle_factor_table_28_imag));
  assign _zz_4041 = ($signed(_zz_388) - $signed(_zz_4042));
  assign _zz_4042 = ($signed(_zz_4043) * $signed(twiddle_factor_table_28_imag));
  assign _zz_4043 = ($signed(data_mid_29_real) + $signed(data_mid_29_imag));
  assign _zz_4044 = fixTo_462_dout;
  assign _zz_4045 = ($signed(_zz_388) + $signed(_zz_4046));
  assign _zz_4046 = ($signed(_zz_4047) * $signed(twiddle_factor_table_28_real));
  assign _zz_4047 = ($signed(data_mid_29_imag) - $signed(data_mid_29_real));
  assign _zz_4048 = fixTo_463_dout;
  assign _zz_4049 = _zz_4050[31 : 0];
  assign _zz_4050 = _zz_4051;
  assign _zz_4051 = ($signed(_zz_4052) >>> _zz_389);
  assign _zz_4052 = _zz_4053;
  assign _zz_4053 = ($signed(_zz_4055) - $signed(_zz_386));
  assign _zz_4054 = ({8'd0,data_mid_13_real} <<< 8);
  assign _zz_4055 = {{8{_zz_4054[23]}}, _zz_4054};
  assign _zz_4056 = fixTo_464_dout;
  assign _zz_4057 = _zz_4058[31 : 0];
  assign _zz_4058 = _zz_4059;
  assign _zz_4059 = ($signed(_zz_4060) >>> _zz_389);
  assign _zz_4060 = _zz_4061;
  assign _zz_4061 = ($signed(_zz_4063) - $signed(_zz_387));
  assign _zz_4062 = ({8'd0,data_mid_13_imag} <<< 8);
  assign _zz_4063 = {{8{_zz_4062[23]}}, _zz_4062};
  assign _zz_4064 = fixTo_465_dout;
  assign _zz_4065 = _zz_4066[31 : 0];
  assign _zz_4066 = _zz_4067;
  assign _zz_4067 = ($signed(_zz_4068) >>> _zz_390);
  assign _zz_4068 = _zz_4069;
  assign _zz_4069 = ($signed(_zz_4071) + $signed(_zz_386));
  assign _zz_4070 = ({8'd0,data_mid_13_real} <<< 8);
  assign _zz_4071 = {{8{_zz_4070[23]}}, _zz_4070};
  assign _zz_4072 = fixTo_466_dout;
  assign _zz_4073 = _zz_4074[31 : 0];
  assign _zz_4074 = _zz_4075;
  assign _zz_4075 = ($signed(_zz_4076) >>> _zz_390);
  assign _zz_4076 = _zz_4077;
  assign _zz_4077 = ($signed(_zz_4079) + $signed(_zz_387));
  assign _zz_4078 = ({8'd0,data_mid_13_imag} <<< 8);
  assign _zz_4079 = {{8{_zz_4078[23]}}, _zz_4078};
  assign _zz_4080 = fixTo_467_dout;
  assign _zz_4081 = ($signed(twiddle_factor_table_29_real) + $signed(twiddle_factor_table_29_imag));
  assign _zz_4082 = ($signed(_zz_393) - $signed(_zz_4083));
  assign _zz_4083 = ($signed(_zz_4084) * $signed(twiddle_factor_table_29_imag));
  assign _zz_4084 = ($signed(data_mid_30_real) + $signed(data_mid_30_imag));
  assign _zz_4085 = fixTo_468_dout;
  assign _zz_4086 = ($signed(_zz_393) + $signed(_zz_4087));
  assign _zz_4087 = ($signed(_zz_4088) * $signed(twiddle_factor_table_29_real));
  assign _zz_4088 = ($signed(data_mid_30_imag) - $signed(data_mid_30_real));
  assign _zz_4089 = fixTo_469_dout;
  assign _zz_4090 = _zz_4091[31 : 0];
  assign _zz_4091 = _zz_4092;
  assign _zz_4092 = ($signed(_zz_4093) >>> _zz_394);
  assign _zz_4093 = _zz_4094;
  assign _zz_4094 = ($signed(_zz_4096) - $signed(_zz_391));
  assign _zz_4095 = ({8'd0,data_mid_14_real} <<< 8);
  assign _zz_4096 = {{8{_zz_4095[23]}}, _zz_4095};
  assign _zz_4097 = fixTo_470_dout;
  assign _zz_4098 = _zz_4099[31 : 0];
  assign _zz_4099 = _zz_4100;
  assign _zz_4100 = ($signed(_zz_4101) >>> _zz_394);
  assign _zz_4101 = _zz_4102;
  assign _zz_4102 = ($signed(_zz_4104) - $signed(_zz_392));
  assign _zz_4103 = ({8'd0,data_mid_14_imag} <<< 8);
  assign _zz_4104 = {{8{_zz_4103[23]}}, _zz_4103};
  assign _zz_4105 = fixTo_471_dout;
  assign _zz_4106 = _zz_4107[31 : 0];
  assign _zz_4107 = _zz_4108;
  assign _zz_4108 = ($signed(_zz_4109) >>> _zz_395);
  assign _zz_4109 = _zz_4110;
  assign _zz_4110 = ($signed(_zz_4112) + $signed(_zz_391));
  assign _zz_4111 = ({8'd0,data_mid_14_real} <<< 8);
  assign _zz_4112 = {{8{_zz_4111[23]}}, _zz_4111};
  assign _zz_4113 = fixTo_472_dout;
  assign _zz_4114 = _zz_4115[31 : 0];
  assign _zz_4115 = _zz_4116;
  assign _zz_4116 = ($signed(_zz_4117) >>> _zz_395);
  assign _zz_4117 = _zz_4118;
  assign _zz_4118 = ($signed(_zz_4120) + $signed(_zz_392));
  assign _zz_4119 = ({8'd0,data_mid_14_imag} <<< 8);
  assign _zz_4120 = {{8{_zz_4119[23]}}, _zz_4119};
  assign _zz_4121 = fixTo_473_dout;
  assign _zz_4122 = ($signed(twiddle_factor_table_30_real) + $signed(twiddle_factor_table_30_imag));
  assign _zz_4123 = ($signed(_zz_398) - $signed(_zz_4124));
  assign _zz_4124 = ($signed(_zz_4125) * $signed(twiddle_factor_table_30_imag));
  assign _zz_4125 = ($signed(data_mid_31_real) + $signed(data_mid_31_imag));
  assign _zz_4126 = fixTo_474_dout;
  assign _zz_4127 = ($signed(_zz_398) + $signed(_zz_4128));
  assign _zz_4128 = ($signed(_zz_4129) * $signed(twiddle_factor_table_30_real));
  assign _zz_4129 = ($signed(data_mid_31_imag) - $signed(data_mid_31_real));
  assign _zz_4130 = fixTo_475_dout;
  assign _zz_4131 = _zz_4132[31 : 0];
  assign _zz_4132 = _zz_4133;
  assign _zz_4133 = ($signed(_zz_4134) >>> _zz_399);
  assign _zz_4134 = _zz_4135;
  assign _zz_4135 = ($signed(_zz_4137) - $signed(_zz_396));
  assign _zz_4136 = ({8'd0,data_mid_15_real} <<< 8);
  assign _zz_4137 = {{8{_zz_4136[23]}}, _zz_4136};
  assign _zz_4138 = fixTo_476_dout;
  assign _zz_4139 = _zz_4140[31 : 0];
  assign _zz_4140 = _zz_4141;
  assign _zz_4141 = ($signed(_zz_4142) >>> _zz_399);
  assign _zz_4142 = _zz_4143;
  assign _zz_4143 = ($signed(_zz_4145) - $signed(_zz_397));
  assign _zz_4144 = ({8'd0,data_mid_15_imag} <<< 8);
  assign _zz_4145 = {{8{_zz_4144[23]}}, _zz_4144};
  assign _zz_4146 = fixTo_477_dout;
  assign _zz_4147 = _zz_4148[31 : 0];
  assign _zz_4148 = _zz_4149;
  assign _zz_4149 = ($signed(_zz_4150) >>> _zz_400);
  assign _zz_4150 = _zz_4151;
  assign _zz_4151 = ($signed(_zz_4153) + $signed(_zz_396));
  assign _zz_4152 = ({8'd0,data_mid_15_real} <<< 8);
  assign _zz_4153 = {{8{_zz_4152[23]}}, _zz_4152};
  assign _zz_4154 = fixTo_478_dout;
  assign _zz_4155 = _zz_4156[31 : 0];
  assign _zz_4156 = _zz_4157;
  assign _zz_4157 = ($signed(_zz_4158) >>> _zz_400);
  assign _zz_4158 = _zz_4159;
  assign _zz_4159 = ($signed(_zz_4161) + $signed(_zz_397));
  assign _zz_4160 = ({8'd0,data_mid_15_imag} <<< 8);
  assign _zz_4161 = {{8{_zz_4160[23]}}, _zz_4160};
  assign _zz_4162 = fixTo_479_dout;
  SInt32fixTo31_0_ROUNDTOINF fixTo (
    .din     (_zz_401[31:0]     ), //i
    .dout    (fixTo_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_1 (
    .din     (_zz_402[31:0]       ), //i
    .dout    (fixTo_1_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_2 (
    .din     (_zz_403[31:0]       ), //i
    .dout    (fixTo_2_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_3 (
    .din     (_zz_404[31:0]       ), //i
    .dout    (fixTo_3_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_4 (
    .din     (_zz_405[31:0]       ), //i
    .dout    (fixTo_4_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_5 (
    .din     (_zz_406[31:0]       ), //i
    .dout    (fixTo_5_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_6 (
    .din     (_zz_407[31:0]       ), //i
    .dout    (fixTo_6_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_7 (
    .din     (_zz_408[31:0]       ), //i
    .dout    (fixTo_7_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_8 (
    .din     (_zz_409[31:0]       ), //i
    .dout    (fixTo_8_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_9 (
    .din     (_zz_410[31:0]       ), //i
    .dout    (fixTo_9_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_10 (
    .din     (_zz_411[31:0]        ), //i
    .dout    (fixTo_10_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_11 (
    .din     (_zz_412[31:0]        ), //i
    .dout    (fixTo_11_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_12 (
    .din     (_zz_413[31:0]        ), //i
    .dout    (fixTo_12_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_13 (
    .din     (_zz_414[31:0]        ), //i
    .dout    (fixTo_13_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_14 (
    .din     (_zz_415[31:0]        ), //i
    .dout    (fixTo_14_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_15 (
    .din     (_zz_416[31:0]        ), //i
    .dout    (fixTo_15_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_16 (
    .din     (_zz_417[31:0]        ), //i
    .dout    (fixTo_16_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_17 (
    .din     (_zz_418[31:0]        ), //i
    .dout    (fixTo_17_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_18 (
    .din     (_zz_419[31:0]        ), //i
    .dout    (fixTo_18_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_19 (
    .din     (_zz_420[31:0]        ), //i
    .dout    (fixTo_19_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_20 (
    .din     (_zz_421[31:0]        ), //i
    .dout    (fixTo_20_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_21 (
    .din     (_zz_422[31:0]        ), //i
    .dout    (fixTo_21_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_22 (
    .din     (_zz_423[31:0]        ), //i
    .dout    (fixTo_22_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_23 (
    .din     (_zz_424[31:0]        ), //i
    .dout    (fixTo_23_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_24 (
    .din     (_zz_425[31:0]        ), //i
    .dout    (fixTo_24_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_25 (
    .din     (_zz_426[31:0]        ), //i
    .dout    (fixTo_25_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_26 (
    .din     (_zz_427[31:0]        ), //i
    .dout    (fixTo_26_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_27 (
    .din     (_zz_428[31:0]        ), //i
    .dout    (fixTo_27_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_28 (
    .din     (_zz_429[31:0]        ), //i
    .dout    (fixTo_28_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_29 (
    .din     (_zz_430[31:0]        ), //i
    .dout    (fixTo_29_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_30 (
    .din     (_zz_431[31:0]        ), //i
    .dout    (fixTo_30_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_31 (
    .din     (_zz_432[31:0]        ), //i
    .dout    (fixTo_31_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_32 (
    .din     (_zz_433[31:0]        ), //i
    .dout    (fixTo_32_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_33 (
    .din     (_zz_434[31:0]        ), //i
    .dout    (fixTo_33_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_34 (
    .din     (_zz_435[31:0]        ), //i
    .dout    (fixTo_34_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_35 (
    .din     (_zz_436[31:0]        ), //i
    .dout    (fixTo_35_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_36 (
    .din     (_zz_437[31:0]        ), //i
    .dout    (fixTo_36_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_37 (
    .din     (_zz_438[31:0]        ), //i
    .dout    (fixTo_37_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_38 (
    .din     (_zz_439[31:0]        ), //i
    .dout    (fixTo_38_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_39 (
    .din     (_zz_440[31:0]        ), //i
    .dout    (fixTo_39_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_40 (
    .din     (_zz_441[31:0]        ), //i
    .dout    (fixTo_40_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_41 (
    .din     (_zz_442[31:0]        ), //i
    .dout    (fixTo_41_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_42 (
    .din     (_zz_443[31:0]        ), //i
    .dout    (fixTo_42_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_43 (
    .din     (_zz_444[31:0]        ), //i
    .dout    (fixTo_43_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_44 (
    .din     (_zz_445[31:0]        ), //i
    .dout    (fixTo_44_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_45 (
    .din     (_zz_446[31:0]        ), //i
    .dout    (fixTo_45_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_46 (
    .din     (_zz_447[31:0]        ), //i
    .dout    (fixTo_46_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_47 (
    .din     (_zz_448[31:0]        ), //i
    .dout    (fixTo_47_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_48 (
    .din     (_zz_449[31:0]        ), //i
    .dout    (fixTo_48_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_49 (
    .din     (_zz_450[31:0]        ), //i
    .dout    (fixTo_49_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_50 (
    .din     (_zz_451[31:0]        ), //i
    .dout    (fixTo_50_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_51 (
    .din     (_zz_452[31:0]        ), //i
    .dout    (fixTo_51_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_52 (
    .din     (_zz_453[31:0]        ), //i
    .dout    (fixTo_52_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_53 (
    .din     (_zz_454[31:0]        ), //i
    .dout    (fixTo_53_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_54 (
    .din     (_zz_455[31:0]        ), //i
    .dout    (fixTo_54_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_55 (
    .din     (_zz_456[31:0]        ), //i
    .dout    (fixTo_55_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_56 (
    .din     (_zz_457[31:0]        ), //i
    .dout    (fixTo_56_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_57 (
    .din     (_zz_458[31:0]        ), //i
    .dout    (fixTo_57_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_58 (
    .din     (_zz_459[31:0]        ), //i
    .dout    (fixTo_58_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_59 (
    .din     (_zz_460[31:0]        ), //i
    .dout    (fixTo_59_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_60 (
    .din     (_zz_461[31:0]        ), //i
    .dout    (fixTo_60_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_61 (
    .din     (_zz_462[31:0]        ), //i
    .dout    (fixTo_61_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_62 (
    .din     (_zz_463[31:0]        ), //i
    .dout    (fixTo_62_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_63 (
    .din     (_zz_464[31:0]        ), //i
    .dout    (fixTo_63_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_64 (
    .din     (_zz_465[31:0]        ), //i
    .dout    (fixTo_64_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_65 (
    .din     (_zz_466[31:0]        ), //i
    .dout    (fixTo_65_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_66 (
    .din     (_zz_467[31:0]        ), //i
    .dout    (fixTo_66_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_67 (
    .din     (_zz_468[31:0]        ), //i
    .dout    (fixTo_67_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_68 (
    .din     (_zz_469[31:0]        ), //i
    .dout    (fixTo_68_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_69 (
    .din     (_zz_470[31:0]        ), //i
    .dout    (fixTo_69_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_70 (
    .din     (_zz_471[31:0]        ), //i
    .dout    (fixTo_70_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_71 (
    .din     (_zz_472[31:0]        ), //i
    .dout    (fixTo_71_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_72 (
    .din     (_zz_473[31:0]        ), //i
    .dout    (fixTo_72_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_73 (
    .din     (_zz_474[31:0]        ), //i
    .dout    (fixTo_73_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_74 (
    .din     (_zz_475[31:0]        ), //i
    .dout    (fixTo_74_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_75 (
    .din     (_zz_476[31:0]        ), //i
    .dout    (fixTo_75_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_76 (
    .din     (_zz_477[31:0]        ), //i
    .dout    (fixTo_76_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_77 (
    .din     (_zz_478[31:0]        ), //i
    .dout    (fixTo_77_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_78 (
    .din     (_zz_479[31:0]        ), //i
    .dout    (fixTo_78_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_79 (
    .din     (_zz_480[31:0]        ), //i
    .dout    (fixTo_79_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_80 (
    .din     (_zz_481[31:0]        ), //i
    .dout    (fixTo_80_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_81 (
    .din     (_zz_482[31:0]        ), //i
    .dout    (fixTo_81_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_82 (
    .din     (_zz_483[31:0]        ), //i
    .dout    (fixTo_82_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_83 (
    .din     (_zz_484[31:0]        ), //i
    .dout    (fixTo_83_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_84 (
    .din     (_zz_485[31:0]        ), //i
    .dout    (fixTo_84_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_85 (
    .din     (_zz_486[31:0]        ), //i
    .dout    (fixTo_85_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_86 (
    .din     (_zz_487[31:0]        ), //i
    .dout    (fixTo_86_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_87 (
    .din     (_zz_488[31:0]        ), //i
    .dout    (fixTo_87_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_88 (
    .din     (_zz_489[31:0]        ), //i
    .dout    (fixTo_88_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_89 (
    .din     (_zz_490[31:0]        ), //i
    .dout    (fixTo_89_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_90 (
    .din     (_zz_491[31:0]        ), //i
    .dout    (fixTo_90_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_91 (
    .din     (_zz_492[31:0]        ), //i
    .dout    (fixTo_91_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_92 (
    .din     (_zz_493[31:0]        ), //i
    .dout    (fixTo_92_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_93 (
    .din     (_zz_494[31:0]        ), //i
    .dout    (fixTo_93_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_94 (
    .din     (_zz_495[31:0]        ), //i
    .dout    (fixTo_94_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_95 (
    .din     (_zz_496[31:0]        ), //i
    .dout    (fixTo_95_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_96 (
    .din     (_zz_497[31:0]        ), //i
    .dout    (fixTo_96_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_97 (
    .din     (_zz_498[31:0]        ), //i
    .dout    (fixTo_97_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_98 (
    .din     (_zz_499[31:0]        ), //i
    .dout    (fixTo_98_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_99 (
    .din     (_zz_500[31:0]        ), //i
    .dout    (fixTo_99_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_100 (
    .din     (_zz_501[31:0]         ), //i
    .dout    (fixTo_100_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_101 (
    .din     (_zz_502[31:0]         ), //i
    .dout    (fixTo_101_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_102 (
    .din     (_zz_503[31:0]         ), //i
    .dout    (fixTo_102_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_103 (
    .din     (_zz_504[31:0]         ), //i
    .dout    (fixTo_103_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_104 (
    .din     (_zz_505[31:0]         ), //i
    .dout    (fixTo_104_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_105 (
    .din     (_zz_506[31:0]         ), //i
    .dout    (fixTo_105_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_106 (
    .din     (_zz_507[31:0]         ), //i
    .dout    (fixTo_106_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_107 (
    .din     (_zz_508[31:0]         ), //i
    .dout    (fixTo_107_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_108 (
    .din     (_zz_509[31:0]         ), //i
    .dout    (fixTo_108_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_109 (
    .din     (_zz_510[31:0]         ), //i
    .dout    (fixTo_109_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_110 (
    .din     (_zz_511[31:0]         ), //i
    .dout    (fixTo_110_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_111 (
    .din     (_zz_512[31:0]         ), //i
    .dout    (fixTo_111_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_112 (
    .din     (_zz_513[31:0]         ), //i
    .dout    (fixTo_112_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_113 (
    .din     (_zz_514[31:0]         ), //i
    .dout    (fixTo_113_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_114 (
    .din     (_zz_515[31:0]         ), //i
    .dout    (fixTo_114_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_115 (
    .din     (_zz_516[31:0]         ), //i
    .dout    (fixTo_115_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_116 (
    .din     (_zz_517[31:0]         ), //i
    .dout    (fixTo_116_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_117 (
    .din     (_zz_518[31:0]         ), //i
    .dout    (fixTo_117_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_118 (
    .din     (_zz_519[31:0]         ), //i
    .dout    (fixTo_118_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_119 (
    .din     (_zz_520[31:0]         ), //i
    .dout    (fixTo_119_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_120 (
    .din     (_zz_521[31:0]         ), //i
    .dout    (fixTo_120_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_121 (
    .din     (_zz_522[31:0]         ), //i
    .dout    (fixTo_121_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_122 (
    .din     (_zz_523[31:0]         ), //i
    .dout    (fixTo_122_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_123 (
    .din     (_zz_524[31:0]         ), //i
    .dout    (fixTo_123_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_124 (
    .din     (_zz_525[31:0]         ), //i
    .dout    (fixTo_124_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_125 (
    .din     (_zz_526[31:0]         ), //i
    .dout    (fixTo_125_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_126 (
    .din     (_zz_527[31:0]         ), //i
    .dout    (fixTo_126_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_127 (
    .din     (_zz_528[31:0]         ), //i
    .dout    (fixTo_127_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_128 (
    .din     (_zz_529[31:0]         ), //i
    .dout    (fixTo_128_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_129 (
    .din     (_zz_530[31:0]         ), //i
    .dout    (fixTo_129_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_130 (
    .din     (_zz_531[31:0]         ), //i
    .dout    (fixTo_130_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_131 (
    .din     (_zz_532[31:0]         ), //i
    .dout    (fixTo_131_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_132 (
    .din     (_zz_533[31:0]         ), //i
    .dout    (fixTo_132_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_133 (
    .din     (_zz_534[31:0]         ), //i
    .dout    (fixTo_133_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_134 (
    .din     (_zz_535[31:0]         ), //i
    .dout    (fixTo_134_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_135 (
    .din     (_zz_536[31:0]         ), //i
    .dout    (fixTo_135_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_136 (
    .din     (_zz_537[31:0]         ), //i
    .dout    (fixTo_136_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_137 (
    .din     (_zz_538[31:0]         ), //i
    .dout    (fixTo_137_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_138 (
    .din     (_zz_539[31:0]         ), //i
    .dout    (fixTo_138_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_139 (
    .din     (_zz_540[31:0]         ), //i
    .dout    (fixTo_139_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_140 (
    .din     (_zz_541[31:0]         ), //i
    .dout    (fixTo_140_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_141 (
    .din     (_zz_542[31:0]         ), //i
    .dout    (fixTo_141_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_142 (
    .din     (_zz_543[31:0]         ), //i
    .dout    (fixTo_142_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_143 (
    .din     (_zz_544[31:0]         ), //i
    .dout    (fixTo_143_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_144 (
    .din     (_zz_545[31:0]         ), //i
    .dout    (fixTo_144_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_145 (
    .din     (_zz_546[31:0]         ), //i
    .dout    (fixTo_145_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_146 (
    .din     (_zz_547[31:0]         ), //i
    .dout    (fixTo_146_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_147 (
    .din     (_zz_548[31:0]         ), //i
    .dout    (fixTo_147_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_148 (
    .din     (_zz_549[31:0]         ), //i
    .dout    (fixTo_148_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_149 (
    .din     (_zz_550[31:0]         ), //i
    .dout    (fixTo_149_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_150 (
    .din     (_zz_551[31:0]         ), //i
    .dout    (fixTo_150_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_151 (
    .din     (_zz_552[31:0]         ), //i
    .dout    (fixTo_151_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_152 (
    .din     (_zz_553[31:0]         ), //i
    .dout    (fixTo_152_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_153 (
    .din     (_zz_554[31:0]         ), //i
    .dout    (fixTo_153_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_154 (
    .din     (_zz_555[31:0]         ), //i
    .dout    (fixTo_154_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_155 (
    .din     (_zz_556[31:0]         ), //i
    .dout    (fixTo_155_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_156 (
    .din     (_zz_557[31:0]         ), //i
    .dout    (fixTo_156_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_157 (
    .din     (_zz_558[31:0]         ), //i
    .dout    (fixTo_157_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_158 (
    .din     (_zz_559[31:0]         ), //i
    .dout    (fixTo_158_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_159 (
    .din     (_zz_560[31:0]         ), //i
    .dout    (fixTo_159_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_160 (
    .din     (_zz_561[31:0]         ), //i
    .dout    (fixTo_160_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_161 (
    .din     (_zz_562[31:0]         ), //i
    .dout    (fixTo_161_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_162 (
    .din     (_zz_563[31:0]         ), //i
    .dout    (fixTo_162_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_163 (
    .din     (_zz_564[31:0]         ), //i
    .dout    (fixTo_163_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_164 (
    .din     (_zz_565[31:0]         ), //i
    .dout    (fixTo_164_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_165 (
    .din     (_zz_566[31:0]         ), //i
    .dout    (fixTo_165_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_166 (
    .din     (_zz_567[31:0]         ), //i
    .dout    (fixTo_166_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_167 (
    .din     (_zz_568[31:0]         ), //i
    .dout    (fixTo_167_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_168 (
    .din     (_zz_569[31:0]         ), //i
    .dout    (fixTo_168_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_169 (
    .din     (_zz_570[31:0]         ), //i
    .dout    (fixTo_169_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_170 (
    .din     (_zz_571[31:0]         ), //i
    .dout    (fixTo_170_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_171 (
    .din     (_zz_572[31:0]         ), //i
    .dout    (fixTo_171_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_172 (
    .din     (_zz_573[31:0]         ), //i
    .dout    (fixTo_172_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_173 (
    .din     (_zz_574[31:0]         ), //i
    .dout    (fixTo_173_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_174 (
    .din     (_zz_575[31:0]         ), //i
    .dout    (fixTo_174_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_175 (
    .din     (_zz_576[31:0]         ), //i
    .dout    (fixTo_175_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_176 (
    .din     (_zz_577[31:0]         ), //i
    .dout    (fixTo_176_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_177 (
    .din     (_zz_578[31:0]         ), //i
    .dout    (fixTo_177_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_178 (
    .din     (_zz_579[31:0]         ), //i
    .dout    (fixTo_178_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_179 (
    .din     (_zz_580[31:0]         ), //i
    .dout    (fixTo_179_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_180 (
    .din     (_zz_581[31:0]         ), //i
    .dout    (fixTo_180_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_181 (
    .din     (_zz_582[31:0]         ), //i
    .dout    (fixTo_181_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_182 (
    .din     (_zz_583[31:0]         ), //i
    .dout    (fixTo_182_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_183 (
    .din     (_zz_584[31:0]         ), //i
    .dout    (fixTo_183_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_184 (
    .din     (_zz_585[31:0]         ), //i
    .dout    (fixTo_184_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_185 (
    .din     (_zz_586[31:0]         ), //i
    .dout    (fixTo_185_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_186 (
    .din     (_zz_587[31:0]         ), //i
    .dout    (fixTo_186_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_187 (
    .din     (_zz_588[31:0]         ), //i
    .dout    (fixTo_187_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_188 (
    .din     (_zz_589[31:0]         ), //i
    .dout    (fixTo_188_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_189 (
    .din     (_zz_590[31:0]         ), //i
    .dout    (fixTo_189_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_190 (
    .din     (_zz_591[31:0]         ), //i
    .dout    (fixTo_190_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_191 (
    .din     (_zz_592[31:0]         ), //i
    .dout    (fixTo_191_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_192 (
    .din     (_zz_593[31:0]         ), //i
    .dout    (fixTo_192_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_193 (
    .din     (_zz_594[31:0]         ), //i
    .dout    (fixTo_193_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_194 (
    .din     (_zz_595[31:0]         ), //i
    .dout    (fixTo_194_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_195 (
    .din     (_zz_596[31:0]         ), //i
    .dout    (fixTo_195_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_196 (
    .din     (_zz_597[31:0]         ), //i
    .dout    (fixTo_196_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_197 (
    .din     (_zz_598[31:0]         ), //i
    .dout    (fixTo_197_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_198 (
    .din     (_zz_599[31:0]         ), //i
    .dout    (fixTo_198_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_199 (
    .din     (_zz_600[31:0]         ), //i
    .dout    (fixTo_199_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_200 (
    .din     (_zz_601[31:0]         ), //i
    .dout    (fixTo_200_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_201 (
    .din     (_zz_602[31:0]         ), //i
    .dout    (fixTo_201_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_202 (
    .din     (_zz_603[31:0]         ), //i
    .dout    (fixTo_202_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_203 (
    .din     (_zz_604[31:0]         ), //i
    .dout    (fixTo_203_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_204 (
    .din     (_zz_605[31:0]         ), //i
    .dout    (fixTo_204_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_205 (
    .din     (_zz_606[31:0]         ), //i
    .dout    (fixTo_205_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_206 (
    .din     (_zz_607[31:0]         ), //i
    .dout    (fixTo_206_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_207 (
    .din     (_zz_608[31:0]         ), //i
    .dout    (fixTo_207_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_208 (
    .din     (_zz_609[31:0]         ), //i
    .dout    (fixTo_208_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_209 (
    .din     (_zz_610[31:0]         ), //i
    .dout    (fixTo_209_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_210 (
    .din     (_zz_611[31:0]         ), //i
    .dout    (fixTo_210_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_211 (
    .din     (_zz_612[31:0]         ), //i
    .dout    (fixTo_211_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_212 (
    .din     (_zz_613[31:0]         ), //i
    .dout    (fixTo_212_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_213 (
    .din     (_zz_614[31:0]         ), //i
    .dout    (fixTo_213_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_214 (
    .din     (_zz_615[31:0]         ), //i
    .dout    (fixTo_214_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_215 (
    .din     (_zz_616[31:0]         ), //i
    .dout    (fixTo_215_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_216 (
    .din     (_zz_617[31:0]         ), //i
    .dout    (fixTo_216_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_217 (
    .din     (_zz_618[31:0]         ), //i
    .dout    (fixTo_217_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_218 (
    .din     (_zz_619[31:0]         ), //i
    .dout    (fixTo_218_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_219 (
    .din     (_zz_620[31:0]         ), //i
    .dout    (fixTo_219_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_220 (
    .din     (_zz_621[31:0]         ), //i
    .dout    (fixTo_220_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_221 (
    .din     (_zz_622[31:0]         ), //i
    .dout    (fixTo_221_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_222 (
    .din     (_zz_623[31:0]         ), //i
    .dout    (fixTo_222_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_223 (
    .din     (_zz_624[31:0]         ), //i
    .dout    (fixTo_223_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_224 (
    .din     (_zz_625[31:0]         ), //i
    .dout    (fixTo_224_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_225 (
    .din     (_zz_626[31:0]         ), //i
    .dout    (fixTo_225_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_226 (
    .din     (_zz_627[31:0]         ), //i
    .dout    (fixTo_226_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_227 (
    .din     (_zz_628[31:0]         ), //i
    .dout    (fixTo_227_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_228 (
    .din     (_zz_629[31:0]         ), //i
    .dout    (fixTo_228_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_229 (
    .din     (_zz_630[31:0]         ), //i
    .dout    (fixTo_229_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_230 (
    .din     (_zz_631[31:0]         ), //i
    .dout    (fixTo_230_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_231 (
    .din     (_zz_632[31:0]         ), //i
    .dout    (fixTo_231_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_232 (
    .din     (_zz_633[31:0]         ), //i
    .dout    (fixTo_232_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_233 (
    .din     (_zz_634[31:0]         ), //i
    .dout    (fixTo_233_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_234 (
    .din     (_zz_635[31:0]         ), //i
    .dout    (fixTo_234_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_235 (
    .din     (_zz_636[31:0]         ), //i
    .dout    (fixTo_235_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_236 (
    .din     (_zz_637[31:0]         ), //i
    .dout    (fixTo_236_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_237 (
    .din     (_zz_638[31:0]         ), //i
    .dout    (fixTo_237_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_238 (
    .din     (_zz_639[31:0]         ), //i
    .dout    (fixTo_238_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_239 (
    .din     (_zz_640[31:0]         ), //i
    .dout    (fixTo_239_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_240 (
    .din     (_zz_641[31:0]         ), //i
    .dout    (fixTo_240_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_241 (
    .din     (_zz_642[31:0]         ), //i
    .dout    (fixTo_241_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_242 (
    .din     (_zz_643[31:0]         ), //i
    .dout    (fixTo_242_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_243 (
    .din     (_zz_644[31:0]         ), //i
    .dout    (fixTo_243_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_244 (
    .din     (_zz_645[31:0]         ), //i
    .dout    (fixTo_244_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_245 (
    .din     (_zz_646[31:0]         ), //i
    .dout    (fixTo_245_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_246 (
    .din     (_zz_647[31:0]         ), //i
    .dout    (fixTo_246_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_247 (
    .din     (_zz_648[31:0]         ), //i
    .dout    (fixTo_247_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_248 (
    .din     (_zz_649[31:0]         ), //i
    .dout    (fixTo_248_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_249 (
    .din     (_zz_650[31:0]         ), //i
    .dout    (fixTo_249_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_250 (
    .din     (_zz_651[31:0]         ), //i
    .dout    (fixTo_250_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_251 (
    .din     (_zz_652[31:0]         ), //i
    .dout    (fixTo_251_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_252 (
    .din     (_zz_653[31:0]         ), //i
    .dout    (fixTo_252_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_253 (
    .din     (_zz_654[31:0]         ), //i
    .dout    (fixTo_253_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_254 (
    .din     (_zz_655[31:0]         ), //i
    .dout    (fixTo_254_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_255 (
    .din     (_zz_656[31:0]         ), //i
    .dout    (fixTo_255_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_256 (
    .din     (_zz_657[31:0]         ), //i
    .dout    (fixTo_256_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_257 (
    .din     (_zz_658[31:0]         ), //i
    .dout    (fixTo_257_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_258 (
    .din     (_zz_659[31:0]         ), //i
    .dout    (fixTo_258_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_259 (
    .din     (_zz_660[31:0]         ), //i
    .dout    (fixTo_259_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_260 (
    .din     (_zz_661[31:0]         ), //i
    .dout    (fixTo_260_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_261 (
    .din     (_zz_662[31:0]         ), //i
    .dout    (fixTo_261_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_262 (
    .din     (_zz_663[31:0]         ), //i
    .dout    (fixTo_262_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_263 (
    .din     (_zz_664[31:0]         ), //i
    .dout    (fixTo_263_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_264 (
    .din     (_zz_665[31:0]         ), //i
    .dout    (fixTo_264_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_265 (
    .din     (_zz_666[31:0]         ), //i
    .dout    (fixTo_265_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_266 (
    .din     (_zz_667[31:0]         ), //i
    .dout    (fixTo_266_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_267 (
    .din     (_zz_668[31:0]         ), //i
    .dout    (fixTo_267_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_268 (
    .din     (_zz_669[31:0]         ), //i
    .dout    (fixTo_268_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_269 (
    .din     (_zz_670[31:0]         ), //i
    .dout    (fixTo_269_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_270 (
    .din     (_zz_671[31:0]         ), //i
    .dout    (fixTo_270_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_271 (
    .din     (_zz_672[31:0]         ), //i
    .dout    (fixTo_271_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_272 (
    .din     (_zz_673[31:0]         ), //i
    .dout    (fixTo_272_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_273 (
    .din     (_zz_674[31:0]         ), //i
    .dout    (fixTo_273_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_274 (
    .din     (_zz_675[31:0]         ), //i
    .dout    (fixTo_274_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_275 (
    .din     (_zz_676[31:0]         ), //i
    .dout    (fixTo_275_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_276 (
    .din     (_zz_677[31:0]         ), //i
    .dout    (fixTo_276_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_277 (
    .din     (_zz_678[31:0]         ), //i
    .dout    (fixTo_277_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_278 (
    .din     (_zz_679[31:0]         ), //i
    .dout    (fixTo_278_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_279 (
    .din     (_zz_680[31:0]         ), //i
    .dout    (fixTo_279_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_280 (
    .din     (_zz_681[31:0]         ), //i
    .dout    (fixTo_280_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_281 (
    .din     (_zz_682[31:0]         ), //i
    .dout    (fixTo_281_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_282 (
    .din     (_zz_683[31:0]         ), //i
    .dout    (fixTo_282_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_283 (
    .din     (_zz_684[31:0]         ), //i
    .dout    (fixTo_283_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_284 (
    .din     (_zz_685[31:0]         ), //i
    .dout    (fixTo_284_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_285 (
    .din     (_zz_686[31:0]         ), //i
    .dout    (fixTo_285_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_286 (
    .din     (_zz_687[31:0]         ), //i
    .dout    (fixTo_286_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_287 (
    .din     (_zz_688[31:0]         ), //i
    .dout    (fixTo_287_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_288 (
    .din     (_zz_689[31:0]         ), //i
    .dout    (fixTo_288_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_289 (
    .din     (_zz_690[31:0]         ), //i
    .dout    (fixTo_289_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_290 (
    .din     (_zz_691[31:0]         ), //i
    .dout    (fixTo_290_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_291 (
    .din     (_zz_692[31:0]         ), //i
    .dout    (fixTo_291_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_292 (
    .din     (_zz_693[31:0]         ), //i
    .dout    (fixTo_292_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_293 (
    .din     (_zz_694[31:0]         ), //i
    .dout    (fixTo_293_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_294 (
    .din     (_zz_695[31:0]         ), //i
    .dout    (fixTo_294_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_295 (
    .din     (_zz_696[31:0]         ), //i
    .dout    (fixTo_295_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_296 (
    .din     (_zz_697[31:0]         ), //i
    .dout    (fixTo_296_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_297 (
    .din     (_zz_698[31:0]         ), //i
    .dout    (fixTo_297_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_298 (
    .din     (_zz_699[31:0]         ), //i
    .dout    (fixTo_298_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_299 (
    .din     (_zz_700[31:0]         ), //i
    .dout    (fixTo_299_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_300 (
    .din     (_zz_701[31:0]         ), //i
    .dout    (fixTo_300_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_301 (
    .din     (_zz_702[31:0]         ), //i
    .dout    (fixTo_301_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_302 (
    .din     (_zz_703[31:0]         ), //i
    .dout    (fixTo_302_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_303 (
    .din     (_zz_704[31:0]         ), //i
    .dout    (fixTo_303_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_304 (
    .din     (_zz_705[31:0]         ), //i
    .dout    (fixTo_304_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_305 (
    .din     (_zz_706[31:0]         ), //i
    .dout    (fixTo_305_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_306 (
    .din     (_zz_707[31:0]         ), //i
    .dout    (fixTo_306_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_307 (
    .din     (_zz_708[31:0]         ), //i
    .dout    (fixTo_307_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_308 (
    .din     (_zz_709[31:0]         ), //i
    .dout    (fixTo_308_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_309 (
    .din     (_zz_710[31:0]         ), //i
    .dout    (fixTo_309_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_310 (
    .din     (_zz_711[31:0]         ), //i
    .dout    (fixTo_310_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_311 (
    .din     (_zz_712[31:0]         ), //i
    .dout    (fixTo_311_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_312 (
    .din     (_zz_713[31:0]         ), //i
    .dout    (fixTo_312_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_313 (
    .din     (_zz_714[31:0]         ), //i
    .dout    (fixTo_313_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_314 (
    .din     (_zz_715[31:0]         ), //i
    .dout    (fixTo_314_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_315 (
    .din     (_zz_716[31:0]         ), //i
    .dout    (fixTo_315_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_316 (
    .din     (_zz_717[31:0]         ), //i
    .dout    (fixTo_316_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_317 (
    .din     (_zz_718[31:0]         ), //i
    .dout    (fixTo_317_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_318 (
    .din     (_zz_719[31:0]         ), //i
    .dout    (fixTo_318_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_319 (
    .din     (_zz_720[31:0]         ), //i
    .dout    (fixTo_319_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_320 (
    .din     (_zz_721[31:0]         ), //i
    .dout    (fixTo_320_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_321 (
    .din     (_zz_722[31:0]         ), //i
    .dout    (fixTo_321_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_322 (
    .din     (_zz_723[31:0]         ), //i
    .dout    (fixTo_322_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_323 (
    .din     (_zz_724[31:0]         ), //i
    .dout    (fixTo_323_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_324 (
    .din     (_zz_725[31:0]         ), //i
    .dout    (fixTo_324_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_325 (
    .din     (_zz_726[31:0]         ), //i
    .dout    (fixTo_325_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_326 (
    .din     (_zz_727[31:0]         ), //i
    .dout    (fixTo_326_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_327 (
    .din     (_zz_728[31:0]         ), //i
    .dout    (fixTo_327_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_328 (
    .din     (_zz_729[31:0]         ), //i
    .dout    (fixTo_328_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_329 (
    .din     (_zz_730[31:0]         ), //i
    .dout    (fixTo_329_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_330 (
    .din     (_zz_731[31:0]         ), //i
    .dout    (fixTo_330_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_331 (
    .din     (_zz_732[31:0]         ), //i
    .dout    (fixTo_331_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_332 (
    .din     (_zz_733[31:0]         ), //i
    .dout    (fixTo_332_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_333 (
    .din     (_zz_734[31:0]         ), //i
    .dout    (fixTo_333_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_334 (
    .din     (_zz_735[31:0]         ), //i
    .dout    (fixTo_334_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_335 (
    .din     (_zz_736[31:0]         ), //i
    .dout    (fixTo_335_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_336 (
    .din     (_zz_737[31:0]         ), //i
    .dout    (fixTo_336_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_337 (
    .din     (_zz_738[31:0]         ), //i
    .dout    (fixTo_337_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_338 (
    .din     (_zz_739[31:0]         ), //i
    .dout    (fixTo_338_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_339 (
    .din     (_zz_740[31:0]         ), //i
    .dout    (fixTo_339_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_340 (
    .din     (_zz_741[31:0]         ), //i
    .dout    (fixTo_340_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_341 (
    .din     (_zz_742[31:0]         ), //i
    .dout    (fixTo_341_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_342 (
    .din     (_zz_743[31:0]         ), //i
    .dout    (fixTo_342_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_343 (
    .din     (_zz_744[31:0]         ), //i
    .dout    (fixTo_343_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_344 (
    .din     (_zz_745[31:0]         ), //i
    .dout    (fixTo_344_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_345 (
    .din     (_zz_746[31:0]         ), //i
    .dout    (fixTo_345_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_346 (
    .din     (_zz_747[31:0]         ), //i
    .dout    (fixTo_346_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_347 (
    .din     (_zz_748[31:0]         ), //i
    .dout    (fixTo_347_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_348 (
    .din     (_zz_749[31:0]         ), //i
    .dout    (fixTo_348_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_349 (
    .din     (_zz_750[31:0]         ), //i
    .dout    (fixTo_349_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_350 (
    .din     (_zz_751[31:0]         ), //i
    .dout    (fixTo_350_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_351 (
    .din     (_zz_752[31:0]         ), //i
    .dout    (fixTo_351_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_352 (
    .din     (_zz_753[31:0]         ), //i
    .dout    (fixTo_352_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_353 (
    .din     (_zz_754[31:0]         ), //i
    .dout    (fixTo_353_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_354 (
    .din     (_zz_755[31:0]         ), //i
    .dout    (fixTo_354_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_355 (
    .din     (_zz_756[31:0]         ), //i
    .dout    (fixTo_355_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_356 (
    .din     (_zz_757[31:0]         ), //i
    .dout    (fixTo_356_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_357 (
    .din     (_zz_758[31:0]         ), //i
    .dout    (fixTo_357_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_358 (
    .din     (_zz_759[31:0]         ), //i
    .dout    (fixTo_358_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_359 (
    .din     (_zz_760[31:0]         ), //i
    .dout    (fixTo_359_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_360 (
    .din     (_zz_761[31:0]         ), //i
    .dout    (fixTo_360_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_361 (
    .din     (_zz_762[31:0]         ), //i
    .dout    (fixTo_361_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_362 (
    .din     (_zz_763[31:0]         ), //i
    .dout    (fixTo_362_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_363 (
    .din     (_zz_764[31:0]         ), //i
    .dout    (fixTo_363_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_364 (
    .din     (_zz_765[31:0]         ), //i
    .dout    (fixTo_364_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_365 (
    .din     (_zz_766[31:0]         ), //i
    .dout    (fixTo_365_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_366 (
    .din     (_zz_767[31:0]         ), //i
    .dout    (fixTo_366_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_367 (
    .din     (_zz_768[31:0]         ), //i
    .dout    (fixTo_367_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_368 (
    .din     (_zz_769[31:0]         ), //i
    .dout    (fixTo_368_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_369 (
    .din     (_zz_770[31:0]         ), //i
    .dout    (fixTo_369_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_370 (
    .din     (_zz_771[31:0]         ), //i
    .dout    (fixTo_370_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_371 (
    .din     (_zz_772[31:0]         ), //i
    .dout    (fixTo_371_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_372 (
    .din     (_zz_773[31:0]         ), //i
    .dout    (fixTo_372_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_373 (
    .din     (_zz_774[31:0]         ), //i
    .dout    (fixTo_373_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_374 (
    .din     (_zz_775[31:0]         ), //i
    .dout    (fixTo_374_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_375 (
    .din     (_zz_776[31:0]         ), //i
    .dout    (fixTo_375_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_376 (
    .din     (_zz_777[31:0]         ), //i
    .dout    (fixTo_376_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_377 (
    .din     (_zz_778[31:0]         ), //i
    .dout    (fixTo_377_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_378 (
    .din     (_zz_779[31:0]         ), //i
    .dout    (fixTo_378_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_379 (
    .din     (_zz_780[31:0]         ), //i
    .dout    (fixTo_379_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_380 (
    .din     (_zz_781[31:0]         ), //i
    .dout    (fixTo_380_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_381 (
    .din     (_zz_782[31:0]         ), //i
    .dout    (fixTo_381_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_382 (
    .din     (_zz_783[31:0]         ), //i
    .dout    (fixTo_382_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_383 (
    .din     (_zz_784[31:0]         ), //i
    .dout    (fixTo_383_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_384 (
    .din     (_zz_785[31:0]         ), //i
    .dout    (fixTo_384_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_385 (
    .din     (_zz_786[31:0]         ), //i
    .dout    (fixTo_385_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_386 (
    .din     (_zz_787[31:0]         ), //i
    .dout    (fixTo_386_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_387 (
    .din     (_zz_788[31:0]         ), //i
    .dout    (fixTo_387_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_388 (
    .din     (_zz_789[31:0]         ), //i
    .dout    (fixTo_388_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_389 (
    .din     (_zz_790[31:0]         ), //i
    .dout    (fixTo_389_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_390 (
    .din     (_zz_791[31:0]         ), //i
    .dout    (fixTo_390_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_391 (
    .din     (_zz_792[31:0]         ), //i
    .dout    (fixTo_391_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_392 (
    .din     (_zz_793[31:0]         ), //i
    .dout    (fixTo_392_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_393 (
    .din     (_zz_794[31:0]         ), //i
    .dout    (fixTo_393_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_394 (
    .din     (_zz_795[31:0]         ), //i
    .dout    (fixTo_394_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_395 (
    .din     (_zz_796[31:0]         ), //i
    .dout    (fixTo_395_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_396 (
    .din     (_zz_797[31:0]         ), //i
    .dout    (fixTo_396_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_397 (
    .din     (_zz_798[31:0]         ), //i
    .dout    (fixTo_397_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_398 (
    .din     (_zz_799[31:0]         ), //i
    .dout    (fixTo_398_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_399 (
    .din     (_zz_800[31:0]         ), //i
    .dout    (fixTo_399_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_400 (
    .din     (_zz_801[31:0]         ), //i
    .dout    (fixTo_400_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_401 (
    .din     (_zz_802[31:0]         ), //i
    .dout    (fixTo_401_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_402 (
    .din     (_zz_803[31:0]         ), //i
    .dout    (fixTo_402_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_403 (
    .din     (_zz_804[31:0]         ), //i
    .dout    (fixTo_403_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_404 (
    .din     (_zz_805[31:0]         ), //i
    .dout    (fixTo_404_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_405 (
    .din     (_zz_806[31:0]         ), //i
    .dout    (fixTo_405_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_406 (
    .din     (_zz_807[31:0]         ), //i
    .dout    (fixTo_406_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_407 (
    .din     (_zz_808[31:0]         ), //i
    .dout    (fixTo_407_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_408 (
    .din     (_zz_809[31:0]         ), //i
    .dout    (fixTo_408_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_409 (
    .din     (_zz_810[31:0]         ), //i
    .dout    (fixTo_409_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_410 (
    .din     (_zz_811[31:0]         ), //i
    .dout    (fixTo_410_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_411 (
    .din     (_zz_812[31:0]         ), //i
    .dout    (fixTo_411_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_412 (
    .din     (_zz_813[31:0]         ), //i
    .dout    (fixTo_412_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_413 (
    .din     (_zz_814[31:0]         ), //i
    .dout    (fixTo_413_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_414 (
    .din     (_zz_815[31:0]         ), //i
    .dout    (fixTo_414_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_415 (
    .din     (_zz_816[31:0]         ), //i
    .dout    (fixTo_415_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_416 (
    .din     (_zz_817[31:0]         ), //i
    .dout    (fixTo_416_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_417 (
    .din     (_zz_818[31:0]         ), //i
    .dout    (fixTo_417_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_418 (
    .din     (_zz_819[31:0]         ), //i
    .dout    (fixTo_418_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_419 (
    .din     (_zz_820[31:0]         ), //i
    .dout    (fixTo_419_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_420 (
    .din     (_zz_821[31:0]         ), //i
    .dout    (fixTo_420_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_421 (
    .din     (_zz_822[31:0]         ), //i
    .dout    (fixTo_421_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_422 (
    .din     (_zz_823[31:0]         ), //i
    .dout    (fixTo_422_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_423 (
    .din     (_zz_824[31:0]         ), //i
    .dout    (fixTo_423_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_424 (
    .din     (_zz_825[31:0]         ), //i
    .dout    (fixTo_424_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_425 (
    .din     (_zz_826[31:0]         ), //i
    .dout    (fixTo_425_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_426 (
    .din     (_zz_827[31:0]         ), //i
    .dout    (fixTo_426_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_427 (
    .din     (_zz_828[31:0]         ), //i
    .dout    (fixTo_427_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_428 (
    .din     (_zz_829[31:0]         ), //i
    .dout    (fixTo_428_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_429 (
    .din     (_zz_830[31:0]         ), //i
    .dout    (fixTo_429_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_430 (
    .din     (_zz_831[31:0]         ), //i
    .dout    (fixTo_430_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_431 (
    .din     (_zz_832[31:0]         ), //i
    .dout    (fixTo_431_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_432 (
    .din     (_zz_833[31:0]         ), //i
    .dout    (fixTo_432_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_433 (
    .din     (_zz_834[31:0]         ), //i
    .dout    (fixTo_433_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_434 (
    .din     (_zz_835[31:0]         ), //i
    .dout    (fixTo_434_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_435 (
    .din     (_zz_836[31:0]         ), //i
    .dout    (fixTo_435_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_436 (
    .din     (_zz_837[31:0]         ), //i
    .dout    (fixTo_436_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_437 (
    .din     (_zz_838[31:0]         ), //i
    .dout    (fixTo_437_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_438 (
    .din     (_zz_839[31:0]         ), //i
    .dout    (fixTo_438_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_439 (
    .din     (_zz_840[31:0]         ), //i
    .dout    (fixTo_439_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_440 (
    .din     (_zz_841[31:0]         ), //i
    .dout    (fixTo_440_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_441 (
    .din     (_zz_842[31:0]         ), //i
    .dout    (fixTo_441_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_442 (
    .din     (_zz_843[31:0]         ), //i
    .dout    (fixTo_442_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_443 (
    .din     (_zz_844[31:0]         ), //i
    .dout    (fixTo_443_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_444 (
    .din     (_zz_845[31:0]         ), //i
    .dout    (fixTo_444_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_445 (
    .din     (_zz_846[31:0]         ), //i
    .dout    (fixTo_445_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_446 (
    .din     (_zz_847[31:0]         ), //i
    .dout    (fixTo_446_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_447 (
    .din     (_zz_848[31:0]         ), //i
    .dout    (fixTo_447_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_448 (
    .din     (_zz_849[31:0]         ), //i
    .dout    (fixTo_448_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_449 (
    .din     (_zz_850[31:0]         ), //i
    .dout    (fixTo_449_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_450 (
    .din     (_zz_851[31:0]         ), //i
    .dout    (fixTo_450_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_451 (
    .din     (_zz_852[31:0]         ), //i
    .dout    (fixTo_451_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_452 (
    .din     (_zz_853[31:0]         ), //i
    .dout    (fixTo_452_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_453 (
    .din     (_zz_854[31:0]         ), //i
    .dout    (fixTo_453_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_454 (
    .din     (_zz_855[31:0]         ), //i
    .dout    (fixTo_454_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_455 (
    .din     (_zz_856[31:0]         ), //i
    .dout    (fixTo_455_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_456 (
    .din     (_zz_857[31:0]         ), //i
    .dout    (fixTo_456_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_457 (
    .din     (_zz_858[31:0]         ), //i
    .dout    (fixTo_457_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_458 (
    .din     (_zz_859[31:0]         ), //i
    .dout    (fixTo_458_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_459 (
    .din     (_zz_860[31:0]         ), //i
    .dout    (fixTo_459_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_460 (
    .din     (_zz_861[31:0]         ), //i
    .dout    (fixTo_460_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_461 (
    .din     (_zz_862[31:0]         ), //i
    .dout    (fixTo_461_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_462 (
    .din     (_zz_863[31:0]         ), //i
    .dout    (fixTo_462_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_463 (
    .din     (_zz_864[31:0]         ), //i
    .dout    (fixTo_463_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_464 (
    .din     (_zz_865[31:0]         ), //i
    .dout    (fixTo_464_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_465 (
    .din     (_zz_866[31:0]         ), //i
    .dout    (fixTo_465_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_466 (
    .din     (_zz_867[31:0]         ), //i
    .dout    (fixTo_466_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_467 (
    .din     (_zz_868[31:0]         ), //i
    .dout    (fixTo_467_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_468 (
    .din     (_zz_869[31:0]         ), //i
    .dout    (fixTo_468_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_469 (
    .din     (_zz_870[31:0]         ), //i
    .dout    (fixTo_469_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_470 (
    .din     (_zz_871[31:0]         ), //i
    .dout    (fixTo_470_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_471 (
    .din     (_zz_872[31:0]         ), //i
    .dout    (fixTo_471_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_472 (
    .din     (_zz_873[31:0]         ), //i
    .dout    (fixTo_472_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_473 (
    .din     (_zz_874[31:0]         ), //i
    .dout    (fixTo_473_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_474 (
    .din     (_zz_875[31:0]         ), //i
    .dout    (fixTo_474_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_475 (
    .din     (_zz_876[31:0]         ), //i
    .dout    (fixTo_475_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_476 (
    .din     (_zz_877[31:0]         ), //i
    .dout    (fixTo_476_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_477 (
    .din     (_zz_878[31:0]         ), //i
    .dout    (fixTo_477_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_478 (
    .din     (_zz_879[31:0]         ), //i
    .dout    (fixTo_478_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_479 (
    .din     (_zz_880[31:0]         ), //i
    .dout    (fixTo_479_dout[15:0]  )  //o
  );
  assign twiddle_factor_table_0_real = 16'h0100;
  assign twiddle_factor_table_0_imag = 16'h0;
  assign twiddle_factor_table_1_real = 16'h0100;
  assign twiddle_factor_table_1_imag = 16'h0;
  assign twiddle_factor_table_2_real = 16'h0;
  assign twiddle_factor_table_2_imag = 16'hff00;
  assign twiddle_factor_table_3_real = 16'h0100;
  assign twiddle_factor_table_3_imag = 16'h0;
  assign twiddle_factor_table_4_real = 16'h00b5;
  assign twiddle_factor_table_4_imag = 16'hff4b;
  assign twiddle_factor_table_5_real = 16'h0;
  assign twiddle_factor_table_5_imag = 16'hff00;
  assign twiddle_factor_table_6_real = 16'hff4b;
  assign twiddle_factor_table_6_imag = 16'hff4b;
  assign twiddle_factor_table_7_real = 16'h0100;
  assign twiddle_factor_table_7_imag = 16'h0;
  assign twiddle_factor_table_8_real = 16'h00ec;
  assign twiddle_factor_table_8_imag = 16'hff9f;
  assign twiddle_factor_table_9_real = 16'h00b5;
  assign twiddle_factor_table_9_imag = 16'hff4b;
  assign twiddle_factor_table_10_real = 16'h0061;
  assign twiddle_factor_table_10_imag = 16'hff14;
  assign twiddle_factor_table_11_real = 16'h0;
  assign twiddle_factor_table_11_imag = 16'hff00;
  assign twiddle_factor_table_12_real = 16'hff9f;
  assign twiddle_factor_table_12_imag = 16'hff14;
  assign twiddle_factor_table_13_real = 16'hff4b;
  assign twiddle_factor_table_13_imag = 16'hff4b;
  assign twiddle_factor_table_14_real = 16'hff14;
  assign twiddle_factor_table_14_imag = 16'hff9f;
  assign twiddle_factor_table_15_real = 16'h0100;
  assign twiddle_factor_table_15_imag = 16'h0;
  assign twiddle_factor_table_16_real = 16'h00fb;
  assign twiddle_factor_table_16_imag = 16'hffcf;
  assign twiddle_factor_table_17_real = 16'h00ec;
  assign twiddle_factor_table_17_imag = 16'hff9f;
  assign twiddle_factor_table_18_real = 16'h00d4;
  assign twiddle_factor_table_18_imag = 16'hff72;
  assign twiddle_factor_table_19_real = 16'h00b5;
  assign twiddle_factor_table_19_imag = 16'hff4b;
  assign twiddle_factor_table_20_real = 16'h008e;
  assign twiddle_factor_table_20_imag = 16'hff2c;
  assign twiddle_factor_table_21_real = 16'h0061;
  assign twiddle_factor_table_21_imag = 16'hff14;
  assign twiddle_factor_table_22_real = 16'h0031;
  assign twiddle_factor_table_22_imag = 16'hff05;
  assign twiddle_factor_table_23_real = 16'h0;
  assign twiddle_factor_table_23_imag = 16'hff00;
  assign twiddle_factor_table_24_real = 16'hffcf;
  assign twiddle_factor_table_24_imag = 16'hff05;
  assign twiddle_factor_table_25_real = 16'hff9f;
  assign twiddle_factor_table_25_imag = 16'hff14;
  assign twiddle_factor_table_26_real = 16'hff72;
  assign twiddle_factor_table_26_imag = 16'hff2c;
  assign twiddle_factor_table_27_real = 16'hff4b;
  assign twiddle_factor_table_27_imag = 16'hff4b;
  assign twiddle_factor_table_28_real = 16'hff2c;
  assign twiddle_factor_table_28_imag = 16'hff72;
  assign twiddle_factor_table_29_real = 16'hff14;
  assign twiddle_factor_table_29_imag = 16'hff9f;
  assign twiddle_factor_table_30_real = 16'hff05;
  assign twiddle_factor_table_30_imag = 16'hffcf;
  assign data_reorder_0_real = data_in_0_real;
  assign data_reorder_0_imag = data_in_0_imag;
  assign data_reorder_16_real = data_in_1_real;
  assign data_reorder_16_imag = data_in_1_imag;
  assign data_reorder_8_real = data_in_2_real;
  assign data_reorder_8_imag = data_in_2_imag;
  assign data_reorder_24_real = data_in_3_real;
  assign data_reorder_24_imag = data_in_3_imag;
  assign data_reorder_4_real = data_in_4_real;
  assign data_reorder_4_imag = data_in_4_imag;
  assign data_reorder_20_real = data_in_5_real;
  assign data_reorder_20_imag = data_in_5_imag;
  assign data_reorder_12_real = data_in_6_real;
  assign data_reorder_12_imag = data_in_6_imag;
  assign data_reorder_28_real = data_in_7_real;
  assign data_reorder_28_imag = data_in_7_imag;
  assign data_reorder_2_real = data_in_8_real;
  assign data_reorder_2_imag = data_in_8_imag;
  assign data_reorder_18_real = data_in_9_real;
  assign data_reorder_18_imag = data_in_9_imag;
  assign data_reorder_10_real = data_in_10_real;
  assign data_reorder_10_imag = data_in_10_imag;
  assign data_reorder_26_real = data_in_11_real;
  assign data_reorder_26_imag = data_in_11_imag;
  assign data_reorder_6_real = data_in_12_real;
  assign data_reorder_6_imag = data_in_12_imag;
  assign data_reorder_22_real = data_in_13_real;
  assign data_reorder_22_imag = data_in_13_imag;
  assign data_reorder_14_real = data_in_14_real;
  assign data_reorder_14_imag = data_in_14_imag;
  assign data_reorder_30_real = data_in_15_real;
  assign data_reorder_30_imag = data_in_15_imag;
  assign data_reorder_1_real = data_in_16_real;
  assign data_reorder_1_imag = data_in_16_imag;
  assign data_reorder_17_real = data_in_17_real;
  assign data_reorder_17_imag = data_in_17_imag;
  assign data_reorder_9_real = data_in_18_real;
  assign data_reorder_9_imag = data_in_18_imag;
  assign data_reorder_25_real = data_in_19_real;
  assign data_reorder_25_imag = data_in_19_imag;
  assign data_reorder_5_real = data_in_20_real;
  assign data_reorder_5_imag = data_in_20_imag;
  assign data_reorder_21_real = data_in_21_real;
  assign data_reorder_21_imag = data_in_21_imag;
  assign data_reorder_13_real = data_in_22_real;
  assign data_reorder_13_imag = data_in_22_imag;
  assign data_reorder_29_real = data_in_23_real;
  assign data_reorder_29_imag = data_in_23_imag;
  assign data_reorder_3_real = data_in_24_real;
  assign data_reorder_3_imag = data_in_24_imag;
  assign data_reorder_19_real = data_in_25_real;
  assign data_reorder_19_imag = data_in_25_imag;
  assign data_reorder_11_real = data_in_26_real;
  assign data_reorder_11_imag = data_in_26_imag;
  assign data_reorder_27_real = data_in_27_real;
  assign data_reorder_27_imag = data_in_27_imag;
  assign data_reorder_7_real = data_in_28_real;
  assign data_reorder_7_imag = data_in_28_imag;
  assign data_reorder_23_real = data_in_29_real;
  assign data_reorder_23_imag = data_in_29_imag;
  assign data_reorder_15_real = data_in_30_real;
  assign data_reorder_15_imag = data_in_30_imag;
  assign data_reorder_31_real = data_in_31_real;
  assign data_reorder_31_imag = data_in_31_imag;
  always @ (*) begin
    current_level_willIncrement = 1'b0;
    if(null_cond_period)begin
      current_level_willIncrement = 1'b1;
    end
  end

  assign current_level_willClear = 1'b0;
  assign current_level_willOverflowIfInc = (current_level_value == 3'b101);
  assign current_level_willOverflow = (current_level_willOverflowIfInc && current_level_willIncrement);
  always @ (*) begin
    if(current_level_willOverflow)begin
      current_level_valueNext = 3'b000;
    end else begin
      current_level_valueNext = (current_level_value + _zz_882);
    end
    if(current_level_willClear)begin
      current_level_valueNext = 3'b000;
    end
  end

  assign null_cond_period = (io_data_in_valid_regNext || null_cond_period_minus_1);
  assign _zz_3 = ($signed(_zz_883) * $signed(data_mid_1_real));
  assign _zz_401 = _zz_884;
  assign _zz_1 = _zz_887[31 : 0];
  assign _zz_402 = _zz_888;
  assign _zz_2 = _zz_891[31 : 0];
  assign _zz_4 = 1'b1;
  assign _zz_403 = _zz_892;
  assign _zz_404 = _zz_900;
  assign _zz_5 = 1'b1;
  assign _zz_405 = _zz_908;
  assign _zz_406 = _zz_916;
  assign _zz_8 = ($signed(_zz_924) * $signed(data_mid_3_real));
  assign _zz_407 = _zz_925;
  assign _zz_6 = _zz_928[31 : 0];
  assign _zz_408 = _zz_929;
  assign _zz_7 = _zz_932[31 : 0];
  assign _zz_9 = 1'b1;
  assign _zz_409 = _zz_933;
  assign _zz_410 = _zz_941;
  assign _zz_10 = 1'b1;
  assign _zz_411 = _zz_949;
  assign _zz_412 = _zz_957;
  assign _zz_13 = ($signed(_zz_965) * $signed(data_mid_5_real));
  assign _zz_413 = _zz_966;
  assign _zz_11 = _zz_969[31 : 0];
  assign _zz_414 = _zz_970;
  assign _zz_12 = _zz_973[31 : 0];
  assign _zz_14 = 1'b1;
  assign _zz_415 = _zz_974;
  assign _zz_416 = _zz_982;
  assign _zz_15 = 1'b1;
  assign _zz_417 = _zz_990;
  assign _zz_418 = _zz_998;
  assign _zz_18 = ($signed(_zz_1006) * $signed(data_mid_7_real));
  assign _zz_419 = _zz_1007;
  assign _zz_16 = _zz_1010[31 : 0];
  assign _zz_420 = _zz_1011;
  assign _zz_17 = _zz_1014[31 : 0];
  assign _zz_19 = 1'b1;
  assign _zz_421 = _zz_1015;
  assign _zz_422 = _zz_1023;
  assign _zz_20 = 1'b1;
  assign _zz_423 = _zz_1031;
  assign _zz_424 = _zz_1039;
  assign _zz_23 = ($signed(_zz_1047) * $signed(data_mid_9_real));
  assign _zz_425 = _zz_1048;
  assign _zz_21 = _zz_1051[31 : 0];
  assign _zz_426 = _zz_1052;
  assign _zz_22 = _zz_1055[31 : 0];
  assign _zz_24 = 1'b1;
  assign _zz_427 = _zz_1056;
  assign _zz_428 = _zz_1064;
  assign _zz_25 = 1'b1;
  assign _zz_429 = _zz_1072;
  assign _zz_430 = _zz_1080;
  assign _zz_28 = ($signed(_zz_1088) * $signed(data_mid_11_real));
  assign _zz_431 = _zz_1089;
  assign _zz_26 = _zz_1092[31 : 0];
  assign _zz_432 = _zz_1093;
  assign _zz_27 = _zz_1096[31 : 0];
  assign _zz_29 = 1'b1;
  assign _zz_433 = _zz_1097;
  assign _zz_434 = _zz_1105;
  assign _zz_30 = 1'b1;
  assign _zz_435 = _zz_1113;
  assign _zz_436 = _zz_1121;
  assign _zz_33 = ($signed(_zz_1129) * $signed(data_mid_13_real));
  assign _zz_437 = _zz_1130;
  assign _zz_31 = _zz_1133[31 : 0];
  assign _zz_438 = _zz_1134;
  assign _zz_32 = _zz_1137[31 : 0];
  assign _zz_34 = 1'b1;
  assign _zz_439 = _zz_1138;
  assign _zz_440 = _zz_1146;
  assign _zz_35 = 1'b1;
  assign _zz_441 = _zz_1154;
  assign _zz_442 = _zz_1162;
  assign _zz_38 = ($signed(_zz_1170) * $signed(data_mid_15_real));
  assign _zz_443 = _zz_1171;
  assign _zz_36 = _zz_1174[31 : 0];
  assign _zz_444 = _zz_1175;
  assign _zz_37 = _zz_1178[31 : 0];
  assign _zz_39 = 1'b1;
  assign _zz_445 = _zz_1179;
  assign _zz_446 = _zz_1187;
  assign _zz_40 = 1'b1;
  assign _zz_447 = _zz_1195;
  assign _zz_448 = _zz_1203;
  assign _zz_43 = ($signed(_zz_1211) * $signed(data_mid_17_real));
  assign _zz_449 = _zz_1212;
  assign _zz_41 = _zz_1215[31 : 0];
  assign _zz_450 = _zz_1216;
  assign _zz_42 = _zz_1219[31 : 0];
  assign _zz_44 = 1'b1;
  assign _zz_451 = _zz_1220;
  assign _zz_452 = _zz_1228;
  assign _zz_45 = 1'b1;
  assign _zz_453 = _zz_1236;
  assign _zz_454 = _zz_1244;
  assign _zz_48 = ($signed(_zz_1252) * $signed(data_mid_19_real));
  assign _zz_455 = _zz_1253;
  assign _zz_46 = _zz_1256[31 : 0];
  assign _zz_456 = _zz_1257;
  assign _zz_47 = _zz_1260[31 : 0];
  assign _zz_49 = 1'b1;
  assign _zz_457 = _zz_1261;
  assign _zz_458 = _zz_1269;
  assign _zz_50 = 1'b1;
  assign _zz_459 = _zz_1277;
  assign _zz_460 = _zz_1285;
  assign _zz_53 = ($signed(_zz_1293) * $signed(data_mid_21_real));
  assign _zz_461 = _zz_1294;
  assign _zz_51 = _zz_1297[31 : 0];
  assign _zz_462 = _zz_1298;
  assign _zz_52 = _zz_1301[31 : 0];
  assign _zz_54 = 1'b1;
  assign _zz_463 = _zz_1302;
  assign _zz_464 = _zz_1310;
  assign _zz_55 = 1'b1;
  assign _zz_465 = _zz_1318;
  assign _zz_466 = _zz_1326;
  assign _zz_58 = ($signed(_zz_1334) * $signed(data_mid_23_real));
  assign _zz_467 = _zz_1335;
  assign _zz_56 = _zz_1338[31 : 0];
  assign _zz_468 = _zz_1339;
  assign _zz_57 = _zz_1342[31 : 0];
  assign _zz_59 = 1'b1;
  assign _zz_469 = _zz_1343;
  assign _zz_470 = _zz_1351;
  assign _zz_60 = 1'b1;
  assign _zz_471 = _zz_1359;
  assign _zz_472 = _zz_1367;
  assign _zz_63 = ($signed(_zz_1375) * $signed(data_mid_25_real));
  assign _zz_473 = _zz_1376;
  assign _zz_61 = _zz_1379[31 : 0];
  assign _zz_474 = _zz_1380;
  assign _zz_62 = _zz_1383[31 : 0];
  assign _zz_64 = 1'b1;
  assign _zz_475 = _zz_1384;
  assign _zz_476 = _zz_1392;
  assign _zz_65 = 1'b1;
  assign _zz_477 = _zz_1400;
  assign _zz_478 = _zz_1408;
  assign _zz_68 = ($signed(_zz_1416) * $signed(data_mid_27_real));
  assign _zz_479 = _zz_1417;
  assign _zz_66 = _zz_1420[31 : 0];
  assign _zz_480 = _zz_1421;
  assign _zz_67 = _zz_1424[31 : 0];
  assign _zz_69 = 1'b1;
  assign _zz_481 = _zz_1425;
  assign _zz_482 = _zz_1433;
  assign _zz_70 = 1'b1;
  assign _zz_483 = _zz_1441;
  assign _zz_484 = _zz_1449;
  assign _zz_73 = ($signed(_zz_1457) * $signed(data_mid_29_real));
  assign _zz_485 = _zz_1458;
  assign _zz_71 = _zz_1461[31 : 0];
  assign _zz_486 = _zz_1462;
  assign _zz_72 = _zz_1465[31 : 0];
  assign _zz_74 = 1'b1;
  assign _zz_487 = _zz_1466;
  assign _zz_488 = _zz_1474;
  assign _zz_75 = 1'b1;
  assign _zz_489 = _zz_1482;
  assign _zz_490 = _zz_1490;
  assign _zz_78 = ($signed(_zz_1498) * $signed(data_mid_31_real));
  assign _zz_491 = _zz_1499;
  assign _zz_76 = _zz_1502[31 : 0];
  assign _zz_492 = _zz_1503;
  assign _zz_77 = _zz_1506[31 : 0];
  assign _zz_79 = 1'b1;
  assign _zz_493 = _zz_1507;
  assign _zz_494 = _zz_1515;
  assign _zz_80 = 1'b1;
  assign _zz_495 = _zz_1523;
  assign _zz_496 = _zz_1531;
  assign _zz_83 = ($signed(_zz_1539) * $signed(data_mid_2_real));
  assign _zz_497 = _zz_1540;
  assign _zz_81 = _zz_1543[31 : 0];
  assign _zz_498 = _zz_1544;
  assign _zz_82 = _zz_1547[31 : 0];
  assign _zz_84 = 1'b1;
  assign _zz_499 = _zz_1548;
  assign _zz_500 = _zz_1556;
  assign _zz_85 = 1'b1;
  assign _zz_501 = _zz_1564;
  assign _zz_502 = _zz_1572;
  assign _zz_88 = ($signed(_zz_1580) * $signed(data_mid_3_real));
  assign _zz_503 = _zz_1581;
  assign _zz_86 = _zz_1584[31 : 0];
  assign _zz_504 = _zz_1585;
  assign _zz_87 = _zz_1588[31 : 0];
  assign _zz_89 = 1'b1;
  assign _zz_505 = _zz_1589;
  assign _zz_506 = _zz_1597;
  assign _zz_90 = 1'b1;
  assign _zz_507 = _zz_1605;
  assign _zz_508 = _zz_1613;
  assign _zz_93 = ($signed(_zz_1621) * $signed(data_mid_6_real));
  assign _zz_509 = _zz_1622;
  assign _zz_91 = _zz_1625[31 : 0];
  assign _zz_510 = _zz_1626;
  assign _zz_92 = _zz_1629[31 : 0];
  assign _zz_94 = 1'b1;
  assign _zz_511 = _zz_1630;
  assign _zz_512 = _zz_1638;
  assign _zz_95 = 1'b1;
  assign _zz_513 = _zz_1646;
  assign _zz_514 = _zz_1654;
  assign _zz_98 = ($signed(_zz_1662) * $signed(data_mid_7_real));
  assign _zz_515 = _zz_1663;
  assign _zz_96 = _zz_1666[31 : 0];
  assign _zz_516 = _zz_1667;
  assign _zz_97 = _zz_1670[31 : 0];
  assign _zz_99 = 1'b1;
  assign _zz_517 = _zz_1671;
  assign _zz_518 = _zz_1679;
  assign _zz_100 = 1'b1;
  assign _zz_519 = _zz_1687;
  assign _zz_520 = _zz_1695;
  assign _zz_103 = ($signed(_zz_1703) * $signed(data_mid_10_real));
  assign _zz_521 = _zz_1704;
  assign _zz_101 = _zz_1707[31 : 0];
  assign _zz_522 = _zz_1708;
  assign _zz_102 = _zz_1711[31 : 0];
  assign _zz_104 = 1'b1;
  assign _zz_523 = _zz_1712;
  assign _zz_524 = _zz_1720;
  assign _zz_105 = 1'b1;
  assign _zz_525 = _zz_1728;
  assign _zz_526 = _zz_1736;
  assign _zz_108 = ($signed(_zz_1744) * $signed(data_mid_11_real));
  assign _zz_527 = _zz_1745;
  assign _zz_106 = _zz_1748[31 : 0];
  assign _zz_528 = _zz_1749;
  assign _zz_107 = _zz_1752[31 : 0];
  assign _zz_109 = 1'b1;
  assign _zz_529 = _zz_1753;
  assign _zz_530 = _zz_1761;
  assign _zz_110 = 1'b1;
  assign _zz_531 = _zz_1769;
  assign _zz_532 = _zz_1777;
  assign _zz_113 = ($signed(_zz_1785) * $signed(data_mid_14_real));
  assign _zz_533 = _zz_1786;
  assign _zz_111 = _zz_1789[31 : 0];
  assign _zz_534 = _zz_1790;
  assign _zz_112 = _zz_1793[31 : 0];
  assign _zz_114 = 1'b1;
  assign _zz_535 = _zz_1794;
  assign _zz_536 = _zz_1802;
  assign _zz_115 = 1'b1;
  assign _zz_537 = _zz_1810;
  assign _zz_538 = _zz_1818;
  assign _zz_118 = ($signed(_zz_1826) * $signed(data_mid_15_real));
  assign _zz_539 = _zz_1827;
  assign _zz_116 = _zz_1830[31 : 0];
  assign _zz_540 = _zz_1831;
  assign _zz_117 = _zz_1834[31 : 0];
  assign _zz_119 = 1'b1;
  assign _zz_541 = _zz_1835;
  assign _zz_542 = _zz_1843;
  assign _zz_120 = 1'b1;
  assign _zz_543 = _zz_1851;
  assign _zz_544 = _zz_1859;
  assign _zz_123 = ($signed(_zz_1867) * $signed(data_mid_18_real));
  assign _zz_545 = _zz_1868;
  assign _zz_121 = _zz_1871[31 : 0];
  assign _zz_546 = _zz_1872;
  assign _zz_122 = _zz_1875[31 : 0];
  assign _zz_124 = 1'b1;
  assign _zz_547 = _zz_1876;
  assign _zz_548 = _zz_1884;
  assign _zz_125 = 1'b1;
  assign _zz_549 = _zz_1892;
  assign _zz_550 = _zz_1900;
  assign _zz_128 = ($signed(_zz_1908) * $signed(data_mid_19_real));
  assign _zz_551 = _zz_1909;
  assign _zz_126 = _zz_1912[31 : 0];
  assign _zz_552 = _zz_1913;
  assign _zz_127 = _zz_1916[31 : 0];
  assign _zz_129 = 1'b1;
  assign _zz_553 = _zz_1917;
  assign _zz_554 = _zz_1925;
  assign _zz_130 = 1'b1;
  assign _zz_555 = _zz_1933;
  assign _zz_556 = _zz_1941;
  assign _zz_133 = ($signed(_zz_1949) * $signed(data_mid_22_real));
  assign _zz_557 = _zz_1950;
  assign _zz_131 = _zz_1953[31 : 0];
  assign _zz_558 = _zz_1954;
  assign _zz_132 = _zz_1957[31 : 0];
  assign _zz_134 = 1'b1;
  assign _zz_559 = _zz_1958;
  assign _zz_560 = _zz_1966;
  assign _zz_135 = 1'b1;
  assign _zz_561 = _zz_1974;
  assign _zz_562 = _zz_1982;
  assign _zz_138 = ($signed(_zz_1990) * $signed(data_mid_23_real));
  assign _zz_563 = _zz_1991;
  assign _zz_136 = _zz_1994[31 : 0];
  assign _zz_564 = _zz_1995;
  assign _zz_137 = _zz_1998[31 : 0];
  assign _zz_139 = 1'b1;
  assign _zz_565 = _zz_1999;
  assign _zz_566 = _zz_2007;
  assign _zz_140 = 1'b1;
  assign _zz_567 = _zz_2015;
  assign _zz_568 = _zz_2023;
  assign _zz_143 = ($signed(_zz_2031) * $signed(data_mid_26_real));
  assign _zz_569 = _zz_2032;
  assign _zz_141 = _zz_2035[31 : 0];
  assign _zz_570 = _zz_2036;
  assign _zz_142 = _zz_2039[31 : 0];
  assign _zz_144 = 1'b1;
  assign _zz_571 = _zz_2040;
  assign _zz_572 = _zz_2048;
  assign _zz_145 = 1'b1;
  assign _zz_573 = _zz_2056;
  assign _zz_574 = _zz_2064;
  assign _zz_148 = ($signed(_zz_2072) * $signed(data_mid_27_real));
  assign _zz_575 = _zz_2073;
  assign _zz_146 = _zz_2076[31 : 0];
  assign _zz_576 = _zz_2077;
  assign _zz_147 = _zz_2080[31 : 0];
  assign _zz_149 = 1'b1;
  assign _zz_577 = _zz_2081;
  assign _zz_578 = _zz_2089;
  assign _zz_150 = 1'b1;
  assign _zz_579 = _zz_2097;
  assign _zz_580 = _zz_2105;
  assign _zz_153 = ($signed(_zz_2113) * $signed(data_mid_30_real));
  assign _zz_581 = _zz_2114;
  assign _zz_151 = _zz_2117[31 : 0];
  assign _zz_582 = _zz_2118;
  assign _zz_152 = _zz_2121[31 : 0];
  assign _zz_154 = 1'b1;
  assign _zz_583 = _zz_2122;
  assign _zz_584 = _zz_2130;
  assign _zz_155 = 1'b1;
  assign _zz_585 = _zz_2138;
  assign _zz_586 = _zz_2146;
  assign _zz_158 = ($signed(_zz_2154) * $signed(data_mid_31_real));
  assign _zz_587 = _zz_2155;
  assign _zz_156 = _zz_2158[31 : 0];
  assign _zz_588 = _zz_2159;
  assign _zz_157 = _zz_2162[31 : 0];
  assign _zz_159 = 1'b1;
  assign _zz_589 = _zz_2163;
  assign _zz_590 = _zz_2171;
  assign _zz_160 = 1'b1;
  assign _zz_591 = _zz_2179;
  assign _zz_592 = _zz_2187;
  assign _zz_163 = ($signed(_zz_2195) * $signed(data_mid_4_real));
  assign _zz_593 = _zz_2196;
  assign _zz_161 = _zz_2199[31 : 0];
  assign _zz_594 = _zz_2200;
  assign _zz_162 = _zz_2203[31 : 0];
  assign _zz_164 = 1'b1;
  assign _zz_595 = _zz_2204;
  assign _zz_596 = _zz_2212;
  assign _zz_165 = 1'b1;
  assign _zz_597 = _zz_2220;
  assign _zz_598 = _zz_2228;
  assign _zz_168 = ($signed(_zz_2236) * $signed(data_mid_5_real));
  assign _zz_599 = _zz_2237;
  assign _zz_166 = _zz_2240[31 : 0];
  assign _zz_600 = _zz_2241;
  assign _zz_167 = _zz_2244[31 : 0];
  assign _zz_169 = 1'b1;
  assign _zz_601 = _zz_2245;
  assign _zz_602 = _zz_2253;
  assign _zz_170 = 1'b1;
  assign _zz_603 = _zz_2261;
  assign _zz_604 = _zz_2269;
  assign _zz_173 = ($signed(_zz_2277) * $signed(data_mid_6_real));
  assign _zz_605 = _zz_2278;
  assign _zz_171 = _zz_2281[31 : 0];
  assign _zz_606 = _zz_2282;
  assign _zz_172 = _zz_2285[31 : 0];
  assign _zz_174 = 1'b1;
  assign _zz_607 = _zz_2286;
  assign _zz_608 = _zz_2294;
  assign _zz_175 = 1'b1;
  assign _zz_609 = _zz_2302;
  assign _zz_610 = _zz_2310;
  assign _zz_178 = ($signed(_zz_2318) * $signed(data_mid_7_real));
  assign _zz_611 = _zz_2319;
  assign _zz_176 = _zz_2322[31 : 0];
  assign _zz_612 = _zz_2323;
  assign _zz_177 = _zz_2326[31 : 0];
  assign _zz_179 = 1'b1;
  assign _zz_613 = _zz_2327;
  assign _zz_614 = _zz_2335;
  assign _zz_180 = 1'b1;
  assign _zz_615 = _zz_2343;
  assign _zz_616 = _zz_2351;
  assign _zz_183 = ($signed(_zz_2359) * $signed(data_mid_12_real));
  assign _zz_617 = _zz_2360;
  assign _zz_181 = _zz_2363[31 : 0];
  assign _zz_618 = _zz_2364;
  assign _zz_182 = _zz_2367[31 : 0];
  assign _zz_184 = 1'b1;
  assign _zz_619 = _zz_2368;
  assign _zz_620 = _zz_2376;
  assign _zz_185 = 1'b1;
  assign _zz_621 = _zz_2384;
  assign _zz_622 = _zz_2392;
  assign _zz_188 = ($signed(_zz_2400) * $signed(data_mid_13_real));
  assign _zz_623 = _zz_2401;
  assign _zz_186 = _zz_2404[31 : 0];
  assign _zz_624 = _zz_2405;
  assign _zz_187 = _zz_2408[31 : 0];
  assign _zz_189 = 1'b1;
  assign _zz_625 = _zz_2409;
  assign _zz_626 = _zz_2417;
  assign _zz_190 = 1'b1;
  assign _zz_627 = _zz_2425;
  assign _zz_628 = _zz_2433;
  assign _zz_193 = ($signed(_zz_2441) * $signed(data_mid_14_real));
  assign _zz_629 = _zz_2442;
  assign _zz_191 = _zz_2445[31 : 0];
  assign _zz_630 = _zz_2446;
  assign _zz_192 = _zz_2449[31 : 0];
  assign _zz_194 = 1'b1;
  assign _zz_631 = _zz_2450;
  assign _zz_632 = _zz_2458;
  assign _zz_195 = 1'b1;
  assign _zz_633 = _zz_2466;
  assign _zz_634 = _zz_2474;
  assign _zz_198 = ($signed(_zz_2482) * $signed(data_mid_15_real));
  assign _zz_635 = _zz_2483;
  assign _zz_196 = _zz_2486[31 : 0];
  assign _zz_636 = _zz_2487;
  assign _zz_197 = _zz_2490[31 : 0];
  assign _zz_199 = 1'b1;
  assign _zz_637 = _zz_2491;
  assign _zz_638 = _zz_2499;
  assign _zz_200 = 1'b1;
  assign _zz_639 = _zz_2507;
  assign _zz_640 = _zz_2515;
  assign _zz_203 = ($signed(_zz_2523) * $signed(data_mid_20_real));
  assign _zz_641 = _zz_2524;
  assign _zz_201 = _zz_2527[31 : 0];
  assign _zz_642 = _zz_2528;
  assign _zz_202 = _zz_2531[31 : 0];
  assign _zz_204 = 1'b1;
  assign _zz_643 = _zz_2532;
  assign _zz_644 = _zz_2540;
  assign _zz_205 = 1'b1;
  assign _zz_645 = _zz_2548;
  assign _zz_646 = _zz_2556;
  assign _zz_208 = ($signed(_zz_2564) * $signed(data_mid_21_real));
  assign _zz_647 = _zz_2565;
  assign _zz_206 = _zz_2568[31 : 0];
  assign _zz_648 = _zz_2569;
  assign _zz_207 = _zz_2572[31 : 0];
  assign _zz_209 = 1'b1;
  assign _zz_649 = _zz_2573;
  assign _zz_650 = _zz_2581;
  assign _zz_210 = 1'b1;
  assign _zz_651 = _zz_2589;
  assign _zz_652 = _zz_2597;
  assign _zz_213 = ($signed(_zz_2605) * $signed(data_mid_22_real));
  assign _zz_653 = _zz_2606;
  assign _zz_211 = _zz_2609[31 : 0];
  assign _zz_654 = _zz_2610;
  assign _zz_212 = _zz_2613[31 : 0];
  assign _zz_214 = 1'b1;
  assign _zz_655 = _zz_2614;
  assign _zz_656 = _zz_2622;
  assign _zz_215 = 1'b1;
  assign _zz_657 = _zz_2630;
  assign _zz_658 = _zz_2638;
  assign _zz_218 = ($signed(_zz_2646) * $signed(data_mid_23_real));
  assign _zz_659 = _zz_2647;
  assign _zz_216 = _zz_2650[31 : 0];
  assign _zz_660 = _zz_2651;
  assign _zz_217 = _zz_2654[31 : 0];
  assign _zz_219 = 1'b1;
  assign _zz_661 = _zz_2655;
  assign _zz_662 = _zz_2663;
  assign _zz_220 = 1'b1;
  assign _zz_663 = _zz_2671;
  assign _zz_664 = _zz_2679;
  assign _zz_223 = ($signed(_zz_2687) * $signed(data_mid_28_real));
  assign _zz_665 = _zz_2688;
  assign _zz_221 = _zz_2691[31 : 0];
  assign _zz_666 = _zz_2692;
  assign _zz_222 = _zz_2695[31 : 0];
  assign _zz_224 = 1'b1;
  assign _zz_667 = _zz_2696;
  assign _zz_668 = _zz_2704;
  assign _zz_225 = 1'b1;
  assign _zz_669 = _zz_2712;
  assign _zz_670 = _zz_2720;
  assign _zz_228 = ($signed(_zz_2728) * $signed(data_mid_29_real));
  assign _zz_671 = _zz_2729;
  assign _zz_226 = _zz_2732[31 : 0];
  assign _zz_672 = _zz_2733;
  assign _zz_227 = _zz_2736[31 : 0];
  assign _zz_229 = 1'b1;
  assign _zz_673 = _zz_2737;
  assign _zz_674 = _zz_2745;
  assign _zz_230 = 1'b1;
  assign _zz_675 = _zz_2753;
  assign _zz_676 = _zz_2761;
  assign _zz_233 = ($signed(_zz_2769) * $signed(data_mid_30_real));
  assign _zz_677 = _zz_2770;
  assign _zz_231 = _zz_2773[31 : 0];
  assign _zz_678 = _zz_2774;
  assign _zz_232 = _zz_2777[31 : 0];
  assign _zz_234 = 1'b1;
  assign _zz_679 = _zz_2778;
  assign _zz_680 = _zz_2786;
  assign _zz_235 = 1'b1;
  assign _zz_681 = _zz_2794;
  assign _zz_682 = _zz_2802;
  assign _zz_238 = ($signed(_zz_2810) * $signed(data_mid_31_real));
  assign _zz_683 = _zz_2811;
  assign _zz_236 = _zz_2814[31 : 0];
  assign _zz_684 = _zz_2815;
  assign _zz_237 = _zz_2818[31 : 0];
  assign _zz_239 = 1'b1;
  assign _zz_685 = _zz_2819;
  assign _zz_686 = _zz_2827;
  assign _zz_240 = 1'b1;
  assign _zz_687 = _zz_2835;
  assign _zz_688 = _zz_2843;
  assign _zz_243 = ($signed(_zz_2851) * $signed(data_mid_8_real));
  assign _zz_689 = _zz_2852;
  assign _zz_241 = _zz_2855[31 : 0];
  assign _zz_690 = _zz_2856;
  assign _zz_242 = _zz_2859[31 : 0];
  assign _zz_244 = 1'b1;
  assign _zz_691 = _zz_2860;
  assign _zz_692 = _zz_2868;
  assign _zz_245 = 1'b1;
  assign _zz_693 = _zz_2876;
  assign _zz_694 = _zz_2884;
  assign _zz_248 = ($signed(_zz_2892) * $signed(data_mid_9_real));
  assign _zz_695 = _zz_2893;
  assign _zz_246 = _zz_2896[31 : 0];
  assign _zz_696 = _zz_2897;
  assign _zz_247 = _zz_2900[31 : 0];
  assign _zz_249 = 1'b1;
  assign _zz_697 = _zz_2901;
  assign _zz_698 = _zz_2909;
  assign _zz_250 = 1'b1;
  assign _zz_699 = _zz_2917;
  assign _zz_700 = _zz_2925;
  assign _zz_253 = ($signed(_zz_2933) * $signed(data_mid_10_real));
  assign _zz_701 = _zz_2934;
  assign _zz_251 = _zz_2937[31 : 0];
  assign _zz_702 = _zz_2938;
  assign _zz_252 = _zz_2941[31 : 0];
  assign _zz_254 = 1'b1;
  assign _zz_703 = _zz_2942;
  assign _zz_704 = _zz_2950;
  assign _zz_255 = 1'b1;
  assign _zz_705 = _zz_2958;
  assign _zz_706 = _zz_2966;
  assign _zz_258 = ($signed(_zz_2974) * $signed(data_mid_11_real));
  assign _zz_707 = _zz_2975;
  assign _zz_256 = _zz_2978[31 : 0];
  assign _zz_708 = _zz_2979;
  assign _zz_257 = _zz_2982[31 : 0];
  assign _zz_259 = 1'b1;
  assign _zz_709 = _zz_2983;
  assign _zz_710 = _zz_2991;
  assign _zz_260 = 1'b1;
  assign _zz_711 = _zz_2999;
  assign _zz_712 = _zz_3007;
  assign _zz_263 = ($signed(_zz_3015) * $signed(data_mid_12_real));
  assign _zz_713 = _zz_3016;
  assign _zz_261 = _zz_3019[31 : 0];
  assign _zz_714 = _zz_3020;
  assign _zz_262 = _zz_3023[31 : 0];
  assign _zz_264 = 1'b1;
  assign _zz_715 = _zz_3024;
  assign _zz_716 = _zz_3032;
  assign _zz_265 = 1'b1;
  assign _zz_717 = _zz_3040;
  assign _zz_718 = _zz_3048;
  assign _zz_268 = ($signed(_zz_3056) * $signed(data_mid_13_real));
  assign _zz_719 = _zz_3057;
  assign _zz_266 = _zz_3060[31 : 0];
  assign _zz_720 = _zz_3061;
  assign _zz_267 = _zz_3064[31 : 0];
  assign _zz_269 = 1'b1;
  assign _zz_721 = _zz_3065;
  assign _zz_722 = _zz_3073;
  assign _zz_270 = 1'b1;
  assign _zz_723 = _zz_3081;
  assign _zz_724 = _zz_3089;
  assign _zz_273 = ($signed(_zz_3097) * $signed(data_mid_14_real));
  assign _zz_725 = _zz_3098;
  assign _zz_271 = _zz_3101[31 : 0];
  assign _zz_726 = _zz_3102;
  assign _zz_272 = _zz_3105[31 : 0];
  assign _zz_274 = 1'b1;
  assign _zz_727 = _zz_3106;
  assign _zz_728 = _zz_3114;
  assign _zz_275 = 1'b1;
  assign _zz_729 = _zz_3122;
  assign _zz_730 = _zz_3130;
  assign _zz_278 = ($signed(_zz_3138) * $signed(data_mid_15_real));
  assign _zz_731 = _zz_3139;
  assign _zz_276 = _zz_3142[31 : 0];
  assign _zz_732 = _zz_3143;
  assign _zz_277 = _zz_3146[31 : 0];
  assign _zz_279 = 1'b1;
  assign _zz_733 = _zz_3147;
  assign _zz_734 = _zz_3155;
  assign _zz_280 = 1'b1;
  assign _zz_735 = _zz_3163;
  assign _zz_736 = _zz_3171;
  assign _zz_283 = ($signed(_zz_3179) * $signed(data_mid_24_real));
  assign _zz_737 = _zz_3180;
  assign _zz_281 = _zz_3183[31 : 0];
  assign _zz_738 = _zz_3184;
  assign _zz_282 = _zz_3187[31 : 0];
  assign _zz_284 = 1'b1;
  assign _zz_739 = _zz_3188;
  assign _zz_740 = _zz_3196;
  assign _zz_285 = 1'b1;
  assign _zz_741 = _zz_3204;
  assign _zz_742 = _zz_3212;
  assign _zz_288 = ($signed(_zz_3220) * $signed(data_mid_25_real));
  assign _zz_743 = _zz_3221;
  assign _zz_286 = _zz_3224[31 : 0];
  assign _zz_744 = _zz_3225;
  assign _zz_287 = _zz_3228[31 : 0];
  assign _zz_289 = 1'b1;
  assign _zz_745 = _zz_3229;
  assign _zz_746 = _zz_3237;
  assign _zz_290 = 1'b1;
  assign _zz_747 = _zz_3245;
  assign _zz_748 = _zz_3253;
  assign _zz_293 = ($signed(_zz_3261) * $signed(data_mid_26_real));
  assign _zz_749 = _zz_3262;
  assign _zz_291 = _zz_3265[31 : 0];
  assign _zz_750 = _zz_3266;
  assign _zz_292 = _zz_3269[31 : 0];
  assign _zz_294 = 1'b1;
  assign _zz_751 = _zz_3270;
  assign _zz_752 = _zz_3278;
  assign _zz_295 = 1'b1;
  assign _zz_753 = _zz_3286;
  assign _zz_754 = _zz_3294;
  assign _zz_298 = ($signed(_zz_3302) * $signed(data_mid_27_real));
  assign _zz_755 = _zz_3303;
  assign _zz_296 = _zz_3306[31 : 0];
  assign _zz_756 = _zz_3307;
  assign _zz_297 = _zz_3310[31 : 0];
  assign _zz_299 = 1'b1;
  assign _zz_757 = _zz_3311;
  assign _zz_758 = _zz_3319;
  assign _zz_300 = 1'b1;
  assign _zz_759 = _zz_3327;
  assign _zz_760 = _zz_3335;
  assign _zz_303 = ($signed(_zz_3343) * $signed(data_mid_28_real));
  assign _zz_761 = _zz_3344;
  assign _zz_301 = _zz_3347[31 : 0];
  assign _zz_762 = _zz_3348;
  assign _zz_302 = _zz_3351[31 : 0];
  assign _zz_304 = 1'b1;
  assign _zz_763 = _zz_3352;
  assign _zz_764 = _zz_3360;
  assign _zz_305 = 1'b1;
  assign _zz_765 = _zz_3368;
  assign _zz_766 = _zz_3376;
  assign _zz_308 = ($signed(_zz_3384) * $signed(data_mid_29_real));
  assign _zz_767 = _zz_3385;
  assign _zz_306 = _zz_3388[31 : 0];
  assign _zz_768 = _zz_3389;
  assign _zz_307 = _zz_3392[31 : 0];
  assign _zz_309 = 1'b1;
  assign _zz_769 = _zz_3393;
  assign _zz_770 = _zz_3401;
  assign _zz_310 = 1'b1;
  assign _zz_771 = _zz_3409;
  assign _zz_772 = _zz_3417;
  assign _zz_313 = ($signed(_zz_3425) * $signed(data_mid_30_real));
  assign _zz_773 = _zz_3426;
  assign _zz_311 = _zz_3429[31 : 0];
  assign _zz_774 = _zz_3430;
  assign _zz_312 = _zz_3433[31 : 0];
  assign _zz_314 = 1'b1;
  assign _zz_775 = _zz_3434;
  assign _zz_776 = _zz_3442;
  assign _zz_315 = 1'b1;
  assign _zz_777 = _zz_3450;
  assign _zz_778 = _zz_3458;
  assign _zz_318 = ($signed(_zz_3466) * $signed(data_mid_31_real));
  assign _zz_779 = _zz_3467;
  assign _zz_316 = _zz_3470[31 : 0];
  assign _zz_780 = _zz_3471;
  assign _zz_317 = _zz_3474[31 : 0];
  assign _zz_319 = 1'b1;
  assign _zz_781 = _zz_3475;
  assign _zz_782 = _zz_3483;
  assign _zz_320 = 1'b1;
  assign _zz_783 = _zz_3491;
  assign _zz_784 = _zz_3499;
  assign _zz_323 = ($signed(_zz_3507) * $signed(data_mid_16_real));
  assign _zz_785 = _zz_3508;
  assign _zz_321 = _zz_3511[31 : 0];
  assign _zz_786 = _zz_3512;
  assign _zz_322 = _zz_3515[31 : 0];
  assign _zz_324 = 1'b1;
  assign _zz_787 = _zz_3516;
  assign _zz_788 = _zz_3524;
  assign _zz_325 = 1'b1;
  assign _zz_789 = _zz_3532;
  assign _zz_790 = _zz_3540;
  assign _zz_328 = ($signed(_zz_3548) * $signed(data_mid_17_real));
  assign _zz_791 = _zz_3549;
  assign _zz_326 = _zz_3552[31 : 0];
  assign _zz_792 = _zz_3553;
  assign _zz_327 = _zz_3556[31 : 0];
  assign _zz_329 = 1'b1;
  assign _zz_793 = _zz_3557;
  assign _zz_794 = _zz_3565;
  assign _zz_330 = 1'b1;
  assign _zz_795 = _zz_3573;
  assign _zz_796 = _zz_3581;
  assign _zz_333 = ($signed(_zz_3589) * $signed(data_mid_18_real));
  assign _zz_797 = _zz_3590;
  assign _zz_331 = _zz_3593[31 : 0];
  assign _zz_798 = _zz_3594;
  assign _zz_332 = _zz_3597[31 : 0];
  assign _zz_334 = 1'b1;
  assign _zz_799 = _zz_3598;
  assign _zz_800 = _zz_3606;
  assign _zz_335 = 1'b1;
  assign _zz_801 = _zz_3614;
  assign _zz_802 = _zz_3622;
  assign _zz_338 = ($signed(_zz_3630) * $signed(data_mid_19_real));
  assign _zz_803 = _zz_3631;
  assign _zz_336 = _zz_3634[31 : 0];
  assign _zz_804 = _zz_3635;
  assign _zz_337 = _zz_3638[31 : 0];
  assign _zz_339 = 1'b1;
  assign _zz_805 = _zz_3639;
  assign _zz_806 = _zz_3647;
  assign _zz_340 = 1'b1;
  assign _zz_807 = _zz_3655;
  assign _zz_808 = _zz_3663;
  assign _zz_343 = ($signed(_zz_3671) * $signed(data_mid_20_real));
  assign _zz_809 = _zz_3672;
  assign _zz_341 = _zz_3675[31 : 0];
  assign _zz_810 = _zz_3676;
  assign _zz_342 = _zz_3679[31 : 0];
  assign _zz_344 = 1'b1;
  assign _zz_811 = _zz_3680;
  assign _zz_812 = _zz_3688;
  assign _zz_345 = 1'b1;
  assign _zz_813 = _zz_3696;
  assign _zz_814 = _zz_3704;
  assign _zz_348 = ($signed(_zz_3712) * $signed(data_mid_21_real));
  assign _zz_815 = _zz_3713;
  assign _zz_346 = _zz_3716[31 : 0];
  assign _zz_816 = _zz_3717;
  assign _zz_347 = _zz_3720[31 : 0];
  assign _zz_349 = 1'b1;
  assign _zz_817 = _zz_3721;
  assign _zz_818 = _zz_3729;
  assign _zz_350 = 1'b1;
  assign _zz_819 = _zz_3737;
  assign _zz_820 = _zz_3745;
  assign _zz_353 = ($signed(_zz_3753) * $signed(data_mid_22_real));
  assign _zz_821 = _zz_3754;
  assign _zz_351 = _zz_3757[31 : 0];
  assign _zz_822 = _zz_3758;
  assign _zz_352 = _zz_3761[31 : 0];
  assign _zz_354 = 1'b1;
  assign _zz_823 = _zz_3762;
  assign _zz_824 = _zz_3770;
  assign _zz_355 = 1'b1;
  assign _zz_825 = _zz_3778;
  assign _zz_826 = _zz_3786;
  assign _zz_358 = ($signed(_zz_3794) * $signed(data_mid_23_real));
  assign _zz_827 = _zz_3795;
  assign _zz_356 = _zz_3798[31 : 0];
  assign _zz_828 = _zz_3799;
  assign _zz_357 = _zz_3802[31 : 0];
  assign _zz_359 = 1'b1;
  assign _zz_829 = _zz_3803;
  assign _zz_830 = _zz_3811;
  assign _zz_360 = 1'b1;
  assign _zz_831 = _zz_3819;
  assign _zz_832 = _zz_3827;
  assign _zz_363 = ($signed(_zz_3835) * $signed(data_mid_24_real));
  assign _zz_833 = _zz_3836;
  assign _zz_361 = _zz_3839[31 : 0];
  assign _zz_834 = _zz_3840;
  assign _zz_362 = _zz_3843[31 : 0];
  assign _zz_364 = 1'b1;
  assign _zz_835 = _zz_3844;
  assign _zz_836 = _zz_3852;
  assign _zz_365 = 1'b1;
  assign _zz_837 = _zz_3860;
  assign _zz_838 = _zz_3868;
  assign _zz_368 = ($signed(_zz_3876) * $signed(data_mid_25_real));
  assign _zz_839 = _zz_3877;
  assign _zz_366 = _zz_3880[31 : 0];
  assign _zz_840 = _zz_3881;
  assign _zz_367 = _zz_3884[31 : 0];
  assign _zz_369 = 1'b1;
  assign _zz_841 = _zz_3885;
  assign _zz_842 = _zz_3893;
  assign _zz_370 = 1'b1;
  assign _zz_843 = _zz_3901;
  assign _zz_844 = _zz_3909;
  assign _zz_373 = ($signed(_zz_3917) * $signed(data_mid_26_real));
  assign _zz_845 = _zz_3918;
  assign _zz_371 = _zz_3921[31 : 0];
  assign _zz_846 = _zz_3922;
  assign _zz_372 = _zz_3925[31 : 0];
  assign _zz_374 = 1'b1;
  assign _zz_847 = _zz_3926;
  assign _zz_848 = _zz_3934;
  assign _zz_375 = 1'b1;
  assign _zz_849 = _zz_3942;
  assign _zz_850 = _zz_3950;
  assign _zz_378 = ($signed(_zz_3958) * $signed(data_mid_27_real));
  assign _zz_851 = _zz_3959;
  assign _zz_376 = _zz_3962[31 : 0];
  assign _zz_852 = _zz_3963;
  assign _zz_377 = _zz_3966[31 : 0];
  assign _zz_379 = 1'b1;
  assign _zz_853 = _zz_3967;
  assign _zz_854 = _zz_3975;
  assign _zz_380 = 1'b1;
  assign _zz_855 = _zz_3983;
  assign _zz_856 = _zz_3991;
  assign _zz_383 = ($signed(_zz_3999) * $signed(data_mid_28_real));
  assign _zz_857 = _zz_4000;
  assign _zz_381 = _zz_4003[31 : 0];
  assign _zz_858 = _zz_4004;
  assign _zz_382 = _zz_4007[31 : 0];
  assign _zz_384 = 1'b1;
  assign _zz_859 = _zz_4008;
  assign _zz_860 = _zz_4016;
  assign _zz_385 = 1'b1;
  assign _zz_861 = _zz_4024;
  assign _zz_862 = _zz_4032;
  assign _zz_388 = ($signed(_zz_4040) * $signed(data_mid_29_real));
  assign _zz_863 = _zz_4041;
  assign _zz_386 = _zz_4044[31 : 0];
  assign _zz_864 = _zz_4045;
  assign _zz_387 = _zz_4048[31 : 0];
  assign _zz_389 = 1'b1;
  assign _zz_865 = _zz_4049;
  assign _zz_866 = _zz_4057;
  assign _zz_390 = 1'b1;
  assign _zz_867 = _zz_4065;
  assign _zz_868 = _zz_4073;
  assign _zz_393 = ($signed(_zz_4081) * $signed(data_mid_30_real));
  assign _zz_869 = _zz_4082;
  assign _zz_391 = _zz_4085[31 : 0];
  assign _zz_870 = _zz_4086;
  assign _zz_392 = _zz_4089[31 : 0];
  assign _zz_394 = 1'b1;
  assign _zz_871 = _zz_4090;
  assign _zz_872 = _zz_4098;
  assign _zz_395 = 1'b1;
  assign _zz_873 = _zz_4106;
  assign _zz_874 = _zz_4114;
  assign _zz_398 = ($signed(_zz_4122) * $signed(data_mid_31_real));
  assign _zz_875 = _zz_4123;
  assign _zz_396 = _zz_4126[31 : 0];
  assign _zz_876 = _zz_4127;
  assign _zz_397 = _zz_4130[31 : 0];
  assign _zz_399 = 1'b1;
  assign _zz_877 = _zz_4131;
  assign _zz_878 = _zz_4139;
  assign _zz_400 = 1'b1;
  assign _zz_879 = _zz_4147;
  assign _zz_880 = _zz_4155;
  assign sdata_out_valid = current_level_willOverflow_regNext;
  assign sdata_out_payload_0_real = data_mid_0_real;
  assign sdata_out_payload_0_imag = data_mid_0_imag;
  assign sdata_out_payload_1_real = data_mid_1_real;
  assign sdata_out_payload_1_imag = data_mid_1_imag;
  assign sdata_out_payload_2_real = data_mid_2_real;
  assign sdata_out_payload_2_imag = data_mid_2_imag;
  assign sdata_out_payload_3_real = data_mid_3_real;
  assign sdata_out_payload_3_imag = data_mid_3_imag;
  assign sdata_out_payload_4_real = data_mid_4_real;
  assign sdata_out_payload_4_imag = data_mid_4_imag;
  assign sdata_out_payload_5_real = data_mid_5_real;
  assign sdata_out_payload_5_imag = data_mid_5_imag;
  assign sdata_out_payload_6_real = data_mid_6_real;
  assign sdata_out_payload_6_imag = data_mid_6_imag;
  assign sdata_out_payload_7_real = data_mid_7_real;
  assign sdata_out_payload_7_imag = data_mid_7_imag;
  assign sdata_out_payload_8_real = data_mid_8_real;
  assign sdata_out_payload_8_imag = data_mid_8_imag;
  assign sdata_out_payload_9_real = data_mid_9_real;
  assign sdata_out_payload_9_imag = data_mid_9_imag;
  assign sdata_out_payload_10_real = data_mid_10_real;
  assign sdata_out_payload_10_imag = data_mid_10_imag;
  assign sdata_out_payload_11_real = data_mid_11_real;
  assign sdata_out_payload_11_imag = data_mid_11_imag;
  assign sdata_out_payload_12_real = data_mid_12_real;
  assign sdata_out_payload_12_imag = data_mid_12_imag;
  assign sdata_out_payload_13_real = data_mid_13_real;
  assign sdata_out_payload_13_imag = data_mid_13_imag;
  assign sdata_out_payload_14_real = data_mid_14_real;
  assign sdata_out_payload_14_imag = data_mid_14_imag;
  assign sdata_out_payload_15_real = data_mid_15_real;
  assign sdata_out_payload_15_imag = data_mid_15_imag;
  assign sdata_out_payload_16_real = data_mid_16_real;
  assign sdata_out_payload_16_imag = data_mid_16_imag;
  assign sdata_out_payload_17_real = data_mid_17_real;
  assign sdata_out_payload_17_imag = data_mid_17_imag;
  assign sdata_out_payload_18_real = data_mid_18_real;
  assign sdata_out_payload_18_imag = data_mid_18_imag;
  assign sdata_out_payload_19_real = data_mid_19_real;
  assign sdata_out_payload_19_imag = data_mid_19_imag;
  assign sdata_out_payload_20_real = data_mid_20_real;
  assign sdata_out_payload_20_imag = data_mid_20_imag;
  assign sdata_out_payload_21_real = data_mid_21_real;
  assign sdata_out_payload_21_imag = data_mid_21_imag;
  assign sdata_out_payload_22_real = data_mid_22_real;
  assign sdata_out_payload_22_imag = data_mid_22_imag;
  assign sdata_out_payload_23_real = data_mid_23_real;
  assign sdata_out_payload_23_imag = data_mid_23_imag;
  assign sdata_out_payload_24_real = data_mid_24_real;
  assign sdata_out_payload_24_imag = data_mid_24_imag;
  assign sdata_out_payload_25_real = data_mid_25_real;
  assign sdata_out_payload_25_imag = data_mid_25_imag;
  assign sdata_out_payload_26_real = data_mid_26_real;
  assign sdata_out_payload_26_imag = data_mid_26_imag;
  assign sdata_out_payload_27_real = data_mid_27_real;
  assign sdata_out_payload_27_imag = data_mid_27_imag;
  assign sdata_out_payload_28_real = data_mid_28_real;
  assign sdata_out_payload_28_imag = data_mid_28_imag;
  assign sdata_out_payload_29_real = data_mid_29_real;
  assign sdata_out_payload_29_imag = data_mid_29_imag;
  assign sdata_out_payload_30_real = data_mid_30_real;
  assign sdata_out_payload_30_imag = data_mid_30_imag;
  assign sdata_out_payload_31_real = data_mid_31_real;
  assign sdata_out_payload_31_imag = data_mid_31_imag;
  always @ (posedge clk) begin
    if(io_data_in_valid)begin
      data_in_0_real <= io_data_in_payload_0_real;
      data_in_0_imag <= io_data_in_payload_0_imag;
      data_in_1_real <= io_data_in_payload_1_real;
      data_in_1_imag <= io_data_in_payload_1_imag;
      data_in_2_real <= io_data_in_payload_2_real;
      data_in_2_imag <= io_data_in_payload_2_imag;
      data_in_3_real <= io_data_in_payload_3_real;
      data_in_3_imag <= io_data_in_payload_3_imag;
      data_in_4_real <= io_data_in_payload_4_real;
      data_in_4_imag <= io_data_in_payload_4_imag;
      data_in_5_real <= io_data_in_payload_5_real;
      data_in_5_imag <= io_data_in_payload_5_imag;
      data_in_6_real <= io_data_in_payload_6_real;
      data_in_6_imag <= io_data_in_payload_6_imag;
      data_in_7_real <= io_data_in_payload_7_real;
      data_in_7_imag <= io_data_in_payload_7_imag;
      data_in_8_real <= io_data_in_payload_8_real;
      data_in_8_imag <= io_data_in_payload_8_imag;
      data_in_9_real <= io_data_in_payload_9_real;
      data_in_9_imag <= io_data_in_payload_9_imag;
      data_in_10_real <= io_data_in_payload_10_real;
      data_in_10_imag <= io_data_in_payload_10_imag;
      data_in_11_real <= io_data_in_payload_11_real;
      data_in_11_imag <= io_data_in_payload_11_imag;
      data_in_12_real <= io_data_in_payload_12_real;
      data_in_12_imag <= io_data_in_payload_12_imag;
      data_in_13_real <= io_data_in_payload_13_real;
      data_in_13_imag <= io_data_in_payload_13_imag;
      data_in_14_real <= io_data_in_payload_14_real;
      data_in_14_imag <= io_data_in_payload_14_imag;
      data_in_15_real <= io_data_in_payload_15_real;
      data_in_15_imag <= io_data_in_payload_15_imag;
      data_in_16_real <= io_data_in_payload_16_real;
      data_in_16_imag <= io_data_in_payload_16_imag;
      data_in_17_real <= io_data_in_payload_17_real;
      data_in_17_imag <= io_data_in_payload_17_imag;
      data_in_18_real <= io_data_in_payload_18_real;
      data_in_18_imag <= io_data_in_payload_18_imag;
      data_in_19_real <= io_data_in_payload_19_real;
      data_in_19_imag <= io_data_in_payload_19_imag;
      data_in_20_real <= io_data_in_payload_20_real;
      data_in_20_imag <= io_data_in_payload_20_imag;
      data_in_21_real <= io_data_in_payload_21_real;
      data_in_21_imag <= io_data_in_payload_21_imag;
      data_in_22_real <= io_data_in_payload_22_real;
      data_in_22_imag <= io_data_in_payload_22_imag;
      data_in_23_real <= io_data_in_payload_23_real;
      data_in_23_imag <= io_data_in_payload_23_imag;
      data_in_24_real <= io_data_in_payload_24_real;
      data_in_24_imag <= io_data_in_payload_24_imag;
      data_in_25_real <= io_data_in_payload_25_real;
      data_in_25_imag <= io_data_in_payload_25_imag;
      data_in_26_real <= io_data_in_payload_26_real;
      data_in_26_imag <= io_data_in_payload_26_imag;
      data_in_27_real <= io_data_in_payload_27_real;
      data_in_27_imag <= io_data_in_payload_27_imag;
      data_in_28_real <= io_data_in_payload_28_real;
      data_in_28_imag <= io_data_in_payload_28_imag;
      data_in_29_real <= io_data_in_payload_29_real;
      data_in_29_imag <= io_data_in_payload_29_imag;
      data_in_30_real <= io_data_in_payload_30_real;
      data_in_30_imag <= io_data_in_payload_30_imag;
      data_in_31_real <= io_data_in_payload_31_real;
      data_in_31_imag <= io_data_in_payload_31_imag;
    end
    if((current_level_value == 3'b000))begin
      data_mid_0_real <= data_reorder_0_real;
      data_mid_0_imag <= data_reorder_0_imag;
      data_mid_1_real <= data_reorder_1_real;
      data_mid_1_imag <= data_reorder_1_imag;
      data_mid_2_real <= data_reorder_2_real;
      data_mid_2_imag <= data_reorder_2_imag;
      data_mid_3_real <= data_reorder_3_real;
      data_mid_3_imag <= data_reorder_3_imag;
      data_mid_4_real <= data_reorder_4_real;
      data_mid_4_imag <= data_reorder_4_imag;
      data_mid_5_real <= data_reorder_5_real;
      data_mid_5_imag <= data_reorder_5_imag;
      data_mid_6_real <= data_reorder_6_real;
      data_mid_6_imag <= data_reorder_6_imag;
      data_mid_7_real <= data_reorder_7_real;
      data_mid_7_imag <= data_reorder_7_imag;
      data_mid_8_real <= data_reorder_8_real;
      data_mid_8_imag <= data_reorder_8_imag;
      data_mid_9_real <= data_reorder_9_real;
      data_mid_9_imag <= data_reorder_9_imag;
      data_mid_10_real <= data_reorder_10_real;
      data_mid_10_imag <= data_reorder_10_imag;
      data_mid_11_real <= data_reorder_11_real;
      data_mid_11_imag <= data_reorder_11_imag;
      data_mid_12_real <= data_reorder_12_real;
      data_mid_12_imag <= data_reorder_12_imag;
      data_mid_13_real <= data_reorder_13_real;
      data_mid_13_imag <= data_reorder_13_imag;
      data_mid_14_real <= data_reorder_14_real;
      data_mid_14_imag <= data_reorder_14_imag;
      data_mid_15_real <= data_reorder_15_real;
      data_mid_15_imag <= data_reorder_15_imag;
      data_mid_16_real <= data_reorder_16_real;
      data_mid_16_imag <= data_reorder_16_imag;
      data_mid_17_real <= data_reorder_17_real;
      data_mid_17_imag <= data_reorder_17_imag;
      data_mid_18_real <= data_reorder_18_real;
      data_mid_18_imag <= data_reorder_18_imag;
      data_mid_19_real <= data_reorder_19_real;
      data_mid_19_imag <= data_reorder_19_imag;
      data_mid_20_real <= data_reorder_20_real;
      data_mid_20_imag <= data_reorder_20_imag;
      data_mid_21_real <= data_reorder_21_real;
      data_mid_21_imag <= data_reorder_21_imag;
      data_mid_22_real <= data_reorder_22_real;
      data_mid_22_imag <= data_reorder_22_imag;
      data_mid_23_real <= data_reorder_23_real;
      data_mid_23_imag <= data_reorder_23_imag;
      data_mid_24_real <= data_reorder_24_real;
      data_mid_24_imag <= data_reorder_24_imag;
      data_mid_25_real <= data_reorder_25_real;
      data_mid_25_imag <= data_reorder_25_imag;
      data_mid_26_real <= data_reorder_26_real;
      data_mid_26_imag <= data_reorder_26_imag;
      data_mid_27_real <= data_reorder_27_real;
      data_mid_27_imag <= data_reorder_27_imag;
      data_mid_28_real <= data_reorder_28_real;
      data_mid_28_imag <= data_reorder_28_imag;
      data_mid_29_real <= data_reorder_29_real;
      data_mid_29_imag <= data_reorder_29_imag;
      data_mid_30_real <= data_reorder_30_real;
      data_mid_30_imag <= data_reorder_30_imag;
      data_mid_31_real <= data_reorder_31_real;
      data_mid_31_imag <= data_reorder_31_imag;
    end else begin
      if((current_level_value == 3'b001))begin
        data_mid_1_real <= _zz_899[15 : 0];
        data_mid_1_imag <= _zz_907[15 : 0];
        data_mid_0_real <= _zz_915[15 : 0];
        data_mid_0_imag <= _zz_923[15 : 0];
      end
      if((current_level_value == 3'b001))begin
        data_mid_3_real <= _zz_940[15 : 0];
        data_mid_3_imag <= _zz_948[15 : 0];
        data_mid_2_real <= _zz_956[15 : 0];
        data_mid_2_imag <= _zz_964[15 : 0];
      end
      if((current_level_value == 3'b001))begin
        data_mid_5_real <= _zz_981[15 : 0];
        data_mid_5_imag <= _zz_989[15 : 0];
        data_mid_4_real <= _zz_997[15 : 0];
        data_mid_4_imag <= _zz_1005[15 : 0];
      end
      if((current_level_value == 3'b001))begin
        data_mid_7_real <= _zz_1022[15 : 0];
        data_mid_7_imag <= _zz_1030[15 : 0];
        data_mid_6_real <= _zz_1038[15 : 0];
        data_mid_6_imag <= _zz_1046[15 : 0];
      end
      if((current_level_value == 3'b001))begin
        data_mid_9_real <= _zz_1063[15 : 0];
        data_mid_9_imag <= _zz_1071[15 : 0];
        data_mid_8_real <= _zz_1079[15 : 0];
        data_mid_8_imag <= _zz_1087[15 : 0];
      end
      if((current_level_value == 3'b001))begin
        data_mid_11_real <= _zz_1104[15 : 0];
        data_mid_11_imag <= _zz_1112[15 : 0];
        data_mid_10_real <= _zz_1120[15 : 0];
        data_mid_10_imag <= _zz_1128[15 : 0];
      end
      if((current_level_value == 3'b001))begin
        data_mid_13_real <= _zz_1145[15 : 0];
        data_mid_13_imag <= _zz_1153[15 : 0];
        data_mid_12_real <= _zz_1161[15 : 0];
        data_mid_12_imag <= _zz_1169[15 : 0];
      end
      if((current_level_value == 3'b001))begin
        data_mid_15_real <= _zz_1186[15 : 0];
        data_mid_15_imag <= _zz_1194[15 : 0];
        data_mid_14_real <= _zz_1202[15 : 0];
        data_mid_14_imag <= _zz_1210[15 : 0];
      end
      if((current_level_value == 3'b001))begin
        data_mid_17_real <= _zz_1227[15 : 0];
        data_mid_17_imag <= _zz_1235[15 : 0];
        data_mid_16_real <= _zz_1243[15 : 0];
        data_mid_16_imag <= _zz_1251[15 : 0];
      end
      if((current_level_value == 3'b001))begin
        data_mid_19_real <= _zz_1268[15 : 0];
        data_mid_19_imag <= _zz_1276[15 : 0];
        data_mid_18_real <= _zz_1284[15 : 0];
        data_mid_18_imag <= _zz_1292[15 : 0];
      end
      if((current_level_value == 3'b001))begin
        data_mid_21_real <= _zz_1309[15 : 0];
        data_mid_21_imag <= _zz_1317[15 : 0];
        data_mid_20_real <= _zz_1325[15 : 0];
        data_mid_20_imag <= _zz_1333[15 : 0];
      end
      if((current_level_value == 3'b001))begin
        data_mid_23_real <= _zz_1350[15 : 0];
        data_mid_23_imag <= _zz_1358[15 : 0];
        data_mid_22_real <= _zz_1366[15 : 0];
        data_mid_22_imag <= _zz_1374[15 : 0];
      end
      if((current_level_value == 3'b001))begin
        data_mid_25_real <= _zz_1391[15 : 0];
        data_mid_25_imag <= _zz_1399[15 : 0];
        data_mid_24_real <= _zz_1407[15 : 0];
        data_mid_24_imag <= _zz_1415[15 : 0];
      end
      if((current_level_value == 3'b001))begin
        data_mid_27_real <= _zz_1432[15 : 0];
        data_mid_27_imag <= _zz_1440[15 : 0];
        data_mid_26_real <= _zz_1448[15 : 0];
        data_mid_26_imag <= _zz_1456[15 : 0];
      end
      if((current_level_value == 3'b001))begin
        data_mid_29_real <= _zz_1473[15 : 0];
        data_mid_29_imag <= _zz_1481[15 : 0];
        data_mid_28_real <= _zz_1489[15 : 0];
        data_mid_28_imag <= _zz_1497[15 : 0];
      end
      if((current_level_value == 3'b001))begin
        data_mid_31_real <= _zz_1514[15 : 0];
        data_mid_31_imag <= _zz_1522[15 : 0];
        data_mid_30_real <= _zz_1530[15 : 0];
        data_mid_30_imag <= _zz_1538[15 : 0];
      end
      if((current_level_value == 3'b010))begin
        data_mid_2_real <= _zz_1555[15 : 0];
        data_mid_2_imag <= _zz_1563[15 : 0];
        data_mid_0_real <= _zz_1571[15 : 0];
        data_mid_0_imag <= _zz_1579[15 : 0];
      end
      if((current_level_value == 3'b010))begin
        data_mid_3_real <= _zz_1596[15 : 0];
        data_mid_3_imag <= _zz_1604[15 : 0];
        data_mid_1_real <= _zz_1612[15 : 0];
        data_mid_1_imag <= _zz_1620[15 : 0];
      end
      if((current_level_value == 3'b010))begin
        data_mid_6_real <= _zz_1637[15 : 0];
        data_mid_6_imag <= _zz_1645[15 : 0];
        data_mid_4_real <= _zz_1653[15 : 0];
        data_mid_4_imag <= _zz_1661[15 : 0];
      end
      if((current_level_value == 3'b010))begin
        data_mid_7_real <= _zz_1678[15 : 0];
        data_mid_7_imag <= _zz_1686[15 : 0];
        data_mid_5_real <= _zz_1694[15 : 0];
        data_mid_5_imag <= _zz_1702[15 : 0];
      end
      if((current_level_value == 3'b010))begin
        data_mid_10_real <= _zz_1719[15 : 0];
        data_mid_10_imag <= _zz_1727[15 : 0];
        data_mid_8_real <= _zz_1735[15 : 0];
        data_mid_8_imag <= _zz_1743[15 : 0];
      end
      if((current_level_value == 3'b010))begin
        data_mid_11_real <= _zz_1760[15 : 0];
        data_mid_11_imag <= _zz_1768[15 : 0];
        data_mid_9_real <= _zz_1776[15 : 0];
        data_mid_9_imag <= _zz_1784[15 : 0];
      end
      if((current_level_value == 3'b010))begin
        data_mid_14_real <= _zz_1801[15 : 0];
        data_mid_14_imag <= _zz_1809[15 : 0];
        data_mid_12_real <= _zz_1817[15 : 0];
        data_mid_12_imag <= _zz_1825[15 : 0];
      end
      if((current_level_value == 3'b010))begin
        data_mid_15_real <= _zz_1842[15 : 0];
        data_mid_15_imag <= _zz_1850[15 : 0];
        data_mid_13_real <= _zz_1858[15 : 0];
        data_mid_13_imag <= _zz_1866[15 : 0];
      end
      if((current_level_value == 3'b010))begin
        data_mid_18_real <= _zz_1883[15 : 0];
        data_mid_18_imag <= _zz_1891[15 : 0];
        data_mid_16_real <= _zz_1899[15 : 0];
        data_mid_16_imag <= _zz_1907[15 : 0];
      end
      if((current_level_value == 3'b010))begin
        data_mid_19_real <= _zz_1924[15 : 0];
        data_mid_19_imag <= _zz_1932[15 : 0];
        data_mid_17_real <= _zz_1940[15 : 0];
        data_mid_17_imag <= _zz_1948[15 : 0];
      end
      if((current_level_value == 3'b010))begin
        data_mid_22_real <= _zz_1965[15 : 0];
        data_mid_22_imag <= _zz_1973[15 : 0];
        data_mid_20_real <= _zz_1981[15 : 0];
        data_mid_20_imag <= _zz_1989[15 : 0];
      end
      if((current_level_value == 3'b010))begin
        data_mid_23_real <= _zz_2006[15 : 0];
        data_mid_23_imag <= _zz_2014[15 : 0];
        data_mid_21_real <= _zz_2022[15 : 0];
        data_mid_21_imag <= _zz_2030[15 : 0];
      end
      if((current_level_value == 3'b010))begin
        data_mid_26_real <= _zz_2047[15 : 0];
        data_mid_26_imag <= _zz_2055[15 : 0];
        data_mid_24_real <= _zz_2063[15 : 0];
        data_mid_24_imag <= _zz_2071[15 : 0];
      end
      if((current_level_value == 3'b010))begin
        data_mid_27_real <= _zz_2088[15 : 0];
        data_mid_27_imag <= _zz_2096[15 : 0];
        data_mid_25_real <= _zz_2104[15 : 0];
        data_mid_25_imag <= _zz_2112[15 : 0];
      end
      if((current_level_value == 3'b010))begin
        data_mid_30_real <= _zz_2129[15 : 0];
        data_mid_30_imag <= _zz_2137[15 : 0];
        data_mid_28_real <= _zz_2145[15 : 0];
        data_mid_28_imag <= _zz_2153[15 : 0];
      end
      if((current_level_value == 3'b010))begin
        data_mid_31_real <= _zz_2170[15 : 0];
        data_mid_31_imag <= _zz_2178[15 : 0];
        data_mid_29_real <= _zz_2186[15 : 0];
        data_mid_29_imag <= _zz_2194[15 : 0];
      end
      if((current_level_value == 3'b011))begin
        data_mid_4_real <= _zz_2211[15 : 0];
        data_mid_4_imag <= _zz_2219[15 : 0];
        data_mid_0_real <= _zz_2227[15 : 0];
        data_mid_0_imag <= _zz_2235[15 : 0];
      end
      if((current_level_value == 3'b011))begin
        data_mid_5_real <= _zz_2252[15 : 0];
        data_mid_5_imag <= _zz_2260[15 : 0];
        data_mid_1_real <= _zz_2268[15 : 0];
        data_mid_1_imag <= _zz_2276[15 : 0];
      end
      if((current_level_value == 3'b011))begin
        data_mid_6_real <= _zz_2293[15 : 0];
        data_mid_6_imag <= _zz_2301[15 : 0];
        data_mid_2_real <= _zz_2309[15 : 0];
        data_mid_2_imag <= _zz_2317[15 : 0];
      end
      if((current_level_value == 3'b011))begin
        data_mid_7_real <= _zz_2334[15 : 0];
        data_mid_7_imag <= _zz_2342[15 : 0];
        data_mid_3_real <= _zz_2350[15 : 0];
        data_mid_3_imag <= _zz_2358[15 : 0];
      end
      if((current_level_value == 3'b011))begin
        data_mid_12_real <= _zz_2375[15 : 0];
        data_mid_12_imag <= _zz_2383[15 : 0];
        data_mid_8_real <= _zz_2391[15 : 0];
        data_mid_8_imag <= _zz_2399[15 : 0];
      end
      if((current_level_value == 3'b011))begin
        data_mid_13_real <= _zz_2416[15 : 0];
        data_mid_13_imag <= _zz_2424[15 : 0];
        data_mid_9_real <= _zz_2432[15 : 0];
        data_mid_9_imag <= _zz_2440[15 : 0];
      end
      if((current_level_value == 3'b011))begin
        data_mid_14_real <= _zz_2457[15 : 0];
        data_mid_14_imag <= _zz_2465[15 : 0];
        data_mid_10_real <= _zz_2473[15 : 0];
        data_mid_10_imag <= _zz_2481[15 : 0];
      end
      if((current_level_value == 3'b011))begin
        data_mid_15_real <= _zz_2498[15 : 0];
        data_mid_15_imag <= _zz_2506[15 : 0];
        data_mid_11_real <= _zz_2514[15 : 0];
        data_mid_11_imag <= _zz_2522[15 : 0];
      end
      if((current_level_value == 3'b011))begin
        data_mid_20_real <= _zz_2539[15 : 0];
        data_mid_20_imag <= _zz_2547[15 : 0];
        data_mid_16_real <= _zz_2555[15 : 0];
        data_mid_16_imag <= _zz_2563[15 : 0];
      end
      if((current_level_value == 3'b011))begin
        data_mid_21_real <= _zz_2580[15 : 0];
        data_mid_21_imag <= _zz_2588[15 : 0];
        data_mid_17_real <= _zz_2596[15 : 0];
        data_mid_17_imag <= _zz_2604[15 : 0];
      end
      if((current_level_value == 3'b011))begin
        data_mid_22_real <= _zz_2621[15 : 0];
        data_mid_22_imag <= _zz_2629[15 : 0];
        data_mid_18_real <= _zz_2637[15 : 0];
        data_mid_18_imag <= _zz_2645[15 : 0];
      end
      if((current_level_value == 3'b011))begin
        data_mid_23_real <= _zz_2662[15 : 0];
        data_mid_23_imag <= _zz_2670[15 : 0];
        data_mid_19_real <= _zz_2678[15 : 0];
        data_mid_19_imag <= _zz_2686[15 : 0];
      end
      if((current_level_value == 3'b011))begin
        data_mid_28_real <= _zz_2703[15 : 0];
        data_mid_28_imag <= _zz_2711[15 : 0];
        data_mid_24_real <= _zz_2719[15 : 0];
        data_mid_24_imag <= _zz_2727[15 : 0];
      end
      if((current_level_value == 3'b011))begin
        data_mid_29_real <= _zz_2744[15 : 0];
        data_mid_29_imag <= _zz_2752[15 : 0];
        data_mid_25_real <= _zz_2760[15 : 0];
        data_mid_25_imag <= _zz_2768[15 : 0];
      end
      if((current_level_value == 3'b011))begin
        data_mid_30_real <= _zz_2785[15 : 0];
        data_mid_30_imag <= _zz_2793[15 : 0];
        data_mid_26_real <= _zz_2801[15 : 0];
        data_mid_26_imag <= _zz_2809[15 : 0];
      end
      if((current_level_value == 3'b011))begin
        data_mid_31_real <= _zz_2826[15 : 0];
        data_mid_31_imag <= _zz_2834[15 : 0];
        data_mid_27_real <= _zz_2842[15 : 0];
        data_mid_27_imag <= _zz_2850[15 : 0];
      end
      if((current_level_value == 3'b100))begin
        data_mid_8_real <= _zz_2867[15 : 0];
        data_mid_8_imag <= _zz_2875[15 : 0];
        data_mid_0_real <= _zz_2883[15 : 0];
        data_mid_0_imag <= _zz_2891[15 : 0];
      end
      if((current_level_value == 3'b100))begin
        data_mid_9_real <= _zz_2908[15 : 0];
        data_mid_9_imag <= _zz_2916[15 : 0];
        data_mid_1_real <= _zz_2924[15 : 0];
        data_mid_1_imag <= _zz_2932[15 : 0];
      end
      if((current_level_value == 3'b100))begin
        data_mid_10_real <= _zz_2949[15 : 0];
        data_mid_10_imag <= _zz_2957[15 : 0];
        data_mid_2_real <= _zz_2965[15 : 0];
        data_mid_2_imag <= _zz_2973[15 : 0];
      end
      if((current_level_value == 3'b100))begin
        data_mid_11_real <= _zz_2990[15 : 0];
        data_mid_11_imag <= _zz_2998[15 : 0];
        data_mid_3_real <= _zz_3006[15 : 0];
        data_mid_3_imag <= _zz_3014[15 : 0];
      end
      if((current_level_value == 3'b100))begin
        data_mid_12_real <= _zz_3031[15 : 0];
        data_mid_12_imag <= _zz_3039[15 : 0];
        data_mid_4_real <= _zz_3047[15 : 0];
        data_mid_4_imag <= _zz_3055[15 : 0];
      end
      if((current_level_value == 3'b100))begin
        data_mid_13_real <= _zz_3072[15 : 0];
        data_mid_13_imag <= _zz_3080[15 : 0];
        data_mid_5_real <= _zz_3088[15 : 0];
        data_mid_5_imag <= _zz_3096[15 : 0];
      end
      if((current_level_value == 3'b100))begin
        data_mid_14_real <= _zz_3113[15 : 0];
        data_mid_14_imag <= _zz_3121[15 : 0];
        data_mid_6_real <= _zz_3129[15 : 0];
        data_mid_6_imag <= _zz_3137[15 : 0];
      end
      if((current_level_value == 3'b100))begin
        data_mid_15_real <= _zz_3154[15 : 0];
        data_mid_15_imag <= _zz_3162[15 : 0];
        data_mid_7_real <= _zz_3170[15 : 0];
        data_mid_7_imag <= _zz_3178[15 : 0];
      end
      if((current_level_value == 3'b100))begin
        data_mid_24_real <= _zz_3195[15 : 0];
        data_mid_24_imag <= _zz_3203[15 : 0];
        data_mid_16_real <= _zz_3211[15 : 0];
        data_mid_16_imag <= _zz_3219[15 : 0];
      end
      if((current_level_value == 3'b100))begin
        data_mid_25_real <= _zz_3236[15 : 0];
        data_mid_25_imag <= _zz_3244[15 : 0];
        data_mid_17_real <= _zz_3252[15 : 0];
        data_mid_17_imag <= _zz_3260[15 : 0];
      end
      if((current_level_value == 3'b100))begin
        data_mid_26_real <= _zz_3277[15 : 0];
        data_mid_26_imag <= _zz_3285[15 : 0];
        data_mid_18_real <= _zz_3293[15 : 0];
        data_mid_18_imag <= _zz_3301[15 : 0];
      end
      if((current_level_value == 3'b100))begin
        data_mid_27_real <= _zz_3318[15 : 0];
        data_mid_27_imag <= _zz_3326[15 : 0];
        data_mid_19_real <= _zz_3334[15 : 0];
        data_mid_19_imag <= _zz_3342[15 : 0];
      end
      if((current_level_value == 3'b100))begin
        data_mid_28_real <= _zz_3359[15 : 0];
        data_mid_28_imag <= _zz_3367[15 : 0];
        data_mid_20_real <= _zz_3375[15 : 0];
        data_mid_20_imag <= _zz_3383[15 : 0];
      end
      if((current_level_value == 3'b100))begin
        data_mid_29_real <= _zz_3400[15 : 0];
        data_mid_29_imag <= _zz_3408[15 : 0];
        data_mid_21_real <= _zz_3416[15 : 0];
        data_mid_21_imag <= _zz_3424[15 : 0];
      end
      if((current_level_value == 3'b100))begin
        data_mid_30_real <= _zz_3441[15 : 0];
        data_mid_30_imag <= _zz_3449[15 : 0];
        data_mid_22_real <= _zz_3457[15 : 0];
        data_mid_22_imag <= _zz_3465[15 : 0];
      end
      if((current_level_value == 3'b100))begin
        data_mid_31_real <= _zz_3482[15 : 0];
        data_mid_31_imag <= _zz_3490[15 : 0];
        data_mid_23_real <= _zz_3498[15 : 0];
        data_mid_23_imag <= _zz_3506[15 : 0];
      end
      if((current_level_value == 3'b101))begin
        data_mid_16_real <= _zz_3523[15 : 0];
        data_mid_16_imag <= _zz_3531[15 : 0];
        data_mid_0_real <= _zz_3539[15 : 0];
        data_mid_0_imag <= _zz_3547[15 : 0];
      end
      if((current_level_value == 3'b101))begin
        data_mid_17_real <= _zz_3564[15 : 0];
        data_mid_17_imag <= _zz_3572[15 : 0];
        data_mid_1_real <= _zz_3580[15 : 0];
        data_mid_1_imag <= _zz_3588[15 : 0];
      end
      if((current_level_value == 3'b101))begin
        data_mid_18_real <= _zz_3605[15 : 0];
        data_mid_18_imag <= _zz_3613[15 : 0];
        data_mid_2_real <= _zz_3621[15 : 0];
        data_mid_2_imag <= _zz_3629[15 : 0];
      end
      if((current_level_value == 3'b101))begin
        data_mid_19_real <= _zz_3646[15 : 0];
        data_mid_19_imag <= _zz_3654[15 : 0];
        data_mid_3_real <= _zz_3662[15 : 0];
        data_mid_3_imag <= _zz_3670[15 : 0];
      end
      if((current_level_value == 3'b101))begin
        data_mid_20_real <= _zz_3687[15 : 0];
        data_mid_20_imag <= _zz_3695[15 : 0];
        data_mid_4_real <= _zz_3703[15 : 0];
        data_mid_4_imag <= _zz_3711[15 : 0];
      end
      if((current_level_value == 3'b101))begin
        data_mid_21_real <= _zz_3728[15 : 0];
        data_mid_21_imag <= _zz_3736[15 : 0];
        data_mid_5_real <= _zz_3744[15 : 0];
        data_mid_5_imag <= _zz_3752[15 : 0];
      end
      if((current_level_value == 3'b101))begin
        data_mid_22_real <= _zz_3769[15 : 0];
        data_mid_22_imag <= _zz_3777[15 : 0];
        data_mid_6_real <= _zz_3785[15 : 0];
        data_mid_6_imag <= _zz_3793[15 : 0];
      end
      if((current_level_value == 3'b101))begin
        data_mid_23_real <= _zz_3810[15 : 0];
        data_mid_23_imag <= _zz_3818[15 : 0];
        data_mid_7_real <= _zz_3826[15 : 0];
        data_mid_7_imag <= _zz_3834[15 : 0];
      end
      if((current_level_value == 3'b101))begin
        data_mid_24_real <= _zz_3851[15 : 0];
        data_mid_24_imag <= _zz_3859[15 : 0];
        data_mid_8_real <= _zz_3867[15 : 0];
        data_mid_8_imag <= _zz_3875[15 : 0];
      end
      if((current_level_value == 3'b101))begin
        data_mid_25_real <= _zz_3892[15 : 0];
        data_mid_25_imag <= _zz_3900[15 : 0];
        data_mid_9_real <= _zz_3908[15 : 0];
        data_mid_9_imag <= _zz_3916[15 : 0];
      end
      if((current_level_value == 3'b101))begin
        data_mid_26_real <= _zz_3933[15 : 0];
        data_mid_26_imag <= _zz_3941[15 : 0];
        data_mid_10_real <= _zz_3949[15 : 0];
        data_mid_10_imag <= _zz_3957[15 : 0];
      end
      if((current_level_value == 3'b101))begin
        data_mid_27_real <= _zz_3974[15 : 0];
        data_mid_27_imag <= _zz_3982[15 : 0];
        data_mid_11_real <= _zz_3990[15 : 0];
        data_mid_11_imag <= _zz_3998[15 : 0];
      end
      if((current_level_value == 3'b101))begin
        data_mid_28_real <= _zz_4015[15 : 0];
        data_mid_28_imag <= _zz_4023[15 : 0];
        data_mid_12_real <= _zz_4031[15 : 0];
        data_mid_12_imag <= _zz_4039[15 : 0];
      end
      if((current_level_value == 3'b101))begin
        data_mid_29_real <= _zz_4056[15 : 0];
        data_mid_29_imag <= _zz_4064[15 : 0];
        data_mid_13_real <= _zz_4072[15 : 0];
        data_mid_13_imag <= _zz_4080[15 : 0];
      end
      if((current_level_value == 3'b101))begin
        data_mid_30_real <= _zz_4097[15 : 0];
        data_mid_30_imag <= _zz_4105[15 : 0];
        data_mid_14_real <= _zz_4113[15 : 0];
        data_mid_14_imag <= _zz_4121[15 : 0];
      end
      if((current_level_value == 3'b101))begin
        data_mid_31_real <= _zz_4138[15 : 0];
        data_mid_31_imag <= _zz_4146[15 : 0];
        data_mid_15_real <= _zz_4154[15 : 0];
        data_mid_15_imag <= _zz_4162[15 : 0];
      end
    end
  end

  always @ (posedge clk or posedge reset) begin
    if (reset) begin
      io_data_in_valid_regNext <= 1'b0;
      current_level_value <= 3'b000;
      null_cond_period_minus_1 <= 1'b0;
      current_level_willOverflow_regNext <= 1'b0;
    end else begin
      io_data_in_valid_regNext <= io_data_in_valid;
      current_level_value <= current_level_valueNext;
      if(io_data_in_valid_regNext)begin
        null_cond_period_minus_1 <= 1'b1;
      end else begin
        if(current_level_willOverflow)begin
          null_cond_period_minus_1 <= 1'b0;
        end
      end
      current_level_willOverflow_regNext <= current_level_willOverflow;
    end
  end


endmodule

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

module SInt32fixTo23_8_ROUNDTOINF (
  input      [31:0]   din,
  output     [15:0]   dout
);
  wire       [32:0]   _zz_9;
  wire       [32:0]   _zz_10;
  wire       [7:0]    _zz_11;
  wire       [24:0]   _zz_12;
  wire       [24:0]   _zz_13;
  wire       [32:0]   _zz_14;
  wire       [32:0]   _zz_15;
  wire       [32:0]   _zz_16;
  wire       [9:0]    _zz_17;
  wire       [8:0]    _zz_18;
  reg        [24:0]   _zz_1;
  wire       [31:0]   _zz_2;
  wire       [31:0]   _zz_3;
  wire       [31:0]   _zz_4;
  wire       [32:0]   _zz_5;
  wire       [31:0]   _zz_6;
  reg        [24:0]   _zz_7;
  reg        [15:0]   _zz_8;

  assign _zz_9 = {_zz_4[31],_zz_4};
  assign _zz_10 = {_zz_3[31],_zz_3};
  assign _zz_11 = _zz_5[7 : 0];
  assign _zz_12 = _zz_5[32 : 8];
  assign _zz_13 = 25'h0000001;
  assign _zz_14 = ($signed(_zz_15) + $signed(_zz_16));
  assign _zz_15 = {_zz_6[31],_zz_6};
  assign _zz_16 = {_zz_2[31],_zz_2};
  assign _zz_17 = _zz_1[24 : 15];
  assign _zz_18 = _zz_1[23 : 15];
  assign _zz_2 = {{24'h0,1'b1},7'h0};
  assign _zz_3 = {25'h1ffffff,7'h0};
  assign _zz_4 = din[31 : 0];
  assign _zz_5 = ($signed(_zz_9) + $signed(_zz_10));
  assign _zz_6 = din[31 : 0];
  always @ (*) begin
    if((_zz_11 != 8'h0))begin
      _zz_7 = ($signed(_zz_12) + $signed(_zz_13));
    end else begin
      _zz_7 = _zz_5[32 : 8];
    end
  end

  always @ (*) begin
    if(_zz_5[32])begin
      _zz_1 = _zz_7;
    end else begin
      _zz_1 = (_zz_14 >>> 8);
    end
  end

  always @ (*) begin
    if(_zz_1[24])begin
      if((! (_zz_17 == 10'h3ff)))begin
        _zz_8 = 16'h8000;
      end else begin
        _zz_8 = _zz_1[15 : 0];
      end
    end else begin
      if((_zz_18 != 9'h0))begin
        _zz_8 = 16'h7fff;
      end else begin
        _zz_8 = _zz_1[15 : 0];
      end
    end
  end

  assign dout = _zz_8;

endmodule

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

module SInt32fixTo31_0_ROUNDTOINF (
  input      [31:0]   din,
  output     [31:0]   dout
);

  assign dout = din;

endmodule
