// Generator : SpinalHDL v1.4.0    git head : ecb5a80b713566f417ea3ea061f9969e73770a7f
// Date      : 20/05/2020, 17:00:35
// Component : CoefLoadUnit



module CoefLoadUnit (
  input               _zz_1_,
  output              _zz_2_,
  input      [31:0]   _zz_3_,
  input      [3:0]    _zz_4_,
  input      [7:0]    _zz_5_,
  input      [1:0]    _zz_6_,
  input               _zz_7_,
  output              _zz_8_,
  input      [31:0]   _zz_9_,
  output              _zz_10_,
  output     [3:0]    _zz_11_,
  output     [1:0]    _zz_12_,
  output              io_coef_out_valid,
  output     [15:0]   io_coef_out_payload_0_0_0_real,
  output     [15:0]   io_coef_out_payload_0_0_0_imag,
  output     [15:0]   io_coef_out_payload_0_0_1_real,
  output     [15:0]   io_coef_out_payload_0_0_1_imag,
  output     [15:0]   io_coef_out_payload_0_0_2_real,
  output     [15:0]   io_coef_out_payload_0_0_2_imag,
  output     [15:0]   io_coef_out_payload_0_0_3_real,
  output     [15:0]   io_coef_out_payload_0_0_3_imag,
  output     [15:0]   io_coef_out_payload_0_0_4_real,
  output     [15:0]   io_coef_out_payload_0_0_4_imag,
  output     [15:0]   io_coef_out_payload_0_0_5_real,
  output     [15:0]   io_coef_out_payload_0_0_5_imag,
  output     [15:0]   io_coef_out_payload_0_0_6_real,
  output     [15:0]   io_coef_out_payload_0_0_6_imag,
  output     [15:0]   io_coef_out_payload_0_0_7_real,
  output     [15:0]   io_coef_out_payload_0_0_7_imag,
  output     [15:0]   io_coef_out_payload_0_0_8_real,
  output     [15:0]   io_coef_out_payload_0_0_8_imag,
  output     [15:0]   io_coef_out_payload_0_0_9_real,
  output     [15:0]   io_coef_out_payload_0_0_9_imag,
  output     [15:0]   io_coef_out_payload_0_0_10_real,
  output     [15:0]   io_coef_out_payload_0_0_10_imag,
  output     [15:0]   io_coef_out_payload_0_0_11_real,
  output     [15:0]   io_coef_out_payload_0_0_11_imag,
  output     [15:0]   io_coef_out_payload_0_0_12_real,
  output     [15:0]   io_coef_out_payload_0_0_12_imag,
  output     [15:0]   io_coef_out_payload_0_0_13_real,
  output     [15:0]   io_coef_out_payload_0_0_13_imag,
  output     [15:0]   io_coef_out_payload_0_0_14_real,
  output     [15:0]   io_coef_out_payload_0_0_14_imag,
  output     [15:0]   io_coef_out_payload_0_0_15_real,
  output     [15:0]   io_coef_out_payload_0_0_15_imag,
  output     [15:0]   io_coef_out_payload_0_0_16_real,
  output     [15:0]   io_coef_out_payload_0_0_16_imag,
  output     [15:0]   io_coef_out_payload_0_0_17_real,
  output     [15:0]   io_coef_out_payload_0_0_17_imag,
  output     [15:0]   io_coef_out_payload_0_0_18_real,
  output     [15:0]   io_coef_out_payload_0_0_18_imag,
  output     [15:0]   io_coef_out_payload_0_0_19_real,
  output     [15:0]   io_coef_out_payload_0_0_19_imag,
  output     [15:0]   io_coef_out_payload_0_0_20_real,
  output     [15:0]   io_coef_out_payload_0_0_20_imag,
  output     [15:0]   io_coef_out_payload_0_0_21_real,
  output     [15:0]   io_coef_out_payload_0_0_21_imag,
  output     [15:0]   io_coef_out_payload_0_0_22_real,
  output     [15:0]   io_coef_out_payload_0_0_22_imag,
  output     [15:0]   io_coef_out_payload_0_0_23_real,
  output     [15:0]   io_coef_out_payload_0_0_23_imag,
  output     [15:0]   io_coef_out_payload_0_0_24_real,
  output     [15:0]   io_coef_out_payload_0_0_24_imag,
  output     [15:0]   io_coef_out_payload_0_0_25_real,
  output     [15:0]   io_coef_out_payload_0_0_25_imag,
  output     [15:0]   io_coef_out_payload_0_0_26_real,
  output     [15:0]   io_coef_out_payload_0_0_26_imag,
  output     [15:0]   io_coef_out_payload_0_0_27_real,
  output     [15:0]   io_coef_out_payload_0_0_27_imag,
  output     [15:0]   io_coef_out_payload_0_0_28_real,
  output     [15:0]   io_coef_out_payload_0_0_28_imag,
  output     [15:0]   io_coef_out_payload_0_0_29_real,
  output     [15:0]   io_coef_out_payload_0_0_29_imag,
  output     [15:0]   io_coef_out_payload_0_0_30_real,
  output     [15:0]   io_coef_out_payload_0_0_30_imag,
  output     [15:0]   io_coef_out_payload_0_0_31_real,
  output     [15:0]   io_coef_out_payload_0_0_31_imag,
  output     [15:0]   io_coef_out_payload_0_0_32_real,
  output     [15:0]   io_coef_out_payload_0_0_32_imag,
  output     [15:0]   io_coef_out_payload_0_0_33_real,
  output     [15:0]   io_coef_out_payload_0_0_33_imag,
  output     [15:0]   io_coef_out_payload_0_0_34_real,
  output     [15:0]   io_coef_out_payload_0_0_34_imag,
  output     [15:0]   io_coef_out_payload_0_0_35_real,
  output     [15:0]   io_coef_out_payload_0_0_35_imag,
  output     [15:0]   io_coef_out_payload_0_0_36_real,
  output     [15:0]   io_coef_out_payload_0_0_36_imag,
  output     [15:0]   io_coef_out_payload_0_0_37_real,
  output     [15:0]   io_coef_out_payload_0_0_37_imag,
  output     [15:0]   io_coef_out_payload_0_0_38_real,
  output     [15:0]   io_coef_out_payload_0_0_38_imag,
  output     [15:0]   io_coef_out_payload_0_0_39_real,
  output     [15:0]   io_coef_out_payload_0_0_39_imag,
  output     [15:0]   io_coef_out_payload_0_0_40_real,
  output     [15:0]   io_coef_out_payload_0_0_40_imag,
  output     [15:0]   io_coef_out_payload_0_0_41_real,
  output     [15:0]   io_coef_out_payload_0_0_41_imag,
  output     [15:0]   io_coef_out_payload_0_0_42_real,
  output     [15:0]   io_coef_out_payload_0_0_42_imag,
  output     [15:0]   io_coef_out_payload_0_0_43_real,
  output     [15:0]   io_coef_out_payload_0_0_43_imag,
  output     [15:0]   io_coef_out_payload_0_0_44_real,
  output     [15:0]   io_coef_out_payload_0_0_44_imag,
  output     [15:0]   io_coef_out_payload_0_0_45_real,
  output     [15:0]   io_coef_out_payload_0_0_45_imag,
  output     [15:0]   io_coef_out_payload_0_0_46_real,
  output     [15:0]   io_coef_out_payload_0_0_46_imag,
  output     [15:0]   io_coef_out_payload_0_0_47_real,
  output     [15:0]   io_coef_out_payload_0_0_47_imag,
  output     [15:0]   io_coef_out_payload_0_0_48_real,
  output     [15:0]   io_coef_out_payload_0_0_48_imag,
  output     [15:0]   io_coef_out_payload_0_0_49_real,
  output     [15:0]   io_coef_out_payload_0_0_49_imag,
  output     [15:0]   io_coef_out_payload_0_1_0_real,
  output     [15:0]   io_coef_out_payload_0_1_0_imag,
  output     [15:0]   io_coef_out_payload_0_1_1_real,
  output     [15:0]   io_coef_out_payload_0_1_1_imag,
  output     [15:0]   io_coef_out_payload_0_1_2_real,
  output     [15:0]   io_coef_out_payload_0_1_2_imag,
  output     [15:0]   io_coef_out_payload_0_1_3_real,
  output     [15:0]   io_coef_out_payload_0_1_3_imag,
  output     [15:0]   io_coef_out_payload_0_1_4_real,
  output     [15:0]   io_coef_out_payload_0_1_4_imag,
  output     [15:0]   io_coef_out_payload_0_1_5_real,
  output     [15:0]   io_coef_out_payload_0_1_5_imag,
  output     [15:0]   io_coef_out_payload_0_1_6_real,
  output     [15:0]   io_coef_out_payload_0_1_6_imag,
  output     [15:0]   io_coef_out_payload_0_1_7_real,
  output     [15:0]   io_coef_out_payload_0_1_7_imag,
  output     [15:0]   io_coef_out_payload_0_1_8_real,
  output     [15:0]   io_coef_out_payload_0_1_8_imag,
  output     [15:0]   io_coef_out_payload_0_1_9_real,
  output     [15:0]   io_coef_out_payload_0_1_9_imag,
  output     [15:0]   io_coef_out_payload_0_1_10_real,
  output     [15:0]   io_coef_out_payload_0_1_10_imag,
  output     [15:0]   io_coef_out_payload_0_1_11_real,
  output     [15:0]   io_coef_out_payload_0_1_11_imag,
  output     [15:0]   io_coef_out_payload_0_1_12_real,
  output     [15:0]   io_coef_out_payload_0_1_12_imag,
  output     [15:0]   io_coef_out_payload_0_1_13_real,
  output     [15:0]   io_coef_out_payload_0_1_13_imag,
  output     [15:0]   io_coef_out_payload_0_1_14_real,
  output     [15:0]   io_coef_out_payload_0_1_14_imag,
  output     [15:0]   io_coef_out_payload_0_1_15_real,
  output     [15:0]   io_coef_out_payload_0_1_15_imag,
  output     [15:0]   io_coef_out_payload_0_1_16_real,
  output     [15:0]   io_coef_out_payload_0_1_16_imag,
  output     [15:0]   io_coef_out_payload_0_1_17_real,
  output     [15:0]   io_coef_out_payload_0_1_17_imag,
  output     [15:0]   io_coef_out_payload_0_1_18_real,
  output     [15:0]   io_coef_out_payload_0_1_18_imag,
  output     [15:0]   io_coef_out_payload_0_1_19_real,
  output     [15:0]   io_coef_out_payload_0_1_19_imag,
  output     [15:0]   io_coef_out_payload_0_1_20_real,
  output     [15:0]   io_coef_out_payload_0_1_20_imag,
  output     [15:0]   io_coef_out_payload_0_1_21_real,
  output     [15:0]   io_coef_out_payload_0_1_21_imag,
  output     [15:0]   io_coef_out_payload_0_1_22_real,
  output     [15:0]   io_coef_out_payload_0_1_22_imag,
  output     [15:0]   io_coef_out_payload_0_1_23_real,
  output     [15:0]   io_coef_out_payload_0_1_23_imag,
  output     [15:0]   io_coef_out_payload_0_1_24_real,
  output     [15:0]   io_coef_out_payload_0_1_24_imag,
  output     [15:0]   io_coef_out_payload_0_1_25_real,
  output     [15:0]   io_coef_out_payload_0_1_25_imag,
  output     [15:0]   io_coef_out_payload_0_1_26_real,
  output     [15:0]   io_coef_out_payload_0_1_26_imag,
  output     [15:0]   io_coef_out_payload_0_1_27_real,
  output     [15:0]   io_coef_out_payload_0_1_27_imag,
  output     [15:0]   io_coef_out_payload_0_1_28_real,
  output     [15:0]   io_coef_out_payload_0_1_28_imag,
  output     [15:0]   io_coef_out_payload_0_1_29_real,
  output     [15:0]   io_coef_out_payload_0_1_29_imag,
  output     [15:0]   io_coef_out_payload_0_1_30_real,
  output     [15:0]   io_coef_out_payload_0_1_30_imag,
  output     [15:0]   io_coef_out_payload_0_1_31_real,
  output     [15:0]   io_coef_out_payload_0_1_31_imag,
  output     [15:0]   io_coef_out_payload_0_1_32_real,
  output     [15:0]   io_coef_out_payload_0_1_32_imag,
  output     [15:0]   io_coef_out_payload_0_1_33_real,
  output     [15:0]   io_coef_out_payload_0_1_33_imag,
  output     [15:0]   io_coef_out_payload_0_1_34_real,
  output     [15:0]   io_coef_out_payload_0_1_34_imag,
  output     [15:0]   io_coef_out_payload_0_1_35_real,
  output     [15:0]   io_coef_out_payload_0_1_35_imag,
  output     [15:0]   io_coef_out_payload_0_1_36_real,
  output     [15:0]   io_coef_out_payload_0_1_36_imag,
  output     [15:0]   io_coef_out_payload_0_1_37_real,
  output     [15:0]   io_coef_out_payload_0_1_37_imag,
  output     [15:0]   io_coef_out_payload_0_1_38_real,
  output     [15:0]   io_coef_out_payload_0_1_38_imag,
  output     [15:0]   io_coef_out_payload_0_1_39_real,
  output     [15:0]   io_coef_out_payload_0_1_39_imag,
  output     [15:0]   io_coef_out_payload_0_1_40_real,
  output     [15:0]   io_coef_out_payload_0_1_40_imag,
  output     [15:0]   io_coef_out_payload_0_1_41_real,
  output     [15:0]   io_coef_out_payload_0_1_41_imag,
  output     [15:0]   io_coef_out_payload_0_1_42_real,
  output     [15:0]   io_coef_out_payload_0_1_42_imag,
  output     [15:0]   io_coef_out_payload_0_1_43_real,
  output     [15:0]   io_coef_out_payload_0_1_43_imag,
  output     [15:0]   io_coef_out_payload_0_1_44_real,
  output     [15:0]   io_coef_out_payload_0_1_44_imag,
  output     [15:0]   io_coef_out_payload_0_1_45_real,
  output     [15:0]   io_coef_out_payload_0_1_45_imag,
  output     [15:0]   io_coef_out_payload_0_1_46_real,
  output     [15:0]   io_coef_out_payload_0_1_46_imag,
  output     [15:0]   io_coef_out_payload_0_1_47_real,
  output     [15:0]   io_coef_out_payload_0_1_47_imag,
  output     [15:0]   io_coef_out_payload_0_1_48_real,
  output     [15:0]   io_coef_out_payload_0_1_48_imag,
  output     [15:0]   io_coef_out_payload_0_1_49_real,
  output     [15:0]   io_coef_out_payload_0_1_49_imag,
  output     [15:0]   io_coef_out_payload_0_2_0_real,
  output     [15:0]   io_coef_out_payload_0_2_0_imag,
  output     [15:0]   io_coef_out_payload_0_2_1_real,
  output     [15:0]   io_coef_out_payload_0_2_1_imag,
  output     [15:0]   io_coef_out_payload_0_2_2_real,
  output     [15:0]   io_coef_out_payload_0_2_2_imag,
  output     [15:0]   io_coef_out_payload_0_2_3_real,
  output     [15:0]   io_coef_out_payload_0_2_3_imag,
  output     [15:0]   io_coef_out_payload_0_2_4_real,
  output     [15:0]   io_coef_out_payload_0_2_4_imag,
  output     [15:0]   io_coef_out_payload_0_2_5_real,
  output     [15:0]   io_coef_out_payload_0_2_5_imag,
  output     [15:0]   io_coef_out_payload_0_2_6_real,
  output     [15:0]   io_coef_out_payload_0_2_6_imag,
  output     [15:0]   io_coef_out_payload_0_2_7_real,
  output     [15:0]   io_coef_out_payload_0_2_7_imag,
  output     [15:0]   io_coef_out_payload_0_2_8_real,
  output     [15:0]   io_coef_out_payload_0_2_8_imag,
  output     [15:0]   io_coef_out_payload_0_2_9_real,
  output     [15:0]   io_coef_out_payload_0_2_9_imag,
  output     [15:0]   io_coef_out_payload_0_2_10_real,
  output     [15:0]   io_coef_out_payload_0_2_10_imag,
  output     [15:0]   io_coef_out_payload_0_2_11_real,
  output     [15:0]   io_coef_out_payload_0_2_11_imag,
  output     [15:0]   io_coef_out_payload_0_2_12_real,
  output     [15:0]   io_coef_out_payload_0_2_12_imag,
  output     [15:0]   io_coef_out_payload_0_2_13_real,
  output     [15:0]   io_coef_out_payload_0_2_13_imag,
  output     [15:0]   io_coef_out_payload_0_2_14_real,
  output     [15:0]   io_coef_out_payload_0_2_14_imag,
  output     [15:0]   io_coef_out_payload_0_2_15_real,
  output     [15:0]   io_coef_out_payload_0_2_15_imag,
  output     [15:0]   io_coef_out_payload_0_2_16_real,
  output     [15:0]   io_coef_out_payload_0_2_16_imag,
  output     [15:0]   io_coef_out_payload_0_2_17_real,
  output     [15:0]   io_coef_out_payload_0_2_17_imag,
  output     [15:0]   io_coef_out_payload_0_2_18_real,
  output     [15:0]   io_coef_out_payload_0_2_18_imag,
  output     [15:0]   io_coef_out_payload_0_2_19_real,
  output     [15:0]   io_coef_out_payload_0_2_19_imag,
  output     [15:0]   io_coef_out_payload_0_2_20_real,
  output     [15:0]   io_coef_out_payload_0_2_20_imag,
  output     [15:0]   io_coef_out_payload_0_2_21_real,
  output     [15:0]   io_coef_out_payload_0_2_21_imag,
  output     [15:0]   io_coef_out_payload_0_2_22_real,
  output     [15:0]   io_coef_out_payload_0_2_22_imag,
  output     [15:0]   io_coef_out_payload_0_2_23_real,
  output     [15:0]   io_coef_out_payload_0_2_23_imag,
  output     [15:0]   io_coef_out_payload_0_2_24_real,
  output     [15:0]   io_coef_out_payload_0_2_24_imag,
  output     [15:0]   io_coef_out_payload_0_2_25_real,
  output     [15:0]   io_coef_out_payload_0_2_25_imag,
  output     [15:0]   io_coef_out_payload_0_2_26_real,
  output     [15:0]   io_coef_out_payload_0_2_26_imag,
  output     [15:0]   io_coef_out_payload_0_2_27_real,
  output     [15:0]   io_coef_out_payload_0_2_27_imag,
  output     [15:0]   io_coef_out_payload_0_2_28_real,
  output     [15:0]   io_coef_out_payload_0_2_28_imag,
  output     [15:0]   io_coef_out_payload_0_2_29_real,
  output     [15:0]   io_coef_out_payload_0_2_29_imag,
  output     [15:0]   io_coef_out_payload_0_2_30_real,
  output     [15:0]   io_coef_out_payload_0_2_30_imag,
  output     [15:0]   io_coef_out_payload_0_2_31_real,
  output     [15:0]   io_coef_out_payload_0_2_31_imag,
  output     [15:0]   io_coef_out_payload_0_2_32_real,
  output     [15:0]   io_coef_out_payload_0_2_32_imag,
  output     [15:0]   io_coef_out_payload_0_2_33_real,
  output     [15:0]   io_coef_out_payload_0_2_33_imag,
  output     [15:0]   io_coef_out_payload_0_2_34_real,
  output     [15:0]   io_coef_out_payload_0_2_34_imag,
  output     [15:0]   io_coef_out_payload_0_2_35_real,
  output     [15:0]   io_coef_out_payload_0_2_35_imag,
  output     [15:0]   io_coef_out_payload_0_2_36_real,
  output     [15:0]   io_coef_out_payload_0_2_36_imag,
  output     [15:0]   io_coef_out_payload_0_2_37_real,
  output     [15:0]   io_coef_out_payload_0_2_37_imag,
  output     [15:0]   io_coef_out_payload_0_2_38_real,
  output     [15:0]   io_coef_out_payload_0_2_38_imag,
  output     [15:0]   io_coef_out_payload_0_2_39_real,
  output     [15:0]   io_coef_out_payload_0_2_39_imag,
  output     [15:0]   io_coef_out_payload_0_2_40_real,
  output     [15:0]   io_coef_out_payload_0_2_40_imag,
  output     [15:0]   io_coef_out_payload_0_2_41_real,
  output     [15:0]   io_coef_out_payload_0_2_41_imag,
  output     [15:0]   io_coef_out_payload_0_2_42_real,
  output     [15:0]   io_coef_out_payload_0_2_42_imag,
  output     [15:0]   io_coef_out_payload_0_2_43_real,
  output     [15:0]   io_coef_out_payload_0_2_43_imag,
  output     [15:0]   io_coef_out_payload_0_2_44_real,
  output     [15:0]   io_coef_out_payload_0_2_44_imag,
  output     [15:0]   io_coef_out_payload_0_2_45_real,
  output     [15:0]   io_coef_out_payload_0_2_45_imag,
  output     [15:0]   io_coef_out_payload_0_2_46_real,
  output     [15:0]   io_coef_out_payload_0_2_46_imag,
  output     [15:0]   io_coef_out_payload_0_2_47_real,
  output     [15:0]   io_coef_out_payload_0_2_47_imag,
  output     [15:0]   io_coef_out_payload_0_2_48_real,
  output     [15:0]   io_coef_out_payload_0_2_48_imag,
  output     [15:0]   io_coef_out_payload_0_2_49_real,
  output     [15:0]   io_coef_out_payload_0_2_49_imag,
  output     [15:0]   io_coef_out_payload_0_3_0_real,
  output     [15:0]   io_coef_out_payload_0_3_0_imag,
  output     [15:0]   io_coef_out_payload_0_3_1_real,
  output     [15:0]   io_coef_out_payload_0_3_1_imag,
  output     [15:0]   io_coef_out_payload_0_3_2_real,
  output     [15:0]   io_coef_out_payload_0_3_2_imag,
  output     [15:0]   io_coef_out_payload_0_3_3_real,
  output     [15:0]   io_coef_out_payload_0_3_3_imag,
  output     [15:0]   io_coef_out_payload_0_3_4_real,
  output     [15:0]   io_coef_out_payload_0_3_4_imag,
  output     [15:0]   io_coef_out_payload_0_3_5_real,
  output     [15:0]   io_coef_out_payload_0_3_5_imag,
  output     [15:0]   io_coef_out_payload_0_3_6_real,
  output     [15:0]   io_coef_out_payload_0_3_6_imag,
  output     [15:0]   io_coef_out_payload_0_3_7_real,
  output     [15:0]   io_coef_out_payload_0_3_7_imag,
  output     [15:0]   io_coef_out_payload_0_3_8_real,
  output     [15:0]   io_coef_out_payload_0_3_8_imag,
  output     [15:0]   io_coef_out_payload_0_3_9_real,
  output     [15:0]   io_coef_out_payload_0_3_9_imag,
  output     [15:0]   io_coef_out_payload_0_3_10_real,
  output     [15:0]   io_coef_out_payload_0_3_10_imag,
  output     [15:0]   io_coef_out_payload_0_3_11_real,
  output     [15:0]   io_coef_out_payload_0_3_11_imag,
  output     [15:0]   io_coef_out_payload_0_3_12_real,
  output     [15:0]   io_coef_out_payload_0_3_12_imag,
  output     [15:0]   io_coef_out_payload_0_3_13_real,
  output     [15:0]   io_coef_out_payload_0_3_13_imag,
  output     [15:0]   io_coef_out_payload_0_3_14_real,
  output     [15:0]   io_coef_out_payload_0_3_14_imag,
  output     [15:0]   io_coef_out_payload_0_3_15_real,
  output     [15:0]   io_coef_out_payload_0_3_15_imag,
  output     [15:0]   io_coef_out_payload_0_3_16_real,
  output     [15:0]   io_coef_out_payload_0_3_16_imag,
  output     [15:0]   io_coef_out_payload_0_3_17_real,
  output     [15:0]   io_coef_out_payload_0_3_17_imag,
  output     [15:0]   io_coef_out_payload_0_3_18_real,
  output     [15:0]   io_coef_out_payload_0_3_18_imag,
  output     [15:0]   io_coef_out_payload_0_3_19_real,
  output     [15:0]   io_coef_out_payload_0_3_19_imag,
  output     [15:0]   io_coef_out_payload_0_3_20_real,
  output     [15:0]   io_coef_out_payload_0_3_20_imag,
  output     [15:0]   io_coef_out_payload_0_3_21_real,
  output     [15:0]   io_coef_out_payload_0_3_21_imag,
  output     [15:0]   io_coef_out_payload_0_3_22_real,
  output     [15:0]   io_coef_out_payload_0_3_22_imag,
  output     [15:0]   io_coef_out_payload_0_3_23_real,
  output     [15:0]   io_coef_out_payload_0_3_23_imag,
  output     [15:0]   io_coef_out_payload_0_3_24_real,
  output     [15:0]   io_coef_out_payload_0_3_24_imag,
  output     [15:0]   io_coef_out_payload_0_3_25_real,
  output     [15:0]   io_coef_out_payload_0_3_25_imag,
  output     [15:0]   io_coef_out_payload_0_3_26_real,
  output     [15:0]   io_coef_out_payload_0_3_26_imag,
  output     [15:0]   io_coef_out_payload_0_3_27_real,
  output     [15:0]   io_coef_out_payload_0_3_27_imag,
  output     [15:0]   io_coef_out_payload_0_3_28_real,
  output     [15:0]   io_coef_out_payload_0_3_28_imag,
  output     [15:0]   io_coef_out_payload_0_3_29_real,
  output     [15:0]   io_coef_out_payload_0_3_29_imag,
  output     [15:0]   io_coef_out_payload_0_3_30_real,
  output     [15:0]   io_coef_out_payload_0_3_30_imag,
  output     [15:0]   io_coef_out_payload_0_3_31_real,
  output     [15:0]   io_coef_out_payload_0_3_31_imag,
  output     [15:0]   io_coef_out_payload_0_3_32_real,
  output     [15:0]   io_coef_out_payload_0_3_32_imag,
  output     [15:0]   io_coef_out_payload_0_3_33_real,
  output     [15:0]   io_coef_out_payload_0_3_33_imag,
  output     [15:0]   io_coef_out_payload_0_3_34_real,
  output     [15:0]   io_coef_out_payload_0_3_34_imag,
  output     [15:0]   io_coef_out_payload_0_3_35_real,
  output     [15:0]   io_coef_out_payload_0_3_35_imag,
  output     [15:0]   io_coef_out_payload_0_3_36_real,
  output     [15:0]   io_coef_out_payload_0_3_36_imag,
  output     [15:0]   io_coef_out_payload_0_3_37_real,
  output     [15:0]   io_coef_out_payload_0_3_37_imag,
  output     [15:0]   io_coef_out_payload_0_3_38_real,
  output     [15:0]   io_coef_out_payload_0_3_38_imag,
  output     [15:0]   io_coef_out_payload_0_3_39_real,
  output     [15:0]   io_coef_out_payload_0_3_39_imag,
  output     [15:0]   io_coef_out_payload_0_3_40_real,
  output     [15:0]   io_coef_out_payload_0_3_40_imag,
  output     [15:0]   io_coef_out_payload_0_3_41_real,
  output     [15:0]   io_coef_out_payload_0_3_41_imag,
  output     [15:0]   io_coef_out_payload_0_3_42_real,
  output     [15:0]   io_coef_out_payload_0_3_42_imag,
  output     [15:0]   io_coef_out_payload_0_3_43_real,
  output     [15:0]   io_coef_out_payload_0_3_43_imag,
  output     [15:0]   io_coef_out_payload_0_3_44_real,
  output     [15:0]   io_coef_out_payload_0_3_44_imag,
  output     [15:0]   io_coef_out_payload_0_3_45_real,
  output     [15:0]   io_coef_out_payload_0_3_45_imag,
  output     [15:0]   io_coef_out_payload_0_3_46_real,
  output     [15:0]   io_coef_out_payload_0_3_46_imag,
  output     [15:0]   io_coef_out_payload_0_3_47_real,
  output     [15:0]   io_coef_out_payload_0_3_47_imag,
  output     [15:0]   io_coef_out_payload_0_3_48_real,
  output     [15:0]   io_coef_out_payload_0_3_48_imag,
  output     [15:0]   io_coef_out_payload_0_3_49_real,
  output     [15:0]   io_coef_out_payload_0_3_49_imag,
  output     [15:0]   io_coef_out_payload_0_4_0_real,
  output     [15:0]   io_coef_out_payload_0_4_0_imag,
  output     [15:0]   io_coef_out_payload_0_4_1_real,
  output     [15:0]   io_coef_out_payload_0_4_1_imag,
  output     [15:0]   io_coef_out_payload_0_4_2_real,
  output     [15:0]   io_coef_out_payload_0_4_2_imag,
  output     [15:0]   io_coef_out_payload_0_4_3_real,
  output     [15:0]   io_coef_out_payload_0_4_3_imag,
  output     [15:0]   io_coef_out_payload_0_4_4_real,
  output     [15:0]   io_coef_out_payload_0_4_4_imag,
  output     [15:0]   io_coef_out_payload_0_4_5_real,
  output     [15:0]   io_coef_out_payload_0_4_5_imag,
  output     [15:0]   io_coef_out_payload_0_4_6_real,
  output     [15:0]   io_coef_out_payload_0_4_6_imag,
  output     [15:0]   io_coef_out_payload_0_4_7_real,
  output     [15:0]   io_coef_out_payload_0_4_7_imag,
  output     [15:0]   io_coef_out_payload_0_4_8_real,
  output     [15:0]   io_coef_out_payload_0_4_8_imag,
  output     [15:0]   io_coef_out_payload_0_4_9_real,
  output     [15:0]   io_coef_out_payload_0_4_9_imag,
  output     [15:0]   io_coef_out_payload_0_4_10_real,
  output     [15:0]   io_coef_out_payload_0_4_10_imag,
  output     [15:0]   io_coef_out_payload_0_4_11_real,
  output     [15:0]   io_coef_out_payload_0_4_11_imag,
  output     [15:0]   io_coef_out_payload_0_4_12_real,
  output     [15:0]   io_coef_out_payload_0_4_12_imag,
  output     [15:0]   io_coef_out_payload_0_4_13_real,
  output     [15:0]   io_coef_out_payload_0_4_13_imag,
  output     [15:0]   io_coef_out_payload_0_4_14_real,
  output     [15:0]   io_coef_out_payload_0_4_14_imag,
  output     [15:0]   io_coef_out_payload_0_4_15_real,
  output     [15:0]   io_coef_out_payload_0_4_15_imag,
  output     [15:0]   io_coef_out_payload_0_4_16_real,
  output     [15:0]   io_coef_out_payload_0_4_16_imag,
  output     [15:0]   io_coef_out_payload_0_4_17_real,
  output     [15:0]   io_coef_out_payload_0_4_17_imag,
  output     [15:0]   io_coef_out_payload_0_4_18_real,
  output     [15:0]   io_coef_out_payload_0_4_18_imag,
  output     [15:0]   io_coef_out_payload_0_4_19_real,
  output     [15:0]   io_coef_out_payload_0_4_19_imag,
  output     [15:0]   io_coef_out_payload_0_4_20_real,
  output     [15:0]   io_coef_out_payload_0_4_20_imag,
  output     [15:0]   io_coef_out_payload_0_4_21_real,
  output     [15:0]   io_coef_out_payload_0_4_21_imag,
  output     [15:0]   io_coef_out_payload_0_4_22_real,
  output     [15:0]   io_coef_out_payload_0_4_22_imag,
  output     [15:0]   io_coef_out_payload_0_4_23_real,
  output     [15:0]   io_coef_out_payload_0_4_23_imag,
  output     [15:0]   io_coef_out_payload_0_4_24_real,
  output     [15:0]   io_coef_out_payload_0_4_24_imag,
  output     [15:0]   io_coef_out_payload_0_4_25_real,
  output     [15:0]   io_coef_out_payload_0_4_25_imag,
  output     [15:0]   io_coef_out_payload_0_4_26_real,
  output     [15:0]   io_coef_out_payload_0_4_26_imag,
  output     [15:0]   io_coef_out_payload_0_4_27_real,
  output     [15:0]   io_coef_out_payload_0_4_27_imag,
  output     [15:0]   io_coef_out_payload_0_4_28_real,
  output     [15:0]   io_coef_out_payload_0_4_28_imag,
  output     [15:0]   io_coef_out_payload_0_4_29_real,
  output     [15:0]   io_coef_out_payload_0_4_29_imag,
  output     [15:0]   io_coef_out_payload_0_4_30_real,
  output     [15:0]   io_coef_out_payload_0_4_30_imag,
  output     [15:0]   io_coef_out_payload_0_4_31_real,
  output     [15:0]   io_coef_out_payload_0_4_31_imag,
  output     [15:0]   io_coef_out_payload_0_4_32_real,
  output     [15:0]   io_coef_out_payload_0_4_32_imag,
  output     [15:0]   io_coef_out_payload_0_4_33_real,
  output     [15:0]   io_coef_out_payload_0_4_33_imag,
  output     [15:0]   io_coef_out_payload_0_4_34_real,
  output     [15:0]   io_coef_out_payload_0_4_34_imag,
  output     [15:0]   io_coef_out_payload_0_4_35_real,
  output     [15:0]   io_coef_out_payload_0_4_35_imag,
  output     [15:0]   io_coef_out_payload_0_4_36_real,
  output     [15:0]   io_coef_out_payload_0_4_36_imag,
  output     [15:0]   io_coef_out_payload_0_4_37_real,
  output     [15:0]   io_coef_out_payload_0_4_37_imag,
  output     [15:0]   io_coef_out_payload_0_4_38_real,
  output     [15:0]   io_coef_out_payload_0_4_38_imag,
  output     [15:0]   io_coef_out_payload_0_4_39_real,
  output     [15:0]   io_coef_out_payload_0_4_39_imag,
  output     [15:0]   io_coef_out_payload_0_4_40_real,
  output     [15:0]   io_coef_out_payload_0_4_40_imag,
  output     [15:0]   io_coef_out_payload_0_4_41_real,
  output     [15:0]   io_coef_out_payload_0_4_41_imag,
  output     [15:0]   io_coef_out_payload_0_4_42_real,
  output     [15:0]   io_coef_out_payload_0_4_42_imag,
  output     [15:0]   io_coef_out_payload_0_4_43_real,
  output     [15:0]   io_coef_out_payload_0_4_43_imag,
  output     [15:0]   io_coef_out_payload_0_4_44_real,
  output     [15:0]   io_coef_out_payload_0_4_44_imag,
  output     [15:0]   io_coef_out_payload_0_4_45_real,
  output     [15:0]   io_coef_out_payload_0_4_45_imag,
  output     [15:0]   io_coef_out_payload_0_4_46_real,
  output     [15:0]   io_coef_out_payload_0_4_46_imag,
  output     [15:0]   io_coef_out_payload_0_4_47_real,
  output     [15:0]   io_coef_out_payload_0_4_47_imag,
  output     [15:0]   io_coef_out_payload_0_4_48_real,
  output     [15:0]   io_coef_out_payload_0_4_48_imag,
  output     [15:0]   io_coef_out_payload_0_4_49_real,
  output     [15:0]   io_coef_out_payload_0_4_49_imag,
  output     [15:0]   io_coef_out_payload_0_5_0_real,
  output     [15:0]   io_coef_out_payload_0_5_0_imag,
  output     [15:0]   io_coef_out_payload_0_5_1_real,
  output     [15:0]   io_coef_out_payload_0_5_1_imag,
  output     [15:0]   io_coef_out_payload_0_5_2_real,
  output     [15:0]   io_coef_out_payload_0_5_2_imag,
  output     [15:0]   io_coef_out_payload_0_5_3_real,
  output     [15:0]   io_coef_out_payload_0_5_3_imag,
  output     [15:0]   io_coef_out_payload_0_5_4_real,
  output     [15:0]   io_coef_out_payload_0_5_4_imag,
  output     [15:0]   io_coef_out_payload_0_5_5_real,
  output     [15:0]   io_coef_out_payload_0_5_5_imag,
  output     [15:0]   io_coef_out_payload_0_5_6_real,
  output     [15:0]   io_coef_out_payload_0_5_6_imag,
  output     [15:0]   io_coef_out_payload_0_5_7_real,
  output     [15:0]   io_coef_out_payload_0_5_7_imag,
  output     [15:0]   io_coef_out_payload_0_5_8_real,
  output     [15:0]   io_coef_out_payload_0_5_8_imag,
  output     [15:0]   io_coef_out_payload_0_5_9_real,
  output     [15:0]   io_coef_out_payload_0_5_9_imag,
  output     [15:0]   io_coef_out_payload_0_5_10_real,
  output     [15:0]   io_coef_out_payload_0_5_10_imag,
  output     [15:0]   io_coef_out_payload_0_5_11_real,
  output     [15:0]   io_coef_out_payload_0_5_11_imag,
  output     [15:0]   io_coef_out_payload_0_5_12_real,
  output     [15:0]   io_coef_out_payload_0_5_12_imag,
  output     [15:0]   io_coef_out_payload_0_5_13_real,
  output     [15:0]   io_coef_out_payload_0_5_13_imag,
  output     [15:0]   io_coef_out_payload_0_5_14_real,
  output     [15:0]   io_coef_out_payload_0_5_14_imag,
  output     [15:0]   io_coef_out_payload_0_5_15_real,
  output     [15:0]   io_coef_out_payload_0_5_15_imag,
  output     [15:0]   io_coef_out_payload_0_5_16_real,
  output     [15:0]   io_coef_out_payload_0_5_16_imag,
  output     [15:0]   io_coef_out_payload_0_5_17_real,
  output     [15:0]   io_coef_out_payload_0_5_17_imag,
  output     [15:0]   io_coef_out_payload_0_5_18_real,
  output     [15:0]   io_coef_out_payload_0_5_18_imag,
  output     [15:0]   io_coef_out_payload_0_5_19_real,
  output     [15:0]   io_coef_out_payload_0_5_19_imag,
  output     [15:0]   io_coef_out_payload_0_5_20_real,
  output     [15:0]   io_coef_out_payload_0_5_20_imag,
  output     [15:0]   io_coef_out_payload_0_5_21_real,
  output     [15:0]   io_coef_out_payload_0_5_21_imag,
  output     [15:0]   io_coef_out_payload_0_5_22_real,
  output     [15:0]   io_coef_out_payload_0_5_22_imag,
  output     [15:0]   io_coef_out_payload_0_5_23_real,
  output     [15:0]   io_coef_out_payload_0_5_23_imag,
  output     [15:0]   io_coef_out_payload_0_5_24_real,
  output     [15:0]   io_coef_out_payload_0_5_24_imag,
  output     [15:0]   io_coef_out_payload_0_5_25_real,
  output     [15:0]   io_coef_out_payload_0_5_25_imag,
  output     [15:0]   io_coef_out_payload_0_5_26_real,
  output     [15:0]   io_coef_out_payload_0_5_26_imag,
  output     [15:0]   io_coef_out_payload_0_5_27_real,
  output     [15:0]   io_coef_out_payload_0_5_27_imag,
  output     [15:0]   io_coef_out_payload_0_5_28_real,
  output     [15:0]   io_coef_out_payload_0_5_28_imag,
  output     [15:0]   io_coef_out_payload_0_5_29_real,
  output     [15:0]   io_coef_out_payload_0_5_29_imag,
  output     [15:0]   io_coef_out_payload_0_5_30_real,
  output     [15:0]   io_coef_out_payload_0_5_30_imag,
  output     [15:0]   io_coef_out_payload_0_5_31_real,
  output     [15:0]   io_coef_out_payload_0_5_31_imag,
  output     [15:0]   io_coef_out_payload_0_5_32_real,
  output     [15:0]   io_coef_out_payload_0_5_32_imag,
  output     [15:0]   io_coef_out_payload_0_5_33_real,
  output     [15:0]   io_coef_out_payload_0_5_33_imag,
  output     [15:0]   io_coef_out_payload_0_5_34_real,
  output     [15:0]   io_coef_out_payload_0_5_34_imag,
  output     [15:0]   io_coef_out_payload_0_5_35_real,
  output     [15:0]   io_coef_out_payload_0_5_35_imag,
  output     [15:0]   io_coef_out_payload_0_5_36_real,
  output     [15:0]   io_coef_out_payload_0_5_36_imag,
  output     [15:0]   io_coef_out_payload_0_5_37_real,
  output     [15:0]   io_coef_out_payload_0_5_37_imag,
  output     [15:0]   io_coef_out_payload_0_5_38_real,
  output     [15:0]   io_coef_out_payload_0_5_38_imag,
  output     [15:0]   io_coef_out_payload_0_5_39_real,
  output     [15:0]   io_coef_out_payload_0_5_39_imag,
  output     [15:0]   io_coef_out_payload_0_5_40_real,
  output     [15:0]   io_coef_out_payload_0_5_40_imag,
  output     [15:0]   io_coef_out_payload_0_5_41_real,
  output     [15:0]   io_coef_out_payload_0_5_41_imag,
  output     [15:0]   io_coef_out_payload_0_5_42_real,
  output     [15:0]   io_coef_out_payload_0_5_42_imag,
  output     [15:0]   io_coef_out_payload_0_5_43_real,
  output     [15:0]   io_coef_out_payload_0_5_43_imag,
  output     [15:0]   io_coef_out_payload_0_5_44_real,
  output     [15:0]   io_coef_out_payload_0_5_44_imag,
  output     [15:0]   io_coef_out_payload_0_5_45_real,
  output     [15:0]   io_coef_out_payload_0_5_45_imag,
  output     [15:0]   io_coef_out_payload_0_5_46_real,
  output     [15:0]   io_coef_out_payload_0_5_46_imag,
  output     [15:0]   io_coef_out_payload_0_5_47_real,
  output     [15:0]   io_coef_out_payload_0_5_47_imag,
  output     [15:0]   io_coef_out_payload_0_5_48_real,
  output     [15:0]   io_coef_out_payload_0_5_48_imag,
  output     [15:0]   io_coef_out_payload_0_5_49_real,
  output     [15:0]   io_coef_out_payload_0_5_49_imag,
  output     [15:0]   io_coef_out_payload_0_6_0_real,
  output     [15:0]   io_coef_out_payload_0_6_0_imag,
  output     [15:0]   io_coef_out_payload_0_6_1_real,
  output     [15:0]   io_coef_out_payload_0_6_1_imag,
  output     [15:0]   io_coef_out_payload_0_6_2_real,
  output     [15:0]   io_coef_out_payload_0_6_2_imag,
  output     [15:0]   io_coef_out_payload_0_6_3_real,
  output     [15:0]   io_coef_out_payload_0_6_3_imag,
  output     [15:0]   io_coef_out_payload_0_6_4_real,
  output     [15:0]   io_coef_out_payload_0_6_4_imag,
  output     [15:0]   io_coef_out_payload_0_6_5_real,
  output     [15:0]   io_coef_out_payload_0_6_5_imag,
  output     [15:0]   io_coef_out_payload_0_6_6_real,
  output     [15:0]   io_coef_out_payload_0_6_6_imag,
  output     [15:0]   io_coef_out_payload_0_6_7_real,
  output     [15:0]   io_coef_out_payload_0_6_7_imag,
  output     [15:0]   io_coef_out_payload_0_6_8_real,
  output     [15:0]   io_coef_out_payload_0_6_8_imag,
  output     [15:0]   io_coef_out_payload_0_6_9_real,
  output     [15:0]   io_coef_out_payload_0_6_9_imag,
  output     [15:0]   io_coef_out_payload_0_6_10_real,
  output     [15:0]   io_coef_out_payload_0_6_10_imag,
  output     [15:0]   io_coef_out_payload_0_6_11_real,
  output     [15:0]   io_coef_out_payload_0_6_11_imag,
  output     [15:0]   io_coef_out_payload_0_6_12_real,
  output     [15:0]   io_coef_out_payload_0_6_12_imag,
  output     [15:0]   io_coef_out_payload_0_6_13_real,
  output     [15:0]   io_coef_out_payload_0_6_13_imag,
  output     [15:0]   io_coef_out_payload_0_6_14_real,
  output     [15:0]   io_coef_out_payload_0_6_14_imag,
  output     [15:0]   io_coef_out_payload_0_6_15_real,
  output     [15:0]   io_coef_out_payload_0_6_15_imag,
  output     [15:0]   io_coef_out_payload_0_6_16_real,
  output     [15:0]   io_coef_out_payload_0_6_16_imag,
  output     [15:0]   io_coef_out_payload_0_6_17_real,
  output     [15:0]   io_coef_out_payload_0_6_17_imag,
  output     [15:0]   io_coef_out_payload_0_6_18_real,
  output     [15:0]   io_coef_out_payload_0_6_18_imag,
  output     [15:0]   io_coef_out_payload_0_6_19_real,
  output     [15:0]   io_coef_out_payload_0_6_19_imag,
  output     [15:0]   io_coef_out_payload_0_6_20_real,
  output     [15:0]   io_coef_out_payload_0_6_20_imag,
  output     [15:0]   io_coef_out_payload_0_6_21_real,
  output     [15:0]   io_coef_out_payload_0_6_21_imag,
  output     [15:0]   io_coef_out_payload_0_6_22_real,
  output     [15:0]   io_coef_out_payload_0_6_22_imag,
  output     [15:0]   io_coef_out_payload_0_6_23_real,
  output     [15:0]   io_coef_out_payload_0_6_23_imag,
  output     [15:0]   io_coef_out_payload_0_6_24_real,
  output     [15:0]   io_coef_out_payload_0_6_24_imag,
  output     [15:0]   io_coef_out_payload_0_6_25_real,
  output     [15:0]   io_coef_out_payload_0_6_25_imag,
  output     [15:0]   io_coef_out_payload_0_6_26_real,
  output     [15:0]   io_coef_out_payload_0_6_26_imag,
  output     [15:0]   io_coef_out_payload_0_6_27_real,
  output     [15:0]   io_coef_out_payload_0_6_27_imag,
  output     [15:0]   io_coef_out_payload_0_6_28_real,
  output     [15:0]   io_coef_out_payload_0_6_28_imag,
  output     [15:0]   io_coef_out_payload_0_6_29_real,
  output     [15:0]   io_coef_out_payload_0_6_29_imag,
  output     [15:0]   io_coef_out_payload_0_6_30_real,
  output     [15:0]   io_coef_out_payload_0_6_30_imag,
  output     [15:0]   io_coef_out_payload_0_6_31_real,
  output     [15:0]   io_coef_out_payload_0_6_31_imag,
  output     [15:0]   io_coef_out_payload_0_6_32_real,
  output     [15:0]   io_coef_out_payload_0_6_32_imag,
  output     [15:0]   io_coef_out_payload_0_6_33_real,
  output     [15:0]   io_coef_out_payload_0_6_33_imag,
  output     [15:0]   io_coef_out_payload_0_6_34_real,
  output     [15:0]   io_coef_out_payload_0_6_34_imag,
  output     [15:0]   io_coef_out_payload_0_6_35_real,
  output     [15:0]   io_coef_out_payload_0_6_35_imag,
  output     [15:0]   io_coef_out_payload_0_6_36_real,
  output     [15:0]   io_coef_out_payload_0_6_36_imag,
  output     [15:0]   io_coef_out_payload_0_6_37_real,
  output     [15:0]   io_coef_out_payload_0_6_37_imag,
  output     [15:0]   io_coef_out_payload_0_6_38_real,
  output     [15:0]   io_coef_out_payload_0_6_38_imag,
  output     [15:0]   io_coef_out_payload_0_6_39_real,
  output     [15:0]   io_coef_out_payload_0_6_39_imag,
  output     [15:0]   io_coef_out_payload_0_6_40_real,
  output     [15:0]   io_coef_out_payload_0_6_40_imag,
  output     [15:0]   io_coef_out_payload_0_6_41_real,
  output     [15:0]   io_coef_out_payload_0_6_41_imag,
  output     [15:0]   io_coef_out_payload_0_6_42_real,
  output     [15:0]   io_coef_out_payload_0_6_42_imag,
  output     [15:0]   io_coef_out_payload_0_6_43_real,
  output     [15:0]   io_coef_out_payload_0_6_43_imag,
  output     [15:0]   io_coef_out_payload_0_6_44_real,
  output     [15:0]   io_coef_out_payload_0_6_44_imag,
  output     [15:0]   io_coef_out_payload_0_6_45_real,
  output     [15:0]   io_coef_out_payload_0_6_45_imag,
  output     [15:0]   io_coef_out_payload_0_6_46_real,
  output     [15:0]   io_coef_out_payload_0_6_46_imag,
  output     [15:0]   io_coef_out_payload_0_6_47_real,
  output     [15:0]   io_coef_out_payload_0_6_47_imag,
  output     [15:0]   io_coef_out_payload_0_6_48_real,
  output     [15:0]   io_coef_out_payload_0_6_48_imag,
  output     [15:0]   io_coef_out_payload_0_6_49_real,
  output     [15:0]   io_coef_out_payload_0_6_49_imag,
  output     [15:0]   io_coef_out_payload_0_7_0_real,
  output     [15:0]   io_coef_out_payload_0_7_0_imag,
  output     [15:0]   io_coef_out_payload_0_7_1_real,
  output     [15:0]   io_coef_out_payload_0_7_1_imag,
  output     [15:0]   io_coef_out_payload_0_7_2_real,
  output     [15:0]   io_coef_out_payload_0_7_2_imag,
  output     [15:0]   io_coef_out_payload_0_7_3_real,
  output     [15:0]   io_coef_out_payload_0_7_3_imag,
  output     [15:0]   io_coef_out_payload_0_7_4_real,
  output     [15:0]   io_coef_out_payload_0_7_4_imag,
  output     [15:0]   io_coef_out_payload_0_7_5_real,
  output     [15:0]   io_coef_out_payload_0_7_5_imag,
  output     [15:0]   io_coef_out_payload_0_7_6_real,
  output     [15:0]   io_coef_out_payload_0_7_6_imag,
  output     [15:0]   io_coef_out_payload_0_7_7_real,
  output     [15:0]   io_coef_out_payload_0_7_7_imag,
  output     [15:0]   io_coef_out_payload_0_7_8_real,
  output     [15:0]   io_coef_out_payload_0_7_8_imag,
  output     [15:0]   io_coef_out_payload_0_7_9_real,
  output     [15:0]   io_coef_out_payload_0_7_9_imag,
  output     [15:0]   io_coef_out_payload_0_7_10_real,
  output     [15:0]   io_coef_out_payload_0_7_10_imag,
  output     [15:0]   io_coef_out_payload_0_7_11_real,
  output     [15:0]   io_coef_out_payload_0_7_11_imag,
  output     [15:0]   io_coef_out_payload_0_7_12_real,
  output     [15:0]   io_coef_out_payload_0_7_12_imag,
  output     [15:0]   io_coef_out_payload_0_7_13_real,
  output     [15:0]   io_coef_out_payload_0_7_13_imag,
  output     [15:0]   io_coef_out_payload_0_7_14_real,
  output     [15:0]   io_coef_out_payload_0_7_14_imag,
  output     [15:0]   io_coef_out_payload_0_7_15_real,
  output     [15:0]   io_coef_out_payload_0_7_15_imag,
  output     [15:0]   io_coef_out_payload_0_7_16_real,
  output     [15:0]   io_coef_out_payload_0_7_16_imag,
  output     [15:0]   io_coef_out_payload_0_7_17_real,
  output     [15:0]   io_coef_out_payload_0_7_17_imag,
  output     [15:0]   io_coef_out_payload_0_7_18_real,
  output     [15:0]   io_coef_out_payload_0_7_18_imag,
  output     [15:0]   io_coef_out_payload_0_7_19_real,
  output     [15:0]   io_coef_out_payload_0_7_19_imag,
  output     [15:0]   io_coef_out_payload_0_7_20_real,
  output     [15:0]   io_coef_out_payload_0_7_20_imag,
  output     [15:0]   io_coef_out_payload_0_7_21_real,
  output     [15:0]   io_coef_out_payload_0_7_21_imag,
  output     [15:0]   io_coef_out_payload_0_7_22_real,
  output     [15:0]   io_coef_out_payload_0_7_22_imag,
  output     [15:0]   io_coef_out_payload_0_7_23_real,
  output     [15:0]   io_coef_out_payload_0_7_23_imag,
  output     [15:0]   io_coef_out_payload_0_7_24_real,
  output     [15:0]   io_coef_out_payload_0_7_24_imag,
  output     [15:0]   io_coef_out_payload_0_7_25_real,
  output     [15:0]   io_coef_out_payload_0_7_25_imag,
  output     [15:0]   io_coef_out_payload_0_7_26_real,
  output     [15:0]   io_coef_out_payload_0_7_26_imag,
  output     [15:0]   io_coef_out_payload_0_7_27_real,
  output     [15:0]   io_coef_out_payload_0_7_27_imag,
  output     [15:0]   io_coef_out_payload_0_7_28_real,
  output     [15:0]   io_coef_out_payload_0_7_28_imag,
  output     [15:0]   io_coef_out_payload_0_7_29_real,
  output     [15:0]   io_coef_out_payload_0_7_29_imag,
  output     [15:0]   io_coef_out_payload_0_7_30_real,
  output     [15:0]   io_coef_out_payload_0_7_30_imag,
  output     [15:0]   io_coef_out_payload_0_7_31_real,
  output     [15:0]   io_coef_out_payload_0_7_31_imag,
  output     [15:0]   io_coef_out_payload_0_7_32_real,
  output     [15:0]   io_coef_out_payload_0_7_32_imag,
  output     [15:0]   io_coef_out_payload_0_7_33_real,
  output     [15:0]   io_coef_out_payload_0_7_33_imag,
  output     [15:0]   io_coef_out_payload_0_7_34_real,
  output     [15:0]   io_coef_out_payload_0_7_34_imag,
  output     [15:0]   io_coef_out_payload_0_7_35_real,
  output     [15:0]   io_coef_out_payload_0_7_35_imag,
  output     [15:0]   io_coef_out_payload_0_7_36_real,
  output     [15:0]   io_coef_out_payload_0_7_36_imag,
  output     [15:0]   io_coef_out_payload_0_7_37_real,
  output     [15:0]   io_coef_out_payload_0_7_37_imag,
  output     [15:0]   io_coef_out_payload_0_7_38_real,
  output     [15:0]   io_coef_out_payload_0_7_38_imag,
  output     [15:0]   io_coef_out_payload_0_7_39_real,
  output     [15:0]   io_coef_out_payload_0_7_39_imag,
  output     [15:0]   io_coef_out_payload_0_7_40_real,
  output     [15:0]   io_coef_out_payload_0_7_40_imag,
  output     [15:0]   io_coef_out_payload_0_7_41_real,
  output     [15:0]   io_coef_out_payload_0_7_41_imag,
  output     [15:0]   io_coef_out_payload_0_7_42_real,
  output     [15:0]   io_coef_out_payload_0_7_42_imag,
  output     [15:0]   io_coef_out_payload_0_7_43_real,
  output     [15:0]   io_coef_out_payload_0_7_43_imag,
  output     [15:0]   io_coef_out_payload_0_7_44_real,
  output     [15:0]   io_coef_out_payload_0_7_44_imag,
  output     [15:0]   io_coef_out_payload_0_7_45_real,
  output     [15:0]   io_coef_out_payload_0_7_45_imag,
  output     [15:0]   io_coef_out_payload_0_7_46_real,
  output     [15:0]   io_coef_out_payload_0_7_46_imag,
  output     [15:0]   io_coef_out_payload_0_7_47_real,
  output     [15:0]   io_coef_out_payload_0_7_47_imag,
  output     [15:0]   io_coef_out_payload_0_7_48_real,
  output     [15:0]   io_coef_out_payload_0_7_48_imag,
  output     [15:0]   io_coef_out_payload_0_7_49_real,
  output     [15:0]   io_coef_out_payload_0_7_49_imag,
  output     [15:0]   io_coef_out_payload_0_8_0_real,
  output     [15:0]   io_coef_out_payload_0_8_0_imag,
  output     [15:0]   io_coef_out_payload_0_8_1_real,
  output     [15:0]   io_coef_out_payload_0_8_1_imag,
  output     [15:0]   io_coef_out_payload_0_8_2_real,
  output     [15:0]   io_coef_out_payload_0_8_2_imag,
  output     [15:0]   io_coef_out_payload_0_8_3_real,
  output     [15:0]   io_coef_out_payload_0_8_3_imag,
  output     [15:0]   io_coef_out_payload_0_8_4_real,
  output     [15:0]   io_coef_out_payload_0_8_4_imag,
  output     [15:0]   io_coef_out_payload_0_8_5_real,
  output     [15:0]   io_coef_out_payload_0_8_5_imag,
  output     [15:0]   io_coef_out_payload_0_8_6_real,
  output     [15:0]   io_coef_out_payload_0_8_6_imag,
  output     [15:0]   io_coef_out_payload_0_8_7_real,
  output     [15:0]   io_coef_out_payload_0_8_7_imag,
  output     [15:0]   io_coef_out_payload_0_8_8_real,
  output     [15:0]   io_coef_out_payload_0_8_8_imag,
  output     [15:0]   io_coef_out_payload_0_8_9_real,
  output     [15:0]   io_coef_out_payload_0_8_9_imag,
  output     [15:0]   io_coef_out_payload_0_8_10_real,
  output     [15:0]   io_coef_out_payload_0_8_10_imag,
  output     [15:0]   io_coef_out_payload_0_8_11_real,
  output     [15:0]   io_coef_out_payload_0_8_11_imag,
  output     [15:0]   io_coef_out_payload_0_8_12_real,
  output     [15:0]   io_coef_out_payload_0_8_12_imag,
  output     [15:0]   io_coef_out_payload_0_8_13_real,
  output     [15:0]   io_coef_out_payload_0_8_13_imag,
  output     [15:0]   io_coef_out_payload_0_8_14_real,
  output     [15:0]   io_coef_out_payload_0_8_14_imag,
  output     [15:0]   io_coef_out_payload_0_8_15_real,
  output     [15:0]   io_coef_out_payload_0_8_15_imag,
  output     [15:0]   io_coef_out_payload_0_8_16_real,
  output     [15:0]   io_coef_out_payload_0_8_16_imag,
  output     [15:0]   io_coef_out_payload_0_8_17_real,
  output     [15:0]   io_coef_out_payload_0_8_17_imag,
  output     [15:0]   io_coef_out_payload_0_8_18_real,
  output     [15:0]   io_coef_out_payload_0_8_18_imag,
  output     [15:0]   io_coef_out_payload_0_8_19_real,
  output     [15:0]   io_coef_out_payload_0_8_19_imag,
  output     [15:0]   io_coef_out_payload_0_8_20_real,
  output     [15:0]   io_coef_out_payload_0_8_20_imag,
  output     [15:0]   io_coef_out_payload_0_8_21_real,
  output     [15:0]   io_coef_out_payload_0_8_21_imag,
  output     [15:0]   io_coef_out_payload_0_8_22_real,
  output     [15:0]   io_coef_out_payload_0_8_22_imag,
  output     [15:0]   io_coef_out_payload_0_8_23_real,
  output     [15:0]   io_coef_out_payload_0_8_23_imag,
  output     [15:0]   io_coef_out_payload_0_8_24_real,
  output     [15:0]   io_coef_out_payload_0_8_24_imag,
  output     [15:0]   io_coef_out_payload_0_8_25_real,
  output     [15:0]   io_coef_out_payload_0_8_25_imag,
  output     [15:0]   io_coef_out_payload_0_8_26_real,
  output     [15:0]   io_coef_out_payload_0_8_26_imag,
  output     [15:0]   io_coef_out_payload_0_8_27_real,
  output     [15:0]   io_coef_out_payload_0_8_27_imag,
  output     [15:0]   io_coef_out_payload_0_8_28_real,
  output     [15:0]   io_coef_out_payload_0_8_28_imag,
  output     [15:0]   io_coef_out_payload_0_8_29_real,
  output     [15:0]   io_coef_out_payload_0_8_29_imag,
  output     [15:0]   io_coef_out_payload_0_8_30_real,
  output     [15:0]   io_coef_out_payload_0_8_30_imag,
  output     [15:0]   io_coef_out_payload_0_8_31_real,
  output     [15:0]   io_coef_out_payload_0_8_31_imag,
  output     [15:0]   io_coef_out_payload_0_8_32_real,
  output     [15:0]   io_coef_out_payload_0_8_32_imag,
  output     [15:0]   io_coef_out_payload_0_8_33_real,
  output     [15:0]   io_coef_out_payload_0_8_33_imag,
  output     [15:0]   io_coef_out_payload_0_8_34_real,
  output     [15:0]   io_coef_out_payload_0_8_34_imag,
  output     [15:0]   io_coef_out_payload_0_8_35_real,
  output     [15:0]   io_coef_out_payload_0_8_35_imag,
  output     [15:0]   io_coef_out_payload_0_8_36_real,
  output     [15:0]   io_coef_out_payload_0_8_36_imag,
  output     [15:0]   io_coef_out_payload_0_8_37_real,
  output     [15:0]   io_coef_out_payload_0_8_37_imag,
  output     [15:0]   io_coef_out_payload_0_8_38_real,
  output     [15:0]   io_coef_out_payload_0_8_38_imag,
  output     [15:0]   io_coef_out_payload_0_8_39_real,
  output     [15:0]   io_coef_out_payload_0_8_39_imag,
  output     [15:0]   io_coef_out_payload_0_8_40_real,
  output     [15:0]   io_coef_out_payload_0_8_40_imag,
  output     [15:0]   io_coef_out_payload_0_8_41_real,
  output     [15:0]   io_coef_out_payload_0_8_41_imag,
  output     [15:0]   io_coef_out_payload_0_8_42_real,
  output     [15:0]   io_coef_out_payload_0_8_42_imag,
  output     [15:0]   io_coef_out_payload_0_8_43_real,
  output     [15:0]   io_coef_out_payload_0_8_43_imag,
  output     [15:0]   io_coef_out_payload_0_8_44_real,
  output     [15:0]   io_coef_out_payload_0_8_44_imag,
  output     [15:0]   io_coef_out_payload_0_8_45_real,
  output     [15:0]   io_coef_out_payload_0_8_45_imag,
  output     [15:0]   io_coef_out_payload_0_8_46_real,
  output     [15:0]   io_coef_out_payload_0_8_46_imag,
  output     [15:0]   io_coef_out_payload_0_8_47_real,
  output     [15:0]   io_coef_out_payload_0_8_47_imag,
  output     [15:0]   io_coef_out_payload_0_8_48_real,
  output     [15:0]   io_coef_out_payload_0_8_48_imag,
  output     [15:0]   io_coef_out_payload_0_8_49_real,
  output     [15:0]   io_coef_out_payload_0_8_49_imag,
  output     [15:0]   io_coef_out_payload_0_9_0_real,
  output     [15:0]   io_coef_out_payload_0_9_0_imag,
  output     [15:0]   io_coef_out_payload_0_9_1_real,
  output     [15:0]   io_coef_out_payload_0_9_1_imag,
  output     [15:0]   io_coef_out_payload_0_9_2_real,
  output     [15:0]   io_coef_out_payload_0_9_2_imag,
  output     [15:0]   io_coef_out_payload_0_9_3_real,
  output     [15:0]   io_coef_out_payload_0_9_3_imag,
  output     [15:0]   io_coef_out_payload_0_9_4_real,
  output     [15:0]   io_coef_out_payload_0_9_4_imag,
  output     [15:0]   io_coef_out_payload_0_9_5_real,
  output     [15:0]   io_coef_out_payload_0_9_5_imag,
  output     [15:0]   io_coef_out_payload_0_9_6_real,
  output     [15:0]   io_coef_out_payload_0_9_6_imag,
  output     [15:0]   io_coef_out_payload_0_9_7_real,
  output     [15:0]   io_coef_out_payload_0_9_7_imag,
  output     [15:0]   io_coef_out_payload_0_9_8_real,
  output     [15:0]   io_coef_out_payload_0_9_8_imag,
  output     [15:0]   io_coef_out_payload_0_9_9_real,
  output     [15:0]   io_coef_out_payload_0_9_9_imag,
  output     [15:0]   io_coef_out_payload_0_9_10_real,
  output     [15:0]   io_coef_out_payload_0_9_10_imag,
  output     [15:0]   io_coef_out_payload_0_9_11_real,
  output     [15:0]   io_coef_out_payload_0_9_11_imag,
  output     [15:0]   io_coef_out_payload_0_9_12_real,
  output     [15:0]   io_coef_out_payload_0_9_12_imag,
  output     [15:0]   io_coef_out_payload_0_9_13_real,
  output     [15:0]   io_coef_out_payload_0_9_13_imag,
  output     [15:0]   io_coef_out_payload_0_9_14_real,
  output     [15:0]   io_coef_out_payload_0_9_14_imag,
  output     [15:0]   io_coef_out_payload_0_9_15_real,
  output     [15:0]   io_coef_out_payload_0_9_15_imag,
  output     [15:0]   io_coef_out_payload_0_9_16_real,
  output     [15:0]   io_coef_out_payload_0_9_16_imag,
  output     [15:0]   io_coef_out_payload_0_9_17_real,
  output     [15:0]   io_coef_out_payload_0_9_17_imag,
  output     [15:0]   io_coef_out_payload_0_9_18_real,
  output     [15:0]   io_coef_out_payload_0_9_18_imag,
  output     [15:0]   io_coef_out_payload_0_9_19_real,
  output     [15:0]   io_coef_out_payload_0_9_19_imag,
  output     [15:0]   io_coef_out_payload_0_9_20_real,
  output     [15:0]   io_coef_out_payload_0_9_20_imag,
  output     [15:0]   io_coef_out_payload_0_9_21_real,
  output     [15:0]   io_coef_out_payload_0_9_21_imag,
  output     [15:0]   io_coef_out_payload_0_9_22_real,
  output     [15:0]   io_coef_out_payload_0_9_22_imag,
  output     [15:0]   io_coef_out_payload_0_9_23_real,
  output     [15:0]   io_coef_out_payload_0_9_23_imag,
  output     [15:0]   io_coef_out_payload_0_9_24_real,
  output     [15:0]   io_coef_out_payload_0_9_24_imag,
  output     [15:0]   io_coef_out_payload_0_9_25_real,
  output     [15:0]   io_coef_out_payload_0_9_25_imag,
  output     [15:0]   io_coef_out_payload_0_9_26_real,
  output     [15:0]   io_coef_out_payload_0_9_26_imag,
  output     [15:0]   io_coef_out_payload_0_9_27_real,
  output     [15:0]   io_coef_out_payload_0_9_27_imag,
  output     [15:0]   io_coef_out_payload_0_9_28_real,
  output     [15:0]   io_coef_out_payload_0_9_28_imag,
  output     [15:0]   io_coef_out_payload_0_9_29_real,
  output     [15:0]   io_coef_out_payload_0_9_29_imag,
  output     [15:0]   io_coef_out_payload_0_9_30_real,
  output     [15:0]   io_coef_out_payload_0_9_30_imag,
  output     [15:0]   io_coef_out_payload_0_9_31_real,
  output     [15:0]   io_coef_out_payload_0_9_31_imag,
  output     [15:0]   io_coef_out_payload_0_9_32_real,
  output     [15:0]   io_coef_out_payload_0_9_32_imag,
  output     [15:0]   io_coef_out_payload_0_9_33_real,
  output     [15:0]   io_coef_out_payload_0_9_33_imag,
  output     [15:0]   io_coef_out_payload_0_9_34_real,
  output     [15:0]   io_coef_out_payload_0_9_34_imag,
  output     [15:0]   io_coef_out_payload_0_9_35_real,
  output     [15:0]   io_coef_out_payload_0_9_35_imag,
  output     [15:0]   io_coef_out_payload_0_9_36_real,
  output     [15:0]   io_coef_out_payload_0_9_36_imag,
  output     [15:0]   io_coef_out_payload_0_9_37_real,
  output     [15:0]   io_coef_out_payload_0_9_37_imag,
  output     [15:0]   io_coef_out_payload_0_9_38_real,
  output     [15:0]   io_coef_out_payload_0_9_38_imag,
  output     [15:0]   io_coef_out_payload_0_9_39_real,
  output     [15:0]   io_coef_out_payload_0_9_39_imag,
  output     [15:0]   io_coef_out_payload_0_9_40_real,
  output     [15:0]   io_coef_out_payload_0_9_40_imag,
  output     [15:0]   io_coef_out_payload_0_9_41_real,
  output     [15:0]   io_coef_out_payload_0_9_41_imag,
  output     [15:0]   io_coef_out_payload_0_9_42_real,
  output     [15:0]   io_coef_out_payload_0_9_42_imag,
  output     [15:0]   io_coef_out_payload_0_9_43_real,
  output     [15:0]   io_coef_out_payload_0_9_43_imag,
  output     [15:0]   io_coef_out_payload_0_9_44_real,
  output     [15:0]   io_coef_out_payload_0_9_44_imag,
  output     [15:0]   io_coef_out_payload_0_9_45_real,
  output     [15:0]   io_coef_out_payload_0_9_45_imag,
  output     [15:0]   io_coef_out_payload_0_9_46_real,
  output     [15:0]   io_coef_out_payload_0_9_46_imag,
  output     [15:0]   io_coef_out_payload_0_9_47_real,
  output     [15:0]   io_coef_out_payload_0_9_47_imag,
  output     [15:0]   io_coef_out_payload_0_9_48_real,
  output     [15:0]   io_coef_out_payload_0_9_48_imag,
  output     [15:0]   io_coef_out_payload_0_9_49_real,
  output     [15:0]   io_coef_out_payload_0_9_49_imag,
  output     [15:0]   io_coef_out_payload_0_10_0_real,
  output     [15:0]   io_coef_out_payload_0_10_0_imag,
  output     [15:0]   io_coef_out_payload_0_10_1_real,
  output     [15:0]   io_coef_out_payload_0_10_1_imag,
  output     [15:0]   io_coef_out_payload_0_10_2_real,
  output     [15:0]   io_coef_out_payload_0_10_2_imag,
  output     [15:0]   io_coef_out_payload_0_10_3_real,
  output     [15:0]   io_coef_out_payload_0_10_3_imag,
  output     [15:0]   io_coef_out_payload_0_10_4_real,
  output     [15:0]   io_coef_out_payload_0_10_4_imag,
  output     [15:0]   io_coef_out_payload_0_10_5_real,
  output     [15:0]   io_coef_out_payload_0_10_5_imag,
  output     [15:0]   io_coef_out_payload_0_10_6_real,
  output     [15:0]   io_coef_out_payload_0_10_6_imag,
  output     [15:0]   io_coef_out_payload_0_10_7_real,
  output     [15:0]   io_coef_out_payload_0_10_7_imag,
  output     [15:0]   io_coef_out_payload_0_10_8_real,
  output     [15:0]   io_coef_out_payload_0_10_8_imag,
  output     [15:0]   io_coef_out_payload_0_10_9_real,
  output     [15:0]   io_coef_out_payload_0_10_9_imag,
  output     [15:0]   io_coef_out_payload_0_10_10_real,
  output     [15:0]   io_coef_out_payload_0_10_10_imag,
  output     [15:0]   io_coef_out_payload_0_10_11_real,
  output     [15:0]   io_coef_out_payload_0_10_11_imag,
  output     [15:0]   io_coef_out_payload_0_10_12_real,
  output     [15:0]   io_coef_out_payload_0_10_12_imag,
  output     [15:0]   io_coef_out_payload_0_10_13_real,
  output     [15:0]   io_coef_out_payload_0_10_13_imag,
  output     [15:0]   io_coef_out_payload_0_10_14_real,
  output     [15:0]   io_coef_out_payload_0_10_14_imag,
  output     [15:0]   io_coef_out_payload_0_10_15_real,
  output     [15:0]   io_coef_out_payload_0_10_15_imag,
  output     [15:0]   io_coef_out_payload_0_10_16_real,
  output     [15:0]   io_coef_out_payload_0_10_16_imag,
  output     [15:0]   io_coef_out_payload_0_10_17_real,
  output     [15:0]   io_coef_out_payload_0_10_17_imag,
  output     [15:0]   io_coef_out_payload_0_10_18_real,
  output     [15:0]   io_coef_out_payload_0_10_18_imag,
  output     [15:0]   io_coef_out_payload_0_10_19_real,
  output     [15:0]   io_coef_out_payload_0_10_19_imag,
  output     [15:0]   io_coef_out_payload_0_10_20_real,
  output     [15:0]   io_coef_out_payload_0_10_20_imag,
  output     [15:0]   io_coef_out_payload_0_10_21_real,
  output     [15:0]   io_coef_out_payload_0_10_21_imag,
  output     [15:0]   io_coef_out_payload_0_10_22_real,
  output     [15:0]   io_coef_out_payload_0_10_22_imag,
  output     [15:0]   io_coef_out_payload_0_10_23_real,
  output     [15:0]   io_coef_out_payload_0_10_23_imag,
  output     [15:0]   io_coef_out_payload_0_10_24_real,
  output     [15:0]   io_coef_out_payload_0_10_24_imag,
  output     [15:0]   io_coef_out_payload_0_10_25_real,
  output     [15:0]   io_coef_out_payload_0_10_25_imag,
  output     [15:0]   io_coef_out_payload_0_10_26_real,
  output     [15:0]   io_coef_out_payload_0_10_26_imag,
  output     [15:0]   io_coef_out_payload_0_10_27_real,
  output     [15:0]   io_coef_out_payload_0_10_27_imag,
  output     [15:0]   io_coef_out_payload_0_10_28_real,
  output     [15:0]   io_coef_out_payload_0_10_28_imag,
  output     [15:0]   io_coef_out_payload_0_10_29_real,
  output     [15:0]   io_coef_out_payload_0_10_29_imag,
  output     [15:0]   io_coef_out_payload_0_10_30_real,
  output     [15:0]   io_coef_out_payload_0_10_30_imag,
  output     [15:0]   io_coef_out_payload_0_10_31_real,
  output     [15:0]   io_coef_out_payload_0_10_31_imag,
  output     [15:0]   io_coef_out_payload_0_10_32_real,
  output     [15:0]   io_coef_out_payload_0_10_32_imag,
  output     [15:0]   io_coef_out_payload_0_10_33_real,
  output     [15:0]   io_coef_out_payload_0_10_33_imag,
  output     [15:0]   io_coef_out_payload_0_10_34_real,
  output     [15:0]   io_coef_out_payload_0_10_34_imag,
  output     [15:0]   io_coef_out_payload_0_10_35_real,
  output     [15:0]   io_coef_out_payload_0_10_35_imag,
  output     [15:0]   io_coef_out_payload_0_10_36_real,
  output     [15:0]   io_coef_out_payload_0_10_36_imag,
  output     [15:0]   io_coef_out_payload_0_10_37_real,
  output     [15:0]   io_coef_out_payload_0_10_37_imag,
  output     [15:0]   io_coef_out_payload_0_10_38_real,
  output     [15:0]   io_coef_out_payload_0_10_38_imag,
  output     [15:0]   io_coef_out_payload_0_10_39_real,
  output     [15:0]   io_coef_out_payload_0_10_39_imag,
  output     [15:0]   io_coef_out_payload_0_10_40_real,
  output     [15:0]   io_coef_out_payload_0_10_40_imag,
  output     [15:0]   io_coef_out_payload_0_10_41_real,
  output     [15:0]   io_coef_out_payload_0_10_41_imag,
  output     [15:0]   io_coef_out_payload_0_10_42_real,
  output     [15:0]   io_coef_out_payload_0_10_42_imag,
  output     [15:0]   io_coef_out_payload_0_10_43_real,
  output     [15:0]   io_coef_out_payload_0_10_43_imag,
  output     [15:0]   io_coef_out_payload_0_10_44_real,
  output     [15:0]   io_coef_out_payload_0_10_44_imag,
  output     [15:0]   io_coef_out_payload_0_10_45_real,
  output     [15:0]   io_coef_out_payload_0_10_45_imag,
  output     [15:0]   io_coef_out_payload_0_10_46_real,
  output     [15:0]   io_coef_out_payload_0_10_46_imag,
  output     [15:0]   io_coef_out_payload_0_10_47_real,
  output     [15:0]   io_coef_out_payload_0_10_47_imag,
  output     [15:0]   io_coef_out_payload_0_10_48_real,
  output     [15:0]   io_coef_out_payload_0_10_48_imag,
  output     [15:0]   io_coef_out_payload_0_10_49_real,
  output     [15:0]   io_coef_out_payload_0_10_49_imag,
  output     [15:0]   io_coef_out_payload_0_11_0_real,
  output     [15:0]   io_coef_out_payload_0_11_0_imag,
  output     [15:0]   io_coef_out_payload_0_11_1_real,
  output     [15:0]   io_coef_out_payload_0_11_1_imag,
  output     [15:0]   io_coef_out_payload_0_11_2_real,
  output     [15:0]   io_coef_out_payload_0_11_2_imag,
  output     [15:0]   io_coef_out_payload_0_11_3_real,
  output     [15:0]   io_coef_out_payload_0_11_3_imag,
  output     [15:0]   io_coef_out_payload_0_11_4_real,
  output     [15:0]   io_coef_out_payload_0_11_4_imag,
  output     [15:0]   io_coef_out_payload_0_11_5_real,
  output     [15:0]   io_coef_out_payload_0_11_5_imag,
  output     [15:0]   io_coef_out_payload_0_11_6_real,
  output     [15:0]   io_coef_out_payload_0_11_6_imag,
  output     [15:0]   io_coef_out_payload_0_11_7_real,
  output     [15:0]   io_coef_out_payload_0_11_7_imag,
  output     [15:0]   io_coef_out_payload_0_11_8_real,
  output     [15:0]   io_coef_out_payload_0_11_8_imag,
  output     [15:0]   io_coef_out_payload_0_11_9_real,
  output     [15:0]   io_coef_out_payload_0_11_9_imag,
  output     [15:0]   io_coef_out_payload_0_11_10_real,
  output     [15:0]   io_coef_out_payload_0_11_10_imag,
  output     [15:0]   io_coef_out_payload_0_11_11_real,
  output     [15:0]   io_coef_out_payload_0_11_11_imag,
  output     [15:0]   io_coef_out_payload_0_11_12_real,
  output     [15:0]   io_coef_out_payload_0_11_12_imag,
  output     [15:0]   io_coef_out_payload_0_11_13_real,
  output     [15:0]   io_coef_out_payload_0_11_13_imag,
  output     [15:0]   io_coef_out_payload_0_11_14_real,
  output     [15:0]   io_coef_out_payload_0_11_14_imag,
  output     [15:0]   io_coef_out_payload_0_11_15_real,
  output     [15:0]   io_coef_out_payload_0_11_15_imag,
  output     [15:0]   io_coef_out_payload_0_11_16_real,
  output     [15:0]   io_coef_out_payload_0_11_16_imag,
  output     [15:0]   io_coef_out_payload_0_11_17_real,
  output     [15:0]   io_coef_out_payload_0_11_17_imag,
  output     [15:0]   io_coef_out_payload_0_11_18_real,
  output     [15:0]   io_coef_out_payload_0_11_18_imag,
  output     [15:0]   io_coef_out_payload_0_11_19_real,
  output     [15:0]   io_coef_out_payload_0_11_19_imag,
  output     [15:0]   io_coef_out_payload_0_11_20_real,
  output     [15:0]   io_coef_out_payload_0_11_20_imag,
  output     [15:0]   io_coef_out_payload_0_11_21_real,
  output     [15:0]   io_coef_out_payload_0_11_21_imag,
  output     [15:0]   io_coef_out_payload_0_11_22_real,
  output     [15:0]   io_coef_out_payload_0_11_22_imag,
  output     [15:0]   io_coef_out_payload_0_11_23_real,
  output     [15:0]   io_coef_out_payload_0_11_23_imag,
  output     [15:0]   io_coef_out_payload_0_11_24_real,
  output     [15:0]   io_coef_out_payload_0_11_24_imag,
  output     [15:0]   io_coef_out_payload_0_11_25_real,
  output     [15:0]   io_coef_out_payload_0_11_25_imag,
  output     [15:0]   io_coef_out_payload_0_11_26_real,
  output     [15:0]   io_coef_out_payload_0_11_26_imag,
  output     [15:0]   io_coef_out_payload_0_11_27_real,
  output     [15:0]   io_coef_out_payload_0_11_27_imag,
  output     [15:0]   io_coef_out_payload_0_11_28_real,
  output     [15:0]   io_coef_out_payload_0_11_28_imag,
  output     [15:0]   io_coef_out_payload_0_11_29_real,
  output     [15:0]   io_coef_out_payload_0_11_29_imag,
  output     [15:0]   io_coef_out_payload_0_11_30_real,
  output     [15:0]   io_coef_out_payload_0_11_30_imag,
  output     [15:0]   io_coef_out_payload_0_11_31_real,
  output     [15:0]   io_coef_out_payload_0_11_31_imag,
  output     [15:0]   io_coef_out_payload_0_11_32_real,
  output     [15:0]   io_coef_out_payload_0_11_32_imag,
  output     [15:0]   io_coef_out_payload_0_11_33_real,
  output     [15:0]   io_coef_out_payload_0_11_33_imag,
  output     [15:0]   io_coef_out_payload_0_11_34_real,
  output     [15:0]   io_coef_out_payload_0_11_34_imag,
  output     [15:0]   io_coef_out_payload_0_11_35_real,
  output     [15:0]   io_coef_out_payload_0_11_35_imag,
  output     [15:0]   io_coef_out_payload_0_11_36_real,
  output     [15:0]   io_coef_out_payload_0_11_36_imag,
  output     [15:0]   io_coef_out_payload_0_11_37_real,
  output     [15:0]   io_coef_out_payload_0_11_37_imag,
  output     [15:0]   io_coef_out_payload_0_11_38_real,
  output     [15:0]   io_coef_out_payload_0_11_38_imag,
  output     [15:0]   io_coef_out_payload_0_11_39_real,
  output     [15:0]   io_coef_out_payload_0_11_39_imag,
  output     [15:0]   io_coef_out_payload_0_11_40_real,
  output     [15:0]   io_coef_out_payload_0_11_40_imag,
  output     [15:0]   io_coef_out_payload_0_11_41_real,
  output     [15:0]   io_coef_out_payload_0_11_41_imag,
  output     [15:0]   io_coef_out_payload_0_11_42_real,
  output     [15:0]   io_coef_out_payload_0_11_42_imag,
  output     [15:0]   io_coef_out_payload_0_11_43_real,
  output     [15:0]   io_coef_out_payload_0_11_43_imag,
  output     [15:0]   io_coef_out_payload_0_11_44_real,
  output     [15:0]   io_coef_out_payload_0_11_44_imag,
  output     [15:0]   io_coef_out_payload_0_11_45_real,
  output     [15:0]   io_coef_out_payload_0_11_45_imag,
  output     [15:0]   io_coef_out_payload_0_11_46_real,
  output     [15:0]   io_coef_out_payload_0_11_46_imag,
  output     [15:0]   io_coef_out_payload_0_11_47_real,
  output     [15:0]   io_coef_out_payload_0_11_47_imag,
  output     [15:0]   io_coef_out_payload_0_11_48_real,
  output     [15:0]   io_coef_out_payload_0_11_48_imag,
  output     [15:0]   io_coef_out_payload_0_11_49_real,
  output     [15:0]   io_coef_out_payload_0_11_49_imag,
  output     [15:0]   io_coef_out_payload_0_12_0_real,
  output     [15:0]   io_coef_out_payload_0_12_0_imag,
  output     [15:0]   io_coef_out_payload_0_12_1_real,
  output     [15:0]   io_coef_out_payload_0_12_1_imag,
  output     [15:0]   io_coef_out_payload_0_12_2_real,
  output     [15:0]   io_coef_out_payload_0_12_2_imag,
  output     [15:0]   io_coef_out_payload_0_12_3_real,
  output     [15:0]   io_coef_out_payload_0_12_3_imag,
  output     [15:0]   io_coef_out_payload_0_12_4_real,
  output     [15:0]   io_coef_out_payload_0_12_4_imag,
  output     [15:0]   io_coef_out_payload_0_12_5_real,
  output     [15:0]   io_coef_out_payload_0_12_5_imag,
  output     [15:0]   io_coef_out_payload_0_12_6_real,
  output     [15:0]   io_coef_out_payload_0_12_6_imag,
  output     [15:0]   io_coef_out_payload_0_12_7_real,
  output     [15:0]   io_coef_out_payload_0_12_7_imag,
  output     [15:0]   io_coef_out_payload_0_12_8_real,
  output     [15:0]   io_coef_out_payload_0_12_8_imag,
  output     [15:0]   io_coef_out_payload_0_12_9_real,
  output     [15:0]   io_coef_out_payload_0_12_9_imag,
  output     [15:0]   io_coef_out_payload_0_12_10_real,
  output     [15:0]   io_coef_out_payload_0_12_10_imag,
  output     [15:0]   io_coef_out_payload_0_12_11_real,
  output     [15:0]   io_coef_out_payload_0_12_11_imag,
  output     [15:0]   io_coef_out_payload_0_12_12_real,
  output     [15:0]   io_coef_out_payload_0_12_12_imag,
  output     [15:0]   io_coef_out_payload_0_12_13_real,
  output     [15:0]   io_coef_out_payload_0_12_13_imag,
  output     [15:0]   io_coef_out_payload_0_12_14_real,
  output     [15:0]   io_coef_out_payload_0_12_14_imag,
  output     [15:0]   io_coef_out_payload_0_12_15_real,
  output     [15:0]   io_coef_out_payload_0_12_15_imag,
  output     [15:0]   io_coef_out_payload_0_12_16_real,
  output     [15:0]   io_coef_out_payload_0_12_16_imag,
  output     [15:0]   io_coef_out_payload_0_12_17_real,
  output     [15:0]   io_coef_out_payload_0_12_17_imag,
  output     [15:0]   io_coef_out_payload_0_12_18_real,
  output     [15:0]   io_coef_out_payload_0_12_18_imag,
  output     [15:0]   io_coef_out_payload_0_12_19_real,
  output     [15:0]   io_coef_out_payload_0_12_19_imag,
  output     [15:0]   io_coef_out_payload_0_12_20_real,
  output     [15:0]   io_coef_out_payload_0_12_20_imag,
  output     [15:0]   io_coef_out_payload_0_12_21_real,
  output     [15:0]   io_coef_out_payload_0_12_21_imag,
  output     [15:0]   io_coef_out_payload_0_12_22_real,
  output     [15:0]   io_coef_out_payload_0_12_22_imag,
  output     [15:0]   io_coef_out_payload_0_12_23_real,
  output     [15:0]   io_coef_out_payload_0_12_23_imag,
  output     [15:0]   io_coef_out_payload_0_12_24_real,
  output     [15:0]   io_coef_out_payload_0_12_24_imag,
  output     [15:0]   io_coef_out_payload_0_12_25_real,
  output     [15:0]   io_coef_out_payload_0_12_25_imag,
  output     [15:0]   io_coef_out_payload_0_12_26_real,
  output     [15:0]   io_coef_out_payload_0_12_26_imag,
  output     [15:0]   io_coef_out_payload_0_12_27_real,
  output     [15:0]   io_coef_out_payload_0_12_27_imag,
  output     [15:0]   io_coef_out_payload_0_12_28_real,
  output     [15:0]   io_coef_out_payload_0_12_28_imag,
  output     [15:0]   io_coef_out_payload_0_12_29_real,
  output     [15:0]   io_coef_out_payload_0_12_29_imag,
  output     [15:0]   io_coef_out_payload_0_12_30_real,
  output     [15:0]   io_coef_out_payload_0_12_30_imag,
  output     [15:0]   io_coef_out_payload_0_12_31_real,
  output     [15:0]   io_coef_out_payload_0_12_31_imag,
  output     [15:0]   io_coef_out_payload_0_12_32_real,
  output     [15:0]   io_coef_out_payload_0_12_32_imag,
  output     [15:0]   io_coef_out_payload_0_12_33_real,
  output     [15:0]   io_coef_out_payload_0_12_33_imag,
  output     [15:0]   io_coef_out_payload_0_12_34_real,
  output     [15:0]   io_coef_out_payload_0_12_34_imag,
  output     [15:0]   io_coef_out_payload_0_12_35_real,
  output     [15:0]   io_coef_out_payload_0_12_35_imag,
  output     [15:0]   io_coef_out_payload_0_12_36_real,
  output     [15:0]   io_coef_out_payload_0_12_36_imag,
  output     [15:0]   io_coef_out_payload_0_12_37_real,
  output     [15:0]   io_coef_out_payload_0_12_37_imag,
  output     [15:0]   io_coef_out_payload_0_12_38_real,
  output     [15:0]   io_coef_out_payload_0_12_38_imag,
  output     [15:0]   io_coef_out_payload_0_12_39_real,
  output     [15:0]   io_coef_out_payload_0_12_39_imag,
  output     [15:0]   io_coef_out_payload_0_12_40_real,
  output     [15:0]   io_coef_out_payload_0_12_40_imag,
  output     [15:0]   io_coef_out_payload_0_12_41_real,
  output     [15:0]   io_coef_out_payload_0_12_41_imag,
  output     [15:0]   io_coef_out_payload_0_12_42_real,
  output     [15:0]   io_coef_out_payload_0_12_42_imag,
  output     [15:0]   io_coef_out_payload_0_12_43_real,
  output     [15:0]   io_coef_out_payload_0_12_43_imag,
  output     [15:0]   io_coef_out_payload_0_12_44_real,
  output     [15:0]   io_coef_out_payload_0_12_44_imag,
  output     [15:0]   io_coef_out_payload_0_12_45_real,
  output     [15:0]   io_coef_out_payload_0_12_45_imag,
  output     [15:0]   io_coef_out_payload_0_12_46_real,
  output     [15:0]   io_coef_out_payload_0_12_46_imag,
  output     [15:0]   io_coef_out_payload_0_12_47_real,
  output     [15:0]   io_coef_out_payload_0_12_47_imag,
  output     [15:0]   io_coef_out_payload_0_12_48_real,
  output     [15:0]   io_coef_out_payload_0_12_48_imag,
  output     [15:0]   io_coef_out_payload_0_12_49_real,
  output     [15:0]   io_coef_out_payload_0_12_49_imag,
  output     [15:0]   io_coef_out_payload_0_13_0_real,
  output     [15:0]   io_coef_out_payload_0_13_0_imag,
  output     [15:0]   io_coef_out_payload_0_13_1_real,
  output     [15:0]   io_coef_out_payload_0_13_1_imag,
  output     [15:0]   io_coef_out_payload_0_13_2_real,
  output     [15:0]   io_coef_out_payload_0_13_2_imag,
  output     [15:0]   io_coef_out_payload_0_13_3_real,
  output     [15:0]   io_coef_out_payload_0_13_3_imag,
  output     [15:0]   io_coef_out_payload_0_13_4_real,
  output     [15:0]   io_coef_out_payload_0_13_4_imag,
  output     [15:0]   io_coef_out_payload_0_13_5_real,
  output     [15:0]   io_coef_out_payload_0_13_5_imag,
  output     [15:0]   io_coef_out_payload_0_13_6_real,
  output     [15:0]   io_coef_out_payload_0_13_6_imag,
  output     [15:0]   io_coef_out_payload_0_13_7_real,
  output     [15:0]   io_coef_out_payload_0_13_7_imag,
  output     [15:0]   io_coef_out_payload_0_13_8_real,
  output     [15:0]   io_coef_out_payload_0_13_8_imag,
  output     [15:0]   io_coef_out_payload_0_13_9_real,
  output     [15:0]   io_coef_out_payload_0_13_9_imag,
  output     [15:0]   io_coef_out_payload_0_13_10_real,
  output     [15:0]   io_coef_out_payload_0_13_10_imag,
  output     [15:0]   io_coef_out_payload_0_13_11_real,
  output     [15:0]   io_coef_out_payload_0_13_11_imag,
  output     [15:0]   io_coef_out_payload_0_13_12_real,
  output     [15:0]   io_coef_out_payload_0_13_12_imag,
  output     [15:0]   io_coef_out_payload_0_13_13_real,
  output     [15:0]   io_coef_out_payload_0_13_13_imag,
  output     [15:0]   io_coef_out_payload_0_13_14_real,
  output     [15:0]   io_coef_out_payload_0_13_14_imag,
  output     [15:0]   io_coef_out_payload_0_13_15_real,
  output     [15:0]   io_coef_out_payload_0_13_15_imag,
  output     [15:0]   io_coef_out_payload_0_13_16_real,
  output     [15:0]   io_coef_out_payload_0_13_16_imag,
  output     [15:0]   io_coef_out_payload_0_13_17_real,
  output     [15:0]   io_coef_out_payload_0_13_17_imag,
  output     [15:0]   io_coef_out_payload_0_13_18_real,
  output     [15:0]   io_coef_out_payload_0_13_18_imag,
  output     [15:0]   io_coef_out_payload_0_13_19_real,
  output     [15:0]   io_coef_out_payload_0_13_19_imag,
  output     [15:0]   io_coef_out_payload_0_13_20_real,
  output     [15:0]   io_coef_out_payload_0_13_20_imag,
  output     [15:0]   io_coef_out_payload_0_13_21_real,
  output     [15:0]   io_coef_out_payload_0_13_21_imag,
  output     [15:0]   io_coef_out_payload_0_13_22_real,
  output     [15:0]   io_coef_out_payload_0_13_22_imag,
  output     [15:0]   io_coef_out_payload_0_13_23_real,
  output     [15:0]   io_coef_out_payload_0_13_23_imag,
  output     [15:0]   io_coef_out_payload_0_13_24_real,
  output     [15:0]   io_coef_out_payload_0_13_24_imag,
  output     [15:0]   io_coef_out_payload_0_13_25_real,
  output     [15:0]   io_coef_out_payload_0_13_25_imag,
  output     [15:0]   io_coef_out_payload_0_13_26_real,
  output     [15:0]   io_coef_out_payload_0_13_26_imag,
  output     [15:0]   io_coef_out_payload_0_13_27_real,
  output     [15:0]   io_coef_out_payload_0_13_27_imag,
  output     [15:0]   io_coef_out_payload_0_13_28_real,
  output     [15:0]   io_coef_out_payload_0_13_28_imag,
  output     [15:0]   io_coef_out_payload_0_13_29_real,
  output     [15:0]   io_coef_out_payload_0_13_29_imag,
  output     [15:0]   io_coef_out_payload_0_13_30_real,
  output     [15:0]   io_coef_out_payload_0_13_30_imag,
  output     [15:0]   io_coef_out_payload_0_13_31_real,
  output     [15:0]   io_coef_out_payload_0_13_31_imag,
  output     [15:0]   io_coef_out_payload_0_13_32_real,
  output     [15:0]   io_coef_out_payload_0_13_32_imag,
  output     [15:0]   io_coef_out_payload_0_13_33_real,
  output     [15:0]   io_coef_out_payload_0_13_33_imag,
  output     [15:0]   io_coef_out_payload_0_13_34_real,
  output     [15:0]   io_coef_out_payload_0_13_34_imag,
  output     [15:0]   io_coef_out_payload_0_13_35_real,
  output     [15:0]   io_coef_out_payload_0_13_35_imag,
  output     [15:0]   io_coef_out_payload_0_13_36_real,
  output     [15:0]   io_coef_out_payload_0_13_36_imag,
  output     [15:0]   io_coef_out_payload_0_13_37_real,
  output     [15:0]   io_coef_out_payload_0_13_37_imag,
  output     [15:0]   io_coef_out_payload_0_13_38_real,
  output     [15:0]   io_coef_out_payload_0_13_38_imag,
  output     [15:0]   io_coef_out_payload_0_13_39_real,
  output     [15:0]   io_coef_out_payload_0_13_39_imag,
  output     [15:0]   io_coef_out_payload_0_13_40_real,
  output     [15:0]   io_coef_out_payload_0_13_40_imag,
  output     [15:0]   io_coef_out_payload_0_13_41_real,
  output     [15:0]   io_coef_out_payload_0_13_41_imag,
  output     [15:0]   io_coef_out_payload_0_13_42_real,
  output     [15:0]   io_coef_out_payload_0_13_42_imag,
  output     [15:0]   io_coef_out_payload_0_13_43_real,
  output     [15:0]   io_coef_out_payload_0_13_43_imag,
  output     [15:0]   io_coef_out_payload_0_13_44_real,
  output     [15:0]   io_coef_out_payload_0_13_44_imag,
  output     [15:0]   io_coef_out_payload_0_13_45_real,
  output     [15:0]   io_coef_out_payload_0_13_45_imag,
  output     [15:0]   io_coef_out_payload_0_13_46_real,
  output     [15:0]   io_coef_out_payload_0_13_46_imag,
  output     [15:0]   io_coef_out_payload_0_13_47_real,
  output     [15:0]   io_coef_out_payload_0_13_47_imag,
  output     [15:0]   io_coef_out_payload_0_13_48_real,
  output     [15:0]   io_coef_out_payload_0_13_48_imag,
  output     [15:0]   io_coef_out_payload_0_13_49_real,
  output     [15:0]   io_coef_out_payload_0_13_49_imag,
  output     [15:0]   io_coef_out_payload_0_14_0_real,
  output     [15:0]   io_coef_out_payload_0_14_0_imag,
  output     [15:0]   io_coef_out_payload_0_14_1_real,
  output     [15:0]   io_coef_out_payload_0_14_1_imag,
  output     [15:0]   io_coef_out_payload_0_14_2_real,
  output     [15:0]   io_coef_out_payload_0_14_2_imag,
  output     [15:0]   io_coef_out_payload_0_14_3_real,
  output     [15:0]   io_coef_out_payload_0_14_3_imag,
  output     [15:0]   io_coef_out_payload_0_14_4_real,
  output     [15:0]   io_coef_out_payload_0_14_4_imag,
  output     [15:0]   io_coef_out_payload_0_14_5_real,
  output     [15:0]   io_coef_out_payload_0_14_5_imag,
  output     [15:0]   io_coef_out_payload_0_14_6_real,
  output     [15:0]   io_coef_out_payload_0_14_6_imag,
  output     [15:0]   io_coef_out_payload_0_14_7_real,
  output     [15:0]   io_coef_out_payload_0_14_7_imag,
  output     [15:0]   io_coef_out_payload_0_14_8_real,
  output     [15:0]   io_coef_out_payload_0_14_8_imag,
  output     [15:0]   io_coef_out_payload_0_14_9_real,
  output     [15:0]   io_coef_out_payload_0_14_9_imag,
  output     [15:0]   io_coef_out_payload_0_14_10_real,
  output     [15:0]   io_coef_out_payload_0_14_10_imag,
  output     [15:0]   io_coef_out_payload_0_14_11_real,
  output     [15:0]   io_coef_out_payload_0_14_11_imag,
  output     [15:0]   io_coef_out_payload_0_14_12_real,
  output     [15:0]   io_coef_out_payload_0_14_12_imag,
  output     [15:0]   io_coef_out_payload_0_14_13_real,
  output     [15:0]   io_coef_out_payload_0_14_13_imag,
  output     [15:0]   io_coef_out_payload_0_14_14_real,
  output     [15:0]   io_coef_out_payload_0_14_14_imag,
  output     [15:0]   io_coef_out_payload_0_14_15_real,
  output     [15:0]   io_coef_out_payload_0_14_15_imag,
  output     [15:0]   io_coef_out_payload_0_14_16_real,
  output     [15:0]   io_coef_out_payload_0_14_16_imag,
  output     [15:0]   io_coef_out_payload_0_14_17_real,
  output     [15:0]   io_coef_out_payload_0_14_17_imag,
  output     [15:0]   io_coef_out_payload_0_14_18_real,
  output     [15:0]   io_coef_out_payload_0_14_18_imag,
  output     [15:0]   io_coef_out_payload_0_14_19_real,
  output     [15:0]   io_coef_out_payload_0_14_19_imag,
  output     [15:0]   io_coef_out_payload_0_14_20_real,
  output     [15:0]   io_coef_out_payload_0_14_20_imag,
  output     [15:0]   io_coef_out_payload_0_14_21_real,
  output     [15:0]   io_coef_out_payload_0_14_21_imag,
  output     [15:0]   io_coef_out_payload_0_14_22_real,
  output     [15:0]   io_coef_out_payload_0_14_22_imag,
  output     [15:0]   io_coef_out_payload_0_14_23_real,
  output     [15:0]   io_coef_out_payload_0_14_23_imag,
  output     [15:0]   io_coef_out_payload_0_14_24_real,
  output     [15:0]   io_coef_out_payload_0_14_24_imag,
  output     [15:0]   io_coef_out_payload_0_14_25_real,
  output     [15:0]   io_coef_out_payload_0_14_25_imag,
  output     [15:0]   io_coef_out_payload_0_14_26_real,
  output     [15:0]   io_coef_out_payload_0_14_26_imag,
  output     [15:0]   io_coef_out_payload_0_14_27_real,
  output     [15:0]   io_coef_out_payload_0_14_27_imag,
  output     [15:0]   io_coef_out_payload_0_14_28_real,
  output     [15:0]   io_coef_out_payload_0_14_28_imag,
  output     [15:0]   io_coef_out_payload_0_14_29_real,
  output     [15:0]   io_coef_out_payload_0_14_29_imag,
  output     [15:0]   io_coef_out_payload_0_14_30_real,
  output     [15:0]   io_coef_out_payload_0_14_30_imag,
  output     [15:0]   io_coef_out_payload_0_14_31_real,
  output     [15:0]   io_coef_out_payload_0_14_31_imag,
  output     [15:0]   io_coef_out_payload_0_14_32_real,
  output     [15:0]   io_coef_out_payload_0_14_32_imag,
  output     [15:0]   io_coef_out_payload_0_14_33_real,
  output     [15:0]   io_coef_out_payload_0_14_33_imag,
  output     [15:0]   io_coef_out_payload_0_14_34_real,
  output     [15:0]   io_coef_out_payload_0_14_34_imag,
  output     [15:0]   io_coef_out_payload_0_14_35_real,
  output     [15:0]   io_coef_out_payload_0_14_35_imag,
  output     [15:0]   io_coef_out_payload_0_14_36_real,
  output     [15:0]   io_coef_out_payload_0_14_36_imag,
  output     [15:0]   io_coef_out_payload_0_14_37_real,
  output     [15:0]   io_coef_out_payload_0_14_37_imag,
  output     [15:0]   io_coef_out_payload_0_14_38_real,
  output     [15:0]   io_coef_out_payload_0_14_38_imag,
  output     [15:0]   io_coef_out_payload_0_14_39_real,
  output     [15:0]   io_coef_out_payload_0_14_39_imag,
  output     [15:0]   io_coef_out_payload_0_14_40_real,
  output     [15:0]   io_coef_out_payload_0_14_40_imag,
  output     [15:0]   io_coef_out_payload_0_14_41_real,
  output     [15:0]   io_coef_out_payload_0_14_41_imag,
  output     [15:0]   io_coef_out_payload_0_14_42_real,
  output     [15:0]   io_coef_out_payload_0_14_42_imag,
  output     [15:0]   io_coef_out_payload_0_14_43_real,
  output     [15:0]   io_coef_out_payload_0_14_43_imag,
  output     [15:0]   io_coef_out_payload_0_14_44_real,
  output     [15:0]   io_coef_out_payload_0_14_44_imag,
  output     [15:0]   io_coef_out_payload_0_14_45_real,
  output     [15:0]   io_coef_out_payload_0_14_45_imag,
  output     [15:0]   io_coef_out_payload_0_14_46_real,
  output     [15:0]   io_coef_out_payload_0_14_46_imag,
  output     [15:0]   io_coef_out_payload_0_14_47_real,
  output     [15:0]   io_coef_out_payload_0_14_47_imag,
  output     [15:0]   io_coef_out_payload_0_14_48_real,
  output     [15:0]   io_coef_out_payload_0_14_48_imag,
  output     [15:0]   io_coef_out_payload_0_14_49_real,
  output     [15:0]   io_coef_out_payload_0_14_49_imag,
  output     [15:0]   io_coef_out_payload_0_15_0_real,
  output     [15:0]   io_coef_out_payload_0_15_0_imag,
  output     [15:0]   io_coef_out_payload_0_15_1_real,
  output     [15:0]   io_coef_out_payload_0_15_1_imag,
  output     [15:0]   io_coef_out_payload_0_15_2_real,
  output     [15:0]   io_coef_out_payload_0_15_2_imag,
  output     [15:0]   io_coef_out_payload_0_15_3_real,
  output     [15:0]   io_coef_out_payload_0_15_3_imag,
  output     [15:0]   io_coef_out_payload_0_15_4_real,
  output     [15:0]   io_coef_out_payload_0_15_4_imag,
  output     [15:0]   io_coef_out_payload_0_15_5_real,
  output     [15:0]   io_coef_out_payload_0_15_5_imag,
  output     [15:0]   io_coef_out_payload_0_15_6_real,
  output     [15:0]   io_coef_out_payload_0_15_6_imag,
  output     [15:0]   io_coef_out_payload_0_15_7_real,
  output     [15:0]   io_coef_out_payload_0_15_7_imag,
  output     [15:0]   io_coef_out_payload_0_15_8_real,
  output     [15:0]   io_coef_out_payload_0_15_8_imag,
  output     [15:0]   io_coef_out_payload_0_15_9_real,
  output     [15:0]   io_coef_out_payload_0_15_9_imag,
  output     [15:0]   io_coef_out_payload_0_15_10_real,
  output     [15:0]   io_coef_out_payload_0_15_10_imag,
  output     [15:0]   io_coef_out_payload_0_15_11_real,
  output     [15:0]   io_coef_out_payload_0_15_11_imag,
  output     [15:0]   io_coef_out_payload_0_15_12_real,
  output     [15:0]   io_coef_out_payload_0_15_12_imag,
  output     [15:0]   io_coef_out_payload_0_15_13_real,
  output     [15:0]   io_coef_out_payload_0_15_13_imag,
  output     [15:0]   io_coef_out_payload_0_15_14_real,
  output     [15:0]   io_coef_out_payload_0_15_14_imag,
  output     [15:0]   io_coef_out_payload_0_15_15_real,
  output     [15:0]   io_coef_out_payload_0_15_15_imag,
  output     [15:0]   io_coef_out_payload_0_15_16_real,
  output     [15:0]   io_coef_out_payload_0_15_16_imag,
  output     [15:0]   io_coef_out_payload_0_15_17_real,
  output     [15:0]   io_coef_out_payload_0_15_17_imag,
  output     [15:0]   io_coef_out_payload_0_15_18_real,
  output     [15:0]   io_coef_out_payload_0_15_18_imag,
  output     [15:0]   io_coef_out_payload_0_15_19_real,
  output     [15:0]   io_coef_out_payload_0_15_19_imag,
  output     [15:0]   io_coef_out_payload_0_15_20_real,
  output     [15:0]   io_coef_out_payload_0_15_20_imag,
  output     [15:0]   io_coef_out_payload_0_15_21_real,
  output     [15:0]   io_coef_out_payload_0_15_21_imag,
  output     [15:0]   io_coef_out_payload_0_15_22_real,
  output     [15:0]   io_coef_out_payload_0_15_22_imag,
  output     [15:0]   io_coef_out_payload_0_15_23_real,
  output     [15:0]   io_coef_out_payload_0_15_23_imag,
  output     [15:0]   io_coef_out_payload_0_15_24_real,
  output     [15:0]   io_coef_out_payload_0_15_24_imag,
  output     [15:0]   io_coef_out_payload_0_15_25_real,
  output     [15:0]   io_coef_out_payload_0_15_25_imag,
  output     [15:0]   io_coef_out_payload_0_15_26_real,
  output     [15:0]   io_coef_out_payload_0_15_26_imag,
  output     [15:0]   io_coef_out_payload_0_15_27_real,
  output     [15:0]   io_coef_out_payload_0_15_27_imag,
  output     [15:0]   io_coef_out_payload_0_15_28_real,
  output     [15:0]   io_coef_out_payload_0_15_28_imag,
  output     [15:0]   io_coef_out_payload_0_15_29_real,
  output     [15:0]   io_coef_out_payload_0_15_29_imag,
  output     [15:0]   io_coef_out_payload_0_15_30_real,
  output     [15:0]   io_coef_out_payload_0_15_30_imag,
  output     [15:0]   io_coef_out_payload_0_15_31_real,
  output     [15:0]   io_coef_out_payload_0_15_31_imag,
  output     [15:0]   io_coef_out_payload_0_15_32_real,
  output     [15:0]   io_coef_out_payload_0_15_32_imag,
  output     [15:0]   io_coef_out_payload_0_15_33_real,
  output     [15:0]   io_coef_out_payload_0_15_33_imag,
  output     [15:0]   io_coef_out_payload_0_15_34_real,
  output     [15:0]   io_coef_out_payload_0_15_34_imag,
  output     [15:0]   io_coef_out_payload_0_15_35_real,
  output     [15:0]   io_coef_out_payload_0_15_35_imag,
  output     [15:0]   io_coef_out_payload_0_15_36_real,
  output     [15:0]   io_coef_out_payload_0_15_36_imag,
  output     [15:0]   io_coef_out_payload_0_15_37_real,
  output     [15:0]   io_coef_out_payload_0_15_37_imag,
  output     [15:0]   io_coef_out_payload_0_15_38_real,
  output     [15:0]   io_coef_out_payload_0_15_38_imag,
  output     [15:0]   io_coef_out_payload_0_15_39_real,
  output     [15:0]   io_coef_out_payload_0_15_39_imag,
  output     [15:0]   io_coef_out_payload_0_15_40_real,
  output     [15:0]   io_coef_out_payload_0_15_40_imag,
  output     [15:0]   io_coef_out_payload_0_15_41_real,
  output     [15:0]   io_coef_out_payload_0_15_41_imag,
  output     [15:0]   io_coef_out_payload_0_15_42_real,
  output     [15:0]   io_coef_out_payload_0_15_42_imag,
  output     [15:0]   io_coef_out_payload_0_15_43_real,
  output     [15:0]   io_coef_out_payload_0_15_43_imag,
  output     [15:0]   io_coef_out_payload_0_15_44_real,
  output     [15:0]   io_coef_out_payload_0_15_44_imag,
  output     [15:0]   io_coef_out_payload_0_15_45_real,
  output     [15:0]   io_coef_out_payload_0_15_45_imag,
  output     [15:0]   io_coef_out_payload_0_15_46_real,
  output     [15:0]   io_coef_out_payload_0_15_46_imag,
  output     [15:0]   io_coef_out_payload_0_15_47_real,
  output     [15:0]   io_coef_out_payload_0_15_47_imag,
  output     [15:0]   io_coef_out_payload_0_15_48_real,
  output     [15:0]   io_coef_out_payload_0_15_48_imag,
  output     [15:0]   io_coef_out_payload_0_15_49_real,
  output     [15:0]   io_coef_out_payload_0_15_49_imag,
  output     [15:0]   io_coef_out_payload_0_16_0_real,
  output     [15:0]   io_coef_out_payload_0_16_0_imag,
  output     [15:0]   io_coef_out_payload_0_16_1_real,
  output     [15:0]   io_coef_out_payload_0_16_1_imag,
  output     [15:0]   io_coef_out_payload_0_16_2_real,
  output     [15:0]   io_coef_out_payload_0_16_2_imag,
  output     [15:0]   io_coef_out_payload_0_16_3_real,
  output     [15:0]   io_coef_out_payload_0_16_3_imag,
  output     [15:0]   io_coef_out_payload_0_16_4_real,
  output     [15:0]   io_coef_out_payload_0_16_4_imag,
  output     [15:0]   io_coef_out_payload_0_16_5_real,
  output     [15:0]   io_coef_out_payload_0_16_5_imag,
  output     [15:0]   io_coef_out_payload_0_16_6_real,
  output     [15:0]   io_coef_out_payload_0_16_6_imag,
  output     [15:0]   io_coef_out_payload_0_16_7_real,
  output     [15:0]   io_coef_out_payload_0_16_7_imag,
  output     [15:0]   io_coef_out_payload_0_16_8_real,
  output     [15:0]   io_coef_out_payload_0_16_8_imag,
  output     [15:0]   io_coef_out_payload_0_16_9_real,
  output     [15:0]   io_coef_out_payload_0_16_9_imag,
  output     [15:0]   io_coef_out_payload_0_16_10_real,
  output     [15:0]   io_coef_out_payload_0_16_10_imag,
  output     [15:0]   io_coef_out_payload_0_16_11_real,
  output     [15:0]   io_coef_out_payload_0_16_11_imag,
  output     [15:0]   io_coef_out_payload_0_16_12_real,
  output     [15:0]   io_coef_out_payload_0_16_12_imag,
  output     [15:0]   io_coef_out_payload_0_16_13_real,
  output     [15:0]   io_coef_out_payload_0_16_13_imag,
  output     [15:0]   io_coef_out_payload_0_16_14_real,
  output     [15:0]   io_coef_out_payload_0_16_14_imag,
  output     [15:0]   io_coef_out_payload_0_16_15_real,
  output     [15:0]   io_coef_out_payload_0_16_15_imag,
  output     [15:0]   io_coef_out_payload_0_16_16_real,
  output     [15:0]   io_coef_out_payload_0_16_16_imag,
  output     [15:0]   io_coef_out_payload_0_16_17_real,
  output     [15:0]   io_coef_out_payload_0_16_17_imag,
  output     [15:0]   io_coef_out_payload_0_16_18_real,
  output     [15:0]   io_coef_out_payload_0_16_18_imag,
  output     [15:0]   io_coef_out_payload_0_16_19_real,
  output     [15:0]   io_coef_out_payload_0_16_19_imag,
  output     [15:0]   io_coef_out_payload_0_16_20_real,
  output     [15:0]   io_coef_out_payload_0_16_20_imag,
  output     [15:0]   io_coef_out_payload_0_16_21_real,
  output     [15:0]   io_coef_out_payload_0_16_21_imag,
  output     [15:0]   io_coef_out_payload_0_16_22_real,
  output     [15:0]   io_coef_out_payload_0_16_22_imag,
  output     [15:0]   io_coef_out_payload_0_16_23_real,
  output     [15:0]   io_coef_out_payload_0_16_23_imag,
  output     [15:0]   io_coef_out_payload_0_16_24_real,
  output     [15:0]   io_coef_out_payload_0_16_24_imag,
  output     [15:0]   io_coef_out_payload_0_16_25_real,
  output     [15:0]   io_coef_out_payload_0_16_25_imag,
  output     [15:0]   io_coef_out_payload_0_16_26_real,
  output     [15:0]   io_coef_out_payload_0_16_26_imag,
  output     [15:0]   io_coef_out_payload_0_16_27_real,
  output     [15:0]   io_coef_out_payload_0_16_27_imag,
  output     [15:0]   io_coef_out_payload_0_16_28_real,
  output     [15:0]   io_coef_out_payload_0_16_28_imag,
  output     [15:0]   io_coef_out_payload_0_16_29_real,
  output     [15:0]   io_coef_out_payload_0_16_29_imag,
  output     [15:0]   io_coef_out_payload_0_16_30_real,
  output     [15:0]   io_coef_out_payload_0_16_30_imag,
  output     [15:0]   io_coef_out_payload_0_16_31_real,
  output     [15:0]   io_coef_out_payload_0_16_31_imag,
  output     [15:0]   io_coef_out_payload_0_16_32_real,
  output     [15:0]   io_coef_out_payload_0_16_32_imag,
  output     [15:0]   io_coef_out_payload_0_16_33_real,
  output     [15:0]   io_coef_out_payload_0_16_33_imag,
  output     [15:0]   io_coef_out_payload_0_16_34_real,
  output     [15:0]   io_coef_out_payload_0_16_34_imag,
  output     [15:0]   io_coef_out_payload_0_16_35_real,
  output     [15:0]   io_coef_out_payload_0_16_35_imag,
  output     [15:0]   io_coef_out_payload_0_16_36_real,
  output     [15:0]   io_coef_out_payload_0_16_36_imag,
  output     [15:0]   io_coef_out_payload_0_16_37_real,
  output     [15:0]   io_coef_out_payload_0_16_37_imag,
  output     [15:0]   io_coef_out_payload_0_16_38_real,
  output     [15:0]   io_coef_out_payload_0_16_38_imag,
  output     [15:0]   io_coef_out_payload_0_16_39_real,
  output     [15:0]   io_coef_out_payload_0_16_39_imag,
  output     [15:0]   io_coef_out_payload_0_16_40_real,
  output     [15:0]   io_coef_out_payload_0_16_40_imag,
  output     [15:0]   io_coef_out_payload_0_16_41_real,
  output     [15:0]   io_coef_out_payload_0_16_41_imag,
  output     [15:0]   io_coef_out_payload_0_16_42_real,
  output     [15:0]   io_coef_out_payload_0_16_42_imag,
  output     [15:0]   io_coef_out_payload_0_16_43_real,
  output     [15:0]   io_coef_out_payload_0_16_43_imag,
  output     [15:0]   io_coef_out_payload_0_16_44_real,
  output     [15:0]   io_coef_out_payload_0_16_44_imag,
  output     [15:0]   io_coef_out_payload_0_16_45_real,
  output     [15:0]   io_coef_out_payload_0_16_45_imag,
  output     [15:0]   io_coef_out_payload_0_16_46_real,
  output     [15:0]   io_coef_out_payload_0_16_46_imag,
  output     [15:0]   io_coef_out_payload_0_16_47_real,
  output     [15:0]   io_coef_out_payload_0_16_47_imag,
  output     [15:0]   io_coef_out_payload_0_16_48_real,
  output     [15:0]   io_coef_out_payload_0_16_48_imag,
  output     [15:0]   io_coef_out_payload_0_16_49_real,
  output     [15:0]   io_coef_out_payload_0_16_49_imag,
  output     [15:0]   io_coef_out_payload_0_17_0_real,
  output     [15:0]   io_coef_out_payload_0_17_0_imag,
  output     [15:0]   io_coef_out_payload_0_17_1_real,
  output     [15:0]   io_coef_out_payload_0_17_1_imag,
  output     [15:0]   io_coef_out_payload_0_17_2_real,
  output     [15:0]   io_coef_out_payload_0_17_2_imag,
  output     [15:0]   io_coef_out_payload_0_17_3_real,
  output     [15:0]   io_coef_out_payload_0_17_3_imag,
  output     [15:0]   io_coef_out_payload_0_17_4_real,
  output     [15:0]   io_coef_out_payload_0_17_4_imag,
  output     [15:0]   io_coef_out_payload_0_17_5_real,
  output     [15:0]   io_coef_out_payload_0_17_5_imag,
  output     [15:0]   io_coef_out_payload_0_17_6_real,
  output     [15:0]   io_coef_out_payload_0_17_6_imag,
  output     [15:0]   io_coef_out_payload_0_17_7_real,
  output     [15:0]   io_coef_out_payload_0_17_7_imag,
  output     [15:0]   io_coef_out_payload_0_17_8_real,
  output     [15:0]   io_coef_out_payload_0_17_8_imag,
  output     [15:0]   io_coef_out_payload_0_17_9_real,
  output     [15:0]   io_coef_out_payload_0_17_9_imag,
  output     [15:0]   io_coef_out_payload_0_17_10_real,
  output     [15:0]   io_coef_out_payload_0_17_10_imag,
  output     [15:0]   io_coef_out_payload_0_17_11_real,
  output     [15:0]   io_coef_out_payload_0_17_11_imag,
  output     [15:0]   io_coef_out_payload_0_17_12_real,
  output     [15:0]   io_coef_out_payload_0_17_12_imag,
  output     [15:0]   io_coef_out_payload_0_17_13_real,
  output     [15:0]   io_coef_out_payload_0_17_13_imag,
  output     [15:0]   io_coef_out_payload_0_17_14_real,
  output     [15:0]   io_coef_out_payload_0_17_14_imag,
  output     [15:0]   io_coef_out_payload_0_17_15_real,
  output     [15:0]   io_coef_out_payload_0_17_15_imag,
  output     [15:0]   io_coef_out_payload_0_17_16_real,
  output     [15:0]   io_coef_out_payload_0_17_16_imag,
  output     [15:0]   io_coef_out_payload_0_17_17_real,
  output     [15:0]   io_coef_out_payload_0_17_17_imag,
  output     [15:0]   io_coef_out_payload_0_17_18_real,
  output     [15:0]   io_coef_out_payload_0_17_18_imag,
  output     [15:0]   io_coef_out_payload_0_17_19_real,
  output     [15:0]   io_coef_out_payload_0_17_19_imag,
  output     [15:0]   io_coef_out_payload_0_17_20_real,
  output     [15:0]   io_coef_out_payload_0_17_20_imag,
  output     [15:0]   io_coef_out_payload_0_17_21_real,
  output     [15:0]   io_coef_out_payload_0_17_21_imag,
  output     [15:0]   io_coef_out_payload_0_17_22_real,
  output     [15:0]   io_coef_out_payload_0_17_22_imag,
  output     [15:0]   io_coef_out_payload_0_17_23_real,
  output     [15:0]   io_coef_out_payload_0_17_23_imag,
  output     [15:0]   io_coef_out_payload_0_17_24_real,
  output     [15:0]   io_coef_out_payload_0_17_24_imag,
  output     [15:0]   io_coef_out_payload_0_17_25_real,
  output     [15:0]   io_coef_out_payload_0_17_25_imag,
  output     [15:0]   io_coef_out_payload_0_17_26_real,
  output     [15:0]   io_coef_out_payload_0_17_26_imag,
  output     [15:0]   io_coef_out_payload_0_17_27_real,
  output     [15:0]   io_coef_out_payload_0_17_27_imag,
  output     [15:0]   io_coef_out_payload_0_17_28_real,
  output     [15:0]   io_coef_out_payload_0_17_28_imag,
  output     [15:0]   io_coef_out_payload_0_17_29_real,
  output     [15:0]   io_coef_out_payload_0_17_29_imag,
  output     [15:0]   io_coef_out_payload_0_17_30_real,
  output     [15:0]   io_coef_out_payload_0_17_30_imag,
  output     [15:0]   io_coef_out_payload_0_17_31_real,
  output     [15:0]   io_coef_out_payload_0_17_31_imag,
  output     [15:0]   io_coef_out_payload_0_17_32_real,
  output     [15:0]   io_coef_out_payload_0_17_32_imag,
  output     [15:0]   io_coef_out_payload_0_17_33_real,
  output     [15:0]   io_coef_out_payload_0_17_33_imag,
  output     [15:0]   io_coef_out_payload_0_17_34_real,
  output     [15:0]   io_coef_out_payload_0_17_34_imag,
  output     [15:0]   io_coef_out_payload_0_17_35_real,
  output     [15:0]   io_coef_out_payload_0_17_35_imag,
  output     [15:0]   io_coef_out_payload_0_17_36_real,
  output     [15:0]   io_coef_out_payload_0_17_36_imag,
  output     [15:0]   io_coef_out_payload_0_17_37_real,
  output     [15:0]   io_coef_out_payload_0_17_37_imag,
  output     [15:0]   io_coef_out_payload_0_17_38_real,
  output     [15:0]   io_coef_out_payload_0_17_38_imag,
  output     [15:0]   io_coef_out_payload_0_17_39_real,
  output     [15:0]   io_coef_out_payload_0_17_39_imag,
  output     [15:0]   io_coef_out_payload_0_17_40_real,
  output     [15:0]   io_coef_out_payload_0_17_40_imag,
  output     [15:0]   io_coef_out_payload_0_17_41_real,
  output     [15:0]   io_coef_out_payload_0_17_41_imag,
  output     [15:0]   io_coef_out_payload_0_17_42_real,
  output     [15:0]   io_coef_out_payload_0_17_42_imag,
  output     [15:0]   io_coef_out_payload_0_17_43_real,
  output     [15:0]   io_coef_out_payload_0_17_43_imag,
  output     [15:0]   io_coef_out_payload_0_17_44_real,
  output     [15:0]   io_coef_out_payload_0_17_44_imag,
  output     [15:0]   io_coef_out_payload_0_17_45_real,
  output     [15:0]   io_coef_out_payload_0_17_45_imag,
  output     [15:0]   io_coef_out_payload_0_17_46_real,
  output     [15:0]   io_coef_out_payload_0_17_46_imag,
  output     [15:0]   io_coef_out_payload_0_17_47_real,
  output     [15:0]   io_coef_out_payload_0_17_47_imag,
  output     [15:0]   io_coef_out_payload_0_17_48_real,
  output     [15:0]   io_coef_out_payload_0_17_48_imag,
  output     [15:0]   io_coef_out_payload_0_17_49_real,
  output     [15:0]   io_coef_out_payload_0_17_49_imag,
  output     [15:0]   io_coef_out_payload_0_18_0_real,
  output     [15:0]   io_coef_out_payload_0_18_0_imag,
  output     [15:0]   io_coef_out_payload_0_18_1_real,
  output     [15:0]   io_coef_out_payload_0_18_1_imag,
  output     [15:0]   io_coef_out_payload_0_18_2_real,
  output     [15:0]   io_coef_out_payload_0_18_2_imag,
  output     [15:0]   io_coef_out_payload_0_18_3_real,
  output     [15:0]   io_coef_out_payload_0_18_3_imag,
  output     [15:0]   io_coef_out_payload_0_18_4_real,
  output     [15:0]   io_coef_out_payload_0_18_4_imag,
  output     [15:0]   io_coef_out_payload_0_18_5_real,
  output     [15:0]   io_coef_out_payload_0_18_5_imag,
  output     [15:0]   io_coef_out_payload_0_18_6_real,
  output     [15:0]   io_coef_out_payload_0_18_6_imag,
  output     [15:0]   io_coef_out_payload_0_18_7_real,
  output     [15:0]   io_coef_out_payload_0_18_7_imag,
  output     [15:0]   io_coef_out_payload_0_18_8_real,
  output     [15:0]   io_coef_out_payload_0_18_8_imag,
  output     [15:0]   io_coef_out_payload_0_18_9_real,
  output     [15:0]   io_coef_out_payload_0_18_9_imag,
  output     [15:0]   io_coef_out_payload_0_18_10_real,
  output     [15:0]   io_coef_out_payload_0_18_10_imag,
  output     [15:0]   io_coef_out_payload_0_18_11_real,
  output     [15:0]   io_coef_out_payload_0_18_11_imag,
  output     [15:0]   io_coef_out_payload_0_18_12_real,
  output     [15:0]   io_coef_out_payload_0_18_12_imag,
  output     [15:0]   io_coef_out_payload_0_18_13_real,
  output     [15:0]   io_coef_out_payload_0_18_13_imag,
  output     [15:0]   io_coef_out_payload_0_18_14_real,
  output     [15:0]   io_coef_out_payload_0_18_14_imag,
  output     [15:0]   io_coef_out_payload_0_18_15_real,
  output     [15:0]   io_coef_out_payload_0_18_15_imag,
  output     [15:0]   io_coef_out_payload_0_18_16_real,
  output     [15:0]   io_coef_out_payload_0_18_16_imag,
  output     [15:0]   io_coef_out_payload_0_18_17_real,
  output     [15:0]   io_coef_out_payload_0_18_17_imag,
  output     [15:0]   io_coef_out_payload_0_18_18_real,
  output     [15:0]   io_coef_out_payload_0_18_18_imag,
  output     [15:0]   io_coef_out_payload_0_18_19_real,
  output     [15:0]   io_coef_out_payload_0_18_19_imag,
  output     [15:0]   io_coef_out_payload_0_18_20_real,
  output     [15:0]   io_coef_out_payload_0_18_20_imag,
  output     [15:0]   io_coef_out_payload_0_18_21_real,
  output     [15:0]   io_coef_out_payload_0_18_21_imag,
  output     [15:0]   io_coef_out_payload_0_18_22_real,
  output     [15:0]   io_coef_out_payload_0_18_22_imag,
  output     [15:0]   io_coef_out_payload_0_18_23_real,
  output     [15:0]   io_coef_out_payload_0_18_23_imag,
  output     [15:0]   io_coef_out_payload_0_18_24_real,
  output     [15:0]   io_coef_out_payload_0_18_24_imag,
  output     [15:0]   io_coef_out_payload_0_18_25_real,
  output     [15:0]   io_coef_out_payload_0_18_25_imag,
  output     [15:0]   io_coef_out_payload_0_18_26_real,
  output     [15:0]   io_coef_out_payload_0_18_26_imag,
  output     [15:0]   io_coef_out_payload_0_18_27_real,
  output     [15:0]   io_coef_out_payload_0_18_27_imag,
  output     [15:0]   io_coef_out_payload_0_18_28_real,
  output     [15:0]   io_coef_out_payload_0_18_28_imag,
  output     [15:0]   io_coef_out_payload_0_18_29_real,
  output     [15:0]   io_coef_out_payload_0_18_29_imag,
  output     [15:0]   io_coef_out_payload_0_18_30_real,
  output     [15:0]   io_coef_out_payload_0_18_30_imag,
  output     [15:0]   io_coef_out_payload_0_18_31_real,
  output     [15:0]   io_coef_out_payload_0_18_31_imag,
  output     [15:0]   io_coef_out_payload_0_18_32_real,
  output     [15:0]   io_coef_out_payload_0_18_32_imag,
  output     [15:0]   io_coef_out_payload_0_18_33_real,
  output     [15:0]   io_coef_out_payload_0_18_33_imag,
  output     [15:0]   io_coef_out_payload_0_18_34_real,
  output     [15:0]   io_coef_out_payload_0_18_34_imag,
  output     [15:0]   io_coef_out_payload_0_18_35_real,
  output     [15:0]   io_coef_out_payload_0_18_35_imag,
  output     [15:0]   io_coef_out_payload_0_18_36_real,
  output     [15:0]   io_coef_out_payload_0_18_36_imag,
  output     [15:0]   io_coef_out_payload_0_18_37_real,
  output     [15:0]   io_coef_out_payload_0_18_37_imag,
  output     [15:0]   io_coef_out_payload_0_18_38_real,
  output     [15:0]   io_coef_out_payload_0_18_38_imag,
  output     [15:0]   io_coef_out_payload_0_18_39_real,
  output     [15:0]   io_coef_out_payload_0_18_39_imag,
  output     [15:0]   io_coef_out_payload_0_18_40_real,
  output     [15:0]   io_coef_out_payload_0_18_40_imag,
  output     [15:0]   io_coef_out_payload_0_18_41_real,
  output     [15:0]   io_coef_out_payload_0_18_41_imag,
  output     [15:0]   io_coef_out_payload_0_18_42_real,
  output     [15:0]   io_coef_out_payload_0_18_42_imag,
  output     [15:0]   io_coef_out_payload_0_18_43_real,
  output     [15:0]   io_coef_out_payload_0_18_43_imag,
  output     [15:0]   io_coef_out_payload_0_18_44_real,
  output     [15:0]   io_coef_out_payload_0_18_44_imag,
  output     [15:0]   io_coef_out_payload_0_18_45_real,
  output     [15:0]   io_coef_out_payload_0_18_45_imag,
  output     [15:0]   io_coef_out_payload_0_18_46_real,
  output     [15:0]   io_coef_out_payload_0_18_46_imag,
  output     [15:0]   io_coef_out_payload_0_18_47_real,
  output     [15:0]   io_coef_out_payload_0_18_47_imag,
  output     [15:0]   io_coef_out_payload_0_18_48_real,
  output     [15:0]   io_coef_out_payload_0_18_48_imag,
  output     [15:0]   io_coef_out_payload_0_18_49_real,
  output     [15:0]   io_coef_out_payload_0_18_49_imag,
  output     [15:0]   io_coef_out_payload_0_19_0_real,
  output     [15:0]   io_coef_out_payload_0_19_0_imag,
  output     [15:0]   io_coef_out_payload_0_19_1_real,
  output     [15:0]   io_coef_out_payload_0_19_1_imag,
  output     [15:0]   io_coef_out_payload_0_19_2_real,
  output     [15:0]   io_coef_out_payload_0_19_2_imag,
  output     [15:0]   io_coef_out_payload_0_19_3_real,
  output     [15:0]   io_coef_out_payload_0_19_3_imag,
  output     [15:0]   io_coef_out_payload_0_19_4_real,
  output     [15:0]   io_coef_out_payload_0_19_4_imag,
  output     [15:0]   io_coef_out_payload_0_19_5_real,
  output     [15:0]   io_coef_out_payload_0_19_5_imag,
  output     [15:0]   io_coef_out_payload_0_19_6_real,
  output     [15:0]   io_coef_out_payload_0_19_6_imag,
  output     [15:0]   io_coef_out_payload_0_19_7_real,
  output     [15:0]   io_coef_out_payload_0_19_7_imag,
  output     [15:0]   io_coef_out_payload_0_19_8_real,
  output     [15:0]   io_coef_out_payload_0_19_8_imag,
  output     [15:0]   io_coef_out_payload_0_19_9_real,
  output     [15:0]   io_coef_out_payload_0_19_9_imag,
  output     [15:0]   io_coef_out_payload_0_19_10_real,
  output     [15:0]   io_coef_out_payload_0_19_10_imag,
  output     [15:0]   io_coef_out_payload_0_19_11_real,
  output     [15:0]   io_coef_out_payload_0_19_11_imag,
  output     [15:0]   io_coef_out_payload_0_19_12_real,
  output     [15:0]   io_coef_out_payload_0_19_12_imag,
  output     [15:0]   io_coef_out_payload_0_19_13_real,
  output     [15:0]   io_coef_out_payload_0_19_13_imag,
  output     [15:0]   io_coef_out_payload_0_19_14_real,
  output     [15:0]   io_coef_out_payload_0_19_14_imag,
  output     [15:0]   io_coef_out_payload_0_19_15_real,
  output     [15:0]   io_coef_out_payload_0_19_15_imag,
  output     [15:0]   io_coef_out_payload_0_19_16_real,
  output     [15:0]   io_coef_out_payload_0_19_16_imag,
  output     [15:0]   io_coef_out_payload_0_19_17_real,
  output     [15:0]   io_coef_out_payload_0_19_17_imag,
  output     [15:0]   io_coef_out_payload_0_19_18_real,
  output     [15:0]   io_coef_out_payload_0_19_18_imag,
  output     [15:0]   io_coef_out_payload_0_19_19_real,
  output     [15:0]   io_coef_out_payload_0_19_19_imag,
  output     [15:0]   io_coef_out_payload_0_19_20_real,
  output     [15:0]   io_coef_out_payload_0_19_20_imag,
  output     [15:0]   io_coef_out_payload_0_19_21_real,
  output     [15:0]   io_coef_out_payload_0_19_21_imag,
  output     [15:0]   io_coef_out_payload_0_19_22_real,
  output     [15:0]   io_coef_out_payload_0_19_22_imag,
  output     [15:0]   io_coef_out_payload_0_19_23_real,
  output     [15:0]   io_coef_out_payload_0_19_23_imag,
  output     [15:0]   io_coef_out_payload_0_19_24_real,
  output     [15:0]   io_coef_out_payload_0_19_24_imag,
  output     [15:0]   io_coef_out_payload_0_19_25_real,
  output     [15:0]   io_coef_out_payload_0_19_25_imag,
  output     [15:0]   io_coef_out_payload_0_19_26_real,
  output     [15:0]   io_coef_out_payload_0_19_26_imag,
  output     [15:0]   io_coef_out_payload_0_19_27_real,
  output     [15:0]   io_coef_out_payload_0_19_27_imag,
  output     [15:0]   io_coef_out_payload_0_19_28_real,
  output     [15:0]   io_coef_out_payload_0_19_28_imag,
  output     [15:0]   io_coef_out_payload_0_19_29_real,
  output     [15:0]   io_coef_out_payload_0_19_29_imag,
  output     [15:0]   io_coef_out_payload_0_19_30_real,
  output     [15:0]   io_coef_out_payload_0_19_30_imag,
  output     [15:0]   io_coef_out_payload_0_19_31_real,
  output     [15:0]   io_coef_out_payload_0_19_31_imag,
  output     [15:0]   io_coef_out_payload_0_19_32_real,
  output     [15:0]   io_coef_out_payload_0_19_32_imag,
  output     [15:0]   io_coef_out_payload_0_19_33_real,
  output     [15:0]   io_coef_out_payload_0_19_33_imag,
  output     [15:0]   io_coef_out_payload_0_19_34_real,
  output     [15:0]   io_coef_out_payload_0_19_34_imag,
  output     [15:0]   io_coef_out_payload_0_19_35_real,
  output     [15:0]   io_coef_out_payload_0_19_35_imag,
  output     [15:0]   io_coef_out_payload_0_19_36_real,
  output     [15:0]   io_coef_out_payload_0_19_36_imag,
  output     [15:0]   io_coef_out_payload_0_19_37_real,
  output     [15:0]   io_coef_out_payload_0_19_37_imag,
  output     [15:0]   io_coef_out_payload_0_19_38_real,
  output     [15:0]   io_coef_out_payload_0_19_38_imag,
  output     [15:0]   io_coef_out_payload_0_19_39_real,
  output     [15:0]   io_coef_out_payload_0_19_39_imag,
  output     [15:0]   io_coef_out_payload_0_19_40_real,
  output     [15:0]   io_coef_out_payload_0_19_40_imag,
  output     [15:0]   io_coef_out_payload_0_19_41_real,
  output     [15:0]   io_coef_out_payload_0_19_41_imag,
  output     [15:0]   io_coef_out_payload_0_19_42_real,
  output     [15:0]   io_coef_out_payload_0_19_42_imag,
  output     [15:0]   io_coef_out_payload_0_19_43_real,
  output     [15:0]   io_coef_out_payload_0_19_43_imag,
  output     [15:0]   io_coef_out_payload_0_19_44_real,
  output     [15:0]   io_coef_out_payload_0_19_44_imag,
  output     [15:0]   io_coef_out_payload_0_19_45_real,
  output     [15:0]   io_coef_out_payload_0_19_45_imag,
  output     [15:0]   io_coef_out_payload_0_19_46_real,
  output     [15:0]   io_coef_out_payload_0_19_46_imag,
  output     [15:0]   io_coef_out_payload_0_19_47_real,
  output     [15:0]   io_coef_out_payload_0_19_47_imag,
  output     [15:0]   io_coef_out_payload_0_19_48_real,
  output     [15:0]   io_coef_out_payload_0_19_48_imag,
  output     [15:0]   io_coef_out_payload_0_19_49_real,
  output     [15:0]   io_coef_out_payload_0_19_49_imag,
  output     [15:0]   io_coef_out_payload_0_20_0_real,
  output     [15:0]   io_coef_out_payload_0_20_0_imag,
  output     [15:0]   io_coef_out_payload_0_20_1_real,
  output     [15:0]   io_coef_out_payload_0_20_1_imag,
  output     [15:0]   io_coef_out_payload_0_20_2_real,
  output     [15:0]   io_coef_out_payload_0_20_2_imag,
  output     [15:0]   io_coef_out_payload_0_20_3_real,
  output     [15:0]   io_coef_out_payload_0_20_3_imag,
  output     [15:0]   io_coef_out_payload_0_20_4_real,
  output     [15:0]   io_coef_out_payload_0_20_4_imag,
  output     [15:0]   io_coef_out_payload_0_20_5_real,
  output     [15:0]   io_coef_out_payload_0_20_5_imag,
  output     [15:0]   io_coef_out_payload_0_20_6_real,
  output     [15:0]   io_coef_out_payload_0_20_6_imag,
  output     [15:0]   io_coef_out_payload_0_20_7_real,
  output     [15:0]   io_coef_out_payload_0_20_7_imag,
  output     [15:0]   io_coef_out_payload_0_20_8_real,
  output     [15:0]   io_coef_out_payload_0_20_8_imag,
  output     [15:0]   io_coef_out_payload_0_20_9_real,
  output     [15:0]   io_coef_out_payload_0_20_9_imag,
  output     [15:0]   io_coef_out_payload_0_20_10_real,
  output     [15:0]   io_coef_out_payload_0_20_10_imag,
  output     [15:0]   io_coef_out_payload_0_20_11_real,
  output     [15:0]   io_coef_out_payload_0_20_11_imag,
  output     [15:0]   io_coef_out_payload_0_20_12_real,
  output     [15:0]   io_coef_out_payload_0_20_12_imag,
  output     [15:0]   io_coef_out_payload_0_20_13_real,
  output     [15:0]   io_coef_out_payload_0_20_13_imag,
  output     [15:0]   io_coef_out_payload_0_20_14_real,
  output     [15:0]   io_coef_out_payload_0_20_14_imag,
  output     [15:0]   io_coef_out_payload_0_20_15_real,
  output     [15:0]   io_coef_out_payload_0_20_15_imag,
  output     [15:0]   io_coef_out_payload_0_20_16_real,
  output     [15:0]   io_coef_out_payload_0_20_16_imag,
  output     [15:0]   io_coef_out_payload_0_20_17_real,
  output     [15:0]   io_coef_out_payload_0_20_17_imag,
  output     [15:0]   io_coef_out_payload_0_20_18_real,
  output     [15:0]   io_coef_out_payload_0_20_18_imag,
  output     [15:0]   io_coef_out_payload_0_20_19_real,
  output     [15:0]   io_coef_out_payload_0_20_19_imag,
  output     [15:0]   io_coef_out_payload_0_20_20_real,
  output     [15:0]   io_coef_out_payload_0_20_20_imag,
  output     [15:0]   io_coef_out_payload_0_20_21_real,
  output     [15:0]   io_coef_out_payload_0_20_21_imag,
  output     [15:0]   io_coef_out_payload_0_20_22_real,
  output     [15:0]   io_coef_out_payload_0_20_22_imag,
  output     [15:0]   io_coef_out_payload_0_20_23_real,
  output     [15:0]   io_coef_out_payload_0_20_23_imag,
  output     [15:0]   io_coef_out_payload_0_20_24_real,
  output     [15:0]   io_coef_out_payload_0_20_24_imag,
  output     [15:0]   io_coef_out_payload_0_20_25_real,
  output     [15:0]   io_coef_out_payload_0_20_25_imag,
  output     [15:0]   io_coef_out_payload_0_20_26_real,
  output     [15:0]   io_coef_out_payload_0_20_26_imag,
  output     [15:0]   io_coef_out_payload_0_20_27_real,
  output     [15:0]   io_coef_out_payload_0_20_27_imag,
  output     [15:0]   io_coef_out_payload_0_20_28_real,
  output     [15:0]   io_coef_out_payload_0_20_28_imag,
  output     [15:0]   io_coef_out_payload_0_20_29_real,
  output     [15:0]   io_coef_out_payload_0_20_29_imag,
  output     [15:0]   io_coef_out_payload_0_20_30_real,
  output     [15:0]   io_coef_out_payload_0_20_30_imag,
  output     [15:0]   io_coef_out_payload_0_20_31_real,
  output     [15:0]   io_coef_out_payload_0_20_31_imag,
  output     [15:0]   io_coef_out_payload_0_20_32_real,
  output     [15:0]   io_coef_out_payload_0_20_32_imag,
  output     [15:0]   io_coef_out_payload_0_20_33_real,
  output     [15:0]   io_coef_out_payload_0_20_33_imag,
  output     [15:0]   io_coef_out_payload_0_20_34_real,
  output     [15:0]   io_coef_out_payload_0_20_34_imag,
  output     [15:0]   io_coef_out_payload_0_20_35_real,
  output     [15:0]   io_coef_out_payload_0_20_35_imag,
  output     [15:0]   io_coef_out_payload_0_20_36_real,
  output     [15:0]   io_coef_out_payload_0_20_36_imag,
  output     [15:0]   io_coef_out_payload_0_20_37_real,
  output     [15:0]   io_coef_out_payload_0_20_37_imag,
  output     [15:0]   io_coef_out_payload_0_20_38_real,
  output     [15:0]   io_coef_out_payload_0_20_38_imag,
  output     [15:0]   io_coef_out_payload_0_20_39_real,
  output     [15:0]   io_coef_out_payload_0_20_39_imag,
  output     [15:0]   io_coef_out_payload_0_20_40_real,
  output     [15:0]   io_coef_out_payload_0_20_40_imag,
  output     [15:0]   io_coef_out_payload_0_20_41_real,
  output     [15:0]   io_coef_out_payload_0_20_41_imag,
  output     [15:0]   io_coef_out_payload_0_20_42_real,
  output     [15:0]   io_coef_out_payload_0_20_42_imag,
  output     [15:0]   io_coef_out_payload_0_20_43_real,
  output     [15:0]   io_coef_out_payload_0_20_43_imag,
  output     [15:0]   io_coef_out_payload_0_20_44_real,
  output     [15:0]   io_coef_out_payload_0_20_44_imag,
  output     [15:0]   io_coef_out_payload_0_20_45_real,
  output     [15:0]   io_coef_out_payload_0_20_45_imag,
  output     [15:0]   io_coef_out_payload_0_20_46_real,
  output     [15:0]   io_coef_out_payload_0_20_46_imag,
  output     [15:0]   io_coef_out_payload_0_20_47_real,
  output     [15:0]   io_coef_out_payload_0_20_47_imag,
  output     [15:0]   io_coef_out_payload_0_20_48_real,
  output     [15:0]   io_coef_out_payload_0_20_48_imag,
  output     [15:0]   io_coef_out_payload_0_20_49_real,
  output     [15:0]   io_coef_out_payload_0_20_49_imag,
  output     [15:0]   io_coef_out_payload_0_21_0_real,
  output     [15:0]   io_coef_out_payload_0_21_0_imag,
  output     [15:0]   io_coef_out_payload_0_21_1_real,
  output     [15:0]   io_coef_out_payload_0_21_1_imag,
  output     [15:0]   io_coef_out_payload_0_21_2_real,
  output     [15:0]   io_coef_out_payload_0_21_2_imag,
  output     [15:0]   io_coef_out_payload_0_21_3_real,
  output     [15:0]   io_coef_out_payload_0_21_3_imag,
  output     [15:0]   io_coef_out_payload_0_21_4_real,
  output     [15:0]   io_coef_out_payload_0_21_4_imag,
  output     [15:0]   io_coef_out_payload_0_21_5_real,
  output     [15:0]   io_coef_out_payload_0_21_5_imag,
  output     [15:0]   io_coef_out_payload_0_21_6_real,
  output     [15:0]   io_coef_out_payload_0_21_6_imag,
  output     [15:0]   io_coef_out_payload_0_21_7_real,
  output     [15:0]   io_coef_out_payload_0_21_7_imag,
  output     [15:0]   io_coef_out_payload_0_21_8_real,
  output     [15:0]   io_coef_out_payload_0_21_8_imag,
  output     [15:0]   io_coef_out_payload_0_21_9_real,
  output     [15:0]   io_coef_out_payload_0_21_9_imag,
  output     [15:0]   io_coef_out_payload_0_21_10_real,
  output     [15:0]   io_coef_out_payload_0_21_10_imag,
  output     [15:0]   io_coef_out_payload_0_21_11_real,
  output     [15:0]   io_coef_out_payload_0_21_11_imag,
  output     [15:0]   io_coef_out_payload_0_21_12_real,
  output     [15:0]   io_coef_out_payload_0_21_12_imag,
  output     [15:0]   io_coef_out_payload_0_21_13_real,
  output     [15:0]   io_coef_out_payload_0_21_13_imag,
  output     [15:0]   io_coef_out_payload_0_21_14_real,
  output     [15:0]   io_coef_out_payload_0_21_14_imag,
  output     [15:0]   io_coef_out_payload_0_21_15_real,
  output     [15:0]   io_coef_out_payload_0_21_15_imag,
  output     [15:0]   io_coef_out_payload_0_21_16_real,
  output     [15:0]   io_coef_out_payload_0_21_16_imag,
  output     [15:0]   io_coef_out_payload_0_21_17_real,
  output     [15:0]   io_coef_out_payload_0_21_17_imag,
  output     [15:0]   io_coef_out_payload_0_21_18_real,
  output     [15:0]   io_coef_out_payload_0_21_18_imag,
  output     [15:0]   io_coef_out_payload_0_21_19_real,
  output     [15:0]   io_coef_out_payload_0_21_19_imag,
  output     [15:0]   io_coef_out_payload_0_21_20_real,
  output     [15:0]   io_coef_out_payload_0_21_20_imag,
  output     [15:0]   io_coef_out_payload_0_21_21_real,
  output     [15:0]   io_coef_out_payload_0_21_21_imag,
  output     [15:0]   io_coef_out_payload_0_21_22_real,
  output     [15:0]   io_coef_out_payload_0_21_22_imag,
  output     [15:0]   io_coef_out_payload_0_21_23_real,
  output     [15:0]   io_coef_out_payload_0_21_23_imag,
  output     [15:0]   io_coef_out_payload_0_21_24_real,
  output     [15:0]   io_coef_out_payload_0_21_24_imag,
  output     [15:0]   io_coef_out_payload_0_21_25_real,
  output     [15:0]   io_coef_out_payload_0_21_25_imag,
  output     [15:0]   io_coef_out_payload_0_21_26_real,
  output     [15:0]   io_coef_out_payload_0_21_26_imag,
  output     [15:0]   io_coef_out_payload_0_21_27_real,
  output     [15:0]   io_coef_out_payload_0_21_27_imag,
  output     [15:0]   io_coef_out_payload_0_21_28_real,
  output     [15:0]   io_coef_out_payload_0_21_28_imag,
  output     [15:0]   io_coef_out_payload_0_21_29_real,
  output     [15:0]   io_coef_out_payload_0_21_29_imag,
  output     [15:0]   io_coef_out_payload_0_21_30_real,
  output     [15:0]   io_coef_out_payload_0_21_30_imag,
  output     [15:0]   io_coef_out_payload_0_21_31_real,
  output     [15:0]   io_coef_out_payload_0_21_31_imag,
  output     [15:0]   io_coef_out_payload_0_21_32_real,
  output     [15:0]   io_coef_out_payload_0_21_32_imag,
  output     [15:0]   io_coef_out_payload_0_21_33_real,
  output     [15:0]   io_coef_out_payload_0_21_33_imag,
  output     [15:0]   io_coef_out_payload_0_21_34_real,
  output     [15:0]   io_coef_out_payload_0_21_34_imag,
  output     [15:0]   io_coef_out_payload_0_21_35_real,
  output     [15:0]   io_coef_out_payload_0_21_35_imag,
  output     [15:0]   io_coef_out_payload_0_21_36_real,
  output     [15:0]   io_coef_out_payload_0_21_36_imag,
  output     [15:0]   io_coef_out_payload_0_21_37_real,
  output     [15:0]   io_coef_out_payload_0_21_37_imag,
  output     [15:0]   io_coef_out_payload_0_21_38_real,
  output     [15:0]   io_coef_out_payload_0_21_38_imag,
  output     [15:0]   io_coef_out_payload_0_21_39_real,
  output     [15:0]   io_coef_out_payload_0_21_39_imag,
  output     [15:0]   io_coef_out_payload_0_21_40_real,
  output     [15:0]   io_coef_out_payload_0_21_40_imag,
  output     [15:0]   io_coef_out_payload_0_21_41_real,
  output     [15:0]   io_coef_out_payload_0_21_41_imag,
  output     [15:0]   io_coef_out_payload_0_21_42_real,
  output     [15:0]   io_coef_out_payload_0_21_42_imag,
  output     [15:0]   io_coef_out_payload_0_21_43_real,
  output     [15:0]   io_coef_out_payload_0_21_43_imag,
  output     [15:0]   io_coef_out_payload_0_21_44_real,
  output     [15:0]   io_coef_out_payload_0_21_44_imag,
  output     [15:0]   io_coef_out_payload_0_21_45_real,
  output     [15:0]   io_coef_out_payload_0_21_45_imag,
  output     [15:0]   io_coef_out_payload_0_21_46_real,
  output     [15:0]   io_coef_out_payload_0_21_46_imag,
  output     [15:0]   io_coef_out_payload_0_21_47_real,
  output     [15:0]   io_coef_out_payload_0_21_47_imag,
  output     [15:0]   io_coef_out_payload_0_21_48_real,
  output     [15:0]   io_coef_out_payload_0_21_48_imag,
  output     [15:0]   io_coef_out_payload_0_21_49_real,
  output     [15:0]   io_coef_out_payload_0_21_49_imag,
  output     [15:0]   io_coef_out_payload_0_22_0_real,
  output     [15:0]   io_coef_out_payload_0_22_0_imag,
  output     [15:0]   io_coef_out_payload_0_22_1_real,
  output     [15:0]   io_coef_out_payload_0_22_1_imag,
  output     [15:0]   io_coef_out_payload_0_22_2_real,
  output     [15:0]   io_coef_out_payload_0_22_2_imag,
  output     [15:0]   io_coef_out_payload_0_22_3_real,
  output     [15:0]   io_coef_out_payload_0_22_3_imag,
  output     [15:0]   io_coef_out_payload_0_22_4_real,
  output     [15:0]   io_coef_out_payload_0_22_4_imag,
  output     [15:0]   io_coef_out_payload_0_22_5_real,
  output     [15:0]   io_coef_out_payload_0_22_5_imag,
  output     [15:0]   io_coef_out_payload_0_22_6_real,
  output     [15:0]   io_coef_out_payload_0_22_6_imag,
  output     [15:0]   io_coef_out_payload_0_22_7_real,
  output     [15:0]   io_coef_out_payload_0_22_7_imag,
  output     [15:0]   io_coef_out_payload_0_22_8_real,
  output     [15:0]   io_coef_out_payload_0_22_8_imag,
  output     [15:0]   io_coef_out_payload_0_22_9_real,
  output     [15:0]   io_coef_out_payload_0_22_9_imag,
  output     [15:0]   io_coef_out_payload_0_22_10_real,
  output     [15:0]   io_coef_out_payload_0_22_10_imag,
  output     [15:0]   io_coef_out_payload_0_22_11_real,
  output     [15:0]   io_coef_out_payload_0_22_11_imag,
  output     [15:0]   io_coef_out_payload_0_22_12_real,
  output     [15:0]   io_coef_out_payload_0_22_12_imag,
  output     [15:0]   io_coef_out_payload_0_22_13_real,
  output     [15:0]   io_coef_out_payload_0_22_13_imag,
  output     [15:0]   io_coef_out_payload_0_22_14_real,
  output     [15:0]   io_coef_out_payload_0_22_14_imag,
  output     [15:0]   io_coef_out_payload_0_22_15_real,
  output     [15:0]   io_coef_out_payload_0_22_15_imag,
  output     [15:0]   io_coef_out_payload_0_22_16_real,
  output     [15:0]   io_coef_out_payload_0_22_16_imag,
  output     [15:0]   io_coef_out_payload_0_22_17_real,
  output     [15:0]   io_coef_out_payload_0_22_17_imag,
  output     [15:0]   io_coef_out_payload_0_22_18_real,
  output     [15:0]   io_coef_out_payload_0_22_18_imag,
  output     [15:0]   io_coef_out_payload_0_22_19_real,
  output     [15:0]   io_coef_out_payload_0_22_19_imag,
  output     [15:0]   io_coef_out_payload_0_22_20_real,
  output     [15:0]   io_coef_out_payload_0_22_20_imag,
  output     [15:0]   io_coef_out_payload_0_22_21_real,
  output     [15:0]   io_coef_out_payload_0_22_21_imag,
  output     [15:0]   io_coef_out_payload_0_22_22_real,
  output     [15:0]   io_coef_out_payload_0_22_22_imag,
  output     [15:0]   io_coef_out_payload_0_22_23_real,
  output     [15:0]   io_coef_out_payload_0_22_23_imag,
  output     [15:0]   io_coef_out_payload_0_22_24_real,
  output     [15:0]   io_coef_out_payload_0_22_24_imag,
  output     [15:0]   io_coef_out_payload_0_22_25_real,
  output     [15:0]   io_coef_out_payload_0_22_25_imag,
  output     [15:0]   io_coef_out_payload_0_22_26_real,
  output     [15:0]   io_coef_out_payload_0_22_26_imag,
  output     [15:0]   io_coef_out_payload_0_22_27_real,
  output     [15:0]   io_coef_out_payload_0_22_27_imag,
  output     [15:0]   io_coef_out_payload_0_22_28_real,
  output     [15:0]   io_coef_out_payload_0_22_28_imag,
  output     [15:0]   io_coef_out_payload_0_22_29_real,
  output     [15:0]   io_coef_out_payload_0_22_29_imag,
  output     [15:0]   io_coef_out_payload_0_22_30_real,
  output     [15:0]   io_coef_out_payload_0_22_30_imag,
  output     [15:0]   io_coef_out_payload_0_22_31_real,
  output     [15:0]   io_coef_out_payload_0_22_31_imag,
  output     [15:0]   io_coef_out_payload_0_22_32_real,
  output     [15:0]   io_coef_out_payload_0_22_32_imag,
  output     [15:0]   io_coef_out_payload_0_22_33_real,
  output     [15:0]   io_coef_out_payload_0_22_33_imag,
  output     [15:0]   io_coef_out_payload_0_22_34_real,
  output     [15:0]   io_coef_out_payload_0_22_34_imag,
  output     [15:0]   io_coef_out_payload_0_22_35_real,
  output     [15:0]   io_coef_out_payload_0_22_35_imag,
  output     [15:0]   io_coef_out_payload_0_22_36_real,
  output     [15:0]   io_coef_out_payload_0_22_36_imag,
  output     [15:0]   io_coef_out_payload_0_22_37_real,
  output     [15:0]   io_coef_out_payload_0_22_37_imag,
  output     [15:0]   io_coef_out_payload_0_22_38_real,
  output     [15:0]   io_coef_out_payload_0_22_38_imag,
  output     [15:0]   io_coef_out_payload_0_22_39_real,
  output     [15:0]   io_coef_out_payload_0_22_39_imag,
  output     [15:0]   io_coef_out_payload_0_22_40_real,
  output     [15:0]   io_coef_out_payload_0_22_40_imag,
  output     [15:0]   io_coef_out_payload_0_22_41_real,
  output     [15:0]   io_coef_out_payload_0_22_41_imag,
  output     [15:0]   io_coef_out_payload_0_22_42_real,
  output     [15:0]   io_coef_out_payload_0_22_42_imag,
  output     [15:0]   io_coef_out_payload_0_22_43_real,
  output     [15:0]   io_coef_out_payload_0_22_43_imag,
  output     [15:0]   io_coef_out_payload_0_22_44_real,
  output     [15:0]   io_coef_out_payload_0_22_44_imag,
  output     [15:0]   io_coef_out_payload_0_22_45_real,
  output     [15:0]   io_coef_out_payload_0_22_45_imag,
  output     [15:0]   io_coef_out_payload_0_22_46_real,
  output     [15:0]   io_coef_out_payload_0_22_46_imag,
  output     [15:0]   io_coef_out_payload_0_22_47_real,
  output     [15:0]   io_coef_out_payload_0_22_47_imag,
  output     [15:0]   io_coef_out_payload_0_22_48_real,
  output     [15:0]   io_coef_out_payload_0_22_48_imag,
  output     [15:0]   io_coef_out_payload_0_22_49_real,
  output     [15:0]   io_coef_out_payload_0_22_49_imag,
  output     [15:0]   io_coef_out_payload_0_23_0_real,
  output     [15:0]   io_coef_out_payload_0_23_0_imag,
  output     [15:0]   io_coef_out_payload_0_23_1_real,
  output     [15:0]   io_coef_out_payload_0_23_1_imag,
  output     [15:0]   io_coef_out_payload_0_23_2_real,
  output     [15:0]   io_coef_out_payload_0_23_2_imag,
  output     [15:0]   io_coef_out_payload_0_23_3_real,
  output     [15:0]   io_coef_out_payload_0_23_3_imag,
  output     [15:0]   io_coef_out_payload_0_23_4_real,
  output     [15:0]   io_coef_out_payload_0_23_4_imag,
  output     [15:0]   io_coef_out_payload_0_23_5_real,
  output     [15:0]   io_coef_out_payload_0_23_5_imag,
  output     [15:0]   io_coef_out_payload_0_23_6_real,
  output     [15:0]   io_coef_out_payload_0_23_6_imag,
  output     [15:0]   io_coef_out_payload_0_23_7_real,
  output     [15:0]   io_coef_out_payload_0_23_7_imag,
  output     [15:0]   io_coef_out_payload_0_23_8_real,
  output     [15:0]   io_coef_out_payload_0_23_8_imag,
  output     [15:0]   io_coef_out_payload_0_23_9_real,
  output     [15:0]   io_coef_out_payload_0_23_9_imag,
  output     [15:0]   io_coef_out_payload_0_23_10_real,
  output     [15:0]   io_coef_out_payload_0_23_10_imag,
  output     [15:0]   io_coef_out_payload_0_23_11_real,
  output     [15:0]   io_coef_out_payload_0_23_11_imag,
  output     [15:0]   io_coef_out_payload_0_23_12_real,
  output     [15:0]   io_coef_out_payload_0_23_12_imag,
  output     [15:0]   io_coef_out_payload_0_23_13_real,
  output     [15:0]   io_coef_out_payload_0_23_13_imag,
  output     [15:0]   io_coef_out_payload_0_23_14_real,
  output     [15:0]   io_coef_out_payload_0_23_14_imag,
  output     [15:0]   io_coef_out_payload_0_23_15_real,
  output     [15:0]   io_coef_out_payload_0_23_15_imag,
  output     [15:0]   io_coef_out_payload_0_23_16_real,
  output     [15:0]   io_coef_out_payload_0_23_16_imag,
  output     [15:0]   io_coef_out_payload_0_23_17_real,
  output     [15:0]   io_coef_out_payload_0_23_17_imag,
  output     [15:0]   io_coef_out_payload_0_23_18_real,
  output     [15:0]   io_coef_out_payload_0_23_18_imag,
  output     [15:0]   io_coef_out_payload_0_23_19_real,
  output     [15:0]   io_coef_out_payload_0_23_19_imag,
  output     [15:0]   io_coef_out_payload_0_23_20_real,
  output     [15:0]   io_coef_out_payload_0_23_20_imag,
  output     [15:0]   io_coef_out_payload_0_23_21_real,
  output     [15:0]   io_coef_out_payload_0_23_21_imag,
  output     [15:0]   io_coef_out_payload_0_23_22_real,
  output     [15:0]   io_coef_out_payload_0_23_22_imag,
  output     [15:0]   io_coef_out_payload_0_23_23_real,
  output     [15:0]   io_coef_out_payload_0_23_23_imag,
  output     [15:0]   io_coef_out_payload_0_23_24_real,
  output     [15:0]   io_coef_out_payload_0_23_24_imag,
  output     [15:0]   io_coef_out_payload_0_23_25_real,
  output     [15:0]   io_coef_out_payload_0_23_25_imag,
  output     [15:0]   io_coef_out_payload_0_23_26_real,
  output     [15:0]   io_coef_out_payload_0_23_26_imag,
  output     [15:0]   io_coef_out_payload_0_23_27_real,
  output     [15:0]   io_coef_out_payload_0_23_27_imag,
  output     [15:0]   io_coef_out_payload_0_23_28_real,
  output     [15:0]   io_coef_out_payload_0_23_28_imag,
  output     [15:0]   io_coef_out_payload_0_23_29_real,
  output     [15:0]   io_coef_out_payload_0_23_29_imag,
  output     [15:0]   io_coef_out_payload_0_23_30_real,
  output     [15:0]   io_coef_out_payload_0_23_30_imag,
  output     [15:0]   io_coef_out_payload_0_23_31_real,
  output     [15:0]   io_coef_out_payload_0_23_31_imag,
  output     [15:0]   io_coef_out_payload_0_23_32_real,
  output     [15:0]   io_coef_out_payload_0_23_32_imag,
  output     [15:0]   io_coef_out_payload_0_23_33_real,
  output     [15:0]   io_coef_out_payload_0_23_33_imag,
  output     [15:0]   io_coef_out_payload_0_23_34_real,
  output     [15:0]   io_coef_out_payload_0_23_34_imag,
  output     [15:0]   io_coef_out_payload_0_23_35_real,
  output     [15:0]   io_coef_out_payload_0_23_35_imag,
  output     [15:0]   io_coef_out_payload_0_23_36_real,
  output     [15:0]   io_coef_out_payload_0_23_36_imag,
  output     [15:0]   io_coef_out_payload_0_23_37_real,
  output     [15:0]   io_coef_out_payload_0_23_37_imag,
  output     [15:0]   io_coef_out_payload_0_23_38_real,
  output     [15:0]   io_coef_out_payload_0_23_38_imag,
  output     [15:0]   io_coef_out_payload_0_23_39_real,
  output     [15:0]   io_coef_out_payload_0_23_39_imag,
  output     [15:0]   io_coef_out_payload_0_23_40_real,
  output     [15:0]   io_coef_out_payload_0_23_40_imag,
  output     [15:0]   io_coef_out_payload_0_23_41_real,
  output     [15:0]   io_coef_out_payload_0_23_41_imag,
  output     [15:0]   io_coef_out_payload_0_23_42_real,
  output     [15:0]   io_coef_out_payload_0_23_42_imag,
  output     [15:0]   io_coef_out_payload_0_23_43_real,
  output     [15:0]   io_coef_out_payload_0_23_43_imag,
  output     [15:0]   io_coef_out_payload_0_23_44_real,
  output     [15:0]   io_coef_out_payload_0_23_44_imag,
  output     [15:0]   io_coef_out_payload_0_23_45_real,
  output     [15:0]   io_coef_out_payload_0_23_45_imag,
  output     [15:0]   io_coef_out_payload_0_23_46_real,
  output     [15:0]   io_coef_out_payload_0_23_46_imag,
  output     [15:0]   io_coef_out_payload_0_23_47_real,
  output     [15:0]   io_coef_out_payload_0_23_47_imag,
  output     [15:0]   io_coef_out_payload_0_23_48_real,
  output     [15:0]   io_coef_out_payload_0_23_48_imag,
  output     [15:0]   io_coef_out_payload_0_23_49_real,
  output     [15:0]   io_coef_out_payload_0_23_49_imag,
  output     [15:0]   io_coef_out_payload_0_24_0_real,
  output     [15:0]   io_coef_out_payload_0_24_0_imag,
  output     [15:0]   io_coef_out_payload_0_24_1_real,
  output     [15:0]   io_coef_out_payload_0_24_1_imag,
  output     [15:0]   io_coef_out_payload_0_24_2_real,
  output     [15:0]   io_coef_out_payload_0_24_2_imag,
  output     [15:0]   io_coef_out_payload_0_24_3_real,
  output     [15:0]   io_coef_out_payload_0_24_3_imag,
  output     [15:0]   io_coef_out_payload_0_24_4_real,
  output     [15:0]   io_coef_out_payload_0_24_4_imag,
  output     [15:0]   io_coef_out_payload_0_24_5_real,
  output     [15:0]   io_coef_out_payload_0_24_5_imag,
  output     [15:0]   io_coef_out_payload_0_24_6_real,
  output     [15:0]   io_coef_out_payload_0_24_6_imag,
  output     [15:0]   io_coef_out_payload_0_24_7_real,
  output     [15:0]   io_coef_out_payload_0_24_7_imag,
  output     [15:0]   io_coef_out_payload_0_24_8_real,
  output     [15:0]   io_coef_out_payload_0_24_8_imag,
  output     [15:0]   io_coef_out_payload_0_24_9_real,
  output     [15:0]   io_coef_out_payload_0_24_9_imag,
  output     [15:0]   io_coef_out_payload_0_24_10_real,
  output     [15:0]   io_coef_out_payload_0_24_10_imag,
  output     [15:0]   io_coef_out_payload_0_24_11_real,
  output     [15:0]   io_coef_out_payload_0_24_11_imag,
  output     [15:0]   io_coef_out_payload_0_24_12_real,
  output     [15:0]   io_coef_out_payload_0_24_12_imag,
  output     [15:0]   io_coef_out_payload_0_24_13_real,
  output     [15:0]   io_coef_out_payload_0_24_13_imag,
  output     [15:0]   io_coef_out_payload_0_24_14_real,
  output     [15:0]   io_coef_out_payload_0_24_14_imag,
  output     [15:0]   io_coef_out_payload_0_24_15_real,
  output     [15:0]   io_coef_out_payload_0_24_15_imag,
  output     [15:0]   io_coef_out_payload_0_24_16_real,
  output     [15:0]   io_coef_out_payload_0_24_16_imag,
  output     [15:0]   io_coef_out_payload_0_24_17_real,
  output     [15:0]   io_coef_out_payload_0_24_17_imag,
  output     [15:0]   io_coef_out_payload_0_24_18_real,
  output     [15:0]   io_coef_out_payload_0_24_18_imag,
  output     [15:0]   io_coef_out_payload_0_24_19_real,
  output     [15:0]   io_coef_out_payload_0_24_19_imag,
  output     [15:0]   io_coef_out_payload_0_24_20_real,
  output     [15:0]   io_coef_out_payload_0_24_20_imag,
  output     [15:0]   io_coef_out_payload_0_24_21_real,
  output     [15:0]   io_coef_out_payload_0_24_21_imag,
  output     [15:0]   io_coef_out_payload_0_24_22_real,
  output     [15:0]   io_coef_out_payload_0_24_22_imag,
  output     [15:0]   io_coef_out_payload_0_24_23_real,
  output     [15:0]   io_coef_out_payload_0_24_23_imag,
  output     [15:0]   io_coef_out_payload_0_24_24_real,
  output     [15:0]   io_coef_out_payload_0_24_24_imag,
  output     [15:0]   io_coef_out_payload_0_24_25_real,
  output     [15:0]   io_coef_out_payload_0_24_25_imag,
  output     [15:0]   io_coef_out_payload_0_24_26_real,
  output     [15:0]   io_coef_out_payload_0_24_26_imag,
  output     [15:0]   io_coef_out_payload_0_24_27_real,
  output     [15:0]   io_coef_out_payload_0_24_27_imag,
  output     [15:0]   io_coef_out_payload_0_24_28_real,
  output     [15:0]   io_coef_out_payload_0_24_28_imag,
  output     [15:0]   io_coef_out_payload_0_24_29_real,
  output     [15:0]   io_coef_out_payload_0_24_29_imag,
  output     [15:0]   io_coef_out_payload_0_24_30_real,
  output     [15:0]   io_coef_out_payload_0_24_30_imag,
  output     [15:0]   io_coef_out_payload_0_24_31_real,
  output     [15:0]   io_coef_out_payload_0_24_31_imag,
  output     [15:0]   io_coef_out_payload_0_24_32_real,
  output     [15:0]   io_coef_out_payload_0_24_32_imag,
  output     [15:0]   io_coef_out_payload_0_24_33_real,
  output     [15:0]   io_coef_out_payload_0_24_33_imag,
  output     [15:0]   io_coef_out_payload_0_24_34_real,
  output     [15:0]   io_coef_out_payload_0_24_34_imag,
  output     [15:0]   io_coef_out_payload_0_24_35_real,
  output     [15:0]   io_coef_out_payload_0_24_35_imag,
  output     [15:0]   io_coef_out_payload_0_24_36_real,
  output     [15:0]   io_coef_out_payload_0_24_36_imag,
  output     [15:0]   io_coef_out_payload_0_24_37_real,
  output     [15:0]   io_coef_out_payload_0_24_37_imag,
  output     [15:0]   io_coef_out_payload_0_24_38_real,
  output     [15:0]   io_coef_out_payload_0_24_38_imag,
  output     [15:0]   io_coef_out_payload_0_24_39_real,
  output     [15:0]   io_coef_out_payload_0_24_39_imag,
  output     [15:0]   io_coef_out_payload_0_24_40_real,
  output     [15:0]   io_coef_out_payload_0_24_40_imag,
  output     [15:0]   io_coef_out_payload_0_24_41_real,
  output     [15:0]   io_coef_out_payload_0_24_41_imag,
  output     [15:0]   io_coef_out_payload_0_24_42_real,
  output     [15:0]   io_coef_out_payload_0_24_42_imag,
  output     [15:0]   io_coef_out_payload_0_24_43_real,
  output     [15:0]   io_coef_out_payload_0_24_43_imag,
  output     [15:0]   io_coef_out_payload_0_24_44_real,
  output     [15:0]   io_coef_out_payload_0_24_44_imag,
  output     [15:0]   io_coef_out_payload_0_24_45_real,
  output     [15:0]   io_coef_out_payload_0_24_45_imag,
  output     [15:0]   io_coef_out_payload_0_24_46_real,
  output     [15:0]   io_coef_out_payload_0_24_46_imag,
  output     [15:0]   io_coef_out_payload_0_24_47_real,
  output     [15:0]   io_coef_out_payload_0_24_47_imag,
  output     [15:0]   io_coef_out_payload_0_24_48_real,
  output     [15:0]   io_coef_out_payload_0_24_48_imag,
  output     [15:0]   io_coef_out_payload_0_24_49_real,
  output     [15:0]   io_coef_out_payload_0_24_49_imag,
  output     [15:0]   io_coef_out_payload_0_25_0_real,
  output     [15:0]   io_coef_out_payload_0_25_0_imag,
  output     [15:0]   io_coef_out_payload_0_25_1_real,
  output     [15:0]   io_coef_out_payload_0_25_1_imag,
  output     [15:0]   io_coef_out_payload_0_25_2_real,
  output     [15:0]   io_coef_out_payload_0_25_2_imag,
  output     [15:0]   io_coef_out_payload_0_25_3_real,
  output     [15:0]   io_coef_out_payload_0_25_3_imag,
  output     [15:0]   io_coef_out_payload_0_25_4_real,
  output     [15:0]   io_coef_out_payload_0_25_4_imag,
  output     [15:0]   io_coef_out_payload_0_25_5_real,
  output     [15:0]   io_coef_out_payload_0_25_5_imag,
  output     [15:0]   io_coef_out_payload_0_25_6_real,
  output     [15:0]   io_coef_out_payload_0_25_6_imag,
  output     [15:0]   io_coef_out_payload_0_25_7_real,
  output     [15:0]   io_coef_out_payload_0_25_7_imag,
  output     [15:0]   io_coef_out_payload_0_25_8_real,
  output     [15:0]   io_coef_out_payload_0_25_8_imag,
  output     [15:0]   io_coef_out_payload_0_25_9_real,
  output     [15:0]   io_coef_out_payload_0_25_9_imag,
  output     [15:0]   io_coef_out_payload_0_25_10_real,
  output     [15:0]   io_coef_out_payload_0_25_10_imag,
  output     [15:0]   io_coef_out_payload_0_25_11_real,
  output     [15:0]   io_coef_out_payload_0_25_11_imag,
  output     [15:0]   io_coef_out_payload_0_25_12_real,
  output     [15:0]   io_coef_out_payload_0_25_12_imag,
  output     [15:0]   io_coef_out_payload_0_25_13_real,
  output     [15:0]   io_coef_out_payload_0_25_13_imag,
  output     [15:0]   io_coef_out_payload_0_25_14_real,
  output     [15:0]   io_coef_out_payload_0_25_14_imag,
  output     [15:0]   io_coef_out_payload_0_25_15_real,
  output     [15:0]   io_coef_out_payload_0_25_15_imag,
  output     [15:0]   io_coef_out_payload_0_25_16_real,
  output     [15:0]   io_coef_out_payload_0_25_16_imag,
  output     [15:0]   io_coef_out_payload_0_25_17_real,
  output     [15:0]   io_coef_out_payload_0_25_17_imag,
  output     [15:0]   io_coef_out_payload_0_25_18_real,
  output     [15:0]   io_coef_out_payload_0_25_18_imag,
  output     [15:0]   io_coef_out_payload_0_25_19_real,
  output     [15:0]   io_coef_out_payload_0_25_19_imag,
  output     [15:0]   io_coef_out_payload_0_25_20_real,
  output     [15:0]   io_coef_out_payload_0_25_20_imag,
  output     [15:0]   io_coef_out_payload_0_25_21_real,
  output     [15:0]   io_coef_out_payload_0_25_21_imag,
  output     [15:0]   io_coef_out_payload_0_25_22_real,
  output     [15:0]   io_coef_out_payload_0_25_22_imag,
  output     [15:0]   io_coef_out_payload_0_25_23_real,
  output     [15:0]   io_coef_out_payload_0_25_23_imag,
  output     [15:0]   io_coef_out_payload_0_25_24_real,
  output     [15:0]   io_coef_out_payload_0_25_24_imag,
  output     [15:0]   io_coef_out_payload_0_25_25_real,
  output     [15:0]   io_coef_out_payload_0_25_25_imag,
  output     [15:0]   io_coef_out_payload_0_25_26_real,
  output     [15:0]   io_coef_out_payload_0_25_26_imag,
  output     [15:0]   io_coef_out_payload_0_25_27_real,
  output     [15:0]   io_coef_out_payload_0_25_27_imag,
  output     [15:0]   io_coef_out_payload_0_25_28_real,
  output     [15:0]   io_coef_out_payload_0_25_28_imag,
  output     [15:0]   io_coef_out_payload_0_25_29_real,
  output     [15:0]   io_coef_out_payload_0_25_29_imag,
  output     [15:0]   io_coef_out_payload_0_25_30_real,
  output     [15:0]   io_coef_out_payload_0_25_30_imag,
  output     [15:0]   io_coef_out_payload_0_25_31_real,
  output     [15:0]   io_coef_out_payload_0_25_31_imag,
  output     [15:0]   io_coef_out_payload_0_25_32_real,
  output     [15:0]   io_coef_out_payload_0_25_32_imag,
  output     [15:0]   io_coef_out_payload_0_25_33_real,
  output     [15:0]   io_coef_out_payload_0_25_33_imag,
  output     [15:0]   io_coef_out_payload_0_25_34_real,
  output     [15:0]   io_coef_out_payload_0_25_34_imag,
  output     [15:0]   io_coef_out_payload_0_25_35_real,
  output     [15:0]   io_coef_out_payload_0_25_35_imag,
  output     [15:0]   io_coef_out_payload_0_25_36_real,
  output     [15:0]   io_coef_out_payload_0_25_36_imag,
  output     [15:0]   io_coef_out_payload_0_25_37_real,
  output     [15:0]   io_coef_out_payload_0_25_37_imag,
  output     [15:0]   io_coef_out_payload_0_25_38_real,
  output     [15:0]   io_coef_out_payload_0_25_38_imag,
  output     [15:0]   io_coef_out_payload_0_25_39_real,
  output     [15:0]   io_coef_out_payload_0_25_39_imag,
  output     [15:0]   io_coef_out_payload_0_25_40_real,
  output     [15:0]   io_coef_out_payload_0_25_40_imag,
  output     [15:0]   io_coef_out_payload_0_25_41_real,
  output     [15:0]   io_coef_out_payload_0_25_41_imag,
  output     [15:0]   io_coef_out_payload_0_25_42_real,
  output     [15:0]   io_coef_out_payload_0_25_42_imag,
  output     [15:0]   io_coef_out_payload_0_25_43_real,
  output     [15:0]   io_coef_out_payload_0_25_43_imag,
  output     [15:0]   io_coef_out_payload_0_25_44_real,
  output     [15:0]   io_coef_out_payload_0_25_44_imag,
  output     [15:0]   io_coef_out_payload_0_25_45_real,
  output     [15:0]   io_coef_out_payload_0_25_45_imag,
  output     [15:0]   io_coef_out_payload_0_25_46_real,
  output     [15:0]   io_coef_out_payload_0_25_46_imag,
  output     [15:0]   io_coef_out_payload_0_25_47_real,
  output     [15:0]   io_coef_out_payload_0_25_47_imag,
  output     [15:0]   io_coef_out_payload_0_25_48_real,
  output     [15:0]   io_coef_out_payload_0_25_48_imag,
  output     [15:0]   io_coef_out_payload_0_25_49_real,
  output     [15:0]   io_coef_out_payload_0_25_49_imag,
  output     [15:0]   io_coef_out_payload_0_26_0_real,
  output     [15:0]   io_coef_out_payload_0_26_0_imag,
  output     [15:0]   io_coef_out_payload_0_26_1_real,
  output     [15:0]   io_coef_out_payload_0_26_1_imag,
  output     [15:0]   io_coef_out_payload_0_26_2_real,
  output     [15:0]   io_coef_out_payload_0_26_2_imag,
  output     [15:0]   io_coef_out_payload_0_26_3_real,
  output     [15:0]   io_coef_out_payload_0_26_3_imag,
  output     [15:0]   io_coef_out_payload_0_26_4_real,
  output     [15:0]   io_coef_out_payload_0_26_4_imag,
  output     [15:0]   io_coef_out_payload_0_26_5_real,
  output     [15:0]   io_coef_out_payload_0_26_5_imag,
  output     [15:0]   io_coef_out_payload_0_26_6_real,
  output     [15:0]   io_coef_out_payload_0_26_6_imag,
  output     [15:0]   io_coef_out_payload_0_26_7_real,
  output     [15:0]   io_coef_out_payload_0_26_7_imag,
  output     [15:0]   io_coef_out_payload_0_26_8_real,
  output     [15:0]   io_coef_out_payload_0_26_8_imag,
  output     [15:0]   io_coef_out_payload_0_26_9_real,
  output     [15:0]   io_coef_out_payload_0_26_9_imag,
  output     [15:0]   io_coef_out_payload_0_26_10_real,
  output     [15:0]   io_coef_out_payload_0_26_10_imag,
  output     [15:0]   io_coef_out_payload_0_26_11_real,
  output     [15:0]   io_coef_out_payload_0_26_11_imag,
  output     [15:0]   io_coef_out_payload_0_26_12_real,
  output     [15:0]   io_coef_out_payload_0_26_12_imag,
  output     [15:0]   io_coef_out_payload_0_26_13_real,
  output     [15:0]   io_coef_out_payload_0_26_13_imag,
  output     [15:0]   io_coef_out_payload_0_26_14_real,
  output     [15:0]   io_coef_out_payload_0_26_14_imag,
  output     [15:0]   io_coef_out_payload_0_26_15_real,
  output     [15:0]   io_coef_out_payload_0_26_15_imag,
  output     [15:0]   io_coef_out_payload_0_26_16_real,
  output     [15:0]   io_coef_out_payload_0_26_16_imag,
  output     [15:0]   io_coef_out_payload_0_26_17_real,
  output     [15:0]   io_coef_out_payload_0_26_17_imag,
  output     [15:0]   io_coef_out_payload_0_26_18_real,
  output     [15:0]   io_coef_out_payload_0_26_18_imag,
  output     [15:0]   io_coef_out_payload_0_26_19_real,
  output     [15:0]   io_coef_out_payload_0_26_19_imag,
  output     [15:0]   io_coef_out_payload_0_26_20_real,
  output     [15:0]   io_coef_out_payload_0_26_20_imag,
  output     [15:0]   io_coef_out_payload_0_26_21_real,
  output     [15:0]   io_coef_out_payload_0_26_21_imag,
  output     [15:0]   io_coef_out_payload_0_26_22_real,
  output     [15:0]   io_coef_out_payload_0_26_22_imag,
  output     [15:0]   io_coef_out_payload_0_26_23_real,
  output     [15:0]   io_coef_out_payload_0_26_23_imag,
  output     [15:0]   io_coef_out_payload_0_26_24_real,
  output     [15:0]   io_coef_out_payload_0_26_24_imag,
  output     [15:0]   io_coef_out_payload_0_26_25_real,
  output     [15:0]   io_coef_out_payload_0_26_25_imag,
  output     [15:0]   io_coef_out_payload_0_26_26_real,
  output     [15:0]   io_coef_out_payload_0_26_26_imag,
  output     [15:0]   io_coef_out_payload_0_26_27_real,
  output     [15:0]   io_coef_out_payload_0_26_27_imag,
  output     [15:0]   io_coef_out_payload_0_26_28_real,
  output     [15:0]   io_coef_out_payload_0_26_28_imag,
  output     [15:0]   io_coef_out_payload_0_26_29_real,
  output     [15:0]   io_coef_out_payload_0_26_29_imag,
  output     [15:0]   io_coef_out_payload_0_26_30_real,
  output     [15:0]   io_coef_out_payload_0_26_30_imag,
  output     [15:0]   io_coef_out_payload_0_26_31_real,
  output     [15:0]   io_coef_out_payload_0_26_31_imag,
  output     [15:0]   io_coef_out_payload_0_26_32_real,
  output     [15:0]   io_coef_out_payload_0_26_32_imag,
  output     [15:0]   io_coef_out_payload_0_26_33_real,
  output     [15:0]   io_coef_out_payload_0_26_33_imag,
  output     [15:0]   io_coef_out_payload_0_26_34_real,
  output     [15:0]   io_coef_out_payload_0_26_34_imag,
  output     [15:0]   io_coef_out_payload_0_26_35_real,
  output     [15:0]   io_coef_out_payload_0_26_35_imag,
  output     [15:0]   io_coef_out_payload_0_26_36_real,
  output     [15:0]   io_coef_out_payload_0_26_36_imag,
  output     [15:0]   io_coef_out_payload_0_26_37_real,
  output     [15:0]   io_coef_out_payload_0_26_37_imag,
  output     [15:0]   io_coef_out_payload_0_26_38_real,
  output     [15:0]   io_coef_out_payload_0_26_38_imag,
  output     [15:0]   io_coef_out_payload_0_26_39_real,
  output     [15:0]   io_coef_out_payload_0_26_39_imag,
  output     [15:0]   io_coef_out_payload_0_26_40_real,
  output     [15:0]   io_coef_out_payload_0_26_40_imag,
  output     [15:0]   io_coef_out_payload_0_26_41_real,
  output     [15:0]   io_coef_out_payload_0_26_41_imag,
  output     [15:0]   io_coef_out_payload_0_26_42_real,
  output     [15:0]   io_coef_out_payload_0_26_42_imag,
  output     [15:0]   io_coef_out_payload_0_26_43_real,
  output     [15:0]   io_coef_out_payload_0_26_43_imag,
  output     [15:0]   io_coef_out_payload_0_26_44_real,
  output     [15:0]   io_coef_out_payload_0_26_44_imag,
  output     [15:0]   io_coef_out_payload_0_26_45_real,
  output     [15:0]   io_coef_out_payload_0_26_45_imag,
  output     [15:0]   io_coef_out_payload_0_26_46_real,
  output     [15:0]   io_coef_out_payload_0_26_46_imag,
  output     [15:0]   io_coef_out_payload_0_26_47_real,
  output     [15:0]   io_coef_out_payload_0_26_47_imag,
  output     [15:0]   io_coef_out_payload_0_26_48_real,
  output     [15:0]   io_coef_out_payload_0_26_48_imag,
  output     [15:0]   io_coef_out_payload_0_26_49_real,
  output     [15:0]   io_coef_out_payload_0_26_49_imag,
  output     [15:0]   io_coef_out_payload_0_27_0_real,
  output     [15:0]   io_coef_out_payload_0_27_0_imag,
  output     [15:0]   io_coef_out_payload_0_27_1_real,
  output     [15:0]   io_coef_out_payload_0_27_1_imag,
  output     [15:0]   io_coef_out_payload_0_27_2_real,
  output     [15:0]   io_coef_out_payload_0_27_2_imag,
  output     [15:0]   io_coef_out_payload_0_27_3_real,
  output     [15:0]   io_coef_out_payload_0_27_3_imag,
  output     [15:0]   io_coef_out_payload_0_27_4_real,
  output     [15:0]   io_coef_out_payload_0_27_4_imag,
  output     [15:0]   io_coef_out_payload_0_27_5_real,
  output     [15:0]   io_coef_out_payload_0_27_5_imag,
  output     [15:0]   io_coef_out_payload_0_27_6_real,
  output     [15:0]   io_coef_out_payload_0_27_6_imag,
  output     [15:0]   io_coef_out_payload_0_27_7_real,
  output     [15:0]   io_coef_out_payload_0_27_7_imag,
  output     [15:0]   io_coef_out_payload_0_27_8_real,
  output     [15:0]   io_coef_out_payload_0_27_8_imag,
  output     [15:0]   io_coef_out_payload_0_27_9_real,
  output     [15:0]   io_coef_out_payload_0_27_9_imag,
  output     [15:0]   io_coef_out_payload_0_27_10_real,
  output     [15:0]   io_coef_out_payload_0_27_10_imag,
  output     [15:0]   io_coef_out_payload_0_27_11_real,
  output     [15:0]   io_coef_out_payload_0_27_11_imag,
  output     [15:0]   io_coef_out_payload_0_27_12_real,
  output     [15:0]   io_coef_out_payload_0_27_12_imag,
  output     [15:0]   io_coef_out_payload_0_27_13_real,
  output     [15:0]   io_coef_out_payload_0_27_13_imag,
  output     [15:0]   io_coef_out_payload_0_27_14_real,
  output     [15:0]   io_coef_out_payload_0_27_14_imag,
  output     [15:0]   io_coef_out_payload_0_27_15_real,
  output     [15:0]   io_coef_out_payload_0_27_15_imag,
  output     [15:0]   io_coef_out_payload_0_27_16_real,
  output     [15:0]   io_coef_out_payload_0_27_16_imag,
  output     [15:0]   io_coef_out_payload_0_27_17_real,
  output     [15:0]   io_coef_out_payload_0_27_17_imag,
  output     [15:0]   io_coef_out_payload_0_27_18_real,
  output     [15:0]   io_coef_out_payload_0_27_18_imag,
  output     [15:0]   io_coef_out_payload_0_27_19_real,
  output     [15:0]   io_coef_out_payload_0_27_19_imag,
  output     [15:0]   io_coef_out_payload_0_27_20_real,
  output     [15:0]   io_coef_out_payload_0_27_20_imag,
  output     [15:0]   io_coef_out_payload_0_27_21_real,
  output     [15:0]   io_coef_out_payload_0_27_21_imag,
  output     [15:0]   io_coef_out_payload_0_27_22_real,
  output     [15:0]   io_coef_out_payload_0_27_22_imag,
  output     [15:0]   io_coef_out_payload_0_27_23_real,
  output     [15:0]   io_coef_out_payload_0_27_23_imag,
  output     [15:0]   io_coef_out_payload_0_27_24_real,
  output     [15:0]   io_coef_out_payload_0_27_24_imag,
  output     [15:0]   io_coef_out_payload_0_27_25_real,
  output     [15:0]   io_coef_out_payload_0_27_25_imag,
  output     [15:0]   io_coef_out_payload_0_27_26_real,
  output     [15:0]   io_coef_out_payload_0_27_26_imag,
  output     [15:0]   io_coef_out_payload_0_27_27_real,
  output     [15:0]   io_coef_out_payload_0_27_27_imag,
  output     [15:0]   io_coef_out_payload_0_27_28_real,
  output     [15:0]   io_coef_out_payload_0_27_28_imag,
  output     [15:0]   io_coef_out_payload_0_27_29_real,
  output     [15:0]   io_coef_out_payload_0_27_29_imag,
  output     [15:0]   io_coef_out_payload_0_27_30_real,
  output     [15:0]   io_coef_out_payload_0_27_30_imag,
  output     [15:0]   io_coef_out_payload_0_27_31_real,
  output     [15:0]   io_coef_out_payload_0_27_31_imag,
  output     [15:0]   io_coef_out_payload_0_27_32_real,
  output     [15:0]   io_coef_out_payload_0_27_32_imag,
  output     [15:0]   io_coef_out_payload_0_27_33_real,
  output     [15:0]   io_coef_out_payload_0_27_33_imag,
  output     [15:0]   io_coef_out_payload_0_27_34_real,
  output     [15:0]   io_coef_out_payload_0_27_34_imag,
  output     [15:0]   io_coef_out_payload_0_27_35_real,
  output     [15:0]   io_coef_out_payload_0_27_35_imag,
  output     [15:0]   io_coef_out_payload_0_27_36_real,
  output     [15:0]   io_coef_out_payload_0_27_36_imag,
  output     [15:0]   io_coef_out_payload_0_27_37_real,
  output     [15:0]   io_coef_out_payload_0_27_37_imag,
  output     [15:0]   io_coef_out_payload_0_27_38_real,
  output     [15:0]   io_coef_out_payload_0_27_38_imag,
  output     [15:0]   io_coef_out_payload_0_27_39_real,
  output     [15:0]   io_coef_out_payload_0_27_39_imag,
  output     [15:0]   io_coef_out_payload_0_27_40_real,
  output     [15:0]   io_coef_out_payload_0_27_40_imag,
  output     [15:0]   io_coef_out_payload_0_27_41_real,
  output     [15:0]   io_coef_out_payload_0_27_41_imag,
  output     [15:0]   io_coef_out_payload_0_27_42_real,
  output     [15:0]   io_coef_out_payload_0_27_42_imag,
  output     [15:0]   io_coef_out_payload_0_27_43_real,
  output     [15:0]   io_coef_out_payload_0_27_43_imag,
  output     [15:0]   io_coef_out_payload_0_27_44_real,
  output     [15:0]   io_coef_out_payload_0_27_44_imag,
  output     [15:0]   io_coef_out_payload_0_27_45_real,
  output     [15:0]   io_coef_out_payload_0_27_45_imag,
  output     [15:0]   io_coef_out_payload_0_27_46_real,
  output     [15:0]   io_coef_out_payload_0_27_46_imag,
  output     [15:0]   io_coef_out_payload_0_27_47_real,
  output     [15:0]   io_coef_out_payload_0_27_47_imag,
  output     [15:0]   io_coef_out_payload_0_27_48_real,
  output     [15:0]   io_coef_out_payload_0_27_48_imag,
  output     [15:0]   io_coef_out_payload_0_27_49_real,
  output     [15:0]   io_coef_out_payload_0_27_49_imag,
  output     [15:0]   io_coef_out_payload_0_28_0_real,
  output     [15:0]   io_coef_out_payload_0_28_0_imag,
  output     [15:0]   io_coef_out_payload_0_28_1_real,
  output     [15:0]   io_coef_out_payload_0_28_1_imag,
  output     [15:0]   io_coef_out_payload_0_28_2_real,
  output     [15:0]   io_coef_out_payload_0_28_2_imag,
  output     [15:0]   io_coef_out_payload_0_28_3_real,
  output     [15:0]   io_coef_out_payload_0_28_3_imag,
  output     [15:0]   io_coef_out_payload_0_28_4_real,
  output     [15:0]   io_coef_out_payload_0_28_4_imag,
  output     [15:0]   io_coef_out_payload_0_28_5_real,
  output     [15:0]   io_coef_out_payload_0_28_5_imag,
  output     [15:0]   io_coef_out_payload_0_28_6_real,
  output     [15:0]   io_coef_out_payload_0_28_6_imag,
  output     [15:0]   io_coef_out_payload_0_28_7_real,
  output     [15:0]   io_coef_out_payload_0_28_7_imag,
  output     [15:0]   io_coef_out_payload_0_28_8_real,
  output     [15:0]   io_coef_out_payload_0_28_8_imag,
  output     [15:0]   io_coef_out_payload_0_28_9_real,
  output     [15:0]   io_coef_out_payload_0_28_9_imag,
  output     [15:0]   io_coef_out_payload_0_28_10_real,
  output     [15:0]   io_coef_out_payload_0_28_10_imag,
  output     [15:0]   io_coef_out_payload_0_28_11_real,
  output     [15:0]   io_coef_out_payload_0_28_11_imag,
  output     [15:0]   io_coef_out_payload_0_28_12_real,
  output     [15:0]   io_coef_out_payload_0_28_12_imag,
  output     [15:0]   io_coef_out_payload_0_28_13_real,
  output     [15:0]   io_coef_out_payload_0_28_13_imag,
  output     [15:0]   io_coef_out_payload_0_28_14_real,
  output     [15:0]   io_coef_out_payload_0_28_14_imag,
  output     [15:0]   io_coef_out_payload_0_28_15_real,
  output     [15:0]   io_coef_out_payload_0_28_15_imag,
  output     [15:0]   io_coef_out_payload_0_28_16_real,
  output     [15:0]   io_coef_out_payload_0_28_16_imag,
  output     [15:0]   io_coef_out_payload_0_28_17_real,
  output     [15:0]   io_coef_out_payload_0_28_17_imag,
  output     [15:0]   io_coef_out_payload_0_28_18_real,
  output     [15:0]   io_coef_out_payload_0_28_18_imag,
  output     [15:0]   io_coef_out_payload_0_28_19_real,
  output     [15:0]   io_coef_out_payload_0_28_19_imag,
  output     [15:0]   io_coef_out_payload_0_28_20_real,
  output     [15:0]   io_coef_out_payload_0_28_20_imag,
  output     [15:0]   io_coef_out_payload_0_28_21_real,
  output     [15:0]   io_coef_out_payload_0_28_21_imag,
  output     [15:0]   io_coef_out_payload_0_28_22_real,
  output     [15:0]   io_coef_out_payload_0_28_22_imag,
  output     [15:0]   io_coef_out_payload_0_28_23_real,
  output     [15:0]   io_coef_out_payload_0_28_23_imag,
  output     [15:0]   io_coef_out_payload_0_28_24_real,
  output     [15:0]   io_coef_out_payload_0_28_24_imag,
  output     [15:0]   io_coef_out_payload_0_28_25_real,
  output     [15:0]   io_coef_out_payload_0_28_25_imag,
  output     [15:0]   io_coef_out_payload_0_28_26_real,
  output     [15:0]   io_coef_out_payload_0_28_26_imag,
  output     [15:0]   io_coef_out_payload_0_28_27_real,
  output     [15:0]   io_coef_out_payload_0_28_27_imag,
  output     [15:0]   io_coef_out_payload_0_28_28_real,
  output     [15:0]   io_coef_out_payload_0_28_28_imag,
  output     [15:0]   io_coef_out_payload_0_28_29_real,
  output     [15:0]   io_coef_out_payload_0_28_29_imag,
  output     [15:0]   io_coef_out_payload_0_28_30_real,
  output     [15:0]   io_coef_out_payload_0_28_30_imag,
  output     [15:0]   io_coef_out_payload_0_28_31_real,
  output     [15:0]   io_coef_out_payload_0_28_31_imag,
  output     [15:0]   io_coef_out_payload_0_28_32_real,
  output     [15:0]   io_coef_out_payload_0_28_32_imag,
  output     [15:0]   io_coef_out_payload_0_28_33_real,
  output     [15:0]   io_coef_out_payload_0_28_33_imag,
  output     [15:0]   io_coef_out_payload_0_28_34_real,
  output     [15:0]   io_coef_out_payload_0_28_34_imag,
  output     [15:0]   io_coef_out_payload_0_28_35_real,
  output     [15:0]   io_coef_out_payload_0_28_35_imag,
  output     [15:0]   io_coef_out_payload_0_28_36_real,
  output     [15:0]   io_coef_out_payload_0_28_36_imag,
  output     [15:0]   io_coef_out_payload_0_28_37_real,
  output     [15:0]   io_coef_out_payload_0_28_37_imag,
  output     [15:0]   io_coef_out_payload_0_28_38_real,
  output     [15:0]   io_coef_out_payload_0_28_38_imag,
  output     [15:0]   io_coef_out_payload_0_28_39_real,
  output     [15:0]   io_coef_out_payload_0_28_39_imag,
  output     [15:0]   io_coef_out_payload_0_28_40_real,
  output     [15:0]   io_coef_out_payload_0_28_40_imag,
  output     [15:0]   io_coef_out_payload_0_28_41_real,
  output     [15:0]   io_coef_out_payload_0_28_41_imag,
  output     [15:0]   io_coef_out_payload_0_28_42_real,
  output     [15:0]   io_coef_out_payload_0_28_42_imag,
  output     [15:0]   io_coef_out_payload_0_28_43_real,
  output     [15:0]   io_coef_out_payload_0_28_43_imag,
  output     [15:0]   io_coef_out_payload_0_28_44_real,
  output     [15:0]   io_coef_out_payload_0_28_44_imag,
  output     [15:0]   io_coef_out_payload_0_28_45_real,
  output     [15:0]   io_coef_out_payload_0_28_45_imag,
  output     [15:0]   io_coef_out_payload_0_28_46_real,
  output     [15:0]   io_coef_out_payload_0_28_46_imag,
  output     [15:0]   io_coef_out_payload_0_28_47_real,
  output     [15:0]   io_coef_out_payload_0_28_47_imag,
  output     [15:0]   io_coef_out_payload_0_28_48_real,
  output     [15:0]   io_coef_out_payload_0_28_48_imag,
  output     [15:0]   io_coef_out_payload_0_28_49_real,
  output     [15:0]   io_coef_out_payload_0_28_49_imag,
  output     [15:0]   io_coef_out_payload_0_29_0_real,
  output     [15:0]   io_coef_out_payload_0_29_0_imag,
  output     [15:0]   io_coef_out_payload_0_29_1_real,
  output     [15:0]   io_coef_out_payload_0_29_1_imag,
  output     [15:0]   io_coef_out_payload_0_29_2_real,
  output     [15:0]   io_coef_out_payload_0_29_2_imag,
  output     [15:0]   io_coef_out_payload_0_29_3_real,
  output     [15:0]   io_coef_out_payload_0_29_3_imag,
  output     [15:0]   io_coef_out_payload_0_29_4_real,
  output     [15:0]   io_coef_out_payload_0_29_4_imag,
  output     [15:0]   io_coef_out_payload_0_29_5_real,
  output     [15:0]   io_coef_out_payload_0_29_5_imag,
  output     [15:0]   io_coef_out_payload_0_29_6_real,
  output     [15:0]   io_coef_out_payload_0_29_6_imag,
  output     [15:0]   io_coef_out_payload_0_29_7_real,
  output     [15:0]   io_coef_out_payload_0_29_7_imag,
  output     [15:0]   io_coef_out_payload_0_29_8_real,
  output     [15:0]   io_coef_out_payload_0_29_8_imag,
  output     [15:0]   io_coef_out_payload_0_29_9_real,
  output     [15:0]   io_coef_out_payload_0_29_9_imag,
  output     [15:0]   io_coef_out_payload_0_29_10_real,
  output     [15:0]   io_coef_out_payload_0_29_10_imag,
  output     [15:0]   io_coef_out_payload_0_29_11_real,
  output     [15:0]   io_coef_out_payload_0_29_11_imag,
  output     [15:0]   io_coef_out_payload_0_29_12_real,
  output     [15:0]   io_coef_out_payload_0_29_12_imag,
  output     [15:0]   io_coef_out_payload_0_29_13_real,
  output     [15:0]   io_coef_out_payload_0_29_13_imag,
  output     [15:0]   io_coef_out_payload_0_29_14_real,
  output     [15:0]   io_coef_out_payload_0_29_14_imag,
  output     [15:0]   io_coef_out_payload_0_29_15_real,
  output     [15:0]   io_coef_out_payload_0_29_15_imag,
  output     [15:0]   io_coef_out_payload_0_29_16_real,
  output     [15:0]   io_coef_out_payload_0_29_16_imag,
  output     [15:0]   io_coef_out_payload_0_29_17_real,
  output     [15:0]   io_coef_out_payload_0_29_17_imag,
  output     [15:0]   io_coef_out_payload_0_29_18_real,
  output     [15:0]   io_coef_out_payload_0_29_18_imag,
  output     [15:0]   io_coef_out_payload_0_29_19_real,
  output     [15:0]   io_coef_out_payload_0_29_19_imag,
  output     [15:0]   io_coef_out_payload_0_29_20_real,
  output     [15:0]   io_coef_out_payload_0_29_20_imag,
  output     [15:0]   io_coef_out_payload_0_29_21_real,
  output     [15:0]   io_coef_out_payload_0_29_21_imag,
  output     [15:0]   io_coef_out_payload_0_29_22_real,
  output     [15:0]   io_coef_out_payload_0_29_22_imag,
  output     [15:0]   io_coef_out_payload_0_29_23_real,
  output     [15:0]   io_coef_out_payload_0_29_23_imag,
  output     [15:0]   io_coef_out_payload_0_29_24_real,
  output     [15:0]   io_coef_out_payload_0_29_24_imag,
  output     [15:0]   io_coef_out_payload_0_29_25_real,
  output     [15:0]   io_coef_out_payload_0_29_25_imag,
  output     [15:0]   io_coef_out_payload_0_29_26_real,
  output     [15:0]   io_coef_out_payload_0_29_26_imag,
  output     [15:0]   io_coef_out_payload_0_29_27_real,
  output     [15:0]   io_coef_out_payload_0_29_27_imag,
  output     [15:0]   io_coef_out_payload_0_29_28_real,
  output     [15:0]   io_coef_out_payload_0_29_28_imag,
  output     [15:0]   io_coef_out_payload_0_29_29_real,
  output     [15:0]   io_coef_out_payload_0_29_29_imag,
  output     [15:0]   io_coef_out_payload_0_29_30_real,
  output     [15:0]   io_coef_out_payload_0_29_30_imag,
  output     [15:0]   io_coef_out_payload_0_29_31_real,
  output     [15:0]   io_coef_out_payload_0_29_31_imag,
  output     [15:0]   io_coef_out_payload_0_29_32_real,
  output     [15:0]   io_coef_out_payload_0_29_32_imag,
  output     [15:0]   io_coef_out_payload_0_29_33_real,
  output     [15:0]   io_coef_out_payload_0_29_33_imag,
  output     [15:0]   io_coef_out_payload_0_29_34_real,
  output     [15:0]   io_coef_out_payload_0_29_34_imag,
  output     [15:0]   io_coef_out_payload_0_29_35_real,
  output     [15:0]   io_coef_out_payload_0_29_35_imag,
  output     [15:0]   io_coef_out_payload_0_29_36_real,
  output     [15:0]   io_coef_out_payload_0_29_36_imag,
  output     [15:0]   io_coef_out_payload_0_29_37_real,
  output     [15:0]   io_coef_out_payload_0_29_37_imag,
  output     [15:0]   io_coef_out_payload_0_29_38_real,
  output     [15:0]   io_coef_out_payload_0_29_38_imag,
  output     [15:0]   io_coef_out_payload_0_29_39_real,
  output     [15:0]   io_coef_out_payload_0_29_39_imag,
  output     [15:0]   io_coef_out_payload_0_29_40_real,
  output     [15:0]   io_coef_out_payload_0_29_40_imag,
  output     [15:0]   io_coef_out_payload_0_29_41_real,
  output     [15:0]   io_coef_out_payload_0_29_41_imag,
  output     [15:0]   io_coef_out_payload_0_29_42_real,
  output     [15:0]   io_coef_out_payload_0_29_42_imag,
  output     [15:0]   io_coef_out_payload_0_29_43_real,
  output     [15:0]   io_coef_out_payload_0_29_43_imag,
  output     [15:0]   io_coef_out_payload_0_29_44_real,
  output     [15:0]   io_coef_out_payload_0_29_44_imag,
  output     [15:0]   io_coef_out_payload_0_29_45_real,
  output     [15:0]   io_coef_out_payload_0_29_45_imag,
  output     [15:0]   io_coef_out_payload_0_29_46_real,
  output     [15:0]   io_coef_out_payload_0_29_46_imag,
  output     [15:0]   io_coef_out_payload_0_29_47_real,
  output     [15:0]   io_coef_out_payload_0_29_47_imag,
  output     [15:0]   io_coef_out_payload_0_29_48_real,
  output     [15:0]   io_coef_out_payload_0_29_48_imag,
  output     [15:0]   io_coef_out_payload_0_29_49_real,
  output     [15:0]   io_coef_out_payload_0_29_49_imag,
  output     [15:0]   io_coef_out_payload_0_30_0_real,
  output     [15:0]   io_coef_out_payload_0_30_0_imag,
  output     [15:0]   io_coef_out_payload_0_30_1_real,
  output     [15:0]   io_coef_out_payload_0_30_1_imag,
  output     [15:0]   io_coef_out_payload_0_30_2_real,
  output     [15:0]   io_coef_out_payload_0_30_2_imag,
  output     [15:0]   io_coef_out_payload_0_30_3_real,
  output     [15:0]   io_coef_out_payload_0_30_3_imag,
  output     [15:0]   io_coef_out_payload_0_30_4_real,
  output     [15:0]   io_coef_out_payload_0_30_4_imag,
  output     [15:0]   io_coef_out_payload_0_30_5_real,
  output     [15:0]   io_coef_out_payload_0_30_5_imag,
  output     [15:0]   io_coef_out_payload_0_30_6_real,
  output     [15:0]   io_coef_out_payload_0_30_6_imag,
  output     [15:0]   io_coef_out_payload_0_30_7_real,
  output     [15:0]   io_coef_out_payload_0_30_7_imag,
  output     [15:0]   io_coef_out_payload_0_30_8_real,
  output     [15:0]   io_coef_out_payload_0_30_8_imag,
  output     [15:0]   io_coef_out_payload_0_30_9_real,
  output     [15:0]   io_coef_out_payload_0_30_9_imag,
  output     [15:0]   io_coef_out_payload_0_30_10_real,
  output     [15:0]   io_coef_out_payload_0_30_10_imag,
  output     [15:0]   io_coef_out_payload_0_30_11_real,
  output     [15:0]   io_coef_out_payload_0_30_11_imag,
  output     [15:0]   io_coef_out_payload_0_30_12_real,
  output     [15:0]   io_coef_out_payload_0_30_12_imag,
  output     [15:0]   io_coef_out_payload_0_30_13_real,
  output     [15:0]   io_coef_out_payload_0_30_13_imag,
  output     [15:0]   io_coef_out_payload_0_30_14_real,
  output     [15:0]   io_coef_out_payload_0_30_14_imag,
  output     [15:0]   io_coef_out_payload_0_30_15_real,
  output     [15:0]   io_coef_out_payload_0_30_15_imag,
  output     [15:0]   io_coef_out_payload_0_30_16_real,
  output     [15:0]   io_coef_out_payload_0_30_16_imag,
  output     [15:0]   io_coef_out_payload_0_30_17_real,
  output     [15:0]   io_coef_out_payload_0_30_17_imag,
  output     [15:0]   io_coef_out_payload_0_30_18_real,
  output     [15:0]   io_coef_out_payload_0_30_18_imag,
  output     [15:0]   io_coef_out_payload_0_30_19_real,
  output     [15:0]   io_coef_out_payload_0_30_19_imag,
  output     [15:0]   io_coef_out_payload_0_30_20_real,
  output     [15:0]   io_coef_out_payload_0_30_20_imag,
  output     [15:0]   io_coef_out_payload_0_30_21_real,
  output     [15:0]   io_coef_out_payload_0_30_21_imag,
  output     [15:0]   io_coef_out_payload_0_30_22_real,
  output     [15:0]   io_coef_out_payload_0_30_22_imag,
  output     [15:0]   io_coef_out_payload_0_30_23_real,
  output     [15:0]   io_coef_out_payload_0_30_23_imag,
  output     [15:0]   io_coef_out_payload_0_30_24_real,
  output     [15:0]   io_coef_out_payload_0_30_24_imag,
  output     [15:0]   io_coef_out_payload_0_30_25_real,
  output     [15:0]   io_coef_out_payload_0_30_25_imag,
  output     [15:0]   io_coef_out_payload_0_30_26_real,
  output     [15:0]   io_coef_out_payload_0_30_26_imag,
  output     [15:0]   io_coef_out_payload_0_30_27_real,
  output     [15:0]   io_coef_out_payload_0_30_27_imag,
  output     [15:0]   io_coef_out_payload_0_30_28_real,
  output     [15:0]   io_coef_out_payload_0_30_28_imag,
  output     [15:0]   io_coef_out_payload_0_30_29_real,
  output     [15:0]   io_coef_out_payload_0_30_29_imag,
  output     [15:0]   io_coef_out_payload_0_30_30_real,
  output     [15:0]   io_coef_out_payload_0_30_30_imag,
  output     [15:0]   io_coef_out_payload_0_30_31_real,
  output     [15:0]   io_coef_out_payload_0_30_31_imag,
  output     [15:0]   io_coef_out_payload_0_30_32_real,
  output     [15:0]   io_coef_out_payload_0_30_32_imag,
  output     [15:0]   io_coef_out_payload_0_30_33_real,
  output     [15:0]   io_coef_out_payload_0_30_33_imag,
  output     [15:0]   io_coef_out_payload_0_30_34_real,
  output     [15:0]   io_coef_out_payload_0_30_34_imag,
  output     [15:0]   io_coef_out_payload_0_30_35_real,
  output     [15:0]   io_coef_out_payload_0_30_35_imag,
  output     [15:0]   io_coef_out_payload_0_30_36_real,
  output     [15:0]   io_coef_out_payload_0_30_36_imag,
  output     [15:0]   io_coef_out_payload_0_30_37_real,
  output     [15:0]   io_coef_out_payload_0_30_37_imag,
  output     [15:0]   io_coef_out_payload_0_30_38_real,
  output     [15:0]   io_coef_out_payload_0_30_38_imag,
  output     [15:0]   io_coef_out_payload_0_30_39_real,
  output     [15:0]   io_coef_out_payload_0_30_39_imag,
  output     [15:0]   io_coef_out_payload_0_30_40_real,
  output     [15:0]   io_coef_out_payload_0_30_40_imag,
  output     [15:0]   io_coef_out_payload_0_30_41_real,
  output     [15:0]   io_coef_out_payload_0_30_41_imag,
  output     [15:0]   io_coef_out_payload_0_30_42_real,
  output     [15:0]   io_coef_out_payload_0_30_42_imag,
  output     [15:0]   io_coef_out_payload_0_30_43_real,
  output     [15:0]   io_coef_out_payload_0_30_43_imag,
  output     [15:0]   io_coef_out_payload_0_30_44_real,
  output     [15:0]   io_coef_out_payload_0_30_44_imag,
  output     [15:0]   io_coef_out_payload_0_30_45_real,
  output     [15:0]   io_coef_out_payload_0_30_45_imag,
  output     [15:0]   io_coef_out_payload_0_30_46_real,
  output     [15:0]   io_coef_out_payload_0_30_46_imag,
  output     [15:0]   io_coef_out_payload_0_30_47_real,
  output     [15:0]   io_coef_out_payload_0_30_47_imag,
  output     [15:0]   io_coef_out_payload_0_30_48_real,
  output     [15:0]   io_coef_out_payload_0_30_48_imag,
  output     [15:0]   io_coef_out_payload_0_30_49_real,
  output     [15:0]   io_coef_out_payload_0_30_49_imag,
  output     [15:0]   io_coef_out_payload_0_31_0_real,
  output     [15:0]   io_coef_out_payload_0_31_0_imag,
  output     [15:0]   io_coef_out_payload_0_31_1_real,
  output     [15:0]   io_coef_out_payload_0_31_1_imag,
  output     [15:0]   io_coef_out_payload_0_31_2_real,
  output     [15:0]   io_coef_out_payload_0_31_2_imag,
  output     [15:0]   io_coef_out_payload_0_31_3_real,
  output     [15:0]   io_coef_out_payload_0_31_3_imag,
  output     [15:0]   io_coef_out_payload_0_31_4_real,
  output     [15:0]   io_coef_out_payload_0_31_4_imag,
  output     [15:0]   io_coef_out_payload_0_31_5_real,
  output     [15:0]   io_coef_out_payload_0_31_5_imag,
  output     [15:0]   io_coef_out_payload_0_31_6_real,
  output     [15:0]   io_coef_out_payload_0_31_6_imag,
  output     [15:0]   io_coef_out_payload_0_31_7_real,
  output     [15:0]   io_coef_out_payload_0_31_7_imag,
  output     [15:0]   io_coef_out_payload_0_31_8_real,
  output     [15:0]   io_coef_out_payload_0_31_8_imag,
  output     [15:0]   io_coef_out_payload_0_31_9_real,
  output     [15:0]   io_coef_out_payload_0_31_9_imag,
  output     [15:0]   io_coef_out_payload_0_31_10_real,
  output     [15:0]   io_coef_out_payload_0_31_10_imag,
  output     [15:0]   io_coef_out_payload_0_31_11_real,
  output     [15:0]   io_coef_out_payload_0_31_11_imag,
  output     [15:0]   io_coef_out_payload_0_31_12_real,
  output     [15:0]   io_coef_out_payload_0_31_12_imag,
  output     [15:0]   io_coef_out_payload_0_31_13_real,
  output     [15:0]   io_coef_out_payload_0_31_13_imag,
  output     [15:0]   io_coef_out_payload_0_31_14_real,
  output     [15:0]   io_coef_out_payload_0_31_14_imag,
  output     [15:0]   io_coef_out_payload_0_31_15_real,
  output     [15:0]   io_coef_out_payload_0_31_15_imag,
  output     [15:0]   io_coef_out_payload_0_31_16_real,
  output     [15:0]   io_coef_out_payload_0_31_16_imag,
  output     [15:0]   io_coef_out_payload_0_31_17_real,
  output     [15:0]   io_coef_out_payload_0_31_17_imag,
  output     [15:0]   io_coef_out_payload_0_31_18_real,
  output     [15:0]   io_coef_out_payload_0_31_18_imag,
  output     [15:0]   io_coef_out_payload_0_31_19_real,
  output     [15:0]   io_coef_out_payload_0_31_19_imag,
  output     [15:0]   io_coef_out_payload_0_31_20_real,
  output     [15:0]   io_coef_out_payload_0_31_20_imag,
  output     [15:0]   io_coef_out_payload_0_31_21_real,
  output     [15:0]   io_coef_out_payload_0_31_21_imag,
  output     [15:0]   io_coef_out_payload_0_31_22_real,
  output     [15:0]   io_coef_out_payload_0_31_22_imag,
  output     [15:0]   io_coef_out_payload_0_31_23_real,
  output     [15:0]   io_coef_out_payload_0_31_23_imag,
  output     [15:0]   io_coef_out_payload_0_31_24_real,
  output     [15:0]   io_coef_out_payload_0_31_24_imag,
  output     [15:0]   io_coef_out_payload_0_31_25_real,
  output     [15:0]   io_coef_out_payload_0_31_25_imag,
  output     [15:0]   io_coef_out_payload_0_31_26_real,
  output     [15:0]   io_coef_out_payload_0_31_26_imag,
  output     [15:0]   io_coef_out_payload_0_31_27_real,
  output     [15:0]   io_coef_out_payload_0_31_27_imag,
  output     [15:0]   io_coef_out_payload_0_31_28_real,
  output     [15:0]   io_coef_out_payload_0_31_28_imag,
  output     [15:0]   io_coef_out_payload_0_31_29_real,
  output     [15:0]   io_coef_out_payload_0_31_29_imag,
  output     [15:0]   io_coef_out_payload_0_31_30_real,
  output     [15:0]   io_coef_out_payload_0_31_30_imag,
  output     [15:0]   io_coef_out_payload_0_31_31_real,
  output     [15:0]   io_coef_out_payload_0_31_31_imag,
  output     [15:0]   io_coef_out_payload_0_31_32_real,
  output     [15:0]   io_coef_out_payload_0_31_32_imag,
  output     [15:0]   io_coef_out_payload_0_31_33_real,
  output     [15:0]   io_coef_out_payload_0_31_33_imag,
  output     [15:0]   io_coef_out_payload_0_31_34_real,
  output     [15:0]   io_coef_out_payload_0_31_34_imag,
  output     [15:0]   io_coef_out_payload_0_31_35_real,
  output     [15:0]   io_coef_out_payload_0_31_35_imag,
  output     [15:0]   io_coef_out_payload_0_31_36_real,
  output     [15:0]   io_coef_out_payload_0_31_36_imag,
  output     [15:0]   io_coef_out_payload_0_31_37_real,
  output     [15:0]   io_coef_out_payload_0_31_37_imag,
  output     [15:0]   io_coef_out_payload_0_31_38_real,
  output     [15:0]   io_coef_out_payload_0_31_38_imag,
  output     [15:0]   io_coef_out_payload_0_31_39_real,
  output     [15:0]   io_coef_out_payload_0_31_39_imag,
  output     [15:0]   io_coef_out_payload_0_31_40_real,
  output     [15:0]   io_coef_out_payload_0_31_40_imag,
  output     [15:0]   io_coef_out_payload_0_31_41_real,
  output     [15:0]   io_coef_out_payload_0_31_41_imag,
  output     [15:0]   io_coef_out_payload_0_31_42_real,
  output     [15:0]   io_coef_out_payload_0_31_42_imag,
  output     [15:0]   io_coef_out_payload_0_31_43_real,
  output     [15:0]   io_coef_out_payload_0_31_43_imag,
  output     [15:0]   io_coef_out_payload_0_31_44_real,
  output     [15:0]   io_coef_out_payload_0_31_44_imag,
  output     [15:0]   io_coef_out_payload_0_31_45_real,
  output     [15:0]   io_coef_out_payload_0_31_45_imag,
  output     [15:0]   io_coef_out_payload_0_31_46_real,
  output     [15:0]   io_coef_out_payload_0_31_46_imag,
  output     [15:0]   io_coef_out_payload_0_31_47_real,
  output     [15:0]   io_coef_out_payload_0_31_47_imag,
  output     [15:0]   io_coef_out_payload_0_31_48_real,
  output     [15:0]   io_coef_out_payload_0_31_48_imag,
  output     [15:0]   io_coef_out_payload_0_31_49_real,
  output     [15:0]   io_coef_out_payload_0_31_49_imag,
  output     [15:0]   io_coef_out_payload_0_32_0_real,
  output     [15:0]   io_coef_out_payload_0_32_0_imag,
  output     [15:0]   io_coef_out_payload_0_32_1_real,
  output     [15:0]   io_coef_out_payload_0_32_1_imag,
  output     [15:0]   io_coef_out_payload_0_32_2_real,
  output     [15:0]   io_coef_out_payload_0_32_2_imag,
  output     [15:0]   io_coef_out_payload_0_32_3_real,
  output     [15:0]   io_coef_out_payload_0_32_3_imag,
  output     [15:0]   io_coef_out_payload_0_32_4_real,
  output     [15:0]   io_coef_out_payload_0_32_4_imag,
  output     [15:0]   io_coef_out_payload_0_32_5_real,
  output     [15:0]   io_coef_out_payload_0_32_5_imag,
  output     [15:0]   io_coef_out_payload_0_32_6_real,
  output     [15:0]   io_coef_out_payload_0_32_6_imag,
  output     [15:0]   io_coef_out_payload_0_32_7_real,
  output     [15:0]   io_coef_out_payload_0_32_7_imag,
  output     [15:0]   io_coef_out_payload_0_32_8_real,
  output     [15:0]   io_coef_out_payload_0_32_8_imag,
  output     [15:0]   io_coef_out_payload_0_32_9_real,
  output     [15:0]   io_coef_out_payload_0_32_9_imag,
  output     [15:0]   io_coef_out_payload_0_32_10_real,
  output     [15:0]   io_coef_out_payload_0_32_10_imag,
  output     [15:0]   io_coef_out_payload_0_32_11_real,
  output     [15:0]   io_coef_out_payload_0_32_11_imag,
  output     [15:0]   io_coef_out_payload_0_32_12_real,
  output     [15:0]   io_coef_out_payload_0_32_12_imag,
  output     [15:0]   io_coef_out_payload_0_32_13_real,
  output     [15:0]   io_coef_out_payload_0_32_13_imag,
  output     [15:0]   io_coef_out_payload_0_32_14_real,
  output     [15:0]   io_coef_out_payload_0_32_14_imag,
  output     [15:0]   io_coef_out_payload_0_32_15_real,
  output     [15:0]   io_coef_out_payload_0_32_15_imag,
  output     [15:0]   io_coef_out_payload_0_32_16_real,
  output     [15:0]   io_coef_out_payload_0_32_16_imag,
  output     [15:0]   io_coef_out_payload_0_32_17_real,
  output     [15:0]   io_coef_out_payload_0_32_17_imag,
  output     [15:0]   io_coef_out_payload_0_32_18_real,
  output     [15:0]   io_coef_out_payload_0_32_18_imag,
  output     [15:0]   io_coef_out_payload_0_32_19_real,
  output     [15:0]   io_coef_out_payload_0_32_19_imag,
  output     [15:0]   io_coef_out_payload_0_32_20_real,
  output     [15:0]   io_coef_out_payload_0_32_20_imag,
  output     [15:0]   io_coef_out_payload_0_32_21_real,
  output     [15:0]   io_coef_out_payload_0_32_21_imag,
  output     [15:0]   io_coef_out_payload_0_32_22_real,
  output     [15:0]   io_coef_out_payload_0_32_22_imag,
  output     [15:0]   io_coef_out_payload_0_32_23_real,
  output     [15:0]   io_coef_out_payload_0_32_23_imag,
  output     [15:0]   io_coef_out_payload_0_32_24_real,
  output     [15:0]   io_coef_out_payload_0_32_24_imag,
  output     [15:0]   io_coef_out_payload_0_32_25_real,
  output     [15:0]   io_coef_out_payload_0_32_25_imag,
  output     [15:0]   io_coef_out_payload_0_32_26_real,
  output     [15:0]   io_coef_out_payload_0_32_26_imag,
  output     [15:0]   io_coef_out_payload_0_32_27_real,
  output     [15:0]   io_coef_out_payload_0_32_27_imag,
  output     [15:0]   io_coef_out_payload_0_32_28_real,
  output     [15:0]   io_coef_out_payload_0_32_28_imag,
  output     [15:0]   io_coef_out_payload_0_32_29_real,
  output     [15:0]   io_coef_out_payload_0_32_29_imag,
  output     [15:0]   io_coef_out_payload_0_32_30_real,
  output     [15:0]   io_coef_out_payload_0_32_30_imag,
  output     [15:0]   io_coef_out_payload_0_32_31_real,
  output     [15:0]   io_coef_out_payload_0_32_31_imag,
  output     [15:0]   io_coef_out_payload_0_32_32_real,
  output     [15:0]   io_coef_out_payload_0_32_32_imag,
  output     [15:0]   io_coef_out_payload_0_32_33_real,
  output     [15:0]   io_coef_out_payload_0_32_33_imag,
  output     [15:0]   io_coef_out_payload_0_32_34_real,
  output     [15:0]   io_coef_out_payload_0_32_34_imag,
  output     [15:0]   io_coef_out_payload_0_32_35_real,
  output     [15:0]   io_coef_out_payload_0_32_35_imag,
  output     [15:0]   io_coef_out_payload_0_32_36_real,
  output     [15:0]   io_coef_out_payload_0_32_36_imag,
  output     [15:0]   io_coef_out_payload_0_32_37_real,
  output     [15:0]   io_coef_out_payload_0_32_37_imag,
  output     [15:0]   io_coef_out_payload_0_32_38_real,
  output     [15:0]   io_coef_out_payload_0_32_38_imag,
  output     [15:0]   io_coef_out_payload_0_32_39_real,
  output     [15:0]   io_coef_out_payload_0_32_39_imag,
  output     [15:0]   io_coef_out_payload_0_32_40_real,
  output     [15:0]   io_coef_out_payload_0_32_40_imag,
  output     [15:0]   io_coef_out_payload_0_32_41_real,
  output     [15:0]   io_coef_out_payload_0_32_41_imag,
  output     [15:0]   io_coef_out_payload_0_32_42_real,
  output     [15:0]   io_coef_out_payload_0_32_42_imag,
  output     [15:0]   io_coef_out_payload_0_32_43_real,
  output     [15:0]   io_coef_out_payload_0_32_43_imag,
  output     [15:0]   io_coef_out_payload_0_32_44_real,
  output     [15:0]   io_coef_out_payload_0_32_44_imag,
  output     [15:0]   io_coef_out_payload_0_32_45_real,
  output     [15:0]   io_coef_out_payload_0_32_45_imag,
  output     [15:0]   io_coef_out_payload_0_32_46_real,
  output     [15:0]   io_coef_out_payload_0_32_46_imag,
  output     [15:0]   io_coef_out_payload_0_32_47_real,
  output     [15:0]   io_coef_out_payload_0_32_47_imag,
  output     [15:0]   io_coef_out_payload_0_32_48_real,
  output     [15:0]   io_coef_out_payload_0_32_48_imag,
  output     [15:0]   io_coef_out_payload_0_32_49_real,
  output     [15:0]   io_coef_out_payload_0_32_49_imag,
  output     [15:0]   io_coef_out_payload_0_33_0_real,
  output     [15:0]   io_coef_out_payload_0_33_0_imag,
  output     [15:0]   io_coef_out_payload_0_33_1_real,
  output     [15:0]   io_coef_out_payload_0_33_1_imag,
  output     [15:0]   io_coef_out_payload_0_33_2_real,
  output     [15:0]   io_coef_out_payload_0_33_2_imag,
  output     [15:0]   io_coef_out_payload_0_33_3_real,
  output     [15:0]   io_coef_out_payload_0_33_3_imag,
  output     [15:0]   io_coef_out_payload_0_33_4_real,
  output     [15:0]   io_coef_out_payload_0_33_4_imag,
  output     [15:0]   io_coef_out_payload_0_33_5_real,
  output     [15:0]   io_coef_out_payload_0_33_5_imag,
  output     [15:0]   io_coef_out_payload_0_33_6_real,
  output     [15:0]   io_coef_out_payload_0_33_6_imag,
  output     [15:0]   io_coef_out_payload_0_33_7_real,
  output     [15:0]   io_coef_out_payload_0_33_7_imag,
  output     [15:0]   io_coef_out_payload_0_33_8_real,
  output     [15:0]   io_coef_out_payload_0_33_8_imag,
  output     [15:0]   io_coef_out_payload_0_33_9_real,
  output     [15:0]   io_coef_out_payload_0_33_9_imag,
  output     [15:0]   io_coef_out_payload_0_33_10_real,
  output     [15:0]   io_coef_out_payload_0_33_10_imag,
  output     [15:0]   io_coef_out_payload_0_33_11_real,
  output     [15:0]   io_coef_out_payload_0_33_11_imag,
  output     [15:0]   io_coef_out_payload_0_33_12_real,
  output     [15:0]   io_coef_out_payload_0_33_12_imag,
  output     [15:0]   io_coef_out_payload_0_33_13_real,
  output     [15:0]   io_coef_out_payload_0_33_13_imag,
  output     [15:0]   io_coef_out_payload_0_33_14_real,
  output     [15:0]   io_coef_out_payload_0_33_14_imag,
  output     [15:0]   io_coef_out_payload_0_33_15_real,
  output     [15:0]   io_coef_out_payload_0_33_15_imag,
  output     [15:0]   io_coef_out_payload_0_33_16_real,
  output     [15:0]   io_coef_out_payload_0_33_16_imag,
  output     [15:0]   io_coef_out_payload_0_33_17_real,
  output     [15:0]   io_coef_out_payload_0_33_17_imag,
  output     [15:0]   io_coef_out_payload_0_33_18_real,
  output     [15:0]   io_coef_out_payload_0_33_18_imag,
  output     [15:0]   io_coef_out_payload_0_33_19_real,
  output     [15:0]   io_coef_out_payload_0_33_19_imag,
  output     [15:0]   io_coef_out_payload_0_33_20_real,
  output     [15:0]   io_coef_out_payload_0_33_20_imag,
  output     [15:0]   io_coef_out_payload_0_33_21_real,
  output     [15:0]   io_coef_out_payload_0_33_21_imag,
  output     [15:0]   io_coef_out_payload_0_33_22_real,
  output     [15:0]   io_coef_out_payload_0_33_22_imag,
  output     [15:0]   io_coef_out_payload_0_33_23_real,
  output     [15:0]   io_coef_out_payload_0_33_23_imag,
  output     [15:0]   io_coef_out_payload_0_33_24_real,
  output     [15:0]   io_coef_out_payload_0_33_24_imag,
  output     [15:0]   io_coef_out_payload_0_33_25_real,
  output     [15:0]   io_coef_out_payload_0_33_25_imag,
  output     [15:0]   io_coef_out_payload_0_33_26_real,
  output     [15:0]   io_coef_out_payload_0_33_26_imag,
  output     [15:0]   io_coef_out_payload_0_33_27_real,
  output     [15:0]   io_coef_out_payload_0_33_27_imag,
  output     [15:0]   io_coef_out_payload_0_33_28_real,
  output     [15:0]   io_coef_out_payload_0_33_28_imag,
  output     [15:0]   io_coef_out_payload_0_33_29_real,
  output     [15:0]   io_coef_out_payload_0_33_29_imag,
  output     [15:0]   io_coef_out_payload_0_33_30_real,
  output     [15:0]   io_coef_out_payload_0_33_30_imag,
  output     [15:0]   io_coef_out_payload_0_33_31_real,
  output     [15:0]   io_coef_out_payload_0_33_31_imag,
  output     [15:0]   io_coef_out_payload_0_33_32_real,
  output     [15:0]   io_coef_out_payload_0_33_32_imag,
  output     [15:0]   io_coef_out_payload_0_33_33_real,
  output     [15:0]   io_coef_out_payload_0_33_33_imag,
  output     [15:0]   io_coef_out_payload_0_33_34_real,
  output     [15:0]   io_coef_out_payload_0_33_34_imag,
  output     [15:0]   io_coef_out_payload_0_33_35_real,
  output     [15:0]   io_coef_out_payload_0_33_35_imag,
  output     [15:0]   io_coef_out_payload_0_33_36_real,
  output     [15:0]   io_coef_out_payload_0_33_36_imag,
  output     [15:0]   io_coef_out_payload_0_33_37_real,
  output     [15:0]   io_coef_out_payload_0_33_37_imag,
  output     [15:0]   io_coef_out_payload_0_33_38_real,
  output     [15:0]   io_coef_out_payload_0_33_38_imag,
  output     [15:0]   io_coef_out_payload_0_33_39_real,
  output     [15:0]   io_coef_out_payload_0_33_39_imag,
  output     [15:0]   io_coef_out_payload_0_33_40_real,
  output     [15:0]   io_coef_out_payload_0_33_40_imag,
  output     [15:0]   io_coef_out_payload_0_33_41_real,
  output     [15:0]   io_coef_out_payload_0_33_41_imag,
  output     [15:0]   io_coef_out_payload_0_33_42_real,
  output     [15:0]   io_coef_out_payload_0_33_42_imag,
  output     [15:0]   io_coef_out_payload_0_33_43_real,
  output     [15:0]   io_coef_out_payload_0_33_43_imag,
  output     [15:0]   io_coef_out_payload_0_33_44_real,
  output     [15:0]   io_coef_out_payload_0_33_44_imag,
  output     [15:0]   io_coef_out_payload_0_33_45_real,
  output     [15:0]   io_coef_out_payload_0_33_45_imag,
  output     [15:0]   io_coef_out_payload_0_33_46_real,
  output     [15:0]   io_coef_out_payload_0_33_46_imag,
  output     [15:0]   io_coef_out_payload_0_33_47_real,
  output     [15:0]   io_coef_out_payload_0_33_47_imag,
  output     [15:0]   io_coef_out_payload_0_33_48_real,
  output     [15:0]   io_coef_out_payload_0_33_48_imag,
  output     [15:0]   io_coef_out_payload_0_33_49_real,
  output     [15:0]   io_coef_out_payload_0_33_49_imag,
  output     [15:0]   io_coef_out_payload_0_34_0_real,
  output     [15:0]   io_coef_out_payload_0_34_0_imag,
  output     [15:0]   io_coef_out_payload_0_34_1_real,
  output     [15:0]   io_coef_out_payload_0_34_1_imag,
  output     [15:0]   io_coef_out_payload_0_34_2_real,
  output     [15:0]   io_coef_out_payload_0_34_2_imag,
  output     [15:0]   io_coef_out_payload_0_34_3_real,
  output     [15:0]   io_coef_out_payload_0_34_3_imag,
  output     [15:0]   io_coef_out_payload_0_34_4_real,
  output     [15:0]   io_coef_out_payload_0_34_4_imag,
  output     [15:0]   io_coef_out_payload_0_34_5_real,
  output     [15:0]   io_coef_out_payload_0_34_5_imag,
  output     [15:0]   io_coef_out_payload_0_34_6_real,
  output     [15:0]   io_coef_out_payload_0_34_6_imag,
  output     [15:0]   io_coef_out_payload_0_34_7_real,
  output     [15:0]   io_coef_out_payload_0_34_7_imag,
  output     [15:0]   io_coef_out_payload_0_34_8_real,
  output     [15:0]   io_coef_out_payload_0_34_8_imag,
  output     [15:0]   io_coef_out_payload_0_34_9_real,
  output     [15:0]   io_coef_out_payload_0_34_9_imag,
  output     [15:0]   io_coef_out_payload_0_34_10_real,
  output     [15:0]   io_coef_out_payload_0_34_10_imag,
  output     [15:0]   io_coef_out_payload_0_34_11_real,
  output     [15:0]   io_coef_out_payload_0_34_11_imag,
  output     [15:0]   io_coef_out_payload_0_34_12_real,
  output     [15:0]   io_coef_out_payload_0_34_12_imag,
  output     [15:0]   io_coef_out_payload_0_34_13_real,
  output     [15:0]   io_coef_out_payload_0_34_13_imag,
  output     [15:0]   io_coef_out_payload_0_34_14_real,
  output     [15:0]   io_coef_out_payload_0_34_14_imag,
  output     [15:0]   io_coef_out_payload_0_34_15_real,
  output     [15:0]   io_coef_out_payload_0_34_15_imag,
  output     [15:0]   io_coef_out_payload_0_34_16_real,
  output     [15:0]   io_coef_out_payload_0_34_16_imag,
  output     [15:0]   io_coef_out_payload_0_34_17_real,
  output     [15:0]   io_coef_out_payload_0_34_17_imag,
  output     [15:0]   io_coef_out_payload_0_34_18_real,
  output     [15:0]   io_coef_out_payload_0_34_18_imag,
  output     [15:0]   io_coef_out_payload_0_34_19_real,
  output     [15:0]   io_coef_out_payload_0_34_19_imag,
  output     [15:0]   io_coef_out_payload_0_34_20_real,
  output     [15:0]   io_coef_out_payload_0_34_20_imag,
  output     [15:0]   io_coef_out_payload_0_34_21_real,
  output     [15:0]   io_coef_out_payload_0_34_21_imag,
  output     [15:0]   io_coef_out_payload_0_34_22_real,
  output     [15:0]   io_coef_out_payload_0_34_22_imag,
  output     [15:0]   io_coef_out_payload_0_34_23_real,
  output     [15:0]   io_coef_out_payload_0_34_23_imag,
  output     [15:0]   io_coef_out_payload_0_34_24_real,
  output     [15:0]   io_coef_out_payload_0_34_24_imag,
  output     [15:0]   io_coef_out_payload_0_34_25_real,
  output     [15:0]   io_coef_out_payload_0_34_25_imag,
  output     [15:0]   io_coef_out_payload_0_34_26_real,
  output     [15:0]   io_coef_out_payload_0_34_26_imag,
  output     [15:0]   io_coef_out_payload_0_34_27_real,
  output     [15:0]   io_coef_out_payload_0_34_27_imag,
  output     [15:0]   io_coef_out_payload_0_34_28_real,
  output     [15:0]   io_coef_out_payload_0_34_28_imag,
  output     [15:0]   io_coef_out_payload_0_34_29_real,
  output     [15:0]   io_coef_out_payload_0_34_29_imag,
  output     [15:0]   io_coef_out_payload_0_34_30_real,
  output     [15:0]   io_coef_out_payload_0_34_30_imag,
  output     [15:0]   io_coef_out_payload_0_34_31_real,
  output     [15:0]   io_coef_out_payload_0_34_31_imag,
  output     [15:0]   io_coef_out_payload_0_34_32_real,
  output     [15:0]   io_coef_out_payload_0_34_32_imag,
  output     [15:0]   io_coef_out_payload_0_34_33_real,
  output     [15:0]   io_coef_out_payload_0_34_33_imag,
  output     [15:0]   io_coef_out_payload_0_34_34_real,
  output     [15:0]   io_coef_out_payload_0_34_34_imag,
  output     [15:0]   io_coef_out_payload_0_34_35_real,
  output     [15:0]   io_coef_out_payload_0_34_35_imag,
  output     [15:0]   io_coef_out_payload_0_34_36_real,
  output     [15:0]   io_coef_out_payload_0_34_36_imag,
  output     [15:0]   io_coef_out_payload_0_34_37_real,
  output     [15:0]   io_coef_out_payload_0_34_37_imag,
  output     [15:0]   io_coef_out_payload_0_34_38_real,
  output     [15:0]   io_coef_out_payload_0_34_38_imag,
  output     [15:0]   io_coef_out_payload_0_34_39_real,
  output     [15:0]   io_coef_out_payload_0_34_39_imag,
  output     [15:0]   io_coef_out_payload_0_34_40_real,
  output     [15:0]   io_coef_out_payload_0_34_40_imag,
  output     [15:0]   io_coef_out_payload_0_34_41_real,
  output     [15:0]   io_coef_out_payload_0_34_41_imag,
  output     [15:0]   io_coef_out_payload_0_34_42_real,
  output     [15:0]   io_coef_out_payload_0_34_42_imag,
  output     [15:0]   io_coef_out_payload_0_34_43_real,
  output     [15:0]   io_coef_out_payload_0_34_43_imag,
  output     [15:0]   io_coef_out_payload_0_34_44_real,
  output     [15:0]   io_coef_out_payload_0_34_44_imag,
  output     [15:0]   io_coef_out_payload_0_34_45_real,
  output     [15:0]   io_coef_out_payload_0_34_45_imag,
  output     [15:0]   io_coef_out_payload_0_34_46_real,
  output     [15:0]   io_coef_out_payload_0_34_46_imag,
  output     [15:0]   io_coef_out_payload_0_34_47_real,
  output     [15:0]   io_coef_out_payload_0_34_47_imag,
  output     [15:0]   io_coef_out_payload_0_34_48_real,
  output     [15:0]   io_coef_out_payload_0_34_48_imag,
  output     [15:0]   io_coef_out_payload_0_34_49_real,
  output     [15:0]   io_coef_out_payload_0_34_49_imag,
  output     [15:0]   io_coef_out_payload_0_35_0_real,
  output     [15:0]   io_coef_out_payload_0_35_0_imag,
  output     [15:0]   io_coef_out_payload_0_35_1_real,
  output     [15:0]   io_coef_out_payload_0_35_1_imag,
  output     [15:0]   io_coef_out_payload_0_35_2_real,
  output     [15:0]   io_coef_out_payload_0_35_2_imag,
  output     [15:0]   io_coef_out_payload_0_35_3_real,
  output     [15:0]   io_coef_out_payload_0_35_3_imag,
  output     [15:0]   io_coef_out_payload_0_35_4_real,
  output     [15:0]   io_coef_out_payload_0_35_4_imag,
  output     [15:0]   io_coef_out_payload_0_35_5_real,
  output     [15:0]   io_coef_out_payload_0_35_5_imag,
  output     [15:0]   io_coef_out_payload_0_35_6_real,
  output     [15:0]   io_coef_out_payload_0_35_6_imag,
  output     [15:0]   io_coef_out_payload_0_35_7_real,
  output     [15:0]   io_coef_out_payload_0_35_7_imag,
  output     [15:0]   io_coef_out_payload_0_35_8_real,
  output     [15:0]   io_coef_out_payload_0_35_8_imag,
  output     [15:0]   io_coef_out_payload_0_35_9_real,
  output     [15:0]   io_coef_out_payload_0_35_9_imag,
  output     [15:0]   io_coef_out_payload_0_35_10_real,
  output     [15:0]   io_coef_out_payload_0_35_10_imag,
  output     [15:0]   io_coef_out_payload_0_35_11_real,
  output     [15:0]   io_coef_out_payload_0_35_11_imag,
  output     [15:0]   io_coef_out_payload_0_35_12_real,
  output     [15:0]   io_coef_out_payload_0_35_12_imag,
  output     [15:0]   io_coef_out_payload_0_35_13_real,
  output     [15:0]   io_coef_out_payload_0_35_13_imag,
  output     [15:0]   io_coef_out_payload_0_35_14_real,
  output     [15:0]   io_coef_out_payload_0_35_14_imag,
  output     [15:0]   io_coef_out_payload_0_35_15_real,
  output     [15:0]   io_coef_out_payload_0_35_15_imag,
  output     [15:0]   io_coef_out_payload_0_35_16_real,
  output     [15:0]   io_coef_out_payload_0_35_16_imag,
  output     [15:0]   io_coef_out_payload_0_35_17_real,
  output     [15:0]   io_coef_out_payload_0_35_17_imag,
  output     [15:0]   io_coef_out_payload_0_35_18_real,
  output     [15:0]   io_coef_out_payload_0_35_18_imag,
  output     [15:0]   io_coef_out_payload_0_35_19_real,
  output     [15:0]   io_coef_out_payload_0_35_19_imag,
  output     [15:0]   io_coef_out_payload_0_35_20_real,
  output     [15:0]   io_coef_out_payload_0_35_20_imag,
  output     [15:0]   io_coef_out_payload_0_35_21_real,
  output     [15:0]   io_coef_out_payload_0_35_21_imag,
  output     [15:0]   io_coef_out_payload_0_35_22_real,
  output     [15:0]   io_coef_out_payload_0_35_22_imag,
  output     [15:0]   io_coef_out_payload_0_35_23_real,
  output     [15:0]   io_coef_out_payload_0_35_23_imag,
  output     [15:0]   io_coef_out_payload_0_35_24_real,
  output     [15:0]   io_coef_out_payload_0_35_24_imag,
  output     [15:0]   io_coef_out_payload_0_35_25_real,
  output     [15:0]   io_coef_out_payload_0_35_25_imag,
  output     [15:0]   io_coef_out_payload_0_35_26_real,
  output     [15:0]   io_coef_out_payload_0_35_26_imag,
  output     [15:0]   io_coef_out_payload_0_35_27_real,
  output     [15:0]   io_coef_out_payload_0_35_27_imag,
  output     [15:0]   io_coef_out_payload_0_35_28_real,
  output     [15:0]   io_coef_out_payload_0_35_28_imag,
  output     [15:0]   io_coef_out_payload_0_35_29_real,
  output     [15:0]   io_coef_out_payload_0_35_29_imag,
  output     [15:0]   io_coef_out_payload_0_35_30_real,
  output     [15:0]   io_coef_out_payload_0_35_30_imag,
  output     [15:0]   io_coef_out_payload_0_35_31_real,
  output     [15:0]   io_coef_out_payload_0_35_31_imag,
  output     [15:0]   io_coef_out_payload_0_35_32_real,
  output     [15:0]   io_coef_out_payload_0_35_32_imag,
  output     [15:0]   io_coef_out_payload_0_35_33_real,
  output     [15:0]   io_coef_out_payload_0_35_33_imag,
  output     [15:0]   io_coef_out_payload_0_35_34_real,
  output     [15:0]   io_coef_out_payload_0_35_34_imag,
  output     [15:0]   io_coef_out_payload_0_35_35_real,
  output     [15:0]   io_coef_out_payload_0_35_35_imag,
  output     [15:0]   io_coef_out_payload_0_35_36_real,
  output     [15:0]   io_coef_out_payload_0_35_36_imag,
  output     [15:0]   io_coef_out_payload_0_35_37_real,
  output     [15:0]   io_coef_out_payload_0_35_37_imag,
  output     [15:0]   io_coef_out_payload_0_35_38_real,
  output     [15:0]   io_coef_out_payload_0_35_38_imag,
  output     [15:0]   io_coef_out_payload_0_35_39_real,
  output     [15:0]   io_coef_out_payload_0_35_39_imag,
  output     [15:0]   io_coef_out_payload_0_35_40_real,
  output     [15:0]   io_coef_out_payload_0_35_40_imag,
  output     [15:0]   io_coef_out_payload_0_35_41_real,
  output     [15:0]   io_coef_out_payload_0_35_41_imag,
  output     [15:0]   io_coef_out_payload_0_35_42_real,
  output     [15:0]   io_coef_out_payload_0_35_42_imag,
  output     [15:0]   io_coef_out_payload_0_35_43_real,
  output     [15:0]   io_coef_out_payload_0_35_43_imag,
  output     [15:0]   io_coef_out_payload_0_35_44_real,
  output     [15:0]   io_coef_out_payload_0_35_44_imag,
  output     [15:0]   io_coef_out_payload_0_35_45_real,
  output     [15:0]   io_coef_out_payload_0_35_45_imag,
  output     [15:0]   io_coef_out_payload_0_35_46_real,
  output     [15:0]   io_coef_out_payload_0_35_46_imag,
  output     [15:0]   io_coef_out_payload_0_35_47_real,
  output     [15:0]   io_coef_out_payload_0_35_47_imag,
  output     [15:0]   io_coef_out_payload_0_35_48_real,
  output     [15:0]   io_coef_out_payload_0_35_48_imag,
  output     [15:0]   io_coef_out_payload_0_35_49_real,
  output     [15:0]   io_coef_out_payload_0_35_49_imag,
  output     [15:0]   io_coef_out_payload_0_36_0_real,
  output     [15:0]   io_coef_out_payload_0_36_0_imag,
  output     [15:0]   io_coef_out_payload_0_36_1_real,
  output     [15:0]   io_coef_out_payload_0_36_1_imag,
  output     [15:0]   io_coef_out_payload_0_36_2_real,
  output     [15:0]   io_coef_out_payload_0_36_2_imag,
  output     [15:0]   io_coef_out_payload_0_36_3_real,
  output     [15:0]   io_coef_out_payload_0_36_3_imag,
  output     [15:0]   io_coef_out_payload_0_36_4_real,
  output     [15:0]   io_coef_out_payload_0_36_4_imag,
  output     [15:0]   io_coef_out_payload_0_36_5_real,
  output     [15:0]   io_coef_out_payload_0_36_5_imag,
  output     [15:0]   io_coef_out_payload_0_36_6_real,
  output     [15:0]   io_coef_out_payload_0_36_6_imag,
  output     [15:0]   io_coef_out_payload_0_36_7_real,
  output     [15:0]   io_coef_out_payload_0_36_7_imag,
  output     [15:0]   io_coef_out_payload_0_36_8_real,
  output     [15:0]   io_coef_out_payload_0_36_8_imag,
  output     [15:0]   io_coef_out_payload_0_36_9_real,
  output     [15:0]   io_coef_out_payload_0_36_9_imag,
  output     [15:0]   io_coef_out_payload_0_36_10_real,
  output     [15:0]   io_coef_out_payload_0_36_10_imag,
  output     [15:0]   io_coef_out_payload_0_36_11_real,
  output     [15:0]   io_coef_out_payload_0_36_11_imag,
  output     [15:0]   io_coef_out_payload_0_36_12_real,
  output     [15:0]   io_coef_out_payload_0_36_12_imag,
  output     [15:0]   io_coef_out_payload_0_36_13_real,
  output     [15:0]   io_coef_out_payload_0_36_13_imag,
  output     [15:0]   io_coef_out_payload_0_36_14_real,
  output     [15:0]   io_coef_out_payload_0_36_14_imag,
  output     [15:0]   io_coef_out_payload_0_36_15_real,
  output     [15:0]   io_coef_out_payload_0_36_15_imag,
  output     [15:0]   io_coef_out_payload_0_36_16_real,
  output     [15:0]   io_coef_out_payload_0_36_16_imag,
  output     [15:0]   io_coef_out_payload_0_36_17_real,
  output     [15:0]   io_coef_out_payload_0_36_17_imag,
  output     [15:0]   io_coef_out_payload_0_36_18_real,
  output     [15:0]   io_coef_out_payload_0_36_18_imag,
  output     [15:0]   io_coef_out_payload_0_36_19_real,
  output     [15:0]   io_coef_out_payload_0_36_19_imag,
  output     [15:0]   io_coef_out_payload_0_36_20_real,
  output     [15:0]   io_coef_out_payload_0_36_20_imag,
  output     [15:0]   io_coef_out_payload_0_36_21_real,
  output     [15:0]   io_coef_out_payload_0_36_21_imag,
  output     [15:0]   io_coef_out_payload_0_36_22_real,
  output     [15:0]   io_coef_out_payload_0_36_22_imag,
  output     [15:0]   io_coef_out_payload_0_36_23_real,
  output     [15:0]   io_coef_out_payload_0_36_23_imag,
  output     [15:0]   io_coef_out_payload_0_36_24_real,
  output     [15:0]   io_coef_out_payload_0_36_24_imag,
  output     [15:0]   io_coef_out_payload_0_36_25_real,
  output     [15:0]   io_coef_out_payload_0_36_25_imag,
  output     [15:0]   io_coef_out_payload_0_36_26_real,
  output     [15:0]   io_coef_out_payload_0_36_26_imag,
  output     [15:0]   io_coef_out_payload_0_36_27_real,
  output     [15:0]   io_coef_out_payload_0_36_27_imag,
  output     [15:0]   io_coef_out_payload_0_36_28_real,
  output     [15:0]   io_coef_out_payload_0_36_28_imag,
  output     [15:0]   io_coef_out_payload_0_36_29_real,
  output     [15:0]   io_coef_out_payload_0_36_29_imag,
  output     [15:0]   io_coef_out_payload_0_36_30_real,
  output     [15:0]   io_coef_out_payload_0_36_30_imag,
  output     [15:0]   io_coef_out_payload_0_36_31_real,
  output     [15:0]   io_coef_out_payload_0_36_31_imag,
  output     [15:0]   io_coef_out_payload_0_36_32_real,
  output     [15:0]   io_coef_out_payload_0_36_32_imag,
  output     [15:0]   io_coef_out_payload_0_36_33_real,
  output     [15:0]   io_coef_out_payload_0_36_33_imag,
  output     [15:0]   io_coef_out_payload_0_36_34_real,
  output     [15:0]   io_coef_out_payload_0_36_34_imag,
  output     [15:0]   io_coef_out_payload_0_36_35_real,
  output     [15:0]   io_coef_out_payload_0_36_35_imag,
  output     [15:0]   io_coef_out_payload_0_36_36_real,
  output     [15:0]   io_coef_out_payload_0_36_36_imag,
  output     [15:0]   io_coef_out_payload_0_36_37_real,
  output     [15:0]   io_coef_out_payload_0_36_37_imag,
  output     [15:0]   io_coef_out_payload_0_36_38_real,
  output     [15:0]   io_coef_out_payload_0_36_38_imag,
  output     [15:0]   io_coef_out_payload_0_36_39_real,
  output     [15:0]   io_coef_out_payload_0_36_39_imag,
  output     [15:0]   io_coef_out_payload_0_36_40_real,
  output     [15:0]   io_coef_out_payload_0_36_40_imag,
  output     [15:0]   io_coef_out_payload_0_36_41_real,
  output     [15:0]   io_coef_out_payload_0_36_41_imag,
  output     [15:0]   io_coef_out_payload_0_36_42_real,
  output     [15:0]   io_coef_out_payload_0_36_42_imag,
  output     [15:0]   io_coef_out_payload_0_36_43_real,
  output     [15:0]   io_coef_out_payload_0_36_43_imag,
  output     [15:0]   io_coef_out_payload_0_36_44_real,
  output     [15:0]   io_coef_out_payload_0_36_44_imag,
  output     [15:0]   io_coef_out_payload_0_36_45_real,
  output     [15:0]   io_coef_out_payload_0_36_45_imag,
  output     [15:0]   io_coef_out_payload_0_36_46_real,
  output     [15:0]   io_coef_out_payload_0_36_46_imag,
  output     [15:0]   io_coef_out_payload_0_36_47_real,
  output     [15:0]   io_coef_out_payload_0_36_47_imag,
  output     [15:0]   io_coef_out_payload_0_36_48_real,
  output     [15:0]   io_coef_out_payload_0_36_48_imag,
  output     [15:0]   io_coef_out_payload_0_36_49_real,
  output     [15:0]   io_coef_out_payload_0_36_49_imag,
  output     [15:0]   io_coef_out_payload_0_37_0_real,
  output     [15:0]   io_coef_out_payload_0_37_0_imag,
  output     [15:0]   io_coef_out_payload_0_37_1_real,
  output     [15:0]   io_coef_out_payload_0_37_1_imag,
  output     [15:0]   io_coef_out_payload_0_37_2_real,
  output     [15:0]   io_coef_out_payload_0_37_2_imag,
  output     [15:0]   io_coef_out_payload_0_37_3_real,
  output     [15:0]   io_coef_out_payload_0_37_3_imag,
  output     [15:0]   io_coef_out_payload_0_37_4_real,
  output     [15:0]   io_coef_out_payload_0_37_4_imag,
  output     [15:0]   io_coef_out_payload_0_37_5_real,
  output     [15:0]   io_coef_out_payload_0_37_5_imag,
  output     [15:0]   io_coef_out_payload_0_37_6_real,
  output     [15:0]   io_coef_out_payload_0_37_6_imag,
  output     [15:0]   io_coef_out_payload_0_37_7_real,
  output     [15:0]   io_coef_out_payload_0_37_7_imag,
  output     [15:0]   io_coef_out_payload_0_37_8_real,
  output     [15:0]   io_coef_out_payload_0_37_8_imag,
  output     [15:0]   io_coef_out_payload_0_37_9_real,
  output     [15:0]   io_coef_out_payload_0_37_9_imag,
  output     [15:0]   io_coef_out_payload_0_37_10_real,
  output     [15:0]   io_coef_out_payload_0_37_10_imag,
  output     [15:0]   io_coef_out_payload_0_37_11_real,
  output     [15:0]   io_coef_out_payload_0_37_11_imag,
  output     [15:0]   io_coef_out_payload_0_37_12_real,
  output     [15:0]   io_coef_out_payload_0_37_12_imag,
  output     [15:0]   io_coef_out_payload_0_37_13_real,
  output     [15:0]   io_coef_out_payload_0_37_13_imag,
  output     [15:0]   io_coef_out_payload_0_37_14_real,
  output     [15:0]   io_coef_out_payload_0_37_14_imag,
  output     [15:0]   io_coef_out_payload_0_37_15_real,
  output     [15:0]   io_coef_out_payload_0_37_15_imag,
  output     [15:0]   io_coef_out_payload_0_37_16_real,
  output     [15:0]   io_coef_out_payload_0_37_16_imag,
  output     [15:0]   io_coef_out_payload_0_37_17_real,
  output     [15:0]   io_coef_out_payload_0_37_17_imag,
  output     [15:0]   io_coef_out_payload_0_37_18_real,
  output     [15:0]   io_coef_out_payload_0_37_18_imag,
  output     [15:0]   io_coef_out_payload_0_37_19_real,
  output     [15:0]   io_coef_out_payload_0_37_19_imag,
  output     [15:0]   io_coef_out_payload_0_37_20_real,
  output     [15:0]   io_coef_out_payload_0_37_20_imag,
  output     [15:0]   io_coef_out_payload_0_37_21_real,
  output     [15:0]   io_coef_out_payload_0_37_21_imag,
  output     [15:0]   io_coef_out_payload_0_37_22_real,
  output     [15:0]   io_coef_out_payload_0_37_22_imag,
  output     [15:0]   io_coef_out_payload_0_37_23_real,
  output     [15:0]   io_coef_out_payload_0_37_23_imag,
  output     [15:0]   io_coef_out_payload_0_37_24_real,
  output     [15:0]   io_coef_out_payload_0_37_24_imag,
  output     [15:0]   io_coef_out_payload_0_37_25_real,
  output     [15:0]   io_coef_out_payload_0_37_25_imag,
  output     [15:0]   io_coef_out_payload_0_37_26_real,
  output     [15:0]   io_coef_out_payload_0_37_26_imag,
  output     [15:0]   io_coef_out_payload_0_37_27_real,
  output     [15:0]   io_coef_out_payload_0_37_27_imag,
  output     [15:0]   io_coef_out_payload_0_37_28_real,
  output     [15:0]   io_coef_out_payload_0_37_28_imag,
  output     [15:0]   io_coef_out_payload_0_37_29_real,
  output     [15:0]   io_coef_out_payload_0_37_29_imag,
  output     [15:0]   io_coef_out_payload_0_37_30_real,
  output     [15:0]   io_coef_out_payload_0_37_30_imag,
  output     [15:0]   io_coef_out_payload_0_37_31_real,
  output     [15:0]   io_coef_out_payload_0_37_31_imag,
  output     [15:0]   io_coef_out_payload_0_37_32_real,
  output     [15:0]   io_coef_out_payload_0_37_32_imag,
  output     [15:0]   io_coef_out_payload_0_37_33_real,
  output     [15:0]   io_coef_out_payload_0_37_33_imag,
  output     [15:0]   io_coef_out_payload_0_37_34_real,
  output     [15:0]   io_coef_out_payload_0_37_34_imag,
  output     [15:0]   io_coef_out_payload_0_37_35_real,
  output     [15:0]   io_coef_out_payload_0_37_35_imag,
  output     [15:0]   io_coef_out_payload_0_37_36_real,
  output     [15:0]   io_coef_out_payload_0_37_36_imag,
  output     [15:0]   io_coef_out_payload_0_37_37_real,
  output     [15:0]   io_coef_out_payload_0_37_37_imag,
  output     [15:0]   io_coef_out_payload_0_37_38_real,
  output     [15:0]   io_coef_out_payload_0_37_38_imag,
  output     [15:0]   io_coef_out_payload_0_37_39_real,
  output     [15:0]   io_coef_out_payload_0_37_39_imag,
  output     [15:0]   io_coef_out_payload_0_37_40_real,
  output     [15:0]   io_coef_out_payload_0_37_40_imag,
  output     [15:0]   io_coef_out_payload_0_37_41_real,
  output     [15:0]   io_coef_out_payload_0_37_41_imag,
  output     [15:0]   io_coef_out_payload_0_37_42_real,
  output     [15:0]   io_coef_out_payload_0_37_42_imag,
  output     [15:0]   io_coef_out_payload_0_37_43_real,
  output     [15:0]   io_coef_out_payload_0_37_43_imag,
  output     [15:0]   io_coef_out_payload_0_37_44_real,
  output     [15:0]   io_coef_out_payload_0_37_44_imag,
  output     [15:0]   io_coef_out_payload_0_37_45_real,
  output     [15:0]   io_coef_out_payload_0_37_45_imag,
  output     [15:0]   io_coef_out_payload_0_37_46_real,
  output     [15:0]   io_coef_out_payload_0_37_46_imag,
  output     [15:0]   io_coef_out_payload_0_37_47_real,
  output     [15:0]   io_coef_out_payload_0_37_47_imag,
  output     [15:0]   io_coef_out_payload_0_37_48_real,
  output     [15:0]   io_coef_out_payload_0_37_48_imag,
  output     [15:0]   io_coef_out_payload_0_37_49_real,
  output     [15:0]   io_coef_out_payload_0_37_49_imag,
  output     [15:0]   io_coef_out_payload_0_38_0_real,
  output     [15:0]   io_coef_out_payload_0_38_0_imag,
  output     [15:0]   io_coef_out_payload_0_38_1_real,
  output     [15:0]   io_coef_out_payload_0_38_1_imag,
  output     [15:0]   io_coef_out_payload_0_38_2_real,
  output     [15:0]   io_coef_out_payload_0_38_2_imag,
  output     [15:0]   io_coef_out_payload_0_38_3_real,
  output     [15:0]   io_coef_out_payload_0_38_3_imag,
  output     [15:0]   io_coef_out_payload_0_38_4_real,
  output     [15:0]   io_coef_out_payload_0_38_4_imag,
  output     [15:0]   io_coef_out_payload_0_38_5_real,
  output     [15:0]   io_coef_out_payload_0_38_5_imag,
  output     [15:0]   io_coef_out_payload_0_38_6_real,
  output     [15:0]   io_coef_out_payload_0_38_6_imag,
  output     [15:0]   io_coef_out_payload_0_38_7_real,
  output     [15:0]   io_coef_out_payload_0_38_7_imag,
  output     [15:0]   io_coef_out_payload_0_38_8_real,
  output     [15:0]   io_coef_out_payload_0_38_8_imag,
  output     [15:0]   io_coef_out_payload_0_38_9_real,
  output     [15:0]   io_coef_out_payload_0_38_9_imag,
  output     [15:0]   io_coef_out_payload_0_38_10_real,
  output     [15:0]   io_coef_out_payload_0_38_10_imag,
  output     [15:0]   io_coef_out_payload_0_38_11_real,
  output     [15:0]   io_coef_out_payload_0_38_11_imag,
  output     [15:0]   io_coef_out_payload_0_38_12_real,
  output     [15:0]   io_coef_out_payload_0_38_12_imag,
  output     [15:0]   io_coef_out_payload_0_38_13_real,
  output     [15:0]   io_coef_out_payload_0_38_13_imag,
  output     [15:0]   io_coef_out_payload_0_38_14_real,
  output     [15:0]   io_coef_out_payload_0_38_14_imag,
  output     [15:0]   io_coef_out_payload_0_38_15_real,
  output     [15:0]   io_coef_out_payload_0_38_15_imag,
  output     [15:0]   io_coef_out_payload_0_38_16_real,
  output     [15:0]   io_coef_out_payload_0_38_16_imag,
  output     [15:0]   io_coef_out_payload_0_38_17_real,
  output     [15:0]   io_coef_out_payload_0_38_17_imag,
  output     [15:0]   io_coef_out_payload_0_38_18_real,
  output     [15:0]   io_coef_out_payload_0_38_18_imag,
  output     [15:0]   io_coef_out_payload_0_38_19_real,
  output     [15:0]   io_coef_out_payload_0_38_19_imag,
  output     [15:0]   io_coef_out_payload_0_38_20_real,
  output     [15:0]   io_coef_out_payload_0_38_20_imag,
  output     [15:0]   io_coef_out_payload_0_38_21_real,
  output     [15:0]   io_coef_out_payload_0_38_21_imag,
  output     [15:0]   io_coef_out_payload_0_38_22_real,
  output     [15:0]   io_coef_out_payload_0_38_22_imag,
  output     [15:0]   io_coef_out_payload_0_38_23_real,
  output     [15:0]   io_coef_out_payload_0_38_23_imag,
  output     [15:0]   io_coef_out_payload_0_38_24_real,
  output     [15:0]   io_coef_out_payload_0_38_24_imag,
  output     [15:0]   io_coef_out_payload_0_38_25_real,
  output     [15:0]   io_coef_out_payload_0_38_25_imag,
  output     [15:0]   io_coef_out_payload_0_38_26_real,
  output     [15:0]   io_coef_out_payload_0_38_26_imag,
  output     [15:0]   io_coef_out_payload_0_38_27_real,
  output     [15:0]   io_coef_out_payload_0_38_27_imag,
  output     [15:0]   io_coef_out_payload_0_38_28_real,
  output     [15:0]   io_coef_out_payload_0_38_28_imag,
  output     [15:0]   io_coef_out_payload_0_38_29_real,
  output     [15:0]   io_coef_out_payload_0_38_29_imag,
  output     [15:0]   io_coef_out_payload_0_38_30_real,
  output     [15:0]   io_coef_out_payload_0_38_30_imag,
  output     [15:0]   io_coef_out_payload_0_38_31_real,
  output     [15:0]   io_coef_out_payload_0_38_31_imag,
  output     [15:0]   io_coef_out_payload_0_38_32_real,
  output     [15:0]   io_coef_out_payload_0_38_32_imag,
  output     [15:0]   io_coef_out_payload_0_38_33_real,
  output     [15:0]   io_coef_out_payload_0_38_33_imag,
  output     [15:0]   io_coef_out_payload_0_38_34_real,
  output     [15:0]   io_coef_out_payload_0_38_34_imag,
  output     [15:0]   io_coef_out_payload_0_38_35_real,
  output     [15:0]   io_coef_out_payload_0_38_35_imag,
  output     [15:0]   io_coef_out_payload_0_38_36_real,
  output     [15:0]   io_coef_out_payload_0_38_36_imag,
  output     [15:0]   io_coef_out_payload_0_38_37_real,
  output     [15:0]   io_coef_out_payload_0_38_37_imag,
  output     [15:0]   io_coef_out_payload_0_38_38_real,
  output     [15:0]   io_coef_out_payload_0_38_38_imag,
  output     [15:0]   io_coef_out_payload_0_38_39_real,
  output     [15:0]   io_coef_out_payload_0_38_39_imag,
  output     [15:0]   io_coef_out_payload_0_38_40_real,
  output     [15:0]   io_coef_out_payload_0_38_40_imag,
  output     [15:0]   io_coef_out_payload_0_38_41_real,
  output     [15:0]   io_coef_out_payload_0_38_41_imag,
  output     [15:0]   io_coef_out_payload_0_38_42_real,
  output     [15:0]   io_coef_out_payload_0_38_42_imag,
  output     [15:0]   io_coef_out_payload_0_38_43_real,
  output     [15:0]   io_coef_out_payload_0_38_43_imag,
  output     [15:0]   io_coef_out_payload_0_38_44_real,
  output     [15:0]   io_coef_out_payload_0_38_44_imag,
  output     [15:0]   io_coef_out_payload_0_38_45_real,
  output     [15:0]   io_coef_out_payload_0_38_45_imag,
  output     [15:0]   io_coef_out_payload_0_38_46_real,
  output     [15:0]   io_coef_out_payload_0_38_46_imag,
  output     [15:0]   io_coef_out_payload_0_38_47_real,
  output     [15:0]   io_coef_out_payload_0_38_47_imag,
  output     [15:0]   io_coef_out_payload_0_38_48_real,
  output     [15:0]   io_coef_out_payload_0_38_48_imag,
  output     [15:0]   io_coef_out_payload_0_38_49_real,
  output     [15:0]   io_coef_out_payload_0_38_49_imag,
  output     [15:0]   io_coef_out_payload_0_39_0_real,
  output     [15:0]   io_coef_out_payload_0_39_0_imag,
  output     [15:0]   io_coef_out_payload_0_39_1_real,
  output     [15:0]   io_coef_out_payload_0_39_1_imag,
  output     [15:0]   io_coef_out_payload_0_39_2_real,
  output     [15:0]   io_coef_out_payload_0_39_2_imag,
  output     [15:0]   io_coef_out_payload_0_39_3_real,
  output     [15:0]   io_coef_out_payload_0_39_3_imag,
  output     [15:0]   io_coef_out_payload_0_39_4_real,
  output     [15:0]   io_coef_out_payload_0_39_4_imag,
  output     [15:0]   io_coef_out_payload_0_39_5_real,
  output     [15:0]   io_coef_out_payload_0_39_5_imag,
  output     [15:0]   io_coef_out_payload_0_39_6_real,
  output     [15:0]   io_coef_out_payload_0_39_6_imag,
  output     [15:0]   io_coef_out_payload_0_39_7_real,
  output     [15:0]   io_coef_out_payload_0_39_7_imag,
  output     [15:0]   io_coef_out_payload_0_39_8_real,
  output     [15:0]   io_coef_out_payload_0_39_8_imag,
  output     [15:0]   io_coef_out_payload_0_39_9_real,
  output     [15:0]   io_coef_out_payload_0_39_9_imag,
  output     [15:0]   io_coef_out_payload_0_39_10_real,
  output     [15:0]   io_coef_out_payload_0_39_10_imag,
  output     [15:0]   io_coef_out_payload_0_39_11_real,
  output     [15:0]   io_coef_out_payload_0_39_11_imag,
  output     [15:0]   io_coef_out_payload_0_39_12_real,
  output     [15:0]   io_coef_out_payload_0_39_12_imag,
  output     [15:0]   io_coef_out_payload_0_39_13_real,
  output     [15:0]   io_coef_out_payload_0_39_13_imag,
  output     [15:0]   io_coef_out_payload_0_39_14_real,
  output     [15:0]   io_coef_out_payload_0_39_14_imag,
  output     [15:0]   io_coef_out_payload_0_39_15_real,
  output     [15:0]   io_coef_out_payload_0_39_15_imag,
  output     [15:0]   io_coef_out_payload_0_39_16_real,
  output     [15:0]   io_coef_out_payload_0_39_16_imag,
  output     [15:0]   io_coef_out_payload_0_39_17_real,
  output     [15:0]   io_coef_out_payload_0_39_17_imag,
  output     [15:0]   io_coef_out_payload_0_39_18_real,
  output     [15:0]   io_coef_out_payload_0_39_18_imag,
  output     [15:0]   io_coef_out_payload_0_39_19_real,
  output     [15:0]   io_coef_out_payload_0_39_19_imag,
  output     [15:0]   io_coef_out_payload_0_39_20_real,
  output     [15:0]   io_coef_out_payload_0_39_20_imag,
  output     [15:0]   io_coef_out_payload_0_39_21_real,
  output     [15:0]   io_coef_out_payload_0_39_21_imag,
  output     [15:0]   io_coef_out_payload_0_39_22_real,
  output     [15:0]   io_coef_out_payload_0_39_22_imag,
  output     [15:0]   io_coef_out_payload_0_39_23_real,
  output     [15:0]   io_coef_out_payload_0_39_23_imag,
  output     [15:0]   io_coef_out_payload_0_39_24_real,
  output     [15:0]   io_coef_out_payload_0_39_24_imag,
  output     [15:0]   io_coef_out_payload_0_39_25_real,
  output     [15:0]   io_coef_out_payload_0_39_25_imag,
  output     [15:0]   io_coef_out_payload_0_39_26_real,
  output     [15:0]   io_coef_out_payload_0_39_26_imag,
  output     [15:0]   io_coef_out_payload_0_39_27_real,
  output     [15:0]   io_coef_out_payload_0_39_27_imag,
  output     [15:0]   io_coef_out_payload_0_39_28_real,
  output     [15:0]   io_coef_out_payload_0_39_28_imag,
  output     [15:0]   io_coef_out_payload_0_39_29_real,
  output     [15:0]   io_coef_out_payload_0_39_29_imag,
  output     [15:0]   io_coef_out_payload_0_39_30_real,
  output     [15:0]   io_coef_out_payload_0_39_30_imag,
  output     [15:0]   io_coef_out_payload_0_39_31_real,
  output     [15:0]   io_coef_out_payload_0_39_31_imag,
  output     [15:0]   io_coef_out_payload_0_39_32_real,
  output     [15:0]   io_coef_out_payload_0_39_32_imag,
  output     [15:0]   io_coef_out_payload_0_39_33_real,
  output     [15:0]   io_coef_out_payload_0_39_33_imag,
  output     [15:0]   io_coef_out_payload_0_39_34_real,
  output     [15:0]   io_coef_out_payload_0_39_34_imag,
  output     [15:0]   io_coef_out_payload_0_39_35_real,
  output     [15:0]   io_coef_out_payload_0_39_35_imag,
  output     [15:0]   io_coef_out_payload_0_39_36_real,
  output     [15:0]   io_coef_out_payload_0_39_36_imag,
  output     [15:0]   io_coef_out_payload_0_39_37_real,
  output     [15:0]   io_coef_out_payload_0_39_37_imag,
  output     [15:0]   io_coef_out_payload_0_39_38_real,
  output     [15:0]   io_coef_out_payload_0_39_38_imag,
  output     [15:0]   io_coef_out_payload_0_39_39_real,
  output     [15:0]   io_coef_out_payload_0_39_39_imag,
  output     [15:0]   io_coef_out_payload_0_39_40_real,
  output     [15:0]   io_coef_out_payload_0_39_40_imag,
  output     [15:0]   io_coef_out_payload_0_39_41_real,
  output     [15:0]   io_coef_out_payload_0_39_41_imag,
  output     [15:0]   io_coef_out_payload_0_39_42_real,
  output     [15:0]   io_coef_out_payload_0_39_42_imag,
  output     [15:0]   io_coef_out_payload_0_39_43_real,
  output     [15:0]   io_coef_out_payload_0_39_43_imag,
  output     [15:0]   io_coef_out_payload_0_39_44_real,
  output     [15:0]   io_coef_out_payload_0_39_44_imag,
  output     [15:0]   io_coef_out_payload_0_39_45_real,
  output     [15:0]   io_coef_out_payload_0_39_45_imag,
  output     [15:0]   io_coef_out_payload_0_39_46_real,
  output     [15:0]   io_coef_out_payload_0_39_46_imag,
  output     [15:0]   io_coef_out_payload_0_39_47_real,
  output     [15:0]   io_coef_out_payload_0_39_47_imag,
  output     [15:0]   io_coef_out_payload_0_39_48_real,
  output     [15:0]   io_coef_out_payload_0_39_48_imag,
  output     [15:0]   io_coef_out_payload_0_39_49_real,
  output     [15:0]   io_coef_out_payload_0_39_49_imag,
  output     [15:0]   io_coef_out_payload_0_40_0_real,
  output     [15:0]   io_coef_out_payload_0_40_0_imag,
  output     [15:0]   io_coef_out_payload_0_40_1_real,
  output     [15:0]   io_coef_out_payload_0_40_1_imag,
  output     [15:0]   io_coef_out_payload_0_40_2_real,
  output     [15:0]   io_coef_out_payload_0_40_2_imag,
  output     [15:0]   io_coef_out_payload_0_40_3_real,
  output     [15:0]   io_coef_out_payload_0_40_3_imag,
  output     [15:0]   io_coef_out_payload_0_40_4_real,
  output     [15:0]   io_coef_out_payload_0_40_4_imag,
  output     [15:0]   io_coef_out_payload_0_40_5_real,
  output     [15:0]   io_coef_out_payload_0_40_5_imag,
  output     [15:0]   io_coef_out_payload_0_40_6_real,
  output     [15:0]   io_coef_out_payload_0_40_6_imag,
  output     [15:0]   io_coef_out_payload_0_40_7_real,
  output     [15:0]   io_coef_out_payload_0_40_7_imag,
  output     [15:0]   io_coef_out_payload_0_40_8_real,
  output     [15:0]   io_coef_out_payload_0_40_8_imag,
  output     [15:0]   io_coef_out_payload_0_40_9_real,
  output     [15:0]   io_coef_out_payload_0_40_9_imag,
  output     [15:0]   io_coef_out_payload_0_40_10_real,
  output     [15:0]   io_coef_out_payload_0_40_10_imag,
  output     [15:0]   io_coef_out_payload_0_40_11_real,
  output     [15:0]   io_coef_out_payload_0_40_11_imag,
  output     [15:0]   io_coef_out_payload_0_40_12_real,
  output     [15:0]   io_coef_out_payload_0_40_12_imag,
  output     [15:0]   io_coef_out_payload_0_40_13_real,
  output     [15:0]   io_coef_out_payload_0_40_13_imag,
  output     [15:0]   io_coef_out_payload_0_40_14_real,
  output     [15:0]   io_coef_out_payload_0_40_14_imag,
  output     [15:0]   io_coef_out_payload_0_40_15_real,
  output     [15:0]   io_coef_out_payload_0_40_15_imag,
  output     [15:0]   io_coef_out_payload_0_40_16_real,
  output     [15:0]   io_coef_out_payload_0_40_16_imag,
  output     [15:0]   io_coef_out_payload_0_40_17_real,
  output     [15:0]   io_coef_out_payload_0_40_17_imag,
  output     [15:0]   io_coef_out_payload_0_40_18_real,
  output     [15:0]   io_coef_out_payload_0_40_18_imag,
  output     [15:0]   io_coef_out_payload_0_40_19_real,
  output     [15:0]   io_coef_out_payload_0_40_19_imag,
  output     [15:0]   io_coef_out_payload_0_40_20_real,
  output     [15:0]   io_coef_out_payload_0_40_20_imag,
  output     [15:0]   io_coef_out_payload_0_40_21_real,
  output     [15:0]   io_coef_out_payload_0_40_21_imag,
  output     [15:0]   io_coef_out_payload_0_40_22_real,
  output     [15:0]   io_coef_out_payload_0_40_22_imag,
  output     [15:0]   io_coef_out_payload_0_40_23_real,
  output     [15:0]   io_coef_out_payload_0_40_23_imag,
  output     [15:0]   io_coef_out_payload_0_40_24_real,
  output     [15:0]   io_coef_out_payload_0_40_24_imag,
  output     [15:0]   io_coef_out_payload_0_40_25_real,
  output     [15:0]   io_coef_out_payload_0_40_25_imag,
  output     [15:0]   io_coef_out_payload_0_40_26_real,
  output     [15:0]   io_coef_out_payload_0_40_26_imag,
  output     [15:0]   io_coef_out_payload_0_40_27_real,
  output     [15:0]   io_coef_out_payload_0_40_27_imag,
  output     [15:0]   io_coef_out_payload_0_40_28_real,
  output     [15:0]   io_coef_out_payload_0_40_28_imag,
  output     [15:0]   io_coef_out_payload_0_40_29_real,
  output     [15:0]   io_coef_out_payload_0_40_29_imag,
  output     [15:0]   io_coef_out_payload_0_40_30_real,
  output     [15:0]   io_coef_out_payload_0_40_30_imag,
  output     [15:0]   io_coef_out_payload_0_40_31_real,
  output     [15:0]   io_coef_out_payload_0_40_31_imag,
  output     [15:0]   io_coef_out_payload_0_40_32_real,
  output     [15:0]   io_coef_out_payload_0_40_32_imag,
  output     [15:0]   io_coef_out_payload_0_40_33_real,
  output     [15:0]   io_coef_out_payload_0_40_33_imag,
  output     [15:0]   io_coef_out_payload_0_40_34_real,
  output     [15:0]   io_coef_out_payload_0_40_34_imag,
  output     [15:0]   io_coef_out_payload_0_40_35_real,
  output     [15:0]   io_coef_out_payload_0_40_35_imag,
  output     [15:0]   io_coef_out_payload_0_40_36_real,
  output     [15:0]   io_coef_out_payload_0_40_36_imag,
  output     [15:0]   io_coef_out_payload_0_40_37_real,
  output     [15:0]   io_coef_out_payload_0_40_37_imag,
  output     [15:0]   io_coef_out_payload_0_40_38_real,
  output     [15:0]   io_coef_out_payload_0_40_38_imag,
  output     [15:0]   io_coef_out_payload_0_40_39_real,
  output     [15:0]   io_coef_out_payload_0_40_39_imag,
  output     [15:0]   io_coef_out_payload_0_40_40_real,
  output     [15:0]   io_coef_out_payload_0_40_40_imag,
  output     [15:0]   io_coef_out_payload_0_40_41_real,
  output     [15:0]   io_coef_out_payload_0_40_41_imag,
  output     [15:0]   io_coef_out_payload_0_40_42_real,
  output     [15:0]   io_coef_out_payload_0_40_42_imag,
  output     [15:0]   io_coef_out_payload_0_40_43_real,
  output     [15:0]   io_coef_out_payload_0_40_43_imag,
  output     [15:0]   io_coef_out_payload_0_40_44_real,
  output     [15:0]   io_coef_out_payload_0_40_44_imag,
  output     [15:0]   io_coef_out_payload_0_40_45_real,
  output     [15:0]   io_coef_out_payload_0_40_45_imag,
  output     [15:0]   io_coef_out_payload_0_40_46_real,
  output     [15:0]   io_coef_out_payload_0_40_46_imag,
  output     [15:0]   io_coef_out_payload_0_40_47_real,
  output     [15:0]   io_coef_out_payload_0_40_47_imag,
  output     [15:0]   io_coef_out_payload_0_40_48_real,
  output     [15:0]   io_coef_out_payload_0_40_48_imag,
  output     [15:0]   io_coef_out_payload_0_40_49_real,
  output     [15:0]   io_coef_out_payload_0_40_49_imag,
  output     [15:0]   io_coef_out_payload_0_41_0_real,
  output     [15:0]   io_coef_out_payload_0_41_0_imag,
  output     [15:0]   io_coef_out_payload_0_41_1_real,
  output     [15:0]   io_coef_out_payload_0_41_1_imag,
  output     [15:0]   io_coef_out_payload_0_41_2_real,
  output     [15:0]   io_coef_out_payload_0_41_2_imag,
  output     [15:0]   io_coef_out_payload_0_41_3_real,
  output     [15:0]   io_coef_out_payload_0_41_3_imag,
  output     [15:0]   io_coef_out_payload_0_41_4_real,
  output     [15:0]   io_coef_out_payload_0_41_4_imag,
  output     [15:0]   io_coef_out_payload_0_41_5_real,
  output     [15:0]   io_coef_out_payload_0_41_5_imag,
  output     [15:0]   io_coef_out_payload_0_41_6_real,
  output     [15:0]   io_coef_out_payload_0_41_6_imag,
  output     [15:0]   io_coef_out_payload_0_41_7_real,
  output     [15:0]   io_coef_out_payload_0_41_7_imag,
  output     [15:0]   io_coef_out_payload_0_41_8_real,
  output     [15:0]   io_coef_out_payload_0_41_8_imag,
  output     [15:0]   io_coef_out_payload_0_41_9_real,
  output     [15:0]   io_coef_out_payload_0_41_9_imag,
  output     [15:0]   io_coef_out_payload_0_41_10_real,
  output     [15:0]   io_coef_out_payload_0_41_10_imag,
  output     [15:0]   io_coef_out_payload_0_41_11_real,
  output     [15:0]   io_coef_out_payload_0_41_11_imag,
  output     [15:0]   io_coef_out_payload_0_41_12_real,
  output     [15:0]   io_coef_out_payload_0_41_12_imag,
  output     [15:0]   io_coef_out_payload_0_41_13_real,
  output     [15:0]   io_coef_out_payload_0_41_13_imag,
  output     [15:0]   io_coef_out_payload_0_41_14_real,
  output     [15:0]   io_coef_out_payload_0_41_14_imag,
  output     [15:0]   io_coef_out_payload_0_41_15_real,
  output     [15:0]   io_coef_out_payload_0_41_15_imag,
  output     [15:0]   io_coef_out_payload_0_41_16_real,
  output     [15:0]   io_coef_out_payload_0_41_16_imag,
  output     [15:0]   io_coef_out_payload_0_41_17_real,
  output     [15:0]   io_coef_out_payload_0_41_17_imag,
  output     [15:0]   io_coef_out_payload_0_41_18_real,
  output     [15:0]   io_coef_out_payload_0_41_18_imag,
  output     [15:0]   io_coef_out_payload_0_41_19_real,
  output     [15:0]   io_coef_out_payload_0_41_19_imag,
  output     [15:0]   io_coef_out_payload_0_41_20_real,
  output     [15:0]   io_coef_out_payload_0_41_20_imag,
  output     [15:0]   io_coef_out_payload_0_41_21_real,
  output     [15:0]   io_coef_out_payload_0_41_21_imag,
  output     [15:0]   io_coef_out_payload_0_41_22_real,
  output     [15:0]   io_coef_out_payload_0_41_22_imag,
  output     [15:0]   io_coef_out_payload_0_41_23_real,
  output     [15:0]   io_coef_out_payload_0_41_23_imag,
  output     [15:0]   io_coef_out_payload_0_41_24_real,
  output     [15:0]   io_coef_out_payload_0_41_24_imag,
  output     [15:0]   io_coef_out_payload_0_41_25_real,
  output     [15:0]   io_coef_out_payload_0_41_25_imag,
  output     [15:0]   io_coef_out_payload_0_41_26_real,
  output     [15:0]   io_coef_out_payload_0_41_26_imag,
  output     [15:0]   io_coef_out_payload_0_41_27_real,
  output     [15:0]   io_coef_out_payload_0_41_27_imag,
  output     [15:0]   io_coef_out_payload_0_41_28_real,
  output     [15:0]   io_coef_out_payload_0_41_28_imag,
  output     [15:0]   io_coef_out_payload_0_41_29_real,
  output     [15:0]   io_coef_out_payload_0_41_29_imag,
  output     [15:0]   io_coef_out_payload_0_41_30_real,
  output     [15:0]   io_coef_out_payload_0_41_30_imag,
  output     [15:0]   io_coef_out_payload_0_41_31_real,
  output     [15:0]   io_coef_out_payload_0_41_31_imag,
  output     [15:0]   io_coef_out_payload_0_41_32_real,
  output     [15:0]   io_coef_out_payload_0_41_32_imag,
  output     [15:0]   io_coef_out_payload_0_41_33_real,
  output     [15:0]   io_coef_out_payload_0_41_33_imag,
  output     [15:0]   io_coef_out_payload_0_41_34_real,
  output     [15:0]   io_coef_out_payload_0_41_34_imag,
  output     [15:0]   io_coef_out_payload_0_41_35_real,
  output     [15:0]   io_coef_out_payload_0_41_35_imag,
  output     [15:0]   io_coef_out_payload_0_41_36_real,
  output     [15:0]   io_coef_out_payload_0_41_36_imag,
  output     [15:0]   io_coef_out_payload_0_41_37_real,
  output     [15:0]   io_coef_out_payload_0_41_37_imag,
  output     [15:0]   io_coef_out_payload_0_41_38_real,
  output     [15:0]   io_coef_out_payload_0_41_38_imag,
  output     [15:0]   io_coef_out_payload_0_41_39_real,
  output     [15:0]   io_coef_out_payload_0_41_39_imag,
  output     [15:0]   io_coef_out_payload_0_41_40_real,
  output     [15:0]   io_coef_out_payload_0_41_40_imag,
  output     [15:0]   io_coef_out_payload_0_41_41_real,
  output     [15:0]   io_coef_out_payload_0_41_41_imag,
  output     [15:0]   io_coef_out_payload_0_41_42_real,
  output     [15:0]   io_coef_out_payload_0_41_42_imag,
  output     [15:0]   io_coef_out_payload_0_41_43_real,
  output     [15:0]   io_coef_out_payload_0_41_43_imag,
  output     [15:0]   io_coef_out_payload_0_41_44_real,
  output     [15:0]   io_coef_out_payload_0_41_44_imag,
  output     [15:0]   io_coef_out_payload_0_41_45_real,
  output     [15:0]   io_coef_out_payload_0_41_45_imag,
  output     [15:0]   io_coef_out_payload_0_41_46_real,
  output     [15:0]   io_coef_out_payload_0_41_46_imag,
  output     [15:0]   io_coef_out_payload_0_41_47_real,
  output     [15:0]   io_coef_out_payload_0_41_47_imag,
  output     [15:0]   io_coef_out_payload_0_41_48_real,
  output     [15:0]   io_coef_out_payload_0_41_48_imag,
  output     [15:0]   io_coef_out_payload_0_41_49_real,
  output     [15:0]   io_coef_out_payload_0_41_49_imag,
  output     [15:0]   io_coef_out_payload_0_42_0_real,
  output     [15:0]   io_coef_out_payload_0_42_0_imag,
  output     [15:0]   io_coef_out_payload_0_42_1_real,
  output     [15:0]   io_coef_out_payload_0_42_1_imag,
  output     [15:0]   io_coef_out_payload_0_42_2_real,
  output     [15:0]   io_coef_out_payload_0_42_2_imag,
  output     [15:0]   io_coef_out_payload_0_42_3_real,
  output     [15:0]   io_coef_out_payload_0_42_3_imag,
  output     [15:0]   io_coef_out_payload_0_42_4_real,
  output     [15:0]   io_coef_out_payload_0_42_4_imag,
  output     [15:0]   io_coef_out_payload_0_42_5_real,
  output     [15:0]   io_coef_out_payload_0_42_5_imag,
  output     [15:0]   io_coef_out_payload_0_42_6_real,
  output     [15:0]   io_coef_out_payload_0_42_6_imag,
  output     [15:0]   io_coef_out_payload_0_42_7_real,
  output     [15:0]   io_coef_out_payload_0_42_7_imag,
  output     [15:0]   io_coef_out_payload_0_42_8_real,
  output     [15:0]   io_coef_out_payload_0_42_8_imag,
  output     [15:0]   io_coef_out_payload_0_42_9_real,
  output     [15:0]   io_coef_out_payload_0_42_9_imag,
  output     [15:0]   io_coef_out_payload_0_42_10_real,
  output     [15:0]   io_coef_out_payload_0_42_10_imag,
  output     [15:0]   io_coef_out_payload_0_42_11_real,
  output     [15:0]   io_coef_out_payload_0_42_11_imag,
  output     [15:0]   io_coef_out_payload_0_42_12_real,
  output     [15:0]   io_coef_out_payload_0_42_12_imag,
  output     [15:0]   io_coef_out_payload_0_42_13_real,
  output     [15:0]   io_coef_out_payload_0_42_13_imag,
  output     [15:0]   io_coef_out_payload_0_42_14_real,
  output     [15:0]   io_coef_out_payload_0_42_14_imag,
  output     [15:0]   io_coef_out_payload_0_42_15_real,
  output     [15:0]   io_coef_out_payload_0_42_15_imag,
  output     [15:0]   io_coef_out_payload_0_42_16_real,
  output     [15:0]   io_coef_out_payload_0_42_16_imag,
  output     [15:0]   io_coef_out_payload_0_42_17_real,
  output     [15:0]   io_coef_out_payload_0_42_17_imag,
  output     [15:0]   io_coef_out_payload_0_42_18_real,
  output     [15:0]   io_coef_out_payload_0_42_18_imag,
  output     [15:0]   io_coef_out_payload_0_42_19_real,
  output     [15:0]   io_coef_out_payload_0_42_19_imag,
  output     [15:0]   io_coef_out_payload_0_42_20_real,
  output     [15:0]   io_coef_out_payload_0_42_20_imag,
  output     [15:0]   io_coef_out_payload_0_42_21_real,
  output     [15:0]   io_coef_out_payload_0_42_21_imag,
  output     [15:0]   io_coef_out_payload_0_42_22_real,
  output     [15:0]   io_coef_out_payload_0_42_22_imag,
  output     [15:0]   io_coef_out_payload_0_42_23_real,
  output     [15:0]   io_coef_out_payload_0_42_23_imag,
  output     [15:0]   io_coef_out_payload_0_42_24_real,
  output     [15:0]   io_coef_out_payload_0_42_24_imag,
  output     [15:0]   io_coef_out_payload_0_42_25_real,
  output     [15:0]   io_coef_out_payload_0_42_25_imag,
  output     [15:0]   io_coef_out_payload_0_42_26_real,
  output     [15:0]   io_coef_out_payload_0_42_26_imag,
  output     [15:0]   io_coef_out_payload_0_42_27_real,
  output     [15:0]   io_coef_out_payload_0_42_27_imag,
  output     [15:0]   io_coef_out_payload_0_42_28_real,
  output     [15:0]   io_coef_out_payload_0_42_28_imag,
  output     [15:0]   io_coef_out_payload_0_42_29_real,
  output     [15:0]   io_coef_out_payload_0_42_29_imag,
  output     [15:0]   io_coef_out_payload_0_42_30_real,
  output     [15:0]   io_coef_out_payload_0_42_30_imag,
  output     [15:0]   io_coef_out_payload_0_42_31_real,
  output     [15:0]   io_coef_out_payload_0_42_31_imag,
  output     [15:0]   io_coef_out_payload_0_42_32_real,
  output     [15:0]   io_coef_out_payload_0_42_32_imag,
  output     [15:0]   io_coef_out_payload_0_42_33_real,
  output     [15:0]   io_coef_out_payload_0_42_33_imag,
  output     [15:0]   io_coef_out_payload_0_42_34_real,
  output     [15:0]   io_coef_out_payload_0_42_34_imag,
  output     [15:0]   io_coef_out_payload_0_42_35_real,
  output     [15:0]   io_coef_out_payload_0_42_35_imag,
  output     [15:0]   io_coef_out_payload_0_42_36_real,
  output     [15:0]   io_coef_out_payload_0_42_36_imag,
  output     [15:0]   io_coef_out_payload_0_42_37_real,
  output     [15:0]   io_coef_out_payload_0_42_37_imag,
  output     [15:0]   io_coef_out_payload_0_42_38_real,
  output     [15:0]   io_coef_out_payload_0_42_38_imag,
  output     [15:0]   io_coef_out_payload_0_42_39_real,
  output     [15:0]   io_coef_out_payload_0_42_39_imag,
  output     [15:0]   io_coef_out_payload_0_42_40_real,
  output     [15:0]   io_coef_out_payload_0_42_40_imag,
  output     [15:0]   io_coef_out_payload_0_42_41_real,
  output     [15:0]   io_coef_out_payload_0_42_41_imag,
  output     [15:0]   io_coef_out_payload_0_42_42_real,
  output     [15:0]   io_coef_out_payload_0_42_42_imag,
  output     [15:0]   io_coef_out_payload_0_42_43_real,
  output     [15:0]   io_coef_out_payload_0_42_43_imag,
  output     [15:0]   io_coef_out_payload_0_42_44_real,
  output     [15:0]   io_coef_out_payload_0_42_44_imag,
  output     [15:0]   io_coef_out_payload_0_42_45_real,
  output     [15:0]   io_coef_out_payload_0_42_45_imag,
  output     [15:0]   io_coef_out_payload_0_42_46_real,
  output     [15:0]   io_coef_out_payload_0_42_46_imag,
  output     [15:0]   io_coef_out_payload_0_42_47_real,
  output     [15:0]   io_coef_out_payload_0_42_47_imag,
  output     [15:0]   io_coef_out_payload_0_42_48_real,
  output     [15:0]   io_coef_out_payload_0_42_48_imag,
  output     [15:0]   io_coef_out_payload_0_42_49_real,
  output     [15:0]   io_coef_out_payload_0_42_49_imag,
  output     [15:0]   io_coef_out_payload_0_43_0_real,
  output     [15:0]   io_coef_out_payload_0_43_0_imag,
  output     [15:0]   io_coef_out_payload_0_43_1_real,
  output     [15:0]   io_coef_out_payload_0_43_1_imag,
  output     [15:0]   io_coef_out_payload_0_43_2_real,
  output     [15:0]   io_coef_out_payload_0_43_2_imag,
  output     [15:0]   io_coef_out_payload_0_43_3_real,
  output     [15:0]   io_coef_out_payload_0_43_3_imag,
  output     [15:0]   io_coef_out_payload_0_43_4_real,
  output     [15:0]   io_coef_out_payload_0_43_4_imag,
  output     [15:0]   io_coef_out_payload_0_43_5_real,
  output     [15:0]   io_coef_out_payload_0_43_5_imag,
  output     [15:0]   io_coef_out_payload_0_43_6_real,
  output     [15:0]   io_coef_out_payload_0_43_6_imag,
  output     [15:0]   io_coef_out_payload_0_43_7_real,
  output     [15:0]   io_coef_out_payload_0_43_7_imag,
  output     [15:0]   io_coef_out_payload_0_43_8_real,
  output     [15:0]   io_coef_out_payload_0_43_8_imag,
  output     [15:0]   io_coef_out_payload_0_43_9_real,
  output     [15:0]   io_coef_out_payload_0_43_9_imag,
  output     [15:0]   io_coef_out_payload_0_43_10_real,
  output     [15:0]   io_coef_out_payload_0_43_10_imag,
  output     [15:0]   io_coef_out_payload_0_43_11_real,
  output     [15:0]   io_coef_out_payload_0_43_11_imag,
  output     [15:0]   io_coef_out_payload_0_43_12_real,
  output     [15:0]   io_coef_out_payload_0_43_12_imag,
  output     [15:0]   io_coef_out_payload_0_43_13_real,
  output     [15:0]   io_coef_out_payload_0_43_13_imag,
  output     [15:0]   io_coef_out_payload_0_43_14_real,
  output     [15:0]   io_coef_out_payload_0_43_14_imag,
  output     [15:0]   io_coef_out_payload_0_43_15_real,
  output     [15:0]   io_coef_out_payload_0_43_15_imag,
  output     [15:0]   io_coef_out_payload_0_43_16_real,
  output     [15:0]   io_coef_out_payload_0_43_16_imag,
  output     [15:0]   io_coef_out_payload_0_43_17_real,
  output     [15:0]   io_coef_out_payload_0_43_17_imag,
  output     [15:0]   io_coef_out_payload_0_43_18_real,
  output     [15:0]   io_coef_out_payload_0_43_18_imag,
  output     [15:0]   io_coef_out_payload_0_43_19_real,
  output     [15:0]   io_coef_out_payload_0_43_19_imag,
  output     [15:0]   io_coef_out_payload_0_43_20_real,
  output     [15:0]   io_coef_out_payload_0_43_20_imag,
  output     [15:0]   io_coef_out_payload_0_43_21_real,
  output     [15:0]   io_coef_out_payload_0_43_21_imag,
  output     [15:0]   io_coef_out_payload_0_43_22_real,
  output     [15:0]   io_coef_out_payload_0_43_22_imag,
  output     [15:0]   io_coef_out_payload_0_43_23_real,
  output     [15:0]   io_coef_out_payload_0_43_23_imag,
  output     [15:0]   io_coef_out_payload_0_43_24_real,
  output     [15:0]   io_coef_out_payload_0_43_24_imag,
  output     [15:0]   io_coef_out_payload_0_43_25_real,
  output     [15:0]   io_coef_out_payload_0_43_25_imag,
  output     [15:0]   io_coef_out_payload_0_43_26_real,
  output     [15:0]   io_coef_out_payload_0_43_26_imag,
  output     [15:0]   io_coef_out_payload_0_43_27_real,
  output     [15:0]   io_coef_out_payload_0_43_27_imag,
  output     [15:0]   io_coef_out_payload_0_43_28_real,
  output     [15:0]   io_coef_out_payload_0_43_28_imag,
  output     [15:0]   io_coef_out_payload_0_43_29_real,
  output     [15:0]   io_coef_out_payload_0_43_29_imag,
  output     [15:0]   io_coef_out_payload_0_43_30_real,
  output     [15:0]   io_coef_out_payload_0_43_30_imag,
  output     [15:0]   io_coef_out_payload_0_43_31_real,
  output     [15:0]   io_coef_out_payload_0_43_31_imag,
  output     [15:0]   io_coef_out_payload_0_43_32_real,
  output     [15:0]   io_coef_out_payload_0_43_32_imag,
  output     [15:0]   io_coef_out_payload_0_43_33_real,
  output     [15:0]   io_coef_out_payload_0_43_33_imag,
  output     [15:0]   io_coef_out_payload_0_43_34_real,
  output     [15:0]   io_coef_out_payload_0_43_34_imag,
  output     [15:0]   io_coef_out_payload_0_43_35_real,
  output     [15:0]   io_coef_out_payload_0_43_35_imag,
  output     [15:0]   io_coef_out_payload_0_43_36_real,
  output     [15:0]   io_coef_out_payload_0_43_36_imag,
  output     [15:0]   io_coef_out_payload_0_43_37_real,
  output     [15:0]   io_coef_out_payload_0_43_37_imag,
  output     [15:0]   io_coef_out_payload_0_43_38_real,
  output     [15:0]   io_coef_out_payload_0_43_38_imag,
  output     [15:0]   io_coef_out_payload_0_43_39_real,
  output     [15:0]   io_coef_out_payload_0_43_39_imag,
  output     [15:0]   io_coef_out_payload_0_43_40_real,
  output     [15:0]   io_coef_out_payload_0_43_40_imag,
  output     [15:0]   io_coef_out_payload_0_43_41_real,
  output     [15:0]   io_coef_out_payload_0_43_41_imag,
  output     [15:0]   io_coef_out_payload_0_43_42_real,
  output     [15:0]   io_coef_out_payload_0_43_42_imag,
  output     [15:0]   io_coef_out_payload_0_43_43_real,
  output     [15:0]   io_coef_out_payload_0_43_43_imag,
  output     [15:0]   io_coef_out_payload_0_43_44_real,
  output     [15:0]   io_coef_out_payload_0_43_44_imag,
  output     [15:0]   io_coef_out_payload_0_43_45_real,
  output     [15:0]   io_coef_out_payload_0_43_45_imag,
  output     [15:0]   io_coef_out_payload_0_43_46_real,
  output     [15:0]   io_coef_out_payload_0_43_46_imag,
  output     [15:0]   io_coef_out_payload_0_43_47_real,
  output     [15:0]   io_coef_out_payload_0_43_47_imag,
  output     [15:0]   io_coef_out_payload_0_43_48_real,
  output     [15:0]   io_coef_out_payload_0_43_48_imag,
  output     [15:0]   io_coef_out_payload_0_43_49_real,
  output     [15:0]   io_coef_out_payload_0_43_49_imag,
  output     [15:0]   io_coef_out_payload_0_44_0_real,
  output     [15:0]   io_coef_out_payload_0_44_0_imag,
  output     [15:0]   io_coef_out_payload_0_44_1_real,
  output     [15:0]   io_coef_out_payload_0_44_1_imag,
  output     [15:0]   io_coef_out_payload_0_44_2_real,
  output     [15:0]   io_coef_out_payload_0_44_2_imag,
  output     [15:0]   io_coef_out_payload_0_44_3_real,
  output     [15:0]   io_coef_out_payload_0_44_3_imag,
  output     [15:0]   io_coef_out_payload_0_44_4_real,
  output     [15:0]   io_coef_out_payload_0_44_4_imag,
  output     [15:0]   io_coef_out_payload_0_44_5_real,
  output     [15:0]   io_coef_out_payload_0_44_5_imag,
  output     [15:0]   io_coef_out_payload_0_44_6_real,
  output     [15:0]   io_coef_out_payload_0_44_6_imag,
  output     [15:0]   io_coef_out_payload_0_44_7_real,
  output     [15:0]   io_coef_out_payload_0_44_7_imag,
  output     [15:0]   io_coef_out_payload_0_44_8_real,
  output     [15:0]   io_coef_out_payload_0_44_8_imag,
  output     [15:0]   io_coef_out_payload_0_44_9_real,
  output     [15:0]   io_coef_out_payload_0_44_9_imag,
  output     [15:0]   io_coef_out_payload_0_44_10_real,
  output     [15:0]   io_coef_out_payload_0_44_10_imag,
  output     [15:0]   io_coef_out_payload_0_44_11_real,
  output     [15:0]   io_coef_out_payload_0_44_11_imag,
  output     [15:0]   io_coef_out_payload_0_44_12_real,
  output     [15:0]   io_coef_out_payload_0_44_12_imag,
  output     [15:0]   io_coef_out_payload_0_44_13_real,
  output     [15:0]   io_coef_out_payload_0_44_13_imag,
  output     [15:0]   io_coef_out_payload_0_44_14_real,
  output     [15:0]   io_coef_out_payload_0_44_14_imag,
  output     [15:0]   io_coef_out_payload_0_44_15_real,
  output     [15:0]   io_coef_out_payload_0_44_15_imag,
  output     [15:0]   io_coef_out_payload_0_44_16_real,
  output     [15:0]   io_coef_out_payload_0_44_16_imag,
  output     [15:0]   io_coef_out_payload_0_44_17_real,
  output     [15:0]   io_coef_out_payload_0_44_17_imag,
  output     [15:0]   io_coef_out_payload_0_44_18_real,
  output     [15:0]   io_coef_out_payload_0_44_18_imag,
  output     [15:0]   io_coef_out_payload_0_44_19_real,
  output     [15:0]   io_coef_out_payload_0_44_19_imag,
  output     [15:0]   io_coef_out_payload_0_44_20_real,
  output     [15:0]   io_coef_out_payload_0_44_20_imag,
  output     [15:0]   io_coef_out_payload_0_44_21_real,
  output     [15:0]   io_coef_out_payload_0_44_21_imag,
  output     [15:0]   io_coef_out_payload_0_44_22_real,
  output     [15:0]   io_coef_out_payload_0_44_22_imag,
  output     [15:0]   io_coef_out_payload_0_44_23_real,
  output     [15:0]   io_coef_out_payload_0_44_23_imag,
  output     [15:0]   io_coef_out_payload_0_44_24_real,
  output     [15:0]   io_coef_out_payload_0_44_24_imag,
  output     [15:0]   io_coef_out_payload_0_44_25_real,
  output     [15:0]   io_coef_out_payload_0_44_25_imag,
  output     [15:0]   io_coef_out_payload_0_44_26_real,
  output     [15:0]   io_coef_out_payload_0_44_26_imag,
  output     [15:0]   io_coef_out_payload_0_44_27_real,
  output     [15:0]   io_coef_out_payload_0_44_27_imag,
  output     [15:0]   io_coef_out_payload_0_44_28_real,
  output     [15:0]   io_coef_out_payload_0_44_28_imag,
  output     [15:0]   io_coef_out_payload_0_44_29_real,
  output     [15:0]   io_coef_out_payload_0_44_29_imag,
  output     [15:0]   io_coef_out_payload_0_44_30_real,
  output     [15:0]   io_coef_out_payload_0_44_30_imag,
  output     [15:0]   io_coef_out_payload_0_44_31_real,
  output     [15:0]   io_coef_out_payload_0_44_31_imag,
  output     [15:0]   io_coef_out_payload_0_44_32_real,
  output     [15:0]   io_coef_out_payload_0_44_32_imag,
  output     [15:0]   io_coef_out_payload_0_44_33_real,
  output     [15:0]   io_coef_out_payload_0_44_33_imag,
  output     [15:0]   io_coef_out_payload_0_44_34_real,
  output     [15:0]   io_coef_out_payload_0_44_34_imag,
  output     [15:0]   io_coef_out_payload_0_44_35_real,
  output     [15:0]   io_coef_out_payload_0_44_35_imag,
  output     [15:0]   io_coef_out_payload_0_44_36_real,
  output     [15:0]   io_coef_out_payload_0_44_36_imag,
  output     [15:0]   io_coef_out_payload_0_44_37_real,
  output     [15:0]   io_coef_out_payload_0_44_37_imag,
  output     [15:0]   io_coef_out_payload_0_44_38_real,
  output     [15:0]   io_coef_out_payload_0_44_38_imag,
  output     [15:0]   io_coef_out_payload_0_44_39_real,
  output     [15:0]   io_coef_out_payload_0_44_39_imag,
  output     [15:0]   io_coef_out_payload_0_44_40_real,
  output     [15:0]   io_coef_out_payload_0_44_40_imag,
  output     [15:0]   io_coef_out_payload_0_44_41_real,
  output     [15:0]   io_coef_out_payload_0_44_41_imag,
  output     [15:0]   io_coef_out_payload_0_44_42_real,
  output     [15:0]   io_coef_out_payload_0_44_42_imag,
  output     [15:0]   io_coef_out_payload_0_44_43_real,
  output     [15:0]   io_coef_out_payload_0_44_43_imag,
  output     [15:0]   io_coef_out_payload_0_44_44_real,
  output     [15:0]   io_coef_out_payload_0_44_44_imag,
  output     [15:0]   io_coef_out_payload_0_44_45_real,
  output     [15:0]   io_coef_out_payload_0_44_45_imag,
  output     [15:0]   io_coef_out_payload_0_44_46_real,
  output     [15:0]   io_coef_out_payload_0_44_46_imag,
  output     [15:0]   io_coef_out_payload_0_44_47_real,
  output     [15:0]   io_coef_out_payload_0_44_47_imag,
  output     [15:0]   io_coef_out_payload_0_44_48_real,
  output     [15:0]   io_coef_out_payload_0_44_48_imag,
  output     [15:0]   io_coef_out_payload_0_44_49_real,
  output     [15:0]   io_coef_out_payload_0_44_49_imag,
  output     [15:0]   io_coef_out_payload_0_45_0_real,
  output     [15:0]   io_coef_out_payload_0_45_0_imag,
  output     [15:0]   io_coef_out_payload_0_45_1_real,
  output     [15:0]   io_coef_out_payload_0_45_1_imag,
  output     [15:0]   io_coef_out_payload_0_45_2_real,
  output     [15:0]   io_coef_out_payload_0_45_2_imag,
  output     [15:0]   io_coef_out_payload_0_45_3_real,
  output     [15:0]   io_coef_out_payload_0_45_3_imag,
  output     [15:0]   io_coef_out_payload_0_45_4_real,
  output     [15:0]   io_coef_out_payload_0_45_4_imag,
  output     [15:0]   io_coef_out_payload_0_45_5_real,
  output     [15:0]   io_coef_out_payload_0_45_5_imag,
  output     [15:0]   io_coef_out_payload_0_45_6_real,
  output     [15:0]   io_coef_out_payload_0_45_6_imag,
  output     [15:0]   io_coef_out_payload_0_45_7_real,
  output     [15:0]   io_coef_out_payload_0_45_7_imag,
  output     [15:0]   io_coef_out_payload_0_45_8_real,
  output     [15:0]   io_coef_out_payload_0_45_8_imag,
  output     [15:0]   io_coef_out_payload_0_45_9_real,
  output     [15:0]   io_coef_out_payload_0_45_9_imag,
  output     [15:0]   io_coef_out_payload_0_45_10_real,
  output     [15:0]   io_coef_out_payload_0_45_10_imag,
  output     [15:0]   io_coef_out_payload_0_45_11_real,
  output     [15:0]   io_coef_out_payload_0_45_11_imag,
  output     [15:0]   io_coef_out_payload_0_45_12_real,
  output     [15:0]   io_coef_out_payload_0_45_12_imag,
  output     [15:0]   io_coef_out_payload_0_45_13_real,
  output     [15:0]   io_coef_out_payload_0_45_13_imag,
  output     [15:0]   io_coef_out_payload_0_45_14_real,
  output     [15:0]   io_coef_out_payload_0_45_14_imag,
  output     [15:0]   io_coef_out_payload_0_45_15_real,
  output     [15:0]   io_coef_out_payload_0_45_15_imag,
  output     [15:0]   io_coef_out_payload_0_45_16_real,
  output     [15:0]   io_coef_out_payload_0_45_16_imag,
  output     [15:0]   io_coef_out_payload_0_45_17_real,
  output     [15:0]   io_coef_out_payload_0_45_17_imag,
  output     [15:0]   io_coef_out_payload_0_45_18_real,
  output     [15:0]   io_coef_out_payload_0_45_18_imag,
  output     [15:0]   io_coef_out_payload_0_45_19_real,
  output     [15:0]   io_coef_out_payload_0_45_19_imag,
  output     [15:0]   io_coef_out_payload_0_45_20_real,
  output     [15:0]   io_coef_out_payload_0_45_20_imag,
  output     [15:0]   io_coef_out_payload_0_45_21_real,
  output     [15:0]   io_coef_out_payload_0_45_21_imag,
  output     [15:0]   io_coef_out_payload_0_45_22_real,
  output     [15:0]   io_coef_out_payload_0_45_22_imag,
  output     [15:0]   io_coef_out_payload_0_45_23_real,
  output     [15:0]   io_coef_out_payload_0_45_23_imag,
  output     [15:0]   io_coef_out_payload_0_45_24_real,
  output     [15:0]   io_coef_out_payload_0_45_24_imag,
  output     [15:0]   io_coef_out_payload_0_45_25_real,
  output     [15:0]   io_coef_out_payload_0_45_25_imag,
  output     [15:0]   io_coef_out_payload_0_45_26_real,
  output     [15:0]   io_coef_out_payload_0_45_26_imag,
  output     [15:0]   io_coef_out_payload_0_45_27_real,
  output     [15:0]   io_coef_out_payload_0_45_27_imag,
  output     [15:0]   io_coef_out_payload_0_45_28_real,
  output     [15:0]   io_coef_out_payload_0_45_28_imag,
  output     [15:0]   io_coef_out_payload_0_45_29_real,
  output     [15:0]   io_coef_out_payload_0_45_29_imag,
  output     [15:0]   io_coef_out_payload_0_45_30_real,
  output     [15:0]   io_coef_out_payload_0_45_30_imag,
  output     [15:0]   io_coef_out_payload_0_45_31_real,
  output     [15:0]   io_coef_out_payload_0_45_31_imag,
  output     [15:0]   io_coef_out_payload_0_45_32_real,
  output     [15:0]   io_coef_out_payload_0_45_32_imag,
  output     [15:0]   io_coef_out_payload_0_45_33_real,
  output     [15:0]   io_coef_out_payload_0_45_33_imag,
  output     [15:0]   io_coef_out_payload_0_45_34_real,
  output     [15:0]   io_coef_out_payload_0_45_34_imag,
  output     [15:0]   io_coef_out_payload_0_45_35_real,
  output     [15:0]   io_coef_out_payload_0_45_35_imag,
  output     [15:0]   io_coef_out_payload_0_45_36_real,
  output     [15:0]   io_coef_out_payload_0_45_36_imag,
  output     [15:0]   io_coef_out_payload_0_45_37_real,
  output     [15:0]   io_coef_out_payload_0_45_37_imag,
  output     [15:0]   io_coef_out_payload_0_45_38_real,
  output     [15:0]   io_coef_out_payload_0_45_38_imag,
  output     [15:0]   io_coef_out_payload_0_45_39_real,
  output     [15:0]   io_coef_out_payload_0_45_39_imag,
  output     [15:0]   io_coef_out_payload_0_45_40_real,
  output     [15:0]   io_coef_out_payload_0_45_40_imag,
  output     [15:0]   io_coef_out_payload_0_45_41_real,
  output     [15:0]   io_coef_out_payload_0_45_41_imag,
  output     [15:0]   io_coef_out_payload_0_45_42_real,
  output     [15:0]   io_coef_out_payload_0_45_42_imag,
  output     [15:0]   io_coef_out_payload_0_45_43_real,
  output     [15:0]   io_coef_out_payload_0_45_43_imag,
  output     [15:0]   io_coef_out_payload_0_45_44_real,
  output     [15:0]   io_coef_out_payload_0_45_44_imag,
  output     [15:0]   io_coef_out_payload_0_45_45_real,
  output     [15:0]   io_coef_out_payload_0_45_45_imag,
  output     [15:0]   io_coef_out_payload_0_45_46_real,
  output     [15:0]   io_coef_out_payload_0_45_46_imag,
  output     [15:0]   io_coef_out_payload_0_45_47_real,
  output     [15:0]   io_coef_out_payload_0_45_47_imag,
  output     [15:0]   io_coef_out_payload_0_45_48_real,
  output     [15:0]   io_coef_out_payload_0_45_48_imag,
  output     [15:0]   io_coef_out_payload_0_45_49_real,
  output     [15:0]   io_coef_out_payload_0_45_49_imag,
  output     [15:0]   io_coef_out_payload_0_46_0_real,
  output     [15:0]   io_coef_out_payload_0_46_0_imag,
  output     [15:0]   io_coef_out_payload_0_46_1_real,
  output     [15:0]   io_coef_out_payload_0_46_1_imag,
  output     [15:0]   io_coef_out_payload_0_46_2_real,
  output     [15:0]   io_coef_out_payload_0_46_2_imag,
  output     [15:0]   io_coef_out_payload_0_46_3_real,
  output     [15:0]   io_coef_out_payload_0_46_3_imag,
  output     [15:0]   io_coef_out_payload_0_46_4_real,
  output     [15:0]   io_coef_out_payload_0_46_4_imag,
  output     [15:0]   io_coef_out_payload_0_46_5_real,
  output     [15:0]   io_coef_out_payload_0_46_5_imag,
  output     [15:0]   io_coef_out_payload_0_46_6_real,
  output     [15:0]   io_coef_out_payload_0_46_6_imag,
  output     [15:0]   io_coef_out_payload_0_46_7_real,
  output     [15:0]   io_coef_out_payload_0_46_7_imag,
  output     [15:0]   io_coef_out_payload_0_46_8_real,
  output     [15:0]   io_coef_out_payload_0_46_8_imag,
  output     [15:0]   io_coef_out_payload_0_46_9_real,
  output     [15:0]   io_coef_out_payload_0_46_9_imag,
  output     [15:0]   io_coef_out_payload_0_46_10_real,
  output     [15:0]   io_coef_out_payload_0_46_10_imag,
  output     [15:0]   io_coef_out_payload_0_46_11_real,
  output     [15:0]   io_coef_out_payload_0_46_11_imag,
  output     [15:0]   io_coef_out_payload_0_46_12_real,
  output     [15:0]   io_coef_out_payload_0_46_12_imag,
  output     [15:0]   io_coef_out_payload_0_46_13_real,
  output     [15:0]   io_coef_out_payload_0_46_13_imag,
  output     [15:0]   io_coef_out_payload_0_46_14_real,
  output     [15:0]   io_coef_out_payload_0_46_14_imag,
  output     [15:0]   io_coef_out_payload_0_46_15_real,
  output     [15:0]   io_coef_out_payload_0_46_15_imag,
  output     [15:0]   io_coef_out_payload_0_46_16_real,
  output     [15:0]   io_coef_out_payload_0_46_16_imag,
  output     [15:0]   io_coef_out_payload_0_46_17_real,
  output     [15:0]   io_coef_out_payload_0_46_17_imag,
  output     [15:0]   io_coef_out_payload_0_46_18_real,
  output     [15:0]   io_coef_out_payload_0_46_18_imag,
  output     [15:0]   io_coef_out_payload_0_46_19_real,
  output     [15:0]   io_coef_out_payload_0_46_19_imag,
  output     [15:0]   io_coef_out_payload_0_46_20_real,
  output     [15:0]   io_coef_out_payload_0_46_20_imag,
  output     [15:0]   io_coef_out_payload_0_46_21_real,
  output     [15:0]   io_coef_out_payload_0_46_21_imag,
  output     [15:0]   io_coef_out_payload_0_46_22_real,
  output     [15:0]   io_coef_out_payload_0_46_22_imag,
  output     [15:0]   io_coef_out_payload_0_46_23_real,
  output     [15:0]   io_coef_out_payload_0_46_23_imag,
  output     [15:0]   io_coef_out_payload_0_46_24_real,
  output     [15:0]   io_coef_out_payload_0_46_24_imag,
  output     [15:0]   io_coef_out_payload_0_46_25_real,
  output     [15:0]   io_coef_out_payload_0_46_25_imag,
  output     [15:0]   io_coef_out_payload_0_46_26_real,
  output     [15:0]   io_coef_out_payload_0_46_26_imag,
  output     [15:0]   io_coef_out_payload_0_46_27_real,
  output     [15:0]   io_coef_out_payload_0_46_27_imag,
  output     [15:0]   io_coef_out_payload_0_46_28_real,
  output     [15:0]   io_coef_out_payload_0_46_28_imag,
  output     [15:0]   io_coef_out_payload_0_46_29_real,
  output     [15:0]   io_coef_out_payload_0_46_29_imag,
  output     [15:0]   io_coef_out_payload_0_46_30_real,
  output     [15:0]   io_coef_out_payload_0_46_30_imag,
  output     [15:0]   io_coef_out_payload_0_46_31_real,
  output     [15:0]   io_coef_out_payload_0_46_31_imag,
  output     [15:0]   io_coef_out_payload_0_46_32_real,
  output     [15:0]   io_coef_out_payload_0_46_32_imag,
  output     [15:0]   io_coef_out_payload_0_46_33_real,
  output     [15:0]   io_coef_out_payload_0_46_33_imag,
  output     [15:0]   io_coef_out_payload_0_46_34_real,
  output     [15:0]   io_coef_out_payload_0_46_34_imag,
  output     [15:0]   io_coef_out_payload_0_46_35_real,
  output     [15:0]   io_coef_out_payload_0_46_35_imag,
  output     [15:0]   io_coef_out_payload_0_46_36_real,
  output     [15:0]   io_coef_out_payload_0_46_36_imag,
  output     [15:0]   io_coef_out_payload_0_46_37_real,
  output     [15:0]   io_coef_out_payload_0_46_37_imag,
  output     [15:0]   io_coef_out_payload_0_46_38_real,
  output     [15:0]   io_coef_out_payload_0_46_38_imag,
  output     [15:0]   io_coef_out_payload_0_46_39_real,
  output     [15:0]   io_coef_out_payload_0_46_39_imag,
  output     [15:0]   io_coef_out_payload_0_46_40_real,
  output     [15:0]   io_coef_out_payload_0_46_40_imag,
  output     [15:0]   io_coef_out_payload_0_46_41_real,
  output     [15:0]   io_coef_out_payload_0_46_41_imag,
  output     [15:0]   io_coef_out_payload_0_46_42_real,
  output     [15:0]   io_coef_out_payload_0_46_42_imag,
  output     [15:0]   io_coef_out_payload_0_46_43_real,
  output     [15:0]   io_coef_out_payload_0_46_43_imag,
  output     [15:0]   io_coef_out_payload_0_46_44_real,
  output     [15:0]   io_coef_out_payload_0_46_44_imag,
  output     [15:0]   io_coef_out_payload_0_46_45_real,
  output     [15:0]   io_coef_out_payload_0_46_45_imag,
  output     [15:0]   io_coef_out_payload_0_46_46_real,
  output     [15:0]   io_coef_out_payload_0_46_46_imag,
  output     [15:0]   io_coef_out_payload_0_46_47_real,
  output     [15:0]   io_coef_out_payload_0_46_47_imag,
  output     [15:0]   io_coef_out_payload_0_46_48_real,
  output     [15:0]   io_coef_out_payload_0_46_48_imag,
  output     [15:0]   io_coef_out_payload_0_46_49_real,
  output     [15:0]   io_coef_out_payload_0_46_49_imag,
  output     [15:0]   io_coef_out_payload_0_47_0_real,
  output     [15:0]   io_coef_out_payload_0_47_0_imag,
  output     [15:0]   io_coef_out_payload_0_47_1_real,
  output     [15:0]   io_coef_out_payload_0_47_1_imag,
  output     [15:0]   io_coef_out_payload_0_47_2_real,
  output     [15:0]   io_coef_out_payload_0_47_2_imag,
  output     [15:0]   io_coef_out_payload_0_47_3_real,
  output     [15:0]   io_coef_out_payload_0_47_3_imag,
  output     [15:0]   io_coef_out_payload_0_47_4_real,
  output     [15:0]   io_coef_out_payload_0_47_4_imag,
  output     [15:0]   io_coef_out_payload_0_47_5_real,
  output     [15:0]   io_coef_out_payload_0_47_5_imag,
  output     [15:0]   io_coef_out_payload_0_47_6_real,
  output     [15:0]   io_coef_out_payload_0_47_6_imag,
  output     [15:0]   io_coef_out_payload_0_47_7_real,
  output     [15:0]   io_coef_out_payload_0_47_7_imag,
  output     [15:0]   io_coef_out_payload_0_47_8_real,
  output     [15:0]   io_coef_out_payload_0_47_8_imag,
  output     [15:0]   io_coef_out_payload_0_47_9_real,
  output     [15:0]   io_coef_out_payload_0_47_9_imag,
  output     [15:0]   io_coef_out_payload_0_47_10_real,
  output     [15:0]   io_coef_out_payload_0_47_10_imag,
  output     [15:0]   io_coef_out_payload_0_47_11_real,
  output     [15:0]   io_coef_out_payload_0_47_11_imag,
  output     [15:0]   io_coef_out_payload_0_47_12_real,
  output     [15:0]   io_coef_out_payload_0_47_12_imag,
  output     [15:0]   io_coef_out_payload_0_47_13_real,
  output     [15:0]   io_coef_out_payload_0_47_13_imag,
  output     [15:0]   io_coef_out_payload_0_47_14_real,
  output     [15:0]   io_coef_out_payload_0_47_14_imag,
  output     [15:0]   io_coef_out_payload_0_47_15_real,
  output     [15:0]   io_coef_out_payload_0_47_15_imag,
  output     [15:0]   io_coef_out_payload_0_47_16_real,
  output     [15:0]   io_coef_out_payload_0_47_16_imag,
  output     [15:0]   io_coef_out_payload_0_47_17_real,
  output     [15:0]   io_coef_out_payload_0_47_17_imag,
  output     [15:0]   io_coef_out_payload_0_47_18_real,
  output     [15:0]   io_coef_out_payload_0_47_18_imag,
  output     [15:0]   io_coef_out_payload_0_47_19_real,
  output     [15:0]   io_coef_out_payload_0_47_19_imag,
  output     [15:0]   io_coef_out_payload_0_47_20_real,
  output     [15:0]   io_coef_out_payload_0_47_20_imag,
  output     [15:0]   io_coef_out_payload_0_47_21_real,
  output     [15:0]   io_coef_out_payload_0_47_21_imag,
  output     [15:0]   io_coef_out_payload_0_47_22_real,
  output     [15:0]   io_coef_out_payload_0_47_22_imag,
  output     [15:0]   io_coef_out_payload_0_47_23_real,
  output     [15:0]   io_coef_out_payload_0_47_23_imag,
  output     [15:0]   io_coef_out_payload_0_47_24_real,
  output     [15:0]   io_coef_out_payload_0_47_24_imag,
  output     [15:0]   io_coef_out_payload_0_47_25_real,
  output     [15:0]   io_coef_out_payload_0_47_25_imag,
  output     [15:0]   io_coef_out_payload_0_47_26_real,
  output     [15:0]   io_coef_out_payload_0_47_26_imag,
  output     [15:0]   io_coef_out_payload_0_47_27_real,
  output     [15:0]   io_coef_out_payload_0_47_27_imag,
  output     [15:0]   io_coef_out_payload_0_47_28_real,
  output     [15:0]   io_coef_out_payload_0_47_28_imag,
  output     [15:0]   io_coef_out_payload_0_47_29_real,
  output     [15:0]   io_coef_out_payload_0_47_29_imag,
  output     [15:0]   io_coef_out_payload_0_47_30_real,
  output     [15:0]   io_coef_out_payload_0_47_30_imag,
  output     [15:0]   io_coef_out_payload_0_47_31_real,
  output     [15:0]   io_coef_out_payload_0_47_31_imag,
  output     [15:0]   io_coef_out_payload_0_47_32_real,
  output     [15:0]   io_coef_out_payload_0_47_32_imag,
  output     [15:0]   io_coef_out_payload_0_47_33_real,
  output     [15:0]   io_coef_out_payload_0_47_33_imag,
  output     [15:0]   io_coef_out_payload_0_47_34_real,
  output     [15:0]   io_coef_out_payload_0_47_34_imag,
  output     [15:0]   io_coef_out_payload_0_47_35_real,
  output     [15:0]   io_coef_out_payload_0_47_35_imag,
  output     [15:0]   io_coef_out_payload_0_47_36_real,
  output     [15:0]   io_coef_out_payload_0_47_36_imag,
  output     [15:0]   io_coef_out_payload_0_47_37_real,
  output     [15:0]   io_coef_out_payload_0_47_37_imag,
  output     [15:0]   io_coef_out_payload_0_47_38_real,
  output     [15:0]   io_coef_out_payload_0_47_38_imag,
  output     [15:0]   io_coef_out_payload_0_47_39_real,
  output     [15:0]   io_coef_out_payload_0_47_39_imag,
  output     [15:0]   io_coef_out_payload_0_47_40_real,
  output     [15:0]   io_coef_out_payload_0_47_40_imag,
  output     [15:0]   io_coef_out_payload_0_47_41_real,
  output     [15:0]   io_coef_out_payload_0_47_41_imag,
  output     [15:0]   io_coef_out_payload_0_47_42_real,
  output     [15:0]   io_coef_out_payload_0_47_42_imag,
  output     [15:0]   io_coef_out_payload_0_47_43_real,
  output     [15:0]   io_coef_out_payload_0_47_43_imag,
  output     [15:0]   io_coef_out_payload_0_47_44_real,
  output     [15:0]   io_coef_out_payload_0_47_44_imag,
  output     [15:0]   io_coef_out_payload_0_47_45_real,
  output     [15:0]   io_coef_out_payload_0_47_45_imag,
  output     [15:0]   io_coef_out_payload_0_47_46_real,
  output     [15:0]   io_coef_out_payload_0_47_46_imag,
  output     [15:0]   io_coef_out_payload_0_47_47_real,
  output     [15:0]   io_coef_out_payload_0_47_47_imag,
  output     [15:0]   io_coef_out_payload_0_47_48_real,
  output     [15:0]   io_coef_out_payload_0_47_48_imag,
  output     [15:0]   io_coef_out_payload_0_47_49_real,
  output     [15:0]   io_coef_out_payload_0_47_49_imag,
  output     [15:0]   io_coef_out_payload_0_48_0_real,
  output     [15:0]   io_coef_out_payload_0_48_0_imag,
  output     [15:0]   io_coef_out_payload_0_48_1_real,
  output     [15:0]   io_coef_out_payload_0_48_1_imag,
  output     [15:0]   io_coef_out_payload_0_48_2_real,
  output     [15:0]   io_coef_out_payload_0_48_2_imag,
  output     [15:0]   io_coef_out_payload_0_48_3_real,
  output     [15:0]   io_coef_out_payload_0_48_3_imag,
  output     [15:0]   io_coef_out_payload_0_48_4_real,
  output     [15:0]   io_coef_out_payload_0_48_4_imag,
  output     [15:0]   io_coef_out_payload_0_48_5_real,
  output     [15:0]   io_coef_out_payload_0_48_5_imag,
  output     [15:0]   io_coef_out_payload_0_48_6_real,
  output     [15:0]   io_coef_out_payload_0_48_6_imag,
  output     [15:0]   io_coef_out_payload_0_48_7_real,
  output     [15:0]   io_coef_out_payload_0_48_7_imag,
  output     [15:0]   io_coef_out_payload_0_48_8_real,
  output     [15:0]   io_coef_out_payload_0_48_8_imag,
  output     [15:0]   io_coef_out_payload_0_48_9_real,
  output     [15:0]   io_coef_out_payload_0_48_9_imag,
  output     [15:0]   io_coef_out_payload_0_48_10_real,
  output     [15:0]   io_coef_out_payload_0_48_10_imag,
  output     [15:0]   io_coef_out_payload_0_48_11_real,
  output     [15:0]   io_coef_out_payload_0_48_11_imag,
  output     [15:0]   io_coef_out_payload_0_48_12_real,
  output     [15:0]   io_coef_out_payload_0_48_12_imag,
  output     [15:0]   io_coef_out_payload_0_48_13_real,
  output     [15:0]   io_coef_out_payload_0_48_13_imag,
  output     [15:0]   io_coef_out_payload_0_48_14_real,
  output     [15:0]   io_coef_out_payload_0_48_14_imag,
  output     [15:0]   io_coef_out_payload_0_48_15_real,
  output     [15:0]   io_coef_out_payload_0_48_15_imag,
  output     [15:0]   io_coef_out_payload_0_48_16_real,
  output     [15:0]   io_coef_out_payload_0_48_16_imag,
  output     [15:0]   io_coef_out_payload_0_48_17_real,
  output     [15:0]   io_coef_out_payload_0_48_17_imag,
  output     [15:0]   io_coef_out_payload_0_48_18_real,
  output     [15:0]   io_coef_out_payload_0_48_18_imag,
  output     [15:0]   io_coef_out_payload_0_48_19_real,
  output     [15:0]   io_coef_out_payload_0_48_19_imag,
  output     [15:0]   io_coef_out_payload_0_48_20_real,
  output     [15:0]   io_coef_out_payload_0_48_20_imag,
  output     [15:0]   io_coef_out_payload_0_48_21_real,
  output     [15:0]   io_coef_out_payload_0_48_21_imag,
  output     [15:0]   io_coef_out_payload_0_48_22_real,
  output     [15:0]   io_coef_out_payload_0_48_22_imag,
  output     [15:0]   io_coef_out_payload_0_48_23_real,
  output     [15:0]   io_coef_out_payload_0_48_23_imag,
  output     [15:0]   io_coef_out_payload_0_48_24_real,
  output     [15:0]   io_coef_out_payload_0_48_24_imag,
  output     [15:0]   io_coef_out_payload_0_48_25_real,
  output     [15:0]   io_coef_out_payload_0_48_25_imag,
  output     [15:0]   io_coef_out_payload_0_48_26_real,
  output     [15:0]   io_coef_out_payload_0_48_26_imag,
  output     [15:0]   io_coef_out_payload_0_48_27_real,
  output     [15:0]   io_coef_out_payload_0_48_27_imag,
  output     [15:0]   io_coef_out_payload_0_48_28_real,
  output     [15:0]   io_coef_out_payload_0_48_28_imag,
  output     [15:0]   io_coef_out_payload_0_48_29_real,
  output     [15:0]   io_coef_out_payload_0_48_29_imag,
  output     [15:0]   io_coef_out_payload_0_48_30_real,
  output     [15:0]   io_coef_out_payload_0_48_30_imag,
  output     [15:0]   io_coef_out_payload_0_48_31_real,
  output     [15:0]   io_coef_out_payload_0_48_31_imag,
  output     [15:0]   io_coef_out_payload_0_48_32_real,
  output     [15:0]   io_coef_out_payload_0_48_32_imag,
  output     [15:0]   io_coef_out_payload_0_48_33_real,
  output     [15:0]   io_coef_out_payload_0_48_33_imag,
  output     [15:0]   io_coef_out_payload_0_48_34_real,
  output     [15:0]   io_coef_out_payload_0_48_34_imag,
  output     [15:0]   io_coef_out_payload_0_48_35_real,
  output     [15:0]   io_coef_out_payload_0_48_35_imag,
  output     [15:0]   io_coef_out_payload_0_48_36_real,
  output     [15:0]   io_coef_out_payload_0_48_36_imag,
  output     [15:0]   io_coef_out_payload_0_48_37_real,
  output     [15:0]   io_coef_out_payload_0_48_37_imag,
  output     [15:0]   io_coef_out_payload_0_48_38_real,
  output     [15:0]   io_coef_out_payload_0_48_38_imag,
  output     [15:0]   io_coef_out_payload_0_48_39_real,
  output     [15:0]   io_coef_out_payload_0_48_39_imag,
  output     [15:0]   io_coef_out_payload_0_48_40_real,
  output     [15:0]   io_coef_out_payload_0_48_40_imag,
  output     [15:0]   io_coef_out_payload_0_48_41_real,
  output     [15:0]   io_coef_out_payload_0_48_41_imag,
  output     [15:0]   io_coef_out_payload_0_48_42_real,
  output     [15:0]   io_coef_out_payload_0_48_42_imag,
  output     [15:0]   io_coef_out_payload_0_48_43_real,
  output     [15:0]   io_coef_out_payload_0_48_43_imag,
  output     [15:0]   io_coef_out_payload_0_48_44_real,
  output     [15:0]   io_coef_out_payload_0_48_44_imag,
  output     [15:0]   io_coef_out_payload_0_48_45_real,
  output     [15:0]   io_coef_out_payload_0_48_45_imag,
  output     [15:0]   io_coef_out_payload_0_48_46_real,
  output     [15:0]   io_coef_out_payload_0_48_46_imag,
  output     [15:0]   io_coef_out_payload_0_48_47_real,
  output     [15:0]   io_coef_out_payload_0_48_47_imag,
  output     [15:0]   io_coef_out_payload_0_48_48_real,
  output     [15:0]   io_coef_out_payload_0_48_48_imag,
  output     [15:0]   io_coef_out_payload_0_48_49_real,
  output     [15:0]   io_coef_out_payload_0_48_49_imag,
  output     [15:0]   io_coef_out_payload_0_49_0_real,
  output     [15:0]   io_coef_out_payload_0_49_0_imag,
  output     [15:0]   io_coef_out_payload_0_49_1_real,
  output     [15:0]   io_coef_out_payload_0_49_1_imag,
  output     [15:0]   io_coef_out_payload_0_49_2_real,
  output     [15:0]   io_coef_out_payload_0_49_2_imag,
  output     [15:0]   io_coef_out_payload_0_49_3_real,
  output     [15:0]   io_coef_out_payload_0_49_3_imag,
  output     [15:0]   io_coef_out_payload_0_49_4_real,
  output     [15:0]   io_coef_out_payload_0_49_4_imag,
  output     [15:0]   io_coef_out_payload_0_49_5_real,
  output     [15:0]   io_coef_out_payload_0_49_5_imag,
  output     [15:0]   io_coef_out_payload_0_49_6_real,
  output     [15:0]   io_coef_out_payload_0_49_6_imag,
  output     [15:0]   io_coef_out_payload_0_49_7_real,
  output     [15:0]   io_coef_out_payload_0_49_7_imag,
  output     [15:0]   io_coef_out_payload_0_49_8_real,
  output     [15:0]   io_coef_out_payload_0_49_8_imag,
  output     [15:0]   io_coef_out_payload_0_49_9_real,
  output     [15:0]   io_coef_out_payload_0_49_9_imag,
  output     [15:0]   io_coef_out_payload_0_49_10_real,
  output     [15:0]   io_coef_out_payload_0_49_10_imag,
  output     [15:0]   io_coef_out_payload_0_49_11_real,
  output     [15:0]   io_coef_out_payload_0_49_11_imag,
  output     [15:0]   io_coef_out_payload_0_49_12_real,
  output     [15:0]   io_coef_out_payload_0_49_12_imag,
  output     [15:0]   io_coef_out_payload_0_49_13_real,
  output     [15:0]   io_coef_out_payload_0_49_13_imag,
  output     [15:0]   io_coef_out_payload_0_49_14_real,
  output     [15:0]   io_coef_out_payload_0_49_14_imag,
  output     [15:0]   io_coef_out_payload_0_49_15_real,
  output     [15:0]   io_coef_out_payload_0_49_15_imag,
  output     [15:0]   io_coef_out_payload_0_49_16_real,
  output     [15:0]   io_coef_out_payload_0_49_16_imag,
  output     [15:0]   io_coef_out_payload_0_49_17_real,
  output     [15:0]   io_coef_out_payload_0_49_17_imag,
  output     [15:0]   io_coef_out_payload_0_49_18_real,
  output     [15:0]   io_coef_out_payload_0_49_18_imag,
  output     [15:0]   io_coef_out_payload_0_49_19_real,
  output     [15:0]   io_coef_out_payload_0_49_19_imag,
  output     [15:0]   io_coef_out_payload_0_49_20_real,
  output     [15:0]   io_coef_out_payload_0_49_20_imag,
  output     [15:0]   io_coef_out_payload_0_49_21_real,
  output     [15:0]   io_coef_out_payload_0_49_21_imag,
  output     [15:0]   io_coef_out_payload_0_49_22_real,
  output     [15:0]   io_coef_out_payload_0_49_22_imag,
  output     [15:0]   io_coef_out_payload_0_49_23_real,
  output     [15:0]   io_coef_out_payload_0_49_23_imag,
  output     [15:0]   io_coef_out_payload_0_49_24_real,
  output     [15:0]   io_coef_out_payload_0_49_24_imag,
  output     [15:0]   io_coef_out_payload_0_49_25_real,
  output     [15:0]   io_coef_out_payload_0_49_25_imag,
  output     [15:0]   io_coef_out_payload_0_49_26_real,
  output     [15:0]   io_coef_out_payload_0_49_26_imag,
  output     [15:0]   io_coef_out_payload_0_49_27_real,
  output     [15:0]   io_coef_out_payload_0_49_27_imag,
  output     [15:0]   io_coef_out_payload_0_49_28_real,
  output     [15:0]   io_coef_out_payload_0_49_28_imag,
  output     [15:0]   io_coef_out_payload_0_49_29_real,
  output     [15:0]   io_coef_out_payload_0_49_29_imag,
  output     [15:0]   io_coef_out_payload_0_49_30_real,
  output     [15:0]   io_coef_out_payload_0_49_30_imag,
  output     [15:0]   io_coef_out_payload_0_49_31_real,
  output     [15:0]   io_coef_out_payload_0_49_31_imag,
  output     [15:0]   io_coef_out_payload_0_49_32_real,
  output     [15:0]   io_coef_out_payload_0_49_32_imag,
  output     [15:0]   io_coef_out_payload_0_49_33_real,
  output     [15:0]   io_coef_out_payload_0_49_33_imag,
  output     [15:0]   io_coef_out_payload_0_49_34_real,
  output     [15:0]   io_coef_out_payload_0_49_34_imag,
  output     [15:0]   io_coef_out_payload_0_49_35_real,
  output     [15:0]   io_coef_out_payload_0_49_35_imag,
  output     [15:0]   io_coef_out_payload_0_49_36_real,
  output     [15:0]   io_coef_out_payload_0_49_36_imag,
  output     [15:0]   io_coef_out_payload_0_49_37_real,
  output     [15:0]   io_coef_out_payload_0_49_37_imag,
  output     [15:0]   io_coef_out_payload_0_49_38_real,
  output     [15:0]   io_coef_out_payload_0_49_38_imag,
  output     [15:0]   io_coef_out_payload_0_49_39_real,
  output     [15:0]   io_coef_out_payload_0_49_39_imag,
  output     [15:0]   io_coef_out_payload_0_49_40_real,
  output     [15:0]   io_coef_out_payload_0_49_40_imag,
  output     [15:0]   io_coef_out_payload_0_49_41_real,
  output     [15:0]   io_coef_out_payload_0_49_41_imag,
  output     [15:0]   io_coef_out_payload_0_49_42_real,
  output     [15:0]   io_coef_out_payload_0_49_42_imag,
  output     [15:0]   io_coef_out_payload_0_49_43_real,
  output     [15:0]   io_coef_out_payload_0_49_43_imag,
  output     [15:0]   io_coef_out_payload_0_49_44_real,
  output     [15:0]   io_coef_out_payload_0_49_44_imag,
  output     [15:0]   io_coef_out_payload_0_49_45_real,
  output     [15:0]   io_coef_out_payload_0_49_45_imag,
  output     [15:0]   io_coef_out_payload_0_49_46_real,
  output     [15:0]   io_coef_out_payload_0_49_46_imag,
  output     [15:0]   io_coef_out_payload_0_49_47_real,
  output     [15:0]   io_coef_out_payload_0_49_47_imag,
  output     [15:0]   io_coef_out_payload_0_49_48_real,
  output     [15:0]   io_coef_out_payload_0_49_48_imag,
  output     [15:0]   io_coef_out_payload_0_49_49_real,
  output     [15:0]   io_coef_out_payload_0_49_49_imag,
  input               clk,
  input               reset 
);
  reg        [11:0]   _zz_4433_;
  reg        [15:0]   _zz_4434_;
  reg        [15:0]   _zz_4435_;
  reg        [15:0]   _zz_4436_;
  reg        [15:0]   _zz_4437_;
  reg        [15:0]   _zz_4438_;
  reg        [15:0]   _zz_4439_;
  reg        [15:0]   _zz_4440_;
  reg        [15:0]   _zz_4441_;
  reg        [15:0]   _zz_4442_;
  reg        [15:0]   _zz_4443_;
  reg        [15:0]   _zz_4444_;
  reg        [15:0]   _zz_4445_;
  reg        [15:0]   _zz_4446_;
  reg        [15:0]   _zz_4447_;
  reg        [15:0]   _zz_4448_;
  reg        [15:0]   _zz_4449_;
  reg        [15:0]   _zz_4450_;
  reg        [15:0]   _zz_4451_;
  reg        [15:0]   _zz_4452_;
  reg        [15:0]   _zz_4453_;
  reg        [15:0]   _zz_4454_;
  reg        [15:0]   _zz_4455_;
  reg        [15:0]   _zz_4456_;
  reg        [15:0]   _zz_4457_;
  reg        [15:0]   _zz_4458_;
  reg        [15:0]   _zz_4459_;
  reg        [15:0]   _zz_4460_;
  reg        [15:0]   _zz_4461_;
  reg        [15:0]   _zz_4462_;
  reg        [15:0]   _zz_4463_;
  reg        [15:0]   _zz_4464_;
  reg        [15:0]   _zz_4465_;
  reg        [15:0]   _zz_4466_;
  reg        [15:0]   _zz_4467_;
  reg        [15:0]   _zz_4468_;
  reg        [15:0]   _zz_4469_;
  reg        [15:0]   _zz_4470_;
  reg        [15:0]   _zz_4471_;
  reg        [15:0]   _zz_4472_;
  reg        [15:0]   _zz_4473_;
  reg        [15:0]   _zz_4474_;
  reg        [15:0]   _zz_4475_;
  reg        [15:0]   _zz_4476_;
  reg        [15:0]   _zz_4477_;
  reg        [15:0]   _zz_4478_;
  reg        [15:0]   _zz_4479_;
  reg        [15:0]   _zz_4480_;
  reg        [15:0]   _zz_4481_;
  reg        [15:0]   _zz_4482_;
  reg        [15:0]   _zz_4483_;
  reg        [15:0]   _zz_4484_;
  reg        [15:0]   _zz_4485_;
  reg        [15:0]   _zz_4486_;
  reg        [15:0]   _zz_4487_;
  reg        [15:0]   _zz_4488_;
  reg        [15:0]   _zz_4489_;
  reg        [15:0]   _zz_4490_;
  reg        [15:0]   _zz_4491_;
  reg        [15:0]   _zz_4492_;
  reg        [15:0]   _zz_4493_;
  reg        [15:0]   _zz_4494_;
  reg        [15:0]   _zz_4495_;
  reg        [15:0]   _zz_4496_;
  reg        [15:0]   _zz_4497_;
  reg        [15:0]   _zz_4498_;
  reg        [15:0]   _zz_4499_;
  reg        [15:0]   _zz_4500_;
  reg        [15:0]   _zz_4501_;
  reg        [15:0]   _zz_4502_;
  reg        [15:0]   _zz_4503_;
  reg        [15:0]   _zz_4504_;
  reg        [15:0]   _zz_4505_;
  reg        [15:0]   _zz_4506_;
  reg        [15:0]   _zz_4507_;
  reg        [15:0]   _zz_4508_;
  reg        [15:0]   _zz_4509_;
  reg        [15:0]   _zz_4510_;
  reg        [15:0]   _zz_4511_;
  reg        [15:0]   _zz_4512_;
  reg        [15:0]   _zz_4513_;
  reg        [15:0]   _zz_4514_;
  reg        [15:0]   _zz_4515_;
  reg        [15:0]   _zz_4516_;
  reg        [15:0]   _zz_4517_;
  reg        [15:0]   _zz_4518_;
  reg        [15:0]   _zz_4519_;
  reg        [15:0]   _zz_4520_;
  reg        [15:0]   _zz_4521_;
  reg        [15:0]   _zz_4522_;
  reg        [15:0]   _zz_4523_;
  reg        [15:0]   _zz_4524_;
  reg        [15:0]   _zz_4525_;
  reg        [15:0]   _zz_4526_;
  reg        [15:0]   _zz_4527_;
  reg        [15:0]   _zz_4528_;
  reg        [15:0]   _zz_4529_;
  reg        [15:0]   _zz_4530_;
  reg        [15:0]   _zz_4531_;
  reg        [15:0]   _zz_4532_;
  reg        [15:0]   _zz_4533_;
  reg        [15:0]   _zz_4534_;
  reg        [15:0]   _zz_4535_;
  reg        [15:0]   _zz_4536_;
  reg        [15:0]   _zz_4537_;
  reg        [15:0]   _zz_4538_;
  reg        [15:0]   _zz_4539_;
  reg        [15:0]   _zz_4540_;
  reg        [15:0]   _zz_4541_;
  reg        [15:0]   _zz_4542_;
  reg        [15:0]   _zz_4543_;
  reg        [15:0]   _zz_4544_;
  reg        [15:0]   _zz_4545_;
  reg        [15:0]   _zz_4546_;
  reg        [15:0]   _zz_4547_;
  reg        [15:0]   _zz_4548_;
  reg        [15:0]   _zz_4549_;
  reg        [15:0]   _zz_4550_;
  reg        [15:0]   _zz_4551_;
  reg        [15:0]   _zz_4552_;
  reg        [15:0]   _zz_4553_;
  reg        [15:0]   _zz_4554_;
  reg        [15:0]   _zz_4555_;
  reg        [15:0]   _zz_4556_;
  reg        [15:0]   _zz_4557_;
  reg        [15:0]   _zz_4558_;
  reg        [15:0]   _zz_4559_;
  reg        [15:0]   _zz_4560_;
  reg        [15:0]   _zz_4561_;
  wire       [11:0]   _zz_4562_;
  wire       [11:0]   _zz_4563_;
  wire       [11:0]   _zz_4564_;
  wire       [0:0]    _zz_4565_;
  wire       [31:0]   _zz_4566_;
  wire       [31:0]   _zz_4567_;
  wire       [31:0]   _zz_4568_;
  wire       [31:0]   _zz_4569_;
  wire       [31:0]   _zz_4570_;
  wire       [31:0]   _zz_4571_;
  wire       [31:0]   _zz_4572_;
  wire       [31:0]   _zz_4573_;
  wire       [31:0]   _zz_4574_;
  wire       [31:0]   _zz_4575_;
  wire       [31:0]   _zz_4576_;
  wire       [31:0]   _zz_4577_;
  wire       [31:0]   _zz_4578_;
  wire       [31:0]   _zz_4579_;
  wire       [31:0]   _zz_4580_;
  wire       [31:0]   _zz_4581_;
  wire       [31:0]   _zz_4582_;
  wire       [31:0]   _zz_4583_;
  wire       [31:0]   _zz_4584_;
  wire       [31:0]   _zz_4585_;
  wire       [31:0]   _zz_4586_;
  wire       [31:0]   _zz_4587_;
  wire       [31:0]   _zz_4588_;
  wire       [31:0]   _zz_4589_;
  wire       [31:0]   _zz_4590_;
  wire       [31:0]   _zz_4591_;
  wire       [31:0]   _zz_4592_;
  wire       [31:0]   _zz_4593_;
  wire       [31:0]   _zz_4594_;
  wire       [31:0]   _zz_4595_;
  wire       [31:0]   _zz_4596_;
  wire       [31:0]   _zz_4597_;
  wire       [31:0]   _zz_4598_;
  wire       [31:0]   _zz_4599_;
  wire       [31:0]   _zz_4600_;
  wire       [31:0]   _zz_4601_;
  wire       [31:0]   _zz_4602_;
  wire       [31:0]   _zz_4603_;
  wire       [31:0]   _zz_4604_;
  wire       [31:0]   _zz_4605_;
  wire       [31:0]   _zz_4606_;
  wire       [31:0]   _zz_4607_;
  wire       [31:0]   _zz_4608_;
  wire       [31:0]   _zz_4609_;
  wire       [31:0]   _zz_4610_;
  wire       [31:0]   _zz_4611_;
  wire       [31:0]   _zz_4612_;
  wire       [31:0]   _zz_4613_;
  wire       [31:0]   _zz_4614_;
  wire       [31:0]   _zz_4615_;
  wire       [31:0]   _zz_4616_;
  wire       [31:0]   _zz_4617_;
  wire       [31:0]   _zz_4618_;
  wire       [31:0]   _zz_4619_;
  wire       [31:0]   _zz_4620_;
  wire       [31:0]   _zz_4621_;
  wire       [31:0]   _zz_4622_;
  wire       [31:0]   _zz_4623_;
  wire       [31:0]   _zz_4624_;
  wire       [31:0]   _zz_4625_;
  wire       [31:0]   _zz_4626_;
  wire       [31:0]   _zz_4627_;
  wire       [31:0]   _zz_4628_;
  wire       [31:0]   _zz_4629_;
  reg        [31:0]   _zz_13_;
  reg        [7:0]    _zz_14_;
  reg        [3:0]    _zz_15_;
  reg                 transfer_done;
  reg        [15:0]   int_reg_array_0_0_real;
  reg        [15:0]   int_reg_array_0_0_imag;
  reg        [15:0]   int_reg_array_0_1_real;
  reg        [15:0]   int_reg_array_0_1_imag;
  reg        [15:0]   int_reg_array_0_2_real;
  reg        [15:0]   int_reg_array_0_2_imag;
  reg        [15:0]   int_reg_array_0_3_real;
  reg        [15:0]   int_reg_array_0_3_imag;
  reg        [15:0]   int_reg_array_0_4_real;
  reg        [15:0]   int_reg_array_0_4_imag;
  reg        [15:0]   int_reg_array_0_5_real;
  reg        [15:0]   int_reg_array_0_5_imag;
  reg        [15:0]   int_reg_array_0_6_real;
  reg        [15:0]   int_reg_array_0_6_imag;
  reg        [15:0]   int_reg_array_0_7_real;
  reg        [15:0]   int_reg_array_0_7_imag;
  reg        [15:0]   int_reg_array_0_8_real;
  reg        [15:0]   int_reg_array_0_8_imag;
  reg        [15:0]   int_reg_array_0_9_real;
  reg        [15:0]   int_reg_array_0_9_imag;
  reg        [15:0]   int_reg_array_0_10_real;
  reg        [15:0]   int_reg_array_0_10_imag;
  reg        [15:0]   int_reg_array_0_11_real;
  reg        [15:0]   int_reg_array_0_11_imag;
  reg        [15:0]   int_reg_array_0_12_real;
  reg        [15:0]   int_reg_array_0_12_imag;
  reg        [15:0]   int_reg_array_0_13_real;
  reg        [15:0]   int_reg_array_0_13_imag;
  reg        [15:0]   int_reg_array_0_14_real;
  reg        [15:0]   int_reg_array_0_14_imag;
  reg        [15:0]   int_reg_array_0_15_real;
  reg        [15:0]   int_reg_array_0_15_imag;
  reg        [15:0]   int_reg_array_0_16_real;
  reg        [15:0]   int_reg_array_0_16_imag;
  reg        [15:0]   int_reg_array_0_17_real;
  reg        [15:0]   int_reg_array_0_17_imag;
  reg        [15:0]   int_reg_array_0_18_real;
  reg        [15:0]   int_reg_array_0_18_imag;
  reg        [15:0]   int_reg_array_0_19_real;
  reg        [15:0]   int_reg_array_0_19_imag;
  reg        [15:0]   int_reg_array_0_20_real;
  reg        [15:0]   int_reg_array_0_20_imag;
  reg        [15:0]   int_reg_array_0_21_real;
  reg        [15:0]   int_reg_array_0_21_imag;
  reg        [15:0]   int_reg_array_0_22_real;
  reg        [15:0]   int_reg_array_0_22_imag;
  reg        [15:0]   int_reg_array_0_23_real;
  reg        [15:0]   int_reg_array_0_23_imag;
  reg        [15:0]   int_reg_array_0_24_real;
  reg        [15:0]   int_reg_array_0_24_imag;
  reg        [15:0]   int_reg_array_0_25_real;
  reg        [15:0]   int_reg_array_0_25_imag;
  reg        [15:0]   int_reg_array_0_26_real;
  reg        [15:0]   int_reg_array_0_26_imag;
  reg        [15:0]   int_reg_array_0_27_real;
  reg        [15:0]   int_reg_array_0_27_imag;
  reg        [15:0]   int_reg_array_0_28_real;
  reg        [15:0]   int_reg_array_0_28_imag;
  reg        [15:0]   int_reg_array_0_29_real;
  reg        [15:0]   int_reg_array_0_29_imag;
  reg        [15:0]   int_reg_array_0_30_real;
  reg        [15:0]   int_reg_array_0_30_imag;
  reg        [15:0]   int_reg_array_0_31_real;
  reg        [15:0]   int_reg_array_0_31_imag;
  reg        [15:0]   int_reg_array_0_32_real;
  reg        [15:0]   int_reg_array_0_32_imag;
  reg        [15:0]   int_reg_array_0_33_real;
  reg        [15:0]   int_reg_array_0_33_imag;
  reg        [15:0]   int_reg_array_0_34_real;
  reg        [15:0]   int_reg_array_0_34_imag;
  reg        [15:0]   int_reg_array_0_35_real;
  reg        [15:0]   int_reg_array_0_35_imag;
  reg        [15:0]   int_reg_array_0_36_real;
  reg        [15:0]   int_reg_array_0_36_imag;
  reg        [15:0]   int_reg_array_0_37_real;
  reg        [15:0]   int_reg_array_0_37_imag;
  reg        [15:0]   int_reg_array_0_38_real;
  reg        [15:0]   int_reg_array_0_38_imag;
  reg        [15:0]   int_reg_array_0_39_real;
  reg        [15:0]   int_reg_array_0_39_imag;
  reg        [15:0]   int_reg_array_0_40_real;
  reg        [15:0]   int_reg_array_0_40_imag;
  reg        [15:0]   int_reg_array_0_41_real;
  reg        [15:0]   int_reg_array_0_41_imag;
  reg        [15:0]   int_reg_array_0_42_real;
  reg        [15:0]   int_reg_array_0_42_imag;
  reg        [15:0]   int_reg_array_0_43_real;
  reg        [15:0]   int_reg_array_0_43_imag;
  reg        [15:0]   int_reg_array_0_44_real;
  reg        [15:0]   int_reg_array_0_44_imag;
  reg        [15:0]   int_reg_array_0_45_real;
  reg        [15:0]   int_reg_array_0_45_imag;
  reg        [15:0]   int_reg_array_0_46_real;
  reg        [15:0]   int_reg_array_0_46_imag;
  reg        [15:0]   int_reg_array_0_47_real;
  reg        [15:0]   int_reg_array_0_47_imag;
  reg        [15:0]   int_reg_array_0_48_real;
  reg        [15:0]   int_reg_array_0_48_imag;
  reg        [15:0]   int_reg_array_0_49_real;
  reg        [15:0]   int_reg_array_0_49_imag;
  reg        [15:0]   int_reg_array_0_50_real;
  reg        [15:0]   int_reg_array_0_50_imag;
  reg        [15:0]   int_reg_array_0_51_real;
  reg        [15:0]   int_reg_array_0_51_imag;
  reg        [15:0]   int_reg_array_0_52_real;
  reg        [15:0]   int_reg_array_0_52_imag;
  reg        [15:0]   int_reg_array_0_53_real;
  reg        [15:0]   int_reg_array_0_53_imag;
  reg        [15:0]   int_reg_array_0_54_real;
  reg        [15:0]   int_reg_array_0_54_imag;
  reg        [15:0]   int_reg_array_0_55_real;
  reg        [15:0]   int_reg_array_0_55_imag;
  reg        [15:0]   int_reg_array_0_56_real;
  reg        [15:0]   int_reg_array_0_56_imag;
  reg        [15:0]   int_reg_array_0_57_real;
  reg        [15:0]   int_reg_array_0_57_imag;
  reg        [15:0]   int_reg_array_0_58_real;
  reg        [15:0]   int_reg_array_0_58_imag;
  reg        [15:0]   int_reg_array_0_59_real;
  reg        [15:0]   int_reg_array_0_59_imag;
  reg        [15:0]   int_reg_array_0_60_real;
  reg        [15:0]   int_reg_array_0_60_imag;
  reg        [15:0]   int_reg_array_0_61_real;
  reg        [15:0]   int_reg_array_0_61_imag;
  reg        [15:0]   int_reg_array_0_62_real;
  reg        [15:0]   int_reg_array_0_62_imag;
  reg        [15:0]   int_reg_array_0_63_real;
  reg        [15:0]   int_reg_array_0_63_imag;
  reg        [15:0]   int_reg_array_33_0_real;
  reg        [15:0]   int_reg_array_33_0_imag;
  reg        [15:0]   int_reg_array_33_1_real;
  reg        [15:0]   int_reg_array_33_1_imag;
  reg        [15:0]   int_reg_array_33_2_real;
  reg        [15:0]   int_reg_array_33_2_imag;
  reg        [15:0]   int_reg_array_33_3_real;
  reg        [15:0]   int_reg_array_33_3_imag;
  reg        [15:0]   int_reg_array_33_4_real;
  reg        [15:0]   int_reg_array_33_4_imag;
  reg        [15:0]   int_reg_array_33_5_real;
  reg        [15:0]   int_reg_array_33_5_imag;
  reg        [15:0]   int_reg_array_33_6_real;
  reg        [15:0]   int_reg_array_33_6_imag;
  reg        [15:0]   int_reg_array_33_7_real;
  reg        [15:0]   int_reg_array_33_7_imag;
  reg        [15:0]   int_reg_array_33_8_real;
  reg        [15:0]   int_reg_array_33_8_imag;
  reg        [15:0]   int_reg_array_33_9_real;
  reg        [15:0]   int_reg_array_33_9_imag;
  reg        [15:0]   int_reg_array_33_10_real;
  reg        [15:0]   int_reg_array_33_10_imag;
  reg        [15:0]   int_reg_array_33_11_real;
  reg        [15:0]   int_reg_array_33_11_imag;
  reg        [15:0]   int_reg_array_33_12_real;
  reg        [15:0]   int_reg_array_33_12_imag;
  reg        [15:0]   int_reg_array_33_13_real;
  reg        [15:0]   int_reg_array_33_13_imag;
  reg        [15:0]   int_reg_array_33_14_real;
  reg        [15:0]   int_reg_array_33_14_imag;
  reg        [15:0]   int_reg_array_33_15_real;
  reg        [15:0]   int_reg_array_33_15_imag;
  reg        [15:0]   int_reg_array_33_16_real;
  reg        [15:0]   int_reg_array_33_16_imag;
  reg        [15:0]   int_reg_array_33_17_real;
  reg        [15:0]   int_reg_array_33_17_imag;
  reg        [15:0]   int_reg_array_33_18_real;
  reg        [15:0]   int_reg_array_33_18_imag;
  reg        [15:0]   int_reg_array_33_19_real;
  reg        [15:0]   int_reg_array_33_19_imag;
  reg        [15:0]   int_reg_array_33_20_real;
  reg        [15:0]   int_reg_array_33_20_imag;
  reg        [15:0]   int_reg_array_33_21_real;
  reg        [15:0]   int_reg_array_33_21_imag;
  reg        [15:0]   int_reg_array_33_22_real;
  reg        [15:0]   int_reg_array_33_22_imag;
  reg        [15:0]   int_reg_array_33_23_real;
  reg        [15:0]   int_reg_array_33_23_imag;
  reg        [15:0]   int_reg_array_33_24_real;
  reg        [15:0]   int_reg_array_33_24_imag;
  reg        [15:0]   int_reg_array_33_25_real;
  reg        [15:0]   int_reg_array_33_25_imag;
  reg        [15:0]   int_reg_array_33_26_real;
  reg        [15:0]   int_reg_array_33_26_imag;
  reg        [15:0]   int_reg_array_33_27_real;
  reg        [15:0]   int_reg_array_33_27_imag;
  reg        [15:0]   int_reg_array_33_28_real;
  reg        [15:0]   int_reg_array_33_28_imag;
  reg        [15:0]   int_reg_array_33_29_real;
  reg        [15:0]   int_reg_array_33_29_imag;
  reg        [15:0]   int_reg_array_33_30_real;
  reg        [15:0]   int_reg_array_33_30_imag;
  reg        [15:0]   int_reg_array_33_31_real;
  reg        [15:0]   int_reg_array_33_31_imag;
  reg        [15:0]   int_reg_array_33_32_real;
  reg        [15:0]   int_reg_array_33_32_imag;
  reg        [15:0]   int_reg_array_33_33_real;
  reg        [15:0]   int_reg_array_33_33_imag;
  reg        [15:0]   int_reg_array_33_34_real;
  reg        [15:0]   int_reg_array_33_34_imag;
  reg        [15:0]   int_reg_array_33_35_real;
  reg        [15:0]   int_reg_array_33_35_imag;
  reg        [15:0]   int_reg_array_33_36_real;
  reg        [15:0]   int_reg_array_33_36_imag;
  reg        [15:0]   int_reg_array_33_37_real;
  reg        [15:0]   int_reg_array_33_37_imag;
  reg        [15:0]   int_reg_array_33_38_real;
  reg        [15:0]   int_reg_array_33_38_imag;
  reg        [15:0]   int_reg_array_33_39_real;
  reg        [15:0]   int_reg_array_33_39_imag;
  reg        [15:0]   int_reg_array_33_40_real;
  reg        [15:0]   int_reg_array_33_40_imag;
  reg        [15:0]   int_reg_array_33_41_real;
  reg        [15:0]   int_reg_array_33_41_imag;
  reg        [15:0]   int_reg_array_33_42_real;
  reg        [15:0]   int_reg_array_33_42_imag;
  reg        [15:0]   int_reg_array_33_43_real;
  reg        [15:0]   int_reg_array_33_43_imag;
  reg        [15:0]   int_reg_array_33_44_real;
  reg        [15:0]   int_reg_array_33_44_imag;
  reg        [15:0]   int_reg_array_33_45_real;
  reg        [15:0]   int_reg_array_33_45_imag;
  reg        [15:0]   int_reg_array_33_46_real;
  reg        [15:0]   int_reg_array_33_46_imag;
  reg        [15:0]   int_reg_array_33_47_real;
  reg        [15:0]   int_reg_array_33_47_imag;
  reg        [15:0]   int_reg_array_33_48_real;
  reg        [15:0]   int_reg_array_33_48_imag;
  reg        [15:0]   int_reg_array_33_49_real;
  reg        [15:0]   int_reg_array_33_49_imag;
  reg        [15:0]   int_reg_array_33_50_real;
  reg        [15:0]   int_reg_array_33_50_imag;
  reg        [15:0]   int_reg_array_33_51_real;
  reg        [15:0]   int_reg_array_33_51_imag;
  reg        [15:0]   int_reg_array_33_52_real;
  reg        [15:0]   int_reg_array_33_52_imag;
  reg        [15:0]   int_reg_array_33_53_real;
  reg        [15:0]   int_reg_array_33_53_imag;
  reg        [15:0]   int_reg_array_33_54_real;
  reg        [15:0]   int_reg_array_33_54_imag;
  reg        [15:0]   int_reg_array_33_55_real;
  reg        [15:0]   int_reg_array_33_55_imag;
  reg        [15:0]   int_reg_array_33_56_real;
  reg        [15:0]   int_reg_array_33_56_imag;
  reg        [15:0]   int_reg_array_33_57_real;
  reg        [15:0]   int_reg_array_33_57_imag;
  reg        [15:0]   int_reg_array_33_58_real;
  reg        [15:0]   int_reg_array_33_58_imag;
  reg        [15:0]   int_reg_array_33_59_real;
  reg        [15:0]   int_reg_array_33_59_imag;
  reg        [15:0]   int_reg_array_33_60_real;
  reg        [15:0]   int_reg_array_33_60_imag;
  reg        [15:0]   int_reg_array_33_61_real;
  reg        [15:0]   int_reg_array_33_61_imag;
  reg        [15:0]   int_reg_array_33_62_real;
  reg        [15:0]   int_reg_array_33_62_imag;
  reg        [15:0]   int_reg_array_33_63_real;
  reg        [15:0]   int_reg_array_33_63_imag;
  reg        [15:0]   int_reg_array_38_0_real;
  reg        [15:0]   int_reg_array_38_0_imag;
  reg        [15:0]   int_reg_array_38_1_real;
  reg        [15:0]   int_reg_array_38_1_imag;
  reg        [15:0]   int_reg_array_38_2_real;
  reg        [15:0]   int_reg_array_38_2_imag;
  reg        [15:0]   int_reg_array_38_3_real;
  reg        [15:0]   int_reg_array_38_3_imag;
  reg        [15:0]   int_reg_array_38_4_real;
  reg        [15:0]   int_reg_array_38_4_imag;
  reg        [15:0]   int_reg_array_38_5_real;
  reg        [15:0]   int_reg_array_38_5_imag;
  reg        [15:0]   int_reg_array_38_6_real;
  reg        [15:0]   int_reg_array_38_6_imag;
  reg        [15:0]   int_reg_array_38_7_real;
  reg        [15:0]   int_reg_array_38_7_imag;
  reg        [15:0]   int_reg_array_38_8_real;
  reg        [15:0]   int_reg_array_38_8_imag;
  reg        [15:0]   int_reg_array_38_9_real;
  reg        [15:0]   int_reg_array_38_9_imag;
  reg        [15:0]   int_reg_array_38_10_real;
  reg        [15:0]   int_reg_array_38_10_imag;
  reg        [15:0]   int_reg_array_38_11_real;
  reg        [15:0]   int_reg_array_38_11_imag;
  reg        [15:0]   int_reg_array_38_12_real;
  reg        [15:0]   int_reg_array_38_12_imag;
  reg        [15:0]   int_reg_array_38_13_real;
  reg        [15:0]   int_reg_array_38_13_imag;
  reg        [15:0]   int_reg_array_38_14_real;
  reg        [15:0]   int_reg_array_38_14_imag;
  reg        [15:0]   int_reg_array_38_15_real;
  reg        [15:0]   int_reg_array_38_15_imag;
  reg        [15:0]   int_reg_array_38_16_real;
  reg        [15:0]   int_reg_array_38_16_imag;
  reg        [15:0]   int_reg_array_38_17_real;
  reg        [15:0]   int_reg_array_38_17_imag;
  reg        [15:0]   int_reg_array_38_18_real;
  reg        [15:0]   int_reg_array_38_18_imag;
  reg        [15:0]   int_reg_array_38_19_real;
  reg        [15:0]   int_reg_array_38_19_imag;
  reg        [15:0]   int_reg_array_38_20_real;
  reg        [15:0]   int_reg_array_38_20_imag;
  reg        [15:0]   int_reg_array_38_21_real;
  reg        [15:0]   int_reg_array_38_21_imag;
  reg        [15:0]   int_reg_array_38_22_real;
  reg        [15:0]   int_reg_array_38_22_imag;
  reg        [15:0]   int_reg_array_38_23_real;
  reg        [15:0]   int_reg_array_38_23_imag;
  reg        [15:0]   int_reg_array_38_24_real;
  reg        [15:0]   int_reg_array_38_24_imag;
  reg        [15:0]   int_reg_array_38_25_real;
  reg        [15:0]   int_reg_array_38_25_imag;
  reg        [15:0]   int_reg_array_38_26_real;
  reg        [15:0]   int_reg_array_38_26_imag;
  reg        [15:0]   int_reg_array_38_27_real;
  reg        [15:0]   int_reg_array_38_27_imag;
  reg        [15:0]   int_reg_array_38_28_real;
  reg        [15:0]   int_reg_array_38_28_imag;
  reg        [15:0]   int_reg_array_38_29_real;
  reg        [15:0]   int_reg_array_38_29_imag;
  reg        [15:0]   int_reg_array_38_30_real;
  reg        [15:0]   int_reg_array_38_30_imag;
  reg        [15:0]   int_reg_array_38_31_real;
  reg        [15:0]   int_reg_array_38_31_imag;
  reg        [15:0]   int_reg_array_38_32_real;
  reg        [15:0]   int_reg_array_38_32_imag;
  reg        [15:0]   int_reg_array_38_33_real;
  reg        [15:0]   int_reg_array_38_33_imag;
  reg        [15:0]   int_reg_array_38_34_real;
  reg        [15:0]   int_reg_array_38_34_imag;
  reg        [15:0]   int_reg_array_38_35_real;
  reg        [15:0]   int_reg_array_38_35_imag;
  reg        [15:0]   int_reg_array_38_36_real;
  reg        [15:0]   int_reg_array_38_36_imag;
  reg        [15:0]   int_reg_array_38_37_real;
  reg        [15:0]   int_reg_array_38_37_imag;
  reg        [15:0]   int_reg_array_38_38_real;
  reg        [15:0]   int_reg_array_38_38_imag;
  reg        [15:0]   int_reg_array_38_39_real;
  reg        [15:0]   int_reg_array_38_39_imag;
  reg        [15:0]   int_reg_array_38_40_real;
  reg        [15:0]   int_reg_array_38_40_imag;
  reg        [15:0]   int_reg_array_38_41_real;
  reg        [15:0]   int_reg_array_38_41_imag;
  reg        [15:0]   int_reg_array_38_42_real;
  reg        [15:0]   int_reg_array_38_42_imag;
  reg        [15:0]   int_reg_array_38_43_real;
  reg        [15:0]   int_reg_array_38_43_imag;
  reg        [15:0]   int_reg_array_38_44_real;
  reg        [15:0]   int_reg_array_38_44_imag;
  reg        [15:0]   int_reg_array_38_45_real;
  reg        [15:0]   int_reg_array_38_45_imag;
  reg        [15:0]   int_reg_array_38_46_real;
  reg        [15:0]   int_reg_array_38_46_imag;
  reg        [15:0]   int_reg_array_38_47_real;
  reg        [15:0]   int_reg_array_38_47_imag;
  reg        [15:0]   int_reg_array_38_48_real;
  reg        [15:0]   int_reg_array_38_48_imag;
  reg        [15:0]   int_reg_array_38_49_real;
  reg        [15:0]   int_reg_array_38_49_imag;
  reg        [15:0]   int_reg_array_38_50_real;
  reg        [15:0]   int_reg_array_38_50_imag;
  reg        [15:0]   int_reg_array_38_51_real;
  reg        [15:0]   int_reg_array_38_51_imag;
  reg        [15:0]   int_reg_array_38_52_real;
  reg        [15:0]   int_reg_array_38_52_imag;
  reg        [15:0]   int_reg_array_38_53_real;
  reg        [15:0]   int_reg_array_38_53_imag;
  reg        [15:0]   int_reg_array_38_54_real;
  reg        [15:0]   int_reg_array_38_54_imag;
  reg        [15:0]   int_reg_array_38_55_real;
  reg        [15:0]   int_reg_array_38_55_imag;
  reg        [15:0]   int_reg_array_38_56_real;
  reg        [15:0]   int_reg_array_38_56_imag;
  reg        [15:0]   int_reg_array_38_57_real;
  reg        [15:0]   int_reg_array_38_57_imag;
  reg        [15:0]   int_reg_array_38_58_real;
  reg        [15:0]   int_reg_array_38_58_imag;
  reg        [15:0]   int_reg_array_38_59_real;
  reg        [15:0]   int_reg_array_38_59_imag;
  reg        [15:0]   int_reg_array_38_60_real;
  reg        [15:0]   int_reg_array_38_60_imag;
  reg        [15:0]   int_reg_array_38_61_real;
  reg        [15:0]   int_reg_array_38_61_imag;
  reg        [15:0]   int_reg_array_38_62_real;
  reg        [15:0]   int_reg_array_38_62_imag;
  reg        [15:0]   int_reg_array_38_63_real;
  reg        [15:0]   int_reg_array_38_63_imag;
  reg        [15:0]   int_reg_array_41_0_real;
  reg        [15:0]   int_reg_array_41_0_imag;
  reg        [15:0]   int_reg_array_41_1_real;
  reg        [15:0]   int_reg_array_41_1_imag;
  reg        [15:0]   int_reg_array_41_2_real;
  reg        [15:0]   int_reg_array_41_2_imag;
  reg        [15:0]   int_reg_array_41_3_real;
  reg        [15:0]   int_reg_array_41_3_imag;
  reg        [15:0]   int_reg_array_41_4_real;
  reg        [15:0]   int_reg_array_41_4_imag;
  reg        [15:0]   int_reg_array_41_5_real;
  reg        [15:0]   int_reg_array_41_5_imag;
  reg        [15:0]   int_reg_array_41_6_real;
  reg        [15:0]   int_reg_array_41_6_imag;
  reg        [15:0]   int_reg_array_41_7_real;
  reg        [15:0]   int_reg_array_41_7_imag;
  reg        [15:0]   int_reg_array_41_8_real;
  reg        [15:0]   int_reg_array_41_8_imag;
  reg        [15:0]   int_reg_array_41_9_real;
  reg        [15:0]   int_reg_array_41_9_imag;
  reg        [15:0]   int_reg_array_41_10_real;
  reg        [15:0]   int_reg_array_41_10_imag;
  reg        [15:0]   int_reg_array_41_11_real;
  reg        [15:0]   int_reg_array_41_11_imag;
  reg        [15:0]   int_reg_array_41_12_real;
  reg        [15:0]   int_reg_array_41_12_imag;
  reg        [15:0]   int_reg_array_41_13_real;
  reg        [15:0]   int_reg_array_41_13_imag;
  reg        [15:0]   int_reg_array_41_14_real;
  reg        [15:0]   int_reg_array_41_14_imag;
  reg        [15:0]   int_reg_array_41_15_real;
  reg        [15:0]   int_reg_array_41_15_imag;
  reg        [15:0]   int_reg_array_41_16_real;
  reg        [15:0]   int_reg_array_41_16_imag;
  reg        [15:0]   int_reg_array_41_17_real;
  reg        [15:0]   int_reg_array_41_17_imag;
  reg        [15:0]   int_reg_array_41_18_real;
  reg        [15:0]   int_reg_array_41_18_imag;
  reg        [15:0]   int_reg_array_41_19_real;
  reg        [15:0]   int_reg_array_41_19_imag;
  reg        [15:0]   int_reg_array_41_20_real;
  reg        [15:0]   int_reg_array_41_20_imag;
  reg        [15:0]   int_reg_array_41_21_real;
  reg        [15:0]   int_reg_array_41_21_imag;
  reg        [15:0]   int_reg_array_41_22_real;
  reg        [15:0]   int_reg_array_41_22_imag;
  reg        [15:0]   int_reg_array_41_23_real;
  reg        [15:0]   int_reg_array_41_23_imag;
  reg        [15:0]   int_reg_array_41_24_real;
  reg        [15:0]   int_reg_array_41_24_imag;
  reg        [15:0]   int_reg_array_41_25_real;
  reg        [15:0]   int_reg_array_41_25_imag;
  reg        [15:0]   int_reg_array_41_26_real;
  reg        [15:0]   int_reg_array_41_26_imag;
  reg        [15:0]   int_reg_array_41_27_real;
  reg        [15:0]   int_reg_array_41_27_imag;
  reg        [15:0]   int_reg_array_41_28_real;
  reg        [15:0]   int_reg_array_41_28_imag;
  reg        [15:0]   int_reg_array_41_29_real;
  reg        [15:0]   int_reg_array_41_29_imag;
  reg        [15:0]   int_reg_array_41_30_real;
  reg        [15:0]   int_reg_array_41_30_imag;
  reg        [15:0]   int_reg_array_41_31_real;
  reg        [15:0]   int_reg_array_41_31_imag;
  reg        [15:0]   int_reg_array_41_32_real;
  reg        [15:0]   int_reg_array_41_32_imag;
  reg        [15:0]   int_reg_array_41_33_real;
  reg        [15:0]   int_reg_array_41_33_imag;
  reg        [15:0]   int_reg_array_41_34_real;
  reg        [15:0]   int_reg_array_41_34_imag;
  reg        [15:0]   int_reg_array_41_35_real;
  reg        [15:0]   int_reg_array_41_35_imag;
  reg        [15:0]   int_reg_array_41_36_real;
  reg        [15:0]   int_reg_array_41_36_imag;
  reg        [15:0]   int_reg_array_41_37_real;
  reg        [15:0]   int_reg_array_41_37_imag;
  reg        [15:0]   int_reg_array_41_38_real;
  reg        [15:0]   int_reg_array_41_38_imag;
  reg        [15:0]   int_reg_array_41_39_real;
  reg        [15:0]   int_reg_array_41_39_imag;
  reg        [15:0]   int_reg_array_41_40_real;
  reg        [15:0]   int_reg_array_41_40_imag;
  reg        [15:0]   int_reg_array_41_41_real;
  reg        [15:0]   int_reg_array_41_41_imag;
  reg        [15:0]   int_reg_array_41_42_real;
  reg        [15:0]   int_reg_array_41_42_imag;
  reg        [15:0]   int_reg_array_41_43_real;
  reg        [15:0]   int_reg_array_41_43_imag;
  reg        [15:0]   int_reg_array_41_44_real;
  reg        [15:0]   int_reg_array_41_44_imag;
  reg        [15:0]   int_reg_array_41_45_real;
  reg        [15:0]   int_reg_array_41_45_imag;
  reg        [15:0]   int_reg_array_41_46_real;
  reg        [15:0]   int_reg_array_41_46_imag;
  reg        [15:0]   int_reg_array_41_47_real;
  reg        [15:0]   int_reg_array_41_47_imag;
  reg        [15:0]   int_reg_array_41_48_real;
  reg        [15:0]   int_reg_array_41_48_imag;
  reg        [15:0]   int_reg_array_41_49_real;
  reg        [15:0]   int_reg_array_41_49_imag;
  reg        [15:0]   int_reg_array_41_50_real;
  reg        [15:0]   int_reg_array_41_50_imag;
  reg        [15:0]   int_reg_array_41_51_real;
  reg        [15:0]   int_reg_array_41_51_imag;
  reg        [15:0]   int_reg_array_41_52_real;
  reg        [15:0]   int_reg_array_41_52_imag;
  reg        [15:0]   int_reg_array_41_53_real;
  reg        [15:0]   int_reg_array_41_53_imag;
  reg        [15:0]   int_reg_array_41_54_real;
  reg        [15:0]   int_reg_array_41_54_imag;
  reg        [15:0]   int_reg_array_41_55_real;
  reg        [15:0]   int_reg_array_41_55_imag;
  reg        [15:0]   int_reg_array_41_56_real;
  reg        [15:0]   int_reg_array_41_56_imag;
  reg        [15:0]   int_reg_array_41_57_real;
  reg        [15:0]   int_reg_array_41_57_imag;
  reg        [15:0]   int_reg_array_41_58_real;
  reg        [15:0]   int_reg_array_41_58_imag;
  reg        [15:0]   int_reg_array_41_59_real;
  reg        [15:0]   int_reg_array_41_59_imag;
  reg        [15:0]   int_reg_array_41_60_real;
  reg        [15:0]   int_reg_array_41_60_imag;
  reg        [15:0]   int_reg_array_41_61_real;
  reg        [15:0]   int_reg_array_41_61_imag;
  reg        [15:0]   int_reg_array_41_62_real;
  reg        [15:0]   int_reg_array_41_62_imag;
  reg        [15:0]   int_reg_array_41_63_real;
  reg        [15:0]   int_reg_array_41_63_imag;
  reg        [15:0]   int_reg_array_49_0_real;
  reg        [15:0]   int_reg_array_49_0_imag;
  reg        [15:0]   int_reg_array_49_1_real;
  reg        [15:0]   int_reg_array_49_1_imag;
  reg        [15:0]   int_reg_array_49_2_real;
  reg        [15:0]   int_reg_array_49_2_imag;
  reg        [15:0]   int_reg_array_49_3_real;
  reg        [15:0]   int_reg_array_49_3_imag;
  reg        [15:0]   int_reg_array_49_4_real;
  reg        [15:0]   int_reg_array_49_4_imag;
  reg        [15:0]   int_reg_array_49_5_real;
  reg        [15:0]   int_reg_array_49_5_imag;
  reg        [15:0]   int_reg_array_49_6_real;
  reg        [15:0]   int_reg_array_49_6_imag;
  reg        [15:0]   int_reg_array_49_7_real;
  reg        [15:0]   int_reg_array_49_7_imag;
  reg        [15:0]   int_reg_array_49_8_real;
  reg        [15:0]   int_reg_array_49_8_imag;
  reg        [15:0]   int_reg_array_49_9_real;
  reg        [15:0]   int_reg_array_49_9_imag;
  reg        [15:0]   int_reg_array_49_10_real;
  reg        [15:0]   int_reg_array_49_10_imag;
  reg        [15:0]   int_reg_array_49_11_real;
  reg        [15:0]   int_reg_array_49_11_imag;
  reg        [15:0]   int_reg_array_49_12_real;
  reg        [15:0]   int_reg_array_49_12_imag;
  reg        [15:0]   int_reg_array_49_13_real;
  reg        [15:0]   int_reg_array_49_13_imag;
  reg        [15:0]   int_reg_array_49_14_real;
  reg        [15:0]   int_reg_array_49_14_imag;
  reg        [15:0]   int_reg_array_49_15_real;
  reg        [15:0]   int_reg_array_49_15_imag;
  reg        [15:0]   int_reg_array_49_16_real;
  reg        [15:0]   int_reg_array_49_16_imag;
  reg        [15:0]   int_reg_array_49_17_real;
  reg        [15:0]   int_reg_array_49_17_imag;
  reg        [15:0]   int_reg_array_49_18_real;
  reg        [15:0]   int_reg_array_49_18_imag;
  reg        [15:0]   int_reg_array_49_19_real;
  reg        [15:0]   int_reg_array_49_19_imag;
  reg        [15:0]   int_reg_array_49_20_real;
  reg        [15:0]   int_reg_array_49_20_imag;
  reg        [15:0]   int_reg_array_49_21_real;
  reg        [15:0]   int_reg_array_49_21_imag;
  reg        [15:0]   int_reg_array_49_22_real;
  reg        [15:0]   int_reg_array_49_22_imag;
  reg        [15:0]   int_reg_array_49_23_real;
  reg        [15:0]   int_reg_array_49_23_imag;
  reg        [15:0]   int_reg_array_49_24_real;
  reg        [15:0]   int_reg_array_49_24_imag;
  reg        [15:0]   int_reg_array_49_25_real;
  reg        [15:0]   int_reg_array_49_25_imag;
  reg        [15:0]   int_reg_array_49_26_real;
  reg        [15:0]   int_reg_array_49_26_imag;
  reg        [15:0]   int_reg_array_49_27_real;
  reg        [15:0]   int_reg_array_49_27_imag;
  reg        [15:0]   int_reg_array_49_28_real;
  reg        [15:0]   int_reg_array_49_28_imag;
  reg        [15:0]   int_reg_array_49_29_real;
  reg        [15:0]   int_reg_array_49_29_imag;
  reg        [15:0]   int_reg_array_49_30_real;
  reg        [15:0]   int_reg_array_49_30_imag;
  reg        [15:0]   int_reg_array_49_31_real;
  reg        [15:0]   int_reg_array_49_31_imag;
  reg        [15:0]   int_reg_array_49_32_real;
  reg        [15:0]   int_reg_array_49_32_imag;
  reg        [15:0]   int_reg_array_49_33_real;
  reg        [15:0]   int_reg_array_49_33_imag;
  reg        [15:0]   int_reg_array_49_34_real;
  reg        [15:0]   int_reg_array_49_34_imag;
  reg        [15:0]   int_reg_array_49_35_real;
  reg        [15:0]   int_reg_array_49_35_imag;
  reg        [15:0]   int_reg_array_49_36_real;
  reg        [15:0]   int_reg_array_49_36_imag;
  reg        [15:0]   int_reg_array_49_37_real;
  reg        [15:0]   int_reg_array_49_37_imag;
  reg        [15:0]   int_reg_array_49_38_real;
  reg        [15:0]   int_reg_array_49_38_imag;
  reg        [15:0]   int_reg_array_49_39_real;
  reg        [15:0]   int_reg_array_49_39_imag;
  reg        [15:0]   int_reg_array_49_40_real;
  reg        [15:0]   int_reg_array_49_40_imag;
  reg        [15:0]   int_reg_array_49_41_real;
  reg        [15:0]   int_reg_array_49_41_imag;
  reg        [15:0]   int_reg_array_49_42_real;
  reg        [15:0]   int_reg_array_49_42_imag;
  reg        [15:0]   int_reg_array_49_43_real;
  reg        [15:0]   int_reg_array_49_43_imag;
  reg        [15:0]   int_reg_array_49_44_real;
  reg        [15:0]   int_reg_array_49_44_imag;
  reg        [15:0]   int_reg_array_49_45_real;
  reg        [15:0]   int_reg_array_49_45_imag;
  reg        [15:0]   int_reg_array_49_46_real;
  reg        [15:0]   int_reg_array_49_46_imag;
  reg        [15:0]   int_reg_array_49_47_real;
  reg        [15:0]   int_reg_array_49_47_imag;
  reg        [15:0]   int_reg_array_49_48_real;
  reg        [15:0]   int_reg_array_49_48_imag;
  reg        [15:0]   int_reg_array_49_49_real;
  reg        [15:0]   int_reg_array_49_49_imag;
  reg        [15:0]   int_reg_array_49_50_real;
  reg        [15:0]   int_reg_array_49_50_imag;
  reg        [15:0]   int_reg_array_49_51_real;
  reg        [15:0]   int_reg_array_49_51_imag;
  reg        [15:0]   int_reg_array_49_52_real;
  reg        [15:0]   int_reg_array_49_52_imag;
  reg        [15:0]   int_reg_array_49_53_real;
  reg        [15:0]   int_reg_array_49_53_imag;
  reg        [15:0]   int_reg_array_49_54_real;
  reg        [15:0]   int_reg_array_49_54_imag;
  reg        [15:0]   int_reg_array_49_55_real;
  reg        [15:0]   int_reg_array_49_55_imag;
  reg        [15:0]   int_reg_array_49_56_real;
  reg        [15:0]   int_reg_array_49_56_imag;
  reg        [15:0]   int_reg_array_49_57_real;
  reg        [15:0]   int_reg_array_49_57_imag;
  reg        [15:0]   int_reg_array_49_58_real;
  reg        [15:0]   int_reg_array_49_58_imag;
  reg        [15:0]   int_reg_array_49_59_real;
  reg        [15:0]   int_reg_array_49_59_imag;
  reg        [15:0]   int_reg_array_49_60_real;
  reg        [15:0]   int_reg_array_49_60_imag;
  reg        [15:0]   int_reg_array_49_61_real;
  reg        [15:0]   int_reg_array_49_61_imag;
  reg        [15:0]   int_reg_array_49_62_real;
  reg        [15:0]   int_reg_array_49_62_imag;
  reg        [15:0]   int_reg_array_49_63_real;
  reg        [15:0]   int_reg_array_49_63_imag;
  reg        [15:0]   int_reg_array_40_0_real;
  reg        [15:0]   int_reg_array_40_0_imag;
  reg        [15:0]   int_reg_array_40_1_real;
  reg        [15:0]   int_reg_array_40_1_imag;
  reg        [15:0]   int_reg_array_40_2_real;
  reg        [15:0]   int_reg_array_40_2_imag;
  reg        [15:0]   int_reg_array_40_3_real;
  reg        [15:0]   int_reg_array_40_3_imag;
  reg        [15:0]   int_reg_array_40_4_real;
  reg        [15:0]   int_reg_array_40_4_imag;
  reg        [15:0]   int_reg_array_40_5_real;
  reg        [15:0]   int_reg_array_40_5_imag;
  reg        [15:0]   int_reg_array_40_6_real;
  reg        [15:0]   int_reg_array_40_6_imag;
  reg        [15:0]   int_reg_array_40_7_real;
  reg        [15:0]   int_reg_array_40_7_imag;
  reg        [15:0]   int_reg_array_40_8_real;
  reg        [15:0]   int_reg_array_40_8_imag;
  reg        [15:0]   int_reg_array_40_9_real;
  reg        [15:0]   int_reg_array_40_9_imag;
  reg        [15:0]   int_reg_array_40_10_real;
  reg        [15:0]   int_reg_array_40_10_imag;
  reg        [15:0]   int_reg_array_40_11_real;
  reg        [15:0]   int_reg_array_40_11_imag;
  reg        [15:0]   int_reg_array_40_12_real;
  reg        [15:0]   int_reg_array_40_12_imag;
  reg        [15:0]   int_reg_array_40_13_real;
  reg        [15:0]   int_reg_array_40_13_imag;
  reg        [15:0]   int_reg_array_40_14_real;
  reg        [15:0]   int_reg_array_40_14_imag;
  reg        [15:0]   int_reg_array_40_15_real;
  reg        [15:0]   int_reg_array_40_15_imag;
  reg        [15:0]   int_reg_array_40_16_real;
  reg        [15:0]   int_reg_array_40_16_imag;
  reg        [15:0]   int_reg_array_40_17_real;
  reg        [15:0]   int_reg_array_40_17_imag;
  reg        [15:0]   int_reg_array_40_18_real;
  reg        [15:0]   int_reg_array_40_18_imag;
  reg        [15:0]   int_reg_array_40_19_real;
  reg        [15:0]   int_reg_array_40_19_imag;
  reg        [15:0]   int_reg_array_40_20_real;
  reg        [15:0]   int_reg_array_40_20_imag;
  reg        [15:0]   int_reg_array_40_21_real;
  reg        [15:0]   int_reg_array_40_21_imag;
  reg        [15:0]   int_reg_array_40_22_real;
  reg        [15:0]   int_reg_array_40_22_imag;
  reg        [15:0]   int_reg_array_40_23_real;
  reg        [15:0]   int_reg_array_40_23_imag;
  reg        [15:0]   int_reg_array_40_24_real;
  reg        [15:0]   int_reg_array_40_24_imag;
  reg        [15:0]   int_reg_array_40_25_real;
  reg        [15:0]   int_reg_array_40_25_imag;
  reg        [15:0]   int_reg_array_40_26_real;
  reg        [15:0]   int_reg_array_40_26_imag;
  reg        [15:0]   int_reg_array_40_27_real;
  reg        [15:0]   int_reg_array_40_27_imag;
  reg        [15:0]   int_reg_array_40_28_real;
  reg        [15:0]   int_reg_array_40_28_imag;
  reg        [15:0]   int_reg_array_40_29_real;
  reg        [15:0]   int_reg_array_40_29_imag;
  reg        [15:0]   int_reg_array_40_30_real;
  reg        [15:0]   int_reg_array_40_30_imag;
  reg        [15:0]   int_reg_array_40_31_real;
  reg        [15:0]   int_reg_array_40_31_imag;
  reg        [15:0]   int_reg_array_40_32_real;
  reg        [15:0]   int_reg_array_40_32_imag;
  reg        [15:0]   int_reg_array_40_33_real;
  reg        [15:0]   int_reg_array_40_33_imag;
  reg        [15:0]   int_reg_array_40_34_real;
  reg        [15:0]   int_reg_array_40_34_imag;
  reg        [15:0]   int_reg_array_40_35_real;
  reg        [15:0]   int_reg_array_40_35_imag;
  reg        [15:0]   int_reg_array_40_36_real;
  reg        [15:0]   int_reg_array_40_36_imag;
  reg        [15:0]   int_reg_array_40_37_real;
  reg        [15:0]   int_reg_array_40_37_imag;
  reg        [15:0]   int_reg_array_40_38_real;
  reg        [15:0]   int_reg_array_40_38_imag;
  reg        [15:0]   int_reg_array_40_39_real;
  reg        [15:0]   int_reg_array_40_39_imag;
  reg        [15:0]   int_reg_array_40_40_real;
  reg        [15:0]   int_reg_array_40_40_imag;
  reg        [15:0]   int_reg_array_40_41_real;
  reg        [15:0]   int_reg_array_40_41_imag;
  reg        [15:0]   int_reg_array_40_42_real;
  reg        [15:0]   int_reg_array_40_42_imag;
  reg        [15:0]   int_reg_array_40_43_real;
  reg        [15:0]   int_reg_array_40_43_imag;
  reg        [15:0]   int_reg_array_40_44_real;
  reg        [15:0]   int_reg_array_40_44_imag;
  reg        [15:0]   int_reg_array_40_45_real;
  reg        [15:0]   int_reg_array_40_45_imag;
  reg        [15:0]   int_reg_array_40_46_real;
  reg        [15:0]   int_reg_array_40_46_imag;
  reg        [15:0]   int_reg_array_40_47_real;
  reg        [15:0]   int_reg_array_40_47_imag;
  reg        [15:0]   int_reg_array_40_48_real;
  reg        [15:0]   int_reg_array_40_48_imag;
  reg        [15:0]   int_reg_array_40_49_real;
  reg        [15:0]   int_reg_array_40_49_imag;
  reg        [15:0]   int_reg_array_40_50_real;
  reg        [15:0]   int_reg_array_40_50_imag;
  reg        [15:0]   int_reg_array_40_51_real;
  reg        [15:0]   int_reg_array_40_51_imag;
  reg        [15:0]   int_reg_array_40_52_real;
  reg        [15:0]   int_reg_array_40_52_imag;
  reg        [15:0]   int_reg_array_40_53_real;
  reg        [15:0]   int_reg_array_40_53_imag;
  reg        [15:0]   int_reg_array_40_54_real;
  reg        [15:0]   int_reg_array_40_54_imag;
  reg        [15:0]   int_reg_array_40_55_real;
  reg        [15:0]   int_reg_array_40_55_imag;
  reg        [15:0]   int_reg_array_40_56_real;
  reg        [15:0]   int_reg_array_40_56_imag;
  reg        [15:0]   int_reg_array_40_57_real;
  reg        [15:0]   int_reg_array_40_57_imag;
  reg        [15:0]   int_reg_array_40_58_real;
  reg        [15:0]   int_reg_array_40_58_imag;
  reg        [15:0]   int_reg_array_40_59_real;
  reg        [15:0]   int_reg_array_40_59_imag;
  reg        [15:0]   int_reg_array_40_60_real;
  reg        [15:0]   int_reg_array_40_60_imag;
  reg        [15:0]   int_reg_array_40_61_real;
  reg        [15:0]   int_reg_array_40_61_imag;
  reg        [15:0]   int_reg_array_40_62_real;
  reg        [15:0]   int_reg_array_40_62_imag;
  reg        [15:0]   int_reg_array_40_63_real;
  reg        [15:0]   int_reg_array_40_63_imag;
  reg        [15:0]   int_reg_array_14_0_real;
  reg        [15:0]   int_reg_array_14_0_imag;
  reg        [15:0]   int_reg_array_14_1_real;
  reg        [15:0]   int_reg_array_14_1_imag;
  reg        [15:0]   int_reg_array_14_2_real;
  reg        [15:0]   int_reg_array_14_2_imag;
  reg        [15:0]   int_reg_array_14_3_real;
  reg        [15:0]   int_reg_array_14_3_imag;
  reg        [15:0]   int_reg_array_14_4_real;
  reg        [15:0]   int_reg_array_14_4_imag;
  reg        [15:0]   int_reg_array_14_5_real;
  reg        [15:0]   int_reg_array_14_5_imag;
  reg        [15:0]   int_reg_array_14_6_real;
  reg        [15:0]   int_reg_array_14_6_imag;
  reg        [15:0]   int_reg_array_14_7_real;
  reg        [15:0]   int_reg_array_14_7_imag;
  reg        [15:0]   int_reg_array_14_8_real;
  reg        [15:0]   int_reg_array_14_8_imag;
  reg        [15:0]   int_reg_array_14_9_real;
  reg        [15:0]   int_reg_array_14_9_imag;
  reg        [15:0]   int_reg_array_14_10_real;
  reg        [15:0]   int_reg_array_14_10_imag;
  reg        [15:0]   int_reg_array_14_11_real;
  reg        [15:0]   int_reg_array_14_11_imag;
  reg        [15:0]   int_reg_array_14_12_real;
  reg        [15:0]   int_reg_array_14_12_imag;
  reg        [15:0]   int_reg_array_14_13_real;
  reg        [15:0]   int_reg_array_14_13_imag;
  reg        [15:0]   int_reg_array_14_14_real;
  reg        [15:0]   int_reg_array_14_14_imag;
  reg        [15:0]   int_reg_array_14_15_real;
  reg        [15:0]   int_reg_array_14_15_imag;
  reg        [15:0]   int_reg_array_14_16_real;
  reg        [15:0]   int_reg_array_14_16_imag;
  reg        [15:0]   int_reg_array_14_17_real;
  reg        [15:0]   int_reg_array_14_17_imag;
  reg        [15:0]   int_reg_array_14_18_real;
  reg        [15:0]   int_reg_array_14_18_imag;
  reg        [15:0]   int_reg_array_14_19_real;
  reg        [15:0]   int_reg_array_14_19_imag;
  reg        [15:0]   int_reg_array_14_20_real;
  reg        [15:0]   int_reg_array_14_20_imag;
  reg        [15:0]   int_reg_array_14_21_real;
  reg        [15:0]   int_reg_array_14_21_imag;
  reg        [15:0]   int_reg_array_14_22_real;
  reg        [15:0]   int_reg_array_14_22_imag;
  reg        [15:0]   int_reg_array_14_23_real;
  reg        [15:0]   int_reg_array_14_23_imag;
  reg        [15:0]   int_reg_array_14_24_real;
  reg        [15:0]   int_reg_array_14_24_imag;
  reg        [15:0]   int_reg_array_14_25_real;
  reg        [15:0]   int_reg_array_14_25_imag;
  reg        [15:0]   int_reg_array_14_26_real;
  reg        [15:0]   int_reg_array_14_26_imag;
  reg        [15:0]   int_reg_array_14_27_real;
  reg        [15:0]   int_reg_array_14_27_imag;
  reg        [15:0]   int_reg_array_14_28_real;
  reg        [15:0]   int_reg_array_14_28_imag;
  reg        [15:0]   int_reg_array_14_29_real;
  reg        [15:0]   int_reg_array_14_29_imag;
  reg        [15:0]   int_reg_array_14_30_real;
  reg        [15:0]   int_reg_array_14_30_imag;
  reg        [15:0]   int_reg_array_14_31_real;
  reg        [15:0]   int_reg_array_14_31_imag;
  reg        [15:0]   int_reg_array_14_32_real;
  reg        [15:0]   int_reg_array_14_32_imag;
  reg        [15:0]   int_reg_array_14_33_real;
  reg        [15:0]   int_reg_array_14_33_imag;
  reg        [15:0]   int_reg_array_14_34_real;
  reg        [15:0]   int_reg_array_14_34_imag;
  reg        [15:0]   int_reg_array_14_35_real;
  reg        [15:0]   int_reg_array_14_35_imag;
  reg        [15:0]   int_reg_array_14_36_real;
  reg        [15:0]   int_reg_array_14_36_imag;
  reg        [15:0]   int_reg_array_14_37_real;
  reg        [15:0]   int_reg_array_14_37_imag;
  reg        [15:0]   int_reg_array_14_38_real;
  reg        [15:0]   int_reg_array_14_38_imag;
  reg        [15:0]   int_reg_array_14_39_real;
  reg        [15:0]   int_reg_array_14_39_imag;
  reg        [15:0]   int_reg_array_14_40_real;
  reg        [15:0]   int_reg_array_14_40_imag;
  reg        [15:0]   int_reg_array_14_41_real;
  reg        [15:0]   int_reg_array_14_41_imag;
  reg        [15:0]   int_reg_array_14_42_real;
  reg        [15:0]   int_reg_array_14_42_imag;
  reg        [15:0]   int_reg_array_14_43_real;
  reg        [15:0]   int_reg_array_14_43_imag;
  reg        [15:0]   int_reg_array_14_44_real;
  reg        [15:0]   int_reg_array_14_44_imag;
  reg        [15:0]   int_reg_array_14_45_real;
  reg        [15:0]   int_reg_array_14_45_imag;
  reg        [15:0]   int_reg_array_14_46_real;
  reg        [15:0]   int_reg_array_14_46_imag;
  reg        [15:0]   int_reg_array_14_47_real;
  reg        [15:0]   int_reg_array_14_47_imag;
  reg        [15:0]   int_reg_array_14_48_real;
  reg        [15:0]   int_reg_array_14_48_imag;
  reg        [15:0]   int_reg_array_14_49_real;
  reg        [15:0]   int_reg_array_14_49_imag;
  reg        [15:0]   int_reg_array_14_50_real;
  reg        [15:0]   int_reg_array_14_50_imag;
  reg        [15:0]   int_reg_array_14_51_real;
  reg        [15:0]   int_reg_array_14_51_imag;
  reg        [15:0]   int_reg_array_14_52_real;
  reg        [15:0]   int_reg_array_14_52_imag;
  reg        [15:0]   int_reg_array_14_53_real;
  reg        [15:0]   int_reg_array_14_53_imag;
  reg        [15:0]   int_reg_array_14_54_real;
  reg        [15:0]   int_reg_array_14_54_imag;
  reg        [15:0]   int_reg_array_14_55_real;
  reg        [15:0]   int_reg_array_14_55_imag;
  reg        [15:0]   int_reg_array_14_56_real;
  reg        [15:0]   int_reg_array_14_56_imag;
  reg        [15:0]   int_reg_array_14_57_real;
  reg        [15:0]   int_reg_array_14_57_imag;
  reg        [15:0]   int_reg_array_14_58_real;
  reg        [15:0]   int_reg_array_14_58_imag;
  reg        [15:0]   int_reg_array_14_59_real;
  reg        [15:0]   int_reg_array_14_59_imag;
  reg        [15:0]   int_reg_array_14_60_real;
  reg        [15:0]   int_reg_array_14_60_imag;
  reg        [15:0]   int_reg_array_14_61_real;
  reg        [15:0]   int_reg_array_14_61_imag;
  reg        [15:0]   int_reg_array_14_62_real;
  reg        [15:0]   int_reg_array_14_62_imag;
  reg        [15:0]   int_reg_array_14_63_real;
  reg        [15:0]   int_reg_array_14_63_imag;
  reg        [15:0]   int_reg_array_19_0_real;
  reg        [15:0]   int_reg_array_19_0_imag;
  reg        [15:0]   int_reg_array_19_1_real;
  reg        [15:0]   int_reg_array_19_1_imag;
  reg        [15:0]   int_reg_array_19_2_real;
  reg        [15:0]   int_reg_array_19_2_imag;
  reg        [15:0]   int_reg_array_19_3_real;
  reg        [15:0]   int_reg_array_19_3_imag;
  reg        [15:0]   int_reg_array_19_4_real;
  reg        [15:0]   int_reg_array_19_4_imag;
  reg        [15:0]   int_reg_array_19_5_real;
  reg        [15:0]   int_reg_array_19_5_imag;
  reg        [15:0]   int_reg_array_19_6_real;
  reg        [15:0]   int_reg_array_19_6_imag;
  reg        [15:0]   int_reg_array_19_7_real;
  reg        [15:0]   int_reg_array_19_7_imag;
  reg        [15:0]   int_reg_array_19_8_real;
  reg        [15:0]   int_reg_array_19_8_imag;
  reg        [15:0]   int_reg_array_19_9_real;
  reg        [15:0]   int_reg_array_19_9_imag;
  reg        [15:0]   int_reg_array_19_10_real;
  reg        [15:0]   int_reg_array_19_10_imag;
  reg        [15:0]   int_reg_array_19_11_real;
  reg        [15:0]   int_reg_array_19_11_imag;
  reg        [15:0]   int_reg_array_19_12_real;
  reg        [15:0]   int_reg_array_19_12_imag;
  reg        [15:0]   int_reg_array_19_13_real;
  reg        [15:0]   int_reg_array_19_13_imag;
  reg        [15:0]   int_reg_array_19_14_real;
  reg        [15:0]   int_reg_array_19_14_imag;
  reg        [15:0]   int_reg_array_19_15_real;
  reg        [15:0]   int_reg_array_19_15_imag;
  reg        [15:0]   int_reg_array_19_16_real;
  reg        [15:0]   int_reg_array_19_16_imag;
  reg        [15:0]   int_reg_array_19_17_real;
  reg        [15:0]   int_reg_array_19_17_imag;
  reg        [15:0]   int_reg_array_19_18_real;
  reg        [15:0]   int_reg_array_19_18_imag;
  reg        [15:0]   int_reg_array_19_19_real;
  reg        [15:0]   int_reg_array_19_19_imag;
  reg        [15:0]   int_reg_array_19_20_real;
  reg        [15:0]   int_reg_array_19_20_imag;
  reg        [15:0]   int_reg_array_19_21_real;
  reg        [15:0]   int_reg_array_19_21_imag;
  reg        [15:0]   int_reg_array_19_22_real;
  reg        [15:0]   int_reg_array_19_22_imag;
  reg        [15:0]   int_reg_array_19_23_real;
  reg        [15:0]   int_reg_array_19_23_imag;
  reg        [15:0]   int_reg_array_19_24_real;
  reg        [15:0]   int_reg_array_19_24_imag;
  reg        [15:0]   int_reg_array_19_25_real;
  reg        [15:0]   int_reg_array_19_25_imag;
  reg        [15:0]   int_reg_array_19_26_real;
  reg        [15:0]   int_reg_array_19_26_imag;
  reg        [15:0]   int_reg_array_19_27_real;
  reg        [15:0]   int_reg_array_19_27_imag;
  reg        [15:0]   int_reg_array_19_28_real;
  reg        [15:0]   int_reg_array_19_28_imag;
  reg        [15:0]   int_reg_array_19_29_real;
  reg        [15:0]   int_reg_array_19_29_imag;
  reg        [15:0]   int_reg_array_19_30_real;
  reg        [15:0]   int_reg_array_19_30_imag;
  reg        [15:0]   int_reg_array_19_31_real;
  reg        [15:0]   int_reg_array_19_31_imag;
  reg        [15:0]   int_reg_array_19_32_real;
  reg        [15:0]   int_reg_array_19_32_imag;
  reg        [15:0]   int_reg_array_19_33_real;
  reg        [15:0]   int_reg_array_19_33_imag;
  reg        [15:0]   int_reg_array_19_34_real;
  reg        [15:0]   int_reg_array_19_34_imag;
  reg        [15:0]   int_reg_array_19_35_real;
  reg        [15:0]   int_reg_array_19_35_imag;
  reg        [15:0]   int_reg_array_19_36_real;
  reg        [15:0]   int_reg_array_19_36_imag;
  reg        [15:0]   int_reg_array_19_37_real;
  reg        [15:0]   int_reg_array_19_37_imag;
  reg        [15:0]   int_reg_array_19_38_real;
  reg        [15:0]   int_reg_array_19_38_imag;
  reg        [15:0]   int_reg_array_19_39_real;
  reg        [15:0]   int_reg_array_19_39_imag;
  reg        [15:0]   int_reg_array_19_40_real;
  reg        [15:0]   int_reg_array_19_40_imag;
  reg        [15:0]   int_reg_array_19_41_real;
  reg        [15:0]   int_reg_array_19_41_imag;
  reg        [15:0]   int_reg_array_19_42_real;
  reg        [15:0]   int_reg_array_19_42_imag;
  reg        [15:0]   int_reg_array_19_43_real;
  reg        [15:0]   int_reg_array_19_43_imag;
  reg        [15:0]   int_reg_array_19_44_real;
  reg        [15:0]   int_reg_array_19_44_imag;
  reg        [15:0]   int_reg_array_19_45_real;
  reg        [15:0]   int_reg_array_19_45_imag;
  reg        [15:0]   int_reg_array_19_46_real;
  reg        [15:0]   int_reg_array_19_46_imag;
  reg        [15:0]   int_reg_array_19_47_real;
  reg        [15:0]   int_reg_array_19_47_imag;
  reg        [15:0]   int_reg_array_19_48_real;
  reg        [15:0]   int_reg_array_19_48_imag;
  reg        [15:0]   int_reg_array_19_49_real;
  reg        [15:0]   int_reg_array_19_49_imag;
  reg        [15:0]   int_reg_array_19_50_real;
  reg        [15:0]   int_reg_array_19_50_imag;
  reg        [15:0]   int_reg_array_19_51_real;
  reg        [15:0]   int_reg_array_19_51_imag;
  reg        [15:0]   int_reg_array_19_52_real;
  reg        [15:0]   int_reg_array_19_52_imag;
  reg        [15:0]   int_reg_array_19_53_real;
  reg        [15:0]   int_reg_array_19_53_imag;
  reg        [15:0]   int_reg_array_19_54_real;
  reg        [15:0]   int_reg_array_19_54_imag;
  reg        [15:0]   int_reg_array_19_55_real;
  reg        [15:0]   int_reg_array_19_55_imag;
  reg        [15:0]   int_reg_array_19_56_real;
  reg        [15:0]   int_reg_array_19_56_imag;
  reg        [15:0]   int_reg_array_19_57_real;
  reg        [15:0]   int_reg_array_19_57_imag;
  reg        [15:0]   int_reg_array_19_58_real;
  reg        [15:0]   int_reg_array_19_58_imag;
  reg        [15:0]   int_reg_array_19_59_real;
  reg        [15:0]   int_reg_array_19_59_imag;
  reg        [15:0]   int_reg_array_19_60_real;
  reg        [15:0]   int_reg_array_19_60_imag;
  reg        [15:0]   int_reg_array_19_61_real;
  reg        [15:0]   int_reg_array_19_61_imag;
  reg        [15:0]   int_reg_array_19_62_real;
  reg        [15:0]   int_reg_array_19_62_imag;
  reg        [15:0]   int_reg_array_19_63_real;
  reg        [15:0]   int_reg_array_19_63_imag;
  reg        [15:0]   int_reg_array_15_0_real;
  reg        [15:0]   int_reg_array_15_0_imag;
  reg        [15:0]   int_reg_array_15_1_real;
  reg        [15:0]   int_reg_array_15_1_imag;
  reg        [15:0]   int_reg_array_15_2_real;
  reg        [15:0]   int_reg_array_15_2_imag;
  reg        [15:0]   int_reg_array_15_3_real;
  reg        [15:0]   int_reg_array_15_3_imag;
  reg        [15:0]   int_reg_array_15_4_real;
  reg        [15:0]   int_reg_array_15_4_imag;
  reg        [15:0]   int_reg_array_15_5_real;
  reg        [15:0]   int_reg_array_15_5_imag;
  reg        [15:0]   int_reg_array_15_6_real;
  reg        [15:0]   int_reg_array_15_6_imag;
  reg        [15:0]   int_reg_array_15_7_real;
  reg        [15:0]   int_reg_array_15_7_imag;
  reg        [15:0]   int_reg_array_15_8_real;
  reg        [15:0]   int_reg_array_15_8_imag;
  reg        [15:0]   int_reg_array_15_9_real;
  reg        [15:0]   int_reg_array_15_9_imag;
  reg        [15:0]   int_reg_array_15_10_real;
  reg        [15:0]   int_reg_array_15_10_imag;
  reg        [15:0]   int_reg_array_15_11_real;
  reg        [15:0]   int_reg_array_15_11_imag;
  reg        [15:0]   int_reg_array_15_12_real;
  reg        [15:0]   int_reg_array_15_12_imag;
  reg        [15:0]   int_reg_array_15_13_real;
  reg        [15:0]   int_reg_array_15_13_imag;
  reg        [15:0]   int_reg_array_15_14_real;
  reg        [15:0]   int_reg_array_15_14_imag;
  reg        [15:0]   int_reg_array_15_15_real;
  reg        [15:0]   int_reg_array_15_15_imag;
  reg        [15:0]   int_reg_array_15_16_real;
  reg        [15:0]   int_reg_array_15_16_imag;
  reg        [15:0]   int_reg_array_15_17_real;
  reg        [15:0]   int_reg_array_15_17_imag;
  reg        [15:0]   int_reg_array_15_18_real;
  reg        [15:0]   int_reg_array_15_18_imag;
  reg        [15:0]   int_reg_array_15_19_real;
  reg        [15:0]   int_reg_array_15_19_imag;
  reg        [15:0]   int_reg_array_15_20_real;
  reg        [15:0]   int_reg_array_15_20_imag;
  reg        [15:0]   int_reg_array_15_21_real;
  reg        [15:0]   int_reg_array_15_21_imag;
  reg        [15:0]   int_reg_array_15_22_real;
  reg        [15:0]   int_reg_array_15_22_imag;
  reg        [15:0]   int_reg_array_15_23_real;
  reg        [15:0]   int_reg_array_15_23_imag;
  reg        [15:0]   int_reg_array_15_24_real;
  reg        [15:0]   int_reg_array_15_24_imag;
  reg        [15:0]   int_reg_array_15_25_real;
  reg        [15:0]   int_reg_array_15_25_imag;
  reg        [15:0]   int_reg_array_15_26_real;
  reg        [15:0]   int_reg_array_15_26_imag;
  reg        [15:0]   int_reg_array_15_27_real;
  reg        [15:0]   int_reg_array_15_27_imag;
  reg        [15:0]   int_reg_array_15_28_real;
  reg        [15:0]   int_reg_array_15_28_imag;
  reg        [15:0]   int_reg_array_15_29_real;
  reg        [15:0]   int_reg_array_15_29_imag;
  reg        [15:0]   int_reg_array_15_30_real;
  reg        [15:0]   int_reg_array_15_30_imag;
  reg        [15:0]   int_reg_array_15_31_real;
  reg        [15:0]   int_reg_array_15_31_imag;
  reg        [15:0]   int_reg_array_15_32_real;
  reg        [15:0]   int_reg_array_15_32_imag;
  reg        [15:0]   int_reg_array_15_33_real;
  reg        [15:0]   int_reg_array_15_33_imag;
  reg        [15:0]   int_reg_array_15_34_real;
  reg        [15:0]   int_reg_array_15_34_imag;
  reg        [15:0]   int_reg_array_15_35_real;
  reg        [15:0]   int_reg_array_15_35_imag;
  reg        [15:0]   int_reg_array_15_36_real;
  reg        [15:0]   int_reg_array_15_36_imag;
  reg        [15:0]   int_reg_array_15_37_real;
  reg        [15:0]   int_reg_array_15_37_imag;
  reg        [15:0]   int_reg_array_15_38_real;
  reg        [15:0]   int_reg_array_15_38_imag;
  reg        [15:0]   int_reg_array_15_39_real;
  reg        [15:0]   int_reg_array_15_39_imag;
  reg        [15:0]   int_reg_array_15_40_real;
  reg        [15:0]   int_reg_array_15_40_imag;
  reg        [15:0]   int_reg_array_15_41_real;
  reg        [15:0]   int_reg_array_15_41_imag;
  reg        [15:0]   int_reg_array_15_42_real;
  reg        [15:0]   int_reg_array_15_42_imag;
  reg        [15:0]   int_reg_array_15_43_real;
  reg        [15:0]   int_reg_array_15_43_imag;
  reg        [15:0]   int_reg_array_15_44_real;
  reg        [15:0]   int_reg_array_15_44_imag;
  reg        [15:0]   int_reg_array_15_45_real;
  reg        [15:0]   int_reg_array_15_45_imag;
  reg        [15:0]   int_reg_array_15_46_real;
  reg        [15:0]   int_reg_array_15_46_imag;
  reg        [15:0]   int_reg_array_15_47_real;
  reg        [15:0]   int_reg_array_15_47_imag;
  reg        [15:0]   int_reg_array_15_48_real;
  reg        [15:0]   int_reg_array_15_48_imag;
  reg        [15:0]   int_reg_array_15_49_real;
  reg        [15:0]   int_reg_array_15_49_imag;
  reg        [15:0]   int_reg_array_15_50_real;
  reg        [15:0]   int_reg_array_15_50_imag;
  reg        [15:0]   int_reg_array_15_51_real;
  reg        [15:0]   int_reg_array_15_51_imag;
  reg        [15:0]   int_reg_array_15_52_real;
  reg        [15:0]   int_reg_array_15_52_imag;
  reg        [15:0]   int_reg_array_15_53_real;
  reg        [15:0]   int_reg_array_15_53_imag;
  reg        [15:0]   int_reg_array_15_54_real;
  reg        [15:0]   int_reg_array_15_54_imag;
  reg        [15:0]   int_reg_array_15_55_real;
  reg        [15:0]   int_reg_array_15_55_imag;
  reg        [15:0]   int_reg_array_15_56_real;
  reg        [15:0]   int_reg_array_15_56_imag;
  reg        [15:0]   int_reg_array_15_57_real;
  reg        [15:0]   int_reg_array_15_57_imag;
  reg        [15:0]   int_reg_array_15_58_real;
  reg        [15:0]   int_reg_array_15_58_imag;
  reg        [15:0]   int_reg_array_15_59_real;
  reg        [15:0]   int_reg_array_15_59_imag;
  reg        [15:0]   int_reg_array_15_60_real;
  reg        [15:0]   int_reg_array_15_60_imag;
  reg        [15:0]   int_reg_array_15_61_real;
  reg        [15:0]   int_reg_array_15_61_imag;
  reg        [15:0]   int_reg_array_15_62_real;
  reg        [15:0]   int_reg_array_15_62_imag;
  reg        [15:0]   int_reg_array_15_63_real;
  reg        [15:0]   int_reg_array_15_63_imag;
  reg        [15:0]   int_reg_array_35_0_real;
  reg        [15:0]   int_reg_array_35_0_imag;
  reg        [15:0]   int_reg_array_35_1_real;
  reg        [15:0]   int_reg_array_35_1_imag;
  reg        [15:0]   int_reg_array_35_2_real;
  reg        [15:0]   int_reg_array_35_2_imag;
  reg        [15:0]   int_reg_array_35_3_real;
  reg        [15:0]   int_reg_array_35_3_imag;
  reg        [15:0]   int_reg_array_35_4_real;
  reg        [15:0]   int_reg_array_35_4_imag;
  reg        [15:0]   int_reg_array_35_5_real;
  reg        [15:0]   int_reg_array_35_5_imag;
  reg        [15:0]   int_reg_array_35_6_real;
  reg        [15:0]   int_reg_array_35_6_imag;
  reg        [15:0]   int_reg_array_35_7_real;
  reg        [15:0]   int_reg_array_35_7_imag;
  reg        [15:0]   int_reg_array_35_8_real;
  reg        [15:0]   int_reg_array_35_8_imag;
  reg        [15:0]   int_reg_array_35_9_real;
  reg        [15:0]   int_reg_array_35_9_imag;
  reg        [15:0]   int_reg_array_35_10_real;
  reg        [15:0]   int_reg_array_35_10_imag;
  reg        [15:0]   int_reg_array_35_11_real;
  reg        [15:0]   int_reg_array_35_11_imag;
  reg        [15:0]   int_reg_array_35_12_real;
  reg        [15:0]   int_reg_array_35_12_imag;
  reg        [15:0]   int_reg_array_35_13_real;
  reg        [15:0]   int_reg_array_35_13_imag;
  reg        [15:0]   int_reg_array_35_14_real;
  reg        [15:0]   int_reg_array_35_14_imag;
  reg        [15:0]   int_reg_array_35_15_real;
  reg        [15:0]   int_reg_array_35_15_imag;
  reg        [15:0]   int_reg_array_35_16_real;
  reg        [15:0]   int_reg_array_35_16_imag;
  reg        [15:0]   int_reg_array_35_17_real;
  reg        [15:0]   int_reg_array_35_17_imag;
  reg        [15:0]   int_reg_array_35_18_real;
  reg        [15:0]   int_reg_array_35_18_imag;
  reg        [15:0]   int_reg_array_35_19_real;
  reg        [15:0]   int_reg_array_35_19_imag;
  reg        [15:0]   int_reg_array_35_20_real;
  reg        [15:0]   int_reg_array_35_20_imag;
  reg        [15:0]   int_reg_array_35_21_real;
  reg        [15:0]   int_reg_array_35_21_imag;
  reg        [15:0]   int_reg_array_35_22_real;
  reg        [15:0]   int_reg_array_35_22_imag;
  reg        [15:0]   int_reg_array_35_23_real;
  reg        [15:0]   int_reg_array_35_23_imag;
  reg        [15:0]   int_reg_array_35_24_real;
  reg        [15:0]   int_reg_array_35_24_imag;
  reg        [15:0]   int_reg_array_35_25_real;
  reg        [15:0]   int_reg_array_35_25_imag;
  reg        [15:0]   int_reg_array_35_26_real;
  reg        [15:0]   int_reg_array_35_26_imag;
  reg        [15:0]   int_reg_array_35_27_real;
  reg        [15:0]   int_reg_array_35_27_imag;
  reg        [15:0]   int_reg_array_35_28_real;
  reg        [15:0]   int_reg_array_35_28_imag;
  reg        [15:0]   int_reg_array_35_29_real;
  reg        [15:0]   int_reg_array_35_29_imag;
  reg        [15:0]   int_reg_array_35_30_real;
  reg        [15:0]   int_reg_array_35_30_imag;
  reg        [15:0]   int_reg_array_35_31_real;
  reg        [15:0]   int_reg_array_35_31_imag;
  reg        [15:0]   int_reg_array_35_32_real;
  reg        [15:0]   int_reg_array_35_32_imag;
  reg        [15:0]   int_reg_array_35_33_real;
  reg        [15:0]   int_reg_array_35_33_imag;
  reg        [15:0]   int_reg_array_35_34_real;
  reg        [15:0]   int_reg_array_35_34_imag;
  reg        [15:0]   int_reg_array_35_35_real;
  reg        [15:0]   int_reg_array_35_35_imag;
  reg        [15:0]   int_reg_array_35_36_real;
  reg        [15:0]   int_reg_array_35_36_imag;
  reg        [15:0]   int_reg_array_35_37_real;
  reg        [15:0]   int_reg_array_35_37_imag;
  reg        [15:0]   int_reg_array_35_38_real;
  reg        [15:0]   int_reg_array_35_38_imag;
  reg        [15:0]   int_reg_array_35_39_real;
  reg        [15:0]   int_reg_array_35_39_imag;
  reg        [15:0]   int_reg_array_35_40_real;
  reg        [15:0]   int_reg_array_35_40_imag;
  reg        [15:0]   int_reg_array_35_41_real;
  reg        [15:0]   int_reg_array_35_41_imag;
  reg        [15:0]   int_reg_array_35_42_real;
  reg        [15:0]   int_reg_array_35_42_imag;
  reg        [15:0]   int_reg_array_35_43_real;
  reg        [15:0]   int_reg_array_35_43_imag;
  reg        [15:0]   int_reg_array_35_44_real;
  reg        [15:0]   int_reg_array_35_44_imag;
  reg        [15:0]   int_reg_array_35_45_real;
  reg        [15:0]   int_reg_array_35_45_imag;
  reg        [15:0]   int_reg_array_35_46_real;
  reg        [15:0]   int_reg_array_35_46_imag;
  reg        [15:0]   int_reg_array_35_47_real;
  reg        [15:0]   int_reg_array_35_47_imag;
  reg        [15:0]   int_reg_array_35_48_real;
  reg        [15:0]   int_reg_array_35_48_imag;
  reg        [15:0]   int_reg_array_35_49_real;
  reg        [15:0]   int_reg_array_35_49_imag;
  reg        [15:0]   int_reg_array_35_50_real;
  reg        [15:0]   int_reg_array_35_50_imag;
  reg        [15:0]   int_reg_array_35_51_real;
  reg        [15:0]   int_reg_array_35_51_imag;
  reg        [15:0]   int_reg_array_35_52_real;
  reg        [15:0]   int_reg_array_35_52_imag;
  reg        [15:0]   int_reg_array_35_53_real;
  reg        [15:0]   int_reg_array_35_53_imag;
  reg        [15:0]   int_reg_array_35_54_real;
  reg        [15:0]   int_reg_array_35_54_imag;
  reg        [15:0]   int_reg_array_35_55_real;
  reg        [15:0]   int_reg_array_35_55_imag;
  reg        [15:0]   int_reg_array_35_56_real;
  reg        [15:0]   int_reg_array_35_56_imag;
  reg        [15:0]   int_reg_array_35_57_real;
  reg        [15:0]   int_reg_array_35_57_imag;
  reg        [15:0]   int_reg_array_35_58_real;
  reg        [15:0]   int_reg_array_35_58_imag;
  reg        [15:0]   int_reg_array_35_59_real;
  reg        [15:0]   int_reg_array_35_59_imag;
  reg        [15:0]   int_reg_array_35_60_real;
  reg        [15:0]   int_reg_array_35_60_imag;
  reg        [15:0]   int_reg_array_35_61_real;
  reg        [15:0]   int_reg_array_35_61_imag;
  reg        [15:0]   int_reg_array_35_62_real;
  reg        [15:0]   int_reg_array_35_62_imag;
  reg        [15:0]   int_reg_array_35_63_real;
  reg        [15:0]   int_reg_array_35_63_imag;
  reg        [15:0]   int_reg_array_45_0_real;
  reg        [15:0]   int_reg_array_45_0_imag;
  reg        [15:0]   int_reg_array_45_1_real;
  reg        [15:0]   int_reg_array_45_1_imag;
  reg        [15:0]   int_reg_array_45_2_real;
  reg        [15:0]   int_reg_array_45_2_imag;
  reg        [15:0]   int_reg_array_45_3_real;
  reg        [15:0]   int_reg_array_45_3_imag;
  reg        [15:0]   int_reg_array_45_4_real;
  reg        [15:0]   int_reg_array_45_4_imag;
  reg        [15:0]   int_reg_array_45_5_real;
  reg        [15:0]   int_reg_array_45_5_imag;
  reg        [15:0]   int_reg_array_45_6_real;
  reg        [15:0]   int_reg_array_45_6_imag;
  reg        [15:0]   int_reg_array_45_7_real;
  reg        [15:0]   int_reg_array_45_7_imag;
  reg        [15:0]   int_reg_array_45_8_real;
  reg        [15:0]   int_reg_array_45_8_imag;
  reg        [15:0]   int_reg_array_45_9_real;
  reg        [15:0]   int_reg_array_45_9_imag;
  reg        [15:0]   int_reg_array_45_10_real;
  reg        [15:0]   int_reg_array_45_10_imag;
  reg        [15:0]   int_reg_array_45_11_real;
  reg        [15:0]   int_reg_array_45_11_imag;
  reg        [15:0]   int_reg_array_45_12_real;
  reg        [15:0]   int_reg_array_45_12_imag;
  reg        [15:0]   int_reg_array_45_13_real;
  reg        [15:0]   int_reg_array_45_13_imag;
  reg        [15:0]   int_reg_array_45_14_real;
  reg        [15:0]   int_reg_array_45_14_imag;
  reg        [15:0]   int_reg_array_45_15_real;
  reg        [15:0]   int_reg_array_45_15_imag;
  reg        [15:0]   int_reg_array_45_16_real;
  reg        [15:0]   int_reg_array_45_16_imag;
  reg        [15:0]   int_reg_array_45_17_real;
  reg        [15:0]   int_reg_array_45_17_imag;
  reg        [15:0]   int_reg_array_45_18_real;
  reg        [15:0]   int_reg_array_45_18_imag;
  reg        [15:0]   int_reg_array_45_19_real;
  reg        [15:0]   int_reg_array_45_19_imag;
  reg        [15:0]   int_reg_array_45_20_real;
  reg        [15:0]   int_reg_array_45_20_imag;
  reg        [15:0]   int_reg_array_45_21_real;
  reg        [15:0]   int_reg_array_45_21_imag;
  reg        [15:0]   int_reg_array_45_22_real;
  reg        [15:0]   int_reg_array_45_22_imag;
  reg        [15:0]   int_reg_array_45_23_real;
  reg        [15:0]   int_reg_array_45_23_imag;
  reg        [15:0]   int_reg_array_45_24_real;
  reg        [15:0]   int_reg_array_45_24_imag;
  reg        [15:0]   int_reg_array_45_25_real;
  reg        [15:0]   int_reg_array_45_25_imag;
  reg        [15:0]   int_reg_array_45_26_real;
  reg        [15:0]   int_reg_array_45_26_imag;
  reg        [15:0]   int_reg_array_45_27_real;
  reg        [15:0]   int_reg_array_45_27_imag;
  reg        [15:0]   int_reg_array_45_28_real;
  reg        [15:0]   int_reg_array_45_28_imag;
  reg        [15:0]   int_reg_array_45_29_real;
  reg        [15:0]   int_reg_array_45_29_imag;
  reg        [15:0]   int_reg_array_45_30_real;
  reg        [15:0]   int_reg_array_45_30_imag;
  reg        [15:0]   int_reg_array_45_31_real;
  reg        [15:0]   int_reg_array_45_31_imag;
  reg        [15:0]   int_reg_array_45_32_real;
  reg        [15:0]   int_reg_array_45_32_imag;
  reg        [15:0]   int_reg_array_45_33_real;
  reg        [15:0]   int_reg_array_45_33_imag;
  reg        [15:0]   int_reg_array_45_34_real;
  reg        [15:0]   int_reg_array_45_34_imag;
  reg        [15:0]   int_reg_array_45_35_real;
  reg        [15:0]   int_reg_array_45_35_imag;
  reg        [15:0]   int_reg_array_45_36_real;
  reg        [15:0]   int_reg_array_45_36_imag;
  reg        [15:0]   int_reg_array_45_37_real;
  reg        [15:0]   int_reg_array_45_37_imag;
  reg        [15:0]   int_reg_array_45_38_real;
  reg        [15:0]   int_reg_array_45_38_imag;
  reg        [15:0]   int_reg_array_45_39_real;
  reg        [15:0]   int_reg_array_45_39_imag;
  reg        [15:0]   int_reg_array_45_40_real;
  reg        [15:0]   int_reg_array_45_40_imag;
  reg        [15:0]   int_reg_array_45_41_real;
  reg        [15:0]   int_reg_array_45_41_imag;
  reg        [15:0]   int_reg_array_45_42_real;
  reg        [15:0]   int_reg_array_45_42_imag;
  reg        [15:0]   int_reg_array_45_43_real;
  reg        [15:0]   int_reg_array_45_43_imag;
  reg        [15:0]   int_reg_array_45_44_real;
  reg        [15:0]   int_reg_array_45_44_imag;
  reg        [15:0]   int_reg_array_45_45_real;
  reg        [15:0]   int_reg_array_45_45_imag;
  reg        [15:0]   int_reg_array_45_46_real;
  reg        [15:0]   int_reg_array_45_46_imag;
  reg        [15:0]   int_reg_array_45_47_real;
  reg        [15:0]   int_reg_array_45_47_imag;
  reg        [15:0]   int_reg_array_45_48_real;
  reg        [15:0]   int_reg_array_45_48_imag;
  reg        [15:0]   int_reg_array_45_49_real;
  reg        [15:0]   int_reg_array_45_49_imag;
  reg        [15:0]   int_reg_array_45_50_real;
  reg        [15:0]   int_reg_array_45_50_imag;
  reg        [15:0]   int_reg_array_45_51_real;
  reg        [15:0]   int_reg_array_45_51_imag;
  reg        [15:0]   int_reg_array_45_52_real;
  reg        [15:0]   int_reg_array_45_52_imag;
  reg        [15:0]   int_reg_array_45_53_real;
  reg        [15:0]   int_reg_array_45_53_imag;
  reg        [15:0]   int_reg_array_45_54_real;
  reg        [15:0]   int_reg_array_45_54_imag;
  reg        [15:0]   int_reg_array_45_55_real;
  reg        [15:0]   int_reg_array_45_55_imag;
  reg        [15:0]   int_reg_array_45_56_real;
  reg        [15:0]   int_reg_array_45_56_imag;
  reg        [15:0]   int_reg_array_45_57_real;
  reg        [15:0]   int_reg_array_45_57_imag;
  reg        [15:0]   int_reg_array_45_58_real;
  reg        [15:0]   int_reg_array_45_58_imag;
  reg        [15:0]   int_reg_array_45_59_real;
  reg        [15:0]   int_reg_array_45_59_imag;
  reg        [15:0]   int_reg_array_45_60_real;
  reg        [15:0]   int_reg_array_45_60_imag;
  reg        [15:0]   int_reg_array_45_61_real;
  reg        [15:0]   int_reg_array_45_61_imag;
  reg        [15:0]   int_reg_array_45_62_real;
  reg        [15:0]   int_reg_array_45_62_imag;
  reg        [15:0]   int_reg_array_45_63_real;
  reg        [15:0]   int_reg_array_45_63_imag;
  reg        [15:0]   int_reg_array_8_0_real;
  reg        [15:0]   int_reg_array_8_0_imag;
  reg        [15:0]   int_reg_array_8_1_real;
  reg        [15:0]   int_reg_array_8_1_imag;
  reg        [15:0]   int_reg_array_8_2_real;
  reg        [15:0]   int_reg_array_8_2_imag;
  reg        [15:0]   int_reg_array_8_3_real;
  reg        [15:0]   int_reg_array_8_3_imag;
  reg        [15:0]   int_reg_array_8_4_real;
  reg        [15:0]   int_reg_array_8_4_imag;
  reg        [15:0]   int_reg_array_8_5_real;
  reg        [15:0]   int_reg_array_8_5_imag;
  reg        [15:0]   int_reg_array_8_6_real;
  reg        [15:0]   int_reg_array_8_6_imag;
  reg        [15:0]   int_reg_array_8_7_real;
  reg        [15:0]   int_reg_array_8_7_imag;
  reg        [15:0]   int_reg_array_8_8_real;
  reg        [15:0]   int_reg_array_8_8_imag;
  reg        [15:0]   int_reg_array_8_9_real;
  reg        [15:0]   int_reg_array_8_9_imag;
  reg        [15:0]   int_reg_array_8_10_real;
  reg        [15:0]   int_reg_array_8_10_imag;
  reg        [15:0]   int_reg_array_8_11_real;
  reg        [15:0]   int_reg_array_8_11_imag;
  reg        [15:0]   int_reg_array_8_12_real;
  reg        [15:0]   int_reg_array_8_12_imag;
  reg        [15:0]   int_reg_array_8_13_real;
  reg        [15:0]   int_reg_array_8_13_imag;
  reg        [15:0]   int_reg_array_8_14_real;
  reg        [15:0]   int_reg_array_8_14_imag;
  reg        [15:0]   int_reg_array_8_15_real;
  reg        [15:0]   int_reg_array_8_15_imag;
  reg        [15:0]   int_reg_array_8_16_real;
  reg        [15:0]   int_reg_array_8_16_imag;
  reg        [15:0]   int_reg_array_8_17_real;
  reg        [15:0]   int_reg_array_8_17_imag;
  reg        [15:0]   int_reg_array_8_18_real;
  reg        [15:0]   int_reg_array_8_18_imag;
  reg        [15:0]   int_reg_array_8_19_real;
  reg        [15:0]   int_reg_array_8_19_imag;
  reg        [15:0]   int_reg_array_8_20_real;
  reg        [15:0]   int_reg_array_8_20_imag;
  reg        [15:0]   int_reg_array_8_21_real;
  reg        [15:0]   int_reg_array_8_21_imag;
  reg        [15:0]   int_reg_array_8_22_real;
  reg        [15:0]   int_reg_array_8_22_imag;
  reg        [15:0]   int_reg_array_8_23_real;
  reg        [15:0]   int_reg_array_8_23_imag;
  reg        [15:0]   int_reg_array_8_24_real;
  reg        [15:0]   int_reg_array_8_24_imag;
  reg        [15:0]   int_reg_array_8_25_real;
  reg        [15:0]   int_reg_array_8_25_imag;
  reg        [15:0]   int_reg_array_8_26_real;
  reg        [15:0]   int_reg_array_8_26_imag;
  reg        [15:0]   int_reg_array_8_27_real;
  reg        [15:0]   int_reg_array_8_27_imag;
  reg        [15:0]   int_reg_array_8_28_real;
  reg        [15:0]   int_reg_array_8_28_imag;
  reg        [15:0]   int_reg_array_8_29_real;
  reg        [15:0]   int_reg_array_8_29_imag;
  reg        [15:0]   int_reg_array_8_30_real;
  reg        [15:0]   int_reg_array_8_30_imag;
  reg        [15:0]   int_reg_array_8_31_real;
  reg        [15:0]   int_reg_array_8_31_imag;
  reg        [15:0]   int_reg_array_8_32_real;
  reg        [15:0]   int_reg_array_8_32_imag;
  reg        [15:0]   int_reg_array_8_33_real;
  reg        [15:0]   int_reg_array_8_33_imag;
  reg        [15:0]   int_reg_array_8_34_real;
  reg        [15:0]   int_reg_array_8_34_imag;
  reg        [15:0]   int_reg_array_8_35_real;
  reg        [15:0]   int_reg_array_8_35_imag;
  reg        [15:0]   int_reg_array_8_36_real;
  reg        [15:0]   int_reg_array_8_36_imag;
  reg        [15:0]   int_reg_array_8_37_real;
  reg        [15:0]   int_reg_array_8_37_imag;
  reg        [15:0]   int_reg_array_8_38_real;
  reg        [15:0]   int_reg_array_8_38_imag;
  reg        [15:0]   int_reg_array_8_39_real;
  reg        [15:0]   int_reg_array_8_39_imag;
  reg        [15:0]   int_reg_array_8_40_real;
  reg        [15:0]   int_reg_array_8_40_imag;
  reg        [15:0]   int_reg_array_8_41_real;
  reg        [15:0]   int_reg_array_8_41_imag;
  reg        [15:0]   int_reg_array_8_42_real;
  reg        [15:0]   int_reg_array_8_42_imag;
  reg        [15:0]   int_reg_array_8_43_real;
  reg        [15:0]   int_reg_array_8_43_imag;
  reg        [15:0]   int_reg_array_8_44_real;
  reg        [15:0]   int_reg_array_8_44_imag;
  reg        [15:0]   int_reg_array_8_45_real;
  reg        [15:0]   int_reg_array_8_45_imag;
  reg        [15:0]   int_reg_array_8_46_real;
  reg        [15:0]   int_reg_array_8_46_imag;
  reg        [15:0]   int_reg_array_8_47_real;
  reg        [15:0]   int_reg_array_8_47_imag;
  reg        [15:0]   int_reg_array_8_48_real;
  reg        [15:0]   int_reg_array_8_48_imag;
  reg        [15:0]   int_reg_array_8_49_real;
  reg        [15:0]   int_reg_array_8_49_imag;
  reg        [15:0]   int_reg_array_8_50_real;
  reg        [15:0]   int_reg_array_8_50_imag;
  reg        [15:0]   int_reg_array_8_51_real;
  reg        [15:0]   int_reg_array_8_51_imag;
  reg        [15:0]   int_reg_array_8_52_real;
  reg        [15:0]   int_reg_array_8_52_imag;
  reg        [15:0]   int_reg_array_8_53_real;
  reg        [15:0]   int_reg_array_8_53_imag;
  reg        [15:0]   int_reg_array_8_54_real;
  reg        [15:0]   int_reg_array_8_54_imag;
  reg        [15:0]   int_reg_array_8_55_real;
  reg        [15:0]   int_reg_array_8_55_imag;
  reg        [15:0]   int_reg_array_8_56_real;
  reg        [15:0]   int_reg_array_8_56_imag;
  reg        [15:0]   int_reg_array_8_57_real;
  reg        [15:0]   int_reg_array_8_57_imag;
  reg        [15:0]   int_reg_array_8_58_real;
  reg        [15:0]   int_reg_array_8_58_imag;
  reg        [15:0]   int_reg_array_8_59_real;
  reg        [15:0]   int_reg_array_8_59_imag;
  reg        [15:0]   int_reg_array_8_60_real;
  reg        [15:0]   int_reg_array_8_60_imag;
  reg        [15:0]   int_reg_array_8_61_real;
  reg        [15:0]   int_reg_array_8_61_imag;
  reg        [15:0]   int_reg_array_8_62_real;
  reg        [15:0]   int_reg_array_8_62_imag;
  reg        [15:0]   int_reg_array_8_63_real;
  reg        [15:0]   int_reg_array_8_63_imag;
  reg        [15:0]   int_reg_array_58_0_real;
  reg        [15:0]   int_reg_array_58_0_imag;
  reg        [15:0]   int_reg_array_58_1_real;
  reg        [15:0]   int_reg_array_58_1_imag;
  reg        [15:0]   int_reg_array_58_2_real;
  reg        [15:0]   int_reg_array_58_2_imag;
  reg        [15:0]   int_reg_array_58_3_real;
  reg        [15:0]   int_reg_array_58_3_imag;
  reg        [15:0]   int_reg_array_58_4_real;
  reg        [15:0]   int_reg_array_58_4_imag;
  reg        [15:0]   int_reg_array_58_5_real;
  reg        [15:0]   int_reg_array_58_5_imag;
  reg        [15:0]   int_reg_array_58_6_real;
  reg        [15:0]   int_reg_array_58_6_imag;
  reg        [15:0]   int_reg_array_58_7_real;
  reg        [15:0]   int_reg_array_58_7_imag;
  reg        [15:0]   int_reg_array_58_8_real;
  reg        [15:0]   int_reg_array_58_8_imag;
  reg        [15:0]   int_reg_array_58_9_real;
  reg        [15:0]   int_reg_array_58_9_imag;
  reg        [15:0]   int_reg_array_58_10_real;
  reg        [15:0]   int_reg_array_58_10_imag;
  reg        [15:0]   int_reg_array_58_11_real;
  reg        [15:0]   int_reg_array_58_11_imag;
  reg        [15:0]   int_reg_array_58_12_real;
  reg        [15:0]   int_reg_array_58_12_imag;
  reg        [15:0]   int_reg_array_58_13_real;
  reg        [15:0]   int_reg_array_58_13_imag;
  reg        [15:0]   int_reg_array_58_14_real;
  reg        [15:0]   int_reg_array_58_14_imag;
  reg        [15:0]   int_reg_array_58_15_real;
  reg        [15:0]   int_reg_array_58_15_imag;
  reg        [15:0]   int_reg_array_58_16_real;
  reg        [15:0]   int_reg_array_58_16_imag;
  reg        [15:0]   int_reg_array_58_17_real;
  reg        [15:0]   int_reg_array_58_17_imag;
  reg        [15:0]   int_reg_array_58_18_real;
  reg        [15:0]   int_reg_array_58_18_imag;
  reg        [15:0]   int_reg_array_58_19_real;
  reg        [15:0]   int_reg_array_58_19_imag;
  reg        [15:0]   int_reg_array_58_20_real;
  reg        [15:0]   int_reg_array_58_20_imag;
  reg        [15:0]   int_reg_array_58_21_real;
  reg        [15:0]   int_reg_array_58_21_imag;
  reg        [15:0]   int_reg_array_58_22_real;
  reg        [15:0]   int_reg_array_58_22_imag;
  reg        [15:0]   int_reg_array_58_23_real;
  reg        [15:0]   int_reg_array_58_23_imag;
  reg        [15:0]   int_reg_array_58_24_real;
  reg        [15:0]   int_reg_array_58_24_imag;
  reg        [15:0]   int_reg_array_58_25_real;
  reg        [15:0]   int_reg_array_58_25_imag;
  reg        [15:0]   int_reg_array_58_26_real;
  reg        [15:0]   int_reg_array_58_26_imag;
  reg        [15:0]   int_reg_array_58_27_real;
  reg        [15:0]   int_reg_array_58_27_imag;
  reg        [15:0]   int_reg_array_58_28_real;
  reg        [15:0]   int_reg_array_58_28_imag;
  reg        [15:0]   int_reg_array_58_29_real;
  reg        [15:0]   int_reg_array_58_29_imag;
  reg        [15:0]   int_reg_array_58_30_real;
  reg        [15:0]   int_reg_array_58_30_imag;
  reg        [15:0]   int_reg_array_58_31_real;
  reg        [15:0]   int_reg_array_58_31_imag;
  reg        [15:0]   int_reg_array_58_32_real;
  reg        [15:0]   int_reg_array_58_32_imag;
  reg        [15:0]   int_reg_array_58_33_real;
  reg        [15:0]   int_reg_array_58_33_imag;
  reg        [15:0]   int_reg_array_58_34_real;
  reg        [15:0]   int_reg_array_58_34_imag;
  reg        [15:0]   int_reg_array_58_35_real;
  reg        [15:0]   int_reg_array_58_35_imag;
  reg        [15:0]   int_reg_array_58_36_real;
  reg        [15:0]   int_reg_array_58_36_imag;
  reg        [15:0]   int_reg_array_58_37_real;
  reg        [15:0]   int_reg_array_58_37_imag;
  reg        [15:0]   int_reg_array_58_38_real;
  reg        [15:0]   int_reg_array_58_38_imag;
  reg        [15:0]   int_reg_array_58_39_real;
  reg        [15:0]   int_reg_array_58_39_imag;
  reg        [15:0]   int_reg_array_58_40_real;
  reg        [15:0]   int_reg_array_58_40_imag;
  reg        [15:0]   int_reg_array_58_41_real;
  reg        [15:0]   int_reg_array_58_41_imag;
  reg        [15:0]   int_reg_array_58_42_real;
  reg        [15:0]   int_reg_array_58_42_imag;
  reg        [15:0]   int_reg_array_58_43_real;
  reg        [15:0]   int_reg_array_58_43_imag;
  reg        [15:0]   int_reg_array_58_44_real;
  reg        [15:0]   int_reg_array_58_44_imag;
  reg        [15:0]   int_reg_array_58_45_real;
  reg        [15:0]   int_reg_array_58_45_imag;
  reg        [15:0]   int_reg_array_58_46_real;
  reg        [15:0]   int_reg_array_58_46_imag;
  reg        [15:0]   int_reg_array_58_47_real;
  reg        [15:0]   int_reg_array_58_47_imag;
  reg        [15:0]   int_reg_array_58_48_real;
  reg        [15:0]   int_reg_array_58_48_imag;
  reg        [15:0]   int_reg_array_58_49_real;
  reg        [15:0]   int_reg_array_58_49_imag;
  reg        [15:0]   int_reg_array_58_50_real;
  reg        [15:0]   int_reg_array_58_50_imag;
  reg        [15:0]   int_reg_array_58_51_real;
  reg        [15:0]   int_reg_array_58_51_imag;
  reg        [15:0]   int_reg_array_58_52_real;
  reg        [15:0]   int_reg_array_58_52_imag;
  reg        [15:0]   int_reg_array_58_53_real;
  reg        [15:0]   int_reg_array_58_53_imag;
  reg        [15:0]   int_reg_array_58_54_real;
  reg        [15:0]   int_reg_array_58_54_imag;
  reg        [15:0]   int_reg_array_58_55_real;
  reg        [15:0]   int_reg_array_58_55_imag;
  reg        [15:0]   int_reg_array_58_56_real;
  reg        [15:0]   int_reg_array_58_56_imag;
  reg        [15:0]   int_reg_array_58_57_real;
  reg        [15:0]   int_reg_array_58_57_imag;
  reg        [15:0]   int_reg_array_58_58_real;
  reg        [15:0]   int_reg_array_58_58_imag;
  reg        [15:0]   int_reg_array_58_59_real;
  reg        [15:0]   int_reg_array_58_59_imag;
  reg        [15:0]   int_reg_array_58_60_real;
  reg        [15:0]   int_reg_array_58_60_imag;
  reg        [15:0]   int_reg_array_58_61_real;
  reg        [15:0]   int_reg_array_58_61_imag;
  reg        [15:0]   int_reg_array_58_62_real;
  reg        [15:0]   int_reg_array_58_62_imag;
  reg        [15:0]   int_reg_array_58_63_real;
  reg        [15:0]   int_reg_array_58_63_imag;
  reg        [15:0]   int_reg_array_42_0_real;
  reg        [15:0]   int_reg_array_42_0_imag;
  reg        [15:0]   int_reg_array_42_1_real;
  reg        [15:0]   int_reg_array_42_1_imag;
  reg        [15:0]   int_reg_array_42_2_real;
  reg        [15:0]   int_reg_array_42_2_imag;
  reg        [15:0]   int_reg_array_42_3_real;
  reg        [15:0]   int_reg_array_42_3_imag;
  reg        [15:0]   int_reg_array_42_4_real;
  reg        [15:0]   int_reg_array_42_4_imag;
  reg        [15:0]   int_reg_array_42_5_real;
  reg        [15:0]   int_reg_array_42_5_imag;
  reg        [15:0]   int_reg_array_42_6_real;
  reg        [15:0]   int_reg_array_42_6_imag;
  reg        [15:0]   int_reg_array_42_7_real;
  reg        [15:0]   int_reg_array_42_7_imag;
  reg        [15:0]   int_reg_array_42_8_real;
  reg        [15:0]   int_reg_array_42_8_imag;
  reg        [15:0]   int_reg_array_42_9_real;
  reg        [15:0]   int_reg_array_42_9_imag;
  reg        [15:0]   int_reg_array_42_10_real;
  reg        [15:0]   int_reg_array_42_10_imag;
  reg        [15:0]   int_reg_array_42_11_real;
  reg        [15:0]   int_reg_array_42_11_imag;
  reg        [15:0]   int_reg_array_42_12_real;
  reg        [15:0]   int_reg_array_42_12_imag;
  reg        [15:0]   int_reg_array_42_13_real;
  reg        [15:0]   int_reg_array_42_13_imag;
  reg        [15:0]   int_reg_array_42_14_real;
  reg        [15:0]   int_reg_array_42_14_imag;
  reg        [15:0]   int_reg_array_42_15_real;
  reg        [15:0]   int_reg_array_42_15_imag;
  reg        [15:0]   int_reg_array_42_16_real;
  reg        [15:0]   int_reg_array_42_16_imag;
  reg        [15:0]   int_reg_array_42_17_real;
  reg        [15:0]   int_reg_array_42_17_imag;
  reg        [15:0]   int_reg_array_42_18_real;
  reg        [15:0]   int_reg_array_42_18_imag;
  reg        [15:0]   int_reg_array_42_19_real;
  reg        [15:0]   int_reg_array_42_19_imag;
  reg        [15:0]   int_reg_array_42_20_real;
  reg        [15:0]   int_reg_array_42_20_imag;
  reg        [15:0]   int_reg_array_42_21_real;
  reg        [15:0]   int_reg_array_42_21_imag;
  reg        [15:0]   int_reg_array_42_22_real;
  reg        [15:0]   int_reg_array_42_22_imag;
  reg        [15:0]   int_reg_array_42_23_real;
  reg        [15:0]   int_reg_array_42_23_imag;
  reg        [15:0]   int_reg_array_42_24_real;
  reg        [15:0]   int_reg_array_42_24_imag;
  reg        [15:0]   int_reg_array_42_25_real;
  reg        [15:0]   int_reg_array_42_25_imag;
  reg        [15:0]   int_reg_array_42_26_real;
  reg        [15:0]   int_reg_array_42_26_imag;
  reg        [15:0]   int_reg_array_42_27_real;
  reg        [15:0]   int_reg_array_42_27_imag;
  reg        [15:0]   int_reg_array_42_28_real;
  reg        [15:0]   int_reg_array_42_28_imag;
  reg        [15:0]   int_reg_array_42_29_real;
  reg        [15:0]   int_reg_array_42_29_imag;
  reg        [15:0]   int_reg_array_42_30_real;
  reg        [15:0]   int_reg_array_42_30_imag;
  reg        [15:0]   int_reg_array_42_31_real;
  reg        [15:0]   int_reg_array_42_31_imag;
  reg        [15:0]   int_reg_array_42_32_real;
  reg        [15:0]   int_reg_array_42_32_imag;
  reg        [15:0]   int_reg_array_42_33_real;
  reg        [15:0]   int_reg_array_42_33_imag;
  reg        [15:0]   int_reg_array_42_34_real;
  reg        [15:0]   int_reg_array_42_34_imag;
  reg        [15:0]   int_reg_array_42_35_real;
  reg        [15:0]   int_reg_array_42_35_imag;
  reg        [15:0]   int_reg_array_42_36_real;
  reg        [15:0]   int_reg_array_42_36_imag;
  reg        [15:0]   int_reg_array_42_37_real;
  reg        [15:0]   int_reg_array_42_37_imag;
  reg        [15:0]   int_reg_array_42_38_real;
  reg        [15:0]   int_reg_array_42_38_imag;
  reg        [15:0]   int_reg_array_42_39_real;
  reg        [15:0]   int_reg_array_42_39_imag;
  reg        [15:0]   int_reg_array_42_40_real;
  reg        [15:0]   int_reg_array_42_40_imag;
  reg        [15:0]   int_reg_array_42_41_real;
  reg        [15:0]   int_reg_array_42_41_imag;
  reg        [15:0]   int_reg_array_42_42_real;
  reg        [15:0]   int_reg_array_42_42_imag;
  reg        [15:0]   int_reg_array_42_43_real;
  reg        [15:0]   int_reg_array_42_43_imag;
  reg        [15:0]   int_reg_array_42_44_real;
  reg        [15:0]   int_reg_array_42_44_imag;
  reg        [15:0]   int_reg_array_42_45_real;
  reg        [15:0]   int_reg_array_42_45_imag;
  reg        [15:0]   int_reg_array_42_46_real;
  reg        [15:0]   int_reg_array_42_46_imag;
  reg        [15:0]   int_reg_array_42_47_real;
  reg        [15:0]   int_reg_array_42_47_imag;
  reg        [15:0]   int_reg_array_42_48_real;
  reg        [15:0]   int_reg_array_42_48_imag;
  reg        [15:0]   int_reg_array_42_49_real;
  reg        [15:0]   int_reg_array_42_49_imag;
  reg        [15:0]   int_reg_array_42_50_real;
  reg        [15:0]   int_reg_array_42_50_imag;
  reg        [15:0]   int_reg_array_42_51_real;
  reg        [15:0]   int_reg_array_42_51_imag;
  reg        [15:0]   int_reg_array_42_52_real;
  reg        [15:0]   int_reg_array_42_52_imag;
  reg        [15:0]   int_reg_array_42_53_real;
  reg        [15:0]   int_reg_array_42_53_imag;
  reg        [15:0]   int_reg_array_42_54_real;
  reg        [15:0]   int_reg_array_42_54_imag;
  reg        [15:0]   int_reg_array_42_55_real;
  reg        [15:0]   int_reg_array_42_55_imag;
  reg        [15:0]   int_reg_array_42_56_real;
  reg        [15:0]   int_reg_array_42_56_imag;
  reg        [15:0]   int_reg_array_42_57_real;
  reg        [15:0]   int_reg_array_42_57_imag;
  reg        [15:0]   int_reg_array_42_58_real;
  reg        [15:0]   int_reg_array_42_58_imag;
  reg        [15:0]   int_reg_array_42_59_real;
  reg        [15:0]   int_reg_array_42_59_imag;
  reg        [15:0]   int_reg_array_42_60_real;
  reg        [15:0]   int_reg_array_42_60_imag;
  reg        [15:0]   int_reg_array_42_61_real;
  reg        [15:0]   int_reg_array_42_61_imag;
  reg        [15:0]   int_reg_array_42_62_real;
  reg        [15:0]   int_reg_array_42_62_imag;
  reg        [15:0]   int_reg_array_42_63_real;
  reg        [15:0]   int_reg_array_42_63_imag;
  reg        [15:0]   int_reg_array_24_0_real;
  reg        [15:0]   int_reg_array_24_0_imag;
  reg        [15:0]   int_reg_array_24_1_real;
  reg        [15:0]   int_reg_array_24_1_imag;
  reg        [15:0]   int_reg_array_24_2_real;
  reg        [15:0]   int_reg_array_24_2_imag;
  reg        [15:0]   int_reg_array_24_3_real;
  reg        [15:0]   int_reg_array_24_3_imag;
  reg        [15:0]   int_reg_array_24_4_real;
  reg        [15:0]   int_reg_array_24_4_imag;
  reg        [15:0]   int_reg_array_24_5_real;
  reg        [15:0]   int_reg_array_24_5_imag;
  reg        [15:0]   int_reg_array_24_6_real;
  reg        [15:0]   int_reg_array_24_6_imag;
  reg        [15:0]   int_reg_array_24_7_real;
  reg        [15:0]   int_reg_array_24_7_imag;
  reg        [15:0]   int_reg_array_24_8_real;
  reg        [15:0]   int_reg_array_24_8_imag;
  reg        [15:0]   int_reg_array_24_9_real;
  reg        [15:0]   int_reg_array_24_9_imag;
  reg        [15:0]   int_reg_array_24_10_real;
  reg        [15:0]   int_reg_array_24_10_imag;
  reg        [15:0]   int_reg_array_24_11_real;
  reg        [15:0]   int_reg_array_24_11_imag;
  reg        [15:0]   int_reg_array_24_12_real;
  reg        [15:0]   int_reg_array_24_12_imag;
  reg        [15:0]   int_reg_array_24_13_real;
  reg        [15:0]   int_reg_array_24_13_imag;
  reg        [15:0]   int_reg_array_24_14_real;
  reg        [15:0]   int_reg_array_24_14_imag;
  reg        [15:0]   int_reg_array_24_15_real;
  reg        [15:0]   int_reg_array_24_15_imag;
  reg        [15:0]   int_reg_array_24_16_real;
  reg        [15:0]   int_reg_array_24_16_imag;
  reg        [15:0]   int_reg_array_24_17_real;
  reg        [15:0]   int_reg_array_24_17_imag;
  reg        [15:0]   int_reg_array_24_18_real;
  reg        [15:0]   int_reg_array_24_18_imag;
  reg        [15:0]   int_reg_array_24_19_real;
  reg        [15:0]   int_reg_array_24_19_imag;
  reg        [15:0]   int_reg_array_24_20_real;
  reg        [15:0]   int_reg_array_24_20_imag;
  reg        [15:0]   int_reg_array_24_21_real;
  reg        [15:0]   int_reg_array_24_21_imag;
  reg        [15:0]   int_reg_array_24_22_real;
  reg        [15:0]   int_reg_array_24_22_imag;
  reg        [15:0]   int_reg_array_24_23_real;
  reg        [15:0]   int_reg_array_24_23_imag;
  reg        [15:0]   int_reg_array_24_24_real;
  reg        [15:0]   int_reg_array_24_24_imag;
  reg        [15:0]   int_reg_array_24_25_real;
  reg        [15:0]   int_reg_array_24_25_imag;
  reg        [15:0]   int_reg_array_24_26_real;
  reg        [15:0]   int_reg_array_24_26_imag;
  reg        [15:0]   int_reg_array_24_27_real;
  reg        [15:0]   int_reg_array_24_27_imag;
  reg        [15:0]   int_reg_array_24_28_real;
  reg        [15:0]   int_reg_array_24_28_imag;
  reg        [15:0]   int_reg_array_24_29_real;
  reg        [15:0]   int_reg_array_24_29_imag;
  reg        [15:0]   int_reg_array_24_30_real;
  reg        [15:0]   int_reg_array_24_30_imag;
  reg        [15:0]   int_reg_array_24_31_real;
  reg        [15:0]   int_reg_array_24_31_imag;
  reg        [15:0]   int_reg_array_24_32_real;
  reg        [15:0]   int_reg_array_24_32_imag;
  reg        [15:0]   int_reg_array_24_33_real;
  reg        [15:0]   int_reg_array_24_33_imag;
  reg        [15:0]   int_reg_array_24_34_real;
  reg        [15:0]   int_reg_array_24_34_imag;
  reg        [15:0]   int_reg_array_24_35_real;
  reg        [15:0]   int_reg_array_24_35_imag;
  reg        [15:0]   int_reg_array_24_36_real;
  reg        [15:0]   int_reg_array_24_36_imag;
  reg        [15:0]   int_reg_array_24_37_real;
  reg        [15:0]   int_reg_array_24_37_imag;
  reg        [15:0]   int_reg_array_24_38_real;
  reg        [15:0]   int_reg_array_24_38_imag;
  reg        [15:0]   int_reg_array_24_39_real;
  reg        [15:0]   int_reg_array_24_39_imag;
  reg        [15:0]   int_reg_array_24_40_real;
  reg        [15:0]   int_reg_array_24_40_imag;
  reg        [15:0]   int_reg_array_24_41_real;
  reg        [15:0]   int_reg_array_24_41_imag;
  reg        [15:0]   int_reg_array_24_42_real;
  reg        [15:0]   int_reg_array_24_42_imag;
  reg        [15:0]   int_reg_array_24_43_real;
  reg        [15:0]   int_reg_array_24_43_imag;
  reg        [15:0]   int_reg_array_24_44_real;
  reg        [15:0]   int_reg_array_24_44_imag;
  reg        [15:0]   int_reg_array_24_45_real;
  reg        [15:0]   int_reg_array_24_45_imag;
  reg        [15:0]   int_reg_array_24_46_real;
  reg        [15:0]   int_reg_array_24_46_imag;
  reg        [15:0]   int_reg_array_24_47_real;
  reg        [15:0]   int_reg_array_24_47_imag;
  reg        [15:0]   int_reg_array_24_48_real;
  reg        [15:0]   int_reg_array_24_48_imag;
  reg        [15:0]   int_reg_array_24_49_real;
  reg        [15:0]   int_reg_array_24_49_imag;
  reg        [15:0]   int_reg_array_24_50_real;
  reg        [15:0]   int_reg_array_24_50_imag;
  reg        [15:0]   int_reg_array_24_51_real;
  reg        [15:0]   int_reg_array_24_51_imag;
  reg        [15:0]   int_reg_array_24_52_real;
  reg        [15:0]   int_reg_array_24_52_imag;
  reg        [15:0]   int_reg_array_24_53_real;
  reg        [15:0]   int_reg_array_24_53_imag;
  reg        [15:0]   int_reg_array_24_54_real;
  reg        [15:0]   int_reg_array_24_54_imag;
  reg        [15:0]   int_reg_array_24_55_real;
  reg        [15:0]   int_reg_array_24_55_imag;
  reg        [15:0]   int_reg_array_24_56_real;
  reg        [15:0]   int_reg_array_24_56_imag;
  reg        [15:0]   int_reg_array_24_57_real;
  reg        [15:0]   int_reg_array_24_57_imag;
  reg        [15:0]   int_reg_array_24_58_real;
  reg        [15:0]   int_reg_array_24_58_imag;
  reg        [15:0]   int_reg_array_24_59_real;
  reg        [15:0]   int_reg_array_24_59_imag;
  reg        [15:0]   int_reg_array_24_60_real;
  reg        [15:0]   int_reg_array_24_60_imag;
  reg        [15:0]   int_reg_array_24_61_real;
  reg        [15:0]   int_reg_array_24_61_imag;
  reg        [15:0]   int_reg_array_24_62_real;
  reg        [15:0]   int_reg_array_24_62_imag;
  reg        [15:0]   int_reg_array_24_63_real;
  reg        [15:0]   int_reg_array_24_63_imag;
  reg        [15:0]   int_reg_array_61_0_real;
  reg        [15:0]   int_reg_array_61_0_imag;
  reg        [15:0]   int_reg_array_61_1_real;
  reg        [15:0]   int_reg_array_61_1_imag;
  reg        [15:0]   int_reg_array_61_2_real;
  reg        [15:0]   int_reg_array_61_2_imag;
  reg        [15:0]   int_reg_array_61_3_real;
  reg        [15:0]   int_reg_array_61_3_imag;
  reg        [15:0]   int_reg_array_61_4_real;
  reg        [15:0]   int_reg_array_61_4_imag;
  reg        [15:0]   int_reg_array_61_5_real;
  reg        [15:0]   int_reg_array_61_5_imag;
  reg        [15:0]   int_reg_array_61_6_real;
  reg        [15:0]   int_reg_array_61_6_imag;
  reg        [15:0]   int_reg_array_61_7_real;
  reg        [15:0]   int_reg_array_61_7_imag;
  reg        [15:0]   int_reg_array_61_8_real;
  reg        [15:0]   int_reg_array_61_8_imag;
  reg        [15:0]   int_reg_array_61_9_real;
  reg        [15:0]   int_reg_array_61_9_imag;
  reg        [15:0]   int_reg_array_61_10_real;
  reg        [15:0]   int_reg_array_61_10_imag;
  reg        [15:0]   int_reg_array_61_11_real;
  reg        [15:0]   int_reg_array_61_11_imag;
  reg        [15:0]   int_reg_array_61_12_real;
  reg        [15:0]   int_reg_array_61_12_imag;
  reg        [15:0]   int_reg_array_61_13_real;
  reg        [15:0]   int_reg_array_61_13_imag;
  reg        [15:0]   int_reg_array_61_14_real;
  reg        [15:0]   int_reg_array_61_14_imag;
  reg        [15:0]   int_reg_array_61_15_real;
  reg        [15:0]   int_reg_array_61_15_imag;
  reg        [15:0]   int_reg_array_61_16_real;
  reg        [15:0]   int_reg_array_61_16_imag;
  reg        [15:0]   int_reg_array_61_17_real;
  reg        [15:0]   int_reg_array_61_17_imag;
  reg        [15:0]   int_reg_array_61_18_real;
  reg        [15:0]   int_reg_array_61_18_imag;
  reg        [15:0]   int_reg_array_61_19_real;
  reg        [15:0]   int_reg_array_61_19_imag;
  reg        [15:0]   int_reg_array_61_20_real;
  reg        [15:0]   int_reg_array_61_20_imag;
  reg        [15:0]   int_reg_array_61_21_real;
  reg        [15:0]   int_reg_array_61_21_imag;
  reg        [15:0]   int_reg_array_61_22_real;
  reg        [15:0]   int_reg_array_61_22_imag;
  reg        [15:0]   int_reg_array_61_23_real;
  reg        [15:0]   int_reg_array_61_23_imag;
  reg        [15:0]   int_reg_array_61_24_real;
  reg        [15:0]   int_reg_array_61_24_imag;
  reg        [15:0]   int_reg_array_61_25_real;
  reg        [15:0]   int_reg_array_61_25_imag;
  reg        [15:0]   int_reg_array_61_26_real;
  reg        [15:0]   int_reg_array_61_26_imag;
  reg        [15:0]   int_reg_array_61_27_real;
  reg        [15:0]   int_reg_array_61_27_imag;
  reg        [15:0]   int_reg_array_61_28_real;
  reg        [15:0]   int_reg_array_61_28_imag;
  reg        [15:0]   int_reg_array_61_29_real;
  reg        [15:0]   int_reg_array_61_29_imag;
  reg        [15:0]   int_reg_array_61_30_real;
  reg        [15:0]   int_reg_array_61_30_imag;
  reg        [15:0]   int_reg_array_61_31_real;
  reg        [15:0]   int_reg_array_61_31_imag;
  reg        [15:0]   int_reg_array_61_32_real;
  reg        [15:0]   int_reg_array_61_32_imag;
  reg        [15:0]   int_reg_array_61_33_real;
  reg        [15:0]   int_reg_array_61_33_imag;
  reg        [15:0]   int_reg_array_61_34_real;
  reg        [15:0]   int_reg_array_61_34_imag;
  reg        [15:0]   int_reg_array_61_35_real;
  reg        [15:0]   int_reg_array_61_35_imag;
  reg        [15:0]   int_reg_array_61_36_real;
  reg        [15:0]   int_reg_array_61_36_imag;
  reg        [15:0]   int_reg_array_61_37_real;
  reg        [15:0]   int_reg_array_61_37_imag;
  reg        [15:0]   int_reg_array_61_38_real;
  reg        [15:0]   int_reg_array_61_38_imag;
  reg        [15:0]   int_reg_array_61_39_real;
  reg        [15:0]   int_reg_array_61_39_imag;
  reg        [15:0]   int_reg_array_61_40_real;
  reg        [15:0]   int_reg_array_61_40_imag;
  reg        [15:0]   int_reg_array_61_41_real;
  reg        [15:0]   int_reg_array_61_41_imag;
  reg        [15:0]   int_reg_array_61_42_real;
  reg        [15:0]   int_reg_array_61_42_imag;
  reg        [15:0]   int_reg_array_61_43_real;
  reg        [15:0]   int_reg_array_61_43_imag;
  reg        [15:0]   int_reg_array_61_44_real;
  reg        [15:0]   int_reg_array_61_44_imag;
  reg        [15:0]   int_reg_array_61_45_real;
  reg        [15:0]   int_reg_array_61_45_imag;
  reg        [15:0]   int_reg_array_61_46_real;
  reg        [15:0]   int_reg_array_61_46_imag;
  reg        [15:0]   int_reg_array_61_47_real;
  reg        [15:0]   int_reg_array_61_47_imag;
  reg        [15:0]   int_reg_array_61_48_real;
  reg        [15:0]   int_reg_array_61_48_imag;
  reg        [15:0]   int_reg_array_61_49_real;
  reg        [15:0]   int_reg_array_61_49_imag;
  reg        [15:0]   int_reg_array_61_50_real;
  reg        [15:0]   int_reg_array_61_50_imag;
  reg        [15:0]   int_reg_array_61_51_real;
  reg        [15:0]   int_reg_array_61_51_imag;
  reg        [15:0]   int_reg_array_61_52_real;
  reg        [15:0]   int_reg_array_61_52_imag;
  reg        [15:0]   int_reg_array_61_53_real;
  reg        [15:0]   int_reg_array_61_53_imag;
  reg        [15:0]   int_reg_array_61_54_real;
  reg        [15:0]   int_reg_array_61_54_imag;
  reg        [15:0]   int_reg_array_61_55_real;
  reg        [15:0]   int_reg_array_61_55_imag;
  reg        [15:0]   int_reg_array_61_56_real;
  reg        [15:0]   int_reg_array_61_56_imag;
  reg        [15:0]   int_reg_array_61_57_real;
  reg        [15:0]   int_reg_array_61_57_imag;
  reg        [15:0]   int_reg_array_61_58_real;
  reg        [15:0]   int_reg_array_61_58_imag;
  reg        [15:0]   int_reg_array_61_59_real;
  reg        [15:0]   int_reg_array_61_59_imag;
  reg        [15:0]   int_reg_array_61_60_real;
  reg        [15:0]   int_reg_array_61_60_imag;
  reg        [15:0]   int_reg_array_61_61_real;
  reg        [15:0]   int_reg_array_61_61_imag;
  reg        [15:0]   int_reg_array_61_62_real;
  reg        [15:0]   int_reg_array_61_62_imag;
  reg        [15:0]   int_reg_array_61_63_real;
  reg        [15:0]   int_reg_array_61_63_imag;
  reg        [15:0]   int_reg_array_28_0_real;
  reg        [15:0]   int_reg_array_28_0_imag;
  reg        [15:0]   int_reg_array_28_1_real;
  reg        [15:0]   int_reg_array_28_1_imag;
  reg        [15:0]   int_reg_array_28_2_real;
  reg        [15:0]   int_reg_array_28_2_imag;
  reg        [15:0]   int_reg_array_28_3_real;
  reg        [15:0]   int_reg_array_28_3_imag;
  reg        [15:0]   int_reg_array_28_4_real;
  reg        [15:0]   int_reg_array_28_4_imag;
  reg        [15:0]   int_reg_array_28_5_real;
  reg        [15:0]   int_reg_array_28_5_imag;
  reg        [15:0]   int_reg_array_28_6_real;
  reg        [15:0]   int_reg_array_28_6_imag;
  reg        [15:0]   int_reg_array_28_7_real;
  reg        [15:0]   int_reg_array_28_7_imag;
  reg        [15:0]   int_reg_array_28_8_real;
  reg        [15:0]   int_reg_array_28_8_imag;
  reg        [15:0]   int_reg_array_28_9_real;
  reg        [15:0]   int_reg_array_28_9_imag;
  reg        [15:0]   int_reg_array_28_10_real;
  reg        [15:0]   int_reg_array_28_10_imag;
  reg        [15:0]   int_reg_array_28_11_real;
  reg        [15:0]   int_reg_array_28_11_imag;
  reg        [15:0]   int_reg_array_28_12_real;
  reg        [15:0]   int_reg_array_28_12_imag;
  reg        [15:0]   int_reg_array_28_13_real;
  reg        [15:0]   int_reg_array_28_13_imag;
  reg        [15:0]   int_reg_array_28_14_real;
  reg        [15:0]   int_reg_array_28_14_imag;
  reg        [15:0]   int_reg_array_28_15_real;
  reg        [15:0]   int_reg_array_28_15_imag;
  reg        [15:0]   int_reg_array_28_16_real;
  reg        [15:0]   int_reg_array_28_16_imag;
  reg        [15:0]   int_reg_array_28_17_real;
  reg        [15:0]   int_reg_array_28_17_imag;
  reg        [15:0]   int_reg_array_28_18_real;
  reg        [15:0]   int_reg_array_28_18_imag;
  reg        [15:0]   int_reg_array_28_19_real;
  reg        [15:0]   int_reg_array_28_19_imag;
  reg        [15:0]   int_reg_array_28_20_real;
  reg        [15:0]   int_reg_array_28_20_imag;
  reg        [15:0]   int_reg_array_28_21_real;
  reg        [15:0]   int_reg_array_28_21_imag;
  reg        [15:0]   int_reg_array_28_22_real;
  reg        [15:0]   int_reg_array_28_22_imag;
  reg        [15:0]   int_reg_array_28_23_real;
  reg        [15:0]   int_reg_array_28_23_imag;
  reg        [15:0]   int_reg_array_28_24_real;
  reg        [15:0]   int_reg_array_28_24_imag;
  reg        [15:0]   int_reg_array_28_25_real;
  reg        [15:0]   int_reg_array_28_25_imag;
  reg        [15:0]   int_reg_array_28_26_real;
  reg        [15:0]   int_reg_array_28_26_imag;
  reg        [15:0]   int_reg_array_28_27_real;
  reg        [15:0]   int_reg_array_28_27_imag;
  reg        [15:0]   int_reg_array_28_28_real;
  reg        [15:0]   int_reg_array_28_28_imag;
  reg        [15:0]   int_reg_array_28_29_real;
  reg        [15:0]   int_reg_array_28_29_imag;
  reg        [15:0]   int_reg_array_28_30_real;
  reg        [15:0]   int_reg_array_28_30_imag;
  reg        [15:0]   int_reg_array_28_31_real;
  reg        [15:0]   int_reg_array_28_31_imag;
  reg        [15:0]   int_reg_array_28_32_real;
  reg        [15:0]   int_reg_array_28_32_imag;
  reg        [15:0]   int_reg_array_28_33_real;
  reg        [15:0]   int_reg_array_28_33_imag;
  reg        [15:0]   int_reg_array_28_34_real;
  reg        [15:0]   int_reg_array_28_34_imag;
  reg        [15:0]   int_reg_array_28_35_real;
  reg        [15:0]   int_reg_array_28_35_imag;
  reg        [15:0]   int_reg_array_28_36_real;
  reg        [15:0]   int_reg_array_28_36_imag;
  reg        [15:0]   int_reg_array_28_37_real;
  reg        [15:0]   int_reg_array_28_37_imag;
  reg        [15:0]   int_reg_array_28_38_real;
  reg        [15:0]   int_reg_array_28_38_imag;
  reg        [15:0]   int_reg_array_28_39_real;
  reg        [15:0]   int_reg_array_28_39_imag;
  reg        [15:0]   int_reg_array_28_40_real;
  reg        [15:0]   int_reg_array_28_40_imag;
  reg        [15:0]   int_reg_array_28_41_real;
  reg        [15:0]   int_reg_array_28_41_imag;
  reg        [15:0]   int_reg_array_28_42_real;
  reg        [15:0]   int_reg_array_28_42_imag;
  reg        [15:0]   int_reg_array_28_43_real;
  reg        [15:0]   int_reg_array_28_43_imag;
  reg        [15:0]   int_reg_array_28_44_real;
  reg        [15:0]   int_reg_array_28_44_imag;
  reg        [15:0]   int_reg_array_28_45_real;
  reg        [15:0]   int_reg_array_28_45_imag;
  reg        [15:0]   int_reg_array_28_46_real;
  reg        [15:0]   int_reg_array_28_46_imag;
  reg        [15:0]   int_reg_array_28_47_real;
  reg        [15:0]   int_reg_array_28_47_imag;
  reg        [15:0]   int_reg_array_28_48_real;
  reg        [15:0]   int_reg_array_28_48_imag;
  reg        [15:0]   int_reg_array_28_49_real;
  reg        [15:0]   int_reg_array_28_49_imag;
  reg        [15:0]   int_reg_array_28_50_real;
  reg        [15:0]   int_reg_array_28_50_imag;
  reg        [15:0]   int_reg_array_28_51_real;
  reg        [15:0]   int_reg_array_28_51_imag;
  reg        [15:0]   int_reg_array_28_52_real;
  reg        [15:0]   int_reg_array_28_52_imag;
  reg        [15:0]   int_reg_array_28_53_real;
  reg        [15:0]   int_reg_array_28_53_imag;
  reg        [15:0]   int_reg_array_28_54_real;
  reg        [15:0]   int_reg_array_28_54_imag;
  reg        [15:0]   int_reg_array_28_55_real;
  reg        [15:0]   int_reg_array_28_55_imag;
  reg        [15:0]   int_reg_array_28_56_real;
  reg        [15:0]   int_reg_array_28_56_imag;
  reg        [15:0]   int_reg_array_28_57_real;
  reg        [15:0]   int_reg_array_28_57_imag;
  reg        [15:0]   int_reg_array_28_58_real;
  reg        [15:0]   int_reg_array_28_58_imag;
  reg        [15:0]   int_reg_array_28_59_real;
  reg        [15:0]   int_reg_array_28_59_imag;
  reg        [15:0]   int_reg_array_28_60_real;
  reg        [15:0]   int_reg_array_28_60_imag;
  reg        [15:0]   int_reg_array_28_61_real;
  reg        [15:0]   int_reg_array_28_61_imag;
  reg        [15:0]   int_reg_array_28_62_real;
  reg        [15:0]   int_reg_array_28_62_imag;
  reg        [15:0]   int_reg_array_28_63_real;
  reg        [15:0]   int_reg_array_28_63_imag;
  reg        [15:0]   int_reg_array_51_0_real;
  reg        [15:0]   int_reg_array_51_0_imag;
  reg        [15:0]   int_reg_array_51_1_real;
  reg        [15:0]   int_reg_array_51_1_imag;
  reg        [15:0]   int_reg_array_51_2_real;
  reg        [15:0]   int_reg_array_51_2_imag;
  reg        [15:0]   int_reg_array_51_3_real;
  reg        [15:0]   int_reg_array_51_3_imag;
  reg        [15:0]   int_reg_array_51_4_real;
  reg        [15:0]   int_reg_array_51_4_imag;
  reg        [15:0]   int_reg_array_51_5_real;
  reg        [15:0]   int_reg_array_51_5_imag;
  reg        [15:0]   int_reg_array_51_6_real;
  reg        [15:0]   int_reg_array_51_6_imag;
  reg        [15:0]   int_reg_array_51_7_real;
  reg        [15:0]   int_reg_array_51_7_imag;
  reg        [15:0]   int_reg_array_51_8_real;
  reg        [15:0]   int_reg_array_51_8_imag;
  reg        [15:0]   int_reg_array_51_9_real;
  reg        [15:0]   int_reg_array_51_9_imag;
  reg        [15:0]   int_reg_array_51_10_real;
  reg        [15:0]   int_reg_array_51_10_imag;
  reg        [15:0]   int_reg_array_51_11_real;
  reg        [15:0]   int_reg_array_51_11_imag;
  reg        [15:0]   int_reg_array_51_12_real;
  reg        [15:0]   int_reg_array_51_12_imag;
  reg        [15:0]   int_reg_array_51_13_real;
  reg        [15:0]   int_reg_array_51_13_imag;
  reg        [15:0]   int_reg_array_51_14_real;
  reg        [15:0]   int_reg_array_51_14_imag;
  reg        [15:0]   int_reg_array_51_15_real;
  reg        [15:0]   int_reg_array_51_15_imag;
  reg        [15:0]   int_reg_array_51_16_real;
  reg        [15:0]   int_reg_array_51_16_imag;
  reg        [15:0]   int_reg_array_51_17_real;
  reg        [15:0]   int_reg_array_51_17_imag;
  reg        [15:0]   int_reg_array_51_18_real;
  reg        [15:0]   int_reg_array_51_18_imag;
  reg        [15:0]   int_reg_array_51_19_real;
  reg        [15:0]   int_reg_array_51_19_imag;
  reg        [15:0]   int_reg_array_51_20_real;
  reg        [15:0]   int_reg_array_51_20_imag;
  reg        [15:0]   int_reg_array_51_21_real;
  reg        [15:0]   int_reg_array_51_21_imag;
  reg        [15:0]   int_reg_array_51_22_real;
  reg        [15:0]   int_reg_array_51_22_imag;
  reg        [15:0]   int_reg_array_51_23_real;
  reg        [15:0]   int_reg_array_51_23_imag;
  reg        [15:0]   int_reg_array_51_24_real;
  reg        [15:0]   int_reg_array_51_24_imag;
  reg        [15:0]   int_reg_array_51_25_real;
  reg        [15:0]   int_reg_array_51_25_imag;
  reg        [15:0]   int_reg_array_51_26_real;
  reg        [15:0]   int_reg_array_51_26_imag;
  reg        [15:0]   int_reg_array_51_27_real;
  reg        [15:0]   int_reg_array_51_27_imag;
  reg        [15:0]   int_reg_array_51_28_real;
  reg        [15:0]   int_reg_array_51_28_imag;
  reg        [15:0]   int_reg_array_51_29_real;
  reg        [15:0]   int_reg_array_51_29_imag;
  reg        [15:0]   int_reg_array_51_30_real;
  reg        [15:0]   int_reg_array_51_30_imag;
  reg        [15:0]   int_reg_array_51_31_real;
  reg        [15:0]   int_reg_array_51_31_imag;
  reg        [15:0]   int_reg_array_51_32_real;
  reg        [15:0]   int_reg_array_51_32_imag;
  reg        [15:0]   int_reg_array_51_33_real;
  reg        [15:0]   int_reg_array_51_33_imag;
  reg        [15:0]   int_reg_array_51_34_real;
  reg        [15:0]   int_reg_array_51_34_imag;
  reg        [15:0]   int_reg_array_51_35_real;
  reg        [15:0]   int_reg_array_51_35_imag;
  reg        [15:0]   int_reg_array_51_36_real;
  reg        [15:0]   int_reg_array_51_36_imag;
  reg        [15:0]   int_reg_array_51_37_real;
  reg        [15:0]   int_reg_array_51_37_imag;
  reg        [15:0]   int_reg_array_51_38_real;
  reg        [15:0]   int_reg_array_51_38_imag;
  reg        [15:0]   int_reg_array_51_39_real;
  reg        [15:0]   int_reg_array_51_39_imag;
  reg        [15:0]   int_reg_array_51_40_real;
  reg        [15:0]   int_reg_array_51_40_imag;
  reg        [15:0]   int_reg_array_51_41_real;
  reg        [15:0]   int_reg_array_51_41_imag;
  reg        [15:0]   int_reg_array_51_42_real;
  reg        [15:0]   int_reg_array_51_42_imag;
  reg        [15:0]   int_reg_array_51_43_real;
  reg        [15:0]   int_reg_array_51_43_imag;
  reg        [15:0]   int_reg_array_51_44_real;
  reg        [15:0]   int_reg_array_51_44_imag;
  reg        [15:0]   int_reg_array_51_45_real;
  reg        [15:0]   int_reg_array_51_45_imag;
  reg        [15:0]   int_reg_array_51_46_real;
  reg        [15:0]   int_reg_array_51_46_imag;
  reg        [15:0]   int_reg_array_51_47_real;
  reg        [15:0]   int_reg_array_51_47_imag;
  reg        [15:0]   int_reg_array_51_48_real;
  reg        [15:0]   int_reg_array_51_48_imag;
  reg        [15:0]   int_reg_array_51_49_real;
  reg        [15:0]   int_reg_array_51_49_imag;
  reg        [15:0]   int_reg_array_51_50_real;
  reg        [15:0]   int_reg_array_51_50_imag;
  reg        [15:0]   int_reg_array_51_51_real;
  reg        [15:0]   int_reg_array_51_51_imag;
  reg        [15:0]   int_reg_array_51_52_real;
  reg        [15:0]   int_reg_array_51_52_imag;
  reg        [15:0]   int_reg_array_51_53_real;
  reg        [15:0]   int_reg_array_51_53_imag;
  reg        [15:0]   int_reg_array_51_54_real;
  reg        [15:0]   int_reg_array_51_54_imag;
  reg        [15:0]   int_reg_array_51_55_real;
  reg        [15:0]   int_reg_array_51_55_imag;
  reg        [15:0]   int_reg_array_51_56_real;
  reg        [15:0]   int_reg_array_51_56_imag;
  reg        [15:0]   int_reg_array_51_57_real;
  reg        [15:0]   int_reg_array_51_57_imag;
  reg        [15:0]   int_reg_array_51_58_real;
  reg        [15:0]   int_reg_array_51_58_imag;
  reg        [15:0]   int_reg_array_51_59_real;
  reg        [15:0]   int_reg_array_51_59_imag;
  reg        [15:0]   int_reg_array_51_60_real;
  reg        [15:0]   int_reg_array_51_60_imag;
  reg        [15:0]   int_reg_array_51_61_real;
  reg        [15:0]   int_reg_array_51_61_imag;
  reg        [15:0]   int_reg_array_51_62_real;
  reg        [15:0]   int_reg_array_51_62_imag;
  reg        [15:0]   int_reg_array_51_63_real;
  reg        [15:0]   int_reg_array_51_63_imag;
  reg        [15:0]   int_reg_array_63_0_real;
  reg        [15:0]   int_reg_array_63_0_imag;
  reg        [15:0]   int_reg_array_63_1_real;
  reg        [15:0]   int_reg_array_63_1_imag;
  reg        [15:0]   int_reg_array_63_2_real;
  reg        [15:0]   int_reg_array_63_2_imag;
  reg        [15:0]   int_reg_array_63_3_real;
  reg        [15:0]   int_reg_array_63_3_imag;
  reg        [15:0]   int_reg_array_63_4_real;
  reg        [15:0]   int_reg_array_63_4_imag;
  reg        [15:0]   int_reg_array_63_5_real;
  reg        [15:0]   int_reg_array_63_5_imag;
  reg        [15:0]   int_reg_array_63_6_real;
  reg        [15:0]   int_reg_array_63_6_imag;
  reg        [15:0]   int_reg_array_63_7_real;
  reg        [15:0]   int_reg_array_63_7_imag;
  reg        [15:0]   int_reg_array_63_8_real;
  reg        [15:0]   int_reg_array_63_8_imag;
  reg        [15:0]   int_reg_array_63_9_real;
  reg        [15:0]   int_reg_array_63_9_imag;
  reg        [15:0]   int_reg_array_63_10_real;
  reg        [15:0]   int_reg_array_63_10_imag;
  reg        [15:0]   int_reg_array_63_11_real;
  reg        [15:0]   int_reg_array_63_11_imag;
  reg        [15:0]   int_reg_array_63_12_real;
  reg        [15:0]   int_reg_array_63_12_imag;
  reg        [15:0]   int_reg_array_63_13_real;
  reg        [15:0]   int_reg_array_63_13_imag;
  reg        [15:0]   int_reg_array_63_14_real;
  reg        [15:0]   int_reg_array_63_14_imag;
  reg        [15:0]   int_reg_array_63_15_real;
  reg        [15:0]   int_reg_array_63_15_imag;
  reg        [15:0]   int_reg_array_63_16_real;
  reg        [15:0]   int_reg_array_63_16_imag;
  reg        [15:0]   int_reg_array_63_17_real;
  reg        [15:0]   int_reg_array_63_17_imag;
  reg        [15:0]   int_reg_array_63_18_real;
  reg        [15:0]   int_reg_array_63_18_imag;
  reg        [15:0]   int_reg_array_63_19_real;
  reg        [15:0]   int_reg_array_63_19_imag;
  reg        [15:0]   int_reg_array_63_20_real;
  reg        [15:0]   int_reg_array_63_20_imag;
  reg        [15:0]   int_reg_array_63_21_real;
  reg        [15:0]   int_reg_array_63_21_imag;
  reg        [15:0]   int_reg_array_63_22_real;
  reg        [15:0]   int_reg_array_63_22_imag;
  reg        [15:0]   int_reg_array_63_23_real;
  reg        [15:0]   int_reg_array_63_23_imag;
  reg        [15:0]   int_reg_array_63_24_real;
  reg        [15:0]   int_reg_array_63_24_imag;
  reg        [15:0]   int_reg_array_63_25_real;
  reg        [15:0]   int_reg_array_63_25_imag;
  reg        [15:0]   int_reg_array_63_26_real;
  reg        [15:0]   int_reg_array_63_26_imag;
  reg        [15:0]   int_reg_array_63_27_real;
  reg        [15:0]   int_reg_array_63_27_imag;
  reg        [15:0]   int_reg_array_63_28_real;
  reg        [15:0]   int_reg_array_63_28_imag;
  reg        [15:0]   int_reg_array_63_29_real;
  reg        [15:0]   int_reg_array_63_29_imag;
  reg        [15:0]   int_reg_array_63_30_real;
  reg        [15:0]   int_reg_array_63_30_imag;
  reg        [15:0]   int_reg_array_63_31_real;
  reg        [15:0]   int_reg_array_63_31_imag;
  reg        [15:0]   int_reg_array_63_32_real;
  reg        [15:0]   int_reg_array_63_32_imag;
  reg        [15:0]   int_reg_array_63_33_real;
  reg        [15:0]   int_reg_array_63_33_imag;
  reg        [15:0]   int_reg_array_63_34_real;
  reg        [15:0]   int_reg_array_63_34_imag;
  reg        [15:0]   int_reg_array_63_35_real;
  reg        [15:0]   int_reg_array_63_35_imag;
  reg        [15:0]   int_reg_array_63_36_real;
  reg        [15:0]   int_reg_array_63_36_imag;
  reg        [15:0]   int_reg_array_63_37_real;
  reg        [15:0]   int_reg_array_63_37_imag;
  reg        [15:0]   int_reg_array_63_38_real;
  reg        [15:0]   int_reg_array_63_38_imag;
  reg        [15:0]   int_reg_array_63_39_real;
  reg        [15:0]   int_reg_array_63_39_imag;
  reg        [15:0]   int_reg_array_63_40_real;
  reg        [15:0]   int_reg_array_63_40_imag;
  reg        [15:0]   int_reg_array_63_41_real;
  reg        [15:0]   int_reg_array_63_41_imag;
  reg        [15:0]   int_reg_array_63_42_real;
  reg        [15:0]   int_reg_array_63_42_imag;
  reg        [15:0]   int_reg_array_63_43_real;
  reg        [15:0]   int_reg_array_63_43_imag;
  reg        [15:0]   int_reg_array_63_44_real;
  reg        [15:0]   int_reg_array_63_44_imag;
  reg        [15:0]   int_reg_array_63_45_real;
  reg        [15:0]   int_reg_array_63_45_imag;
  reg        [15:0]   int_reg_array_63_46_real;
  reg        [15:0]   int_reg_array_63_46_imag;
  reg        [15:0]   int_reg_array_63_47_real;
  reg        [15:0]   int_reg_array_63_47_imag;
  reg        [15:0]   int_reg_array_63_48_real;
  reg        [15:0]   int_reg_array_63_48_imag;
  reg        [15:0]   int_reg_array_63_49_real;
  reg        [15:0]   int_reg_array_63_49_imag;
  reg        [15:0]   int_reg_array_63_50_real;
  reg        [15:0]   int_reg_array_63_50_imag;
  reg        [15:0]   int_reg_array_63_51_real;
  reg        [15:0]   int_reg_array_63_51_imag;
  reg        [15:0]   int_reg_array_63_52_real;
  reg        [15:0]   int_reg_array_63_52_imag;
  reg        [15:0]   int_reg_array_63_53_real;
  reg        [15:0]   int_reg_array_63_53_imag;
  reg        [15:0]   int_reg_array_63_54_real;
  reg        [15:0]   int_reg_array_63_54_imag;
  reg        [15:0]   int_reg_array_63_55_real;
  reg        [15:0]   int_reg_array_63_55_imag;
  reg        [15:0]   int_reg_array_63_56_real;
  reg        [15:0]   int_reg_array_63_56_imag;
  reg        [15:0]   int_reg_array_63_57_real;
  reg        [15:0]   int_reg_array_63_57_imag;
  reg        [15:0]   int_reg_array_63_58_real;
  reg        [15:0]   int_reg_array_63_58_imag;
  reg        [15:0]   int_reg_array_63_59_real;
  reg        [15:0]   int_reg_array_63_59_imag;
  reg        [15:0]   int_reg_array_63_60_real;
  reg        [15:0]   int_reg_array_63_60_imag;
  reg        [15:0]   int_reg_array_63_61_real;
  reg        [15:0]   int_reg_array_63_61_imag;
  reg        [15:0]   int_reg_array_63_62_real;
  reg        [15:0]   int_reg_array_63_62_imag;
  reg        [15:0]   int_reg_array_63_63_real;
  reg        [15:0]   int_reg_array_63_63_imag;
  reg        [15:0]   int_reg_array_17_0_real;
  reg        [15:0]   int_reg_array_17_0_imag;
  reg        [15:0]   int_reg_array_17_1_real;
  reg        [15:0]   int_reg_array_17_1_imag;
  reg        [15:0]   int_reg_array_17_2_real;
  reg        [15:0]   int_reg_array_17_2_imag;
  reg        [15:0]   int_reg_array_17_3_real;
  reg        [15:0]   int_reg_array_17_3_imag;
  reg        [15:0]   int_reg_array_17_4_real;
  reg        [15:0]   int_reg_array_17_4_imag;
  reg        [15:0]   int_reg_array_17_5_real;
  reg        [15:0]   int_reg_array_17_5_imag;
  reg        [15:0]   int_reg_array_17_6_real;
  reg        [15:0]   int_reg_array_17_6_imag;
  reg        [15:0]   int_reg_array_17_7_real;
  reg        [15:0]   int_reg_array_17_7_imag;
  reg        [15:0]   int_reg_array_17_8_real;
  reg        [15:0]   int_reg_array_17_8_imag;
  reg        [15:0]   int_reg_array_17_9_real;
  reg        [15:0]   int_reg_array_17_9_imag;
  reg        [15:0]   int_reg_array_17_10_real;
  reg        [15:0]   int_reg_array_17_10_imag;
  reg        [15:0]   int_reg_array_17_11_real;
  reg        [15:0]   int_reg_array_17_11_imag;
  reg        [15:0]   int_reg_array_17_12_real;
  reg        [15:0]   int_reg_array_17_12_imag;
  reg        [15:0]   int_reg_array_17_13_real;
  reg        [15:0]   int_reg_array_17_13_imag;
  reg        [15:0]   int_reg_array_17_14_real;
  reg        [15:0]   int_reg_array_17_14_imag;
  reg        [15:0]   int_reg_array_17_15_real;
  reg        [15:0]   int_reg_array_17_15_imag;
  reg        [15:0]   int_reg_array_17_16_real;
  reg        [15:0]   int_reg_array_17_16_imag;
  reg        [15:0]   int_reg_array_17_17_real;
  reg        [15:0]   int_reg_array_17_17_imag;
  reg        [15:0]   int_reg_array_17_18_real;
  reg        [15:0]   int_reg_array_17_18_imag;
  reg        [15:0]   int_reg_array_17_19_real;
  reg        [15:0]   int_reg_array_17_19_imag;
  reg        [15:0]   int_reg_array_17_20_real;
  reg        [15:0]   int_reg_array_17_20_imag;
  reg        [15:0]   int_reg_array_17_21_real;
  reg        [15:0]   int_reg_array_17_21_imag;
  reg        [15:0]   int_reg_array_17_22_real;
  reg        [15:0]   int_reg_array_17_22_imag;
  reg        [15:0]   int_reg_array_17_23_real;
  reg        [15:0]   int_reg_array_17_23_imag;
  reg        [15:0]   int_reg_array_17_24_real;
  reg        [15:0]   int_reg_array_17_24_imag;
  reg        [15:0]   int_reg_array_17_25_real;
  reg        [15:0]   int_reg_array_17_25_imag;
  reg        [15:0]   int_reg_array_17_26_real;
  reg        [15:0]   int_reg_array_17_26_imag;
  reg        [15:0]   int_reg_array_17_27_real;
  reg        [15:0]   int_reg_array_17_27_imag;
  reg        [15:0]   int_reg_array_17_28_real;
  reg        [15:0]   int_reg_array_17_28_imag;
  reg        [15:0]   int_reg_array_17_29_real;
  reg        [15:0]   int_reg_array_17_29_imag;
  reg        [15:0]   int_reg_array_17_30_real;
  reg        [15:0]   int_reg_array_17_30_imag;
  reg        [15:0]   int_reg_array_17_31_real;
  reg        [15:0]   int_reg_array_17_31_imag;
  reg        [15:0]   int_reg_array_17_32_real;
  reg        [15:0]   int_reg_array_17_32_imag;
  reg        [15:0]   int_reg_array_17_33_real;
  reg        [15:0]   int_reg_array_17_33_imag;
  reg        [15:0]   int_reg_array_17_34_real;
  reg        [15:0]   int_reg_array_17_34_imag;
  reg        [15:0]   int_reg_array_17_35_real;
  reg        [15:0]   int_reg_array_17_35_imag;
  reg        [15:0]   int_reg_array_17_36_real;
  reg        [15:0]   int_reg_array_17_36_imag;
  reg        [15:0]   int_reg_array_17_37_real;
  reg        [15:0]   int_reg_array_17_37_imag;
  reg        [15:0]   int_reg_array_17_38_real;
  reg        [15:0]   int_reg_array_17_38_imag;
  reg        [15:0]   int_reg_array_17_39_real;
  reg        [15:0]   int_reg_array_17_39_imag;
  reg        [15:0]   int_reg_array_17_40_real;
  reg        [15:0]   int_reg_array_17_40_imag;
  reg        [15:0]   int_reg_array_17_41_real;
  reg        [15:0]   int_reg_array_17_41_imag;
  reg        [15:0]   int_reg_array_17_42_real;
  reg        [15:0]   int_reg_array_17_42_imag;
  reg        [15:0]   int_reg_array_17_43_real;
  reg        [15:0]   int_reg_array_17_43_imag;
  reg        [15:0]   int_reg_array_17_44_real;
  reg        [15:0]   int_reg_array_17_44_imag;
  reg        [15:0]   int_reg_array_17_45_real;
  reg        [15:0]   int_reg_array_17_45_imag;
  reg        [15:0]   int_reg_array_17_46_real;
  reg        [15:0]   int_reg_array_17_46_imag;
  reg        [15:0]   int_reg_array_17_47_real;
  reg        [15:0]   int_reg_array_17_47_imag;
  reg        [15:0]   int_reg_array_17_48_real;
  reg        [15:0]   int_reg_array_17_48_imag;
  reg        [15:0]   int_reg_array_17_49_real;
  reg        [15:0]   int_reg_array_17_49_imag;
  reg        [15:0]   int_reg_array_17_50_real;
  reg        [15:0]   int_reg_array_17_50_imag;
  reg        [15:0]   int_reg_array_17_51_real;
  reg        [15:0]   int_reg_array_17_51_imag;
  reg        [15:0]   int_reg_array_17_52_real;
  reg        [15:0]   int_reg_array_17_52_imag;
  reg        [15:0]   int_reg_array_17_53_real;
  reg        [15:0]   int_reg_array_17_53_imag;
  reg        [15:0]   int_reg_array_17_54_real;
  reg        [15:0]   int_reg_array_17_54_imag;
  reg        [15:0]   int_reg_array_17_55_real;
  reg        [15:0]   int_reg_array_17_55_imag;
  reg        [15:0]   int_reg_array_17_56_real;
  reg        [15:0]   int_reg_array_17_56_imag;
  reg        [15:0]   int_reg_array_17_57_real;
  reg        [15:0]   int_reg_array_17_57_imag;
  reg        [15:0]   int_reg_array_17_58_real;
  reg        [15:0]   int_reg_array_17_58_imag;
  reg        [15:0]   int_reg_array_17_59_real;
  reg        [15:0]   int_reg_array_17_59_imag;
  reg        [15:0]   int_reg_array_17_60_real;
  reg        [15:0]   int_reg_array_17_60_imag;
  reg        [15:0]   int_reg_array_17_61_real;
  reg        [15:0]   int_reg_array_17_61_imag;
  reg        [15:0]   int_reg_array_17_62_real;
  reg        [15:0]   int_reg_array_17_62_imag;
  reg        [15:0]   int_reg_array_17_63_real;
  reg        [15:0]   int_reg_array_17_63_imag;
  reg        [15:0]   int_reg_array_12_0_real;
  reg        [15:0]   int_reg_array_12_0_imag;
  reg        [15:0]   int_reg_array_12_1_real;
  reg        [15:0]   int_reg_array_12_1_imag;
  reg        [15:0]   int_reg_array_12_2_real;
  reg        [15:0]   int_reg_array_12_2_imag;
  reg        [15:0]   int_reg_array_12_3_real;
  reg        [15:0]   int_reg_array_12_3_imag;
  reg        [15:0]   int_reg_array_12_4_real;
  reg        [15:0]   int_reg_array_12_4_imag;
  reg        [15:0]   int_reg_array_12_5_real;
  reg        [15:0]   int_reg_array_12_5_imag;
  reg        [15:0]   int_reg_array_12_6_real;
  reg        [15:0]   int_reg_array_12_6_imag;
  reg        [15:0]   int_reg_array_12_7_real;
  reg        [15:0]   int_reg_array_12_7_imag;
  reg        [15:0]   int_reg_array_12_8_real;
  reg        [15:0]   int_reg_array_12_8_imag;
  reg        [15:0]   int_reg_array_12_9_real;
  reg        [15:0]   int_reg_array_12_9_imag;
  reg        [15:0]   int_reg_array_12_10_real;
  reg        [15:0]   int_reg_array_12_10_imag;
  reg        [15:0]   int_reg_array_12_11_real;
  reg        [15:0]   int_reg_array_12_11_imag;
  reg        [15:0]   int_reg_array_12_12_real;
  reg        [15:0]   int_reg_array_12_12_imag;
  reg        [15:0]   int_reg_array_12_13_real;
  reg        [15:0]   int_reg_array_12_13_imag;
  reg        [15:0]   int_reg_array_12_14_real;
  reg        [15:0]   int_reg_array_12_14_imag;
  reg        [15:0]   int_reg_array_12_15_real;
  reg        [15:0]   int_reg_array_12_15_imag;
  reg        [15:0]   int_reg_array_12_16_real;
  reg        [15:0]   int_reg_array_12_16_imag;
  reg        [15:0]   int_reg_array_12_17_real;
  reg        [15:0]   int_reg_array_12_17_imag;
  reg        [15:0]   int_reg_array_12_18_real;
  reg        [15:0]   int_reg_array_12_18_imag;
  reg        [15:0]   int_reg_array_12_19_real;
  reg        [15:0]   int_reg_array_12_19_imag;
  reg        [15:0]   int_reg_array_12_20_real;
  reg        [15:0]   int_reg_array_12_20_imag;
  reg        [15:0]   int_reg_array_12_21_real;
  reg        [15:0]   int_reg_array_12_21_imag;
  reg        [15:0]   int_reg_array_12_22_real;
  reg        [15:0]   int_reg_array_12_22_imag;
  reg        [15:0]   int_reg_array_12_23_real;
  reg        [15:0]   int_reg_array_12_23_imag;
  reg        [15:0]   int_reg_array_12_24_real;
  reg        [15:0]   int_reg_array_12_24_imag;
  reg        [15:0]   int_reg_array_12_25_real;
  reg        [15:0]   int_reg_array_12_25_imag;
  reg        [15:0]   int_reg_array_12_26_real;
  reg        [15:0]   int_reg_array_12_26_imag;
  reg        [15:0]   int_reg_array_12_27_real;
  reg        [15:0]   int_reg_array_12_27_imag;
  reg        [15:0]   int_reg_array_12_28_real;
  reg        [15:0]   int_reg_array_12_28_imag;
  reg        [15:0]   int_reg_array_12_29_real;
  reg        [15:0]   int_reg_array_12_29_imag;
  reg        [15:0]   int_reg_array_12_30_real;
  reg        [15:0]   int_reg_array_12_30_imag;
  reg        [15:0]   int_reg_array_12_31_real;
  reg        [15:0]   int_reg_array_12_31_imag;
  reg        [15:0]   int_reg_array_12_32_real;
  reg        [15:0]   int_reg_array_12_32_imag;
  reg        [15:0]   int_reg_array_12_33_real;
  reg        [15:0]   int_reg_array_12_33_imag;
  reg        [15:0]   int_reg_array_12_34_real;
  reg        [15:0]   int_reg_array_12_34_imag;
  reg        [15:0]   int_reg_array_12_35_real;
  reg        [15:0]   int_reg_array_12_35_imag;
  reg        [15:0]   int_reg_array_12_36_real;
  reg        [15:0]   int_reg_array_12_36_imag;
  reg        [15:0]   int_reg_array_12_37_real;
  reg        [15:0]   int_reg_array_12_37_imag;
  reg        [15:0]   int_reg_array_12_38_real;
  reg        [15:0]   int_reg_array_12_38_imag;
  reg        [15:0]   int_reg_array_12_39_real;
  reg        [15:0]   int_reg_array_12_39_imag;
  reg        [15:0]   int_reg_array_12_40_real;
  reg        [15:0]   int_reg_array_12_40_imag;
  reg        [15:0]   int_reg_array_12_41_real;
  reg        [15:0]   int_reg_array_12_41_imag;
  reg        [15:0]   int_reg_array_12_42_real;
  reg        [15:0]   int_reg_array_12_42_imag;
  reg        [15:0]   int_reg_array_12_43_real;
  reg        [15:0]   int_reg_array_12_43_imag;
  reg        [15:0]   int_reg_array_12_44_real;
  reg        [15:0]   int_reg_array_12_44_imag;
  reg        [15:0]   int_reg_array_12_45_real;
  reg        [15:0]   int_reg_array_12_45_imag;
  reg        [15:0]   int_reg_array_12_46_real;
  reg        [15:0]   int_reg_array_12_46_imag;
  reg        [15:0]   int_reg_array_12_47_real;
  reg        [15:0]   int_reg_array_12_47_imag;
  reg        [15:0]   int_reg_array_12_48_real;
  reg        [15:0]   int_reg_array_12_48_imag;
  reg        [15:0]   int_reg_array_12_49_real;
  reg        [15:0]   int_reg_array_12_49_imag;
  reg        [15:0]   int_reg_array_12_50_real;
  reg        [15:0]   int_reg_array_12_50_imag;
  reg        [15:0]   int_reg_array_12_51_real;
  reg        [15:0]   int_reg_array_12_51_imag;
  reg        [15:0]   int_reg_array_12_52_real;
  reg        [15:0]   int_reg_array_12_52_imag;
  reg        [15:0]   int_reg_array_12_53_real;
  reg        [15:0]   int_reg_array_12_53_imag;
  reg        [15:0]   int_reg_array_12_54_real;
  reg        [15:0]   int_reg_array_12_54_imag;
  reg        [15:0]   int_reg_array_12_55_real;
  reg        [15:0]   int_reg_array_12_55_imag;
  reg        [15:0]   int_reg_array_12_56_real;
  reg        [15:0]   int_reg_array_12_56_imag;
  reg        [15:0]   int_reg_array_12_57_real;
  reg        [15:0]   int_reg_array_12_57_imag;
  reg        [15:0]   int_reg_array_12_58_real;
  reg        [15:0]   int_reg_array_12_58_imag;
  reg        [15:0]   int_reg_array_12_59_real;
  reg        [15:0]   int_reg_array_12_59_imag;
  reg        [15:0]   int_reg_array_12_60_real;
  reg        [15:0]   int_reg_array_12_60_imag;
  reg        [15:0]   int_reg_array_12_61_real;
  reg        [15:0]   int_reg_array_12_61_imag;
  reg        [15:0]   int_reg_array_12_62_real;
  reg        [15:0]   int_reg_array_12_62_imag;
  reg        [15:0]   int_reg_array_12_63_real;
  reg        [15:0]   int_reg_array_12_63_imag;
  reg        [15:0]   int_reg_array_52_0_real;
  reg        [15:0]   int_reg_array_52_0_imag;
  reg        [15:0]   int_reg_array_52_1_real;
  reg        [15:0]   int_reg_array_52_1_imag;
  reg        [15:0]   int_reg_array_52_2_real;
  reg        [15:0]   int_reg_array_52_2_imag;
  reg        [15:0]   int_reg_array_52_3_real;
  reg        [15:0]   int_reg_array_52_3_imag;
  reg        [15:0]   int_reg_array_52_4_real;
  reg        [15:0]   int_reg_array_52_4_imag;
  reg        [15:0]   int_reg_array_52_5_real;
  reg        [15:0]   int_reg_array_52_5_imag;
  reg        [15:0]   int_reg_array_52_6_real;
  reg        [15:0]   int_reg_array_52_6_imag;
  reg        [15:0]   int_reg_array_52_7_real;
  reg        [15:0]   int_reg_array_52_7_imag;
  reg        [15:0]   int_reg_array_52_8_real;
  reg        [15:0]   int_reg_array_52_8_imag;
  reg        [15:0]   int_reg_array_52_9_real;
  reg        [15:0]   int_reg_array_52_9_imag;
  reg        [15:0]   int_reg_array_52_10_real;
  reg        [15:0]   int_reg_array_52_10_imag;
  reg        [15:0]   int_reg_array_52_11_real;
  reg        [15:0]   int_reg_array_52_11_imag;
  reg        [15:0]   int_reg_array_52_12_real;
  reg        [15:0]   int_reg_array_52_12_imag;
  reg        [15:0]   int_reg_array_52_13_real;
  reg        [15:0]   int_reg_array_52_13_imag;
  reg        [15:0]   int_reg_array_52_14_real;
  reg        [15:0]   int_reg_array_52_14_imag;
  reg        [15:0]   int_reg_array_52_15_real;
  reg        [15:0]   int_reg_array_52_15_imag;
  reg        [15:0]   int_reg_array_52_16_real;
  reg        [15:0]   int_reg_array_52_16_imag;
  reg        [15:0]   int_reg_array_52_17_real;
  reg        [15:0]   int_reg_array_52_17_imag;
  reg        [15:0]   int_reg_array_52_18_real;
  reg        [15:0]   int_reg_array_52_18_imag;
  reg        [15:0]   int_reg_array_52_19_real;
  reg        [15:0]   int_reg_array_52_19_imag;
  reg        [15:0]   int_reg_array_52_20_real;
  reg        [15:0]   int_reg_array_52_20_imag;
  reg        [15:0]   int_reg_array_52_21_real;
  reg        [15:0]   int_reg_array_52_21_imag;
  reg        [15:0]   int_reg_array_52_22_real;
  reg        [15:0]   int_reg_array_52_22_imag;
  reg        [15:0]   int_reg_array_52_23_real;
  reg        [15:0]   int_reg_array_52_23_imag;
  reg        [15:0]   int_reg_array_52_24_real;
  reg        [15:0]   int_reg_array_52_24_imag;
  reg        [15:0]   int_reg_array_52_25_real;
  reg        [15:0]   int_reg_array_52_25_imag;
  reg        [15:0]   int_reg_array_52_26_real;
  reg        [15:0]   int_reg_array_52_26_imag;
  reg        [15:0]   int_reg_array_52_27_real;
  reg        [15:0]   int_reg_array_52_27_imag;
  reg        [15:0]   int_reg_array_52_28_real;
  reg        [15:0]   int_reg_array_52_28_imag;
  reg        [15:0]   int_reg_array_52_29_real;
  reg        [15:0]   int_reg_array_52_29_imag;
  reg        [15:0]   int_reg_array_52_30_real;
  reg        [15:0]   int_reg_array_52_30_imag;
  reg        [15:0]   int_reg_array_52_31_real;
  reg        [15:0]   int_reg_array_52_31_imag;
  reg        [15:0]   int_reg_array_52_32_real;
  reg        [15:0]   int_reg_array_52_32_imag;
  reg        [15:0]   int_reg_array_52_33_real;
  reg        [15:0]   int_reg_array_52_33_imag;
  reg        [15:0]   int_reg_array_52_34_real;
  reg        [15:0]   int_reg_array_52_34_imag;
  reg        [15:0]   int_reg_array_52_35_real;
  reg        [15:0]   int_reg_array_52_35_imag;
  reg        [15:0]   int_reg_array_52_36_real;
  reg        [15:0]   int_reg_array_52_36_imag;
  reg        [15:0]   int_reg_array_52_37_real;
  reg        [15:0]   int_reg_array_52_37_imag;
  reg        [15:0]   int_reg_array_52_38_real;
  reg        [15:0]   int_reg_array_52_38_imag;
  reg        [15:0]   int_reg_array_52_39_real;
  reg        [15:0]   int_reg_array_52_39_imag;
  reg        [15:0]   int_reg_array_52_40_real;
  reg        [15:0]   int_reg_array_52_40_imag;
  reg        [15:0]   int_reg_array_52_41_real;
  reg        [15:0]   int_reg_array_52_41_imag;
  reg        [15:0]   int_reg_array_52_42_real;
  reg        [15:0]   int_reg_array_52_42_imag;
  reg        [15:0]   int_reg_array_52_43_real;
  reg        [15:0]   int_reg_array_52_43_imag;
  reg        [15:0]   int_reg_array_52_44_real;
  reg        [15:0]   int_reg_array_52_44_imag;
  reg        [15:0]   int_reg_array_52_45_real;
  reg        [15:0]   int_reg_array_52_45_imag;
  reg        [15:0]   int_reg_array_52_46_real;
  reg        [15:0]   int_reg_array_52_46_imag;
  reg        [15:0]   int_reg_array_52_47_real;
  reg        [15:0]   int_reg_array_52_47_imag;
  reg        [15:0]   int_reg_array_52_48_real;
  reg        [15:0]   int_reg_array_52_48_imag;
  reg        [15:0]   int_reg_array_52_49_real;
  reg        [15:0]   int_reg_array_52_49_imag;
  reg        [15:0]   int_reg_array_52_50_real;
  reg        [15:0]   int_reg_array_52_50_imag;
  reg        [15:0]   int_reg_array_52_51_real;
  reg        [15:0]   int_reg_array_52_51_imag;
  reg        [15:0]   int_reg_array_52_52_real;
  reg        [15:0]   int_reg_array_52_52_imag;
  reg        [15:0]   int_reg_array_52_53_real;
  reg        [15:0]   int_reg_array_52_53_imag;
  reg        [15:0]   int_reg_array_52_54_real;
  reg        [15:0]   int_reg_array_52_54_imag;
  reg        [15:0]   int_reg_array_52_55_real;
  reg        [15:0]   int_reg_array_52_55_imag;
  reg        [15:0]   int_reg_array_52_56_real;
  reg        [15:0]   int_reg_array_52_56_imag;
  reg        [15:0]   int_reg_array_52_57_real;
  reg        [15:0]   int_reg_array_52_57_imag;
  reg        [15:0]   int_reg_array_52_58_real;
  reg        [15:0]   int_reg_array_52_58_imag;
  reg        [15:0]   int_reg_array_52_59_real;
  reg        [15:0]   int_reg_array_52_59_imag;
  reg        [15:0]   int_reg_array_52_60_real;
  reg        [15:0]   int_reg_array_52_60_imag;
  reg        [15:0]   int_reg_array_52_61_real;
  reg        [15:0]   int_reg_array_52_61_imag;
  reg        [15:0]   int_reg_array_52_62_real;
  reg        [15:0]   int_reg_array_52_62_imag;
  reg        [15:0]   int_reg_array_52_63_real;
  reg        [15:0]   int_reg_array_52_63_imag;
  reg        [15:0]   int_reg_array_11_0_real;
  reg        [15:0]   int_reg_array_11_0_imag;
  reg        [15:0]   int_reg_array_11_1_real;
  reg        [15:0]   int_reg_array_11_1_imag;
  reg        [15:0]   int_reg_array_11_2_real;
  reg        [15:0]   int_reg_array_11_2_imag;
  reg        [15:0]   int_reg_array_11_3_real;
  reg        [15:0]   int_reg_array_11_3_imag;
  reg        [15:0]   int_reg_array_11_4_real;
  reg        [15:0]   int_reg_array_11_4_imag;
  reg        [15:0]   int_reg_array_11_5_real;
  reg        [15:0]   int_reg_array_11_5_imag;
  reg        [15:0]   int_reg_array_11_6_real;
  reg        [15:0]   int_reg_array_11_6_imag;
  reg        [15:0]   int_reg_array_11_7_real;
  reg        [15:0]   int_reg_array_11_7_imag;
  reg        [15:0]   int_reg_array_11_8_real;
  reg        [15:0]   int_reg_array_11_8_imag;
  reg        [15:0]   int_reg_array_11_9_real;
  reg        [15:0]   int_reg_array_11_9_imag;
  reg        [15:0]   int_reg_array_11_10_real;
  reg        [15:0]   int_reg_array_11_10_imag;
  reg        [15:0]   int_reg_array_11_11_real;
  reg        [15:0]   int_reg_array_11_11_imag;
  reg        [15:0]   int_reg_array_11_12_real;
  reg        [15:0]   int_reg_array_11_12_imag;
  reg        [15:0]   int_reg_array_11_13_real;
  reg        [15:0]   int_reg_array_11_13_imag;
  reg        [15:0]   int_reg_array_11_14_real;
  reg        [15:0]   int_reg_array_11_14_imag;
  reg        [15:0]   int_reg_array_11_15_real;
  reg        [15:0]   int_reg_array_11_15_imag;
  reg        [15:0]   int_reg_array_11_16_real;
  reg        [15:0]   int_reg_array_11_16_imag;
  reg        [15:0]   int_reg_array_11_17_real;
  reg        [15:0]   int_reg_array_11_17_imag;
  reg        [15:0]   int_reg_array_11_18_real;
  reg        [15:0]   int_reg_array_11_18_imag;
  reg        [15:0]   int_reg_array_11_19_real;
  reg        [15:0]   int_reg_array_11_19_imag;
  reg        [15:0]   int_reg_array_11_20_real;
  reg        [15:0]   int_reg_array_11_20_imag;
  reg        [15:0]   int_reg_array_11_21_real;
  reg        [15:0]   int_reg_array_11_21_imag;
  reg        [15:0]   int_reg_array_11_22_real;
  reg        [15:0]   int_reg_array_11_22_imag;
  reg        [15:0]   int_reg_array_11_23_real;
  reg        [15:0]   int_reg_array_11_23_imag;
  reg        [15:0]   int_reg_array_11_24_real;
  reg        [15:0]   int_reg_array_11_24_imag;
  reg        [15:0]   int_reg_array_11_25_real;
  reg        [15:0]   int_reg_array_11_25_imag;
  reg        [15:0]   int_reg_array_11_26_real;
  reg        [15:0]   int_reg_array_11_26_imag;
  reg        [15:0]   int_reg_array_11_27_real;
  reg        [15:0]   int_reg_array_11_27_imag;
  reg        [15:0]   int_reg_array_11_28_real;
  reg        [15:0]   int_reg_array_11_28_imag;
  reg        [15:0]   int_reg_array_11_29_real;
  reg        [15:0]   int_reg_array_11_29_imag;
  reg        [15:0]   int_reg_array_11_30_real;
  reg        [15:0]   int_reg_array_11_30_imag;
  reg        [15:0]   int_reg_array_11_31_real;
  reg        [15:0]   int_reg_array_11_31_imag;
  reg        [15:0]   int_reg_array_11_32_real;
  reg        [15:0]   int_reg_array_11_32_imag;
  reg        [15:0]   int_reg_array_11_33_real;
  reg        [15:0]   int_reg_array_11_33_imag;
  reg        [15:0]   int_reg_array_11_34_real;
  reg        [15:0]   int_reg_array_11_34_imag;
  reg        [15:0]   int_reg_array_11_35_real;
  reg        [15:0]   int_reg_array_11_35_imag;
  reg        [15:0]   int_reg_array_11_36_real;
  reg        [15:0]   int_reg_array_11_36_imag;
  reg        [15:0]   int_reg_array_11_37_real;
  reg        [15:0]   int_reg_array_11_37_imag;
  reg        [15:0]   int_reg_array_11_38_real;
  reg        [15:0]   int_reg_array_11_38_imag;
  reg        [15:0]   int_reg_array_11_39_real;
  reg        [15:0]   int_reg_array_11_39_imag;
  reg        [15:0]   int_reg_array_11_40_real;
  reg        [15:0]   int_reg_array_11_40_imag;
  reg        [15:0]   int_reg_array_11_41_real;
  reg        [15:0]   int_reg_array_11_41_imag;
  reg        [15:0]   int_reg_array_11_42_real;
  reg        [15:0]   int_reg_array_11_42_imag;
  reg        [15:0]   int_reg_array_11_43_real;
  reg        [15:0]   int_reg_array_11_43_imag;
  reg        [15:0]   int_reg_array_11_44_real;
  reg        [15:0]   int_reg_array_11_44_imag;
  reg        [15:0]   int_reg_array_11_45_real;
  reg        [15:0]   int_reg_array_11_45_imag;
  reg        [15:0]   int_reg_array_11_46_real;
  reg        [15:0]   int_reg_array_11_46_imag;
  reg        [15:0]   int_reg_array_11_47_real;
  reg        [15:0]   int_reg_array_11_47_imag;
  reg        [15:0]   int_reg_array_11_48_real;
  reg        [15:0]   int_reg_array_11_48_imag;
  reg        [15:0]   int_reg_array_11_49_real;
  reg        [15:0]   int_reg_array_11_49_imag;
  reg        [15:0]   int_reg_array_11_50_real;
  reg        [15:0]   int_reg_array_11_50_imag;
  reg        [15:0]   int_reg_array_11_51_real;
  reg        [15:0]   int_reg_array_11_51_imag;
  reg        [15:0]   int_reg_array_11_52_real;
  reg        [15:0]   int_reg_array_11_52_imag;
  reg        [15:0]   int_reg_array_11_53_real;
  reg        [15:0]   int_reg_array_11_53_imag;
  reg        [15:0]   int_reg_array_11_54_real;
  reg        [15:0]   int_reg_array_11_54_imag;
  reg        [15:0]   int_reg_array_11_55_real;
  reg        [15:0]   int_reg_array_11_55_imag;
  reg        [15:0]   int_reg_array_11_56_real;
  reg        [15:0]   int_reg_array_11_56_imag;
  reg        [15:0]   int_reg_array_11_57_real;
  reg        [15:0]   int_reg_array_11_57_imag;
  reg        [15:0]   int_reg_array_11_58_real;
  reg        [15:0]   int_reg_array_11_58_imag;
  reg        [15:0]   int_reg_array_11_59_real;
  reg        [15:0]   int_reg_array_11_59_imag;
  reg        [15:0]   int_reg_array_11_60_real;
  reg        [15:0]   int_reg_array_11_60_imag;
  reg        [15:0]   int_reg_array_11_61_real;
  reg        [15:0]   int_reg_array_11_61_imag;
  reg        [15:0]   int_reg_array_11_62_real;
  reg        [15:0]   int_reg_array_11_62_imag;
  reg        [15:0]   int_reg_array_11_63_real;
  reg        [15:0]   int_reg_array_11_63_imag;
  reg        [15:0]   int_reg_array_5_0_real;
  reg        [15:0]   int_reg_array_5_0_imag;
  reg        [15:0]   int_reg_array_5_1_real;
  reg        [15:0]   int_reg_array_5_1_imag;
  reg        [15:0]   int_reg_array_5_2_real;
  reg        [15:0]   int_reg_array_5_2_imag;
  reg        [15:0]   int_reg_array_5_3_real;
  reg        [15:0]   int_reg_array_5_3_imag;
  reg        [15:0]   int_reg_array_5_4_real;
  reg        [15:0]   int_reg_array_5_4_imag;
  reg        [15:0]   int_reg_array_5_5_real;
  reg        [15:0]   int_reg_array_5_5_imag;
  reg        [15:0]   int_reg_array_5_6_real;
  reg        [15:0]   int_reg_array_5_6_imag;
  reg        [15:0]   int_reg_array_5_7_real;
  reg        [15:0]   int_reg_array_5_7_imag;
  reg        [15:0]   int_reg_array_5_8_real;
  reg        [15:0]   int_reg_array_5_8_imag;
  reg        [15:0]   int_reg_array_5_9_real;
  reg        [15:0]   int_reg_array_5_9_imag;
  reg        [15:0]   int_reg_array_5_10_real;
  reg        [15:0]   int_reg_array_5_10_imag;
  reg        [15:0]   int_reg_array_5_11_real;
  reg        [15:0]   int_reg_array_5_11_imag;
  reg        [15:0]   int_reg_array_5_12_real;
  reg        [15:0]   int_reg_array_5_12_imag;
  reg        [15:0]   int_reg_array_5_13_real;
  reg        [15:0]   int_reg_array_5_13_imag;
  reg        [15:0]   int_reg_array_5_14_real;
  reg        [15:0]   int_reg_array_5_14_imag;
  reg        [15:0]   int_reg_array_5_15_real;
  reg        [15:0]   int_reg_array_5_15_imag;
  reg        [15:0]   int_reg_array_5_16_real;
  reg        [15:0]   int_reg_array_5_16_imag;
  reg        [15:0]   int_reg_array_5_17_real;
  reg        [15:0]   int_reg_array_5_17_imag;
  reg        [15:0]   int_reg_array_5_18_real;
  reg        [15:0]   int_reg_array_5_18_imag;
  reg        [15:0]   int_reg_array_5_19_real;
  reg        [15:0]   int_reg_array_5_19_imag;
  reg        [15:0]   int_reg_array_5_20_real;
  reg        [15:0]   int_reg_array_5_20_imag;
  reg        [15:0]   int_reg_array_5_21_real;
  reg        [15:0]   int_reg_array_5_21_imag;
  reg        [15:0]   int_reg_array_5_22_real;
  reg        [15:0]   int_reg_array_5_22_imag;
  reg        [15:0]   int_reg_array_5_23_real;
  reg        [15:0]   int_reg_array_5_23_imag;
  reg        [15:0]   int_reg_array_5_24_real;
  reg        [15:0]   int_reg_array_5_24_imag;
  reg        [15:0]   int_reg_array_5_25_real;
  reg        [15:0]   int_reg_array_5_25_imag;
  reg        [15:0]   int_reg_array_5_26_real;
  reg        [15:0]   int_reg_array_5_26_imag;
  reg        [15:0]   int_reg_array_5_27_real;
  reg        [15:0]   int_reg_array_5_27_imag;
  reg        [15:0]   int_reg_array_5_28_real;
  reg        [15:0]   int_reg_array_5_28_imag;
  reg        [15:0]   int_reg_array_5_29_real;
  reg        [15:0]   int_reg_array_5_29_imag;
  reg        [15:0]   int_reg_array_5_30_real;
  reg        [15:0]   int_reg_array_5_30_imag;
  reg        [15:0]   int_reg_array_5_31_real;
  reg        [15:0]   int_reg_array_5_31_imag;
  reg        [15:0]   int_reg_array_5_32_real;
  reg        [15:0]   int_reg_array_5_32_imag;
  reg        [15:0]   int_reg_array_5_33_real;
  reg        [15:0]   int_reg_array_5_33_imag;
  reg        [15:0]   int_reg_array_5_34_real;
  reg        [15:0]   int_reg_array_5_34_imag;
  reg        [15:0]   int_reg_array_5_35_real;
  reg        [15:0]   int_reg_array_5_35_imag;
  reg        [15:0]   int_reg_array_5_36_real;
  reg        [15:0]   int_reg_array_5_36_imag;
  reg        [15:0]   int_reg_array_5_37_real;
  reg        [15:0]   int_reg_array_5_37_imag;
  reg        [15:0]   int_reg_array_5_38_real;
  reg        [15:0]   int_reg_array_5_38_imag;
  reg        [15:0]   int_reg_array_5_39_real;
  reg        [15:0]   int_reg_array_5_39_imag;
  reg        [15:0]   int_reg_array_5_40_real;
  reg        [15:0]   int_reg_array_5_40_imag;
  reg        [15:0]   int_reg_array_5_41_real;
  reg        [15:0]   int_reg_array_5_41_imag;
  reg        [15:0]   int_reg_array_5_42_real;
  reg        [15:0]   int_reg_array_5_42_imag;
  reg        [15:0]   int_reg_array_5_43_real;
  reg        [15:0]   int_reg_array_5_43_imag;
  reg        [15:0]   int_reg_array_5_44_real;
  reg        [15:0]   int_reg_array_5_44_imag;
  reg        [15:0]   int_reg_array_5_45_real;
  reg        [15:0]   int_reg_array_5_45_imag;
  reg        [15:0]   int_reg_array_5_46_real;
  reg        [15:0]   int_reg_array_5_46_imag;
  reg        [15:0]   int_reg_array_5_47_real;
  reg        [15:0]   int_reg_array_5_47_imag;
  reg        [15:0]   int_reg_array_5_48_real;
  reg        [15:0]   int_reg_array_5_48_imag;
  reg        [15:0]   int_reg_array_5_49_real;
  reg        [15:0]   int_reg_array_5_49_imag;
  reg        [15:0]   int_reg_array_5_50_real;
  reg        [15:0]   int_reg_array_5_50_imag;
  reg        [15:0]   int_reg_array_5_51_real;
  reg        [15:0]   int_reg_array_5_51_imag;
  reg        [15:0]   int_reg_array_5_52_real;
  reg        [15:0]   int_reg_array_5_52_imag;
  reg        [15:0]   int_reg_array_5_53_real;
  reg        [15:0]   int_reg_array_5_53_imag;
  reg        [15:0]   int_reg_array_5_54_real;
  reg        [15:0]   int_reg_array_5_54_imag;
  reg        [15:0]   int_reg_array_5_55_real;
  reg        [15:0]   int_reg_array_5_55_imag;
  reg        [15:0]   int_reg_array_5_56_real;
  reg        [15:0]   int_reg_array_5_56_imag;
  reg        [15:0]   int_reg_array_5_57_real;
  reg        [15:0]   int_reg_array_5_57_imag;
  reg        [15:0]   int_reg_array_5_58_real;
  reg        [15:0]   int_reg_array_5_58_imag;
  reg        [15:0]   int_reg_array_5_59_real;
  reg        [15:0]   int_reg_array_5_59_imag;
  reg        [15:0]   int_reg_array_5_60_real;
  reg        [15:0]   int_reg_array_5_60_imag;
  reg        [15:0]   int_reg_array_5_61_real;
  reg        [15:0]   int_reg_array_5_61_imag;
  reg        [15:0]   int_reg_array_5_62_real;
  reg        [15:0]   int_reg_array_5_62_imag;
  reg        [15:0]   int_reg_array_5_63_real;
  reg        [15:0]   int_reg_array_5_63_imag;
  reg        [15:0]   int_reg_array_32_0_real;
  reg        [15:0]   int_reg_array_32_0_imag;
  reg        [15:0]   int_reg_array_32_1_real;
  reg        [15:0]   int_reg_array_32_1_imag;
  reg        [15:0]   int_reg_array_32_2_real;
  reg        [15:0]   int_reg_array_32_2_imag;
  reg        [15:0]   int_reg_array_32_3_real;
  reg        [15:0]   int_reg_array_32_3_imag;
  reg        [15:0]   int_reg_array_32_4_real;
  reg        [15:0]   int_reg_array_32_4_imag;
  reg        [15:0]   int_reg_array_32_5_real;
  reg        [15:0]   int_reg_array_32_5_imag;
  reg        [15:0]   int_reg_array_32_6_real;
  reg        [15:0]   int_reg_array_32_6_imag;
  reg        [15:0]   int_reg_array_32_7_real;
  reg        [15:0]   int_reg_array_32_7_imag;
  reg        [15:0]   int_reg_array_32_8_real;
  reg        [15:0]   int_reg_array_32_8_imag;
  reg        [15:0]   int_reg_array_32_9_real;
  reg        [15:0]   int_reg_array_32_9_imag;
  reg        [15:0]   int_reg_array_32_10_real;
  reg        [15:0]   int_reg_array_32_10_imag;
  reg        [15:0]   int_reg_array_32_11_real;
  reg        [15:0]   int_reg_array_32_11_imag;
  reg        [15:0]   int_reg_array_32_12_real;
  reg        [15:0]   int_reg_array_32_12_imag;
  reg        [15:0]   int_reg_array_32_13_real;
  reg        [15:0]   int_reg_array_32_13_imag;
  reg        [15:0]   int_reg_array_32_14_real;
  reg        [15:0]   int_reg_array_32_14_imag;
  reg        [15:0]   int_reg_array_32_15_real;
  reg        [15:0]   int_reg_array_32_15_imag;
  reg        [15:0]   int_reg_array_32_16_real;
  reg        [15:0]   int_reg_array_32_16_imag;
  reg        [15:0]   int_reg_array_32_17_real;
  reg        [15:0]   int_reg_array_32_17_imag;
  reg        [15:0]   int_reg_array_32_18_real;
  reg        [15:0]   int_reg_array_32_18_imag;
  reg        [15:0]   int_reg_array_32_19_real;
  reg        [15:0]   int_reg_array_32_19_imag;
  reg        [15:0]   int_reg_array_32_20_real;
  reg        [15:0]   int_reg_array_32_20_imag;
  reg        [15:0]   int_reg_array_32_21_real;
  reg        [15:0]   int_reg_array_32_21_imag;
  reg        [15:0]   int_reg_array_32_22_real;
  reg        [15:0]   int_reg_array_32_22_imag;
  reg        [15:0]   int_reg_array_32_23_real;
  reg        [15:0]   int_reg_array_32_23_imag;
  reg        [15:0]   int_reg_array_32_24_real;
  reg        [15:0]   int_reg_array_32_24_imag;
  reg        [15:0]   int_reg_array_32_25_real;
  reg        [15:0]   int_reg_array_32_25_imag;
  reg        [15:0]   int_reg_array_32_26_real;
  reg        [15:0]   int_reg_array_32_26_imag;
  reg        [15:0]   int_reg_array_32_27_real;
  reg        [15:0]   int_reg_array_32_27_imag;
  reg        [15:0]   int_reg_array_32_28_real;
  reg        [15:0]   int_reg_array_32_28_imag;
  reg        [15:0]   int_reg_array_32_29_real;
  reg        [15:0]   int_reg_array_32_29_imag;
  reg        [15:0]   int_reg_array_32_30_real;
  reg        [15:0]   int_reg_array_32_30_imag;
  reg        [15:0]   int_reg_array_32_31_real;
  reg        [15:0]   int_reg_array_32_31_imag;
  reg        [15:0]   int_reg_array_32_32_real;
  reg        [15:0]   int_reg_array_32_32_imag;
  reg        [15:0]   int_reg_array_32_33_real;
  reg        [15:0]   int_reg_array_32_33_imag;
  reg        [15:0]   int_reg_array_32_34_real;
  reg        [15:0]   int_reg_array_32_34_imag;
  reg        [15:0]   int_reg_array_32_35_real;
  reg        [15:0]   int_reg_array_32_35_imag;
  reg        [15:0]   int_reg_array_32_36_real;
  reg        [15:0]   int_reg_array_32_36_imag;
  reg        [15:0]   int_reg_array_32_37_real;
  reg        [15:0]   int_reg_array_32_37_imag;
  reg        [15:0]   int_reg_array_32_38_real;
  reg        [15:0]   int_reg_array_32_38_imag;
  reg        [15:0]   int_reg_array_32_39_real;
  reg        [15:0]   int_reg_array_32_39_imag;
  reg        [15:0]   int_reg_array_32_40_real;
  reg        [15:0]   int_reg_array_32_40_imag;
  reg        [15:0]   int_reg_array_32_41_real;
  reg        [15:0]   int_reg_array_32_41_imag;
  reg        [15:0]   int_reg_array_32_42_real;
  reg        [15:0]   int_reg_array_32_42_imag;
  reg        [15:0]   int_reg_array_32_43_real;
  reg        [15:0]   int_reg_array_32_43_imag;
  reg        [15:0]   int_reg_array_32_44_real;
  reg        [15:0]   int_reg_array_32_44_imag;
  reg        [15:0]   int_reg_array_32_45_real;
  reg        [15:0]   int_reg_array_32_45_imag;
  reg        [15:0]   int_reg_array_32_46_real;
  reg        [15:0]   int_reg_array_32_46_imag;
  reg        [15:0]   int_reg_array_32_47_real;
  reg        [15:0]   int_reg_array_32_47_imag;
  reg        [15:0]   int_reg_array_32_48_real;
  reg        [15:0]   int_reg_array_32_48_imag;
  reg        [15:0]   int_reg_array_32_49_real;
  reg        [15:0]   int_reg_array_32_49_imag;
  reg        [15:0]   int_reg_array_32_50_real;
  reg        [15:0]   int_reg_array_32_50_imag;
  reg        [15:0]   int_reg_array_32_51_real;
  reg        [15:0]   int_reg_array_32_51_imag;
  reg        [15:0]   int_reg_array_32_52_real;
  reg        [15:0]   int_reg_array_32_52_imag;
  reg        [15:0]   int_reg_array_32_53_real;
  reg        [15:0]   int_reg_array_32_53_imag;
  reg        [15:0]   int_reg_array_32_54_real;
  reg        [15:0]   int_reg_array_32_54_imag;
  reg        [15:0]   int_reg_array_32_55_real;
  reg        [15:0]   int_reg_array_32_55_imag;
  reg        [15:0]   int_reg_array_32_56_real;
  reg        [15:0]   int_reg_array_32_56_imag;
  reg        [15:0]   int_reg_array_32_57_real;
  reg        [15:0]   int_reg_array_32_57_imag;
  reg        [15:0]   int_reg_array_32_58_real;
  reg        [15:0]   int_reg_array_32_58_imag;
  reg        [15:0]   int_reg_array_32_59_real;
  reg        [15:0]   int_reg_array_32_59_imag;
  reg        [15:0]   int_reg_array_32_60_real;
  reg        [15:0]   int_reg_array_32_60_imag;
  reg        [15:0]   int_reg_array_32_61_real;
  reg        [15:0]   int_reg_array_32_61_imag;
  reg        [15:0]   int_reg_array_32_62_real;
  reg        [15:0]   int_reg_array_32_62_imag;
  reg        [15:0]   int_reg_array_32_63_real;
  reg        [15:0]   int_reg_array_32_63_imag;
  reg        [15:0]   int_reg_array_37_0_real;
  reg        [15:0]   int_reg_array_37_0_imag;
  reg        [15:0]   int_reg_array_37_1_real;
  reg        [15:0]   int_reg_array_37_1_imag;
  reg        [15:0]   int_reg_array_37_2_real;
  reg        [15:0]   int_reg_array_37_2_imag;
  reg        [15:0]   int_reg_array_37_3_real;
  reg        [15:0]   int_reg_array_37_3_imag;
  reg        [15:0]   int_reg_array_37_4_real;
  reg        [15:0]   int_reg_array_37_4_imag;
  reg        [15:0]   int_reg_array_37_5_real;
  reg        [15:0]   int_reg_array_37_5_imag;
  reg        [15:0]   int_reg_array_37_6_real;
  reg        [15:0]   int_reg_array_37_6_imag;
  reg        [15:0]   int_reg_array_37_7_real;
  reg        [15:0]   int_reg_array_37_7_imag;
  reg        [15:0]   int_reg_array_37_8_real;
  reg        [15:0]   int_reg_array_37_8_imag;
  reg        [15:0]   int_reg_array_37_9_real;
  reg        [15:0]   int_reg_array_37_9_imag;
  reg        [15:0]   int_reg_array_37_10_real;
  reg        [15:0]   int_reg_array_37_10_imag;
  reg        [15:0]   int_reg_array_37_11_real;
  reg        [15:0]   int_reg_array_37_11_imag;
  reg        [15:0]   int_reg_array_37_12_real;
  reg        [15:0]   int_reg_array_37_12_imag;
  reg        [15:0]   int_reg_array_37_13_real;
  reg        [15:0]   int_reg_array_37_13_imag;
  reg        [15:0]   int_reg_array_37_14_real;
  reg        [15:0]   int_reg_array_37_14_imag;
  reg        [15:0]   int_reg_array_37_15_real;
  reg        [15:0]   int_reg_array_37_15_imag;
  reg        [15:0]   int_reg_array_37_16_real;
  reg        [15:0]   int_reg_array_37_16_imag;
  reg        [15:0]   int_reg_array_37_17_real;
  reg        [15:0]   int_reg_array_37_17_imag;
  reg        [15:0]   int_reg_array_37_18_real;
  reg        [15:0]   int_reg_array_37_18_imag;
  reg        [15:0]   int_reg_array_37_19_real;
  reg        [15:0]   int_reg_array_37_19_imag;
  reg        [15:0]   int_reg_array_37_20_real;
  reg        [15:0]   int_reg_array_37_20_imag;
  reg        [15:0]   int_reg_array_37_21_real;
  reg        [15:0]   int_reg_array_37_21_imag;
  reg        [15:0]   int_reg_array_37_22_real;
  reg        [15:0]   int_reg_array_37_22_imag;
  reg        [15:0]   int_reg_array_37_23_real;
  reg        [15:0]   int_reg_array_37_23_imag;
  reg        [15:0]   int_reg_array_37_24_real;
  reg        [15:0]   int_reg_array_37_24_imag;
  reg        [15:0]   int_reg_array_37_25_real;
  reg        [15:0]   int_reg_array_37_25_imag;
  reg        [15:0]   int_reg_array_37_26_real;
  reg        [15:0]   int_reg_array_37_26_imag;
  reg        [15:0]   int_reg_array_37_27_real;
  reg        [15:0]   int_reg_array_37_27_imag;
  reg        [15:0]   int_reg_array_37_28_real;
  reg        [15:0]   int_reg_array_37_28_imag;
  reg        [15:0]   int_reg_array_37_29_real;
  reg        [15:0]   int_reg_array_37_29_imag;
  reg        [15:0]   int_reg_array_37_30_real;
  reg        [15:0]   int_reg_array_37_30_imag;
  reg        [15:0]   int_reg_array_37_31_real;
  reg        [15:0]   int_reg_array_37_31_imag;
  reg        [15:0]   int_reg_array_37_32_real;
  reg        [15:0]   int_reg_array_37_32_imag;
  reg        [15:0]   int_reg_array_37_33_real;
  reg        [15:0]   int_reg_array_37_33_imag;
  reg        [15:0]   int_reg_array_37_34_real;
  reg        [15:0]   int_reg_array_37_34_imag;
  reg        [15:0]   int_reg_array_37_35_real;
  reg        [15:0]   int_reg_array_37_35_imag;
  reg        [15:0]   int_reg_array_37_36_real;
  reg        [15:0]   int_reg_array_37_36_imag;
  reg        [15:0]   int_reg_array_37_37_real;
  reg        [15:0]   int_reg_array_37_37_imag;
  reg        [15:0]   int_reg_array_37_38_real;
  reg        [15:0]   int_reg_array_37_38_imag;
  reg        [15:0]   int_reg_array_37_39_real;
  reg        [15:0]   int_reg_array_37_39_imag;
  reg        [15:0]   int_reg_array_37_40_real;
  reg        [15:0]   int_reg_array_37_40_imag;
  reg        [15:0]   int_reg_array_37_41_real;
  reg        [15:0]   int_reg_array_37_41_imag;
  reg        [15:0]   int_reg_array_37_42_real;
  reg        [15:0]   int_reg_array_37_42_imag;
  reg        [15:0]   int_reg_array_37_43_real;
  reg        [15:0]   int_reg_array_37_43_imag;
  reg        [15:0]   int_reg_array_37_44_real;
  reg        [15:0]   int_reg_array_37_44_imag;
  reg        [15:0]   int_reg_array_37_45_real;
  reg        [15:0]   int_reg_array_37_45_imag;
  reg        [15:0]   int_reg_array_37_46_real;
  reg        [15:0]   int_reg_array_37_46_imag;
  reg        [15:0]   int_reg_array_37_47_real;
  reg        [15:0]   int_reg_array_37_47_imag;
  reg        [15:0]   int_reg_array_37_48_real;
  reg        [15:0]   int_reg_array_37_48_imag;
  reg        [15:0]   int_reg_array_37_49_real;
  reg        [15:0]   int_reg_array_37_49_imag;
  reg        [15:0]   int_reg_array_37_50_real;
  reg        [15:0]   int_reg_array_37_50_imag;
  reg        [15:0]   int_reg_array_37_51_real;
  reg        [15:0]   int_reg_array_37_51_imag;
  reg        [15:0]   int_reg_array_37_52_real;
  reg        [15:0]   int_reg_array_37_52_imag;
  reg        [15:0]   int_reg_array_37_53_real;
  reg        [15:0]   int_reg_array_37_53_imag;
  reg        [15:0]   int_reg_array_37_54_real;
  reg        [15:0]   int_reg_array_37_54_imag;
  reg        [15:0]   int_reg_array_37_55_real;
  reg        [15:0]   int_reg_array_37_55_imag;
  reg        [15:0]   int_reg_array_37_56_real;
  reg        [15:0]   int_reg_array_37_56_imag;
  reg        [15:0]   int_reg_array_37_57_real;
  reg        [15:0]   int_reg_array_37_57_imag;
  reg        [15:0]   int_reg_array_37_58_real;
  reg        [15:0]   int_reg_array_37_58_imag;
  reg        [15:0]   int_reg_array_37_59_real;
  reg        [15:0]   int_reg_array_37_59_imag;
  reg        [15:0]   int_reg_array_37_60_real;
  reg        [15:0]   int_reg_array_37_60_imag;
  reg        [15:0]   int_reg_array_37_61_real;
  reg        [15:0]   int_reg_array_37_61_imag;
  reg        [15:0]   int_reg_array_37_62_real;
  reg        [15:0]   int_reg_array_37_62_imag;
  reg        [15:0]   int_reg_array_37_63_real;
  reg        [15:0]   int_reg_array_37_63_imag;
  reg        [15:0]   int_reg_array_27_0_real;
  reg        [15:0]   int_reg_array_27_0_imag;
  reg        [15:0]   int_reg_array_27_1_real;
  reg        [15:0]   int_reg_array_27_1_imag;
  reg        [15:0]   int_reg_array_27_2_real;
  reg        [15:0]   int_reg_array_27_2_imag;
  reg        [15:0]   int_reg_array_27_3_real;
  reg        [15:0]   int_reg_array_27_3_imag;
  reg        [15:0]   int_reg_array_27_4_real;
  reg        [15:0]   int_reg_array_27_4_imag;
  reg        [15:0]   int_reg_array_27_5_real;
  reg        [15:0]   int_reg_array_27_5_imag;
  reg        [15:0]   int_reg_array_27_6_real;
  reg        [15:0]   int_reg_array_27_6_imag;
  reg        [15:0]   int_reg_array_27_7_real;
  reg        [15:0]   int_reg_array_27_7_imag;
  reg        [15:0]   int_reg_array_27_8_real;
  reg        [15:0]   int_reg_array_27_8_imag;
  reg        [15:0]   int_reg_array_27_9_real;
  reg        [15:0]   int_reg_array_27_9_imag;
  reg        [15:0]   int_reg_array_27_10_real;
  reg        [15:0]   int_reg_array_27_10_imag;
  reg        [15:0]   int_reg_array_27_11_real;
  reg        [15:0]   int_reg_array_27_11_imag;
  reg        [15:0]   int_reg_array_27_12_real;
  reg        [15:0]   int_reg_array_27_12_imag;
  reg        [15:0]   int_reg_array_27_13_real;
  reg        [15:0]   int_reg_array_27_13_imag;
  reg        [15:0]   int_reg_array_27_14_real;
  reg        [15:0]   int_reg_array_27_14_imag;
  reg        [15:0]   int_reg_array_27_15_real;
  reg        [15:0]   int_reg_array_27_15_imag;
  reg        [15:0]   int_reg_array_27_16_real;
  reg        [15:0]   int_reg_array_27_16_imag;
  reg        [15:0]   int_reg_array_27_17_real;
  reg        [15:0]   int_reg_array_27_17_imag;
  reg        [15:0]   int_reg_array_27_18_real;
  reg        [15:0]   int_reg_array_27_18_imag;
  reg        [15:0]   int_reg_array_27_19_real;
  reg        [15:0]   int_reg_array_27_19_imag;
  reg        [15:0]   int_reg_array_27_20_real;
  reg        [15:0]   int_reg_array_27_20_imag;
  reg        [15:0]   int_reg_array_27_21_real;
  reg        [15:0]   int_reg_array_27_21_imag;
  reg        [15:0]   int_reg_array_27_22_real;
  reg        [15:0]   int_reg_array_27_22_imag;
  reg        [15:0]   int_reg_array_27_23_real;
  reg        [15:0]   int_reg_array_27_23_imag;
  reg        [15:0]   int_reg_array_27_24_real;
  reg        [15:0]   int_reg_array_27_24_imag;
  reg        [15:0]   int_reg_array_27_25_real;
  reg        [15:0]   int_reg_array_27_25_imag;
  reg        [15:0]   int_reg_array_27_26_real;
  reg        [15:0]   int_reg_array_27_26_imag;
  reg        [15:0]   int_reg_array_27_27_real;
  reg        [15:0]   int_reg_array_27_27_imag;
  reg        [15:0]   int_reg_array_27_28_real;
  reg        [15:0]   int_reg_array_27_28_imag;
  reg        [15:0]   int_reg_array_27_29_real;
  reg        [15:0]   int_reg_array_27_29_imag;
  reg        [15:0]   int_reg_array_27_30_real;
  reg        [15:0]   int_reg_array_27_30_imag;
  reg        [15:0]   int_reg_array_27_31_real;
  reg        [15:0]   int_reg_array_27_31_imag;
  reg        [15:0]   int_reg_array_27_32_real;
  reg        [15:0]   int_reg_array_27_32_imag;
  reg        [15:0]   int_reg_array_27_33_real;
  reg        [15:0]   int_reg_array_27_33_imag;
  reg        [15:0]   int_reg_array_27_34_real;
  reg        [15:0]   int_reg_array_27_34_imag;
  reg        [15:0]   int_reg_array_27_35_real;
  reg        [15:0]   int_reg_array_27_35_imag;
  reg        [15:0]   int_reg_array_27_36_real;
  reg        [15:0]   int_reg_array_27_36_imag;
  reg        [15:0]   int_reg_array_27_37_real;
  reg        [15:0]   int_reg_array_27_37_imag;
  reg        [15:0]   int_reg_array_27_38_real;
  reg        [15:0]   int_reg_array_27_38_imag;
  reg        [15:0]   int_reg_array_27_39_real;
  reg        [15:0]   int_reg_array_27_39_imag;
  reg        [15:0]   int_reg_array_27_40_real;
  reg        [15:0]   int_reg_array_27_40_imag;
  reg        [15:0]   int_reg_array_27_41_real;
  reg        [15:0]   int_reg_array_27_41_imag;
  reg        [15:0]   int_reg_array_27_42_real;
  reg        [15:0]   int_reg_array_27_42_imag;
  reg        [15:0]   int_reg_array_27_43_real;
  reg        [15:0]   int_reg_array_27_43_imag;
  reg        [15:0]   int_reg_array_27_44_real;
  reg        [15:0]   int_reg_array_27_44_imag;
  reg        [15:0]   int_reg_array_27_45_real;
  reg        [15:0]   int_reg_array_27_45_imag;
  reg        [15:0]   int_reg_array_27_46_real;
  reg        [15:0]   int_reg_array_27_46_imag;
  reg        [15:0]   int_reg_array_27_47_real;
  reg        [15:0]   int_reg_array_27_47_imag;
  reg        [15:0]   int_reg_array_27_48_real;
  reg        [15:0]   int_reg_array_27_48_imag;
  reg        [15:0]   int_reg_array_27_49_real;
  reg        [15:0]   int_reg_array_27_49_imag;
  reg        [15:0]   int_reg_array_27_50_real;
  reg        [15:0]   int_reg_array_27_50_imag;
  reg        [15:0]   int_reg_array_27_51_real;
  reg        [15:0]   int_reg_array_27_51_imag;
  reg        [15:0]   int_reg_array_27_52_real;
  reg        [15:0]   int_reg_array_27_52_imag;
  reg        [15:0]   int_reg_array_27_53_real;
  reg        [15:0]   int_reg_array_27_53_imag;
  reg        [15:0]   int_reg_array_27_54_real;
  reg        [15:0]   int_reg_array_27_54_imag;
  reg        [15:0]   int_reg_array_27_55_real;
  reg        [15:0]   int_reg_array_27_55_imag;
  reg        [15:0]   int_reg_array_27_56_real;
  reg        [15:0]   int_reg_array_27_56_imag;
  reg        [15:0]   int_reg_array_27_57_real;
  reg        [15:0]   int_reg_array_27_57_imag;
  reg        [15:0]   int_reg_array_27_58_real;
  reg        [15:0]   int_reg_array_27_58_imag;
  reg        [15:0]   int_reg_array_27_59_real;
  reg        [15:0]   int_reg_array_27_59_imag;
  reg        [15:0]   int_reg_array_27_60_real;
  reg        [15:0]   int_reg_array_27_60_imag;
  reg        [15:0]   int_reg_array_27_61_real;
  reg        [15:0]   int_reg_array_27_61_imag;
  reg        [15:0]   int_reg_array_27_62_real;
  reg        [15:0]   int_reg_array_27_62_imag;
  reg        [15:0]   int_reg_array_27_63_real;
  reg        [15:0]   int_reg_array_27_63_imag;
  reg        [15:0]   int_reg_array_16_0_real;
  reg        [15:0]   int_reg_array_16_0_imag;
  reg        [15:0]   int_reg_array_16_1_real;
  reg        [15:0]   int_reg_array_16_1_imag;
  reg        [15:0]   int_reg_array_16_2_real;
  reg        [15:0]   int_reg_array_16_2_imag;
  reg        [15:0]   int_reg_array_16_3_real;
  reg        [15:0]   int_reg_array_16_3_imag;
  reg        [15:0]   int_reg_array_16_4_real;
  reg        [15:0]   int_reg_array_16_4_imag;
  reg        [15:0]   int_reg_array_16_5_real;
  reg        [15:0]   int_reg_array_16_5_imag;
  reg        [15:0]   int_reg_array_16_6_real;
  reg        [15:0]   int_reg_array_16_6_imag;
  reg        [15:0]   int_reg_array_16_7_real;
  reg        [15:0]   int_reg_array_16_7_imag;
  reg        [15:0]   int_reg_array_16_8_real;
  reg        [15:0]   int_reg_array_16_8_imag;
  reg        [15:0]   int_reg_array_16_9_real;
  reg        [15:0]   int_reg_array_16_9_imag;
  reg        [15:0]   int_reg_array_16_10_real;
  reg        [15:0]   int_reg_array_16_10_imag;
  reg        [15:0]   int_reg_array_16_11_real;
  reg        [15:0]   int_reg_array_16_11_imag;
  reg        [15:0]   int_reg_array_16_12_real;
  reg        [15:0]   int_reg_array_16_12_imag;
  reg        [15:0]   int_reg_array_16_13_real;
  reg        [15:0]   int_reg_array_16_13_imag;
  reg        [15:0]   int_reg_array_16_14_real;
  reg        [15:0]   int_reg_array_16_14_imag;
  reg        [15:0]   int_reg_array_16_15_real;
  reg        [15:0]   int_reg_array_16_15_imag;
  reg        [15:0]   int_reg_array_16_16_real;
  reg        [15:0]   int_reg_array_16_16_imag;
  reg        [15:0]   int_reg_array_16_17_real;
  reg        [15:0]   int_reg_array_16_17_imag;
  reg        [15:0]   int_reg_array_16_18_real;
  reg        [15:0]   int_reg_array_16_18_imag;
  reg        [15:0]   int_reg_array_16_19_real;
  reg        [15:0]   int_reg_array_16_19_imag;
  reg        [15:0]   int_reg_array_16_20_real;
  reg        [15:0]   int_reg_array_16_20_imag;
  reg        [15:0]   int_reg_array_16_21_real;
  reg        [15:0]   int_reg_array_16_21_imag;
  reg        [15:0]   int_reg_array_16_22_real;
  reg        [15:0]   int_reg_array_16_22_imag;
  reg        [15:0]   int_reg_array_16_23_real;
  reg        [15:0]   int_reg_array_16_23_imag;
  reg        [15:0]   int_reg_array_16_24_real;
  reg        [15:0]   int_reg_array_16_24_imag;
  reg        [15:0]   int_reg_array_16_25_real;
  reg        [15:0]   int_reg_array_16_25_imag;
  reg        [15:0]   int_reg_array_16_26_real;
  reg        [15:0]   int_reg_array_16_26_imag;
  reg        [15:0]   int_reg_array_16_27_real;
  reg        [15:0]   int_reg_array_16_27_imag;
  reg        [15:0]   int_reg_array_16_28_real;
  reg        [15:0]   int_reg_array_16_28_imag;
  reg        [15:0]   int_reg_array_16_29_real;
  reg        [15:0]   int_reg_array_16_29_imag;
  reg        [15:0]   int_reg_array_16_30_real;
  reg        [15:0]   int_reg_array_16_30_imag;
  reg        [15:0]   int_reg_array_16_31_real;
  reg        [15:0]   int_reg_array_16_31_imag;
  reg        [15:0]   int_reg_array_16_32_real;
  reg        [15:0]   int_reg_array_16_32_imag;
  reg        [15:0]   int_reg_array_16_33_real;
  reg        [15:0]   int_reg_array_16_33_imag;
  reg        [15:0]   int_reg_array_16_34_real;
  reg        [15:0]   int_reg_array_16_34_imag;
  reg        [15:0]   int_reg_array_16_35_real;
  reg        [15:0]   int_reg_array_16_35_imag;
  reg        [15:0]   int_reg_array_16_36_real;
  reg        [15:0]   int_reg_array_16_36_imag;
  reg        [15:0]   int_reg_array_16_37_real;
  reg        [15:0]   int_reg_array_16_37_imag;
  reg        [15:0]   int_reg_array_16_38_real;
  reg        [15:0]   int_reg_array_16_38_imag;
  reg        [15:0]   int_reg_array_16_39_real;
  reg        [15:0]   int_reg_array_16_39_imag;
  reg        [15:0]   int_reg_array_16_40_real;
  reg        [15:0]   int_reg_array_16_40_imag;
  reg        [15:0]   int_reg_array_16_41_real;
  reg        [15:0]   int_reg_array_16_41_imag;
  reg        [15:0]   int_reg_array_16_42_real;
  reg        [15:0]   int_reg_array_16_42_imag;
  reg        [15:0]   int_reg_array_16_43_real;
  reg        [15:0]   int_reg_array_16_43_imag;
  reg        [15:0]   int_reg_array_16_44_real;
  reg        [15:0]   int_reg_array_16_44_imag;
  reg        [15:0]   int_reg_array_16_45_real;
  reg        [15:0]   int_reg_array_16_45_imag;
  reg        [15:0]   int_reg_array_16_46_real;
  reg        [15:0]   int_reg_array_16_46_imag;
  reg        [15:0]   int_reg_array_16_47_real;
  reg        [15:0]   int_reg_array_16_47_imag;
  reg        [15:0]   int_reg_array_16_48_real;
  reg        [15:0]   int_reg_array_16_48_imag;
  reg        [15:0]   int_reg_array_16_49_real;
  reg        [15:0]   int_reg_array_16_49_imag;
  reg        [15:0]   int_reg_array_16_50_real;
  reg        [15:0]   int_reg_array_16_50_imag;
  reg        [15:0]   int_reg_array_16_51_real;
  reg        [15:0]   int_reg_array_16_51_imag;
  reg        [15:0]   int_reg_array_16_52_real;
  reg        [15:0]   int_reg_array_16_52_imag;
  reg        [15:0]   int_reg_array_16_53_real;
  reg        [15:0]   int_reg_array_16_53_imag;
  reg        [15:0]   int_reg_array_16_54_real;
  reg        [15:0]   int_reg_array_16_54_imag;
  reg        [15:0]   int_reg_array_16_55_real;
  reg        [15:0]   int_reg_array_16_55_imag;
  reg        [15:0]   int_reg_array_16_56_real;
  reg        [15:0]   int_reg_array_16_56_imag;
  reg        [15:0]   int_reg_array_16_57_real;
  reg        [15:0]   int_reg_array_16_57_imag;
  reg        [15:0]   int_reg_array_16_58_real;
  reg        [15:0]   int_reg_array_16_58_imag;
  reg        [15:0]   int_reg_array_16_59_real;
  reg        [15:0]   int_reg_array_16_59_imag;
  reg        [15:0]   int_reg_array_16_60_real;
  reg        [15:0]   int_reg_array_16_60_imag;
  reg        [15:0]   int_reg_array_16_61_real;
  reg        [15:0]   int_reg_array_16_61_imag;
  reg        [15:0]   int_reg_array_16_62_real;
  reg        [15:0]   int_reg_array_16_62_imag;
  reg        [15:0]   int_reg_array_16_63_real;
  reg        [15:0]   int_reg_array_16_63_imag;
  reg        [15:0]   int_reg_array_21_0_real;
  reg        [15:0]   int_reg_array_21_0_imag;
  reg        [15:0]   int_reg_array_21_1_real;
  reg        [15:0]   int_reg_array_21_1_imag;
  reg        [15:0]   int_reg_array_21_2_real;
  reg        [15:0]   int_reg_array_21_2_imag;
  reg        [15:0]   int_reg_array_21_3_real;
  reg        [15:0]   int_reg_array_21_3_imag;
  reg        [15:0]   int_reg_array_21_4_real;
  reg        [15:0]   int_reg_array_21_4_imag;
  reg        [15:0]   int_reg_array_21_5_real;
  reg        [15:0]   int_reg_array_21_5_imag;
  reg        [15:0]   int_reg_array_21_6_real;
  reg        [15:0]   int_reg_array_21_6_imag;
  reg        [15:0]   int_reg_array_21_7_real;
  reg        [15:0]   int_reg_array_21_7_imag;
  reg        [15:0]   int_reg_array_21_8_real;
  reg        [15:0]   int_reg_array_21_8_imag;
  reg        [15:0]   int_reg_array_21_9_real;
  reg        [15:0]   int_reg_array_21_9_imag;
  reg        [15:0]   int_reg_array_21_10_real;
  reg        [15:0]   int_reg_array_21_10_imag;
  reg        [15:0]   int_reg_array_21_11_real;
  reg        [15:0]   int_reg_array_21_11_imag;
  reg        [15:0]   int_reg_array_21_12_real;
  reg        [15:0]   int_reg_array_21_12_imag;
  reg        [15:0]   int_reg_array_21_13_real;
  reg        [15:0]   int_reg_array_21_13_imag;
  reg        [15:0]   int_reg_array_21_14_real;
  reg        [15:0]   int_reg_array_21_14_imag;
  reg        [15:0]   int_reg_array_21_15_real;
  reg        [15:0]   int_reg_array_21_15_imag;
  reg        [15:0]   int_reg_array_21_16_real;
  reg        [15:0]   int_reg_array_21_16_imag;
  reg        [15:0]   int_reg_array_21_17_real;
  reg        [15:0]   int_reg_array_21_17_imag;
  reg        [15:0]   int_reg_array_21_18_real;
  reg        [15:0]   int_reg_array_21_18_imag;
  reg        [15:0]   int_reg_array_21_19_real;
  reg        [15:0]   int_reg_array_21_19_imag;
  reg        [15:0]   int_reg_array_21_20_real;
  reg        [15:0]   int_reg_array_21_20_imag;
  reg        [15:0]   int_reg_array_21_21_real;
  reg        [15:0]   int_reg_array_21_21_imag;
  reg        [15:0]   int_reg_array_21_22_real;
  reg        [15:0]   int_reg_array_21_22_imag;
  reg        [15:0]   int_reg_array_21_23_real;
  reg        [15:0]   int_reg_array_21_23_imag;
  reg        [15:0]   int_reg_array_21_24_real;
  reg        [15:0]   int_reg_array_21_24_imag;
  reg        [15:0]   int_reg_array_21_25_real;
  reg        [15:0]   int_reg_array_21_25_imag;
  reg        [15:0]   int_reg_array_21_26_real;
  reg        [15:0]   int_reg_array_21_26_imag;
  reg        [15:0]   int_reg_array_21_27_real;
  reg        [15:0]   int_reg_array_21_27_imag;
  reg        [15:0]   int_reg_array_21_28_real;
  reg        [15:0]   int_reg_array_21_28_imag;
  reg        [15:0]   int_reg_array_21_29_real;
  reg        [15:0]   int_reg_array_21_29_imag;
  reg        [15:0]   int_reg_array_21_30_real;
  reg        [15:0]   int_reg_array_21_30_imag;
  reg        [15:0]   int_reg_array_21_31_real;
  reg        [15:0]   int_reg_array_21_31_imag;
  reg        [15:0]   int_reg_array_21_32_real;
  reg        [15:0]   int_reg_array_21_32_imag;
  reg        [15:0]   int_reg_array_21_33_real;
  reg        [15:0]   int_reg_array_21_33_imag;
  reg        [15:0]   int_reg_array_21_34_real;
  reg        [15:0]   int_reg_array_21_34_imag;
  reg        [15:0]   int_reg_array_21_35_real;
  reg        [15:0]   int_reg_array_21_35_imag;
  reg        [15:0]   int_reg_array_21_36_real;
  reg        [15:0]   int_reg_array_21_36_imag;
  reg        [15:0]   int_reg_array_21_37_real;
  reg        [15:0]   int_reg_array_21_37_imag;
  reg        [15:0]   int_reg_array_21_38_real;
  reg        [15:0]   int_reg_array_21_38_imag;
  reg        [15:0]   int_reg_array_21_39_real;
  reg        [15:0]   int_reg_array_21_39_imag;
  reg        [15:0]   int_reg_array_21_40_real;
  reg        [15:0]   int_reg_array_21_40_imag;
  reg        [15:0]   int_reg_array_21_41_real;
  reg        [15:0]   int_reg_array_21_41_imag;
  reg        [15:0]   int_reg_array_21_42_real;
  reg        [15:0]   int_reg_array_21_42_imag;
  reg        [15:0]   int_reg_array_21_43_real;
  reg        [15:0]   int_reg_array_21_43_imag;
  reg        [15:0]   int_reg_array_21_44_real;
  reg        [15:0]   int_reg_array_21_44_imag;
  reg        [15:0]   int_reg_array_21_45_real;
  reg        [15:0]   int_reg_array_21_45_imag;
  reg        [15:0]   int_reg_array_21_46_real;
  reg        [15:0]   int_reg_array_21_46_imag;
  reg        [15:0]   int_reg_array_21_47_real;
  reg        [15:0]   int_reg_array_21_47_imag;
  reg        [15:0]   int_reg_array_21_48_real;
  reg        [15:0]   int_reg_array_21_48_imag;
  reg        [15:0]   int_reg_array_21_49_real;
  reg        [15:0]   int_reg_array_21_49_imag;
  reg        [15:0]   int_reg_array_21_50_real;
  reg        [15:0]   int_reg_array_21_50_imag;
  reg        [15:0]   int_reg_array_21_51_real;
  reg        [15:0]   int_reg_array_21_51_imag;
  reg        [15:0]   int_reg_array_21_52_real;
  reg        [15:0]   int_reg_array_21_52_imag;
  reg        [15:0]   int_reg_array_21_53_real;
  reg        [15:0]   int_reg_array_21_53_imag;
  reg        [15:0]   int_reg_array_21_54_real;
  reg        [15:0]   int_reg_array_21_54_imag;
  reg        [15:0]   int_reg_array_21_55_real;
  reg        [15:0]   int_reg_array_21_55_imag;
  reg        [15:0]   int_reg_array_21_56_real;
  reg        [15:0]   int_reg_array_21_56_imag;
  reg        [15:0]   int_reg_array_21_57_real;
  reg        [15:0]   int_reg_array_21_57_imag;
  reg        [15:0]   int_reg_array_21_58_real;
  reg        [15:0]   int_reg_array_21_58_imag;
  reg        [15:0]   int_reg_array_21_59_real;
  reg        [15:0]   int_reg_array_21_59_imag;
  reg        [15:0]   int_reg_array_21_60_real;
  reg        [15:0]   int_reg_array_21_60_imag;
  reg        [15:0]   int_reg_array_21_61_real;
  reg        [15:0]   int_reg_array_21_61_imag;
  reg        [15:0]   int_reg_array_21_62_real;
  reg        [15:0]   int_reg_array_21_62_imag;
  reg        [15:0]   int_reg_array_21_63_real;
  reg        [15:0]   int_reg_array_21_63_imag;
  reg        [15:0]   int_reg_array_46_0_real;
  reg        [15:0]   int_reg_array_46_0_imag;
  reg        [15:0]   int_reg_array_46_1_real;
  reg        [15:0]   int_reg_array_46_1_imag;
  reg        [15:0]   int_reg_array_46_2_real;
  reg        [15:0]   int_reg_array_46_2_imag;
  reg        [15:0]   int_reg_array_46_3_real;
  reg        [15:0]   int_reg_array_46_3_imag;
  reg        [15:0]   int_reg_array_46_4_real;
  reg        [15:0]   int_reg_array_46_4_imag;
  reg        [15:0]   int_reg_array_46_5_real;
  reg        [15:0]   int_reg_array_46_5_imag;
  reg        [15:0]   int_reg_array_46_6_real;
  reg        [15:0]   int_reg_array_46_6_imag;
  reg        [15:0]   int_reg_array_46_7_real;
  reg        [15:0]   int_reg_array_46_7_imag;
  reg        [15:0]   int_reg_array_46_8_real;
  reg        [15:0]   int_reg_array_46_8_imag;
  reg        [15:0]   int_reg_array_46_9_real;
  reg        [15:0]   int_reg_array_46_9_imag;
  reg        [15:0]   int_reg_array_46_10_real;
  reg        [15:0]   int_reg_array_46_10_imag;
  reg        [15:0]   int_reg_array_46_11_real;
  reg        [15:0]   int_reg_array_46_11_imag;
  reg        [15:0]   int_reg_array_46_12_real;
  reg        [15:0]   int_reg_array_46_12_imag;
  reg        [15:0]   int_reg_array_46_13_real;
  reg        [15:0]   int_reg_array_46_13_imag;
  reg        [15:0]   int_reg_array_46_14_real;
  reg        [15:0]   int_reg_array_46_14_imag;
  reg        [15:0]   int_reg_array_46_15_real;
  reg        [15:0]   int_reg_array_46_15_imag;
  reg        [15:0]   int_reg_array_46_16_real;
  reg        [15:0]   int_reg_array_46_16_imag;
  reg        [15:0]   int_reg_array_46_17_real;
  reg        [15:0]   int_reg_array_46_17_imag;
  reg        [15:0]   int_reg_array_46_18_real;
  reg        [15:0]   int_reg_array_46_18_imag;
  reg        [15:0]   int_reg_array_46_19_real;
  reg        [15:0]   int_reg_array_46_19_imag;
  reg        [15:0]   int_reg_array_46_20_real;
  reg        [15:0]   int_reg_array_46_20_imag;
  reg        [15:0]   int_reg_array_46_21_real;
  reg        [15:0]   int_reg_array_46_21_imag;
  reg        [15:0]   int_reg_array_46_22_real;
  reg        [15:0]   int_reg_array_46_22_imag;
  reg        [15:0]   int_reg_array_46_23_real;
  reg        [15:0]   int_reg_array_46_23_imag;
  reg        [15:0]   int_reg_array_46_24_real;
  reg        [15:0]   int_reg_array_46_24_imag;
  reg        [15:0]   int_reg_array_46_25_real;
  reg        [15:0]   int_reg_array_46_25_imag;
  reg        [15:0]   int_reg_array_46_26_real;
  reg        [15:0]   int_reg_array_46_26_imag;
  reg        [15:0]   int_reg_array_46_27_real;
  reg        [15:0]   int_reg_array_46_27_imag;
  reg        [15:0]   int_reg_array_46_28_real;
  reg        [15:0]   int_reg_array_46_28_imag;
  reg        [15:0]   int_reg_array_46_29_real;
  reg        [15:0]   int_reg_array_46_29_imag;
  reg        [15:0]   int_reg_array_46_30_real;
  reg        [15:0]   int_reg_array_46_30_imag;
  reg        [15:0]   int_reg_array_46_31_real;
  reg        [15:0]   int_reg_array_46_31_imag;
  reg        [15:0]   int_reg_array_46_32_real;
  reg        [15:0]   int_reg_array_46_32_imag;
  reg        [15:0]   int_reg_array_46_33_real;
  reg        [15:0]   int_reg_array_46_33_imag;
  reg        [15:0]   int_reg_array_46_34_real;
  reg        [15:0]   int_reg_array_46_34_imag;
  reg        [15:0]   int_reg_array_46_35_real;
  reg        [15:0]   int_reg_array_46_35_imag;
  reg        [15:0]   int_reg_array_46_36_real;
  reg        [15:0]   int_reg_array_46_36_imag;
  reg        [15:0]   int_reg_array_46_37_real;
  reg        [15:0]   int_reg_array_46_37_imag;
  reg        [15:0]   int_reg_array_46_38_real;
  reg        [15:0]   int_reg_array_46_38_imag;
  reg        [15:0]   int_reg_array_46_39_real;
  reg        [15:0]   int_reg_array_46_39_imag;
  reg        [15:0]   int_reg_array_46_40_real;
  reg        [15:0]   int_reg_array_46_40_imag;
  reg        [15:0]   int_reg_array_46_41_real;
  reg        [15:0]   int_reg_array_46_41_imag;
  reg        [15:0]   int_reg_array_46_42_real;
  reg        [15:0]   int_reg_array_46_42_imag;
  reg        [15:0]   int_reg_array_46_43_real;
  reg        [15:0]   int_reg_array_46_43_imag;
  reg        [15:0]   int_reg_array_46_44_real;
  reg        [15:0]   int_reg_array_46_44_imag;
  reg        [15:0]   int_reg_array_46_45_real;
  reg        [15:0]   int_reg_array_46_45_imag;
  reg        [15:0]   int_reg_array_46_46_real;
  reg        [15:0]   int_reg_array_46_46_imag;
  reg        [15:0]   int_reg_array_46_47_real;
  reg        [15:0]   int_reg_array_46_47_imag;
  reg        [15:0]   int_reg_array_46_48_real;
  reg        [15:0]   int_reg_array_46_48_imag;
  reg        [15:0]   int_reg_array_46_49_real;
  reg        [15:0]   int_reg_array_46_49_imag;
  reg        [15:0]   int_reg_array_46_50_real;
  reg        [15:0]   int_reg_array_46_50_imag;
  reg        [15:0]   int_reg_array_46_51_real;
  reg        [15:0]   int_reg_array_46_51_imag;
  reg        [15:0]   int_reg_array_46_52_real;
  reg        [15:0]   int_reg_array_46_52_imag;
  reg        [15:0]   int_reg_array_46_53_real;
  reg        [15:0]   int_reg_array_46_53_imag;
  reg        [15:0]   int_reg_array_46_54_real;
  reg        [15:0]   int_reg_array_46_54_imag;
  reg        [15:0]   int_reg_array_46_55_real;
  reg        [15:0]   int_reg_array_46_55_imag;
  reg        [15:0]   int_reg_array_46_56_real;
  reg        [15:0]   int_reg_array_46_56_imag;
  reg        [15:0]   int_reg_array_46_57_real;
  reg        [15:0]   int_reg_array_46_57_imag;
  reg        [15:0]   int_reg_array_46_58_real;
  reg        [15:0]   int_reg_array_46_58_imag;
  reg        [15:0]   int_reg_array_46_59_real;
  reg        [15:0]   int_reg_array_46_59_imag;
  reg        [15:0]   int_reg_array_46_60_real;
  reg        [15:0]   int_reg_array_46_60_imag;
  reg        [15:0]   int_reg_array_46_61_real;
  reg        [15:0]   int_reg_array_46_61_imag;
  reg        [15:0]   int_reg_array_46_62_real;
  reg        [15:0]   int_reg_array_46_62_imag;
  reg        [15:0]   int_reg_array_46_63_real;
  reg        [15:0]   int_reg_array_46_63_imag;
  reg        [15:0]   int_reg_array_10_0_real;
  reg        [15:0]   int_reg_array_10_0_imag;
  reg        [15:0]   int_reg_array_10_1_real;
  reg        [15:0]   int_reg_array_10_1_imag;
  reg        [15:0]   int_reg_array_10_2_real;
  reg        [15:0]   int_reg_array_10_2_imag;
  reg        [15:0]   int_reg_array_10_3_real;
  reg        [15:0]   int_reg_array_10_3_imag;
  reg        [15:0]   int_reg_array_10_4_real;
  reg        [15:0]   int_reg_array_10_4_imag;
  reg        [15:0]   int_reg_array_10_5_real;
  reg        [15:0]   int_reg_array_10_5_imag;
  reg        [15:0]   int_reg_array_10_6_real;
  reg        [15:0]   int_reg_array_10_6_imag;
  reg        [15:0]   int_reg_array_10_7_real;
  reg        [15:0]   int_reg_array_10_7_imag;
  reg        [15:0]   int_reg_array_10_8_real;
  reg        [15:0]   int_reg_array_10_8_imag;
  reg        [15:0]   int_reg_array_10_9_real;
  reg        [15:0]   int_reg_array_10_9_imag;
  reg        [15:0]   int_reg_array_10_10_real;
  reg        [15:0]   int_reg_array_10_10_imag;
  reg        [15:0]   int_reg_array_10_11_real;
  reg        [15:0]   int_reg_array_10_11_imag;
  reg        [15:0]   int_reg_array_10_12_real;
  reg        [15:0]   int_reg_array_10_12_imag;
  reg        [15:0]   int_reg_array_10_13_real;
  reg        [15:0]   int_reg_array_10_13_imag;
  reg        [15:0]   int_reg_array_10_14_real;
  reg        [15:0]   int_reg_array_10_14_imag;
  reg        [15:0]   int_reg_array_10_15_real;
  reg        [15:0]   int_reg_array_10_15_imag;
  reg        [15:0]   int_reg_array_10_16_real;
  reg        [15:0]   int_reg_array_10_16_imag;
  reg        [15:0]   int_reg_array_10_17_real;
  reg        [15:0]   int_reg_array_10_17_imag;
  reg        [15:0]   int_reg_array_10_18_real;
  reg        [15:0]   int_reg_array_10_18_imag;
  reg        [15:0]   int_reg_array_10_19_real;
  reg        [15:0]   int_reg_array_10_19_imag;
  reg        [15:0]   int_reg_array_10_20_real;
  reg        [15:0]   int_reg_array_10_20_imag;
  reg        [15:0]   int_reg_array_10_21_real;
  reg        [15:0]   int_reg_array_10_21_imag;
  reg        [15:0]   int_reg_array_10_22_real;
  reg        [15:0]   int_reg_array_10_22_imag;
  reg        [15:0]   int_reg_array_10_23_real;
  reg        [15:0]   int_reg_array_10_23_imag;
  reg        [15:0]   int_reg_array_10_24_real;
  reg        [15:0]   int_reg_array_10_24_imag;
  reg        [15:0]   int_reg_array_10_25_real;
  reg        [15:0]   int_reg_array_10_25_imag;
  reg        [15:0]   int_reg_array_10_26_real;
  reg        [15:0]   int_reg_array_10_26_imag;
  reg        [15:0]   int_reg_array_10_27_real;
  reg        [15:0]   int_reg_array_10_27_imag;
  reg        [15:0]   int_reg_array_10_28_real;
  reg        [15:0]   int_reg_array_10_28_imag;
  reg        [15:0]   int_reg_array_10_29_real;
  reg        [15:0]   int_reg_array_10_29_imag;
  reg        [15:0]   int_reg_array_10_30_real;
  reg        [15:0]   int_reg_array_10_30_imag;
  reg        [15:0]   int_reg_array_10_31_real;
  reg        [15:0]   int_reg_array_10_31_imag;
  reg        [15:0]   int_reg_array_10_32_real;
  reg        [15:0]   int_reg_array_10_32_imag;
  reg        [15:0]   int_reg_array_10_33_real;
  reg        [15:0]   int_reg_array_10_33_imag;
  reg        [15:0]   int_reg_array_10_34_real;
  reg        [15:0]   int_reg_array_10_34_imag;
  reg        [15:0]   int_reg_array_10_35_real;
  reg        [15:0]   int_reg_array_10_35_imag;
  reg        [15:0]   int_reg_array_10_36_real;
  reg        [15:0]   int_reg_array_10_36_imag;
  reg        [15:0]   int_reg_array_10_37_real;
  reg        [15:0]   int_reg_array_10_37_imag;
  reg        [15:0]   int_reg_array_10_38_real;
  reg        [15:0]   int_reg_array_10_38_imag;
  reg        [15:0]   int_reg_array_10_39_real;
  reg        [15:0]   int_reg_array_10_39_imag;
  reg        [15:0]   int_reg_array_10_40_real;
  reg        [15:0]   int_reg_array_10_40_imag;
  reg        [15:0]   int_reg_array_10_41_real;
  reg        [15:0]   int_reg_array_10_41_imag;
  reg        [15:0]   int_reg_array_10_42_real;
  reg        [15:0]   int_reg_array_10_42_imag;
  reg        [15:0]   int_reg_array_10_43_real;
  reg        [15:0]   int_reg_array_10_43_imag;
  reg        [15:0]   int_reg_array_10_44_real;
  reg        [15:0]   int_reg_array_10_44_imag;
  reg        [15:0]   int_reg_array_10_45_real;
  reg        [15:0]   int_reg_array_10_45_imag;
  reg        [15:0]   int_reg_array_10_46_real;
  reg        [15:0]   int_reg_array_10_46_imag;
  reg        [15:0]   int_reg_array_10_47_real;
  reg        [15:0]   int_reg_array_10_47_imag;
  reg        [15:0]   int_reg_array_10_48_real;
  reg        [15:0]   int_reg_array_10_48_imag;
  reg        [15:0]   int_reg_array_10_49_real;
  reg        [15:0]   int_reg_array_10_49_imag;
  reg        [15:0]   int_reg_array_10_50_real;
  reg        [15:0]   int_reg_array_10_50_imag;
  reg        [15:0]   int_reg_array_10_51_real;
  reg        [15:0]   int_reg_array_10_51_imag;
  reg        [15:0]   int_reg_array_10_52_real;
  reg        [15:0]   int_reg_array_10_52_imag;
  reg        [15:0]   int_reg_array_10_53_real;
  reg        [15:0]   int_reg_array_10_53_imag;
  reg        [15:0]   int_reg_array_10_54_real;
  reg        [15:0]   int_reg_array_10_54_imag;
  reg        [15:0]   int_reg_array_10_55_real;
  reg        [15:0]   int_reg_array_10_55_imag;
  reg        [15:0]   int_reg_array_10_56_real;
  reg        [15:0]   int_reg_array_10_56_imag;
  reg        [15:0]   int_reg_array_10_57_real;
  reg        [15:0]   int_reg_array_10_57_imag;
  reg        [15:0]   int_reg_array_10_58_real;
  reg        [15:0]   int_reg_array_10_58_imag;
  reg        [15:0]   int_reg_array_10_59_real;
  reg        [15:0]   int_reg_array_10_59_imag;
  reg        [15:0]   int_reg_array_10_60_real;
  reg        [15:0]   int_reg_array_10_60_imag;
  reg        [15:0]   int_reg_array_10_61_real;
  reg        [15:0]   int_reg_array_10_61_imag;
  reg        [15:0]   int_reg_array_10_62_real;
  reg        [15:0]   int_reg_array_10_62_imag;
  reg        [15:0]   int_reg_array_10_63_real;
  reg        [15:0]   int_reg_array_10_63_imag;
  reg        [15:0]   int_reg_array_55_0_real;
  reg        [15:0]   int_reg_array_55_0_imag;
  reg        [15:0]   int_reg_array_55_1_real;
  reg        [15:0]   int_reg_array_55_1_imag;
  reg        [15:0]   int_reg_array_55_2_real;
  reg        [15:0]   int_reg_array_55_2_imag;
  reg        [15:0]   int_reg_array_55_3_real;
  reg        [15:0]   int_reg_array_55_3_imag;
  reg        [15:0]   int_reg_array_55_4_real;
  reg        [15:0]   int_reg_array_55_4_imag;
  reg        [15:0]   int_reg_array_55_5_real;
  reg        [15:0]   int_reg_array_55_5_imag;
  reg        [15:0]   int_reg_array_55_6_real;
  reg        [15:0]   int_reg_array_55_6_imag;
  reg        [15:0]   int_reg_array_55_7_real;
  reg        [15:0]   int_reg_array_55_7_imag;
  reg        [15:0]   int_reg_array_55_8_real;
  reg        [15:0]   int_reg_array_55_8_imag;
  reg        [15:0]   int_reg_array_55_9_real;
  reg        [15:0]   int_reg_array_55_9_imag;
  reg        [15:0]   int_reg_array_55_10_real;
  reg        [15:0]   int_reg_array_55_10_imag;
  reg        [15:0]   int_reg_array_55_11_real;
  reg        [15:0]   int_reg_array_55_11_imag;
  reg        [15:0]   int_reg_array_55_12_real;
  reg        [15:0]   int_reg_array_55_12_imag;
  reg        [15:0]   int_reg_array_55_13_real;
  reg        [15:0]   int_reg_array_55_13_imag;
  reg        [15:0]   int_reg_array_55_14_real;
  reg        [15:0]   int_reg_array_55_14_imag;
  reg        [15:0]   int_reg_array_55_15_real;
  reg        [15:0]   int_reg_array_55_15_imag;
  reg        [15:0]   int_reg_array_55_16_real;
  reg        [15:0]   int_reg_array_55_16_imag;
  reg        [15:0]   int_reg_array_55_17_real;
  reg        [15:0]   int_reg_array_55_17_imag;
  reg        [15:0]   int_reg_array_55_18_real;
  reg        [15:0]   int_reg_array_55_18_imag;
  reg        [15:0]   int_reg_array_55_19_real;
  reg        [15:0]   int_reg_array_55_19_imag;
  reg        [15:0]   int_reg_array_55_20_real;
  reg        [15:0]   int_reg_array_55_20_imag;
  reg        [15:0]   int_reg_array_55_21_real;
  reg        [15:0]   int_reg_array_55_21_imag;
  reg        [15:0]   int_reg_array_55_22_real;
  reg        [15:0]   int_reg_array_55_22_imag;
  reg        [15:0]   int_reg_array_55_23_real;
  reg        [15:0]   int_reg_array_55_23_imag;
  reg        [15:0]   int_reg_array_55_24_real;
  reg        [15:0]   int_reg_array_55_24_imag;
  reg        [15:0]   int_reg_array_55_25_real;
  reg        [15:0]   int_reg_array_55_25_imag;
  reg        [15:0]   int_reg_array_55_26_real;
  reg        [15:0]   int_reg_array_55_26_imag;
  reg        [15:0]   int_reg_array_55_27_real;
  reg        [15:0]   int_reg_array_55_27_imag;
  reg        [15:0]   int_reg_array_55_28_real;
  reg        [15:0]   int_reg_array_55_28_imag;
  reg        [15:0]   int_reg_array_55_29_real;
  reg        [15:0]   int_reg_array_55_29_imag;
  reg        [15:0]   int_reg_array_55_30_real;
  reg        [15:0]   int_reg_array_55_30_imag;
  reg        [15:0]   int_reg_array_55_31_real;
  reg        [15:0]   int_reg_array_55_31_imag;
  reg        [15:0]   int_reg_array_55_32_real;
  reg        [15:0]   int_reg_array_55_32_imag;
  reg        [15:0]   int_reg_array_55_33_real;
  reg        [15:0]   int_reg_array_55_33_imag;
  reg        [15:0]   int_reg_array_55_34_real;
  reg        [15:0]   int_reg_array_55_34_imag;
  reg        [15:0]   int_reg_array_55_35_real;
  reg        [15:0]   int_reg_array_55_35_imag;
  reg        [15:0]   int_reg_array_55_36_real;
  reg        [15:0]   int_reg_array_55_36_imag;
  reg        [15:0]   int_reg_array_55_37_real;
  reg        [15:0]   int_reg_array_55_37_imag;
  reg        [15:0]   int_reg_array_55_38_real;
  reg        [15:0]   int_reg_array_55_38_imag;
  reg        [15:0]   int_reg_array_55_39_real;
  reg        [15:0]   int_reg_array_55_39_imag;
  reg        [15:0]   int_reg_array_55_40_real;
  reg        [15:0]   int_reg_array_55_40_imag;
  reg        [15:0]   int_reg_array_55_41_real;
  reg        [15:0]   int_reg_array_55_41_imag;
  reg        [15:0]   int_reg_array_55_42_real;
  reg        [15:0]   int_reg_array_55_42_imag;
  reg        [15:0]   int_reg_array_55_43_real;
  reg        [15:0]   int_reg_array_55_43_imag;
  reg        [15:0]   int_reg_array_55_44_real;
  reg        [15:0]   int_reg_array_55_44_imag;
  reg        [15:0]   int_reg_array_55_45_real;
  reg        [15:0]   int_reg_array_55_45_imag;
  reg        [15:0]   int_reg_array_55_46_real;
  reg        [15:0]   int_reg_array_55_46_imag;
  reg        [15:0]   int_reg_array_55_47_real;
  reg        [15:0]   int_reg_array_55_47_imag;
  reg        [15:0]   int_reg_array_55_48_real;
  reg        [15:0]   int_reg_array_55_48_imag;
  reg        [15:0]   int_reg_array_55_49_real;
  reg        [15:0]   int_reg_array_55_49_imag;
  reg        [15:0]   int_reg_array_55_50_real;
  reg        [15:0]   int_reg_array_55_50_imag;
  reg        [15:0]   int_reg_array_55_51_real;
  reg        [15:0]   int_reg_array_55_51_imag;
  reg        [15:0]   int_reg_array_55_52_real;
  reg        [15:0]   int_reg_array_55_52_imag;
  reg        [15:0]   int_reg_array_55_53_real;
  reg        [15:0]   int_reg_array_55_53_imag;
  reg        [15:0]   int_reg_array_55_54_real;
  reg        [15:0]   int_reg_array_55_54_imag;
  reg        [15:0]   int_reg_array_55_55_real;
  reg        [15:0]   int_reg_array_55_55_imag;
  reg        [15:0]   int_reg_array_55_56_real;
  reg        [15:0]   int_reg_array_55_56_imag;
  reg        [15:0]   int_reg_array_55_57_real;
  reg        [15:0]   int_reg_array_55_57_imag;
  reg        [15:0]   int_reg_array_55_58_real;
  reg        [15:0]   int_reg_array_55_58_imag;
  reg        [15:0]   int_reg_array_55_59_real;
  reg        [15:0]   int_reg_array_55_59_imag;
  reg        [15:0]   int_reg_array_55_60_real;
  reg        [15:0]   int_reg_array_55_60_imag;
  reg        [15:0]   int_reg_array_55_61_real;
  reg        [15:0]   int_reg_array_55_61_imag;
  reg        [15:0]   int_reg_array_55_62_real;
  reg        [15:0]   int_reg_array_55_62_imag;
  reg        [15:0]   int_reg_array_55_63_real;
  reg        [15:0]   int_reg_array_55_63_imag;
  reg        [15:0]   int_reg_array_25_0_real;
  reg        [15:0]   int_reg_array_25_0_imag;
  reg        [15:0]   int_reg_array_25_1_real;
  reg        [15:0]   int_reg_array_25_1_imag;
  reg        [15:0]   int_reg_array_25_2_real;
  reg        [15:0]   int_reg_array_25_2_imag;
  reg        [15:0]   int_reg_array_25_3_real;
  reg        [15:0]   int_reg_array_25_3_imag;
  reg        [15:0]   int_reg_array_25_4_real;
  reg        [15:0]   int_reg_array_25_4_imag;
  reg        [15:0]   int_reg_array_25_5_real;
  reg        [15:0]   int_reg_array_25_5_imag;
  reg        [15:0]   int_reg_array_25_6_real;
  reg        [15:0]   int_reg_array_25_6_imag;
  reg        [15:0]   int_reg_array_25_7_real;
  reg        [15:0]   int_reg_array_25_7_imag;
  reg        [15:0]   int_reg_array_25_8_real;
  reg        [15:0]   int_reg_array_25_8_imag;
  reg        [15:0]   int_reg_array_25_9_real;
  reg        [15:0]   int_reg_array_25_9_imag;
  reg        [15:0]   int_reg_array_25_10_real;
  reg        [15:0]   int_reg_array_25_10_imag;
  reg        [15:0]   int_reg_array_25_11_real;
  reg        [15:0]   int_reg_array_25_11_imag;
  reg        [15:0]   int_reg_array_25_12_real;
  reg        [15:0]   int_reg_array_25_12_imag;
  reg        [15:0]   int_reg_array_25_13_real;
  reg        [15:0]   int_reg_array_25_13_imag;
  reg        [15:0]   int_reg_array_25_14_real;
  reg        [15:0]   int_reg_array_25_14_imag;
  reg        [15:0]   int_reg_array_25_15_real;
  reg        [15:0]   int_reg_array_25_15_imag;
  reg        [15:0]   int_reg_array_25_16_real;
  reg        [15:0]   int_reg_array_25_16_imag;
  reg        [15:0]   int_reg_array_25_17_real;
  reg        [15:0]   int_reg_array_25_17_imag;
  reg        [15:0]   int_reg_array_25_18_real;
  reg        [15:0]   int_reg_array_25_18_imag;
  reg        [15:0]   int_reg_array_25_19_real;
  reg        [15:0]   int_reg_array_25_19_imag;
  reg        [15:0]   int_reg_array_25_20_real;
  reg        [15:0]   int_reg_array_25_20_imag;
  reg        [15:0]   int_reg_array_25_21_real;
  reg        [15:0]   int_reg_array_25_21_imag;
  reg        [15:0]   int_reg_array_25_22_real;
  reg        [15:0]   int_reg_array_25_22_imag;
  reg        [15:0]   int_reg_array_25_23_real;
  reg        [15:0]   int_reg_array_25_23_imag;
  reg        [15:0]   int_reg_array_25_24_real;
  reg        [15:0]   int_reg_array_25_24_imag;
  reg        [15:0]   int_reg_array_25_25_real;
  reg        [15:0]   int_reg_array_25_25_imag;
  reg        [15:0]   int_reg_array_25_26_real;
  reg        [15:0]   int_reg_array_25_26_imag;
  reg        [15:0]   int_reg_array_25_27_real;
  reg        [15:0]   int_reg_array_25_27_imag;
  reg        [15:0]   int_reg_array_25_28_real;
  reg        [15:0]   int_reg_array_25_28_imag;
  reg        [15:0]   int_reg_array_25_29_real;
  reg        [15:0]   int_reg_array_25_29_imag;
  reg        [15:0]   int_reg_array_25_30_real;
  reg        [15:0]   int_reg_array_25_30_imag;
  reg        [15:0]   int_reg_array_25_31_real;
  reg        [15:0]   int_reg_array_25_31_imag;
  reg        [15:0]   int_reg_array_25_32_real;
  reg        [15:0]   int_reg_array_25_32_imag;
  reg        [15:0]   int_reg_array_25_33_real;
  reg        [15:0]   int_reg_array_25_33_imag;
  reg        [15:0]   int_reg_array_25_34_real;
  reg        [15:0]   int_reg_array_25_34_imag;
  reg        [15:0]   int_reg_array_25_35_real;
  reg        [15:0]   int_reg_array_25_35_imag;
  reg        [15:0]   int_reg_array_25_36_real;
  reg        [15:0]   int_reg_array_25_36_imag;
  reg        [15:0]   int_reg_array_25_37_real;
  reg        [15:0]   int_reg_array_25_37_imag;
  reg        [15:0]   int_reg_array_25_38_real;
  reg        [15:0]   int_reg_array_25_38_imag;
  reg        [15:0]   int_reg_array_25_39_real;
  reg        [15:0]   int_reg_array_25_39_imag;
  reg        [15:0]   int_reg_array_25_40_real;
  reg        [15:0]   int_reg_array_25_40_imag;
  reg        [15:0]   int_reg_array_25_41_real;
  reg        [15:0]   int_reg_array_25_41_imag;
  reg        [15:0]   int_reg_array_25_42_real;
  reg        [15:0]   int_reg_array_25_42_imag;
  reg        [15:0]   int_reg_array_25_43_real;
  reg        [15:0]   int_reg_array_25_43_imag;
  reg        [15:0]   int_reg_array_25_44_real;
  reg        [15:0]   int_reg_array_25_44_imag;
  reg        [15:0]   int_reg_array_25_45_real;
  reg        [15:0]   int_reg_array_25_45_imag;
  reg        [15:0]   int_reg_array_25_46_real;
  reg        [15:0]   int_reg_array_25_46_imag;
  reg        [15:0]   int_reg_array_25_47_real;
  reg        [15:0]   int_reg_array_25_47_imag;
  reg        [15:0]   int_reg_array_25_48_real;
  reg        [15:0]   int_reg_array_25_48_imag;
  reg        [15:0]   int_reg_array_25_49_real;
  reg        [15:0]   int_reg_array_25_49_imag;
  reg        [15:0]   int_reg_array_25_50_real;
  reg        [15:0]   int_reg_array_25_50_imag;
  reg        [15:0]   int_reg_array_25_51_real;
  reg        [15:0]   int_reg_array_25_51_imag;
  reg        [15:0]   int_reg_array_25_52_real;
  reg        [15:0]   int_reg_array_25_52_imag;
  reg        [15:0]   int_reg_array_25_53_real;
  reg        [15:0]   int_reg_array_25_53_imag;
  reg        [15:0]   int_reg_array_25_54_real;
  reg        [15:0]   int_reg_array_25_54_imag;
  reg        [15:0]   int_reg_array_25_55_real;
  reg        [15:0]   int_reg_array_25_55_imag;
  reg        [15:0]   int_reg_array_25_56_real;
  reg        [15:0]   int_reg_array_25_56_imag;
  reg        [15:0]   int_reg_array_25_57_real;
  reg        [15:0]   int_reg_array_25_57_imag;
  reg        [15:0]   int_reg_array_25_58_real;
  reg        [15:0]   int_reg_array_25_58_imag;
  reg        [15:0]   int_reg_array_25_59_real;
  reg        [15:0]   int_reg_array_25_59_imag;
  reg        [15:0]   int_reg_array_25_60_real;
  reg        [15:0]   int_reg_array_25_60_imag;
  reg        [15:0]   int_reg_array_25_61_real;
  reg        [15:0]   int_reg_array_25_61_imag;
  reg        [15:0]   int_reg_array_25_62_real;
  reg        [15:0]   int_reg_array_25_62_imag;
  reg        [15:0]   int_reg_array_25_63_real;
  reg        [15:0]   int_reg_array_25_63_imag;
  reg        [15:0]   int_reg_array_39_0_real;
  reg        [15:0]   int_reg_array_39_0_imag;
  reg        [15:0]   int_reg_array_39_1_real;
  reg        [15:0]   int_reg_array_39_1_imag;
  reg        [15:0]   int_reg_array_39_2_real;
  reg        [15:0]   int_reg_array_39_2_imag;
  reg        [15:0]   int_reg_array_39_3_real;
  reg        [15:0]   int_reg_array_39_3_imag;
  reg        [15:0]   int_reg_array_39_4_real;
  reg        [15:0]   int_reg_array_39_4_imag;
  reg        [15:0]   int_reg_array_39_5_real;
  reg        [15:0]   int_reg_array_39_5_imag;
  reg        [15:0]   int_reg_array_39_6_real;
  reg        [15:0]   int_reg_array_39_6_imag;
  reg        [15:0]   int_reg_array_39_7_real;
  reg        [15:0]   int_reg_array_39_7_imag;
  reg        [15:0]   int_reg_array_39_8_real;
  reg        [15:0]   int_reg_array_39_8_imag;
  reg        [15:0]   int_reg_array_39_9_real;
  reg        [15:0]   int_reg_array_39_9_imag;
  reg        [15:0]   int_reg_array_39_10_real;
  reg        [15:0]   int_reg_array_39_10_imag;
  reg        [15:0]   int_reg_array_39_11_real;
  reg        [15:0]   int_reg_array_39_11_imag;
  reg        [15:0]   int_reg_array_39_12_real;
  reg        [15:0]   int_reg_array_39_12_imag;
  reg        [15:0]   int_reg_array_39_13_real;
  reg        [15:0]   int_reg_array_39_13_imag;
  reg        [15:0]   int_reg_array_39_14_real;
  reg        [15:0]   int_reg_array_39_14_imag;
  reg        [15:0]   int_reg_array_39_15_real;
  reg        [15:0]   int_reg_array_39_15_imag;
  reg        [15:0]   int_reg_array_39_16_real;
  reg        [15:0]   int_reg_array_39_16_imag;
  reg        [15:0]   int_reg_array_39_17_real;
  reg        [15:0]   int_reg_array_39_17_imag;
  reg        [15:0]   int_reg_array_39_18_real;
  reg        [15:0]   int_reg_array_39_18_imag;
  reg        [15:0]   int_reg_array_39_19_real;
  reg        [15:0]   int_reg_array_39_19_imag;
  reg        [15:0]   int_reg_array_39_20_real;
  reg        [15:0]   int_reg_array_39_20_imag;
  reg        [15:0]   int_reg_array_39_21_real;
  reg        [15:0]   int_reg_array_39_21_imag;
  reg        [15:0]   int_reg_array_39_22_real;
  reg        [15:0]   int_reg_array_39_22_imag;
  reg        [15:0]   int_reg_array_39_23_real;
  reg        [15:0]   int_reg_array_39_23_imag;
  reg        [15:0]   int_reg_array_39_24_real;
  reg        [15:0]   int_reg_array_39_24_imag;
  reg        [15:0]   int_reg_array_39_25_real;
  reg        [15:0]   int_reg_array_39_25_imag;
  reg        [15:0]   int_reg_array_39_26_real;
  reg        [15:0]   int_reg_array_39_26_imag;
  reg        [15:0]   int_reg_array_39_27_real;
  reg        [15:0]   int_reg_array_39_27_imag;
  reg        [15:0]   int_reg_array_39_28_real;
  reg        [15:0]   int_reg_array_39_28_imag;
  reg        [15:0]   int_reg_array_39_29_real;
  reg        [15:0]   int_reg_array_39_29_imag;
  reg        [15:0]   int_reg_array_39_30_real;
  reg        [15:0]   int_reg_array_39_30_imag;
  reg        [15:0]   int_reg_array_39_31_real;
  reg        [15:0]   int_reg_array_39_31_imag;
  reg        [15:0]   int_reg_array_39_32_real;
  reg        [15:0]   int_reg_array_39_32_imag;
  reg        [15:0]   int_reg_array_39_33_real;
  reg        [15:0]   int_reg_array_39_33_imag;
  reg        [15:0]   int_reg_array_39_34_real;
  reg        [15:0]   int_reg_array_39_34_imag;
  reg        [15:0]   int_reg_array_39_35_real;
  reg        [15:0]   int_reg_array_39_35_imag;
  reg        [15:0]   int_reg_array_39_36_real;
  reg        [15:0]   int_reg_array_39_36_imag;
  reg        [15:0]   int_reg_array_39_37_real;
  reg        [15:0]   int_reg_array_39_37_imag;
  reg        [15:0]   int_reg_array_39_38_real;
  reg        [15:0]   int_reg_array_39_38_imag;
  reg        [15:0]   int_reg_array_39_39_real;
  reg        [15:0]   int_reg_array_39_39_imag;
  reg        [15:0]   int_reg_array_39_40_real;
  reg        [15:0]   int_reg_array_39_40_imag;
  reg        [15:0]   int_reg_array_39_41_real;
  reg        [15:0]   int_reg_array_39_41_imag;
  reg        [15:0]   int_reg_array_39_42_real;
  reg        [15:0]   int_reg_array_39_42_imag;
  reg        [15:0]   int_reg_array_39_43_real;
  reg        [15:0]   int_reg_array_39_43_imag;
  reg        [15:0]   int_reg_array_39_44_real;
  reg        [15:0]   int_reg_array_39_44_imag;
  reg        [15:0]   int_reg_array_39_45_real;
  reg        [15:0]   int_reg_array_39_45_imag;
  reg        [15:0]   int_reg_array_39_46_real;
  reg        [15:0]   int_reg_array_39_46_imag;
  reg        [15:0]   int_reg_array_39_47_real;
  reg        [15:0]   int_reg_array_39_47_imag;
  reg        [15:0]   int_reg_array_39_48_real;
  reg        [15:0]   int_reg_array_39_48_imag;
  reg        [15:0]   int_reg_array_39_49_real;
  reg        [15:0]   int_reg_array_39_49_imag;
  reg        [15:0]   int_reg_array_39_50_real;
  reg        [15:0]   int_reg_array_39_50_imag;
  reg        [15:0]   int_reg_array_39_51_real;
  reg        [15:0]   int_reg_array_39_51_imag;
  reg        [15:0]   int_reg_array_39_52_real;
  reg        [15:0]   int_reg_array_39_52_imag;
  reg        [15:0]   int_reg_array_39_53_real;
  reg        [15:0]   int_reg_array_39_53_imag;
  reg        [15:0]   int_reg_array_39_54_real;
  reg        [15:0]   int_reg_array_39_54_imag;
  reg        [15:0]   int_reg_array_39_55_real;
  reg        [15:0]   int_reg_array_39_55_imag;
  reg        [15:0]   int_reg_array_39_56_real;
  reg        [15:0]   int_reg_array_39_56_imag;
  reg        [15:0]   int_reg_array_39_57_real;
  reg        [15:0]   int_reg_array_39_57_imag;
  reg        [15:0]   int_reg_array_39_58_real;
  reg        [15:0]   int_reg_array_39_58_imag;
  reg        [15:0]   int_reg_array_39_59_real;
  reg        [15:0]   int_reg_array_39_59_imag;
  reg        [15:0]   int_reg_array_39_60_real;
  reg        [15:0]   int_reg_array_39_60_imag;
  reg        [15:0]   int_reg_array_39_61_real;
  reg        [15:0]   int_reg_array_39_61_imag;
  reg        [15:0]   int_reg_array_39_62_real;
  reg        [15:0]   int_reg_array_39_62_imag;
  reg        [15:0]   int_reg_array_39_63_real;
  reg        [15:0]   int_reg_array_39_63_imag;
  reg        [15:0]   int_reg_array_13_0_real;
  reg        [15:0]   int_reg_array_13_0_imag;
  reg        [15:0]   int_reg_array_13_1_real;
  reg        [15:0]   int_reg_array_13_1_imag;
  reg        [15:0]   int_reg_array_13_2_real;
  reg        [15:0]   int_reg_array_13_2_imag;
  reg        [15:0]   int_reg_array_13_3_real;
  reg        [15:0]   int_reg_array_13_3_imag;
  reg        [15:0]   int_reg_array_13_4_real;
  reg        [15:0]   int_reg_array_13_4_imag;
  reg        [15:0]   int_reg_array_13_5_real;
  reg        [15:0]   int_reg_array_13_5_imag;
  reg        [15:0]   int_reg_array_13_6_real;
  reg        [15:0]   int_reg_array_13_6_imag;
  reg        [15:0]   int_reg_array_13_7_real;
  reg        [15:0]   int_reg_array_13_7_imag;
  reg        [15:0]   int_reg_array_13_8_real;
  reg        [15:0]   int_reg_array_13_8_imag;
  reg        [15:0]   int_reg_array_13_9_real;
  reg        [15:0]   int_reg_array_13_9_imag;
  reg        [15:0]   int_reg_array_13_10_real;
  reg        [15:0]   int_reg_array_13_10_imag;
  reg        [15:0]   int_reg_array_13_11_real;
  reg        [15:0]   int_reg_array_13_11_imag;
  reg        [15:0]   int_reg_array_13_12_real;
  reg        [15:0]   int_reg_array_13_12_imag;
  reg        [15:0]   int_reg_array_13_13_real;
  reg        [15:0]   int_reg_array_13_13_imag;
  reg        [15:0]   int_reg_array_13_14_real;
  reg        [15:0]   int_reg_array_13_14_imag;
  reg        [15:0]   int_reg_array_13_15_real;
  reg        [15:0]   int_reg_array_13_15_imag;
  reg        [15:0]   int_reg_array_13_16_real;
  reg        [15:0]   int_reg_array_13_16_imag;
  reg        [15:0]   int_reg_array_13_17_real;
  reg        [15:0]   int_reg_array_13_17_imag;
  reg        [15:0]   int_reg_array_13_18_real;
  reg        [15:0]   int_reg_array_13_18_imag;
  reg        [15:0]   int_reg_array_13_19_real;
  reg        [15:0]   int_reg_array_13_19_imag;
  reg        [15:0]   int_reg_array_13_20_real;
  reg        [15:0]   int_reg_array_13_20_imag;
  reg        [15:0]   int_reg_array_13_21_real;
  reg        [15:0]   int_reg_array_13_21_imag;
  reg        [15:0]   int_reg_array_13_22_real;
  reg        [15:0]   int_reg_array_13_22_imag;
  reg        [15:0]   int_reg_array_13_23_real;
  reg        [15:0]   int_reg_array_13_23_imag;
  reg        [15:0]   int_reg_array_13_24_real;
  reg        [15:0]   int_reg_array_13_24_imag;
  reg        [15:0]   int_reg_array_13_25_real;
  reg        [15:0]   int_reg_array_13_25_imag;
  reg        [15:0]   int_reg_array_13_26_real;
  reg        [15:0]   int_reg_array_13_26_imag;
  reg        [15:0]   int_reg_array_13_27_real;
  reg        [15:0]   int_reg_array_13_27_imag;
  reg        [15:0]   int_reg_array_13_28_real;
  reg        [15:0]   int_reg_array_13_28_imag;
  reg        [15:0]   int_reg_array_13_29_real;
  reg        [15:0]   int_reg_array_13_29_imag;
  reg        [15:0]   int_reg_array_13_30_real;
  reg        [15:0]   int_reg_array_13_30_imag;
  reg        [15:0]   int_reg_array_13_31_real;
  reg        [15:0]   int_reg_array_13_31_imag;
  reg        [15:0]   int_reg_array_13_32_real;
  reg        [15:0]   int_reg_array_13_32_imag;
  reg        [15:0]   int_reg_array_13_33_real;
  reg        [15:0]   int_reg_array_13_33_imag;
  reg        [15:0]   int_reg_array_13_34_real;
  reg        [15:0]   int_reg_array_13_34_imag;
  reg        [15:0]   int_reg_array_13_35_real;
  reg        [15:0]   int_reg_array_13_35_imag;
  reg        [15:0]   int_reg_array_13_36_real;
  reg        [15:0]   int_reg_array_13_36_imag;
  reg        [15:0]   int_reg_array_13_37_real;
  reg        [15:0]   int_reg_array_13_37_imag;
  reg        [15:0]   int_reg_array_13_38_real;
  reg        [15:0]   int_reg_array_13_38_imag;
  reg        [15:0]   int_reg_array_13_39_real;
  reg        [15:0]   int_reg_array_13_39_imag;
  reg        [15:0]   int_reg_array_13_40_real;
  reg        [15:0]   int_reg_array_13_40_imag;
  reg        [15:0]   int_reg_array_13_41_real;
  reg        [15:0]   int_reg_array_13_41_imag;
  reg        [15:0]   int_reg_array_13_42_real;
  reg        [15:0]   int_reg_array_13_42_imag;
  reg        [15:0]   int_reg_array_13_43_real;
  reg        [15:0]   int_reg_array_13_43_imag;
  reg        [15:0]   int_reg_array_13_44_real;
  reg        [15:0]   int_reg_array_13_44_imag;
  reg        [15:0]   int_reg_array_13_45_real;
  reg        [15:0]   int_reg_array_13_45_imag;
  reg        [15:0]   int_reg_array_13_46_real;
  reg        [15:0]   int_reg_array_13_46_imag;
  reg        [15:0]   int_reg_array_13_47_real;
  reg        [15:0]   int_reg_array_13_47_imag;
  reg        [15:0]   int_reg_array_13_48_real;
  reg        [15:0]   int_reg_array_13_48_imag;
  reg        [15:0]   int_reg_array_13_49_real;
  reg        [15:0]   int_reg_array_13_49_imag;
  reg        [15:0]   int_reg_array_13_50_real;
  reg        [15:0]   int_reg_array_13_50_imag;
  reg        [15:0]   int_reg_array_13_51_real;
  reg        [15:0]   int_reg_array_13_51_imag;
  reg        [15:0]   int_reg_array_13_52_real;
  reg        [15:0]   int_reg_array_13_52_imag;
  reg        [15:0]   int_reg_array_13_53_real;
  reg        [15:0]   int_reg_array_13_53_imag;
  reg        [15:0]   int_reg_array_13_54_real;
  reg        [15:0]   int_reg_array_13_54_imag;
  reg        [15:0]   int_reg_array_13_55_real;
  reg        [15:0]   int_reg_array_13_55_imag;
  reg        [15:0]   int_reg_array_13_56_real;
  reg        [15:0]   int_reg_array_13_56_imag;
  reg        [15:0]   int_reg_array_13_57_real;
  reg        [15:0]   int_reg_array_13_57_imag;
  reg        [15:0]   int_reg_array_13_58_real;
  reg        [15:0]   int_reg_array_13_58_imag;
  reg        [15:0]   int_reg_array_13_59_real;
  reg        [15:0]   int_reg_array_13_59_imag;
  reg        [15:0]   int_reg_array_13_60_real;
  reg        [15:0]   int_reg_array_13_60_imag;
  reg        [15:0]   int_reg_array_13_61_real;
  reg        [15:0]   int_reg_array_13_61_imag;
  reg        [15:0]   int_reg_array_13_62_real;
  reg        [15:0]   int_reg_array_13_62_imag;
  reg        [15:0]   int_reg_array_13_63_real;
  reg        [15:0]   int_reg_array_13_63_imag;
  reg        [15:0]   int_reg_array_53_0_real;
  reg        [15:0]   int_reg_array_53_0_imag;
  reg        [15:0]   int_reg_array_53_1_real;
  reg        [15:0]   int_reg_array_53_1_imag;
  reg        [15:0]   int_reg_array_53_2_real;
  reg        [15:0]   int_reg_array_53_2_imag;
  reg        [15:0]   int_reg_array_53_3_real;
  reg        [15:0]   int_reg_array_53_3_imag;
  reg        [15:0]   int_reg_array_53_4_real;
  reg        [15:0]   int_reg_array_53_4_imag;
  reg        [15:0]   int_reg_array_53_5_real;
  reg        [15:0]   int_reg_array_53_5_imag;
  reg        [15:0]   int_reg_array_53_6_real;
  reg        [15:0]   int_reg_array_53_6_imag;
  reg        [15:0]   int_reg_array_53_7_real;
  reg        [15:0]   int_reg_array_53_7_imag;
  reg        [15:0]   int_reg_array_53_8_real;
  reg        [15:0]   int_reg_array_53_8_imag;
  reg        [15:0]   int_reg_array_53_9_real;
  reg        [15:0]   int_reg_array_53_9_imag;
  reg        [15:0]   int_reg_array_53_10_real;
  reg        [15:0]   int_reg_array_53_10_imag;
  reg        [15:0]   int_reg_array_53_11_real;
  reg        [15:0]   int_reg_array_53_11_imag;
  reg        [15:0]   int_reg_array_53_12_real;
  reg        [15:0]   int_reg_array_53_12_imag;
  reg        [15:0]   int_reg_array_53_13_real;
  reg        [15:0]   int_reg_array_53_13_imag;
  reg        [15:0]   int_reg_array_53_14_real;
  reg        [15:0]   int_reg_array_53_14_imag;
  reg        [15:0]   int_reg_array_53_15_real;
  reg        [15:0]   int_reg_array_53_15_imag;
  reg        [15:0]   int_reg_array_53_16_real;
  reg        [15:0]   int_reg_array_53_16_imag;
  reg        [15:0]   int_reg_array_53_17_real;
  reg        [15:0]   int_reg_array_53_17_imag;
  reg        [15:0]   int_reg_array_53_18_real;
  reg        [15:0]   int_reg_array_53_18_imag;
  reg        [15:0]   int_reg_array_53_19_real;
  reg        [15:0]   int_reg_array_53_19_imag;
  reg        [15:0]   int_reg_array_53_20_real;
  reg        [15:0]   int_reg_array_53_20_imag;
  reg        [15:0]   int_reg_array_53_21_real;
  reg        [15:0]   int_reg_array_53_21_imag;
  reg        [15:0]   int_reg_array_53_22_real;
  reg        [15:0]   int_reg_array_53_22_imag;
  reg        [15:0]   int_reg_array_53_23_real;
  reg        [15:0]   int_reg_array_53_23_imag;
  reg        [15:0]   int_reg_array_53_24_real;
  reg        [15:0]   int_reg_array_53_24_imag;
  reg        [15:0]   int_reg_array_53_25_real;
  reg        [15:0]   int_reg_array_53_25_imag;
  reg        [15:0]   int_reg_array_53_26_real;
  reg        [15:0]   int_reg_array_53_26_imag;
  reg        [15:0]   int_reg_array_53_27_real;
  reg        [15:0]   int_reg_array_53_27_imag;
  reg        [15:0]   int_reg_array_53_28_real;
  reg        [15:0]   int_reg_array_53_28_imag;
  reg        [15:0]   int_reg_array_53_29_real;
  reg        [15:0]   int_reg_array_53_29_imag;
  reg        [15:0]   int_reg_array_53_30_real;
  reg        [15:0]   int_reg_array_53_30_imag;
  reg        [15:0]   int_reg_array_53_31_real;
  reg        [15:0]   int_reg_array_53_31_imag;
  reg        [15:0]   int_reg_array_53_32_real;
  reg        [15:0]   int_reg_array_53_32_imag;
  reg        [15:0]   int_reg_array_53_33_real;
  reg        [15:0]   int_reg_array_53_33_imag;
  reg        [15:0]   int_reg_array_53_34_real;
  reg        [15:0]   int_reg_array_53_34_imag;
  reg        [15:0]   int_reg_array_53_35_real;
  reg        [15:0]   int_reg_array_53_35_imag;
  reg        [15:0]   int_reg_array_53_36_real;
  reg        [15:0]   int_reg_array_53_36_imag;
  reg        [15:0]   int_reg_array_53_37_real;
  reg        [15:0]   int_reg_array_53_37_imag;
  reg        [15:0]   int_reg_array_53_38_real;
  reg        [15:0]   int_reg_array_53_38_imag;
  reg        [15:0]   int_reg_array_53_39_real;
  reg        [15:0]   int_reg_array_53_39_imag;
  reg        [15:0]   int_reg_array_53_40_real;
  reg        [15:0]   int_reg_array_53_40_imag;
  reg        [15:0]   int_reg_array_53_41_real;
  reg        [15:0]   int_reg_array_53_41_imag;
  reg        [15:0]   int_reg_array_53_42_real;
  reg        [15:0]   int_reg_array_53_42_imag;
  reg        [15:0]   int_reg_array_53_43_real;
  reg        [15:0]   int_reg_array_53_43_imag;
  reg        [15:0]   int_reg_array_53_44_real;
  reg        [15:0]   int_reg_array_53_44_imag;
  reg        [15:0]   int_reg_array_53_45_real;
  reg        [15:0]   int_reg_array_53_45_imag;
  reg        [15:0]   int_reg_array_53_46_real;
  reg        [15:0]   int_reg_array_53_46_imag;
  reg        [15:0]   int_reg_array_53_47_real;
  reg        [15:0]   int_reg_array_53_47_imag;
  reg        [15:0]   int_reg_array_53_48_real;
  reg        [15:0]   int_reg_array_53_48_imag;
  reg        [15:0]   int_reg_array_53_49_real;
  reg        [15:0]   int_reg_array_53_49_imag;
  reg        [15:0]   int_reg_array_53_50_real;
  reg        [15:0]   int_reg_array_53_50_imag;
  reg        [15:0]   int_reg_array_53_51_real;
  reg        [15:0]   int_reg_array_53_51_imag;
  reg        [15:0]   int_reg_array_53_52_real;
  reg        [15:0]   int_reg_array_53_52_imag;
  reg        [15:0]   int_reg_array_53_53_real;
  reg        [15:0]   int_reg_array_53_53_imag;
  reg        [15:0]   int_reg_array_53_54_real;
  reg        [15:0]   int_reg_array_53_54_imag;
  reg        [15:0]   int_reg_array_53_55_real;
  reg        [15:0]   int_reg_array_53_55_imag;
  reg        [15:0]   int_reg_array_53_56_real;
  reg        [15:0]   int_reg_array_53_56_imag;
  reg        [15:0]   int_reg_array_53_57_real;
  reg        [15:0]   int_reg_array_53_57_imag;
  reg        [15:0]   int_reg_array_53_58_real;
  reg        [15:0]   int_reg_array_53_58_imag;
  reg        [15:0]   int_reg_array_53_59_real;
  reg        [15:0]   int_reg_array_53_59_imag;
  reg        [15:0]   int_reg_array_53_60_real;
  reg        [15:0]   int_reg_array_53_60_imag;
  reg        [15:0]   int_reg_array_53_61_real;
  reg        [15:0]   int_reg_array_53_61_imag;
  reg        [15:0]   int_reg_array_53_62_real;
  reg        [15:0]   int_reg_array_53_62_imag;
  reg        [15:0]   int_reg_array_53_63_real;
  reg        [15:0]   int_reg_array_53_63_imag;
  reg        [15:0]   int_reg_array_59_0_real;
  reg        [15:0]   int_reg_array_59_0_imag;
  reg        [15:0]   int_reg_array_59_1_real;
  reg        [15:0]   int_reg_array_59_1_imag;
  reg        [15:0]   int_reg_array_59_2_real;
  reg        [15:0]   int_reg_array_59_2_imag;
  reg        [15:0]   int_reg_array_59_3_real;
  reg        [15:0]   int_reg_array_59_3_imag;
  reg        [15:0]   int_reg_array_59_4_real;
  reg        [15:0]   int_reg_array_59_4_imag;
  reg        [15:0]   int_reg_array_59_5_real;
  reg        [15:0]   int_reg_array_59_5_imag;
  reg        [15:0]   int_reg_array_59_6_real;
  reg        [15:0]   int_reg_array_59_6_imag;
  reg        [15:0]   int_reg_array_59_7_real;
  reg        [15:0]   int_reg_array_59_7_imag;
  reg        [15:0]   int_reg_array_59_8_real;
  reg        [15:0]   int_reg_array_59_8_imag;
  reg        [15:0]   int_reg_array_59_9_real;
  reg        [15:0]   int_reg_array_59_9_imag;
  reg        [15:0]   int_reg_array_59_10_real;
  reg        [15:0]   int_reg_array_59_10_imag;
  reg        [15:0]   int_reg_array_59_11_real;
  reg        [15:0]   int_reg_array_59_11_imag;
  reg        [15:0]   int_reg_array_59_12_real;
  reg        [15:0]   int_reg_array_59_12_imag;
  reg        [15:0]   int_reg_array_59_13_real;
  reg        [15:0]   int_reg_array_59_13_imag;
  reg        [15:0]   int_reg_array_59_14_real;
  reg        [15:0]   int_reg_array_59_14_imag;
  reg        [15:0]   int_reg_array_59_15_real;
  reg        [15:0]   int_reg_array_59_15_imag;
  reg        [15:0]   int_reg_array_59_16_real;
  reg        [15:0]   int_reg_array_59_16_imag;
  reg        [15:0]   int_reg_array_59_17_real;
  reg        [15:0]   int_reg_array_59_17_imag;
  reg        [15:0]   int_reg_array_59_18_real;
  reg        [15:0]   int_reg_array_59_18_imag;
  reg        [15:0]   int_reg_array_59_19_real;
  reg        [15:0]   int_reg_array_59_19_imag;
  reg        [15:0]   int_reg_array_59_20_real;
  reg        [15:0]   int_reg_array_59_20_imag;
  reg        [15:0]   int_reg_array_59_21_real;
  reg        [15:0]   int_reg_array_59_21_imag;
  reg        [15:0]   int_reg_array_59_22_real;
  reg        [15:0]   int_reg_array_59_22_imag;
  reg        [15:0]   int_reg_array_59_23_real;
  reg        [15:0]   int_reg_array_59_23_imag;
  reg        [15:0]   int_reg_array_59_24_real;
  reg        [15:0]   int_reg_array_59_24_imag;
  reg        [15:0]   int_reg_array_59_25_real;
  reg        [15:0]   int_reg_array_59_25_imag;
  reg        [15:0]   int_reg_array_59_26_real;
  reg        [15:0]   int_reg_array_59_26_imag;
  reg        [15:0]   int_reg_array_59_27_real;
  reg        [15:0]   int_reg_array_59_27_imag;
  reg        [15:0]   int_reg_array_59_28_real;
  reg        [15:0]   int_reg_array_59_28_imag;
  reg        [15:0]   int_reg_array_59_29_real;
  reg        [15:0]   int_reg_array_59_29_imag;
  reg        [15:0]   int_reg_array_59_30_real;
  reg        [15:0]   int_reg_array_59_30_imag;
  reg        [15:0]   int_reg_array_59_31_real;
  reg        [15:0]   int_reg_array_59_31_imag;
  reg        [15:0]   int_reg_array_59_32_real;
  reg        [15:0]   int_reg_array_59_32_imag;
  reg        [15:0]   int_reg_array_59_33_real;
  reg        [15:0]   int_reg_array_59_33_imag;
  reg        [15:0]   int_reg_array_59_34_real;
  reg        [15:0]   int_reg_array_59_34_imag;
  reg        [15:0]   int_reg_array_59_35_real;
  reg        [15:0]   int_reg_array_59_35_imag;
  reg        [15:0]   int_reg_array_59_36_real;
  reg        [15:0]   int_reg_array_59_36_imag;
  reg        [15:0]   int_reg_array_59_37_real;
  reg        [15:0]   int_reg_array_59_37_imag;
  reg        [15:0]   int_reg_array_59_38_real;
  reg        [15:0]   int_reg_array_59_38_imag;
  reg        [15:0]   int_reg_array_59_39_real;
  reg        [15:0]   int_reg_array_59_39_imag;
  reg        [15:0]   int_reg_array_59_40_real;
  reg        [15:0]   int_reg_array_59_40_imag;
  reg        [15:0]   int_reg_array_59_41_real;
  reg        [15:0]   int_reg_array_59_41_imag;
  reg        [15:0]   int_reg_array_59_42_real;
  reg        [15:0]   int_reg_array_59_42_imag;
  reg        [15:0]   int_reg_array_59_43_real;
  reg        [15:0]   int_reg_array_59_43_imag;
  reg        [15:0]   int_reg_array_59_44_real;
  reg        [15:0]   int_reg_array_59_44_imag;
  reg        [15:0]   int_reg_array_59_45_real;
  reg        [15:0]   int_reg_array_59_45_imag;
  reg        [15:0]   int_reg_array_59_46_real;
  reg        [15:0]   int_reg_array_59_46_imag;
  reg        [15:0]   int_reg_array_59_47_real;
  reg        [15:0]   int_reg_array_59_47_imag;
  reg        [15:0]   int_reg_array_59_48_real;
  reg        [15:0]   int_reg_array_59_48_imag;
  reg        [15:0]   int_reg_array_59_49_real;
  reg        [15:0]   int_reg_array_59_49_imag;
  reg        [15:0]   int_reg_array_59_50_real;
  reg        [15:0]   int_reg_array_59_50_imag;
  reg        [15:0]   int_reg_array_59_51_real;
  reg        [15:0]   int_reg_array_59_51_imag;
  reg        [15:0]   int_reg_array_59_52_real;
  reg        [15:0]   int_reg_array_59_52_imag;
  reg        [15:0]   int_reg_array_59_53_real;
  reg        [15:0]   int_reg_array_59_53_imag;
  reg        [15:0]   int_reg_array_59_54_real;
  reg        [15:0]   int_reg_array_59_54_imag;
  reg        [15:0]   int_reg_array_59_55_real;
  reg        [15:0]   int_reg_array_59_55_imag;
  reg        [15:0]   int_reg_array_59_56_real;
  reg        [15:0]   int_reg_array_59_56_imag;
  reg        [15:0]   int_reg_array_59_57_real;
  reg        [15:0]   int_reg_array_59_57_imag;
  reg        [15:0]   int_reg_array_59_58_real;
  reg        [15:0]   int_reg_array_59_58_imag;
  reg        [15:0]   int_reg_array_59_59_real;
  reg        [15:0]   int_reg_array_59_59_imag;
  reg        [15:0]   int_reg_array_59_60_real;
  reg        [15:0]   int_reg_array_59_60_imag;
  reg        [15:0]   int_reg_array_59_61_real;
  reg        [15:0]   int_reg_array_59_61_imag;
  reg        [15:0]   int_reg_array_59_62_real;
  reg        [15:0]   int_reg_array_59_62_imag;
  reg        [15:0]   int_reg_array_59_63_real;
  reg        [15:0]   int_reg_array_59_63_imag;
  reg        [15:0]   int_reg_array_57_0_real;
  reg        [15:0]   int_reg_array_57_0_imag;
  reg        [15:0]   int_reg_array_57_1_real;
  reg        [15:0]   int_reg_array_57_1_imag;
  reg        [15:0]   int_reg_array_57_2_real;
  reg        [15:0]   int_reg_array_57_2_imag;
  reg        [15:0]   int_reg_array_57_3_real;
  reg        [15:0]   int_reg_array_57_3_imag;
  reg        [15:0]   int_reg_array_57_4_real;
  reg        [15:0]   int_reg_array_57_4_imag;
  reg        [15:0]   int_reg_array_57_5_real;
  reg        [15:0]   int_reg_array_57_5_imag;
  reg        [15:0]   int_reg_array_57_6_real;
  reg        [15:0]   int_reg_array_57_6_imag;
  reg        [15:0]   int_reg_array_57_7_real;
  reg        [15:0]   int_reg_array_57_7_imag;
  reg        [15:0]   int_reg_array_57_8_real;
  reg        [15:0]   int_reg_array_57_8_imag;
  reg        [15:0]   int_reg_array_57_9_real;
  reg        [15:0]   int_reg_array_57_9_imag;
  reg        [15:0]   int_reg_array_57_10_real;
  reg        [15:0]   int_reg_array_57_10_imag;
  reg        [15:0]   int_reg_array_57_11_real;
  reg        [15:0]   int_reg_array_57_11_imag;
  reg        [15:0]   int_reg_array_57_12_real;
  reg        [15:0]   int_reg_array_57_12_imag;
  reg        [15:0]   int_reg_array_57_13_real;
  reg        [15:0]   int_reg_array_57_13_imag;
  reg        [15:0]   int_reg_array_57_14_real;
  reg        [15:0]   int_reg_array_57_14_imag;
  reg        [15:0]   int_reg_array_57_15_real;
  reg        [15:0]   int_reg_array_57_15_imag;
  reg        [15:0]   int_reg_array_57_16_real;
  reg        [15:0]   int_reg_array_57_16_imag;
  reg        [15:0]   int_reg_array_57_17_real;
  reg        [15:0]   int_reg_array_57_17_imag;
  reg        [15:0]   int_reg_array_57_18_real;
  reg        [15:0]   int_reg_array_57_18_imag;
  reg        [15:0]   int_reg_array_57_19_real;
  reg        [15:0]   int_reg_array_57_19_imag;
  reg        [15:0]   int_reg_array_57_20_real;
  reg        [15:0]   int_reg_array_57_20_imag;
  reg        [15:0]   int_reg_array_57_21_real;
  reg        [15:0]   int_reg_array_57_21_imag;
  reg        [15:0]   int_reg_array_57_22_real;
  reg        [15:0]   int_reg_array_57_22_imag;
  reg        [15:0]   int_reg_array_57_23_real;
  reg        [15:0]   int_reg_array_57_23_imag;
  reg        [15:0]   int_reg_array_57_24_real;
  reg        [15:0]   int_reg_array_57_24_imag;
  reg        [15:0]   int_reg_array_57_25_real;
  reg        [15:0]   int_reg_array_57_25_imag;
  reg        [15:0]   int_reg_array_57_26_real;
  reg        [15:0]   int_reg_array_57_26_imag;
  reg        [15:0]   int_reg_array_57_27_real;
  reg        [15:0]   int_reg_array_57_27_imag;
  reg        [15:0]   int_reg_array_57_28_real;
  reg        [15:0]   int_reg_array_57_28_imag;
  reg        [15:0]   int_reg_array_57_29_real;
  reg        [15:0]   int_reg_array_57_29_imag;
  reg        [15:0]   int_reg_array_57_30_real;
  reg        [15:0]   int_reg_array_57_30_imag;
  reg        [15:0]   int_reg_array_57_31_real;
  reg        [15:0]   int_reg_array_57_31_imag;
  reg        [15:0]   int_reg_array_57_32_real;
  reg        [15:0]   int_reg_array_57_32_imag;
  reg        [15:0]   int_reg_array_57_33_real;
  reg        [15:0]   int_reg_array_57_33_imag;
  reg        [15:0]   int_reg_array_57_34_real;
  reg        [15:0]   int_reg_array_57_34_imag;
  reg        [15:0]   int_reg_array_57_35_real;
  reg        [15:0]   int_reg_array_57_35_imag;
  reg        [15:0]   int_reg_array_57_36_real;
  reg        [15:0]   int_reg_array_57_36_imag;
  reg        [15:0]   int_reg_array_57_37_real;
  reg        [15:0]   int_reg_array_57_37_imag;
  reg        [15:0]   int_reg_array_57_38_real;
  reg        [15:0]   int_reg_array_57_38_imag;
  reg        [15:0]   int_reg_array_57_39_real;
  reg        [15:0]   int_reg_array_57_39_imag;
  reg        [15:0]   int_reg_array_57_40_real;
  reg        [15:0]   int_reg_array_57_40_imag;
  reg        [15:0]   int_reg_array_57_41_real;
  reg        [15:0]   int_reg_array_57_41_imag;
  reg        [15:0]   int_reg_array_57_42_real;
  reg        [15:0]   int_reg_array_57_42_imag;
  reg        [15:0]   int_reg_array_57_43_real;
  reg        [15:0]   int_reg_array_57_43_imag;
  reg        [15:0]   int_reg_array_57_44_real;
  reg        [15:0]   int_reg_array_57_44_imag;
  reg        [15:0]   int_reg_array_57_45_real;
  reg        [15:0]   int_reg_array_57_45_imag;
  reg        [15:0]   int_reg_array_57_46_real;
  reg        [15:0]   int_reg_array_57_46_imag;
  reg        [15:0]   int_reg_array_57_47_real;
  reg        [15:0]   int_reg_array_57_47_imag;
  reg        [15:0]   int_reg_array_57_48_real;
  reg        [15:0]   int_reg_array_57_48_imag;
  reg        [15:0]   int_reg_array_57_49_real;
  reg        [15:0]   int_reg_array_57_49_imag;
  reg        [15:0]   int_reg_array_57_50_real;
  reg        [15:0]   int_reg_array_57_50_imag;
  reg        [15:0]   int_reg_array_57_51_real;
  reg        [15:0]   int_reg_array_57_51_imag;
  reg        [15:0]   int_reg_array_57_52_real;
  reg        [15:0]   int_reg_array_57_52_imag;
  reg        [15:0]   int_reg_array_57_53_real;
  reg        [15:0]   int_reg_array_57_53_imag;
  reg        [15:0]   int_reg_array_57_54_real;
  reg        [15:0]   int_reg_array_57_54_imag;
  reg        [15:0]   int_reg_array_57_55_real;
  reg        [15:0]   int_reg_array_57_55_imag;
  reg        [15:0]   int_reg_array_57_56_real;
  reg        [15:0]   int_reg_array_57_56_imag;
  reg        [15:0]   int_reg_array_57_57_real;
  reg        [15:0]   int_reg_array_57_57_imag;
  reg        [15:0]   int_reg_array_57_58_real;
  reg        [15:0]   int_reg_array_57_58_imag;
  reg        [15:0]   int_reg_array_57_59_real;
  reg        [15:0]   int_reg_array_57_59_imag;
  reg        [15:0]   int_reg_array_57_60_real;
  reg        [15:0]   int_reg_array_57_60_imag;
  reg        [15:0]   int_reg_array_57_61_real;
  reg        [15:0]   int_reg_array_57_61_imag;
  reg        [15:0]   int_reg_array_57_62_real;
  reg        [15:0]   int_reg_array_57_62_imag;
  reg        [15:0]   int_reg_array_57_63_real;
  reg        [15:0]   int_reg_array_57_63_imag;
  reg        [15:0]   int_reg_array_29_0_real;
  reg        [15:0]   int_reg_array_29_0_imag;
  reg        [15:0]   int_reg_array_29_1_real;
  reg        [15:0]   int_reg_array_29_1_imag;
  reg        [15:0]   int_reg_array_29_2_real;
  reg        [15:0]   int_reg_array_29_2_imag;
  reg        [15:0]   int_reg_array_29_3_real;
  reg        [15:0]   int_reg_array_29_3_imag;
  reg        [15:0]   int_reg_array_29_4_real;
  reg        [15:0]   int_reg_array_29_4_imag;
  reg        [15:0]   int_reg_array_29_5_real;
  reg        [15:0]   int_reg_array_29_5_imag;
  reg        [15:0]   int_reg_array_29_6_real;
  reg        [15:0]   int_reg_array_29_6_imag;
  reg        [15:0]   int_reg_array_29_7_real;
  reg        [15:0]   int_reg_array_29_7_imag;
  reg        [15:0]   int_reg_array_29_8_real;
  reg        [15:0]   int_reg_array_29_8_imag;
  reg        [15:0]   int_reg_array_29_9_real;
  reg        [15:0]   int_reg_array_29_9_imag;
  reg        [15:0]   int_reg_array_29_10_real;
  reg        [15:0]   int_reg_array_29_10_imag;
  reg        [15:0]   int_reg_array_29_11_real;
  reg        [15:0]   int_reg_array_29_11_imag;
  reg        [15:0]   int_reg_array_29_12_real;
  reg        [15:0]   int_reg_array_29_12_imag;
  reg        [15:0]   int_reg_array_29_13_real;
  reg        [15:0]   int_reg_array_29_13_imag;
  reg        [15:0]   int_reg_array_29_14_real;
  reg        [15:0]   int_reg_array_29_14_imag;
  reg        [15:0]   int_reg_array_29_15_real;
  reg        [15:0]   int_reg_array_29_15_imag;
  reg        [15:0]   int_reg_array_29_16_real;
  reg        [15:0]   int_reg_array_29_16_imag;
  reg        [15:0]   int_reg_array_29_17_real;
  reg        [15:0]   int_reg_array_29_17_imag;
  reg        [15:0]   int_reg_array_29_18_real;
  reg        [15:0]   int_reg_array_29_18_imag;
  reg        [15:0]   int_reg_array_29_19_real;
  reg        [15:0]   int_reg_array_29_19_imag;
  reg        [15:0]   int_reg_array_29_20_real;
  reg        [15:0]   int_reg_array_29_20_imag;
  reg        [15:0]   int_reg_array_29_21_real;
  reg        [15:0]   int_reg_array_29_21_imag;
  reg        [15:0]   int_reg_array_29_22_real;
  reg        [15:0]   int_reg_array_29_22_imag;
  reg        [15:0]   int_reg_array_29_23_real;
  reg        [15:0]   int_reg_array_29_23_imag;
  reg        [15:0]   int_reg_array_29_24_real;
  reg        [15:0]   int_reg_array_29_24_imag;
  reg        [15:0]   int_reg_array_29_25_real;
  reg        [15:0]   int_reg_array_29_25_imag;
  reg        [15:0]   int_reg_array_29_26_real;
  reg        [15:0]   int_reg_array_29_26_imag;
  reg        [15:0]   int_reg_array_29_27_real;
  reg        [15:0]   int_reg_array_29_27_imag;
  reg        [15:0]   int_reg_array_29_28_real;
  reg        [15:0]   int_reg_array_29_28_imag;
  reg        [15:0]   int_reg_array_29_29_real;
  reg        [15:0]   int_reg_array_29_29_imag;
  reg        [15:0]   int_reg_array_29_30_real;
  reg        [15:0]   int_reg_array_29_30_imag;
  reg        [15:0]   int_reg_array_29_31_real;
  reg        [15:0]   int_reg_array_29_31_imag;
  reg        [15:0]   int_reg_array_29_32_real;
  reg        [15:0]   int_reg_array_29_32_imag;
  reg        [15:0]   int_reg_array_29_33_real;
  reg        [15:0]   int_reg_array_29_33_imag;
  reg        [15:0]   int_reg_array_29_34_real;
  reg        [15:0]   int_reg_array_29_34_imag;
  reg        [15:0]   int_reg_array_29_35_real;
  reg        [15:0]   int_reg_array_29_35_imag;
  reg        [15:0]   int_reg_array_29_36_real;
  reg        [15:0]   int_reg_array_29_36_imag;
  reg        [15:0]   int_reg_array_29_37_real;
  reg        [15:0]   int_reg_array_29_37_imag;
  reg        [15:0]   int_reg_array_29_38_real;
  reg        [15:0]   int_reg_array_29_38_imag;
  reg        [15:0]   int_reg_array_29_39_real;
  reg        [15:0]   int_reg_array_29_39_imag;
  reg        [15:0]   int_reg_array_29_40_real;
  reg        [15:0]   int_reg_array_29_40_imag;
  reg        [15:0]   int_reg_array_29_41_real;
  reg        [15:0]   int_reg_array_29_41_imag;
  reg        [15:0]   int_reg_array_29_42_real;
  reg        [15:0]   int_reg_array_29_42_imag;
  reg        [15:0]   int_reg_array_29_43_real;
  reg        [15:0]   int_reg_array_29_43_imag;
  reg        [15:0]   int_reg_array_29_44_real;
  reg        [15:0]   int_reg_array_29_44_imag;
  reg        [15:0]   int_reg_array_29_45_real;
  reg        [15:0]   int_reg_array_29_45_imag;
  reg        [15:0]   int_reg_array_29_46_real;
  reg        [15:0]   int_reg_array_29_46_imag;
  reg        [15:0]   int_reg_array_29_47_real;
  reg        [15:0]   int_reg_array_29_47_imag;
  reg        [15:0]   int_reg_array_29_48_real;
  reg        [15:0]   int_reg_array_29_48_imag;
  reg        [15:0]   int_reg_array_29_49_real;
  reg        [15:0]   int_reg_array_29_49_imag;
  reg        [15:0]   int_reg_array_29_50_real;
  reg        [15:0]   int_reg_array_29_50_imag;
  reg        [15:0]   int_reg_array_29_51_real;
  reg        [15:0]   int_reg_array_29_51_imag;
  reg        [15:0]   int_reg_array_29_52_real;
  reg        [15:0]   int_reg_array_29_52_imag;
  reg        [15:0]   int_reg_array_29_53_real;
  reg        [15:0]   int_reg_array_29_53_imag;
  reg        [15:0]   int_reg_array_29_54_real;
  reg        [15:0]   int_reg_array_29_54_imag;
  reg        [15:0]   int_reg_array_29_55_real;
  reg        [15:0]   int_reg_array_29_55_imag;
  reg        [15:0]   int_reg_array_29_56_real;
  reg        [15:0]   int_reg_array_29_56_imag;
  reg        [15:0]   int_reg_array_29_57_real;
  reg        [15:0]   int_reg_array_29_57_imag;
  reg        [15:0]   int_reg_array_29_58_real;
  reg        [15:0]   int_reg_array_29_58_imag;
  reg        [15:0]   int_reg_array_29_59_real;
  reg        [15:0]   int_reg_array_29_59_imag;
  reg        [15:0]   int_reg_array_29_60_real;
  reg        [15:0]   int_reg_array_29_60_imag;
  reg        [15:0]   int_reg_array_29_61_real;
  reg        [15:0]   int_reg_array_29_61_imag;
  reg        [15:0]   int_reg_array_29_62_real;
  reg        [15:0]   int_reg_array_29_62_imag;
  reg        [15:0]   int_reg_array_29_63_real;
  reg        [15:0]   int_reg_array_29_63_imag;
  reg        [15:0]   int_reg_array_3_0_real;
  reg        [15:0]   int_reg_array_3_0_imag;
  reg        [15:0]   int_reg_array_3_1_real;
  reg        [15:0]   int_reg_array_3_1_imag;
  reg        [15:0]   int_reg_array_3_2_real;
  reg        [15:0]   int_reg_array_3_2_imag;
  reg        [15:0]   int_reg_array_3_3_real;
  reg        [15:0]   int_reg_array_3_3_imag;
  reg        [15:0]   int_reg_array_3_4_real;
  reg        [15:0]   int_reg_array_3_4_imag;
  reg        [15:0]   int_reg_array_3_5_real;
  reg        [15:0]   int_reg_array_3_5_imag;
  reg        [15:0]   int_reg_array_3_6_real;
  reg        [15:0]   int_reg_array_3_6_imag;
  reg        [15:0]   int_reg_array_3_7_real;
  reg        [15:0]   int_reg_array_3_7_imag;
  reg        [15:0]   int_reg_array_3_8_real;
  reg        [15:0]   int_reg_array_3_8_imag;
  reg        [15:0]   int_reg_array_3_9_real;
  reg        [15:0]   int_reg_array_3_9_imag;
  reg        [15:0]   int_reg_array_3_10_real;
  reg        [15:0]   int_reg_array_3_10_imag;
  reg        [15:0]   int_reg_array_3_11_real;
  reg        [15:0]   int_reg_array_3_11_imag;
  reg        [15:0]   int_reg_array_3_12_real;
  reg        [15:0]   int_reg_array_3_12_imag;
  reg        [15:0]   int_reg_array_3_13_real;
  reg        [15:0]   int_reg_array_3_13_imag;
  reg        [15:0]   int_reg_array_3_14_real;
  reg        [15:0]   int_reg_array_3_14_imag;
  reg        [15:0]   int_reg_array_3_15_real;
  reg        [15:0]   int_reg_array_3_15_imag;
  reg        [15:0]   int_reg_array_3_16_real;
  reg        [15:0]   int_reg_array_3_16_imag;
  reg        [15:0]   int_reg_array_3_17_real;
  reg        [15:0]   int_reg_array_3_17_imag;
  reg        [15:0]   int_reg_array_3_18_real;
  reg        [15:0]   int_reg_array_3_18_imag;
  reg        [15:0]   int_reg_array_3_19_real;
  reg        [15:0]   int_reg_array_3_19_imag;
  reg        [15:0]   int_reg_array_3_20_real;
  reg        [15:0]   int_reg_array_3_20_imag;
  reg        [15:0]   int_reg_array_3_21_real;
  reg        [15:0]   int_reg_array_3_21_imag;
  reg        [15:0]   int_reg_array_3_22_real;
  reg        [15:0]   int_reg_array_3_22_imag;
  reg        [15:0]   int_reg_array_3_23_real;
  reg        [15:0]   int_reg_array_3_23_imag;
  reg        [15:0]   int_reg_array_3_24_real;
  reg        [15:0]   int_reg_array_3_24_imag;
  reg        [15:0]   int_reg_array_3_25_real;
  reg        [15:0]   int_reg_array_3_25_imag;
  reg        [15:0]   int_reg_array_3_26_real;
  reg        [15:0]   int_reg_array_3_26_imag;
  reg        [15:0]   int_reg_array_3_27_real;
  reg        [15:0]   int_reg_array_3_27_imag;
  reg        [15:0]   int_reg_array_3_28_real;
  reg        [15:0]   int_reg_array_3_28_imag;
  reg        [15:0]   int_reg_array_3_29_real;
  reg        [15:0]   int_reg_array_3_29_imag;
  reg        [15:0]   int_reg_array_3_30_real;
  reg        [15:0]   int_reg_array_3_30_imag;
  reg        [15:0]   int_reg_array_3_31_real;
  reg        [15:0]   int_reg_array_3_31_imag;
  reg        [15:0]   int_reg_array_3_32_real;
  reg        [15:0]   int_reg_array_3_32_imag;
  reg        [15:0]   int_reg_array_3_33_real;
  reg        [15:0]   int_reg_array_3_33_imag;
  reg        [15:0]   int_reg_array_3_34_real;
  reg        [15:0]   int_reg_array_3_34_imag;
  reg        [15:0]   int_reg_array_3_35_real;
  reg        [15:0]   int_reg_array_3_35_imag;
  reg        [15:0]   int_reg_array_3_36_real;
  reg        [15:0]   int_reg_array_3_36_imag;
  reg        [15:0]   int_reg_array_3_37_real;
  reg        [15:0]   int_reg_array_3_37_imag;
  reg        [15:0]   int_reg_array_3_38_real;
  reg        [15:0]   int_reg_array_3_38_imag;
  reg        [15:0]   int_reg_array_3_39_real;
  reg        [15:0]   int_reg_array_3_39_imag;
  reg        [15:0]   int_reg_array_3_40_real;
  reg        [15:0]   int_reg_array_3_40_imag;
  reg        [15:0]   int_reg_array_3_41_real;
  reg        [15:0]   int_reg_array_3_41_imag;
  reg        [15:0]   int_reg_array_3_42_real;
  reg        [15:0]   int_reg_array_3_42_imag;
  reg        [15:0]   int_reg_array_3_43_real;
  reg        [15:0]   int_reg_array_3_43_imag;
  reg        [15:0]   int_reg_array_3_44_real;
  reg        [15:0]   int_reg_array_3_44_imag;
  reg        [15:0]   int_reg_array_3_45_real;
  reg        [15:0]   int_reg_array_3_45_imag;
  reg        [15:0]   int_reg_array_3_46_real;
  reg        [15:0]   int_reg_array_3_46_imag;
  reg        [15:0]   int_reg_array_3_47_real;
  reg        [15:0]   int_reg_array_3_47_imag;
  reg        [15:0]   int_reg_array_3_48_real;
  reg        [15:0]   int_reg_array_3_48_imag;
  reg        [15:0]   int_reg_array_3_49_real;
  reg        [15:0]   int_reg_array_3_49_imag;
  reg        [15:0]   int_reg_array_3_50_real;
  reg        [15:0]   int_reg_array_3_50_imag;
  reg        [15:0]   int_reg_array_3_51_real;
  reg        [15:0]   int_reg_array_3_51_imag;
  reg        [15:0]   int_reg_array_3_52_real;
  reg        [15:0]   int_reg_array_3_52_imag;
  reg        [15:0]   int_reg_array_3_53_real;
  reg        [15:0]   int_reg_array_3_53_imag;
  reg        [15:0]   int_reg_array_3_54_real;
  reg        [15:0]   int_reg_array_3_54_imag;
  reg        [15:0]   int_reg_array_3_55_real;
  reg        [15:0]   int_reg_array_3_55_imag;
  reg        [15:0]   int_reg_array_3_56_real;
  reg        [15:0]   int_reg_array_3_56_imag;
  reg        [15:0]   int_reg_array_3_57_real;
  reg        [15:0]   int_reg_array_3_57_imag;
  reg        [15:0]   int_reg_array_3_58_real;
  reg        [15:0]   int_reg_array_3_58_imag;
  reg        [15:0]   int_reg_array_3_59_real;
  reg        [15:0]   int_reg_array_3_59_imag;
  reg        [15:0]   int_reg_array_3_60_real;
  reg        [15:0]   int_reg_array_3_60_imag;
  reg        [15:0]   int_reg_array_3_61_real;
  reg        [15:0]   int_reg_array_3_61_imag;
  reg        [15:0]   int_reg_array_3_62_real;
  reg        [15:0]   int_reg_array_3_62_imag;
  reg        [15:0]   int_reg_array_3_63_real;
  reg        [15:0]   int_reg_array_3_63_imag;
  reg        [15:0]   int_reg_array_36_0_real;
  reg        [15:0]   int_reg_array_36_0_imag;
  reg        [15:0]   int_reg_array_36_1_real;
  reg        [15:0]   int_reg_array_36_1_imag;
  reg        [15:0]   int_reg_array_36_2_real;
  reg        [15:0]   int_reg_array_36_2_imag;
  reg        [15:0]   int_reg_array_36_3_real;
  reg        [15:0]   int_reg_array_36_3_imag;
  reg        [15:0]   int_reg_array_36_4_real;
  reg        [15:0]   int_reg_array_36_4_imag;
  reg        [15:0]   int_reg_array_36_5_real;
  reg        [15:0]   int_reg_array_36_5_imag;
  reg        [15:0]   int_reg_array_36_6_real;
  reg        [15:0]   int_reg_array_36_6_imag;
  reg        [15:0]   int_reg_array_36_7_real;
  reg        [15:0]   int_reg_array_36_7_imag;
  reg        [15:0]   int_reg_array_36_8_real;
  reg        [15:0]   int_reg_array_36_8_imag;
  reg        [15:0]   int_reg_array_36_9_real;
  reg        [15:0]   int_reg_array_36_9_imag;
  reg        [15:0]   int_reg_array_36_10_real;
  reg        [15:0]   int_reg_array_36_10_imag;
  reg        [15:0]   int_reg_array_36_11_real;
  reg        [15:0]   int_reg_array_36_11_imag;
  reg        [15:0]   int_reg_array_36_12_real;
  reg        [15:0]   int_reg_array_36_12_imag;
  reg        [15:0]   int_reg_array_36_13_real;
  reg        [15:0]   int_reg_array_36_13_imag;
  reg        [15:0]   int_reg_array_36_14_real;
  reg        [15:0]   int_reg_array_36_14_imag;
  reg        [15:0]   int_reg_array_36_15_real;
  reg        [15:0]   int_reg_array_36_15_imag;
  reg        [15:0]   int_reg_array_36_16_real;
  reg        [15:0]   int_reg_array_36_16_imag;
  reg        [15:0]   int_reg_array_36_17_real;
  reg        [15:0]   int_reg_array_36_17_imag;
  reg        [15:0]   int_reg_array_36_18_real;
  reg        [15:0]   int_reg_array_36_18_imag;
  reg        [15:0]   int_reg_array_36_19_real;
  reg        [15:0]   int_reg_array_36_19_imag;
  reg        [15:0]   int_reg_array_36_20_real;
  reg        [15:0]   int_reg_array_36_20_imag;
  reg        [15:0]   int_reg_array_36_21_real;
  reg        [15:0]   int_reg_array_36_21_imag;
  reg        [15:0]   int_reg_array_36_22_real;
  reg        [15:0]   int_reg_array_36_22_imag;
  reg        [15:0]   int_reg_array_36_23_real;
  reg        [15:0]   int_reg_array_36_23_imag;
  reg        [15:0]   int_reg_array_36_24_real;
  reg        [15:0]   int_reg_array_36_24_imag;
  reg        [15:0]   int_reg_array_36_25_real;
  reg        [15:0]   int_reg_array_36_25_imag;
  reg        [15:0]   int_reg_array_36_26_real;
  reg        [15:0]   int_reg_array_36_26_imag;
  reg        [15:0]   int_reg_array_36_27_real;
  reg        [15:0]   int_reg_array_36_27_imag;
  reg        [15:0]   int_reg_array_36_28_real;
  reg        [15:0]   int_reg_array_36_28_imag;
  reg        [15:0]   int_reg_array_36_29_real;
  reg        [15:0]   int_reg_array_36_29_imag;
  reg        [15:0]   int_reg_array_36_30_real;
  reg        [15:0]   int_reg_array_36_30_imag;
  reg        [15:0]   int_reg_array_36_31_real;
  reg        [15:0]   int_reg_array_36_31_imag;
  reg        [15:0]   int_reg_array_36_32_real;
  reg        [15:0]   int_reg_array_36_32_imag;
  reg        [15:0]   int_reg_array_36_33_real;
  reg        [15:0]   int_reg_array_36_33_imag;
  reg        [15:0]   int_reg_array_36_34_real;
  reg        [15:0]   int_reg_array_36_34_imag;
  reg        [15:0]   int_reg_array_36_35_real;
  reg        [15:0]   int_reg_array_36_35_imag;
  reg        [15:0]   int_reg_array_36_36_real;
  reg        [15:0]   int_reg_array_36_36_imag;
  reg        [15:0]   int_reg_array_36_37_real;
  reg        [15:0]   int_reg_array_36_37_imag;
  reg        [15:0]   int_reg_array_36_38_real;
  reg        [15:0]   int_reg_array_36_38_imag;
  reg        [15:0]   int_reg_array_36_39_real;
  reg        [15:0]   int_reg_array_36_39_imag;
  reg        [15:0]   int_reg_array_36_40_real;
  reg        [15:0]   int_reg_array_36_40_imag;
  reg        [15:0]   int_reg_array_36_41_real;
  reg        [15:0]   int_reg_array_36_41_imag;
  reg        [15:0]   int_reg_array_36_42_real;
  reg        [15:0]   int_reg_array_36_42_imag;
  reg        [15:0]   int_reg_array_36_43_real;
  reg        [15:0]   int_reg_array_36_43_imag;
  reg        [15:0]   int_reg_array_36_44_real;
  reg        [15:0]   int_reg_array_36_44_imag;
  reg        [15:0]   int_reg_array_36_45_real;
  reg        [15:0]   int_reg_array_36_45_imag;
  reg        [15:0]   int_reg_array_36_46_real;
  reg        [15:0]   int_reg_array_36_46_imag;
  reg        [15:0]   int_reg_array_36_47_real;
  reg        [15:0]   int_reg_array_36_47_imag;
  reg        [15:0]   int_reg_array_36_48_real;
  reg        [15:0]   int_reg_array_36_48_imag;
  reg        [15:0]   int_reg_array_36_49_real;
  reg        [15:0]   int_reg_array_36_49_imag;
  reg        [15:0]   int_reg_array_36_50_real;
  reg        [15:0]   int_reg_array_36_50_imag;
  reg        [15:0]   int_reg_array_36_51_real;
  reg        [15:0]   int_reg_array_36_51_imag;
  reg        [15:0]   int_reg_array_36_52_real;
  reg        [15:0]   int_reg_array_36_52_imag;
  reg        [15:0]   int_reg_array_36_53_real;
  reg        [15:0]   int_reg_array_36_53_imag;
  reg        [15:0]   int_reg_array_36_54_real;
  reg        [15:0]   int_reg_array_36_54_imag;
  reg        [15:0]   int_reg_array_36_55_real;
  reg        [15:0]   int_reg_array_36_55_imag;
  reg        [15:0]   int_reg_array_36_56_real;
  reg        [15:0]   int_reg_array_36_56_imag;
  reg        [15:0]   int_reg_array_36_57_real;
  reg        [15:0]   int_reg_array_36_57_imag;
  reg        [15:0]   int_reg_array_36_58_real;
  reg        [15:0]   int_reg_array_36_58_imag;
  reg        [15:0]   int_reg_array_36_59_real;
  reg        [15:0]   int_reg_array_36_59_imag;
  reg        [15:0]   int_reg_array_36_60_real;
  reg        [15:0]   int_reg_array_36_60_imag;
  reg        [15:0]   int_reg_array_36_61_real;
  reg        [15:0]   int_reg_array_36_61_imag;
  reg        [15:0]   int_reg_array_36_62_real;
  reg        [15:0]   int_reg_array_36_62_imag;
  reg        [15:0]   int_reg_array_36_63_real;
  reg        [15:0]   int_reg_array_36_63_imag;
  reg        [15:0]   int_reg_array_7_0_real;
  reg        [15:0]   int_reg_array_7_0_imag;
  reg        [15:0]   int_reg_array_7_1_real;
  reg        [15:0]   int_reg_array_7_1_imag;
  reg        [15:0]   int_reg_array_7_2_real;
  reg        [15:0]   int_reg_array_7_2_imag;
  reg        [15:0]   int_reg_array_7_3_real;
  reg        [15:0]   int_reg_array_7_3_imag;
  reg        [15:0]   int_reg_array_7_4_real;
  reg        [15:0]   int_reg_array_7_4_imag;
  reg        [15:0]   int_reg_array_7_5_real;
  reg        [15:0]   int_reg_array_7_5_imag;
  reg        [15:0]   int_reg_array_7_6_real;
  reg        [15:0]   int_reg_array_7_6_imag;
  reg        [15:0]   int_reg_array_7_7_real;
  reg        [15:0]   int_reg_array_7_7_imag;
  reg        [15:0]   int_reg_array_7_8_real;
  reg        [15:0]   int_reg_array_7_8_imag;
  reg        [15:0]   int_reg_array_7_9_real;
  reg        [15:0]   int_reg_array_7_9_imag;
  reg        [15:0]   int_reg_array_7_10_real;
  reg        [15:0]   int_reg_array_7_10_imag;
  reg        [15:0]   int_reg_array_7_11_real;
  reg        [15:0]   int_reg_array_7_11_imag;
  reg        [15:0]   int_reg_array_7_12_real;
  reg        [15:0]   int_reg_array_7_12_imag;
  reg        [15:0]   int_reg_array_7_13_real;
  reg        [15:0]   int_reg_array_7_13_imag;
  reg        [15:0]   int_reg_array_7_14_real;
  reg        [15:0]   int_reg_array_7_14_imag;
  reg        [15:0]   int_reg_array_7_15_real;
  reg        [15:0]   int_reg_array_7_15_imag;
  reg        [15:0]   int_reg_array_7_16_real;
  reg        [15:0]   int_reg_array_7_16_imag;
  reg        [15:0]   int_reg_array_7_17_real;
  reg        [15:0]   int_reg_array_7_17_imag;
  reg        [15:0]   int_reg_array_7_18_real;
  reg        [15:0]   int_reg_array_7_18_imag;
  reg        [15:0]   int_reg_array_7_19_real;
  reg        [15:0]   int_reg_array_7_19_imag;
  reg        [15:0]   int_reg_array_7_20_real;
  reg        [15:0]   int_reg_array_7_20_imag;
  reg        [15:0]   int_reg_array_7_21_real;
  reg        [15:0]   int_reg_array_7_21_imag;
  reg        [15:0]   int_reg_array_7_22_real;
  reg        [15:0]   int_reg_array_7_22_imag;
  reg        [15:0]   int_reg_array_7_23_real;
  reg        [15:0]   int_reg_array_7_23_imag;
  reg        [15:0]   int_reg_array_7_24_real;
  reg        [15:0]   int_reg_array_7_24_imag;
  reg        [15:0]   int_reg_array_7_25_real;
  reg        [15:0]   int_reg_array_7_25_imag;
  reg        [15:0]   int_reg_array_7_26_real;
  reg        [15:0]   int_reg_array_7_26_imag;
  reg        [15:0]   int_reg_array_7_27_real;
  reg        [15:0]   int_reg_array_7_27_imag;
  reg        [15:0]   int_reg_array_7_28_real;
  reg        [15:0]   int_reg_array_7_28_imag;
  reg        [15:0]   int_reg_array_7_29_real;
  reg        [15:0]   int_reg_array_7_29_imag;
  reg        [15:0]   int_reg_array_7_30_real;
  reg        [15:0]   int_reg_array_7_30_imag;
  reg        [15:0]   int_reg_array_7_31_real;
  reg        [15:0]   int_reg_array_7_31_imag;
  reg        [15:0]   int_reg_array_7_32_real;
  reg        [15:0]   int_reg_array_7_32_imag;
  reg        [15:0]   int_reg_array_7_33_real;
  reg        [15:0]   int_reg_array_7_33_imag;
  reg        [15:0]   int_reg_array_7_34_real;
  reg        [15:0]   int_reg_array_7_34_imag;
  reg        [15:0]   int_reg_array_7_35_real;
  reg        [15:0]   int_reg_array_7_35_imag;
  reg        [15:0]   int_reg_array_7_36_real;
  reg        [15:0]   int_reg_array_7_36_imag;
  reg        [15:0]   int_reg_array_7_37_real;
  reg        [15:0]   int_reg_array_7_37_imag;
  reg        [15:0]   int_reg_array_7_38_real;
  reg        [15:0]   int_reg_array_7_38_imag;
  reg        [15:0]   int_reg_array_7_39_real;
  reg        [15:0]   int_reg_array_7_39_imag;
  reg        [15:0]   int_reg_array_7_40_real;
  reg        [15:0]   int_reg_array_7_40_imag;
  reg        [15:0]   int_reg_array_7_41_real;
  reg        [15:0]   int_reg_array_7_41_imag;
  reg        [15:0]   int_reg_array_7_42_real;
  reg        [15:0]   int_reg_array_7_42_imag;
  reg        [15:0]   int_reg_array_7_43_real;
  reg        [15:0]   int_reg_array_7_43_imag;
  reg        [15:0]   int_reg_array_7_44_real;
  reg        [15:0]   int_reg_array_7_44_imag;
  reg        [15:0]   int_reg_array_7_45_real;
  reg        [15:0]   int_reg_array_7_45_imag;
  reg        [15:0]   int_reg_array_7_46_real;
  reg        [15:0]   int_reg_array_7_46_imag;
  reg        [15:0]   int_reg_array_7_47_real;
  reg        [15:0]   int_reg_array_7_47_imag;
  reg        [15:0]   int_reg_array_7_48_real;
  reg        [15:0]   int_reg_array_7_48_imag;
  reg        [15:0]   int_reg_array_7_49_real;
  reg        [15:0]   int_reg_array_7_49_imag;
  reg        [15:0]   int_reg_array_7_50_real;
  reg        [15:0]   int_reg_array_7_50_imag;
  reg        [15:0]   int_reg_array_7_51_real;
  reg        [15:0]   int_reg_array_7_51_imag;
  reg        [15:0]   int_reg_array_7_52_real;
  reg        [15:0]   int_reg_array_7_52_imag;
  reg        [15:0]   int_reg_array_7_53_real;
  reg        [15:0]   int_reg_array_7_53_imag;
  reg        [15:0]   int_reg_array_7_54_real;
  reg        [15:0]   int_reg_array_7_54_imag;
  reg        [15:0]   int_reg_array_7_55_real;
  reg        [15:0]   int_reg_array_7_55_imag;
  reg        [15:0]   int_reg_array_7_56_real;
  reg        [15:0]   int_reg_array_7_56_imag;
  reg        [15:0]   int_reg_array_7_57_real;
  reg        [15:0]   int_reg_array_7_57_imag;
  reg        [15:0]   int_reg_array_7_58_real;
  reg        [15:0]   int_reg_array_7_58_imag;
  reg        [15:0]   int_reg_array_7_59_real;
  reg        [15:0]   int_reg_array_7_59_imag;
  reg        [15:0]   int_reg_array_7_60_real;
  reg        [15:0]   int_reg_array_7_60_imag;
  reg        [15:0]   int_reg_array_7_61_real;
  reg        [15:0]   int_reg_array_7_61_imag;
  reg        [15:0]   int_reg_array_7_62_real;
  reg        [15:0]   int_reg_array_7_62_imag;
  reg        [15:0]   int_reg_array_7_63_real;
  reg        [15:0]   int_reg_array_7_63_imag;
  reg        [15:0]   int_reg_array_54_0_real;
  reg        [15:0]   int_reg_array_54_0_imag;
  reg        [15:0]   int_reg_array_54_1_real;
  reg        [15:0]   int_reg_array_54_1_imag;
  reg        [15:0]   int_reg_array_54_2_real;
  reg        [15:0]   int_reg_array_54_2_imag;
  reg        [15:0]   int_reg_array_54_3_real;
  reg        [15:0]   int_reg_array_54_3_imag;
  reg        [15:0]   int_reg_array_54_4_real;
  reg        [15:0]   int_reg_array_54_4_imag;
  reg        [15:0]   int_reg_array_54_5_real;
  reg        [15:0]   int_reg_array_54_5_imag;
  reg        [15:0]   int_reg_array_54_6_real;
  reg        [15:0]   int_reg_array_54_6_imag;
  reg        [15:0]   int_reg_array_54_7_real;
  reg        [15:0]   int_reg_array_54_7_imag;
  reg        [15:0]   int_reg_array_54_8_real;
  reg        [15:0]   int_reg_array_54_8_imag;
  reg        [15:0]   int_reg_array_54_9_real;
  reg        [15:0]   int_reg_array_54_9_imag;
  reg        [15:0]   int_reg_array_54_10_real;
  reg        [15:0]   int_reg_array_54_10_imag;
  reg        [15:0]   int_reg_array_54_11_real;
  reg        [15:0]   int_reg_array_54_11_imag;
  reg        [15:0]   int_reg_array_54_12_real;
  reg        [15:0]   int_reg_array_54_12_imag;
  reg        [15:0]   int_reg_array_54_13_real;
  reg        [15:0]   int_reg_array_54_13_imag;
  reg        [15:0]   int_reg_array_54_14_real;
  reg        [15:0]   int_reg_array_54_14_imag;
  reg        [15:0]   int_reg_array_54_15_real;
  reg        [15:0]   int_reg_array_54_15_imag;
  reg        [15:0]   int_reg_array_54_16_real;
  reg        [15:0]   int_reg_array_54_16_imag;
  reg        [15:0]   int_reg_array_54_17_real;
  reg        [15:0]   int_reg_array_54_17_imag;
  reg        [15:0]   int_reg_array_54_18_real;
  reg        [15:0]   int_reg_array_54_18_imag;
  reg        [15:0]   int_reg_array_54_19_real;
  reg        [15:0]   int_reg_array_54_19_imag;
  reg        [15:0]   int_reg_array_54_20_real;
  reg        [15:0]   int_reg_array_54_20_imag;
  reg        [15:0]   int_reg_array_54_21_real;
  reg        [15:0]   int_reg_array_54_21_imag;
  reg        [15:0]   int_reg_array_54_22_real;
  reg        [15:0]   int_reg_array_54_22_imag;
  reg        [15:0]   int_reg_array_54_23_real;
  reg        [15:0]   int_reg_array_54_23_imag;
  reg        [15:0]   int_reg_array_54_24_real;
  reg        [15:0]   int_reg_array_54_24_imag;
  reg        [15:0]   int_reg_array_54_25_real;
  reg        [15:0]   int_reg_array_54_25_imag;
  reg        [15:0]   int_reg_array_54_26_real;
  reg        [15:0]   int_reg_array_54_26_imag;
  reg        [15:0]   int_reg_array_54_27_real;
  reg        [15:0]   int_reg_array_54_27_imag;
  reg        [15:0]   int_reg_array_54_28_real;
  reg        [15:0]   int_reg_array_54_28_imag;
  reg        [15:0]   int_reg_array_54_29_real;
  reg        [15:0]   int_reg_array_54_29_imag;
  reg        [15:0]   int_reg_array_54_30_real;
  reg        [15:0]   int_reg_array_54_30_imag;
  reg        [15:0]   int_reg_array_54_31_real;
  reg        [15:0]   int_reg_array_54_31_imag;
  reg        [15:0]   int_reg_array_54_32_real;
  reg        [15:0]   int_reg_array_54_32_imag;
  reg        [15:0]   int_reg_array_54_33_real;
  reg        [15:0]   int_reg_array_54_33_imag;
  reg        [15:0]   int_reg_array_54_34_real;
  reg        [15:0]   int_reg_array_54_34_imag;
  reg        [15:0]   int_reg_array_54_35_real;
  reg        [15:0]   int_reg_array_54_35_imag;
  reg        [15:0]   int_reg_array_54_36_real;
  reg        [15:0]   int_reg_array_54_36_imag;
  reg        [15:0]   int_reg_array_54_37_real;
  reg        [15:0]   int_reg_array_54_37_imag;
  reg        [15:0]   int_reg_array_54_38_real;
  reg        [15:0]   int_reg_array_54_38_imag;
  reg        [15:0]   int_reg_array_54_39_real;
  reg        [15:0]   int_reg_array_54_39_imag;
  reg        [15:0]   int_reg_array_54_40_real;
  reg        [15:0]   int_reg_array_54_40_imag;
  reg        [15:0]   int_reg_array_54_41_real;
  reg        [15:0]   int_reg_array_54_41_imag;
  reg        [15:0]   int_reg_array_54_42_real;
  reg        [15:0]   int_reg_array_54_42_imag;
  reg        [15:0]   int_reg_array_54_43_real;
  reg        [15:0]   int_reg_array_54_43_imag;
  reg        [15:0]   int_reg_array_54_44_real;
  reg        [15:0]   int_reg_array_54_44_imag;
  reg        [15:0]   int_reg_array_54_45_real;
  reg        [15:0]   int_reg_array_54_45_imag;
  reg        [15:0]   int_reg_array_54_46_real;
  reg        [15:0]   int_reg_array_54_46_imag;
  reg        [15:0]   int_reg_array_54_47_real;
  reg        [15:0]   int_reg_array_54_47_imag;
  reg        [15:0]   int_reg_array_54_48_real;
  reg        [15:0]   int_reg_array_54_48_imag;
  reg        [15:0]   int_reg_array_54_49_real;
  reg        [15:0]   int_reg_array_54_49_imag;
  reg        [15:0]   int_reg_array_54_50_real;
  reg        [15:0]   int_reg_array_54_50_imag;
  reg        [15:0]   int_reg_array_54_51_real;
  reg        [15:0]   int_reg_array_54_51_imag;
  reg        [15:0]   int_reg_array_54_52_real;
  reg        [15:0]   int_reg_array_54_52_imag;
  reg        [15:0]   int_reg_array_54_53_real;
  reg        [15:0]   int_reg_array_54_53_imag;
  reg        [15:0]   int_reg_array_54_54_real;
  reg        [15:0]   int_reg_array_54_54_imag;
  reg        [15:0]   int_reg_array_54_55_real;
  reg        [15:0]   int_reg_array_54_55_imag;
  reg        [15:0]   int_reg_array_54_56_real;
  reg        [15:0]   int_reg_array_54_56_imag;
  reg        [15:0]   int_reg_array_54_57_real;
  reg        [15:0]   int_reg_array_54_57_imag;
  reg        [15:0]   int_reg_array_54_58_real;
  reg        [15:0]   int_reg_array_54_58_imag;
  reg        [15:0]   int_reg_array_54_59_real;
  reg        [15:0]   int_reg_array_54_59_imag;
  reg        [15:0]   int_reg_array_54_60_real;
  reg        [15:0]   int_reg_array_54_60_imag;
  reg        [15:0]   int_reg_array_54_61_real;
  reg        [15:0]   int_reg_array_54_61_imag;
  reg        [15:0]   int_reg_array_54_62_real;
  reg        [15:0]   int_reg_array_54_62_imag;
  reg        [15:0]   int_reg_array_54_63_real;
  reg        [15:0]   int_reg_array_54_63_imag;
  reg        [15:0]   int_reg_array_23_0_real;
  reg        [15:0]   int_reg_array_23_0_imag;
  reg        [15:0]   int_reg_array_23_1_real;
  reg        [15:0]   int_reg_array_23_1_imag;
  reg        [15:0]   int_reg_array_23_2_real;
  reg        [15:0]   int_reg_array_23_2_imag;
  reg        [15:0]   int_reg_array_23_3_real;
  reg        [15:0]   int_reg_array_23_3_imag;
  reg        [15:0]   int_reg_array_23_4_real;
  reg        [15:0]   int_reg_array_23_4_imag;
  reg        [15:0]   int_reg_array_23_5_real;
  reg        [15:0]   int_reg_array_23_5_imag;
  reg        [15:0]   int_reg_array_23_6_real;
  reg        [15:0]   int_reg_array_23_6_imag;
  reg        [15:0]   int_reg_array_23_7_real;
  reg        [15:0]   int_reg_array_23_7_imag;
  reg        [15:0]   int_reg_array_23_8_real;
  reg        [15:0]   int_reg_array_23_8_imag;
  reg        [15:0]   int_reg_array_23_9_real;
  reg        [15:0]   int_reg_array_23_9_imag;
  reg        [15:0]   int_reg_array_23_10_real;
  reg        [15:0]   int_reg_array_23_10_imag;
  reg        [15:0]   int_reg_array_23_11_real;
  reg        [15:0]   int_reg_array_23_11_imag;
  reg        [15:0]   int_reg_array_23_12_real;
  reg        [15:0]   int_reg_array_23_12_imag;
  reg        [15:0]   int_reg_array_23_13_real;
  reg        [15:0]   int_reg_array_23_13_imag;
  reg        [15:0]   int_reg_array_23_14_real;
  reg        [15:0]   int_reg_array_23_14_imag;
  reg        [15:0]   int_reg_array_23_15_real;
  reg        [15:0]   int_reg_array_23_15_imag;
  reg        [15:0]   int_reg_array_23_16_real;
  reg        [15:0]   int_reg_array_23_16_imag;
  reg        [15:0]   int_reg_array_23_17_real;
  reg        [15:0]   int_reg_array_23_17_imag;
  reg        [15:0]   int_reg_array_23_18_real;
  reg        [15:0]   int_reg_array_23_18_imag;
  reg        [15:0]   int_reg_array_23_19_real;
  reg        [15:0]   int_reg_array_23_19_imag;
  reg        [15:0]   int_reg_array_23_20_real;
  reg        [15:0]   int_reg_array_23_20_imag;
  reg        [15:0]   int_reg_array_23_21_real;
  reg        [15:0]   int_reg_array_23_21_imag;
  reg        [15:0]   int_reg_array_23_22_real;
  reg        [15:0]   int_reg_array_23_22_imag;
  reg        [15:0]   int_reg_array_23_23_real;
  reg        [15:0]   int_reg_array_23_23_imag;
  reg        [15:0]   int_reg_array_23_24_real;
  reg        [15:0]   int_reg_array_23_24_imag;
  reg        [15:0]   int_reg_array_23_25_real;
  reg        [15:0]   int_reg_array_23_25_imag;
  reg        [15:0]   int_reg_array_23_26_real;
  reg        [15:0]   int_reg_array_23_26_imag;
  reg        [15:0]   int_reg_array_23_27_real;
  reg        [15:0]   int_reg_array_23_27_imag;
  reg        [15:0]   int_reg_array_23_28_real;
  reg        [15:0]   int_reg_array_23_28_imag;
  reg        [15:0]   int_reg_array_23_29_real;
  reg        [15:0]   int_reg_array_23_29_imag;
  reg        [15:0]   int_reg_array_23_30_real;
  reg        [15:0]   int_reg_array_23_30_imag;
  reg        [15:0]   int_reg_array_23_31_real;
  reg        [15:0]   int_reg_array_23_31_imag;
  reg        [15:0]   int_reg_array_23_32_real;
  reg        [15:0]   int_reg_array_23_32_imag;
  reg        [15:0]   int_reg_array_23_33_real;
  reg        [15:0]   int_reg_array_23_33_imag;
  reg        [15:0]   int_reg_array_23_34_real;
  reg        [15:0]   int_reg_array_23_34_imag;
  reg        [15:0]   int_reg_array_23_35_real;
  reg        [15:0]   int_reg_array_23_35_imag;
  reg        [15:0]   int_reg_array_23_36_real;
  reg        [15:0]   int_reg_array_23_36_imag;
  reg        [15:0]   int_reg_array_23_37_real;
  reg        [15:0]   int_reg_array_23_37_imag;
  reg        [15:0]   int_reg_array_23_38_real;
  reg        [15:0]   int_reg_array_23_38_imag;
  reg        [15:0]   int_reg_array_23_39_real;
  reg        [15:0]   int_reg_array_23_39_imag;
  reg        [15:0]   int_reg_array_23_40_real;
  reg        [15:0]   int_reg_array_23_40_imag;
  reg        [15:0]   int_reg_array_23_41_real;
  reg        [15:0]   int_reg_array_23_41_imag;
  reg        [15:0]   int_reg_array_23_42_real;
  reg        [15:0]   int_reg_array_23_42_imag;
  reg        [15:0]   int_reg_array_23_43_real;
  reg        [15:0]   int_reg_array_23_43_imag;
  reg        [15:0]   int_reg_array_23_44_real;
  reg        [15:0]   int_reg_array_23_44_imag;
  reg        [15:0]   int_reg_array_23_45_real;
  reg        [15:0]   int_reg_array_23_45_imag;
  reg        [15:0]   int_reg_array_23_46_real;
  reg        [15:0]   int_reg_array_23_46_imag;
  reg        [15:0]   int_reg_array_23_47_real;
  reg        [15:0]   int_reg_array_23_47_imag;
  reg        [15:0]   int_reg_array_23_48_real;
  reg        [15:0]   int_reg_array_23_48_imag;
  reg        [15:0]   int_reg_array_23_49_real;
  reg        [15:0]   int_reg_array_23_49_imag;
  reg        [15:0]   int_reg_array_23_50_real;
  reg        [15:0]   int_reg_array_23_50_imag;
  reg        [15:0]   int_reg_array_23_51_real;
  reg        [15:0]   int_reg_array_23_51_imag;
  reg        [15:0]   int_reg_array_23_52_real;
  reg        [15:0]   int_reg_array_23_52_imag;
  reg        [15:0]   int_reg_array_23_53_real;
  reg        [15:0]   int_reg_array_23_53_imag;
  reg        [15:0]   int_reg_array_23_54_real;
  reg        [15:0]   int_reg_array_23_54_imag;
  reg        [15:0]   int_reg_array_23_55_real;
  reg        [15:0]   int_reg_array_23_55_imag;
  reg        [15:0]   int_reg_array_23_56_real;
  reg        [15:0]   int_reg_array_23_56_imag;
  reg        [15:0]   int_reg_array_23_57_real;
  reg        [15:0]   int_reg_array_23_57_imag;
  reg        [15:0]   int_reg_array_23_58_real;
  reg        [15:0]   int_reg_array_23_58_imag;
  reg        [15:0]   int_reg_array_23_59_real;
  reg        [15:0]   int_reg_array_23_59_imag;
  reg        [15:0]   int_reg_array_23_60_real;
  reg        [15:0]   int_reg_array_23_60_imag;
  reg        [15:0]   int_reg_array_23_61_real;
  reg        [15:0]   int_reg_array_23_61_imag;
  reg        [15:0]   int_reg_array_23_62_real;
  reg        [15:0]   int_reg_array_23_62_imag;
  reg        [15:0]   int_reg_array_23_63_real;
  reg        [15:0]   int_reg_array_23_63_imag;
  reg        [15:0]   int_reg_array_4_0_real;
  reg        [15:0]   int_reg_array_4_0_imag;
  reg        [15:0]   int_reg_array_4_1_real;
  reg        [15:0]   int_reg_array_4_1_imag;
  reg        [15:0]   int_reg_array_4_2_real;
  reg        [15:0]   int_reg_array_4_2_imag;
  reg        [15:0]   int_reg_array_4_3_real;
  reg        [15:0]   int_reg_array_4_3_imag;
  reg        [15:0]   int_reg_array_4_4_real;
  reg        [15:0]   int_reg_array_4_4_imag;
  reg        [15:0]   int_reg_array_4_5_real;
  reg        [15:0]   int_reg_array_4_5_imag;
  reg        [15:0]   int_reg_array_4_6_real;
  reg        [15:0]   int_reg_array_4_6_imag;
  reg        [15:0]   int_reg_array_4_7_real;
  reg        [15:0]   int_reg_array_4_7_imag;
  reg        [15:0]   int_reg_array_4_8_real;
  reg        [15:0]   int_reg_array_4_8_imag;
  reg        [15:0]   int_reg_array_4_9_real;
  reg        [15:0]   int_reg_array_4_9_imag;
  reg        [15:0]   int_reg_array_4_10_real;
  reg        [15:0]   int_reg_array_4_10_imag;
  reg        [15:0]   int_reg_array_4_11_real;
  reg        [15:0]   int_reg_array_4_11_imag;
  reg        [15:0]   int_reg_array_4_12_real;
  reg        [15:0]   int_reg_array_4_12_imag;
  reg        [15:0]   int_reg_array_4_13_real;
  reg        [15:0]   int_reg_array_4_13_imag;
  reg        [15:0]   int_reg_array_4_14_real;
  reg        [15:0]   int_reg_array_4_14_imag;
  reg        [15:0]   int_reg_array_4_15_real;
  reg        [15:0]   int_reg_array_4_15_imag;
  reg        [15:0]   int_reg_array_4_16_real;
  reg        [15:0]   int_reg_array_4_16_imag;
  reg        [15:0]   int_reg_array_4_17_real;
  reg        [15:0]   int_reg_array_4_17_imag;
  reg        [15:0]   int_reg_array_4_18_real;
  reg        [15:0]   int_reg_array_4_18_imag;
  reg        [15:0]   int_reg_array_4_19_real;
  reg        [15:0]   int_reg_array_4_19_imag;
  reg        [15:0]   int_reg_array_4_20_real;
  reg        [15:0]   int_reg_array_4_20_imag;
  reg        [15:0]   int_reg_array_4_21_real;
  reg        [15:0]   int_reg_array_4_21_imag;
  reg        [15:0]   int_reg_array_4_22_real;
  reg        [15:0]   int_reg_array_4_22_imag;
  reg        [15:0]   int_reg_array_4_23_real;
  reg        [15:0]   int_reg_array_4_23_imag;
  reg        [15:0]   int_reg_array_4_24_real;
  reg        [15:0]   int_reg_array_4_24_imag;
  reg        [15:0]   int_reg_array_4_25_real;
  reg        [15:0]   int_reg_array_4_25_imag;
  reg        [15:0]   int_reg_array_4_26_real;
  reg        [15:0]   int_reg_array_4_26_imag;
  reg        [15:0]   int_reg_array_4_27_real;
  reg        [15:0]   int_reg_array_4_27_imag;
  reg        [15:0]   int_reg_array_4_28_real;
  reg        [15:0]   int_reg_array_4_28_imag;
  reg        [15:0]   int_reg_array_4_29_real;
  reg        [15:0]   int_reg_array_4_29_imag;
  reg        [15:0]   int_reg_array_4_30_real;
  reg        [15:0]   int_reg_array_4_30_imag;
  reg        [15:0]   int_reg_array_4_31_real;
  reg        [15:0]   int_reg_array_4_31_imag;
  reg        [15:0]   int_reg_array_4_32_real;
  reg        [15:0]   int_reg_array_4_32_imag;
  reg        [15:0]   int_reg_array_4_33_real;
  reg        [15:0]   int_reg_array_4_33_imag;
  reg        [15:0]   int_reg_array_4_34_real;
  reg        [15:0]   int_reg_array_4_34_imag;
  reg        [15:0]   int_reg_array_4_35_real;
  reg        [15:0]   int_reg_array_4_35_imag;
  reg        [15:0]   int_reg_array_4_36_real;
  reg        [15:0]   int_reg_array_4_36_imag;
  reg        [15:0]   int_reg_array_4_37_real;
  reg        [15:0]   int_reg_array_4_37_imag;
  reg        [15:0]   int_reg_array_4_38_real;
  reg        [15:0]   int_reg_array_4_38_imag;
  reg        [15:0]   int_reg_array_4_39_real;
  reg        [15:0]   int_reg_array_4_39_imag;
  reg        [15:0]   int_reg_array_4_40_real;
  reg        [15:0]   int_reg_array_4_40_imag;
  reg        [15:0]   int_reg_array_4_41_real;
  reg        [15:0]   int_reg_array_4_41_imag;
  reg        [15:0]   int_reg_array_4_42_real;
  reg        [15:0]   int_reg_array_4_42_imag;
  reg        [15:0]   int_reg_array_4_43_real;
  reg        [15:0]   int_reg_array_4_43_imag;
  reg        [15:0]   int_reg_array_4_44_real;
  reg        [15:0]   int_reg_array_4_44_imag;
  reg        [15:0]   int_reg_array_4_45_real;
  reg        [15:0]   int_reg_array_4_45_imag;
  reg        [15:0]   int_reg_array_4_46_real;
  reg        [15:0]   int_reg_array_4_46_imag;
  reg        [15:0]   int_reg_array_4_47_real;
  reg        [15:0]   int_reg_array_4_47_imag;
  reg        [15:0]   int_reg_array_4_48_real;
  reg        [15:0]   int_reg_array_4_48_imag;
  reg        [15:0]   int_reg_array_4_49_real;
  reg        [15:0]   int_reg_array_4_49_imag;
  reg        [15:0]   int_reg_array_4_50_real;
  reg        [15:0]   int_reg_array_4_50_imag;
  reg        [15:0]   int_reg_array_4_51_real;
  reg        [15:0]   int_reg_array_4_51_imag;
  reg        [15:0]   int_reg_array_4_52_real;
  reg        [15:0]   int_reg_array_4_52_imag;
  reg        [15:0]   int_reg_array_4_53_real;
  reg        [15:0]   int_reg_array_4_53_imag;
  reg        [15:0]   int_reg_array_4_54_real;
  reg        [15:0]   int_reg_array_4_54_imag;
  reg        [15:0]   int_reg_array_4_55_real;
  reg        [15:0]   int_reg_array_4_55_imag;
  reg        [15:0]   int_reg_array_4_56_real;
  reg        [15:0]   int_reg_array_4_56_imag;
  reg        [15:0]   int_reg_array_4_57_real;
  reg        [15:0]   int_reg_array_4_57_imag;
  reg        [15:0]   int_reg_array_4_58_real;
  reg        [15:0]   int_reg_array_4_58_imag;
  reg        [15:0]   int_reg_array_4_59_real;
  reg        [15:0]   int_reg_array_4_59_imag;
  reg        [15:0]   int_reg_array_4_60_real;
  reg        [15:0]   int_reg_array_4_60_imag;
  reg        [15:0]   int_reg_array_4_61_real;
  reg        [15:0]   int_reg_array_4_61_imag;
  reg        [15:0]   int_reg_array_4_62_real;
  reg        [15:0]   int_reg_array_4_62_imag;
  reg        [15:0]   int_reg_array_4_63_real;
  reg        [15:0]   int_reg_array_4_63_imag;
  reg        [15:0]   int_reg_array_48_0_real;
  reg        [15:0]   int_reg_array_48_0_imag;
  reg        [15:0]   int_reg_array_48_1_real;
  reg        [15:0]   int_reg_array_48_1_imag;
  reg        [15:0]   int_reg_array_48_2_real;
  reg        [15:0]   int_reg_array_48_2_imag;
  reg        [15:0]   int_reg_array_48_3_real;
  reg        [15:0]   int_reg_array_48_3_imag;
  reg        [15:0]   int_reg_array_48_4_real;
  reg        [15:0]   int_reg_array_48_4_imag;
  reg        [15:0]   int_reg_array_48_5_real;
  reg        [15:0]   int_reg_array_48_5_imag;
  reg        [15:0]   int_reg_array_48_6_real;
  reg        [15:0]   int_reg_array_48_6_imag;
  reg        [15:0]   int_reg_array_48_7_real;
  reg        [15:0]   int_reg_array_48_7_imag;
  reg        [15:0]   int_reg_array_48_8_real;
  reg        [15:0]   int_reg_array_48_8_imag;
  reg        [15:0]   int_reg_array_48_9_real;
  reg        [15:0]   int_reg_array_48_9_imag;
  reg        [15:0]   int_reg_array_48_10_real;
  reg        [15:0]   int_reg_array_48_10_imag;
  reg        [15:0]   int_reg_array_48_11_real;
  reg        [15:0]   int_reg_array_48_11_imag;
  reg        [15:0]   int_reg_array_48_12_real;
  reg        [15:0]   int_reg_array_48_12_imag;
  reg        [15:0]   int_reg_array_48_13_real;
  reg        [15:0]   int_reg_array_48_13_imag;
  reg        [15:0]   int_reg_array_48_14_real;
  reg        [15:0]   int_reg_array_48_14_imag;
  reg        [15:0]   int_reg_array_48_15_real;
  reg        [15:0]   int_reg_array_48_15_imag;
  reg        [15:0]   int_reg_array_48_16_real;
  reg        [15:0]   int_reg_array_48_16_imag;
  reg        [15:0]   int_reg_array_48_17_real;
  reg        [15:0]   int_reg_array_48_17_imag;
  reg        [15:0]   int_reg_array_48_18_real;
  reg        [15:0]   int_reg_array_48_18_imag;
  reg        [15:0]   int_reg_array_48_19_real;
  reg        [15:0]   int_reg_array_48_19_imag;
  reg        [15:0]   int_reg_array_48_20_real;
  reg        [15:0]   int_reg_array_48_20_imag;
  reg        [15:0]   int_reg_array_48_21_real;
  reg        [15:0]   int_reg_array_48_21_imag;
  reg        [15:0]   int_reg_array_48_22_real;
  reg        [15:0]   int_reg_array_48_22_imag;
  reg        [15:0]   int_reg_array_48_23_real;
  reg        [15:0]   int_reg_array_48_23_imag;
  reg        [15:0]   int_reg_array_48_24_real;
  reg        [15:0]   int_reg_array_48_24_imag;
  reg        [15:0]   int_reg_array_48_25_real;
  reg        [15:0]   int_reg_array_48_25_imag;
  reg        [15:0]   int_reg_array_48_26_real;
  reg        [15:0]   int_reg_array_48_26_imag;
  reg        [15:0]   int_reg_array_48_27_real;
  reg        [15:0]   int_reg_array_48_27_imag;
  reg        [15:0]   int_reg_array_48_28_real;
  reg        [15:0]   int_reg_array_48_28_imag;
  reg        [15:0]   int_reg_array_48_29_real;
  reg        [15:0]   int_reg_array_48_29_imag;
  reg        [15:0]   int_reg_array_48_30_real;
  reg        [15:0]   int_reg_array_48_30_imag;
  reg        [15:0]   int_reg_array_48_31_real;
  reg        [15:0]   int_reg_array_48_31_imag;
  reg        [15:0]   int_reg_array_48_32_real;
  reg        [15:0]   int_reg_array_48_32_imag;
  reg        [15:0]   int_reg_array_48_33_real;
  reg        [15:0]   int_reg_array_48_33_imag;
  reg        [15:0]   int_reg_array_48_34_real;
  reg        [15:0]   int_reg_array_48_34_imag;
  reg        [15:0]   int_reg_array_48_35_real;
  reg        [15:0]   int_reg_array_48_35_imag;
  reg        [15:0]   int_reg_array_48_36_real;
  reg        [15:0]   int_reg_array_48_36_imag;
  reg        [15:0]   int_reg_array_48_37_real;
  reg        [15:0]   int_reg_array_48_37_imag;
  reg        [15:0]   int_reg_array_48_38_real;
  reg        [15:0]   int_reg_array_48_38_imag;
  reg        [15:0]   int_reg_array_48_39_real;
  reg        [15:0]   int_reg_array_48_39_imag;
  reg        [15:0]   int_reg_array_48_40_real;
  reg        [15:0]   int_reg_array_48_40_imag;
  reg        [15:0]   int_reg_array_48_41_real;
  reg        [15:0]   int_reg_array_48_41_imag;
  reg        [15:0]   int_reg_array_48_42_real;
  reg        [15:0]   int_reg_array_48_42_imag;
  reg        [15:0]   int_reg_array_48_43_real;
  reg        [15:0]   int_reg_array_48_43_imag;
  reg        [15:0]   int_reg_array_48_44_real;
  reg        [15:0]   int_reg_array_48_44_imag;
  reg        [15:0]   int_reg_array_48_45_real;
  reg        [15:0]   int_reg_array_48_45_imag;
  reg        [15:0]   int_reg_array_48_46_real;
  reg        [15:0]   int_reg_array_48_46_imag;
  reg        [15:0]   int_reg_array_48_47_real;
  reg        [15:0]   int_reg_array_48_47_imag;
  reg        [15:0]   int_reg_array_48_48_real;
  reg        [15:0]   int_reg_array_48_48_imag;
  reg        [15:0]   int_reg_array_48_49_real;
  reg        [15:0]   int_reg_array_48_49_imag;
  reg        [15:0]   int_reg_array_48_50_real;
  reg        [15:0]   int_reg_array_48_50_imag;
  reg        [15:0]   int_reg_array_48_51_real;
  reg        [15:0]   int_reg_array_48_51_imag;
  reg        [15:0]   int_reg_array_48_52_real;
  reg        [15:0]   int_reg_array_48_52_imag;
  reg        [15:0]   int_reg_array_48_53_real;
  reg        [15:0]   int_reg_array_48_53_imag;
  reg        [15:0]   int_reg_array_48_54_real;
  reg        [15:0]   int_reg_array_48_54_imag;
  reg        [15:0]   int_reg_array_48_55_real;
  reg        [15:0]   int_reg_array_48_55_imag;
  reg        [15:0]   int_reg_array_48_56_real;
  reg        [15:0]   int_reg_array_48_56_imag;
  reg        [15:0]   int_reg_array_48_57_real;
  reg        [15:0]   int_reg_array_48_57_imag;
  reg        [15:0]   int_reg_array_48_58_real;
  reg        [15:0]   int_reg_array_48_58_imag;
  reg        [15:0]   int_reg_array_48_59_real;
  reg        [15:0]   int_reg_array_48_59_imag;
  reg        [15:0]   int_reg_array_48_60_real;
  reg        [15:0]   int_reg_array_48_60_imag;
  reg        [15:0]   int_reg_array_48_61_real;
  reg        [15:0]   int_reg_array_48_61_imag;
  reg        [15:0]   int_reg_array_48_62_real;
  reg        [15:0]   int_reg_array_48_62_imag;
  reg        [15:0]   int_reg_array_48_63_real;
  reg        [15:0]   int_reg_array_48_63_imag;
  reg        [15:0]   int_reg_array_2_0_real;
  reg        [15:0]   int_reg_array_2_0_imag;
  reg        [15:0]   int_reg_array_2_1_real;
  reg        [15:0]   int_reg_array_2_1_imag;
  reg        [15:0]   int_reg_array_2_2_real;
  reg        [15:0]   int_reg_array_2_2_imag;
  reg        [15:0]   int_reg_array_2_3_real;
  reg        [15:0]   int_reg_array_2_3_imag;
  reg        [15:0]   int_reg_array_2_4_real;
  reg        [15:0]   int_reg_array_2_4_imag;
  reg        [15:0]   int_reg_array_2_5_real;
  reg        [15:0]   int_reg_array_2_5_imag;
  reg        [15:0]   int_reg_array_2_6_real;
  reg        [15:0]   int_reg_array_2_6_imag;
  reg        [15:0]   int_reg_array_2_7_real;
  reg        [15:0]   int_reg_array_2_7_imag;
  reg        [15:0]   int_reg_array_2_8_real;
  reg        [15:0]   int_reg_array_2_8_imag;
  reg        [15:0]   int_reg_array_2_9_real;
  reg        [15:0]   int_reg_array_2_9_imag;
  reg        [15:0]   int_reg_array_2_10_real;
  reg        [15:0]   int_reg_array_2_10_imag;
  reg        [15:0]   int_reg_array_2_11_real;
  reg        [15:0]   int_reg_array_2_11_imag;
  reg        [15:0]   int_reg_array_2_12_real;
  reg        [15:0]   int_reg_array_2_12_imag;
  reg        [15:0]   int_reg_array_2_13_real;
  reg        [15:0]   int_reg_array_2_13_imag;
  reg        [15:0]   int_reg_array_2_14_real;
  reg        [15:0]   int_reg_array_2_14_imag;
  reg        [15:0]   int_reg_array_2_15_real;
  reg        [15:0]   int_reg_array_2_15_imag;
  reg        [15:0]   int_reg_array_2_16_real;
  reg        [15:0]   int_reg_array_2_16_imag;
  reg        [15:0]   int_reg_array_2_17_real;
  reg        [15:0]   int_reg_array_2_17_imag;
  reg        [15:0]   int_reg_array_2_18_real;
  reg        [15:0]   int_reg_array_2_18_imag;
  reg        [15:0]   int_reg_array_2_19_real;
  reg        [15:0]   int_reg_array_2_19_imag;
  reg        [15:0]   int_reg_array_2_20_real;
  reg        [15:0]   int_reg_array_2_20_imag;
  reg        [15:0]   int_reg_array_2_21_real;
  reg        [15:0]   int_reg_array_2_21_imag;
  reg        [15:0]   int_reg_array_2_22_real;
  reg        [15:0]   int_reg_array_2_22_imag;
  reg        [15:0]   int_reg_array_2_23_real;
  reg        [15:0]   int_reg_array_2_23_imag;
  reg        [15:0]   int_reg_array_2_24_real;
  reg        [15:0]   int_reg_array_2_24_imag;
  reg        [15:0]   int_reg_array_2_25_real;
  reg        [15:0]   int_reg_array_2_25_imag;
  reg        [15:0]   int_reg_array_2_26_real;
  reg        [15:0]   int_reg_array_2_26_imag;
  reg        [15:0]   int_reg_array_2_27_real;
  reg        [15:0]   int_reg_array_2_27_imag;
  reg        [15:0]   int_reg_array_2_28_real;
  reg        [15:0]   int_reg_array_2_28_imag;
  reg        [15:0]   int_reg_array_2_29_real;
  reg        [15:0]   int_reg_array_2_29_imag;
  reg        [15:0]   int_reg_array_2_30_real;
  reg        [15:0]   int_reg_array_2_30_imag;
  reg        [15:0]   int_reg_array_2_31_real;
  reg        [15:0]   int_reg_array_2_31_imag;
  reg        [15:0]   int_reg_array_2_32_real;
  reg        [15:0]   int_reg_array_2_32_imag;
  reg        [15:0]   int_reg_array_2_33_real;
  reg        [15:0]   int_reg_array_2_33_imag;
  reg        [15:0]   int_reg_array_2_34_real;
  reg        [15:0]   int_reg_array_2_34_imag;
  reg        [15:0]   int_reg_array_2_35_real;
  reg        [15:0]   int_reg_array_2_35_imag;
  reg        [15:0]   int_reg_array_2_36_real;
  reg        [15:0]   int_reg_array_2_36_imag;
  reg        [15:0]   int_reg_array_2_37_real;
  reg        [15:0]   int_reg_array_2_37_imag;
  reg        [15:0]   int_reg_array_2_38_real;
  reg        [15:0]   int_reg_array_2_38_imag;
  reg        [15:0]   int_reg_array_2_39_real;
  reg        [15:0]   int_reg_array_2_39_imag;
  reg        [15:0]   int_reg_array_2_40_real;
  reg        [15:0]   int_reg_array_2_40_imag;
  reg        [15:0]   int_reg_array_2_41_real;
  reg        [15:0]   int_reg_array_2_41_imag;
  reg        [15:0]   int_reg_array_2_42_real;
  reg        [15:0]   int_reg_array_2_42_imag;
  reg        [15:0]   int_reg_array_2_43_real;
  reg        [15:0]   int_reg_array_2_43_imag;
  reg        [15:0]   int_reg_array_2_44_real;
  reg        [15:0]   int_reg_array_2_44_imag;
  reg        [15:0]   int_reg_array_2_45_real;
  reg        [15:0]   int_reg_array_2_45_imag;
  reg        [15:0]   int_reg_array_2_46_real;
  reg        [15:0]   int_reg_array_2_46_imag;
  reg        [15:0]   int_reg_array_2_47_real;
  reg        [15:0]   int_reg_array_2_47_imag;
  reg        [15:0]   int_reg_array_2_48_real;
  reg        [15:0]   int_reg_array_2_48_imag;
  reg        [15:0]   int_reg_array_2_49_real;
  reg        [15:0]   int_reg_array_2_49_imag;
  reg        [15:0]   int_reg_array_2_50_real;
  reg        [15:0]   int_reg_array_2_50_imag;
  reg        [15:0]   int_reg_array_2_51_real;
  reg        [15:0]   int_reg_array_2_51_imag;
  reg        [15:0]   int_reg_array_2_52_real;
  reg        [15:0]   int_reg_array_2_52_imag;
  reg        [15:0]   int_reg_array_2_53_real;
  reg        [15:0]   int_reg_array_2_53_imag;
  reg        [15:0]   int_reg_array_2_54_real;
  reg        [15:0]   int_reg_array_2_54_imag;
  reg        [15:0]   int_reg_array_2_55_real;
  reg        [15:0]   int_reg_array_2_55_imag;
  reg        [15:0]   int_reg_array_2_56_real;
  reg        [15:0]   int_reg_array_2_56_imag;
  reg        [15:0]   int_reg_array_2_57_real;
  reg        [15:0]   int_reg_array_2_57_imag;
  reg        [15:0]   int_reg_array_2_58_real;
  reg        [15:0]   int_reg_array_2_58_imag;
  reg        [15:0]   int_reg_array_2_59_real;
  reg        [15:0]   int_reg_array_2_59_imag;
  reg        [15:0]   int_reg_array_2_60_real;
  reg        [15:0]   int_reg_array_2_60_imag;
  reg        [15:0]   int_reg_array_2_61_real;
  reg        [15:0]   int_reg_array_2_61_imag;
  reg        [15:0]   int_reg_array_2_62_real;
  reg        [15:0]   int_reg_array_2_62_imag;
  reg        [15:0]   int_reg_array_2_63_real;
  reg        [15:0]   int_reg_array_2_63_imag;
  reg        [15:0]   int_reg_array_62_0_real;
  reg        [15:0]   int_reg_array_62_0_imag;
  reg        [15:0]   int_reg_array_62_1_real;
  reg        [15:0]   int_reg_array_62_1_imag;
  reg        [15:0]   int_reg_array_62_2_real;
  reg        [15:0]   int_reg_array_62_2_imag;
  reg        [15:0]   int_reg_array_62_3_real;
  reg        [15:0]   int_reg_array_62_3_imag;
  reg        [15:0]   int_reg_array_62_4_real;
  reg        [15:0]   int_reg_array_62_4_imag;
  reg        [15:0]   int_reg_array_62_5_real;
  reg        [15:0]   int_reg_array_62_5_imag;
  reg        [15:0]   int_reg_array_62_6_real;
  reg        [15:0]   int_reg_array_62_6_imag;
  reg        [15:0]   int_reg_array_62_7_real;
  reg        [15:0]   int_reg_array_62_7_imag;
  reg        [15:0]   int_reg_array_62_8_real;
  reg        [15:0]   int_reg_array_62_8_imag;
  reg        [15:0]   int_reg_array_62_9_real;
  reg        [15:0]   int_reg_array_62_9_imag;
  reg        [15:0]   int_reg_array_62_10_real;
  reg        [15:0]   int_reg_array_62_10_imag;
  reg        [15:0]   int_reg_array_62_11_real;
  reg        [15:0]   int_reg_array_62_11_imag;
  reg        [15:0]   int_reg_array_62_12_real;
  reg        [15:0]   int_reg_array_62_12_imag;
  reg        [15:0]   int_reg_array_62_13_real;
  reg        [15:0]   int_reg_array_62_13_imag;
  reg        [15:0]   int_reg_array_62_14_real;
  reg        [15:0]   int_reg_array_62_14_imag;
  reg        [15:0]   int_reg_array_62_15_real;
  reg        [15:0]   int_reg_array_62_15_imag;
  reg        [15:0]   int_reg_array_62_16_real;
  reg        [15:0]   int_reg_array_62_16_imag;
  reg        [15:0]   int_reg_array_62_17_real;
  reg        [15:0]   int_reg_array_62_17_imag;
  reg        [15:0]   int_reg_array_62_18_real;
  reg        [15:0]   int_reg_array_62_18_imag;
  reg        [15:0]   int_reg_array_62_19_real;
  reg        [15:0]   int_reg_array_62_19_imag;
  reg        [15:0]   int_reg_array_62_20_real;
  reg        [15:0]   int_reg_array_62_20_imag;
  reg        [15:0]   int_reg_array_62_21_real;
  reg        [15:0]   int_reg_array_62_21_imag;
  reg        [15:0]   int_reg_array_62_22_real;
  reg        [15:0]   int_reg_array_62_22_imag;
  reg        [15:0]   int_reg_array_62_23_real;
  reg        [15:0]   int_reg_array_62_23_imag;
  reg        [15:0]   int_reg_array_62_24_real;
  reg        [15:0]   int_reg_array_62_24_imag;
  reg        [15:0]   int_reg_array_62_25_real;
  reg        [15:0]   int_reg_array_62_25_imag;
  reg        [15:0]   int_reg_array_62_26_real;
  reg        [15:0]   int_reg_array_62_26_imag;
  reg        [15:0]   int_reg_array_62_27_real;
  reg        [15:0]   int_reg_array_62_27_imag;
  reg        [15:0]   int_reg_array_62_28_real;
  reg        [15:0]   int_reg_array_62_28_imag;
  reg        [15:0]   int_reg_array_62_29_real;
  reg        [15:0]   int_reg_array_62_29_imag;
  reg        [15:0]   int_reg_array_62_30_real;
  reg        [15:0]   int_reg_array_62_30_imag;
  reg        [15:0]   int_reg_array_62_31_real;
  reg        [15:0]   int_reg_array_62_31_imag;
  reg        [15:0]   int_reg_array_62_32_real;
  reg        [15:0]   int_reg_array_62_32_imag;
  reg        [15:0]   int_reg_array_62_33_real;
  reg        [15:0]   int_reg_array_62_33_imag;
  reg        [15:0]   int_reg_array_62_34_real;
  reg        [15:0]   int_reg_array_62_34_imag;
  reg        [15:0]   int_reg_array_62_35_real;
  reg        [15:0]   int_reg_array_62_35_imag;
  reg        [15:0]   int_reg_array_62_36_real;
  reg        [15:0]   int_reg_array_62_36_imag;
  reg        [15:0]   int_reg_array_62_37_real;
  reg        [15:0]   int_reg_array_62_37_imag;
  reg        [15:0]   int_reg_array_62_38_real;
  reg        [15:0]   int_reg_array_62_38_imag;
  reg        [15:0]   int_reg_array_62_39_real;
  reg        [15:0]   int_reg_array_62_39_imag;
  reg        [15:0]   int_reg_array_62_40_real;
  reg        [15:0]   int_reg_array_62_40_imag;
  reg        [15:0]   int_reg_array_62_41_real;
  reg        [15:0]   int_reg_array_62_41_imag;
  reg        [15:0]   int_reg_array_62_42_real;
  reg        [15:0]   int_reg_array_62_42_imag;
  reg        [15:0]   int_reg_array_62_43_real;
  reg        [15:0]   int_reg_array_62_43_imag;
  reg        [15:0]   int_reg_array_62_44_real;
  reg        [15:0]   int_reg_array_62_44_imag;
  reg        [15:0]   int_reg_array_62_45_real;
  reg        [15:0]   int_reg_array_62_45_imag;
  reg        [15:0]   int_reg_array_62_46_real;
  reg        [15:0]   int_reg_array_62_46_imag;
  reg        [15:0]   int_reg_array_62_47_real;
  reg        [15:0]   int_reg_array_62_47_imag;
  reg        [15:0]   int_reg_array_62_48_real;
  reg        [15:0]   int_reg_array_62_48_imag;
  reg        [15:0]   int_reg_array_62_49_real;
  reg        [15:0]   int_reg_array_62_49_imag;
  reg        [15:0]   int_reg_array_62_50_real;
  reg        [15:0]   int_reg_array_62_50_imag;
  reg        [15:0]   int_reg_array_62_51_real;
  reg        [15:0]   int_reg_array_62_51_imag;
  reg        [15:0]   int_reg_array_62_52_real;
  reg        [15:0]   int_reg_array_62_52_imag;
  reg        [15:0]   int_reg_array_62_53_real;
  reg        [15:0]   int_reg_array_62_53_imag;
  reg        [15:0]   int_reg_array_62_54_real;
  reg        [15:0]   int_reg_array_62_54_imag;
  reg        [15:0]   int_reg_array_62_55_real;
  reg        [15:0]   int_reg_array_62_55_imag;
  reg        [15:0]   int_reg_array_62_56_real;
  reg        [15:0]   int_reg_array_62_56_imag;
  reg        [15:0]   int_reg_array_62_57_real;
  reg        [15:0]   int_reg_array_62_57_imag;
  reg        [15:0]   int_reg_array_62_58_real;
  reg        [15:0]   int_reg_array_62_58_imag;
  reg        [15:0]   int_reg_array_62_59_real;
  reg        [15:0]   int_reg_array_62_59_imag;
  reg        [15:0]   int_reg_array_62_60_real;
  reg        [15:0]   int_reg_array_62_60_imag;
  reg        [15:0]   int_reg_array_62_61_real;
  reg        [15:0]   int_reg_array_62_61_imag;
  reg        [15:0]   int_reg_array_62_62_real;
  reg        [15:0]   int_reg_array_62_62_imag;
  reg        [15:0]   int_reg_array_62_63_real;
  reg        [15:0]   int_reg_array_62_63_imag;
  reg        [15:0]   int_reg_array_56_0_real;
  reg        [15:0]   int_reg_array_56_0_imag;
  reg        [15:0]   int_reg_array_56_1_real;
  reg        [15:0]   int_reg_array_56_1_imag;
  reg        [15:0]   int_reg_array_56_2_real;
  reg        [15:0]   int_reg_array_56_2_imag;
  reg        [15:0]   int_reg_array_56_3_real;
  reg        [15:0]   int_reg_array_56_3_imag;
  reg        [15:0]   int_reg_array_56_4_real;
  reg        [15:0]   int_reg_array_56_4_imag;
  reg        [15:0]   int_reg_array_56_5_real;
  reg        [15:0]   int_reg_array_56_5_imag;
  reg        [15:0]   int_reg_array_56_6_real;
  reg        [15:0]   int_reg_array_56_6_imag;
  reg        [15:0]   int_reg_array_56_7_real;
  reg        [15:0]   int_reg_array_56_7_imag;
  reg        [15:0]   int_reg_array_56_8_real;
  reg        [15:0]   int_reg_array_56_8_imag;
  reg        [15:0]   int_reg_array_56_9_real;
  reg        [15:0]   int_reg_array_56_9_imag;
  reg        [15:0]   int_reg_array_56_10_real;
  reg        [15:0]   int_reg_array_56_10_imag;
  reg        [15:0]   int_reg_array_56_11_real;
  reg        [15:0]   int_reg_array_56_11_imag;
  reg        [15:0]   int_reg_array_56_12_real;
  reg        [15:0]   int_reg_array_56_12_imag;
  reg        [15:0]   int_reg_array_56_13_real;
  reg        [15:0]   int_reg_array_56_13_imag;
  reg        [15:0]   int_reg_array_56_14_real;
  reg        [15:0]   int_reg_array_56_14_imag;
  reg        [15:0]   int_reg_array_56_15_real;
  reg        [15:0]   int_reg_array_56_15_imag;
  reg        [15:0]   int_reg_array_56_16_real;
  reg        [15:0]   int_reg_array_56_16_imag;
  reg        [15:0]   int_reg_array_56_17_real;
  reg        [15:0]   int_reg_array_56_17_imag;
  reg        [15:0]   int_reg_array_56_18_real;
  reg        [15:0]   int_reg_array_56_18_imag;
  reg        [15:0]   int_reg_array_56_19_real;
  reg        [15:0]   int_reg_array_56_19_imag;
  reg        [15:0]   int_reg_array_56_20_real;
  reg        [15:0]   int_reg_array_56_20_imag;
  reg        [15:0]   int_reg_array_56_21_real;
  reg        [15:0]   int_reg_array_56_21_imag;
  reg        [15:0]   int_reg_array_56_22_real;
  reg        [15:0]   int_reg_array_56_22_imag;
  reg        [15:0]   int_reg_array_56_23_real;
  reg        [15:0]   int_reg_array_56_23_imag;
  reg        [15:0]   int_reg_array_56_24_real;
  reg        [15:0]   int_reg_array_56_24_imag;
  reg        [15:0]   int_reg_array_56_25_real;
  reg        [15:0]   int_reg_array_56_25_imag;
  reg        [15:0]   int_reg_array_56_26_real;
  reg        [15:0]   int_reg_array_56_26_imag;
  reg        [15:0]   int_reg_array_56_27_real;
  reg        [15:0]   int_reg_array_56_27_imag;
  reg        [15:0]   int_reg_array_56_28_real;
  reg        [15:0]   int_reg_array_56_28_imag;
  reg        [15:0]   int_reg_array_56_29_real;
  reg        [15:0]   int_reg_array_56_29_imag;
  reg        [15:0]   int_reg_array_56_30_real;
  reg        [15:0]   int_reg_array_56_30_imag;
  reg        [15:0]   int_reg_array_56_31_real;
  reg        [15:0]   int_reg_array_56_31_imag;
  reg        [15:0]   int_reg_array_56_32_real;
  reg        [15:0]   int_reg_array_56_32_imag;
  reg        [15:0]   int_reg_array_56_33_real;
  reg        [15:0]   int_reg_array_56_33_imag;
  reg        [15:0]   int_reg_array_56_34_real;
  reg        [15:0]   int_reg_array_56_34_imag;
  reg        [15:0]   int_reg_array_56_35_real;
  reg        [15:0]   int_reg_array_56_35_imag;
  reg        [15:0]   int_reg_array_56_36_real;
  reg        [15:0]   int_reg_array_56_36_imag;
  reg        [15:0]   int_reg_array_56_37_real;
  reg        [15:0]   int_reg_array_56_37_imag;
  reg        [15:0]   int_reg_array_56_38_real;
  reg        [15:0]   int_reg_array_56_38_imag;
  reg        [15:0]   int_reg_array_56_39_real;
  reg        [15:0]   int_reg_array_56_39_imag;
  reg        [15:0]   int_reg_array_56_40_real;
  reg        [15:0]   int_reg_array_56_40_imag;
  reg        [15:0]   int_reg_array_56_41_real;
  reg        [15:0]   int_reg_array_56_41_imag;
  reg        [15:0]   int_reg_array_56_42_real;
  reg        [15:0]   int_reg_array_56_42_imag;
  reg        [15:0]   int_reg_array_56_43_real;
  reg        [15:0]   int_reg_array_56_43_imag;
  reg        [15:0]   int_reg_array_56_44_real;
  reg        [15:0]   int_reg_array_56_44_imag;
  reg        [15:0]   int_reg_array_56_45_real;
  reg        [15:0]   int_reg_array_56_45_imag;
  reg        [15:0]   int_reg_array_56_46_real;
  reg        [15:0]   int_reg_array_56_46_imag;
  reg        [15:0]   int_reg_array_56_47_real;
  reg        [15:0]   int_reg_array_56_47_imag;
  reg        [15:0]   int_reg_array_56_48_real;
  reg        [15:0]   int_reg_array_56_48_imag;
  reg        [15:0]   int_reg_array_56_49_real;
  reg        [15:0]   int_reg_array_56_49_imag;
  reg        [15:0]   int_reg_array_56_50_real;
  reg        [15:0]   int_reg_array_56_50_imag;
  reg        [15:0]   int_reg_array_56_51_real;
  reg        [15:0]   int_reg_array_56_51_imag;
  reg        [15:0]   int_reg_array_56_52_real;
  reg        [15:0]   int_reg_array_56_52_imag;
  reg        [15:0]   int_reg_array_56_53_real;
  reg        [15:0]   int_reg_array_56_53_imag;
  reg        [15:0]   int_reg_array_56_54_real;
  reg        [15:0]   int_reg_array_56_54_imag;
  reg        [15:0]   int_reg_array_56_55_real;
  reg        [15:0]   int_reg_array_56_55_imag;
  reg        [15:0]   int_reg_array_56_56_real;
  reg        [15:0]   int_reg_array_56_56_imag;
  reg        [15:0]   int_reg_array_56_57_real;
  reg        [15:0]   int_reg_array_56_57_imag;
  reg        [15:0]   int_reg_array_56_58_real;
  reg        [15:0]   int_reg_array_56_58_imag;
  reg        [15:0]   int_reg_array_56_59_real;
  reg        [15:0]   int_reg_array_56_59_imag;
  reg        [15:0]   int_reg_array_56_60_real;
  reg        [15:0]   int_reg_array_56_60_imag;
  reg        [15:0]   int_reg_array_56_61_real;
  reg        [15:0]   int_reg_array_56_61_imag;
  reg        [15:0]   int_reg_array_56_62_real;
  reg        [15:0]   int_reg_array_56_62_imag;
  reg        [15:0]   int_reg_array_56_63_real;
  reg        [15:0]   int_reg_array_56_63_imag;
  reg        [15:0]   int_reg_array_18_0_real;
  reg        [15:0]   int_reg_array_18_0_imag;
  reg        [15:0]   int_reg_array_18_1_real;
  reg        [15:0]   int_reg_array_18_1_imag;
  reg        [15:0]   int_reg_array_18_2_real;
  reg        [15:0]   int_reg_array_18_2_imag;
  reg        [15:0]   int_reg_array_18_3_real;
  reg        [15:0]   int_reg_array_18_3_imag;
  reg        [15:0]   int_reg_array_18_4_real;
  reg        [15:0]   int_reg_array_18_4_imag;
  reg        [15:0]   int_reg_array_18_5_real;
  reg        [15:0]   int_reg_array_18_5_imag;
  reg        [15:0]   int_reg_array_18_6_real;
  reg        [15:0]   int_reg_array_18_6_imag;
  reg        [15:0]   int_reg_array_18_7_real;
  reg        [15:0]   int_reg_array_18_7_imag;
  reg        [15:0]   int_reg_array_18_8_real;
  reg        [15:0]   int_reg_array_18_8_imag;
  reg        [15:0]   int_reg_array_18_9_real;
  reg        [15:0]   int_reg_array_18_9_imag;
  reg        [15:0]   int_reg_array_18_10_real;
  reg        [15:0]   int_reg_array_18_10_imag;
  reg        [15:0]   int_reg_array_18_11_real;
  reg        [15:0]   int_reg_array_18_11_imag;
  reg        [15:0]   int_reg_array_18_12_real;
  reg        [15:0]   int_reg_array_18_12_imag;
  reg        [15:0]   int_reg_array_18_13_real;
  reg        [15:0]   int_reg_array_18_13_imag;
  reg        [15:0]   int_reg_array_18_14_real;
  reg        [15:0]   int_reg_array_18_14_imag;
  reg        [15:0]   int_reg_array_18_15_real;
  reg        [15:0]   int_reg_array_18_15_imag;
  reg        [15:0]   int_reg_array_18_16_real;
  reg        [15:0]   int_reg_array_18_16_imag;
  reg        [15:0]   int_reg_array_18_17_real;
  reg        [15:0]   int_reg_array_18_17_imag;
  reg        [15:0]   int_reg_array_18_18_real;
  reg        [15:0]   int_reg_array_18_18_imag;
  reg        [15:0]   int_reg_array_18_19_real;
  reg        [15:0]   int_reg_array_18_19_imag;
  reg        [15:0]   int_reg_array_18_20_real;
  reg        [15:0]   int_reg_array_18_20_imag;
  reg        [15:0]   int_reg_array_18_21_real;
  reg        [15:0]   int_reg_array_18_21_imag;
  reg        [15:0]   int_reg_array_18_22_real;
  reg        [15:0]   int_reg_array_18_22_imag;
  reg        [15:0]   int_reg_array_18_23_real;
  reg        [15:0]   int_reg_array_18_23_imag;
  reg        [15:0]   int_reg_array_18_24_real;
  reg        [15:0]   int_reg_array_18_24_imag;
  reg        [15:0]   int_reg_array_18_25_real;
  reg        [15:0]   int_reg_array_18_25_imag;
  reg        [15:0]   int_reg_array_18_26_real;
  reg        [15:0]   int_reg_array_18_26_imag;
  reg        [15:0]   int_reg_array_18_27_real;
  reg        [15:0]   int_reg_array_18_27_imag;
  reg        [15:0]   int_reg_array_18_28_real;
  reg        [15:0]   int_reg_array_18_28_imag;
  reg        [15:0]   int_reg_array_18_29_real;
  reg        [15:0]   int_reg_array_18_29_imag;
  reg        [15:0]   int_reg_array_18_30_real;
  reg        [15:0]   int_reg_array_18_30_imag;
  reg        [15:0]   int_reg_array_18_31_real;
  reg        [15:0]   int_reg_array_18_31_imag;
  reg        [15:0]   int_reg_array_18_32_real;
  reg        [15:0]   int_reg_array_18_32_imag;
  reg        [15:0]   int_reg_array_18_33_real;
  reg        [15:0]   int_reg_array_18_33_imag;
  reg        [15:0]   int_reg_array_18_34_real;
  reg        [15:0]   int_reg_array_18_34_imag;
  reg        [15:0]   int_reg_array_18_35_real;
  reg        [15:0]   int_reg_array_18_35_imag;
  reg        [15:0]   int_reg_array_18_36_real;
  reg        [15:0]   int_reg_array_18_36_imag;
  reg        [15:0]   int_reg_array_18_37_real;
  reg        [15:0]   int_reg_array_18_37_imag;
  reg        [15:0]   int_reg_array_18_38_real;
  reg        [15:0]   int_reg_array_18_38_imag;
  reg        [15:0]   int_reg_array_18_39_real;
  reg        [15:0]   int_reg_array_18_39_imag;
  reg        [15:0]   int_reg_array_18_40_real;
  reg        [15:0]   int_reg_array_18_40_imag;
  reg        [15:0]   int_reg_array_18_41_real;
  reg        [15:0]   int_reg_array_18_41_imag;
  reg        [15:0]   int_reg_array_18_42_real;
  reg        [15:0]   int_reg_array_18_42_imag;
  reg        [15:0]   int_reg_array_18_43_real;
  reg        [15:0]   int_reg_array_18_43_imag;
  reg        [15:0]   int_reg_array_18_44_real;
  reg        [15:0]   int_reg_array_18_44_imag;
  reg        [15:0]   int_reg_array_18_45_real;
  reg        [15:0]   int_reg_array_18_45_imag;
  reg        [15:0]   int_reg_array_18_46_real;
  reg        [15:0]   int_reg_array_18_46_imag;
  reg        [15:0]   int_reg_array_18_47_real;
  reg        [15:0]   int_reg_array_18_47_imag;
  reg        [15:0]   int_reg_array_18_48_real;
  reg        [15:0]   int_reg_array_18_48_imag;
  reg        [15:0]   int_reg_array_18_49_real;
  reg        [15:0]   int_reg_array_18_49_imag;
  reg        [15:0]   int_reg_array_18_50_real;
  reg        [15:0]   int_reg_array_18_50_imag;
  reg        [15:0]   int_reg_array_18_51_real;
  reg        [15:0]   int_reg_array_18_51_imag;
  reg        [15:0]   int_reg_array_18_52_real;
  reg        [15:0]   int_reg_array_18_52_imag;
  reg        [15:0]   int_reg_array_18_53_real;
  reg        [15:0]   int_reg_array_18_53_imag;
  reg        [15:0]   int_reg_array_18_54_real;
  reg        [15:0]   int_reg_array_18_54_imag;
  reg        [15:0]   int_reg_array_18_55_real;
  reg        [15:0]   int_reg_array_18_55_imag;
  reg        [15:0]   int_reg_array_18_56_real;
  reg        [15:0]   int_reg_array_18_56_imag;
  reg        [15:0]   int_reg_array_18_57_real;
  reg        [15:0]   int_reg_array_18_57_imag;
  reg        [15:0]   int_reg_array_18_58_real;
  reg        [15:0]   int_reg_array_18_58_imag;
  reg        [15:0]   int_reg_array_18_59_real;
  reg        [15:0]   int_reg_array_18_59_imag;
  reg        [15:0]   int_reg_array_18_60_real;
  reg        [15:0]   int_reg_array_18_60_imag;
  reg        [15:0]   int_reg_array_18_61_real;
  reg        [15:0]   int_reg_array_18_61_imag;
  reg        [15:0]   int_reg_array_18_62_real;
  reg        [15:0]   int_reg_array_18_62_imag;
  reg        [15:0]   int_reg_array_18_63_real;
  reg        [15:0]   int_reg_array_18_63_imag;
  reg        [15:0]   int_reg_array_6_0_real;
  reg        [15:0]   int_reg_array_6_0_imag;
  reg        [15:0]   int_reg_array_6_1_real;
  reg        [15:0]   int_reg_array_6_1_imag;
  reg        [15:0]   int_reg_array_6_2_real;
  reg        [15:0]   int_reg_array_6_2_imag;
  reg        [15:0]   int_reg_array_6_3_real;
  reg        [15:0]   int_reg_array_6_3_imag;
  reg        [15:0]   int_reg_array_6_4_real;
  reg        [15:0]   int_reg_array_6_4_imag;
  reg        [15:0]   int_reg_array_6_5_real;
  reg        [15:0]   int_reg_array_6_5_imag;
  reg        [15:0]   int_reg_array_6_6_real;
  reg        [15:0]   int_reg_array_6_6_imag;
  reg        [15:0]   int_reg_array_6_7_real;
  reg        [15:0]   int_reg_array_6_7_imag;
  reg        [15:0]   int_reg_array_6_8_real;
  reg        [15:0]   int_reg_array_6_8_imag;
  reg        [15:0]   int_reg_array_6_9_real;
  reg        [15:0]   int_reg_array_6_9_imag;
  reg        [15:0]   int_reg_array_6_10_real;
  reg        [15:0]   int_reg_array_6_10_imag;
  reg        [15:0]   int_reg_array_6_11_real;
  reg        [15:0]   int_reg_array_6_11_imag;
  reg        [15:0]   int_reg_array_6_12_real;
  reg        [15:0]   int_reg_array_6_12_imag;
  reg        [15:0]   int_reg_array_6_13_real;
  reg        [15:0]   int_reg_array_6_13_imag;
  reg        [15:0]   int_reg_array_6_14_real;
  reg        [15:0]   int_reg_array_6_14_imag;
  reg        [15:0]   int_reg_array_6_15_real;
  reg        [15:0]   int_reg_array_6_15_imag;
  reg        [15:0]   int_reg_array_6_16_real;
  reg        [15:0]   int_reg_array_6_16_imag;
  reg        [15:0]   int_reg_array_6_17_real;
  reg        [15:0]   int_reg_array_6_17_imag;
  reg        [15:0]   int_reg_array_6_18_real;
  reg        [15:0]   int_reg_array_6_18_imag;
  reg        [15:0]   int_reg_array_6_19_real;
  reg        [15:0]   int_reg_array_6_19_imag;
  reg        [15:0]   int_reg_array_6_20_real;
  reg        [15:0]   int_reg_array_6_20_imag;
  reg        [15:0]   int_reg_array_6_21_real;
  reg        [15:0]   int_reg_array_6_21_imag;
  reg        [15:0]   int_reg_array_6_22_real;
  reg        [15:0]   int_reg_array_6_22_imag;
  reg        [15:0]   int_reg_array_6_23_real;
  reg        [15:0]   int_reg_array_6_23_imag;
  reg        [15:0]   int_reg_array_6_24_real;
  reg        [15:0]   int_reg_array_6_24_imag;
  reg        [15:0]   int_reg_array_6_25_real;
  reg        [15:0]   int_reg_array_6_25_imag;
  reg        [15:0]   int_reg_array_6_26_real;
  reg        [15:0]   int_reg_array_6_26_imag;
  reg        [15:0]   int_reg_array_6_27_real;
  reg        [15:0]   int_reg_array_6_27_imag;
  reg        [15:0]   int_reg_array_6_28_real;
  reg        [15:0]   int_reg_array_6_28_imag;
  reg        [15:0]   int_reg_array_6_29_real;
  reg        [15:0]   int_reg_array_6_29_imag;
  reg        [15:0]   int_reg_array_6_30_real;
  reg        [15:0]   int_reg_array_6_30_imag;
  reg        [15:0]   int_reg_array_6_31_real;
  reg        [15:0]   int_reg_array_6_31_imag;
  reg        [15:0]   int_reg_array_6_32_real;
  reg        [15:0]   int_reg_array_6_32_imag;
  reg        [15:0]   int_reg_array_6_33_real;
  reg        [15:0]   int_reg_array_6_33_imag;
  reg        [15:0]   int_reg_array_6_34_real;
  reg        [15:0]   int_reg_array_6_34_imag;
  reg        [15:0]   int_reg_array_6_35_real;
  reg        [15:0]   int_reg_array_6_35_imag;
  reg        [15:0]   int_reg_array_6_36_real;
  reg        [15:0]   int_reg_array_6_36_imag;
  reg        [15:0]   int_reg_array_6_37_real;
  reg        [15:0]   int_reg_array_6_37_imag;
  reg        [15:0]   int_reg_array_6_38_real;
  reg        [15:0]   int_reg_array_6_38_imag;
  reg        [15:0]   int_reg_array_6_39_real;
  reg        [15:0]   int_reg_array_6_39_imag;
  reg        [15:0]   int_reg_array_6_40_real;
  reg        [15:0]   int_reg_array_6_40_imag;
  reg        [15:0]   int_reg_array_6_41_real;
  reg        [15:0]   int_reg_array_6_41_imag;
  reg        [15:0]   int_reg_array_6_42_real;
  reg        [15:0]   int_reg_array_6_42_imag;
  reg        [15:0]   int_reg_array_6_43_real;
  reg        [15:0]   int_reg_array_6_43_imag;
  reg        [15:0]   int_reg_array_6_44_real;
  reg        [15:0]   int_reg_array_6_44_imag;
  reg        [15:0]   int_reg_array_6_45_real;
  reg        [15:0]   int_reg_array_6_45_imag;
  reg        [15:0]   int_reg_array_6_46_real;
  reg        [15:0]   int_reg_array_6_46_imag;
  reg        [15:0]   int_reg_array_6_47_real;
  reg        [15:0]   int_reg_array_6_47_imag;
  reg        [15:0]   int_reg_array_6_48_real;
  reg        [15:0]   int_reg_array_6_48_imag;
  reg        [15:0]   int_reg_array_6_49_real;
  reg        [15:0]   int_reg_array_6_49_imag;
  reg        [15:0]   int_reg_array_6_50_real;
  reg        [15:0]   int_reg_array_6_50_imag;
  reg        [15:0]   int_reg_array_6_51_real;
  reg        [15:0]   int_reg_array_6_51_imag;
  reg        [15:0]   int_reg_array_6_52_real;
  reg        [15:0]   int_reg_array_6_52_imag;
  reg        [15:0]   int_reg_array_6_53_real;
  reg        [15:0]   int_reg_array_6_53_imag;
  reg        [15:0]   int_reg_array_6_54_real;
  reg        [15:0]   int_reg_array_6_54_imag;
  reg        [15:0]   int_reg_array_6_55_real;
  reg        [15:0]   int_reg_array_6_55_imag;
  reg        [15:0]   int_reg_array_6_56_real;
  reg        [15:0]   int_reg_array_6_56_imag;
  reg        [15:0]   int_reg_array_6_57_real;
  reg        [15:0]   int_reg_array_6_57_imag;
  reg        [15:0]   int_reg_array_6_58_real;
  reg        [15:0]   int_reg_array_6_58_imag;
  reg        [15:0]   int_reg_array_6_59_real;
  reg        [15:0]   int_reg_array_6_59_imag;
  reg        [15:0]   int_reg_array_6_60_real;
  reg        [15:0]   int_reg_array_6_60_imag;
  reg        [15:0]   int_reg_array_6_61_real;
  reg        [15:0]   int_reg_array_6_61_imag;
  reg        [15:0]   int_reg_array_6_62_real;
  reg        [15:0]   int_reg_array_6_62_imag;
  reg        [15:0]   int_reg_array_6_63_real;
  reg        [15:0]   int_reg_array_6_63_imag;
  reg        [15:0]   int_reg_array_50_0_real;
  reg        [15:0]   int_reg_array_50_0_imag;
  reg        [15:0]   int_reg_array_50_1_real;
  reg        [15:0]   int_reg_array_50_1_imag;
  reg        [15:0]   int_reg_array_50_2_real;
  reg        [15:0]   int_reg_array_50_2_imag;
  reg        [15:0]   int_reg_array_50_3_real;
  reg        [15:0]   int_reg_array_50_3_imag;
  reg        [15:0]   int_reg_array_50_4_real;
  reg        [15:0]   int_reg_array_50_4_imag;
  reg        [15:0]   int_reg_array_50_5_real;
  reg        [15:0]   int_reg_array_50_5_imag;
  reg        [15:0]   int_reg_array_50_6_real;
  reg        [15:0]   int_reg_array_50_6_imag;
  reg        [15:0]   int_reg_array_50_7_real;
  reg        [15:0]   int_reg_array_50_7_imag;
  reg        [15:0]   int_reg_array_50_8_real;
  reg        [15:0]   int_reg_array_50_8_imag;
  reg        [15:0]   int_reg_array_50_9_real;
  reg        [15:0]   int_reg_array_50_9_imag;
  reg        [15:0]   int_reg_array_50_10_real;
  reg        [15:0]   int_reg_array_50_10_imag;
  reg        [15:0]   int_reg_array_50_11_real;
  reg        [15:0]   int_reg_array_50_11_imag;
  reg        [15:0]   int_reg_array_50_12_real;
  reg        [15:0]   int_reg_array_50_12_imag;
  reg        [15:0]   int_reg_array_50_13_real;
  reg        [15:0]   int_reg_array_50_13_imag;
  reg        [15:0]   int_reg_array_50_14_real;
  reg        [15:0]   int_reg_array_50_14_imag;
  reg        [15:0]   int_reg_array_50_15_real;
  reg        [15:0]   int_reg_array_50_15_imag;
  reg        [15:0]   int_reg_array_50_16_real;
  reg        [15:0]   int_reg_array_50_16_imag;
  reg        [15:0]   int_reg_array_50_17_real;
  reg        [15:0]   int_reg_array_50_17_imag;
  reg        [15:0]   int_reg_array_50_18_real;
  reg        [15:0]   int_reg_array_50_18_imag;
  reg        [15:0]   int_reg_array_50_19_real;
  reg        [15:0]   int_reg_array_50_19_imag;
  reg        [15:0]   int_reg_array_50_20_real;
  reg        [15:0]   int_reg_array_50_20_imag;
  reg        [15:0]   int_reg_array_50_21_real;
  reg        [15:0]   int_reg_array_50_21_imag;
  reg        [15:0]   int_reg_array_50_22_real;
  reg        [15:0]   int_reg_array_50_22_imag;
  reg        [15:0]   int_reg_array_50_23_real;
  reg        [15:0]   int_reg_array_50_23_imag;
  reg        [15:0]   int_reg_array_50_24_real;
  reg        [15:0]   int_reg_array_50_24_imag;
  reg        [15:0]   int_reg_array_50_25_real;
  reg        [15:0]   int_reg_array_50_25_imag;
  reg        [15:0]   int_reg_array_50_26_real;
  reg        [15:0]   int_reg_array_50_26_imag;
  reg        [15:0]   int_reg_array_50_27_real;
  reg        [15:0]   int_reg_array_50_27_imag;
  reg        [15:0]   int_reg_array_50_28_real;
  reg        [15:0]   int_reg_array_50_28_imag;
  reg        [15:0]   int_reg_array_50_29_real;
  reg        [15:0]   int_reg_array_50_29_imag;
  reg        [15:0]   int_reg_array_50_30_real;
  reg        [15:0]   int_reg_array_50_30_imag;
  reg        [15:0]   int_reg_array_50_31_real;
  reg        [15:0]   int_reg_array_50_31_imag;
  reg        [15:0]   int_reg_array_50_32_real;
  reg        [15:0]   int_reg_array_50_32_imag;
  reg        [15:0]   int_reg_array_50_33_real;
  reg        [15:0]   int_reg_array_50_33_imag;
  reg        [15:0]   int_reg_array_50_34_real;
  reg        [15:0]   int_reg_array_50_34_imag;
  reg        [15:0]   int_reg_array_50_35_real;
  reg        [15:0]   int_reg_array_50_35_imag;
  reg        [15:0]   int_reg_array_50_36_real;
  reg        [15:0]   int_reg_array_50_36_imag;
  reg        [15:0]   int_reg_array_50_37_real;
  reg        [15:0]   int_reg_array_50_37_imag;
  reg        [15:0]   int_reg_array_50_38_real;
  reg        [15:0]   int_reg_array_50_38_imag;
  reg        [15:0]   int_reg_array_50_39_real;
  reg        [15:0]   int_reg_array_50_39_imag;
  reg        [15:0]   int_reg_array_50_40_real;
  reg        [15:0]   int_reg_array_50_40_imag;
  reg        [15:0]   int_reg_array_50_41_real;
  reg        [15:0]   int_reg_array_50_41_imag;
  reg        [15:0]   int_reg_array_50_42_real;
  reg        [15:0]   int_reg_array_50_42_imag;
  reg        [15:0]   int_reg_array_50_43_real;
  reg        [15:0]   int_reg_array_50_43_imag;
  reg        [15:0]   int_reg_array_50_44_real;
  reg        [15:0]   int_reg_array_50_44_imag;
  reg        [15:0]   int_reg_array_50_45_real;
  reg        [15:0]   int_reg_array_50_45_imag;
  reg        [15:0]   int_reg_array_50_46_real;
  reg        [15:0]   int_reg_array_50_46_imag;
  reg        [15:0]   int_reg_array_50_47_real;
  reg        [15:0]   int_reg_array_50_47_imag;
  reg        [15:0]   int_reg_array_50_48_real;
  reg        [15:0]   int_reg_array_50_48_imag;
  reg        [15:0]   int_reg_array_50_49_real;
  reg        [15:0]   int_reg_array_50_49_imag;
  reg        [15:0]   int_reg_array_50_50_real;
  reg        [15:0]   int_reg_array_50_50_imag;
  reg        [15:0]   int_reg_array_50_51_real;
  reg        [15:0]   int_reg_array_50_51_imag;
  reg        [15:0]   int_reg_array_50_52_real;
  reg        [15:0]   int_reg_array_50_52_imag;
  reg        [15:0]   int_reg_array_50_53_real;
  reg        [15:0]   int_reg_array_50_53_imag;
  reg        [15:0]   int_reg_array_50_54_real;
  reg        [15:0]   int_reg_array_50_54_imag;
  reg        [15:0]   int_reg_array_50_55_real;
  reg        [15:0]   int_reg_array_50_55_imag;
  reg        [15:0]   int_reg_array_50_56_real;
  reg        [15:0]   int_reg_array_50_56_imag;
  reg        [15:0]   int_reg_array_50_57_real;
  reg        [15:0]   int_reg_array_50_57_imag;
  reg        [15:0]   int_reg_array_50_58_real;
  reg        [15:0]   int_reg_array_50_58_imag;
  reg        [15:0]   int_reg_array_50_59_real;
  reg        [15:0]   int_reg_array_50_59_imag;
  reg        [15:0]   int_reg_array_50_60_real;
  reg        [15:0]   int_reg_array_50_60_imag;
  reg        [15:0]   int_reg_array_50_61_real;
  reg        [15:0]   int_reg_array_50_61_imag;
  reg        [15:0]   int_reg_array_50_62_real;
  reg        [15:0]   int_reg_array_50_62_imag;
  reg        [15:0]   int_reg_array_50_63_real;
  reg        [15:0]   int_reg_array_50_63_imag;
  reg        [15:0]   int_reg_array_34_0_real;
  reg        [15:0]   int_reg_array_34_0_imag;
  reg        [15:0]   int_reg_array_34_1_real;
  reg        [15:0]   int_reg_array_34_1_imag;
  reg        [15:0]   int_reg_array_34_2_real;
  reg        [15:0]   int_reg_array_34_2_imag;
  reg        [15:0]   int_reg_array_34_3_real;
  reg        [15:0]   int_reg_array_34_3_imag;
  reg        [15:0]   int_reg_array_34_4_real;
  reg        [15:0]   int_reg_array_34_4_imag;
  reg        [15:0]   int_reg_array_34_5_real;
  reg        [15:0]   int_reg_array_34_5_imag;
  reg        [15:0]   int_reg_array_34_6_real;
  reg        [15:0]   int_reg_array_34_6_imag;
  reg        [15:0]   int_reg_array_34_7_real;
  reg        [15:0]   int_reg_array_34_7_imag;
  reg        [15:0]   int_reg_array_34_8_real;
  reg        [15:0]   int_reg_array_34_8_imag;
  reg        [15:0]   int_reg_array_34_9_real;
  reg        [15:0]   int_reg_array_34_9_imag;
  reg        [15:0]   int_reg_array_34_10_real;
  reg        [15:0]   int_reg_array_34_10_imag;
  reg        [15:0]   int_reg_array_34_11_real;
  reg        [15:0]   int_reg_array_34_11_imag;
  reg        [15:0]   int_reg_array_34_12_real;
  reg        [15:0]   int_reg_array_34_12_imag;
  reg        [15:0]   int_reg_array_34_13_real;
  reg        [15:0]   int_reg_array_34_13_imag;
  reg        [15:0]   int_reg_array_34_14_real;
  reg        [15:0]   int_reg_array_34_14_imag;
  reg        [15:0]   int_reg_array_34_15_real;
  reg        [15:0]   int_reg_array_34_15_imag;
  reg        [15:0]   int_reg_array_34_16_real;
  reg        [15:0]   int_reg_array_34_16_imag;
  reg        [15:0]   int_reg_array_34_17_real;
  reg        [15:0]   int_reg_array_34_17_imag;
  reg        [15:0]   int_reg_array_34_18_real;
  reg        [15:0]   int_reg_array_34_18_imag;
  reg        [15:0]   int_reg_array_34_19_real;
  reg        [15:0]   int_reg_array_34_19_imag;
  reg        [15:0]   int_reg_array_34_20_real;
  reg        [15:0]   int_reg_array_34_20_imag;
  reg        [15:0]   int_reg_array_34_21_real;
  reg        [15:0]   int_reg_array_34_21_imag;
  reg        [15:0]   int_reg_array_34_22_real;
  reg        [15:0]   int_reg_array_34_22_imag;
  reg        [15:0]   int_reg_array_34_23_real;
  reg        [15:0]   int_reg_array_34_23_imag;
  reg        [15:0]   int_reg_array_34_24_real;
  reg        [15:0]   int_reg_array_34_24_imag;
  reg        [15:0]   int_reg_array_34_25_real;
  reg        [15:0]   int_reg_array_34_25_imag;
  reg        [15:0]   int_reg_array_34_26_real;
  reg        [15:0]   int_reg_array_34_26_imag;
  reg        [15:0]   int_reg_array_34_27_real;
  reg        [15:0]   int_reg_array_34_27_imag;
  reg        [15:0]   int_reg_array_34_28_real;
  reg        [15:0]   int_reg_array_34_28_imag;
  reg        [15:0]   int_reg_array_34_29_real;
  reg        [15:0]   int_reg_array_34_29_imag;
  reg        [15:0]   int_reg_array_34_30_real;
  reg        [15:0]   int_reg_array_34_30_imag;
  reg        [15:0]   int_reg_array_34_31_real;
  reg        [15:0]   int_reg_array_34_31_imag;
  reg        [15:0]   int_reg_array_34_32_real;
  reg        [15:0]   int_reg_array_34_32_imag;
  reg        [15:0]   int_reg_array_34_33_real;
  reg        [15:0]   int_reg_array_34_33_imag;
  reg        [15:0]   int_reg_array_34_34_real;
  reg        [15:0]   int_reg_array_34_34_imag;
  reg        [15:0]   int_reg_array_34_35_real;
  reg        [15:0]   int_reg_array_34_35_imag;
  reg        [15:0]   int_reg_array_34_36_real;
  reg        [15:0]   int_reg_array_34_36_imag;
  reg        [15:0]   int_reg_array_34_37_real;
  reg        [15:0]   int_reg_array_34_37_imag;
  reg        [15:0]   int_reg_array_34_38_real;
  reg        [15:0]   int_reg_array_34_38_imag;
  reg        [15:0]   int_reg_array_34_39_real;
  reg        [15:0]   int_reg_array_34_39_imag;
  reg        [15:0]   int_reg_array_34_40_real;
  reg        [15:0]   int_reg_array_34_40_imag;
  reg        [15:0]   int_reg_array_34_41_real;
  reg        [15:0]   int_reg_array_34_41_imag;
  reg        [15:0]   int_reg_array_34_42_real;
  reg        [15:0]   int_reg_array_34_42_imag;
  reg        [15:0]   int_reg_array_34_43_real;
  reg        [15:0]   int_reg_array_34_43_imag;
  reg        [15:0]   int_reg_array_34_44_real;
  reg        [15:0]   int_reg_array_34_44_imag;
  reg        [15:0]   int_reg_array_34_45_real;
  reg        [15:0]   int_reg_array_34_45_imag;
  reg        [15:0]   int_reg_array_34_46_real;
  reg        [15:0]   int_reg_array_34_46_imag;
  reg        [15:0]   int_reg_array_34_47_real;
  reg        [15:0]   int_reg_array_34_47_imag;
  reg        [15:0]   int_reg_array_34_48_real;
  reg        [15:0]   int_reg_array_34_48_imag;
  reg        [15:0]   int_reg_array_34_49_real;
  reg        [15:0]   int_reg_array_34_49_imag;
  reg        [15:0]   int_reg_array_34_50_real;
  reg        [15:0]   int_reg_array_34_50_imag;
  reg        [15:0]   int_reg_array_34_51_real;
  reg        [15:0]   int_reg_array_34_51_imag;
  reg        [15:0]   int_reg_array_34_52_real;
  reg        [15:0]   int_reg_array_34_52_imag;
  reg        [15:0]   int_reg_array_34_53_real;
  reg        [15:0]   int_reg_array_34_53_imag;
  reg        [15:0]   int_reg_array_34_54_real;
  reg        [15:0]   int_reg_array_34_54_imag;
  reg        [15:0]   int_reg_array_34_55_real;
  reg        [15:0]   int_reg_array_34_55_imag;
  reg        [15:0]   int_reg_array_34_56_real;
  reg        [15:0]   int_reg_array_34_56_imag;
  reg        [15:0]   int_reg_array_34_57_real;
  reg        [15:0]   int_reg_array_34_57_imag;
  reg        [15:0]   int_reg_array_34_58_real;
  reg        [15:0]   int_reg_array_34_58_imag;
  reg        [15:0]   int_reg_array_34_59_real;
  reg        [15:0]   int_reg_array_34_59_imag;
  reg        [15:0]   int_reg_array_34_60_real;
  reg        [15:0]   int_reg_array_34_60_imag;
  reg        [15:0]   int_reg_array_34_61_real;
  reg        [15:0]   int_reg_array_34_61_imag;
  reg        [15:0]   int_reg_array_34_62_real;
  reg        [15:0]   int_reg_array_34_62_imag;
  reg        [15:0]   int_reg_array_34_63_real;
  reg        [15:0]   int_reg_array_34_63_imag;
  reg        [15:0]   int_reg_array_44_0_real;
  reg        [15:0]   int_reg_array_44_0_imag;
  reg        [15:0]   int_reg_array_44_1_real;
  reg        [15:0]   int_reg_array_44_1_imag;
  reg        [15:0]   int_reg_array_44_2_real;
  reg        [15:0]   int_reg_array_44_2_imag;
  reg        [15:0]   int_reg_array_44_3_real;
  reg        [15:0]   int_reg_array_44_3_imag;
  reg        [15:0]   int_reg_array_44_4_real;
  reg        [15:0]   int_reg_array_44_4_imag;
  reg        [15:0]   int_reg_array_44_5_real;
  reg        [15:0]   int_reg_array_44_5_imag;
  reg        [15:0]   int_reg_array_44_6_real;
  reg        [15:0]   int_reg_array_44_6_imag;
  reg        [15:0]   int_reg_array_44_7_real;
  reg        [15:0]   int_reg_array_44_7_imag;
  reg        [15:0]   int_reg_array_44_8_real;
  reg        [15:0]   int_reg_array_44_8_imag;
  reg        [15:0]   int_reg_array_44_9_real;
  reg        [15:0]   int_reg_array_44_9_imag;
  reg        [15:0]   int_reg_array_44_10_real;
  reg        [15:0]   int_reg_array_44_10_imag;
  reg        [15:0]   int_reg_array_44_11_real;
  reg        [15:0]   int_reg_array_44_11_imag;
  reg        [15:0]   int_reg_array_44_12_real;
  reg        [15:0]   int_reg_array_44_12_imag;
  reg        [15:0]   int_reg_array_44_13_real;
  reg        [15:0]   int_reg_array_44_13_imag;
  reg        [15:0]   int_reg_array_44_14_real;
  reg        [15:0]   int_reg_array_44_14_imag;
  reg        [15:0]   int_reg_array_44_15_real;
  reg        [15:0]   int_reg_array_44_15_imag;
  reg        [15:0]   int_reg_array_44_16_real;
  reg        [15:0]   int_reg_array_44_16_imag;
  reg        [15:0]   int_reg_array_44_17_real;
  reg        [15:0]   int_reg_array_44_17_imag;
  reg        [15:0]   int_reg_array_44_18_real;
  reg        [15:0]   int_reg_array_44_18_imag;
  reg        [15:0]   int_reg_array_44_19_real;
  reg        [15:0]   int_reg_array_44_19_imag;
  reg        [15:0]   int_reg_array_44_20_real;
  reg        [15:0]   int_reg_array_44_20_imag;
  reg        [15:0]   int_reg_array_44_21_real;
  reg        [15:0]   int_reg_array_44_21_imag;
  reg        [15:0]   int_reg_array_44_22_real;
  reg        [15:0]   int_reg_array_44_22_imag;
  reg        [15:0]   int_reg_array_44_23_real;
  reg        [15:0]   int_reg_array_44_23_imag;
  reg        [15:0]   int_reg_array_44_24_real;
  reg        [15:0]   int_reg_array_44_24_imag;
  reg        [15:0]   int_reg_array_44_25_real;
  reg        [15:0]   int_reg_array_44_25_imag;
  reg        [15:0]   int_reg_array_44_26_real;
  reg        [15:0]   int_reg_array_44_26_imag;
  reg        [15:0]   int_reg_array_44_27_real;
  reg        [15:0]   int_reg_array_44_27_imag;
  reg        [15:0]   int_reg_array_44_28_real;
  reg        [15:0]   int_reg_array_44_28_imag;
  reg        [15:0]   int_reg_array_44_29_real;
  reg        [15:0]   int_reg_array_44_29_imag;
  reg        [15:0]   int_reg_array_44_30_real;
  reg        [15:0]   int_reg_array_44_30_imag;
  reg        [15:0]   int_reg_array_44_31_real;
  reg        [15:0]   int_reg_array_44_31_imag;
  reg        [15:0]   int_reg_array_44_32_real;
  reg        [15:0]   int_reg_array_44_32_imag;
  reg        [15:0]   int_reg_array_44_33_real;
  reg        [15:0]   int_reg_array_44_33_imag;
  reg        [15:0]   int_reg_array_44_34_real;
  reg        [15:0]   int_reg_array_44_34_imag;
  reg        [15:0]   int_reg_array_44_35_real;
  reg        [15:0]   int_reg_array_44_35_imag;
  reg        [15:0]   int_reg_array_44_36_real;
  reg        [15:0]   int_reg_array_44_36_imag;
  reg        [15:0]   int_reg_array_44_37_real;
  reg        [15:0]   int_reg_array_44_37_imag;
  reg        [15:0]   int_reg_array_44_38_real;
  reg        [15:0]   int_reg_array_44_38_imag;
  reg        [15:0]   int_reg_array_44_39_real;
  reg        [15:0]   int_reg_array_44_39_imag;
  reg        [15:0]   int_reg_array_44_40_real;
  reg        [15:0]   int_reg_array_44_40_imag;
  reg        [15:0]   int_reg_array_44_41_real;
  reg        [15:0]   int_reg_array_44_41_imag;
  reg        [15:0]   int_reg_array_44_42_real;
  reg        [15:0]   int_reg_array_44_42_imag;
  reg        [15:0]   int_reg_array_44_43_real;
  reg        [15:0]   int_reg_array_44_43_imag;
  reg        [15:0]   int_reg_array_44_44_real;
  reg        [15:0]   int_reg_array_44_44_imag;
  reg        [15:0]   int_reg_array_44_45_real;
  reg        [15:0]   int_reg_array_44_45_imag;
  reg        [15:0]   int_reg_array_44_46_real;
  reg        [15:0]   int_reg_array_44_46_imag;
  reg        [15:0]   int_reg_array_44_47_real;
  reg        [15:0]   int_reg_array_44_47_imag;
  reg        [15:0]   int_reg_array_44_48_real;
  reg        [15:0]   int_reg_array_44_48_imag;
  reg        [15:0]   int_reg_array_44_49_real;
  reg        [15:0]   int_reg_array_44_49_imag;
  reg        [15:0]   int_reg_array_44_50_real;
  reg        [15:0]   int_reg_array_44_50_imag;
  reg        [15:0]   int_reg_array_44_51_real;
  reg        [15:0]   int_reg_array_44_51_imag;
  reg        [15:0]   int_reg_array_44_52_real;
  reg        [15:0]   int_reg_array_44_52_imag;
  reg        [15:0]   int_reg_array_44_53_real;
  reg        [15:0]   int_reg_array_44_53_imag;
  reg        [15:0]   int_reg_array_44_54_real;
  reg        [15:0]   int_reg_array_44_54_imag;
  reg        [15:0]   int_reg_array_44_55_real;
  reg        [15:0]   int_reg_array_44_55_imag;
  reg        [15:0]   int_reg_array_44_56_real;
  reg        [15:0]   int_reg_array_44_56_imag;
  reg        [15:0]   int_reg_array_44_57_real;
  reg        [15:0]   int_reg_array_44_57_imag;
  reg        [15:0]   int_reg_array_44_58_real;
  reg        [15:0]   int_reg_array_44_58_imag;
  reg        [15:0]   int_reg_array_44_59_real;
  reg        [15:0]   int_reg_array_44_59_imag;
  reg        [15:0]   int_reg_array_44_60_real;
  reg        [15:0]   int_reg_array_44_60_imag;
  reg        [15:0]   int_reg_array_44_61_real;
  reg        [15:0]   int_reg_array_44_61_imag;
  reg        [15:0]   int_reg_array_44_62_real;
  reg        [15:0]   int_reg_array_44_62_imag;
  reg        [15:0]   int_reg_array_44_63_real;
  reg        [15:0]   int_reg_array_44_63_imag;
  reg        [15:0]   int_reg_array_22_0_real;
  reg        [15:0]   int_reg_array_22_0_imag;
  reg        [15:0]   int_reg_array_22_1_real;
  reg        [15:0]   int_reg_array_22_1_imag;
  reg        [15:0]   int_reg_array_22_2_real;
  reg        [15:0]   int_reg_array_22_2_imag;
  reg        [15:0]   int_reg_array_22_3_real;
  reg        [15:0]   int_reg_array_22_3_imag;
  reg        [15:0]   int_reg_array_22_4_real;
  reg        [15:0]   int_reg_array_22_4_imag;
  reg        [15:0]   int_reg_array_22_5_real;
  reg        [15:0]   int_reg_array_22_5_imag;
  reg        [15:0]   int_reg_array_22_6_real;
  reg        [15:0]   int_reg_array_22_6_imag;
  reg        [15:0]   int_reg_array_22_7_real;
  reg        [15:0]   int_reg_array_22_7_imag;
  reg        [15:0]   int_reg_array_22_8_real;
  reg        [15:0]   int_reg_array_22_8_imag;
  reg        [15:0]   int_reg_array_22_9_real;
  reg        [15:0]   int_reg_array_22_9_imag;
  reg        [15:0]   int_reg_array_22_10_real;
  reg        [15:0]   int_reg_array_22_10_imag;
  reg        [15:0]   int_reg_array_22_11_real;
  reg        [15:0]   int_reg_array_22_11_imag;
  reg        [15:0]   int_reg_array_22_12_real;
  reg        [15:0]   int_reg_array_22_12_imag;
  reg        [15:0]   int_reg_array_22_13_real;
  reg        [15:0]   int_reg_array_22_13_imag;
  reg        [15:0]   int_reg_array_22_14_real;
  reg        [15:0]   int_reg_array_22_14_imag;
  reg        [15:0]   int_reg_array_22_15_real;
  reg        [15:0]   int_reg_array_22_15_imag;
  reg        [15:0]   int_reg_array_22_16_real;
  reg        [15:0]   int_reg_array_22_16_imag;
  reg        [15:0]   int_reg_array_22_17_real;
  reg        [15:0]   int_reg_array_22_17_imag;
  reg        [15:0]   int_reg_array_22_18_real;
  reg        [15:0]   int_reg_array_22_18_imag;
  reg        [15:0]   int_reg_array_22_19_real;
  reg        [15:0]   int_reg_array_22_19_imag;
  reg        [15:0]   int_reg_array_22_20_real;
  reg        [15:0]   int_reg_array_22_20_imag;
  reg        [15:0]   int_reg_array_22_21_real;
  reg        [15:0]   int_reg_array_22_21_imag;
  reg        [15:0]   int_reg_array_22_22_real;
  reg        [15:0]   int_reg_array_22_22_imag;
  reg        [15:0]   int_reg_array_22_23_real;
  reg        [15:0]   int_reg_array_22_23_imag;
  reg        [15:0]   int_reg_array_22_24_real;
  reg        [15:0]   int_reg_array_22_24_imag;
  reg        [15:0]   int_reg_array_22_25_real;
  reg        [15:0]   int_reg_array_22_25_imag;
  reg        [15:0]   int_reg_array_22_26_real;
  reg        [15:0]   int_reg_array_22_26_imag;
  reg        [15:0]   int_reg_array_22_27_real;
  reg        [15:0]   int_reg_array_22_27_imag;
  reg        [15:0]   int_reg_array_22_28_real;
  reg        [15:0]   int_reg_array_22_28_imag;
  reg        [15:0]   int_reg_array_22_29_real;
  reg        [15:0]   int_reg_array_22_29_imag;
  reg        [15:0]   int_reg_array_22_30_real;
  reg        [15:0]   int_reg_array_22_30_imag;
  reg        [15:0]   int_reg_array_22_31_real;
  reg        [15:0]   int_reg_array_22_31_imag;
  reg        [15:0]   int_reg_array_22_32_real;
  reg        [15:0]   int_reg_array_22_32_imag;
  reg        [15:0]   int_reg_array_22_33_real;
  reg        [15:0]   int_reg_array_22_33_imag;
  reg        [15:0]   int_reg_array_22_34_real;
  reg        [15:0]   int_reg_array_22_34_imag;
  reg        [15:0]   int_reg_array_22_35_real;
  reg        [15:0]   int_reg_array_22_35_imag;
  reg        [15:0]   int_reg_array_22_36_real;
  reg        [15:0]   int_reg_array_22_36_imag;
  reg        [15:0]   int_reg_array_22_37_real;
  reg        [15:0]   int_reg_array_22_37_imag;
  reg        [15:0]   int_reg_array_22_38_real;
  reg        [15:0]   int_reg_array_22_38_imag;
  reg        [15:0]   int_reg_array_22_39_real;
  reg        [15:0]   int_reg_array_22_39_imag;
  reg        [15:0]   int_reg_array_22_40_real;
  reg        [15:0]   int_reg_array_22_40_imag;
  reg        [15:0]   int_reg_array_22_41_real;
  reg        [15:0]   int_reg_array_22_41_imag;
  reg        [15:0]   int_reg_array_22_42_real;
  reg        [15:0]   int_reg_array_22_42_imag;
  reg        [15:0]   int_reg_array_22_43_real;
  reg        [15:0]   int_reg_array_22_43_imag;
  reg        [15:0]   int_reg_array_22_44_real;
  reg        [15:0]   int_reg_array_22_44_imag;
  reg        [15:0]   int_reg_array_22_45_real;
  reg        [15:0]   int_reg_array_22_45_imag;
  reg        [15:0]   int_reg_array_22_46_real;
  reg        [15:0]   int_reg_array_22_46_imag;
  reg        [15:0]   int_reg_array_22_47_real;
  reg        [15:0]   int_reg_array_22_47_imag;
  reg        [15:0]   int_reg_array_22_48_real;
  reg        [15:0]   int_reg_array_22_48_imag;
  reg        [15:0]   int_reg_array_22_49_real;
  reg        [15:0]   int_reg_array_22_49_imag;
  reg        [15:0]   int_reg_array_22_50_real;
  reg        [15:0]   int_reg_array_22_50_imag;
  reg        [15:0]   int_reg_array_22_51_real;
  reg        [15:0]   int_reg_array_22_51_imag;
  reg        [15:0]   int_reg_array_22_52_real;
  reg        [15:0]   int_reg_array_22_52_imag;
  reg        [15:0]   int_reg_array_22_53_real;
  reg        [15:0]   int_reg_array_22_53_imag;
  reg        [15:0]   int_reg_array_22_54_real;
  reg        [15:0]   int_reg_array_22_54_imag;
  reg        [15:0]   int_reg_array_22_55_real;
  reg        [15:0]   int_reg_array_22_55_imag;
  reg        [15:0]   int_reg_array_22_56_real;
  reg        [15:0]   int_reg_array_22_56_imag;
  reg        [15:0]   int_reg_array_22_57_real;
  reg        [15:0]   int_reg_array_22_57_imag;
  reg        [15:0]   int_reg_array_22_58_real;
  reg        [15:0]   int_reg_array_22_58_imag;
  reg        [15:0]   int_reg_array_22_59_real;
  reg        [15:0]   int_reg_array_22_59_imag;
  reg        [15:0]   int_reg_array_22_60_real;
  reg        [15:0]   int_reg_array_22_60_imag;
  reg        [15:0]   int_reg_array_22_61_real;
  reg        [15:0]   int_reg_array_22_61_imag;
  reg        [15:0]   int_reg_array_22_62_real;
  reg        [15:0]   int_reg_array_22_62_imag;
  reg        [15:0]   int_reg_array_22_63_real;
  reg        [15:0]   int_reg_array_22_63_imag;
  reg        [15:0]   int_reg_array_43_0_real;
  reg        [15:0]   int_reg_array_43_0_imag;
  reg        [15:0]   int_reg_array_43_1_real;
  reg        [15:0]   int_reg_array_43_1_imag;
  reg        [15:0]   int_reg_array_43_2_real;
  reg        [15:0]   int_reg_array_43_2_imag;
  reg        [15:0]   int_reg_array_43_3_real;
  reg        [15:0]   int_reg_array_43_3_imag;
  reg        [15:0]   int_reg_array_43_4_real;
  reg        [15:0]   int_reg_array_43_4_imag;
  reg        [15:0]   int_reg_array_43_5_real;
  reg        [15:0]   int_reg_array_43_5_imag;
  reg        [15:0]   int_reg_array_43_6_real;
  reg        [15:0]   int_reg_array_43_6_imag;
  reg        [15:0]   int_reg_array_43_7_real;
  reg        [15:0]   int_reg_array_43_7_imag;
  reg        [15:0]   int_reg_array_43_8_real;
  reg        [15:0]   int_reg_array_43_8_imag;
  reg        [15:0]   int_reg_array_43_9_real;
  reg        [15:0]   int_reg_array_43_9_imag;
  reg        [15:0]   int_reg_array_43_10_real;
  reg        [15:0]   int_reg_array_43_10_imag;
  reg        [15:0]   int_reg_array_43_11_real;
  reg        [15:0]   int_reg_array_43_11_imag;
  reg        [15:0]   int_reg_array_43_12_real;
  reg        [15:0]   int_reg_array_43_12_imag;
  reg        [15:0]   int_reg_array_43_13_real;
  reg        [15:0]   int_reg_array_43_13_imag;
  reg        [15:0]   int_reg_array_43_14_real;
  reg        [15:0]   int_reg_array_43_14_imag;
  reg        [15:0]   int_reg_array_43_15_real;
  reg        [15:0]   int_reg_array_43_15_imag;
  reg        [15:0]   int_reg_array_43_16_real;
  reg        [15:0]   int_reg_array_43_16_imag;
  reg        [15:0]   int_reg_array_43_17_real;
  reg        [15:0]   int_reg_array_43_17_imag;
  reg        [15:0]   int_reg_array_43_18_real;
  reg        [15:0]   int_reg_array_43_18_imag;
  reg        [15:0]   int_reg_array_43_19_real;
  reg        [15:0]   int_reg_array_43_19_imag;
  reg        [15:0]   int_reg_array_43_20_real;
  reg        [15:0]   int_reg_array_43_20_imag;
  reg        [15:0]   int_reg_array_43_21_real;
  reg        [15:0]   int_reg_array_43_21_imag;
  reg        [15:0]   int_reg_array_43_22_real;
  reg        [15:0]   int_reg_array_43_22_imag;
  reg        [15:0]   int_reg_array_43_23_real;
  reg        [15:0]   int_reg_array_43_23_imag;
  reg        [15:0]   int_reg_array_43_24_real;
  reg        [15:0]   int_reg_array_43_24_imag;
  reg        [15:0]   int_reg_array_43_25_real;
  reg        [15:0]   int_reg_array_43_25_imag;
  reg        [15:0]   int_reg_array_43_26_real;
  reg        [15:0]   int_reg_array_43_26_imag;
  reg        [15:0]   int_reg_array_43_27_real;
  reg        [15:0]   int_reg_array_43_27_imag;
  reg        [15:0]   int_reg_array_43_28_real;
  reg        [15:0]   int_reg_array_43_28_imag;
  reg        [15:0]   int_reg_array_43_29_real;
  reg        [15:0]   int_reg_array_43_29_imag;
  reg        [15:0]   int_reg_array_43_30_real;
  reg        [15:0]   int_reg_array_43_30_imag;
  reg        [15:0]   int_reg_array_43_31_real;
  reg        [15:0]   int_reg_array_43_31_imag;
  reg        [15:0]   int_reg_array_43_32_real;
  reg        [15:0]   int_reg_array_43_32_imag;
  reg        [15:0]   int_reg_array_43_33_real;
  reg        [15:0]   int_reg_array_43_33_imag;
  reg        [15:0]   int_reg_array_43_34_real;
  reg        [15:0]   int_reg_array_43_34_imag;
  reg        [15:0]   int_reg_array_43_35_real;
  reg        [15:0]   int_reg_array_43_35_imag;
  reg        [15:0]   int_reg_array_43_36_real;
  reg        [15:0]   int_reg_array_43_36_imag;
  reg        [15:0]   int_reg_array_43_37_real;
  reg        [15:0]   int_reg_array_43_37_imag;
  reg        [15:0]   int_reg_array_43_38_real;
  reg        [15:0]   int_reg_array_43_38_imag;
  reg        [15:0]   int_reg_array_43_39_real;
  reg        [15:0]   int_reg_array_43_39_imag;
  reg        [15:0]   int_reg_array_43_40_real;
  reg        [15:0]   int_reg_array_43_40_imag;
  reg        [15:0]   int_reg_array_43_41_real;
  reg        [15:0]   int_reg_array_43_41_imag;
  reg        [15:0]   int_reg_array_43_42_real;
  reg        [15:0]   int_reg_array_43_42_imag;
  reg        [15:0]   int_reg_array_43_43_real;
  reg        [15:0]   int_reg_array_43_43_imag;
  reg        [15:0]   int_reg_array_43_44_real;
  reg        [15:0]   int_reg_array_43_44_imag;
  reg        [15:0]   int_reg_array_43_45_real;
  reg        [15:0]   int_reg_array_43_45_imag;
  reg        [15:0]   int_reg_array_43_46_real;
  reg        [15:0]   int_reg_array_43_46_imag;
  reg        [15:0]   int_reg_array_43_47_real;
  reg        [15:0]   int_reg_array_43_47_imag;
  reg        [15:0]   int_reg_array_43_48_real;
  reg        [15:0]   int_reg_array_43_48_imag;
  reg        [15:0]   int_reg_array_43_49_real;
  reg        [15:0]   int_reg_array_43_49_imag;
  reg        [15:0]   int_reg_array_43_50_real;
  reg        [15:0]   int_reg_array_43_50_imag;
  reg        [15:0]   int_reg_array_43_51_real;
  reg        [15:0]   int_reg_array_43_51_imag;
  reg        [15:0]   int_reg_array_43_52_real;
  reg        [15:0]   int_reg_array_43_52_imag;
  reg        [15:0]   int_reg_array_43_53_real;
  reg        [15:0]   int_reg_array_43_53_imag;
  reg        [15:0]   int_reg_array_43_54_real;
  reg        [15:0]   int_reg_array_43_54_imag;
  reg        [15:0]   int_reg_array_43_55_real;
  reg        [15:0]   int_reg_array_43_55_imag;
  reg        [15:0]   int_reg_array_43_56_real;
  reg        [15:0]   int_reg_array_43_56_imag;
  reg        [15:0]   int_reg_array_43_57_real;
  reg        [15:0]   int_reg_array_43_57_imag;
  reg        [15:0]   int_reg_array_43_58_real;
  reg        [15:0]   int_reg_array_43_58_imag;
  reg        [15:0]   int_reg_array_43_59_real;
  reg        [15:0]   int_reg_array_43_59_imag;
  reg        [15:0]   int_reg_array_43_60_real;
  reg        [15:0]   int_reg_array_43_60_imag;
  reg        [15:0]   int_reg_array_43_61_real;
  reg        [15:0]   int_reg_array_43_61_imag;
  reg        [15:0]   int_reg_array_43_62_real;
  reg        [15:0]   int_reg_array_43_62_imag;
  reg        [15:0]   int_reg_array_43_63_real;
  reg        [15:0]   int_reg_array_43_63_imag;
  reg        [15:0]   int_reg_array_30_0_real;
  reg        [15:0]   int_reg_array_30_0_imag;
  reg        [15:0]   int_reg_array_30_1_real;
  reg        [15:0]   int_reg_array_30_1_imag;
  reg        [15:0]   int_reg_array_30_2_real;
  reg        [15:0]   int_reg_array_30_2_imag;
  reg        [15:0]   int_reg_array_30_3_real;
  reg        [15:0]   int_reg_array_30_3_imag;
  reg        [15:0]   int_reg_array_30_4_real;
  reg        [15:0]   int_reg_array_30_4_imag;
  reg        [15:0]   int_reg_array_30_5_real;
  reg        [15:0]   int_reg_array_30_5_imag;
  reg        [15:0]   int_reg_array_30_6_real;
  reg        [15:0]   int_reg_array_30_6_imag;
  reg        [15:0]   int_reg_array_30_7_real;
  reg        [15:0]   int_reg_array_30_7_imag;
  reg        [15:0]   int_reg_array_30_8_real;
  reg        [15:0]   int_reg_array_30_8_imag;
  reg        [15:0]   int_reg_array_30_9_real;
  reg        [15:0]   int_reg_array_30_9_imag;
  reg        [15:0]   int_reg_array_30_10_real;
  reg        [15:0]   int_reg_array_30_10_imag;
  reg        [15:0]   int_reg_array_30_11_real;
  reg        [15:0]   int_reg_array_30_11_imag;
  reg        [15:0]   int_reg_array_30_12_real;
  reg        [15:0]   int_reg_array_30_12_imag;
  reg        [15:0]   int_reg_array_30_13_real;
  reg        [15:0]   int_reg_array_30_13_imag;
  reg        [15:0]   int_reg_array_30_14_real;
  reg        [15:0]   int_reg_array_30_14_imag;
  reg        [15:0]   int_reg_array_30_15_real;
  reg        [15:0]   int_reg_array_30_15_imag;
  reg        [15:0]   int_reg_array_30_16_real;
  reg        [15:0]   int_reg_array_30_16_imag;
  reg        [15:0]   int_reg_array_30_17_real;
  reg        [15:0]   int_reg_array_30_17_imag;
  reg        [15:0]   int_reg_array_30_18_real;
  reg        [15:0]   int_reg_array_30_18_imag;
  reg        [15:0]   int_reg_array_30_19_real;
  reg        [15:0]   int_reg_array_30_19_imag;
  reg        [15:0]   int_reg_array_30_20_real;
  reg        [15:0]   int_reg_array_30_20_imag;
  reg        [15:0]   int_reg_array_30_21_real;
  reg        [15:0]   int_reg_array_30_21_imag;
  reg        [15:0]   int_reg_array_30_22_real;
  reg        [15:0]   int_reg_array_30_22_imag;
  reg        [15:0]   int_reg_array_30_23_real;
  reg        [15:0]   int_reg_array_30_23_imag;
  reg        [15:0]   int_reg_array_30_24_real;
  reg        [15:0]   int_reg_array_30_24_imag;
  reg        [15:0]   int_reg_array_30_25_real;
  reg        [15:0]   int_reg_array_30_25_imag;
  reg        [15:0]   int_reg_array_30_26_real;
  reg        [15:0]   int_reg_array_30_26_imag;
  reg        [15:0]   int_reg_array_30_27_real;
  reg        [15:0]   int_reg_array_30_27_imag;
  reg        [15:0]   int_reg_array_30_28_real;
  reg        [15:0]   int_reg_array_30_28_imag;
  reg        [15:0]   int_reg_array_30_29_real;
  reg        [15:0]   int_reg_array_30_29_imag;
  reg        [15:0]   int_reg_array_30_30_real;
  reg        [15:0]   int_reg_array_30_30_imag;
  reg        [15:0]   int_reg_array_30_31_real;
  reg        [15:0]   int_reg_array_30_31_imag;
  reg        [15:0]   int_reg_array_30_32_real;
  reg        [15:0]   int_reg_array_30_32_imag;
  reg        [15:0]   int_reg_array_30_33_real;
  reg        [15:0]   int_reg_array_30_33_imag;
  reg        [15:0]   int_reg_array_30_34_real;
  reg        [15:0]   int_reg_array_30_34_imag;
  reg        [15:0]   int_reg_array_30_35_real;
  reg        [15:0]   int_reg_array_30_35_imag;
  reg        [15:0]   int_reg_array_30_36_real;
  reg        [15:0]   int_reg_array_30_36_imag;
  reg        [15:0]   int_reg_array_30_37_real;
  reg        [15:0]   int_reg_array_30_37_imag;
  reg        [15:0]   int_reg_array_30_38_real;
  reg        [15:0]   int_reg_array_30_38_imag;
  reg        [15:0]   int_reg_array_30_39_real;
  reg        [15:0]   int_reg_array_30_39_imag;
  reg        [15:0]   int_reg_array_30_40_real;
  reg        [15:0]   int_reg_array_30_40_imag;
  reg        [15:0]   int_reg_array_30_41_real;
  reg        [15:0]   int_reg_array_30_41_imag;
  reg        [15:0]   int_reg_array_30_42_real;
  reg        [15:0]   int_reg_array_30_42_imag;
  reg        [15:0]   int_reg_array_30_43_real;
  reg        [15:0]   int_reg_array_30_43_imag;
  reg        [15:0]   int_reg_array_30_44_real;
  reg        [15:0]   int_reg_array_30_44_imag;
  reg        [15:0]   int_reg_array_30_45_real;
  reg        [15:0]   int_reg_array_30_45_imag;
  reg        [15:0]   int_reg_array_30_46_real;
  reg        [15:0]   int_reg_array_30_46_imag;
  reg        [15:0]   int_reg_array_30_47_real;
  reg        [15:0]   int_reg_array_30_47_imag;
  reg        [15:0]   int_reg_array_30_48_real;
  reg        [15:0]   int_reg_array_30_48_imag;
  reg        [15:0]   int_reg_array_30_49_real;
  reg        [15:0]   int_reg_array_30_49_imag;
  reg        [15:0]   int_reg_array_30_50_real;
  reg        [15:0]   int_reg_array_30_50_imag;
  reg        [15:0]   int_reg_array_30_51_real;
  reg        [15:0]   int_reg_array_30_51_imag;
  reg        [15:0]   int_reg_array_30_52_real;
  reg        [15:0]   int_reg_array_30_52_imag;
  reg        [15:0]   int_reg_array_30_53_real;
  reg        [15:0]   int_reg_array_30_53_imag;
  reg        [15:0]   int_reg_array_30_54_real;
  reg        [15:0]   int_reg_array_30_54_imag;
  reg        [15:0]   int_reg_array_30_55_real;
  reg        [15:0]   int_reg_array_30_55_imag;
  reg        [15:0]   int_reg_array_30_56_real;
  reg        [15:0]   int_reg_array_30_56_imag;
  reg        [15:0]   int_reg_array_30_57_real;
  reg        [15:0]   int_reg_array_30_57_imag;
  reg        [15:0]   int_reg_array_30_58_real;
  reg        [15:0]   int_reg_array_30_58_imag;
  reg        [15:0]   int_reg_array_30_59_real;
  reg        [15:0]   int_reg_array_30_59_imag;
  reg        [15:0]   int_reg_array_30_60_real;
  reg        [15:0]   int_reg_array_30_60_imag;
  reg        [15:0]   int_reg_array_30_61_real;
  reg        [15:0]   int_reg_array_30_61_imag;
  reg        [15:0]   int_reg_array_30_62_real;
  reg        [15:0]   int_reg_array_30_62_imag;
  reg        [15:0]   int_reg_array_30_63_real;
  reg        [15:0]   int_reg_array_30_63_imag;
  reg        [15:0]   int_reg_array_31_0_real;
  reg        [15:0]   int_reg_array_31_0_imag;
  reg        [15:0]   int_reg_array_31_1_real;
  reg        [15:0]   int_reg_array_31_1_imag;
  reg        [15:0]   int_reg_array_31_2_real;
  reg        [15:0]   int_reg_array_31_2_imag;
  reg        [15:0]   int_reg_array_31_3_real;
  reg        [15:0]   int_reg_array_31_3_imag;
  reg        [15:0]   int_reg_array_31_4_real;
  reg        [15:0]   int_reg_array_31_4_imag;
  reg        [15:0]   int_reg_array_31_5_real;
  reg        [15:0]   int_reg_array_31_5_imag;
  reg        [15:0]   int_reg_array_31_6_real;
  reg        [15:0]   int_reg_array_31_6_imag;
  reg        [15:0]   int_reg_array_31_7_real;
  reg        [15:0]   int_reg_array_31_7_imag;
  reg        [15:0]   int_reg_array_31_8_real;
  reg        [15:0]   int_reg_array_31_8_imag;
  reg        [15:0]   int_reg_array_31_9_real;
  reg        [15:0]   int_reg_array_31_9_imag;
  reg        [15:0]   int_reg_array_31_10_real;
  reg        [15:0]   int_reg_array_31_10_imag;
  reg        [15:0]   int_reg_array_31_11_real;
  reg        [15:0]   int_reg_array_31_11_imag;
  reg        [15:0]   int_reg_array_31_12_real;
  reg        [15:0]   int_reg_array_31_12_imag;
  reg        [15:0]   int_reg_array_31_13_real;
  reg        [15:0]   int_reg_array_31_13_imag;
  reg        [15:0]   int_reg_array_31_14_real;
  reg        [15:0]   int_reg_array_31_14_imag;
  reg        [15:0]   int_reg_array_31_15_real;
  reg        [15:0]   int_reg_array_31_15_imag;
  reg        [15:0]   int_reg_array_31_16_real;
  reg        [15:0]   int_reg_array_31_16_imag;
  reg        [15:0]   int_reg_array_31_17_real;
  reg        [15:0]   int_reg_array_31_17_imag;
  reg        [15:0]   int_reg_array_31_18_real;
  reg        [15:0]   int_reg_array_31_18_imag;
  reg        [15:0]   int_reg_array_31_19_real;
  reg        [15:0]   int_reg_array_31_19_imag;
  reg        [15:0]   int_reg_array_31_20_real;
  reg        [15:0]   int_reg_array_31_20_imag;
  reg        [15:0]   int_reg_array_31_21_real;
  reg        [15:0]   int_reg_array_31_21_imag;
  reg        [15:0]   int_reg_array_31_22_real;
  reg        [15:0]   int_reg_array_31_22_imag;
  reg        [15:0]   int_reg_array_31_23_real;
  reg        [15:0]   int_reg_array_31_23_imag;
  reg        [15:0]   int_reg_array_31_24_real;
  reg        [15:0]   int_reg_array_31_24_imag;
  reg        [15:0]   int_reg_array_31_25_real;
  reg        [15:0]   int_reg_array_31_25_imag;
  reg        [15:0]   int_reg_array_31_26_real;
  reg        [15:0]   int_reg_array_31_26_imag;
  reg        [15:0]   int_reg_array_31_27_real;
  reg        [15:0]   int_reg_array_31_27_imag;
  reg        [15:0]   int_reg_array_31_28_real;
  reg        [15:0]   int_reg_array_31_28_imag;
  reg        [15:0]   int_reg_array_31_29_real;
  reg        [15:0]   int_reg_array_31_29_imag;
  reg        [15:0]   int_reg_array_31_30_real;
  reg        [15:0]   int_reg_array_31_30_imag;
  reg        [15:0]   int_reg_array_31_31_real;
  reg        [15:0]   int_reg_array_31_31_imag;
  reg        [15:0]   int_reg_array_31_32_real;
  reg        [15:0]   int_reg_array_31_32_imag;
  reg        [15:0]   int_reg_array_31_33_real;
  reg        [15:0]   int_reg_array_31_33_imag;
  reg        [15:0]   int_reg_array_31_34_real;
  reg        [15:0]   int_reg_array_31_34_imag;
  reg        [15:0]   int_reg_array_31_35_real;
  reg        [15:0]   int_reg_array_31_35_imag;
  reg        [15:0]   int_reg_array_31_36_real;
  reg        [15:0]   int_reg_array_31_36_imag;
  reg        [15:0]   int_reg_array_31_37_real;
  reg        [15:0]   int_reg_array_31_37_imag;
  reg        [15:0]   int_reg_array_31_38_real;
  reg        [15:0]   int_reg_array_31_38_imag;
  reg        [15:0]   int_reg_array_31_39_real;
  reg        [15:0]   int_reg_array_31_39_imag;
  reg        [15:0]   int_reg_array_31_40_real;
  reg        [15:0]   int_reg_array_31_40_imag;
  reg        [15:0]   int_reg_array_31_41_real;
  reg        [15:0]   int_reg_array_31_41_imag;
  reg        [15:0]   int_reg_array_31_42_real;
  reg        [15:0]   int_reg_array_31_42_imag;
  reg        [15:0]   int_reg_array_31_43_real;
  reg        [15:0]   int_reg_array_31_43_imag;
  reg        [15:0]   int_reg_array_31_44_real;
  reg        [15:0]   int_reg_array_31_44_imag;
  reg        [15:0]   int_reg_array_31_45_real;
  reg        [15:0]   int_reg_array_31_45_imag;
  reg        [15:0]   int_reg_array_31_46_real;
  reg        [15:0]   int_reg_array_31_46_imag;
  reg        [15:0]   int_reg_array_31_47_real;
  reg        [15:0]   int_reg_array_31_47_imag;
  reg        [15:0]   int_reg_array_31_48_real;
  reg        [15:0]   int_reg_array_31_48_imag;
  reg        [15:0]   int_reg_array_31_49_real;
  reg        [15:0]   int_reg_array_31_49_imag;
  reg        [15:0]   int_reg_array_31_50_real;
  reg        [15:0]   int_reg_array_31_50_imag;
  reg        [15:0]   int_reg_array_31_51_real;
  reg        [15:0]   int_reg_array_31_51_imag;
  reg        [15:0]   int_reg_array_31_52_real;
  reg        [15:0]   int_reg_array_31_52_imag;
  reg        [15:0]   int_reg_array_31_53_real;
  reg        [15:0]   int_reg_array_31_53_imag;
  reg        [15:0]   int_reg_array_31_54_real;
  reg        [15:0]   int_reg_array_31_54_imag;
  reg        [15:0]   int_reg_array_31_55_real;
  reg        [15:0]   int_reg_array_31_55_imag;
  reg        [15:0]   int_reg_array_31_56_real;
  reg        [15:0]   int_reg_array_31_56_imag;
  reg        [15:0]   int_reg_array_31_57_real;
  reg        [15:0]   int_reg_array_31_57_imag;
  reg        [15:0]   int_reg_array_31_58_real;
  reg        [15:0]   int_reg_array_31_58_imag;
  reg        [15:0]   int_reg_array_31_59_real;
  reg        [15:0]   int_reg_array_31_59_imag;
  reg        [15:0]   int_reg_array_31_60_real;
  reg        [15:0]   int_reg_array_31_60_imag;
  reg        [15:0]   int_reg_array_31_61_real;
  reg        [15:0]   int_reg_array_31_61_imag;
  reg        [15:0]   int_reg_array_31_62_real;
  reg        [15:0]   int_reg_array_31_62_imag;
  reg        [15:0]   int_reg_array_31_63_real;
  reg        [15:0]   int_reg_array_31_63_imag;
  reg        [15:0]   int_reg_array_20_0_real;
  reg        [15:0]   int_reg_array_20_0_imag;
  reg        [15:0]   int_reg_array_20_1_real;
  reg        [15:0]   int_reg_array_20_1_imag;
  reg        [15:0]   int_reg_array_20_2_real;
  reg        [15:0]   int_reg_array_20_2_imag;
  reg        [15:0]   int_reg_array_20_3_real;
  reg        [15:0]   int_reg_array_20_3_imag;
  reg        [15:0]   int_reg_array_20_4_real;
  reg        [15:0]   int_reg_array_20_4_imag;
  reg        [15:0]   int_reg_array_20_5_real;
  reg        [15:0]   int_reg_array_20_5_imag;
  reg        [15:0]   int_reg_array_20_6_real;
  reg        [15:0]   int_reg_array_20_6_imag;
  reg        [15:0]   int_reg_array_20_7_real;
  reg        [15:0]   int_reg_array_20_7_imag;
  reg        [15:0]   int_reg_array_20_8_real;
  reg        [15:0]   int_reg_array_20_8_imag;
  reg        [15:0]   int_reg_array_20_9_real;
  reg        [15:0]   int_reg_array_20_9_imag;
  reg        [15:0]   int_reg_array_20_10_real;
  reg        [15:0]   int_reg_array_20_10_imag;
  reg        [15:0]   int_reg_array_20_11_real;
  reg        [15:0]   int_reg_array_20_11_imag;
  reg        [15:0]   int_reg_array_20_12_real;
  reg        [15:0]   int_reg_array_20_12_imag;
  reg        [15:0]   int_reg_array_20_13_real;
  reg        [15:0]   int_reg_array_20_13_imag;
  reg        [15:0]   int_reg_array_20_14_real;
  reg        [15:0]   int_reg_array_20_14_imag;
  reg        [15:0]   int_reg_array_20_15_real;
  reg        [15:0]   int_reg_array_20_15_imag;
  reg        [15:0]   int_reg_array_20_16_real;
  reg        [15:0]   int_reg_array_20_16_imag;
  reg        [15:0]   int_reg_array_20_17_real;
  reg        [15:0]   int_reg_array_20_17_imag;
  reg        [15:0]   int_reg_array_20_18_real;
  reg        [15:0]   int_reg_array_20_18_imag;
  reg        [15:0]   int_reg_array_20_19_real;
  reg        [15:0]   int_reg_array_20_19_imag;
  reg        [15:0]   int_reg_array_20_20_real;
  reg        [15:0]   int_reg_array_20_20_imag;
  reg        [15:0]   int_reg_array_20_21_real;
  reg        [15:0]   int_reg_array_20_21_imag;
  reg        [15:0]   int_reg_array_20_22_real;
  reg        [15:0]   int_reg_array_20_22_imag;
  reg        [15:0]   int_reg_array_20_23_real;
  reg        [15:0]   int_reg_array_20_23_imag;
  reg        [15:0]   int_reg_array_20_24_real;
  reg        [15:0]   int_reg_array_20_24_imag;
  reg        [15:0]   int_reg_array_20_25_real;
  reg        [15:0]   int_reg_array_20_25_imag;
  reg        [15:0]   int_reg_array_20_26_real;
  reg        [15:0]   int_reg_array_20_26_imag;
  reg        [15:0]   int_reg_array_20_27_real;
  reg        [15:0]   int_reg_array_20_27_imag;
  reg        [15:0]   int_reg_array_20_28_real;
  reg        [15:0]   int_reg_array_20_28_imag;
  reg        [15:0]   int_reg_array_20_29_real;
  reg        [15:0]   int_reg_array_20_29_imag;
  reg        [15:0]   int_reg_array_20_30_real;
  reg        [15:0]   int_reg_array_20_30_imag;
  reg        [15:0]   int_reg_array_20_31_real;
  reg        [15:0]   int_reg_array_20_31_imag;
  reg        [15:0]   int_reg_array_20_32_real;
  reg        [15:0]   int_reg_array_20_32_imag;
  reg        [15:0]   int_reg_array_20_33_real;
  reg        [15:0]   int_reg_array_20_33_imag;
  reg        [15:0]   int_reg_array_20_34_real;
  reg        [15:0]   int_reg_array_20_34_imag;
  reg        [15:0]   int_reg_array_20_35_real;
  reg        [15:0]   int_reg_array_20_35_imag;
  reg        [15:0]   int_reg_array_20_36_real;
  reg        [15:0]   int_reg_array_20_36_imag;
  reg        [15:0]   int_reg_array_20_37_real;
  reg        [15:0]   int_reg_array_20_37_imag;
  reg        [15:0]   int_reg_array_20_38_real;
  reg        [15:0]   int_reg_array_20_38_imag;
  reg        [15:0]   int_reg_array_20_39_real;
  reg        [15:0]   int_reg_array_20_39_imag;
  reg        [15:0]   int_reg_array_20_40_real;
  reg        [15:0]   int_reg_array_20_40_imag;
  reg        [15:0]   int_reg_array_20_41_real;
  reg        [15:0]   int_reg_array_20_41_imag;
  reg        [15:0]   int_reg_array_20_42_real;
  reg        [15:0]   int_reg_array_20_42_imag;
  reg        [15:0]   int_reg_array_20_43_real;
  reg        [15:0]   int_reg_array_20_43_imag;
  reg        [15:0]   int_reg_array_20_44_real;
  reg        [15:0]   int_reg_array_20_44_imag;
  reg        [15:0]   int_reg_array_20_45_real;
  reg        [15:0]   int_reg_array_20_45_imag;
  reg        [15:0]   int_reg_array_20_46_real;
  reg        [15:0]   int_reg_array_20_46_imag;
  reg        [15:0]   int_reg_array_20_47_real;
  reg        [15:0]   int_reg_array_20_47_imag;
  reg        [15:0]   int_reg_array_20_48_real;
  reg        [15:0]   int_reg_array_20_48_imag;
  reg        [15:0]   int_reg_array_20_49_real;
  reg        [15:0]   int_reg_array_20_49_imag;
  reg        [15:0]   int_reg_array_20_50_real;
  reg        [15:0]   int_reg_array_20_50_imag;
  reg        [15:0]   int_reg_array_20_51_real;
  reg        [15:0]   int_reg_array_20_51_imag;
  reg        [15:0]   int_reg_array_20_52_real;
  reg        [15:0]   int_reg_array_20_52_imag;
  reg        [15:0]   int_reg_array_20_53_real;
  reg        [15:0]   int_reg_array_20_53_imag;
  reg        [15:0]   int_reg_array_20_54_real;
  reg        [15:0]   int_reg_array_20_54_imag;
  reg        [15:0]   int_reg_array_20_55_real;
  reg        [15:0]   int_reg_array_20_55_imag;
  reg        [15:0]   int_reg_array_20_56_real;
  reg        [15:0]   int_reg_array_20_56_imag;
  reg        [15:0]   int_reg_array_20_57_real;
  reg        [15:0]   int_reg_array_20_57_imag;
  reg        [15:0]   int_reg_array_20_58_real;
  reg        [15:0]   int_reg_array_20_58_imag;
  reg        [15:0]   int_reg_array_20_59_real;
  reg        [15:0]   int_reg_array_20_59_imag;
  reg        [15:0]   int_reg_array_20_60_real;
  reg        [15:0]   int_reg_array_20_60_imag;
  reg        [15:0]   int_reg_array_20_61_real;
  reg        [15:0]   int_reg_array_20_61_imag;
  reg        [15:0]   int_reg_array_20_62_real;
  reg        [15:0]   int_reg_array_20_62_imag;
  reg        [15:0]   int_reg_array_20_63_real;
  reg        [15:0]   int_reg_array_20_63_imag;
  reg        [15:0]   int_reg_array_47_0_real;
  reg        [15:0]   int_reg_array_47_0_imag;
  reg        [15:0]   int_reg_array_47_1_real;
  reg        [15:0]   int_reg_array_47_1_imag;
  reg        [15:0]   int_reg_array_47_2_real;
  reg        [15:0]   int_reg_array_47_2_imag;
  reg        [15:0]   int_reg_array_47_3_real;
  reg        [15:0]   int_reg_array_47_3_imag;
  reg        [15:0]   int_reg_array_47_4_real;
  reg        [15:0]   int_reg_array_47_4_imag;
  reg        [15:0]   int_reg_array_47_5_real;
  reg        [15:0]   int_reg_array_47_5_imag;
  reg        [15:0]   int_reg_array_47_6_real;
  reg        [15:0]   int_reg_array_47_6_imag;
  reg        [15:0]   int_reg_array_47_7_real;
  reg        [15:0]   int_reg_array_47_7_imag;
  reg        [15:0]   int_reg_array_47_8_real;
  reg        [15:0]   int_reg_array_47_8_imag;
  reg        [15:0]   int_reg_array_47_9_real;
  reg        [15:0]   int_reg_array_47_9_imag;
  reg        [15:0]   int_reg_array_47_10_real;
  reg        [15:0]   int_reg_array_47_10_imag;
  reg        [15:0]   int_reg_array_47_11_real;
  reg        [15:0]   int_reg_array_47_11_imag;
  reg        [15:0]   int_reg_array_47_12_real;
  reg        [15:0]   int_reg_array_47_12_imag;
  reg        [15:0]   int_reg_array_47_13_real;
  reg        [15:0]   int_reg_array_47_13_imag;
  reg        [15:0]   int_reg_array_47_14_real;
  reg        [15:0]   int_reg_array_47_14_imag;
  reg        [15:0]   int_reg_array_47_15_real;
  reg        [15:0]   int_reg_array_47_15_imag;
  reg        [15:0]   int_reg_array_47_16_real;
  reg        [15:0]   int_reg_array_47_16_imag;
  reg        [15:0]   int_reg_array_47_17_real;
  reg        [15:0]   int_reg_array_47_17_imag;
  reg        [15:0]   int_reg_array_47_18_real;
  reg        [15:0]   int_reg_array_47_18_imag;
  reg        [15:0]   int_reg_array_47_19_real;
  reg        [15:0]   int_reg_array_47_19_imag;
  reg        [15:0]   int_reg_array_47_20_real;
  reg        [15:0]   int_reg_array_47_20_imag;
  reg        [15:0]   int_reg_array_47_21_real;
  reg        [15:0]   int_reg_array_47_21_imag;
  reg        [15:0]   int_reg_array_47_22_real;
  reg        [15:0]   int_reg_array_47_22_imag;
  reg        [15:0]   int_reg_array_47_23_real;
  reg        [15:0]   int_reg_array_47_23_imag;
  reg        [15:0]   int_reg_array_47_24_real;
  reg        [15:0]   int_reg_array_47_24_imag;
  reg        [15:0]   int_reg_array_47_25_real;
  reg        [15:0]   int_reg_array_47_25_imag;
  reg        [15:0]   int_reg_array_47_26_real;
  reg        [15:0]   int_reg_array_47_26_imag;
  reg        [15:0]   int_reg_array_47_27_real;
  reg        [15:0]   int_reg_array_47_27_imag;
  reg        [15:0]   int_reg_array_47_28_real;
  reg        [15:0]   int_reg_array_47_28_imag;
  reg        [15:0]   int_reg_array_47_29_real;
  reg        [15:0]   int_reg_array_47_29_imag;
  reg        [15:0]   int_reg_array_47_30_real;
  reg        [15:0]   int_reg_array_47_30_imag;
  reg        [15:0]   int_reg_array_47_31_real;
  reg        [15:0]   int_reg_array_47_31_imag;
  reg        [15:0]   int_reg_array_47_32_real;
  reg        [15:0]   int_reg_array_47_32_imag;
  reg        [15:0]   int_reg_array_47_33_real;
  reg        [15:0]   int_reg_array_47_33_imag;
  reg        [15:0]   int_reg_array_47_34_real;
  reg        [15:0]   int_reg_array_47_34_imag;
  reg        [15:0]   int_reg_array_47_35_real;
  reg        [15:0]   int_reg_array_47_35_imag;
  reg        [15:0]   int_reg_array_47_36_real;
  reg        [15:0]   int_reg_array_47_36_imag;
  reg        [15:0]   int_reg_array_47_37_real;
  reg        [15:0]   int_reg_array_47_37_imag;
  reg        [15:0]   int_reg_array_47_38_real;
  reg        [15:0]   int_reg_array_47_38_imag;
  reg        [15:0]   int_reg_array_47_39_real;
  reg        [15:0]   int_reg_array_47_39_imag;
  reg        [15:0]   int_reg_array_47_40_real;
  reg        [15:0]   int_reg_array_47_40_imag;
  reg        [15:0]   int_reg_array_47_41_real;
  reg        [15:0]   int_reg_array_47_41_imag;
  reg        [15:0]   int_reg_array_47_42_real;
  reg        [15:0]   int_reg_array_47_42_imag;
  reg        [15:0]   int_reg_array_47_43_real;
  reg        [15:0]   int_reg_array_47_43_imag;
  reg        [15:0]   int_reg_array_47_44_real;
  reg        [15:0]   int_reg_array_47_44_imag;
  reg        [15:0]   int_reg_array_47_45_real;
  reg        [15:0]   int_reg_array_47_45_imag;
  reg        [15:0]   int_reg_array_47_46_real;
  reg        [15:0]   int_reg_array_47_46_imag;
  reg        [15:0]   int_reg_array_47_47_real;
  reg        [15:0]   int_reg_array_47_47_imag;
  reg        [15:0]   int_reg_array_47_48_real;
  reg        [15:0]   int_reg_array_47_48_imag;
  reg        [15:0]   int_reg_array_47_49_real;
  reg        [15:0]   int_reg_array_47_49_imag;
  reg        [15:0]   int_reg_array_47_50_real;
  reg        [15:0]   int_reg_array_47_50_imag;
  reg        [15:0]   int_reg_array_47_51_real;
  reg        [15:0]   int_reg_array_47_51_imag;
  reg        [15:0]   int_reg_array_47_52_real;
  reg        [15:0]   int_reg_array_47_52_imag;
  reg        [15:0]   int_reg_array_47_53_real;
  reg        [15:0]   int_reg_array_47_53_imag;
  reg        [15:0]   int_reg_array_47_54_real;
  reg        [15:0]   int_reg_array_47_54_imag;
  reg        [15:0]   int_reg_array_47_55_real;
  reg        [15:0]   int_reg_array_47_55_imag;
  reg        [15:0]   int_reg_array_47_56_real;
  reg        [15:0]   int_reg_array_47_56_imag;
  reg        [15:0]   int_reg_array_47_57_real;
  reg        [15:0]   int_reg_array_47_57_imag;
  reg        [15:0]   int_reg_array_47_58_real;
  reg        [15:0]   int_reg_array_47_58_imag;
  reg        [15:0]   int_reg_array_47_59_real;
  reg        [15:0]   int_reg_array_47_59_imag;
  reg        [15:0]   int_reg_array_47_60_real;
  reg        [15:0]   int_reg_array_47_60_imag;
  reg        [15:0]   int_reg_array_47_61_real;
  reg        [15:0]   int_reg_array_47_61_imag;
  reg        [15:0]   int_reg_array_47_62_real;
  reg        [15:0]   int_reg_array_47_62_imag;
  reg        [15:0]   int_reg_array_47_63_real;
  reg        [15:0]   int_reg_array_47_63_imag;
  reg        [15:0]   int_reg_array_1_0_real;
  reg        [15:0]   int_reg_array_1_0_imag;
  reg        [15:0]   int_reg_array_1_1_real;
  reg        [15:0]   int_reg_array_1_1_imag;
  reg        [15:0]   int_reg_array_1_2_real;
  reg        [15:0]   int_reg_array_1_2_imag;
  reg        [15:0]   int_reg_array_1_3_real;
  reg        [15:0]   int_reg_array_1_3_imag;
  reg        [15:0]   int_reg_array_1_4_real;
  reg        [15:0]   int_reg_array_1_4_imag;
  reg        [15:0]   int_reg_array_1_5_real;
  reg        [15:0]   int_reg_array_1_5_imag;
  reg        [15:0]   int_reg_array_1_6_real;
  reg        [15:0]   int_reg_array_1_6_imag;
  reg        [15:0]   int_reg_array_1_7_real;
  reg        [15:0]   int_reg_array_1_7_imag;
  reg        [15:0]   int_reg_array_1_8_real;
  reg        [15:0]   int_reg_array_1_8_imag;
  reg        [15:0]   int_reg_array_1_9_real;
  reg        [15:0]   int_reg_array_1_9_imag;
  reg        [15:0]   int_reg_array_1_10_real;
  reg        [15:0]   int_reg_array_1_10_imag;
  reg        [15:0]   int_reg_array_1_11_real;
  reg        [15:0]   int_reg_array_1_11_imag;
  reg        [15:0]   int_reg_array_1_12_real;
  reg        [15:0]   int_reg_array_1_12_imag;
  reg        [15:0]   int_reg_array_1_13_real;
  reg        [15:0]   int_reg_array_1_13_imag;
  reg        [15:0]   int_reg_array_1_14_real;
  reg        [15:0]   int_reg_array_1_14_imag;
  reg        [15:0]   int_reg_array_1_15_real;
  reg        [15:0]   int_reg_array_1_15_imag;
  reg        [15:0]   int_reg_array_1_16_real;
  reg        [15:0]   int_reg_array_1_16_imag;
  reg        [15:0]   int_reg_array_1_17_real;
  reg        [15:0]   int_reg_array_1_17_imag;
  reg        [15:0]   int_reg_array_1_18_real;
  reg        [15:0]   int_reg_array_1_18_imag;
  reg        [15:0]   int_reg_array_1_19_real;
  reg        [15:0]   int_reg_array_1_19_imag;
  reg        [15:0]   int_reg_array_1_20_real;
  reg        [15:0]   int_reg_array_1_20_imag;
  reg        [15:0]   int_reg_array_1_21_real;
  reg        [15:0]   int_reg_array_1_21_imag;
  reg        [15:0]   int_reg_array_1_22_real;
  reg        [15:0]   int_reg_array_1_22_imag;
  reg        [15:0]   int_reg_array_1_23_real;
  reg        [15:0]   int_reg_array_1_23_imag;
  reg        [15:0]   int_reg_array_1_24_real;
  reg        [15:0]   int_reg_array_1_24_imag;
  reg        [15:0]   int_reg_array_1_25_real;
  reg        [15:0]   int_reg_array_1_25_imag;
  reg        [15:0]   int_reg_array_1_26_real;
  reg        [15:0]   int_reg_array_1_26_imag;
  reg        [15:0]   int_reg_array_1_27_real;
  reg        [15:0]   int_reg_array_1_27_imag;
  reg        [15:0]   int_reg_array_1_28_real;
  reg        [15:0]   int_reg_array_1_28_imag;
  reg        [15:0]   int_reg_array_1_29_real;
  reg        [15:0]   int_reg_array_1_29_imag;
  reg        [15:0]   int_reg_array_1_30_real;
  reg        [15:0]   int_reg_array_1_30_imag;
  reg        [15:0]   int_reg_array_1_31_real;
  reg        [15:0]   int_reg_array_1_31_imag;
  reg        [15:0]   int_reg_array_1_32_real;
  reg        [15:0]   int_reg_array_1_32_imag;
  reg        [15:0]   int_reg_array_1_33_real;
  reg        [15:0]   int_reg_array_1_33_imag;
  reg        [15:0]   int_reg_array_1_34_real;
  reg        [15:0]   int_reg_array_1_34_imag;
  reg        [15:0]   int_reg_array_1_35_real;
  reg        [15:0]   int_reg_array_1_35_imag;
  reg        [15:0]   int_reg_array_1_36_real;
  reg        [15:0]   int_reg_array_1_36_imag;
  reg        [15:0]   int_reg_array_1_37_real;
  reg        [15:0]   int_reg_array_1_37_imag;
  reg        [15:0]   int_reg_array_1_38_real;
  reg        [15:0]   int_reg_array_1_38_imag;
  reg        [15:0]   int_reg_array_1_39_real;
  reg        [15:0]   int_reg_array_1_39_imag;
  reg        [15:0]   int_reg_array_1_40_real;
  reg        [15:0]   int_reg_array_1_40_imag;
  reg        [15:0]   int_reg_array_1_41_real;
  reg        [15:0]   int_reg_array_1_41_imag;
  reg        [15:0]   int_reg_array_1_42_real;
  reg        [15:0]   int_reg_array_1_42_imag;
  reg        [15:0]   int_reg_array_1_43_real;
  reg        [15:0]   int_reg_array_1_43_imag;
  reg        [15:0]   int_reg_array_1_44_real;
  reg        [15:0]   int_reg_array_1_44_imag;
  reg        [15:0]   int_reg_array_1_45_real;
  reg        [15:0]   int_reg_array_1_45_imag;
  reg        [15:0]   int_reg_array_1_46_real;
  reg        [15:0]   int_reg_array_1_46_imag;
  reg        [15:0]   int_reg_array_1_47_real;
  reg        [15:0]   int_reg_array_1_47_imag;
  reg        [15:0]   int_reg_array_1_48_real;
  reg        [15:0]   int_reg_array_1_48_imag;
  reg        [15:0]   int_reg_array_1_49_real;
  reg        [15:0]   int_reg_array_1_49_imag;
  reg        [15:0]   int_reg_array_1_50_real;
  reg        [15:0]   int_reg_array_1_50_imag;
  reg        [15:0]   int_reg_array_1_51_real;
  reg        [15:0]   int_reg_array_1_51_imag;
  reg        [15:0]   int_reg_array_1_52_real;
  reg        [15:0]   int_reg_array_1_52_imag;
  reg        [15:0]   int_reg_array_1_53_real;
  reg        [15:0]   int_reg_array_1_53_imag;
  reg        [15:0]   int_reg_array_1_54_real;
  reg        [15:0]   int_reg_array_1_54_imag;
  reg        [15:0]   int_reg_array_1_55_real;
  reg        [15:0]   int_reg_array_1_55_imag;
  reg        [15:0]   int_reg_array_1_56_real;
  reg        [15:0]   int_reg_array_1_56_imag;
  reg        [15:0]   int_reg_array_1_57_real;
  reg        [15:0]   int_reg_array_1_57_imag;
  reg        [15:0]   int_reg_array_1_58_real;
  reg        [15:0]   int_reg_array_1_58_imag;
  reg        [15:0]   int_reg_array_1_59_real;
  reg        [15:0]   int_reg_array_1_59_imag;
  reg        [15:0]   int_reg_array_1_60_real;
  reg        [15:0]   int_reg_array_1_60_imag;
  reg        [15:0]   int_reg_array_1_61_real;
  reg        [15:0]   int_reg_array_1_61_imag;
  reg        [15:0]   int_reg_array_1_62_real;
  reg        [15:0]   int_reg_array_1_62_imag;
  reg        [15:0]   int_reg_array_1_63_real;
  reg        [15:0]   int_reg_array_1_63_imag;
  reg        [15:0]   int_reg_array_26_0_real;
  reg        [15:0]   int_reg_array_26_0_imag;
  reg        [15:0]   int_reg_array_26_1_real;
  reg        [15:0]   int_reg_array_26_1_imag;
  reg        [15:0]   int_reg_array_26_2_real;
  reg        [15:0]   int_reg_array_26_2_imag;
  reg        [15:0]   int_reg_array_26_3_real;
  reg        [15:0]   int_reg_array_26_3_imag;
  reg        [15:0]   int_reg_array_26_4_real;
  reg        [15:0]   int_reg_array_26_4_imag;
  reg        [15:0]   int_reg_array_26_5_real;
  reg        [15:0]   int_reg_array_26_5_imag;
  reg        [15:0]   int_reg_array_26_6_real;
  reg        [15:0]   int_reg_array_26_6_imag;
  reg        [15:0]   int_reg_array_26_7_real;
  reg        [15:0]   int_reg_array_26_7_imag;
  reg        [15:0]   int_reg_array_26_8_real;
  reg        [15:0]   int_reg_array_26_8_imag;
  reg        [15:0]   int_reg_array_26_9_real;
  reg        [15:0]   int_reg_array_26_9_imag;
  reg        [15:0]   int_reg_array_26_10_real;
  reg        [15:0]   int_reg_array_26_10_imag;
  reg        [15:0]   int_reg_array_26_11_real;
  reg        [15:0]   int_reg_array_26_11_imag;
  reg        [15:0]   int_reg_array_26_12_real;
  reg        [15:0]   int_reg_array_26_12_imag;
  reg        [15:0]   int_reg_array_26_13_real;
  reg        [15:0]   int_reg_array_26_13_imag;
  reg        [15:0]   int_reg_array_26_14_real;
  reg        [15:0]   int_reg_array_26_14_imag;
  reg        [15:0]   int_reg_array_26_15_real;
  reg        [15:0]   int_reg_array_26_15_imag;
  reg        [15:0]   int_reg_array_26_16_real;
  reg        [15:0]   int_reg_array_26_16_imag;
  reg        [15:0]   int_reg_array_26_17_real;
  reg        [15:0]   int_reg_array_26_17_imag;
  reg        [15:0]   int_reg_array_26_18_real;
  reg        [15:0]   int_reg_array_26_18_imag;
  reg        [15:0]   int_reg_array_26_19_real;
  reg        [15:0]   int_reg_array_26_19_imag;
  reg        [15:0]   int_reg_array_26_20_real;
  reg        [15:0]   int_reg_array_26_20_imag;
  reg        [15:0]   int_reg_array_26_21_real;
  reg        [15:0]   int_reg_array_26_21_imag;
  reg        [15:0]   int_reg_array_26_22_real;
  reg        [15:0]   int_reg_array_26_22_imag;
  reg        [15:0]   int_reg_array_26_23_real;
  reg        [15:0]   int_reg_array_26_23_imag;
  reg        [15:0]   int_reg_array_26_24_real;
  reg        [15:0]   int_reg_array_26_24_imag;
  reg        [15:0]   int_reg_array_26_25_real;
  reg        [15:0]   int_reg_array_26_25_imag;
  reg        [15:0]   int_reg_array_26_26_real;
  reg        [15:0]   int_reg_array_26_26_imag;
  reg        [15:0]   int_reg_array_26_27_real;
  reg        [15:0]   int_reg_array_26_27_imag;
  reg        [15:0]   int_reg_array_26_28_real;
  reg        [15:0]   int_reg_array_26_28_imag;
  reg        [15:0]   int_reg_array_26_29_real;
  reg        [15:0]   int_reg_array_26_29_imag;
  reg        [15:0]   int_reg_array_26_30_real;
  reg        [15:0]   int_reg_array_26_30_imag;
  reg        [15:0]   int_reg_array_26_31_real;
  reg        [15:0]   int_reg_array_26_31_imag;
  reg        [15:0]   int_reg_array_26_32_real;
  reg        [15:0]   int_reg_array_26_32_imag;
  reg        [15:0]   int_reg_array_26_33_real;
  reg        [15:0]   int_reg_array_26_33_imag;
  reg        [15:0]   int_reg_array_26_34_real;
  reg        [15:0]   int_reg_array_26_34_imag;
  reg        [15:0]   int_reg_array_26_35_real;
  reg        [15:0]   int_reg_array_26_35_imag;
  reg        [15:0]   int_reg_array_26_36_real;
  reg        [15:0]   int_reg_array_26_36_imag;
  reg        [15:0]   int_reg_array_26_37_real;
  reg        [15:0]   int_reg_array_26_37_imag;
  reg        [15:0]   int_reg_array_26_38_real;
  reg        [15:0]   int_reg_array_26_38_imag;
  reg        [15:0]   int_reg_array_26_39_real;
  reg        [15:0]   int_reg_array_26_39_imag;
  reg        [15:0]   int_reg_array_26_40_real;
  reg        [15:0]   int_reg_array_26_40_imag;
  reg        [15:0]   int_reg_array_26_41_real;
  reg        [15:0]   int_reg_array_26_41_imag;
  reg        [15:0]   int_reg_array_26_42_real;
  reg        [15:0]   int_reg_array_26_42_imag;
  reg        [15:0]   int_reg_array_26_43_real;
  reg        [15:0]   int_reg_array_26_43_imag;
  reg        [15:0]   int_reg_array_26_44_real;
  reg        [15:0]   int_reg_array_26_44_imag;
  reg        [15:0]   int_reg_array_26_45_real;
  reg        [15:0]   int_reg_array_26_45_imag;
  reg        [15:0]   int_reg_array_26_46_real;
  reg        [15:0]   int_reg_array_26_46_imag;
  reg        [15:0]   int_reg_array_26_47_real;
  reg        [15:0]   int_reg_array_26_47_imag;
  reg        [15:0]   int_reg_array_26_48_real;
  reg        [15:0]   int_reg_array_26_48_imag;
  reg        [15:0]   int_reg_array_26_49_real;
  reg        [15:0]   int_reg_array_26_49_imag;
  reg        [15:0]   int_reg_array_26_50_real;
  reg        [15:0]   int_reg_array_26_50_imag;
  reg        [15:0]   int_reg_array_26_51_real;
  reg        [15:0]   int_reg_array_26_51_imag;
  reg        [15:0]   int_reg_array_26_52_real;
  reg        [15:0]   int_reg_array_26_52_imag;
  reg        [15:0]   int_reg_array_26_53_real;
  reg        [15:0]   int_reg_array_26_53_imag;
  reg        [15:0]   int_reg_array_26_54_real;
  reg        [15:0]   int_reg_array_26_54_imag;
  reg        [15:0]   int_reg_array_26_55_real;
  reg        [15:0]   int_reg_array_26_55_imag;
  reg        [15:0]   int_reg_array_26_56_real;
  reg        [15:0]   int_reg_array_26_56_imag;
  reg        [15:0]   int_reg_array_26_57_real;
  reg        [15:0]   int_reg_array_26_57_imag;
  reg        [15:0]   int_reg_array_26_58_real;
  reg        [15:0]   int_reg_array_26_58_imag;
  reg        [15:0]   int_reg_array_26_59_real;
  reg        [15:0]   int_reg_array_26_59_imag;
  reg        [15:0]   int_reg_array_26_60_real;
  reg        [15:0]   int_reg_array_26_60_imag;
  reg        [15:0]   int_reg_array_26_61_real;
  reg        [15:0]   int_reg_array_26_61_imag;
  reg        [15:0]   int_reg_array_26_62_real;
  reg        [15:0]   int_reg_array_26_62_imag;
  reg        [15:0]   int_reg_array_26_63_real;
  reg        [15:0]   int_reg_array_26_63_imag;
  reg        [15:0]   int_reg_array_9_0_real;
  reg        [15:0]   int_reg_array_9_0_imag;
  reg        [15:0]   int_reg_array_9_1_real;
  reg        [15:0]   int_reg_array_9_1_imag;
  reg        [15:0]   int_reg_array_9_2_real;
  reg        [15:0]   int_reg_array_9_2_imag;
  reg        [15:0]   int_reg_array_9_3_real;
  reg        [15:0]   int_reg_array_9_3_imag;
  reg        [15:0]   int_reg_array_9_4_real;
  reg        [15:0]   int_reg_array_9_4_imag;
  reg        [15:0]   int_reg_array_9_5_real;
  reg        [15:0]   int_reg_array_9_5_imag;
  reg        [15:0]   int_reg_array_9_6_real;
  reg        [15:0]   int_reg_array_9_6_imag;
  reg        [15:0]   int_reg_array_9_7_real;
  reg        [15:0]   int_reg_array_9_7_imag;
  reg        [15:0]   int_reg_array_9_8_real;
  reg        [15:0]   int_reg_array_9_8_imag;
  reg        [15:0]   int_reg_array_9_9_real;
  reg        [15:0]   int_reg_array_9_9_imag;
  reg        [15:0]   int_reg_array_9_10_real;
  reg        [15:0]   int_reg_array_9_10_imag;
  reg        [15:0]   int_reg_array_9_11_real;
  reg        [15:0]   int_reg_array_9_11_imag;
  reg        [15:0]   int_reg_array_9_12_real;
  reg        [15:0]   int_reg_array_9_12_imag;
  reg        [15:0]   int_reg_array_9_13_real;
  reg        [15:0]   int_reg_array_9_13_imag;
  reg        [15:0]   int_reg_array_9_14_real;
  reg        [15:0]   int_reg_array_9_14_imag;
  reg        [15:0]   int_reg_array_9_15_real;
  reg        [15:0]   int_reg_array_9_15_imag;
  reg        [15:0]   int_reg_array_9_16_real;
  reg        [15:0]   int_reg_array_9_16_imag;
  reg        [15:0]   int_reg_array_9_17_real;
  reg        [15:0]   int_reg_array_9_17_imag;
  reg        [15:0]   int_reg_array_9_18_real;
  reg        [15:0]   int_reg_array_9_18_imag;
  reg        [15:0]   int_reg_array_9_19_real;
  reg        [15:0]   int_reg_array_9_19_imag;
  reg        [15:0]   int_reg_array_9_20_real;
  reg        [15:0]   int_reg_array_9_20_imag;
  reg        [15:0]   int_reg_array_9_21_real;
  reg        [15:0]   int_reg_array_9_21_imag;
  reg        [15:0]   int_reg_array_9_22_real;
  reg        [15:0]   int_reg_array_9_22_imag;
  reg        [15:0]   int_reg_array_9_23_real;
  reg        [15:0]   int_reg_array_9_23_imag;
  reg        [15:0]   int_reg_array_9_24_real;
  reg        [15:0]   int_reg_array_9_24_imag;
  reg        [15:0]   int_reg_array_9_25_real;
  reg        [15:0]   int_reg_array_9_25_imag;
  reg        [15:0]   int_reg_array_9_26_real;
  reg        [15:0]   int_reg_array_9_26_imag;
  reg        [15:0]   int_reg_array_9_27_real;
  reg        [15:0]   int_reg_array_9_27_imag;
  reg        [15:0]   int_reg_array_9_28_real;
  reg        [15:0]   int_reg_array_9_28_imag;
  reg        [15:0]   int_reg_array_9_29_real;
  reg        [15:0]   int_reg_array_9_29_imag;
  reg        [15:0]   int_reg_array_9_30_real;
  reg        [15:0]   int_reg_array_9_30_imag;
  reg        [15:0]   int_reg_array_9_31_real;
  reg        [15:0]   int_reg_array_9_31_imag;
  reg        [15:0]   int_reg_array_9_32_real;
  reg        [15:0]   int_reg_array_9_32_imag;
  reg        [15:0]   int_reg_array_9_33_real;
  reg        [15:0]   int_reg_array_9_33_imag;
  reg        [15:0]   int_reg_array_9_34_real;
  reg        [15:0]   int_reg_array_9_34_imag;
  reg        [15:0]   int_reg_array_9_35_real;
  reg        [15:0]   int_reg_array_9_35_imag;
  reg        [15:0]   int_reg_array_9_36_real;
  reg        [15:0]   int_reg_array_9_36_imag;
  reg        [15:0]   int_reg_array_9_37_real;
  reg        [15:0]   int_reg_array_9_37_imag;
  reg        [15:0]   int_reg_array_9_38_real;
  reg        [15:0]   int_reg_array_9_38_imag;
  reg        [15:0]   int_reg_array_9_39_real;
  reg        [15:0]   int_reg_array_9_39_imag;
  reg        [15:0]   int_reg_array_9_40_real;
  reg        [15:0]   int_reg_array_9_40_imag;
  reg        [15:0]   int_reg_array_9_41_real;
  reg        [15:0]   int_reg_array_9_41_imag;
  reg        [15:0]   int_reg_array_9_42_real;
  reg        [15:0]   int_reg_array_9_42_imag;
  reg        [15:0]   int_reg_array_9_43_real;
  reg        [15:0]   int_reg_array_9_43_imag;
  reg        [15:0]   int_reg_array_9_44_real;
  reg        [15:0]   int_reg_array_9_44_imag;
  reg        [15:0]   int_reg_array_9_45_real;
  reg        [15:0]   int_reg_array_9_45_imag;
  reg        [15:0]   int_reg_array_9_46_real;
  reg        [15:0]   int_reg_array_9_46_imag;
  reg        [15:0]   int_reg_array_9_47_real;
  reg        [15:0]   int_reg_array_9_47_imag;
  reg        [15:0]   int_reg_array_9_48_real;
  reg        [15:0]   int_reg_array_9_48_imag;
  reg        [15:0]   int_reg_array_9_49_real;
  reg        [15:0]   int_reg_array_9_49_imag;
  reg        [15:0]   int_reg_array_9_50_real;
  reg        [15:0]   int_reg_array_9_50_imag;
  reg        [15:0]   int_reg_array_9_51_real;
  reg        [15:0]   int_reg_array_9_51_imag;
  reg        [15:0]   int_reg_array_9_52_real;
  reg        [15:0]   int_reg_array_9_52_imag;
  reg        [15:0]   int_reg_array_9_53_real;
  reg        [15:0]   int_reg_array_9_53_imag;
  reg        [15:0]   int_reg_array_9_54_real;
  reg        [15:0]   int_reg_array_9_54_imag;
  reg        [15:0]   int_reg_array_9_55_real;
  reg        [15:0]   int_reg_array_9_55_imag;
  reg        [15:0]   int_reg_array_9_56_real;
  reg        [15:0]   int_reg_array_9_56_imag;
  reg        [15:0]   int_reg_array_9_57_real;
  reg        [15:0]   int_reg_array_9_57_imag;
  reg        [15:0]   int_reg_array_9_58_real;
  reg        [15:0]   int_reg_array_9_58_imag;
  reg        [15:0]   int_reg_array_9_59_real;
  reg        [15:0]   int_reg_array_9_59_imag;
  reg        [15:0]   int_reg_array_9_60_real;
  reg        [15:0]   int_reg_array_9_60_imag;
  reg        [15:0]   int_reg_array_9_61_real;
  reg        [15:0]   int_reg_array_9_61_imag;
  reg        [15:0]   int_reg_array_9_62_real;
  reg        [15:0]   int_reg_array_9_62_imag;
  reg        [15:0]   int_reg_array_9_63_real;
  reg        [15:0]   int_reg_array_9_63_imag;
  reg        [15:0]   int_reg_array_60_0_real;
  reg        [15:0]   int_reg_array_60_0_imag;
  reg        [15:0]   int_reg_array_60_1_real;
  reg        [15:0]   int_reg_array_60_1_imag;
  reg        [15:0]   int_reg_array_60_2_real;
  reg        [15:0]   int_reg_array_60_2_imag;
  reg        [15:0]   int_reg_array_60_3_real;
  reg        [15:0]   int_reg_array_60_3_imag;
  reg        [15:0]   int_reg_array_60_4_real;
  reg        [15:0]   int_reg_array_60_4_imag;
  reg        [15:0]   int_reg_array_60_5_real;
  reg        [15:0]   int_reg_array_60_5_imag;
  reg        [15:0]   int_reg_array_60_6_real;
  reg        [15:0]   int_reg_array_60_6_imag;
  reg        [15:0]   int_reg_array_60_7_real;
  reg        [15:0]   int_reg_array_60_7_imag;
  reg        [15:0]   int_reg_array_60_8_real;
  reg        [15:0]   int_reg_array_60_8_imag;
  reg        [15:0]   int_reg_array_60_9_real;
  reg        [15:0]   int_reg_array_60_9_imag;
  reg        [15:0]   int_reg_array_60_10_real;
  reg        [15:0]   int_reg_array_60_10_imag;
  reg        [15:0]   int_reg_array_60_11_real;
  reg        [15:0]   int_reg_array_60_11_imag;
  reg        [15:0]   int_reg_array_60_12_real;
  reg        [15:0]   int_reg_array_60_12_imag;
  reg        [15:0]   int_reg_array_60_13_real;
  reg        [15:0]   int_reg_array_60_13_imag;
  reg        [15:0]   int_reg_array_60_14_real;
  reg        [15:0]   int_reg_array_60_14_imag;
  reg        [15:0]   int_reg_array_60_15_real;
  reg        [15:0]   int_reg_array_60_15_imag;
  reg        [15:0]   int_reg_array_60_16_real;
  reg        [15:0]   int_reg_array_60_16_imag;
  reg        [15:0]   int_reg_array_60_17_real;
  reg        [15:0]   int_reg_array_60_17_imag;
  reg        [15:0]   int_reg_array_60_18_real;
  reg        [15:0]   int_reg_array_60_18_imag;
  reg        [15:0]   int_reg_array_60_19_real;
  reg        [15:0]   int_reg_array_60_19_imag;
  reg        [15:0]   int_reg_array_60_20_real;
  reg        [15:0]   int_reg_array_60_20_imag;
  reg        [15:0]   int_reg_array_60_21_real;
  reg        [15:0]   int_reg_array_60_21_imag;
  reg        [15:0]   int_reg_array_60_22_real;
  reg        [15:0]   int_reg_array_60_22_imag;
  reg        [15:0]   int_reg_array_60_23_real;
  reg        [15:0]   int_reg_array_60_23_imag;
  reg        [15:0]   int_reg_array_60_24_real;
  reg        [15:0]   int_reg_array_60_24_imag;
  reg        [15:0]   int_reg_array_60_25_real;
  reg        [15:0]   int_reg_array_60_25_imag;
  reg        [15:0]   int_reg_array_60_26_real;
  reg        [15:0]   int_reg_array_60_26_imag;
  reg        [15:0]   int_reg_array_60_27_real;
  reg        [15:0]   int_reg_array_60_27_imag;
  reg        [15:0]   int_reg_array_60_28_real;
  reg        [15:0]   int_reg_array_60_28_imag;
  reg        [15:0]   int_reg_array_60_29_real;
  reg        [15:0]   int_reg_array_60_29_imag;
  reg        [15:0]   int_reg_array_60_30_real;
  reg        [15:0]   int_reg_array_60_30_imag;
  reg        [15:0]   int_reg_array_60_31_real;
  reg        [15:0]   int_reg_array_60_31_imag;
  reg        [15:0]   int_reg_array_60_32_real;
  reg        [15:0]   int_reg_array_60_32_imag;
  reg        [15:0]   int_reg_array_60_33_real;
  reg        [15:0]   int_reg_array_60_33_imag;
  reg        [15:0]   int_reg_array_60_34_real;
  reg        [15:0]   int_reg_array_60_34_imag;
  reg        [15:0]   int_reg_array_60_35_real;
  reg        [15:0]   int_reg_array_60_35_imag;
  reg        [15:0]   int_reg_array_60_36_real;
  reg        [15:0]   int_reg_array_60_36_imag;
  reg        [15:0]   int_reg_array_60_37_real;
  reg        [15:0]   int_reg_array_60_37_imag;
  reg        [15:0]   int_reg_array_60_38_real;
  reg        [15:0]   int_reg_array_60_38_imag;
  reg        [15:0]   int_reg_array_60_39_real;
  reg        [15:0]   int_reg_array_60_39_imag;
  reg        [15:0]   int_reg_array_60_40_real;
  reg        [15:0]   int_reg_array_60_40_imag;
  reg        [15:0]   int_reg_array_60_41_real;
  reg        [15:0]   int_reg_array_60_41_imag;
  reg        [15:0]   int_reg_array_60_42_real;
  reg        [15:0]   int_reg_array_60_42_imag;
  reg        [15:0]   int_reg_array_60_43_real;
  reg        [15:0]   int_reg_array_60_43_imag;
  reg        [15:0]   int_reg_array_60_44_real;
  reg        [15:0]   int_reg_array_60_44_imag;
  reg        [15:0]   int_reg_array_60_45_real;
  reg        [15:0]   int_reg_array_60_45_imag;
  reg        [15:0]   int_reg_array_60_46_real;
  reg        [15:0]   int_reg_array_60_46_imag;
  reg        [15:0]   int_reg_array_60_47_real;
  reg        [15:0]   int_reg_array_60_47_imag;
  reg        [15:0]   int_reg_array_60_48_real;
  reg        [15:0]   int_reg_array_60_48_imag;
  reg        [15:0]   int_reg_array_60_49_real;
  reg        [15:0]   int_reg_array_60_49_imag;
  reg        [15:0]   int_reg_array_60_50_real;
  reg        [15:0]   int_reg_array_60_50_imag;
  reg        [15:0]   int_reg_array_60_51_real;
  reg        [15:0]   int_reg_array_60_51_imag;
  reg        [15:0]   int_reg_array_60_52_real;
  reg        [15:0]   int_reg_array_60_52_imag;
  reg        [15:0]   int_reg_array_60_53_real;
  reg        [15:0]   int_reg_array_60_53_imag;
  reg        [15:0]   int_reg_array_60_54_real;
  reg        [15:0]   int_reg_array_60_54_imag;
  reg        [15:0]   int_reg_array_60_55_real;
  reg        [15:0]   int_reg_array_60_55_imag;
  reg        [15:0]   int_reg_array_60_56_real;
  reg        [15:0]   int_reg_array_60_56_imag;
  reg        [15:0]   int_reg_array_60_57_real;
  reg        [15:0]   int_reg_array_60_57_imag;
  reg        [15:0]   int_reg_array_60_58_real;
  reg        [15:0]   int_reg_array_60_58_imag;
  reg        [15:0]   int_reg_array_60_59_real;
  reg        [15:0]   int_reg_array_60_59_imag;
  reg        [15:0]   int_reg_array_60_60_real;
  reg        [15:0]   int_reg_array_60_60_imag;
  reg        [15:0]   int_reg_array_60_61_real;
  reg        [15:0]   int_reg_array_60_61_imag;
  reg        [15:0]   int_reg_array_60_62_real;
  reg        [15:0]   int_reg_array_60_62_imag;
  reg        [15:0]   int_reg_array_60_63_real;
  reg        [15:0]   int_reg_array_60_63_imag;
  reg        [31:0]   load_data_area_current_addr;
  reg        [31:0]   Axi4Incr_result;
  wire       [19:0]   Axi4Incr_highCat;
  wire       [0:0]    Axi4Incr_sizeValue;
  wire       [11:0]   Axi4Incr_alignMask;
  wire       [11:0]   Axi4Incr_base;
  wire       [11:0]   Axi4Incr_baseIncr;
  reg        [1:0]    _zz_16_;
  wire       [1:0]    Axi4Incr_wrapCase;
  reg        [31:0]   _zz_9__regNext;
  wire       [5:0]    _zz_17_;
  wire       [63:0]   _zz_18_;
  wire                _zz_19_;
  wire                _zz_20_;
  wire                _zz_21_;
  wire                _zz_22_;
  wire                _zz_23_;
  wire                _zz_24_;
  wire                _zz_25_;
  wire                _zz_26_;
  wire                _zz_27_;
  wire                _zz_28_;
  wire                _zz_29_;
  wire                _zz_30_;
  wire                _zz_31_;
  wire                _zz_32_;
  wire                _zz_33_;
  wire                _zz_34_;
  wire                _zz_35_;
  wire                _zz_36_;
  wire                _zz_37_;
  wire                _zz_38_;
  wire                _zz_39_;
  wire                _zz_40_;
  wire                _zz_41_;
  wire                _zz_42_;
  wire                _zz_43_;
  wire                _zz_44_;
  wire                _zz_45_;
  wire                _zz_46_;
  wire                _zz_47_;
  wire                _zz_48_;
  wire                _zz_49_;
  wire                _zz_50_;
  wire                _zz_51_;
  wire                _zz_52_;
  wire                _zz_53_;
  wire                _zz_54_;
  wire                _zz_55_;
  wire                _zz_56_;
  wire                _zz_57_;
  wire                _zz_58_;
  wire                _zz_59_;
  wire                _zz_60_;
  wire                _zz_61_;
  wire                _zz_62_;
  wire                _zz_63_;
  wire                _zz_64_;
  wire                _zz_65_;
  wire                _zz_66_;
  wire                _zz_67_;
  wire                _zz_68_;
  wire                _zz_69_;
  wire                _zz_70_;
  wire                _zz_71_;
  wire                _zz_72_;
  wire                _zz_73_;
  wire                _zz_74_;
  wire                _zz_75_;
  wire                _zz_76_;
  wire                _zz_77_;
  wire                _zz_78_;
  wire                _zz_79_;
  wire                _zz_80_;
  wire                _zz_81_;
  wire                _zz_82_;
  wire       [31:0]   _zz_83_;
  wire       [15:0]   _zz_84_;
  wire       [15:0]   _zz_85_;
  wire       [5:0]    _zz_86_;
  wire       [63:0]   _zz_87_;
  wire                _zz_88_;
  wire                _zz_89_;
  wire                _zz_90_;
  wire                _zz_91_;
  wire                _zz_92_;
  wire                _zz_93_;
  wire                _zz_94_;
  wire                _zz_95_;
  wire                _zz_96_;
  wire                _zz_97_;
  wire                _zz_98_;
  wire                _zz_99_;
  wire                _zz_100_;
  wire                _zz_101_;
  wire                _zz_102_;
  wire                _zz_103_;
  wire                _zz_104_;
  wire                _zz_105_;
  wire                _zz_106_;
  wire                _zz_107_;
  wire                _zz_108_;
  wire                _zz_109_;
  wire                _zz_110_;
  wire                _zz_111_;
  wire                _zz_112_;
  wire                _zz_113_;
  wire                _zz_114_;
  wire                _zz_115_;
  wire                _zz_116_;
  wire                _zz_117_;
  wire                _zz_118_;
  wire                _zz_119_;
  wire                _zz_120_;
  wire                _zz_121_;
  wire                _zz_122_;
  wire                _zz_123_;
  wire                _zz_124_;
  wire                _zz_125_;
  wire                _zz_126_;
  wire                _zz_127_;
  wire                _zz_128_;
  wire                _zz_129_;
  wire                _zz_130_;
  wire                _zz_131_;
  wire                _zz_132_;
  wire                _zz_133_;
  wire                _zz_134_;
  wire                _zz_135_;
  wire                _zz_136_;
  wire                _zz_137_;
  wire                _zz_138_;
  wire                _zz_139_;
  wire                _zz_140_;
  wire                _zz_141_;
  wire                _zz_142_;
  wire                _zz_143_;
  wire                _zz_144_;
  wire                _zz_145_;
  wire                _zz_146_;
  wire                _zz_147_;
  wire                _zz_148_;
  wire                _zz_149_;
  wire                _zz_150_;
  wire                _zz_151_;
  wire       [31:0]   _zz_152_;
  wire       [15:0]   _zz_153_;
  wire       [15:0]   _zz_154_;
  wire       [5:0]    _zz_155_;
  wire       [63:0]   _zz_156_;
  wire                _zz_157_;
  wire                _zz_158_;
  wire                _zz_159_;
  wire                _zz_160_;
  wire                _zz_161_;
  wire                _zz_162_;
  wire                _zz_163_;
  wire                _zz_164_;
  wire                _zz_165_;
  wire                _zz_166_;
  wire                _zz_167_;
  wire                _zz_168_;
  wire                _zz_169_;
  wire                _zz_170_;
  wire                _zz_171_;
  wire                _zz_172_;
  wire                _zz_173_;
  wire                _zz_174_;
  wire                _zz_175_;
  wire                _zz_176_;
  wire                _zz_177_;
  wire                _zz_178_;
  wire                _zz_179_;
  wire                _zz_180_;
  wire                _zz_181_;
  wire                _zz_182_;
  wire                _zz_183_;
  wire                _zz_184_;
  wire                _zz_185_;
  wire                _zz_186_;
  wire                _zz_187_;
  wire                _zz_188_;
  wire                _zz_189_;
  wire                _zz_190_;
  wire                _zz_191_;
  wire                _zz_192_;
  wire                _zz_193_;
  wire                _zz_194_;
  wire                _zz_195_;
  wire                _zz_196_;
  wire                _zz_197_;
  wire                _zz_198_;
  wire                _zz_199_;
  wire                _zz_200_;
  wire                _zz_201_;
  wire                _zz_202_;
  wire                _zz_203_;
  wire                _zz_204_;
  wire                _zz_205_;
  wire                _zz_206_;
  wire                _zz_207_;
  wire                _zz_208_;
  wire                _zz_209_;
  wire                _zz_210_;
  wire                _zz_211_;
  wire                _zz_212_;
  wire                _zz_213_;
  wire                _zz_214_;
  wire                _zz_215_;
  wire                _zz_216_;
  wire                _zz_217_;
  wire                _zz_218_;
  wire                _zz_219_;
  wire                _zz_220_;
  wire       [31:0]   _zz_221_;
  wire       [15:0]   _zz_222_;
  wire       [15:0]   _zz_223_;
  wire       [5:0]    _zz_224_;
  wire       [63:0]   _zz_225_;
  wire                _zz_226_;
  wire                _zz_227_;
  wire                _zz_228_;
  wire                _zz_229_;
  wire                _zz_230_;
  wire                _zz_231_;
  wire                _zz_232_;
  wire                _zz_233_;
  wire                _zz_234_;
  wire                _zz_235_;
  wire                _zz_236_;
  wire                _zz_237_;
  wire                _zz_238_;
  wire                _zz_239_;
  wire                _zz_240_;
  wire                _zz_241_;
  wire                _zz_242_;
  wire                _zz_243_;
  wire                _zz_244_;
  wire                _zz_245_;
  wire                _zz_246_;
  wire                _zz_247_;
  wire                _zz_248_;
  wire                _zz_249_;
  wire                _zz_250_;
  wire                _zz_251_;
  wire                _zz_252_;
  wire                _zz_253_;
  wire                _zz_254_;
  wire                _zz_255_;
  wire                _zz_256_;
  wire                _zz_257_;
  wire                _zz_258_;
  wire                _zz_259_;
  wire                _zz_260_;
  wire                _zz_261_;
  wire                _zz_262_;
  wire                _zz_263_;
  wire                _zz_264_;
  wire                _zz_265_;
  wire                _zz_266_;
  wire                _zz_267_;
  wire                _zz_268_;
  wire                _zz_269_;
  wire                _zz_270_;
  wire                _zz_271_;
  wire                _zz_272_;
  wire                _zz_273_;
  wire                _zz_274_;
  wire                _zz_275_;
  wire                _zz_276_;
  wire                _zz_277_;
  wire                _zz_278_;
  wire                _zz_279_;
  wire                _zz_280_;
  wire                _zz_281_;
  wire                _zz_282_;
  wire                _zz_283_;
  wire                _zz_284_;
  wire                _zz_285_;
  wire                _zz_286_;
  wire                _zz_287_;
  wire                _zz_288_;
  wire                _zz_289_;
  wire       [31:0]   _zz_290_;
  wire       [15:0]   _zz_291_;
  wire       [15:0]   _zz_292_;
  wire       [5:0]    _zz_293_;
  wire       [63:0]   _zz_294_;
  wire                _zz_295_;
  wire                _zz_296_;
  wire                _zz_297_;
  wire                _zz_298_;
  wire                _zz_299_;
  wire                _zz_300_;
  wire                _zz_301_;
  wire                _zz_302_;
  wire                _zz_303_;
  wire                _zz_304_;
  wire                _zz_305_;
  wire                _zz_306_;
  wire                _zz_307_;
  wire                _zz_308_;
  wire                _zz_309_;
  wire                _zz_310_;
  wire                _zz_311_;
  wire                _zz_312_;
  wire                _zz_313_;
  wire                _zz_314_;
  wire                _zz_315_;
  wire                _zz_316_;
  wire                _zz_317_;
  wire                _zz_318_;
  wire                _zz_319_;
  wire                _zz_320_;
  wire                _zz_321_;
  wire                _zz_322_;
  wire                _zz_323_;
  wire                _zz_324_;
  wire                _zz_325_;
  wire                _zz_326_;
  wire                _zz_327_;
  wire                _zz_328_;
  wire                _zz_329_;
  wire                _zz_330_;
  wire                _zz_331_;
  wire                _zz_332_;
  wire                _zz_333_;
  wire                _zz_334_;
  wire                _zz_335_;
  wire                _zz_336_;
  wire                _zz_337_;
  wire                _zz_338_;
  wire                _zz_339_;
  wire                _zz_340_;
  wire                _zz_341_;
  wire                _zz_342_;
  wire                _zz_343_;
  wire                _zz_344_;
  wire                _zz_345_;
  wire                _zz_346_;
  wire                _zz_347_;
  wire                _zz_348_;
  wire                _zz_349_;
  wire                _zz_350_;
  wire                _zz_351_;
  wire                _zz_352_;
  wire                _zz_353_;
  wire                _zz_354_;
  wire                _zz_355_;
  wire                _zz_356_;
  wire                _zz_357_;
  wire                _zz_358_;
  wire       [31:0]   _zz_359_;
  wire       [15:0]   _zz_360_;
  wire       [15:0]   _zz_361_;
  wire       [5:0]    _zz_362_;
  wire       [63:0]   _zz_363_;
  wire                _zz_364_;
  wire                _zz_365_;
  wire                _zz_366_;
  wire                _zz_367_;
  wire                _zz_368_;
  wire                _zz_369_;
  wire                _zz_370_;
  wire                _zz_371_;
  wire                _zz_372_;
  wire                _zz_373_;
  wire                _zz_374_;
  wire                _zz_375_;
  wire                _zz_376_;
  wire                _zz_377_;
  wire                _zz_378_;
  wire                _zz_379_;
  wire                _zz_380_;
  wire                _zz_381_;
  wire                _zz_382_;
  wire                _zz_383_;
  wire                _zz_384_;
  wire                _zz_385_;
  wire                _zz_386_;
  wire                _zz_387_;
  wire                _zz_388_;
  wire                _zz_389_;
  wire                _zz_390_;
  wire                _zz_391_;
  wire                _zz_392_;
  wire                _zz_393_;
  wire                _zz_394_;
  wire                _zz_395_;
  wire                _zz_396_;
  wire                _zz_397_;
  wire                _zz_398_;
  wire                _zz_399_;
  wire                _zz_400_;
  wire                _zz_401_;
  wire                _zz_402_;
  wire                _zz_403_;
  wire                _zz_404_;
  wire                _zz_405_;
  wire                _zz_406_;
  wire                _zz_407_;
  wire                _zz_408_;
  wire                _zz_409_;
  wire                _zz_410_;
  wire                _zz_411_;
  wire                _zz_412_;
  wire                _zz_413_;
  wire                _zz_414_;
  wire                _zz_415_;
  wire                _zz_416_;
  wire                _zz_417_;
  wire                _zz_418_;
  wire                _zz_419_;
  wire                _zz_420_;
  wire                _zz_421_;
  wire                _zz_422_;
  wire                _zz_423_;
  wire                _zz_424_;
  wire                _zz_425_;
  wire                _zz_426_;
  wire                _zz_427_;
  wire       [31:0]   _zz_428_;
  wire       [15:0]   _zz_429_;
  wire       [15:0]   _zz_430_;
  wire       [5:0]    _zz_431_;
  wire       [63:0]   _zz_432_;
  wire                _zz_433_;
  wire                _zz_434_;
  wire                _zz_435_;
  wire                _zz_436_;
  wire                _zz_437_;
  wire                _zz_438_;
  wire                _zz_439_;
  wire                _zz_440_;
  wire                _zz_441_;
  wire                _zz_442_;
  wire                _zz_443_;
  wire                _zz_444_;
  wire                _zz_445_;
  wire                _zz_446_;
  wire                _zz_447_;
  wire                _zz_448_;
  wire                _zz_449_;
  wire                _zz_450_;
  wire                _zz_451_;
  wire                _zz_452_;
  wire                _zz_453_;
  wire                _zz_454_;
  wire                _zz_455_;
  wire                _zz_456_;
  wire                _zz_457_;
  wire                _zz_458_;
  wire                _zz_459_;
  wire                _zz_460_;
  wire                _zz_461_;
  wire                _zz_462_;
  wire                _zz_463_;
  wire                _zz_464_;
  wire                _zz_465_;
  wire                _zz_466_;
  wire                _zz_467_;
  wire                _zz_468_;
  wire                _zz_469_;
  wire                _zz_470_;
  wire                _zz_471_;
  wire                _zz_472_;
  wire                _zz_473_;
  wire                _zz_474_;
  wire                _zz_475_;
  wire                _zz_476_;
  wire                _zz_477_;
  wire                _zz_478_;
  wire                _zz_479_;
  wire                _zz_480_;
  wire                _zz_481_;
  wire                _zz_482_;
  wire                _zz_483_;
  wire                _zz_484_;
  wire                _zz_485_;
  wire                _zz_486_;
  wire                _zz_487_;
  wire                _zz_488_;
  wire                _zz_489_;
  wire                _zz_490_;
  wire                _zz_491_;
  wire                _zz_492_;
  wire                _zz_493_;
  wire                _zz_494_;
  wire                _zz_495_;
  wire                _zz_496_;
  wire       [31:0]   _zz_497_;
  wire       [15:0]   _zz_498_;
  wire       [15:0]   _zz_499_;
  wire       [5:0]    _zz_500_;
  wire       [63:0]   _zz_501_;
  wire                _zz_502_;
  wire                _zz_503_;
  wire                _zz_504_;
  wire                _zz_505_;
  wire                _zz_506_;
  wire                _zz_507_;
  wire                _zz_508_;
  wire                _zz_509_;
  wire                _zz_510_;
  wire                _zz_511_;
  wire                _zz_512_;
  wire                _zz_513_;
  wire                _zz_514_;
  wire                _zz_515_;
  wire                _zz_516_;
  wire                _zz_517_;
  wire                _zz_518_;
  wire                _zz_519_;
  wire                _zz_520_;
  wire                _zz_521_;
  wire                _zz_522_;
  wire                _zz_523_;
  wire                _zz_524_;
  wire                _zz_525_;
  wire                _zz_526_;
  wire                _zz_527_;
  wire                _zz_528_;
  wire                _zz_529_;
  wire                _zz_530_;
  wire                _zz_531_;
  wire                _zz_532_;
  wire                _zz_533_;
  wire                _zz_534_;
  wire                _zz_535_;
  wire                _zz_536_;
  wire                _zz_537_;
  wire                _zz_538_;
  wire                _zz_539_;
  wire                _zz_540_;
  wire                _zz_541_;
  wire                _zz_542_;
  wire                _zz_543_;
  wire                _zz_544_;
  wire                _zz_545_;
  wire                _zz_546_;
  wire                _zz_547_;
  wire                _zz_548_;
  wire                _zz_549_;
  wire                _zz_550_;
  wire                _zz_551_;
  wire                _zz_552_;
  wire                _zz_553_;
  wire                _zz_554_;
  wire                _zz_555_;
  wire                _zz_556_;
  wire                _zz_557_;
  wire                _zz_558_;
  wire                _zz_559_;
  wire                _zz_560_;
  wire                _zz_561_;
  wire                _zz_562_;
  wire                _zz_563_;
  wire                _zz_564_;
  wire                _zz_565_;
  wire       [31:0]   _zz_566_;
  wire       [15:0]   _zz_567_;
  wire       [15:0]   _zz_568_;
  wire       [5:0]    _zz_569_;
  wire       [63:0]   _zz_570_;
  wire                _zz_571_;
  wire                _zz_572_;
  wire                _zz_573_;
  wire                _zz_574_;
  wire                _zz_575_;
  wire                _zz_576_;
  wire                _zz_577_;
  wire                _zz_578_;
  wire                _zz_579_;
  wire                _zz_580_;
  wire                _zz_581_;
  wire                _zz_582_;
  wire                _zz_583_;
  wire                _zz_584_;
  wire                _zz_585_;
  wire                _zz_586_;
  wire                _zz_587_;
  wire                _zz_588_;
  wire                _zz_589_;
  wire                _zz_590_;
  wire                _zz_591_;
  wire                _zz_592_;
  wire                _zz_593_;
  wire                _zz_594_;
  wire                _zz_595_;
  wire                _zz_596_;
  wire                _zz_597_;
  wire                _zz_598_;
  wire                _zz_599_;
  wire                _zz_600_;
  wire                _zz_601_;
  wire                _zz_602_;
  wire                _zz_603_;
  wire                _zz_604_;
  wire                _zz_605_;
  wire                _zz_606_;
  wire                _zz_607_;
  wire                _zz_608_;
  wire                _zz_609_;
  wire                _zz_610_;
  wire                _zz_611_;
  wire                _zz_612_;
  wire                _zz_613_;
  wire                _zz_614_;
  wire                _zz_615_;
  wire                _zz_616_;
  wire                _zz_617_;
  wire                _zz_618_;
  wire                _zz_619_;
  wire                _zz_620_;
  wire                _zz_621_;
  wire                _zz_622_;
  wire                _zz_623_;
  wire                _zz_624_;
  wire                _zz_625_;
  wire                _zz_626_;
  wire                _zz_627_;
  wire                _zz_628_;
  wire                _zz_629_;
  wire                _zz_630_;
  wire                _zz_631_;
  wire                _zz_632_;
  wire                _zz_633_;
  wire                _zz_634_;
  wire       [31:0]   _zz_635_;
  wire       [15:0]   _zz_636_;
  wire       [15:0]   _zz_637_;
  wire       [5:0]    _zz_638_;
  wire       [63:0]   _zz_639_;
  wire                _zz_640_;
  wire                _zz_641_;
  wire                _zz_642_;
  wire                _zz_643_;
  wire                _zz_644_;
  wire                _zz_645_;
  wire                _zz_646_;
  wire                _zz_647_;
  wire                _zz_648_;
  wire                _zz_649_;
  wire                _zz_650_;
  wire                _zz_651_;
  wire                _zz_652_;
  wire                _zz_653_;
  wire                _zz_654_;
  wire                _zz_655_;
  wire                _zz_656_;
  wire                _zz_657_;
  wire                _zz_658_;
  wire                _zz_659_;
  wire                _zz_660_;
  wire                _zz_661_;
  wire                _zz_662_;
  wire                _zz_663_;
  wire                _zz_664_;
  wire                _zz_665_;
  wire                _zz_666_;
  wire                _zz_667_;
  wire                _zz_668_;
  wire                _zz_669_;
  wire                _zz_670_;
  wire                _zz_671_;
  wire                _zz_672_;
  wire                _zz_673_;
  wire                _zz_674_;
  wire                _zz_675_;
  wire                _zz_676_;
  wire                _zz_677_;
  wire                _zz_678_;
  wire                _zz_679_;
  wire                _zz_680_;
  wire                _zz_681_;
  wire                _zz_682_;
  wire                _zz_683_;
  wire                _zz_684_;
  wire                _zz_685_;
  wire                _zz_686_;
  wire                _zz_687_;
  wire                _zz_688_;
  wire                _zz_689_;
  wire                _zz_690_;
  wire                _zz_691_;
  wire                _zz_692_;
  wire                _zz_693_;
  wire                _zz_694_;
  wire                _zz_695_;
  wire                _zz_696_;
  wire                _zz_697_;
  wire                _zz_698_;
  wire                _zz_699_;
  wire                _zz_700_;
  wire                _zz_701_;
  wire                _zz_702_;
  wire                _zz_703_;
  wire       [31:0]   _zz_704_;
  wire       [15:0]   _zz_705_;
  wire       [15:0]   _zz_706_;
  wire       [5:0]    _zz_707_;
  wire       [63:0]   _zz_708_;
  wire                _zz_709_;
  wire                _zz_710_;
  wire                _zz_711_;
  wire                _zz_712_;
  wire                _zz_713_;
  wire                _zz_714_;
  wire                _zz_715_;
  wire                _zz_716_;
  wire                _zz_717_;
  wire                _zz_718_;
  wire                _zz_719_;
  wire                _zz_720_;
  wire                _zz_721_;
  wire                _zz_722_;
  wire                _zz_723_;
  wire                _zz_724_;
  wire                _zz_725_;
  wire                _zz_726_;
  wire                _zz_727_;
  wire                _zz_728_;
  wire                _zz_729_;
  wire                _zz_730_;
  wire                _zz_731_;
  wire                _zz_732_;
  wire                _zz_733_;
  wire                _zz_734_;
  wire                _zz_735_;
  wire                _zz_736_;
  wire                _zz_737_;
  wire                _zz_738_;
  wire                _zz_739_;
  wire                _zz_740_;
  wire                _zz_741_;
  wire                _zz_742_;
  wire                _zz_743_;
  wire                _zz_744_;
  wire                _zz_745_;
  wire                _zz_746_;
  wire                _zz_747_;
  wire                _zz_748_;
  wire                _zz_749_;
  wire                _zz_750_;
  wire                _zz_751_;
  wire                _zz_752_;
  wire                _zz_753_;
  wire                _zz_754_;
  wire                _zz_755_;
  wire                _zz_756_;
  wire                _zz_757_;
  wire                _zz_758_;
  wire                _zz_759_;
  wire                _zz_760_;
  wire                _zz_761_;
  wire                _zz_762_;
  wire                _zz_763_;
  wire                _zz_764_;
  wire                _zz_765_;
  wire                _zz_766_;
  wire                _zz_767_;
  wire                _zz_768_;
  wire                _zz_769_;
  wire                _zz_770_;
  wire                _zz_771_;
  wire                _zz_772_;
  wire       [31:0]   _zz_773_;
  wire       [15:0]   _zz_774_;
  wire       [15:0]   _zz_775_;
  wire       [5:0]    _zz_776_;
  wire       [63:0]   _zz_777_;
  wire                _zz_778_;
  wire                _zz_779_;
  wire                _zz_780_;
  wire                _zz_781_;
  wire                _zz_782_;
  wire                _zz_783_;
  wire                _zz_784_;
  wire                _zz_785_;
  wire                _zz_786_;
  wire                _zz_787_;
  wire                _zz_788_;
  wire                _zz_789_;
  wire                _zz_790_;
  wire                _zz_791_;
  wire                _zz_792_;
  wire                _zz_793_;
  wire                _zz_794_;
  wire                _zz_795_;
  wire                _zz_796_;
  wire                _zz_797_;
  wire                _zz_798_;
  wire                _zz_799_;
  wire                _zz_800_;
  wire                _zz_801_;
  wire                _zz_802_;
  wire                _zz_803_;
  wire                _zz_804_;
  wire                _zz_805_;
  wire                _zz_806_;
  wire                _zz_807_;
  wire                _zz_808_;
  wire                _zz_809_;
  wire                _zz_810_;
  wire                _zz_811_;
  wire                _zz_812_;
  wire                _zz_813_;
  wire                _zz_814_;
  wire                _zz_815_;
  wire                _zz_816_;
  wire                _zz_817_;
  wire                _zz_818_;
  wire                _zz_819_;
  wire                _zz_820_;
  wire                _zz_821_;
  wire                _zz_822_;
  wire                _zz_823_;
  wire                _zz_824_;
  wire                _zz_825_;
  wire                _zz_826_;
  wire                _zz_827_;
  wire                _zz_828_;
  wire                _zz_829_;
  wire                _zz_830_;
  wire                _zz_831_;
  wire                _zz_832_;
  wire                _zz_833_;
  wire                _zz_834_;
  wire                _zz_835_;
  wire                _zz_836_;
  wire                _zz_837_;
  wire                _zz_838_;
  wire                _zz_839_;
  wire                _zz_840_;
  wire                _zz_841_;
  wire       [31:0]   _zz_842_;
  wire       [15:0]   _zz_843_;
  wire       [15:0]   _zz_844_;
  wire       [5:0]    _zz_845_;
  wire       [63:0]   _zz_846_;
  wire                _zz_847_;
  wire                _zz_848_;
  wire                _zz_849_;
  wire                _zz_850_;
  wire                _zz_851_;
  wire                _zz_852_;
  wire                _zz_853_;
  wire                _zz_854_;
  wire                _zz_855_;
  wire                _zz_856_;
  wire                _zz_857_;
  wire                _zz_858_;
  wire                _zz_859_;
  wire                _zz_860_;
  wire                _zz_861_;
  wire                _zz_862_;
  wire                _zz_863_;
  wire                _zz_864_;
  wire                _zz_865_;
  wire                _zz_866_;
  wire                _zz_867_;
  wire                _zz_868_;
  wire                _zz_869_;
  wire                _zz_870_;
  wire                _zz_871_;
  wire                _zz_872_;
  wire                _zz_873_;
  wire                _zz_874_;
  wire                _zz_875_;
  wire                _zz_876_;
  wire                _zz_877_;
  wire                _zz_878_;
  wire                _zz_879_;
  wire                _zz_880_;
  wire                _zz_881_;
  wire                _zz_882_;
  wire                _zz_883_;
  wire                _zz_884_;
  wire                _zz_885_;
  wire                _zz_886_;
  wire                _zz_887_;
  wire                _zz_888_;
  wire                _zz_889_;
  wire                _zz_890_;
  wire                _zz_891_;
  wire                _zz_892_;
  wire                _zz_893_;
  wire                _zz_894_;
  wire                _zz_895_;
  wire                _zz_896_;
  wire                _zz_897_;
  wire                _zz_898_;
  wire                _zz_899_;
  wire                _zz_900_;
  wire                _zz_901_;
  wire                _zz_902_;
  wire                _zz_903_;
  wire                _zz_904_;
  wire                _zz_905_;
  wire                _zz_906_;
  wire                _zz_907_;
  wire                _zz_908_;
  wire                _zz_909_;
  wire                _zz_910_;
  wire       [31:0]   _zz_911_;
  wire       [15:0]   _zz_912_;
  wire       [15:0]   _zz_913_;
  wire       [5:0]    _zz_914_;
  wire       [63:0]   _zz_915_;
  wire                _zz_916_;
  wire                _zz_917_;
  wire                _zz_918_;
  wire                _zz_919_;
  wire                _zz_920_;
  wire                _zz_921_;
  wire                _zz_922_;
  wire                _zz_923_;
  wire                _zz_924_;
  wire                _zz_925_;
  wire                _zz_926_;
  wire                _zz_927_;
  wire                _zz_928_;
  wire                _zz_929_;
  wire                _zz_930_;
  wire                _zz_931_;
  wire                _zz_932_;
  wire                _zz_933_;
  wire                _zz_934_;
  wire                _zz_935_;
  wire                _zz_936_;
  wire                _zz_937_;
  wire                _zz_938_;
  wire                _zz_939_;
  wire                _zz_940_;
  wire                _zz_941_;
  wire                _zz_942_;
  wire                _zz_943_;
  wire                _zz_944_;
  wire                _zz_945_;
  wire                _zz_946_;
  wire                _zz_947_;
  wire                _zz_948_;
  wire                _zz_949_;
  wire                _zz_950_;
  wire                _zz_951_;
  wire                _zz_952_;
  wire                _zz_953_;
  wire                _zz_954_;
  wire                _zz_955_;
  wire                _zz_956_;
  wire                _zz_957_;
  wire                _zz_958_;
  wire                _zz_959_;
  wire                _zz_960_;
  wire                _zz_961_;
  wire                _zz_962_;
  wire                _zz_963_;
  wire                _zz_964_;
  wire                _zz_965_;
  wire                _zz_966_;
  wire                _zz_967_;
  wire                _zz_968_;
  wire                _zz_969_;
  wire                _zz_970_;
  wire                _zz_971_;
  wire                _zz_972_;
  wire                _zz_973_;
  wire                _zz_974_;
  wire                _zz_975_;
  wire                _zz_976_;
  wire                _zz_977_;
  wire                _zz_978_;
  wire                _zz_979_;
  wire       [31:0]   _zz_980_;
  wire       [15:0]   _zz_981_;
  wire       [15:0]   _zz_982_;
  wire       [5:0]    _zz_983_;
  wire       [63:0]   _zz_984_;
  wire                _zz_985_;
  wire                _zz_986_;
  wire                _zz_987_;
  wire                _zz_988_;
  wire                _zz_989_;
  wire                _zz_990_;
  wire                _zz_991_;
  wire                _zz_992_;
  wire                _zz_993_;
  wire                _zz_994_;
  wire                _zz_995_;
  wire                _zz_996_;
  wire                _zz_997_;
  wire                _zz_998_;
  wire                _zz_999_;
  wire                _zz_1000_;
  wire                _zz_1001_;
  wire                _zz_1002_;
  wire                _zz_1003_;
  wire                _zz_1004_;
  wire                _zz_1005_;
  wire                _zz_1006_;
  wire                _zz_1007_;
  wire                _zz_1008_;
  wire                _zz_1009_;
  wire                _zz_1010_;
  wire                _zz_1011_;
  wire                _zz_1012_;
  wire                _zz_1013_;
  wire                _zz_1014_;
  wire                _zz_1015_;
  wire                _zz_1016_;
  wire                _zz_1017_;
  wire                _zz_1018_;
  wire                _zz_1019_;
  wire                _zz_1020_;
  wire                _zz_1021_;
  wire                _zz_1022_;
  wire                _zz_1023_;
  wire                _zz_1024_;
  wire                _zz_1025_;
  wire                _zz_1026_;
  wire                _zz_1027_;
  wire                _zz_1028_;
  wire                _zz_1029_;
  wire                _zz_1030_;
  wire                _zz_1031_;
  wire                _zz_1032_;
  wire                _zz_1033_;
  wire                _zz_1034_;
  wire                _zz_1035_;
  wire                _zz_1036_;
  wire                _zz_1037_;
  wire                _zz_1038_;
  wire                _zz_1039_;
  wire                _zz_1040_;
  wire                _zz_1041_;
  wire                _zz_1042_;
  wire                _zz_1043_;
  wire                _zz_1044_;
  wire                _zz_1045_;
  wire                _zz_1046_;
  wire                _zz_1047_;
  wire                _zz_1048_;
  wire       [31:0]   _zz_1049_;
  wire       [15:0]   _zz_1050_;
  wire       [15:0]   _zz_1051_;
  wire       [5:0]    _zz_1052_;
  wire       [63:0]   _zz_1053_;
  wire                _zz_1054_;
  wire                _zz_1055_;
  wire                _zz_1056_;
  wire                _zz_1057_;
  wire                _zz_1058_;
  wire                _zz_1059_;
  wire                _zz_1060_;
  wire                _zz_1061_;
  wire                _zz_1062_;
  wire                _zz_1063_;
  wire                _zz_1064_;
  wire                _zz_1065_;
  wire                _zz_1066_;
  wire                _zz_1067_;
  wire                _zz_1068_;
  wire                _zz_1069_;
  wire                _zz_1070_;
  wire                _zz_1071_;
  wire                _zz_1072_;
  wire                _zz_1073_;
  wire                _zz_1074_;
  wire                _zz_1075_;
  wire                _zz_1076_;
  wire                _zz_1077_;
  wire                _zz_1078_;
  wire                _zz_1079_;
  wire                _zz_1080_;
  wire                _zz_1081_;
  wire                _zz_1082_;
  wire                _zz_1083_;
  wire                _zz_1084_;
  wire                _zz_1085_;
  wire                _zz_1086_;
  wire                _zz_1087_;
  wire                _zz_1088_;
  wire                _zz_1089_;
  wire                _zz_1090_;
  wire                _zz_1091_;
  wire                _zz_1092_;
  wire                _zz_1093_;
  wire                _zz_1094_;
  wire                _zz_1095_;
  wire                _zz_1096_;
  wire                _zz_1097_;
  wire                _zz_1098_;
  wire                _zz_1099_;
  wire                _zz_1100_;
  wire                _zz_1101_;
  wire                _zz_1102_;
  wire                _zz_1103_;
  wire                _zz_1104_;
  wire                _zz_1105_;
  wire                _zz_1106_;
  wire                _zz_1107_;
  wire                _zz_1108_;
  wire                _zz_1109_;
  wire                _zz_1110_;
  wire                _zz_1111_;
  wire                _zz_1112_;
  wire                _zz_1113_;
  wire                _zz_1114_;
  wire                _zz_1115_;
  wire                _zz_1116_;
  wire                _zz_1117_;
  wire       [31:0]   _zz_1118_;
  wire       [15:0]   _zz_1119_;
  wire       [15:0]   _zz_1120_;
  wire       [5:0]    _zz_1121_;
  wire       [63:0]   _zz_1122_;
  wire                _zz_1123_;
  wire                _zz_1124_;
  wire                _zz_1125_;
  wire                _zz_1126_;
  wire                _zz_1127_;
  wire                _zz_1128_;
  wire                _zz_1129_;
  wire                _zz_1130_;
  wire                _zz_1131_;
  wire                _zz_1132_;
  wire                _zz_1133_;
  wire                _zz_1134_;
  wire                _zz_1135_;
  wire                _zz_1136_;
  wire                _zz_1137_;
  wire                _zz_1138_;
  wire                _zz_1139_;
  wire                _zz_1140_;
  wire                _zz_1141_;
  wire                _zz_1142_;
  wire                _zz_1143_;
  wire                _zz_1144_;
  wire                _zz_1145_;
  wire                _zz_1146_;
  wire                _zz_1147_;
  wire                _zz_1148_;
  wire                _zz_1149_;
  wire                _zz_1150_;
  wire                _zz_1151_;
  wire                _zz_1152_;
  wire                _zz_1153_;
  wire                _zz_1154_;
  wire                _zz_1155_;
  wire                _zz_1156_;
  wire                _zz_1157_;
  wire                _zz_1158_;
  wire                _zz_1159_;
  wire                _zz_1160_;
  wire                _zz_1161_;
  wire                _zz_1162_;
  wire                _zz_1163_;
  wire                _zz_1164_;
  wire                _zz_1165_;
  wire                _zz_1166_;
  wire                _zz_1167_;
  wire                _zz_1168_;
  wire                _zz_1169_;
  wire                _zz_1170_;
  wire                _zz_1171_;
  wire                _zz_1172_;
  wire                _zz_1173_;
  wire                _zz_1174_;
  wire                _zz_1175_;
  wire                _zz_1176_;
  wire                _zz_1177_;
  wire                _zz_1178_;
  wire                _zz_1179_;
  wire                _zz_1180_;
  wire                _zz_1181_;
  wire                _zz_1182_;
  wire                _zz_1183_;
  wire                _zz_1184_;
  wire                _zz_1185_;
  wire                _zz_1186_;
  wire       [31:0]   _zz_1187_;
  wire       [15:0]   _zz_1188_;
  wire       [15:0]   _zz_1189_;
  wire       [5:0]    _zz_1190_;
  wire       [63:0]   _zz_1191_;
  wire                _zz_1192_;
  wire                _zz_1193_;
  wire                _zz_1194_;
  wire                _zz_1195_;
  wire                _zz_1196_;
  wire                _zz_1197_;
  wire                _zz_1198_;
  wire                _zz_1199_;
  wire                _zz_1200_;
  wire                _zz_1201_;
  wire                _zz_1202_;
  wire                _zz_1203_;
  wire                _zz_1204_;
  wire                _zz_1205_;
  wire                _zz_1206_;
  wire                _zz_1207_;
  wire                _zz_1208_;
  wire                _zz_1209_;
  wire                _zz_1210_;
  wire                _zz_1211_;
  wire                _zz_1212_;
  wire                _zz_1213_;
  wire                _zz_1214_;
  wire                _zz_1215_;
  wire                _zz_1216_;
  wire                _zz_1217_;
  wire                _zz_1218_;
  wire                _zz_1219_;
  wire                _zz_1220_;
  wire                _zz_1221_;
  wire                _zz_1222_;
  wire                _zz_1223_;
  wire                _zz_1224_;
  wire                _zz_1225_;
  wire                _zz_1226_;
  wire                _zz_1227_;
  wire                _zz_1228_;
  wire                _zz_1229_;
  wire                _zz_1230_;
  wire                _zz_1231_;
  wire                _zz_1232_;
  wire                _zz_1233_;
  wire                _zz_1234_;
  wire                _zz_1235_;
  wire                _zz_1236_;
  wire                _zz_1237_;
  wire                _zz_1238_;
  wire                _zz_1239_;
  wire                _zz_1240_;
  wire                _zz_1241_;
  wire                _zz_1242_;
  wire                _zz_1243_;
  wire                _zz_1244_;
  wire                _zz_1245_;
  wire                _zz_1246_;
  wire                _zz_1247_;
  wire                _zz_1248_;
  wire                _zz_1249_;
  wire                _zz_1250_;
  wire                _zz_1251_;
  wire                _zz_1252_;
  wire                _zz_1253_;
  wire                _zz_1254_;
  wire                _zz_1255_;
  wire       [31:0]   _zz_1256_;
  wire       [15:0]   _zz_1257_;
  wire       [15:0]   _zz_1258_;
  wire       [5:0]    _zz_1259_;
  wire       [63:0]   _zz_1260_;
  wire                _zz_1261_;
  wire                _zz_1262_;
  wire                _zz_1263_;
  wire                _zz_1264_;
  wire                _zz_1265_;
  wire                _zz_1266_;
  wire                _zz_1267_;
  wire                _zz_1268_;
  wire                _zz_1269_;
  wire                _zz_1270_;
  wire                _zz_1271_;
  wire                _zz_1272_;
  wire                _zz_1273_;
  wire                _zz_1274_;
  wire                _zz_1275_;
  wire                _zz_1276_;
  wire                _zz_1277_;
  wire                _zz_1278_;
  wire                _zz_1279_;
  wire                _zz_1280_;
  wire                _zz_1281_;
  wire                _zz_1282_;
  wire                _zz_1283_;
  wire                _zz_1284_;
  wire                _zz_1285_;
  wire                _zz_1286_;
  wire                _zz_1287_;
  wire                _zz_1288_;
  wire                _zz_1289_;
  wire                _zz_1290_;
  wire                _zz_1291_;
  wire                _zz_1292_;
  wire                _zz_1293_;
  wire                _zz_1294_;
  wire                _zz_1295_;
  wire                _zz_1296_;
  wire                _zz_1297_;
  wire                _zz_1298_;
  wire                _zz_1299_;
  wire                _zz_1300_;
  wire                _zz_1301_;
  wire                _zz_1302_;
  wire                _zz_1303_;
  wire                _zz_1304_;
  wire                _zz_1305_;
  wire                _zz_1306_;
  wire                _zz_1307_;
  wire                _zz_1308_;
  wire                _zz_1309_;
  wire                _zz_1310_;
  wire                _zz_1311_;
  wire                _zz_1312_;
  wire                _zz_1313_;
  wire                _zz_1314_;
  wire                _zz_1315_;
  wire                _zz_1316_;
  wire                _zz_1317_;
  wire                _zz_1318_;
  wire                _zz_1319_;
  wire                _zz_1320_;
  wire                _zz_1321_;
  wire                _zz_1322_;
  wire                _zz_1323_;
  wire                _zz_1324_;
  wire       [31:0]   _zz_1325_;
  wire       [15:0]   _zz_1326_;
  wire       [15:0]   _zz_1327_;
  wire       [5:0]    _zz_1328_;
  wire       [63:0]   _zz_1329_;
  wire                _zz_1330_;
  wire                _zz_1331_;
  wire                _zz_1332_;
  wire                _zz_1333_;
  wire                _zz_1334_;
  wire                _zz_1335_;
  wire                _zz_1336_;
  wire                _zz_1337_;
  wire                _zz_1338_;
  wire                _zz_1339_;
  wire                _zz_1340_;
  wire                _zz_1341_;
  wire                _zz_1342_;
  wire                _zz_1343_;
  wire                _zz_1344_;
  wire                _zz_1345_;
  wire                _zz_1346_;
  wire                _zz_1347_;
  wire                _zz_1348_;
  wire                _zz_1349_;
  wire                _zz_1350_;
  wire                _zz_1351_;
  wire                _zz_1352_;
  wire                _zz_1353_;
  wire                _zz_1354_;
  wire                _zz_1355_;
  wire                _zz_1356_;
  wire                _zz_1357_;
  wire                _zz_1358_;
  wire                _zz_1359_;
  wire                _zz_1360_;
  wire                _zz_1361_;
  wire                _zz_1362_;
  wire                _zz_1363_;
  wire                _zz_1364_;
  wire                _zz_1365_;
  wire                _zz_1366_;
  wire                _zz_1367_;
  wire                _zz_1368_;
  wire                _zz_1369_;
  wire                _zz_1370_;
  wire                _zz_1371_;
  wire                _zz_1372_;
  wire                _zz_1373_;
  wire                _zz_1374_;
  wire                _zz_1375_;
  wire                _zz_1376_;
  wire                _zz_1377_;
  wire                _zz_1378_;
  wire                _zz_1379_;
  wire                _zz_1380_;
  wire                _zz_1381_;
  wire                _zz_1382_;
  wire                _zz_1383_;
  wire                _zz_1384_;
  wire                _zz_1385_;
  wire                _zz_1386_;
  wire                _zz_1387_;
  wire                _zz_1388_;
  wire                _zz_1389_;
  wire                _zz_1390_;
  wire                _zz_1391_;
  wire                _zz_1392_;
  wire                _zz_1393_;
  wire       [31:0]   _zz_1394_;
  wire       [15:0]   _zz_1395_;
  wire       [15:0]   _zz_1396_;
  wire       [5:0]    _zz_1397_;
  wire       [63:0]   _zz_1398_;
  wire                _zz_1399_;
  wire                _zz_1400_;
  wire                _zz_1401_;
  wire                _zz_1402_;
  wire                _zz_1403_;
  wire                _zz_1404_;
  wire                _zz_1405_;
  wire                _zz_1406_;
  wire                _zz_1407_;
  wire                _zz_1408_;
  wire                _zz_1409_;
  wire                _zz_1410_;
  wire                _zz_1411_;
  wire                _zz_1412_;
  wire                _zz_1413_;
  wire                _zz_1414_;
  wire                _zz_1415_;
  wire                _zz_1416_;
  wire                _zz_1417_;
  wire                _zz_1418_;
  wire                _zz_1419_;
  wire                _zz_1420_;
  wire                _zz_1421_;
  wire                _zz_1422_;
  wire                _zz_1423_;
  wire                _zz_1424_;
  wire                _zz_1425_;
  wire                _zz_1426_;
  wire                _zz_1427_;
  wire                _zz_1428_;
  wire                _zz_1429_;
  wire                _zz_1430_;
  wire                _zz_1431_;
  wire                _zz_1432_;
  wire                _zz_1433_;
  wire                _zz_1434_;
  wire                _zz_1435_;
  wire                _zz_1436_;
  wire                _zz_1437_;
  wire                _zz_1438_;
  wire                _zz_1439_;
  wire                _zz_1440_;
  wire                _zz_1441_;
  wire                _zz_1442_;
  wire                _zz_1443_;
  wire                _zz_1444_;
  wire                _zz_1445_;
  wire                _zz_1446_;
  wire                _zz_1447_;
  wire                _zz_1448_;
  wire                _zz_1449_;
  wire                _zz_1450_;
  wire                _zz_1451_;
  wire                _zz_1452_;
  wire                _zz_1453_;
  wire                _zz_1454_;
  wire                _zz_1455_;
  wire                _zz_1456_;
  wire                _zz_1457_;
  wire                _zz_1458_;
  wire                _zz_1459_;
  wire                _zz_1460_;
  wire                _zz_1461_;
  wire                _zz_1462_;
  wire       [31:0]   _zz_1463_;
  wire       [15:0]   _zz_1464_;
  wire       [15:0]   _zz_1465_;
  wire       [5:0]    _zz_1466_;
  wire       [63:0]   _zz_1467_;
  wire                _zz_1468_;
  wire                _zz_1469_;
  wire                _zz_1470_;
  wire                _zz_1471_;
  wire                _zz_1472_;
  wire                _zz_1473_;
  wire                _zz_1474_;
  wire                _zz_1475_;
  wire                _zz_1476_;
  wire                _zz_1477_;
  wire                _zz_1478_;
  wire                _zz_1479_;
  wire                _zz_1480_;
  wire                _zz_1481_;
  wire                _zz_1482_;
  wire                _zz_1483_;
  wire                _zz_1484_;
  wire                _zz_1485_;
  wire                _zz_1486_;
  wire                _zz_1487_;
  wire                _zz_1488_;
  wire                _zz_1489_;
  wire                _zz_1490_;
  wire                _zz_1491_;
  wire                _zz_1492_;
  wire                _zz_1493_;
  wire                _zz_1494_;
  wire                _zz_1495_;
  wire                _zz_1496_;
  wire                _zz_1497_;
  wire                _zz_1498_;
  wire                _zz_1499_;
  wire                _zz_1500_;
  wire                _zz_1501_;
  wire                _zz_1502_;
  wire                _zz_1503_;
  wire                _zz_1504_;
  wire                _zz_1505_;
  wire                _zz_1506_;
  wire                _zz_1507_;
  wire                _zz_1508_;
  wire                _zz_1509_;
  wire                _zz_1510_;
  wire                _zz_1511_;
  wire                _zz_1512_;
  wire                _zz_1513_;
  wire                _zz_1514_;
  wire                _zz_1515_;
  wire                _zz_1516_;
  wire                _zz_1517_;
  wire                _zz_1518_;
  wire                _zz_1519_;
  wire                _zz_1520_;
  wire                _zz_1521_;
  wire                _zz_1522_;
  wire                _zz_1523_;
  wire                _zz_1524_;
  wire                _zz_1525_;
  wire                _zz_1526_;
  wire                _zz_1527_;
  wire                _zz_1528_;
  wire                _zz_1529_;
  wire                _zz_1530_;
  wire                _zz_1531_;
  wire       [31:0]   _zz_1532_;
  wire       [15:0]   _zz_1533_;
  wire       [15:0]   _zz_1534_;
  wire       [5:0]    _zz_1535_;
  wire       [63:0]   _zz_1536_;
  wire                _zz_1537_;
  wire                _zz_1538_;
  wire                _zz_1539_;
  wire                _zz_1540_;
  wire                _zz_1541_;
  wire                _zz_1542_;
  wire                _zz_1543_;
  wire                _zz_1544_;
  wire                _zz_1545_;
  wire                _zz_1546_;
  wire                _zz_1547_;
  wire                _zz_1548_;
  wire                _zz_1549_;
  wire                _zz_1550_;
  wire                _zz_1551_;
  wire                _zz_1552_;
  wire                _zz_1553_;
  wire                _zz_1554_;
  wire                _zz_1555_;
  wire                _zz_1556_;
  wire                _zz_1557_;
  wire                _zz_1558_;
  wire                _zz_1559_;
  wire                _zz_1560_;
  wire                _zz_1561_;
  wire                _zz_1562_;
  wire                _zz_1563_;
  wire                _zz_1564_;
  wire                _zz_1565_;
  wire                _zz_1566_;
  wire                _zz_1567_;
  wire                _zz_1568_;
  wire                _zz_1569_;
  wire                _zz_1570_;
  wire                _zz_1571_;
  wire                _zz_1572_;
  wire                _zz_1573_;
  wire                _zz_1574_;
  wire                _zz_1575_;
  wire                _zz_1576_;
  wire                _zz_1577_;
  wire                _zz_1578_;
  wire                _zz_1579_;
  wire                _zz_1580_;
  wire                _zz_1581_;
  wire                _zz_1582_;
  wire                _zz_1583_;
  wire                _zz_1584_;
  wire                _zz_1585_;
  wire                _zz_1586_;
  wire                _zz_1587_;
  wire                _zz_1588_;
  wire                _zz_1589_;
  wire                _zz_1590_;
  wire                _zz_1591_;
  wire                _zz_1592_;
  wire                _zz_1593_;
  wire                _zz_1594_;
  wire                _zz_1595_;
  wire                _zz_1596_;
  wire                _zz_1597_;
  wire                _zz_1598_;
  wire                _zz_1599_;
  wire                _zz_1600_;
  wire       [31:0]   _zz_1601_;
  wire       [15:0]   _zz_1602_;
  wire       [15:0]   _zz_1603_;
  wire       [5:0]    _zz_1604_;
  wire       [63:0]   _zz_1605_;
  wire                _zz_1606_;
  wire                _zz_1607_;
  wire                _zz_1608_;
  wire                _zz_1609_;
  wire                _zz_1610_;
  wire                _zz_1611_;
  wire                _zz_1612_;
  wire                _zz_1613_;
  wire                _zz_1614_;
  wire                _zz_1615_;
  wire                _zz_1616_;
  wire                _zz_1617_;
  wire                _zz_1618_;
  wire                _zz_1619_;
  wire                _zz_1620_;
  wire                _zz_1621_;
  wire                _zz_1622_;
  wire                _zz_1623_;
  wire                _zz_1624_;
  wire                _zz_1625_;
  wire                _zz_1626_;
  wire                _zz_1627_;
  wire                _zz_1628_;
  wire                _zz_1629_;
  wire                _zz_1630_;
  wire                _zz_1631_;
  wire                _zz_1632_;
  wire                _zz_1633_;
  wire                _zz_1634_;
  wire                _zz_1635_;
  wire                _zz_1636_;
  wire                _zz_1637_;
  wire                _zz_1638_;
  wire                _zz_1639_;
  wire                _zz_1640_;
  wire                _zz_1641_;
  wire                _zz_1642_;
  wire                _zz_1643_;
  wire                _zz_1644_;
  wire                _zz_1645_;
  wire                _zz_1646_;
  wire                _zz_1647_;
  wire                _zz_1648_;
  wire                _zz_1649_;
  wire                _zz_1650_;
  wire                _zz_1651_;
  wire                _zz_1652_;
  wire                _zz_1653_;
  wire                _zz_1654_;
  wire                _zz_1655_;
  wire                _zz_1656_;
  wire                _zz_1657_;
  wire                _zz_1658_;
  wire                _zz_1659_;
  wire                _zz_1660_;
  wire                _zz_1661_;
  wire                _zz_1662_;
  wire                _zz_1663_;
  wire                _zz_1664_;
  wire                _zz_1665_;
  wire                _zz_1666_;
  wire                _zz_1667_;
  wire                _zz_1668_;
  wire                _zz_1669_;
  wire       [31:0]   _zz_1670_;
  wire       [15:0]   _zz_1671_;
  wire       [15:0]   _zz_1672_;
  wire       [5:0]    _zz_1673_;
  wire       [63:0]   _zz_1674_;
  wire                _zz_1675_;
  wire                _zz_1676_;
  wire                _zz_1677_;
  wire                _zz_1678_;
  wire                _zz_1679_;
  wire                _zz_1680_;
  wire                _zz_1681_;
  wire                _zz_1682_;
  wire                _zz_1683_;
  wire                _zz_1684_;
  wire                _zz_1685_;
  wire                _zz_1686_;
  wire                _zz_1687_;
  wire                _zz_1688_;
  wire                _zz_1689_;
  wire                _zz_1690_;
  wire                _zz_1691_;
  wire                _zz_1692_;
  wire                _zz_1693_;
  wire                _zz_1694_;
  wire                _zz_1695_;
  wire                _zz_1696_;
  wire                _zz_1697_;
  wire                _zz_1698_;
  wire                _zz_1699_;
  wire                _zz_1700_;
  wire                _zz_1701_;
  wire                _zz_1702_;
  wire                _zz_1703_;
  wire                _zz_1704_;
  wire                _zz_1705_;
  wire                _zz_1706_;
  wire                _zz_1707_;
  wire                _zz_1708_;
  wire                _zz_1709_;
  wire                _zz_1710_;
  wire                _zz_1711_;
  wire                _zz_1712_;
  wire                _zz_1713_;
  wire                _zz_1714_;
  wire                _zz_1715_;
  wire                _zz_1716_;
  wire                _zz_1717_;
  wire                _zz_1718_;
  wire                _zz_1719_;
  wire                _zz_1720_;
  wire                _zz_1721_;
  wire                _zz_1722_;
  wire                _zz_1723_;
  wire                _zz_1724_;
  wire                _zz_1725_;
  wire                _zz_1726_;
  wire                _zz_1727_;
  wire                _zz_1728_;
  wire                _zz_1729_;
  wire                _zz_1730_;
  wire                _zz_1731_;
  wire                _zz_1732_;
  wire                _zz_1733_;
  wire                _zz_1734_;
  wire                _zz_1735_;
  wire                _zz_1736_;
  wire                _zz_1737_;
  wire                _zz_1738_;
  wire       [31:0]   _zz_1739_;
  wire       [15:0]   _zz_1740_;
  wire       [15:0]   _zz_1741_;
  wire       [5:0]    _zz_1742_;
  wire       [63:0]   _zz_1743_;
  wire                _zz_1744_;
  wire                _zz_1745_;
  wire                _zz_1746_;
  wire                _zz_1747_;
  wire                _zz_1748_;
  wire                _zz_1749_;
  wire                _zz_1750_;
  wire                _zz_1751_;
  wire                _zz_1752_;
  wire                _zz_1753_;
  wire                _zz_1754_;
  wire                _zz_1755_;
  wire                _zz_1756_;
  wire                _zz_1757_;
  wire                _zz_1758_;
  wire                _zz_1759_;
  wire                _zz_1760_;
  wire                _zz_1761_;
  wire                _zz_1762_;
  wire                _zz_1763_;
  wire                _zz_1764_;
  wire                _zz_1765_;
  wire                _zz_1766_;
  wire                _zz_1767_;
  wire                _zz_1768_;
  wire                _zz_1769_;
  wire                _zz_1770_;
  wire                _zz_1771_;
  wire                _zz_1772_;
  wire                _zz_1773_;
  wire                _zz_1774_;
  wire                _zz_1775_;
  wire                _zz_1776_;
  wire                _zz_1777_;
  wire                _zz_1778_;
  wire                _zz_1779_;
  wire                _zz_1780_;
  wire                _zz_1781_;
  wire                _zz_1782_;
  wire                _zz_1783_;
  wire                _zz_1784_;
  wire                _zz_1785_;
  wire                _zz_1786_;
  wire                _zz_1787_;
  wire                _zz_1788_;
  wire                _zz_1789_;
  wire                _zz_1790_;
  wire                _zz_1791_;
  wire                _zz_1792_;
  wire                _zz_1793_;
  wire                _zz_1794_;
  wire                _zz_1795_;
  wire                _zz_1796_;
  wire                _zz_1797_;
  wire                _zz_1798_;
  wire                _zz_1799_;
  wire                _zz_1800_;
  wire                _zz_1801_;
  wire                _zz_1802_;
  wire                _zz_1803_;
  wire                _zz_1804_;
  wire                _zz_1805_;
  wire                _zz_1806_;
  wire                _zz_1807_;
  wire       [31:0]   _zz_1808_;
  wire       [15:0]   _zz_1809_;
  wire       [15:0]   _zz_1810_;
  wire       [5:0]    _zz_1811_;
  wire       [63:0]   _zz_1812_;
  wire                _zz_1813_;
  wire                _zz_1814_;
  wire                _zz_1815_;
  wire                _zz_1816_;
  wire                _zz_1817_;
  wire                _zz_1818_;
  wire                _zz_1819_;
  wire                _zz_1820_;
  wire                _zz_1821_;
  wire                _zz_1822_;
  wire                _zz_1823_;
  wire                _zz_1824_;
  wire                _zz_1825_;
  wire                _zz_1826_;
  wire                _zz_1827_;
  wire                _zz_1828_;
  wire                _zz_1829_;
  wire                _zz_1830_;
  wire                _zz_1831_;
  wire                _zz_1832_;
  wire                _zz_1833_;
  wire                _zz_1834_;
  wire                _zz_1835_;
  wire                _zz_1836_;
  wire                _zz_1837_;
  wire                _zz_1838_;
  wire                _zz_1839_;
  wire                _zz_1840_;
  wire                _zz_1841_;
  wire                _zz_1842_;
  wire                _zz_1843_;
  wire                _zz_1844_;
  wire                _zz_1845_;
  wire                _zz_1846_;
  wire                _zz_1847_;
  wire                _zz_1848_;
  wire                _zz_1849_;
  wire                _zz_1850_;
  wire                _zz_1851_;
  wire                _zz_1852_;
  wire                _zz_1853_;
  wire                _zz_1854_;
  wire                _zz_1855_;
  wire                _zz_1856_;
  wire                _zz_1857_;
  wire                _zz_1858_;
  wire                _zz_1859_;
  wire                _zz_1860_;
  wire                _zz_1861_;
  wire                _zz_1862_;
  wire                _zz_1863_;
  wire                _zz_1864_;
  wire                _zz_1865_;
  wire                _zz_1866_;
  wire                _zz_1867_;
  wire                _zz_1868_;
  wire                _zz_1869_;
  wire                _zz_1870_;
  wire                _zz_1871_;
  wire                _zz_1872_;
  wire                _zz_1873_;
  wire                _zz_1874_;
  wire                _zz_1875_;
  wire                _zz_1876_;
  wire       [31:0]   _zz_1877_;
  wire       [15:0]   _zz_1878_;
  wire       [15:0]   _zz_1879_;
  wire       [5:0]    _zz_1880_;
  wire       [63:0]   _zz_1881_;
  wire                _zz_1882_;
  wire                _zz_1883_;
  wire                _zz_1884_;
  wire                _zz_1885_;
  wire                _zz_1886_;
  wire                _zz_1887_;
  wire                _zz_1888_;
  wire                _zz_1889_;
  wire                _zz_1890_;
  wire                _zz_1891_;
  wire                _zz_1892_;
  wire                _zz_1893_;
  wire                _zz_1894_;
  wire                _zz_1895_;
  wire                _zz_1896_;
  wire                _zz_1897_;
  wire                _zz_1898_;
  wire                _zz_1899_;
  wire                _zz_1900_;
  wire                _zz_1901_;
  wire                _zz_1902_;
  wire                _zz_1903_;
  wire                _zz_1904_;
  wire                _zz_1905_;
  wire                _zz_1906_;
  wire                _zz_1907_;
  wire                _zz_1908_;
  wire                _zz_1909_;
  wire                _zz_1910_;
  wire                _zz_1911_;
  wire                _zz_1912_;
  wire                _zz_1913_;
  wire                _zz_1914_;
  wire                _zz_1915_;
  wire                _zz_1916_;
  wire                _zz_1917_;
  wire                _zz_1918_;
  wire                _zz_1919_;
  wire                _zz_1920_;
  wire                _zz_1921_;
  wire                _zz_1922_;
  wire                _zz_1923_;
  wire                _zz_1924_;
  wire                _zz_1925_;
  wire                _zz_1926_;
  wire                _zz_1927_;
  wire                _zz_1928_;
  wire                _zz_1929_;
  wire                _zz_1930_;
  wire                _zz_1931_;
  wire                _zz_1932_;
  wire                _zz_1933_;
  wire                _zz_1934_;
  wire                _zz_1935_;
  wire                _zz_1936_;
  wire                _zz_1937_;
  wire                _zz_1938_;
  wire                _zz_1939_;
  wire                _zz_1940_;
  wire                _zz_1941_;
  wire                _zz_1942_;
  wire                _zz_1943_;
  wire                _zz_1944_;
  wire                _zz_1945_;
  wire       [31:0]   _zz_1946_;
  wire       [15:0]   _zz_1947_;
  wire       [15:0]   _zz_1948_;
  wire       [5:0]    _zz_1949_;
  wire       [63:0]   _zz_1950_;
  wire                _zz_1951_;
  wire                _zz_1952_;
  wire                _zz_1953_;
  wire                _zz_1954_;
  wire                _zz_1955_;
  wire                _zz_1956_;
  wire                _zz_1957_;
  wire                _zz_1958_;
  wire                _zz_1959_;
  wire                _zz_1960_;
  wire                _zz_1961_;
  wire                _zz_1962_;
  wire                _zz_1963_;
  wire                _zz_1964_;
  wire                _zz_1965_;
  wire                _zz_1966_;
  wire                _zz_1967_;
  wire                _zz_1968_;
  wire                _zz_1969_;
  wire                _zz_1970_;
  wire                _zz_1971_;
  wire                _zz_1972_;
  wire                _zz_1973_;
  wire                _zz_1974_;
  wire                _zz_1975_;
  wire                _zz_1976_;
  wire                _zz_1977_;
  wire                _zz_1978_;
  wire                _zz_1979_;
  wire                _zz_1980_;
  wire                _zz_1981_;
  wire                _zz_1982_;
  wire                _zz_1983_;
  wire                _zz_1984_;
  wire                _zz_1985_;
  wire                _zz_1986_;
  wire                _zz_1987_;
  wire                _zz_1988_;
  wire                _zz_1989_;
  wire                _zz_1990_;
  wire                _zz_1991_;
  wire                _zz_1992_;
  wire                _zz_1993_;
  wire                _zz_1994_;
  wire                _zz_1995_;
  wire                _zz_1996_;
  wire                _zz_1997_;
  wire                _zz_1998_;
  wire                _zz_1999_;
  wire                _zz_2000_;
  wire                _zz_2001_;
  wire                _zz_2002_;
  wire                _zz_2003_;
  wire                _zz_2004_;
  wire                _zz_2005_;
  wire                _zz_2006_;
  wire                _zz_2007_;
  wire                _zz_2008_;
  wire                _zz_2009_;
  wire                _zz_2010_;
  wire                _zz_2011_;
  wire                _zz_2012_;
  wire                _zz_2013_;
  wire                _zz_2014_;
  wire       [31:0]   _zz_2015_;
  wire       [15:0]   _zz_2016_;
  wire       [15:0]   _zz_2017_;
  wire       [5:0]    _zz_2018_;
  wire       [63:0]   _zz_2019_;
  wire                _zz_2020_;
  wire                _zz_2021_;
  wire                _zz_2022_;
  wire                _zz_2023_;
  wire                _zz_2024_;
  wire                _zz_2025_;
  wire                _zz_2026_;
  wire                _zz_2027_;
  wire                _zz_2028_;
  wire                _zz_2029_;
  wire                _zz_2030_;
  wire                _zz_2031_;
  wire                _zz_2032_;
  wire                _zz_2033_;
  wire                _zz_2034_;
  wire                _zz_2035_;
  wire                _zz_2036_;
  wire                _zz_2037_;
  wire                _zz_2038_;
  wire                _zz_2039_;
  wire                _zz_2040_;
  wire                _zz_2041_;
  wire                _zz_2042_;
  wire                _zz_2043_;
  wire                _zz_2044_;
  wire                _zz_2045_;
  wire                _zz_2046_;
  wire                _zz_2047_;
  wire                _zz_2048_;
  wire                _zz_2049_;
  wire                _zz_2050_;
  wire                _zz_2051_;
  wire                _zz_2052_;
  wire                _zz_2053_;
  wire                _zz_2054_;
  wire                _zz_2055_;
  wire                _zz_2056_;
  wire                _zz_2057_;
  wire                _zz_2058_;
  wire                _zz_2059_;
  wire                _zz_2060_;
  wire                _zz_2061_;
  wire                _zz_2062_;
  wire                _zz_2063_;
  wire                _zz_2064_;
  wire                _zz_2065_;
  wire                _zz_2066_;
  wire                _zz_2067_;
  wire                _zz_2068_;
  wire                _zz_2069_;
  wire                _zz_2070_;
  wire                _zz_2071_;
  wire                _zz_2072_;
  wire                _zz_2073_;
  wire                _zz_2074_;
  wire                _zz_2075_;
  wire                _zz_2076_;
  wire                _zz_2077_;
  wire                _zz_2078_;
  wire                _zz_2079_;
  wire                _zz_2080_;
  wire                _zz_2081_;
  wire                _zz_2082_;
  wire                _zz_2083_;
  wire       [31:0]   _zz_2084_;
  wire       [15:0]   _zz_2085_;
  wire       [15:0]   _zz_2086_;
  wire       [5:0]    _zz_2087_;
  wire       [63:0]   _zz_2088_;
  wire                _zz_2089_;
  wire                _zz_2090_;
  wire                _zz_2091_;
  wire                _zz_2092_;
  wire                _zz_2093_;
  wire                _zz_2094_;
  wire                _zz_2095_;
  wire                _zz_2096_;
  wire                _zz_2097_;
  wire                _zz_2098_;
  wire                _zz_2099_;
  wire                _zz_2100_;
  wire                _zz_2101_;
  wire                _zz_2102_;
  wire                _zz_2103_;
  wire                _zz_2104_;
  wire                _zz_2105_;
  wire                _zz_2106_;
  wire                _zz_2107_;
  wire                _zz_2108_;
  wire                _zz_2109_;
  wire                _zz_2110_;
  wire                _zz_2111_;
  wire                _zz_2112_;
  wire                _zz_2113_;
  wire                _zz_2114_;
  wire                _zz_2115_;
  wire                _zz_2116_;
  wire                _zz_2117_;
  wire                _zz_2118_;
  wire                _zz_2119_;
  wire                _zz_2120_;
  wire                _zz_2121_;
  wire                _zz_2122_;
  wire                _zz_2123_;
  wire                _zz_2124_;
  wire                _zz_2125_;
  wire                _zz_2126_;
  wire                _zz_2127_;
  wire                _zz_2128_;
  wire                _zz_2129_;
  wire                _zz_2130_;
  wire                _zz_2131_;
  wire                _zz_2132_;
  wire                _zz_2133_;
  wire                _zz_2134_;
  wire                _zz_2135_;
  wire                _zz_2136_;
  wire                _zz_2137_;
  wire                _zz_2138_;
  wire                _zz_2139_;
  wire                _zz_2140_;
  wire                _zz_2141_;
  wire                _zz_2142_;
  wire                _zz_2143_;
  wire                _zz_2144_;
  wire                _zz_2145_;
  wire                _zz_2146_;
  wire                _zz_2147_;
  wire                _zz_2148_;
  wire                _zz_2149_;
  wire                _zz_2150_;
  wire                _zz_2151_;
  wire                _zz_2152_;
  wire       [31:0]   _zz_2153_;
  wire       [15:0]   _zz_2154_;
  wire       [15:0]   _zz_2155_;
  wire       [5:0]    _zz_2156_;
  wire       [63:0]   _zz_2157_;
  wire                _zz_2158_;
  wire                _zz_2159_;
  wire                _zz_2160_;
  wire                _zz_2161_;
  wire                _zz_2162_;
  wire                _zz_2163_;
  wire                _zz_2164_;
  wire                _zz_2165_;
  wire                _zz_2166_;
  wire                _zz_2167_;
  wire                _zz_2168_;
  wire                _zz_2169_;
  wire                _zz_2170_;
  wire                _zz_2171_;
  wire                _zz_2172_;
  wire                _zz_2173_;
  wire                _zz_2174_;
  wire                _zz_2175_;
  wire                _zz_2176_;
  wire                _zz_2177_;
  wire                _zz_2178_;
  wire                _zz_2179_;
  wire                _zz_2180_;
  wire                _zz_2181_;
  wire                _zz_2182_;
  wire                _zz_2183_;
  wire                _zz_2184_;
  wire                _zz_2185_;
  wire                _zz_2186_;
  wire                _zz_2187_;
  wire                _zz_2188_;
  wire                _zz_2189_;
  wire                _zz_2190_;
  wire                _zz_2191_;
  wire                _zz_2192_;
  wire                _zz_2193_;
  wire                _zz_2194_;
  wire                _zz_2195_;
  wire                _zz_2196_;
  wire                _zz_2197_;
  wire                _zz_2198_;
  wire                _zz_2199_;
  wire                _zz_2200_;
  wire                _zz_2201_;
  wire                _zz_2202_;
  wire                _zz_2203_;
  wire                _zz_2204_;
  wire                _zz_2205_;
  wire                _zz_2206_;
  wire                _zz_2207_;
  wire                _zz_2208_;
  wire                _zz_2209_;
  wire                _zz_2210_;
  wire                _zz_2211_;
  wire                _zz_2212_;
  wire                _zz_2213_;
  wire                _zz_2214_;
  wire                _zz_2215_;
  wire                _zz_2216_;
  wire                _zz_2217_;
  wire                _zz_2218_;
  wire                _zz_2219_;
  wire                _zz_2220_;
  wire                _zz_2221_;
  wire       [31:0]   _zz_2222_;
  wire       [15:0]   _zz_2223_;
  wire       [15:0]   _zz_2224_;
  wire       [5:0]    _zz_2225_;
  wire       [63:0]   _zz_2226_;
  wire                _zz_2227_;
  wire                _zz_2228_;
  wire                _zz_2229_;
  wire                _zz_2230_;
  wire                _zz_2231_;
  wire                _zz_2232_;
  wire                _zz_2233_;
  wire                _zz_2234_;
  wire                _zz_2235_;
  wire                _zz_2236_;
  wire                _zz_2237_;
  wire                _zz_2238_;
  wire                _zz_2239_;
  wire                _zz_2240_;
  wire                _zz_2241_;
  wire                _zz_2242_;
  wire                _zz_2243_;
  wire                _zz_2244_;
  wire                _zz_2245_;
  wire                _zz_2246_;
  wire                _zz_2247_;
  wire                _zz_2248_;
  wire                _zz_2249_;
  wire                _zz_2250_;
  wire                _zz_2251_;
  wire                _zz_2252_;
  wire                _zz_2253_;
  wire                _zz_2254_;
  wire                _zz_2255_;
  wire                _zz_2256_;
  wire                _zz_2257_;
  wire                _zz_2258_;
  wire                _zz_2259_;
  wire                _zz_2260_;
  wire                _zz_2261_;
  wire                _zz_2262_;
  wire                _zz_2263_;
  wire                _zz_2264_;
  wire                _zz_2265_;
  wire                _zz_2266_;
  wire                _zz_2267_;
  wire                _zz_2268_;
  wire                _zz_2269_;
  wire                _zz_2270_;
  wire                _zz_2271_;
  wire                _zz_2272_;
  wire                _zz_2273_;
  wire                _zz_2274_;
  wire                _zz_2275_;
  wire                _zz_2276_;
  wire                _zz_2277_;
  wire                _zz_2278_;
  wire                _zz_2279_;
  wire                _zz_2280_;
  wire                _zz_2281_;
  wire                _zz_2282_;
  wire                _zz_2283_;
  wire                _zz_2284_;
  wire                _zz_2285_;
  wire                _zz_2286_;
  wire                _zz_2287_;
  wire                _zz_2288_;
  wire                _zz_2289_;
  wire                _zz_2290_;
  wire       [31:0]   _zz_2291_;
  wire       [15:0]   _zz_2292_;
  wire       [15:0]   _zz_2293_;
  wire       [5:0]    _zz_2294_;
  wire       [63:0]   _zz_2295_;
  wire                _zz_2296_;
  wire                _zz_2297_;
  wire                _zz_2298_;
  wire                _zz_2299_;
  wire                _zz_2300_;
  wire                _zz_2301_;
  wire                _zz_2302_;
  wire                _zz_2303_;
  wire                _zz_2304_;
  wire                _zz_2305_;
  wire                _zz_2306_;
  wire                _zz_2307_;
  wire                _zz_2308_;
  wire                _zz_2309_;
  wire                _zz_2310_;
  wire                _zz_2311_;
  wire                _zz_2312_;
  wire                _zz_2313_;
  wire                _zz_2314_;
  wire                _zz_2315_;
  wire                _zz_2316_;
  wire                _zz_2317_;
  wire                _zz_2318_;
  wire                _zz_2319_;
  wire                _zz_2320_;
  wire                _zz_2321_;
  wire                _zz_2322_;
  wire                _zz_2323_;
  wire                _zz_2324_;
  wire                _zz_2325_;
  wire                _zz_2326_;
  wire                _zz_2327_;
  wire                _zz_2328_;
  wire                _zz_2329_;
  wire                _zz_2330_;
  wire                _zz_2331_;
  wire                _zz_2332_;
  wire                _zz_2333_;
  wire                _zz_2334_;
  wire                _zz_2335_;
  wire                _zz_2336_;
  wire                _zz_2337_;
  wire                _zz_2338_;
  wire                _zz_2339_;
  wire                _zz_2340_;
  wire                _zz_2341_;
  wire                _zz_2342_;
  wire                _zz_2343_;
  wire                _zz_2344_;
  wire                _zz_2345_;
  wire                _zz_2346_;
  wire                _zz_2347_;
  wire                _zz_2348_;
  wire                _zz_2349_;
  wire                _zz_2350_;
  wire                _zz_2351_;
  wire                _zz_2352_;
  wire                _zz_2353_;
  wire                _zz_2354_;
  wire                _zz_2355_;
  wire                _zz_2356_;
  wire                _zz_2357_;
  wire                _zz_2358_;
  wire                _zz_2359_;
  wire       [31:0]   _zz_2360_;
  wire       [15:0]   _zz_2361_;
  wire       [15:0]   _zz_2362_;
  wire       [5:0]    _zz_2363_;
  wire       [63:0]   _zz_2364_;
  wire                _zz_2365_;
  wire                _zz_2366_;
  wire                _zz_2367_;
  wire                _zz_2368_;
  wire                _zz_2369_;
  wire                _zz_2370_;
  wire                _zz_2371_;
  wire                _zz_2372_;
  wire                _zz_2373_;
  wire                _zz_2374_;
  wire                _zz_2375_;
  wire                _zz_2376_;
  wire                _zz_2377_;
  wire                _zz_2378_;
  wire                _zz_2379_;
  wire                _zz_2380_;
  wire                _zz_2381_;
  wire                _zz_2382_;
  wire                _zz_2383_;
  wire                _zz_2384_;
  wire                _zz_2385_;
  wire                _zz_2386_;
  wire                _zz_2387_;
  wire                _zz_2388_;
  wire                _zz_2389_;
  wire                _zz_2390_;
  wire                _zz_2391_;
  wire                _zz_2392_;
  wire                _zz_2393_;
  wire                _zz_2394_;
  wire                _zz_2395_;
  wire                _zz_2396_;
  wire                _zz_2397_;
  wire                _zz_2398_;
  wire                _zz_2399_;
  wire                _zz_2400_;
  wire                _zz_2401_;
  wire                _zz_2402_;
  wire                _zz_2403_;
  wire                _zz_2404_;
  wire                _zz_2405_;
  wire                _zz_2406_;
  wire                _zz_2407_;
  wire                _zz_2408_;
  wire                _zz_2409_;
  wire                _zz_2410_;
  wire                _zz_2411_;
  wire                _zz_2412_;
  wire                _zz_2413_;
  wire                _zz_2414_;
  wire                _zz_2415_;
  wire                _zz_2416_;
  wire                _zz_2417_;
  wire                _zz_2418_;
  wire                _zz_2419_;
  wire                _zz_2420_;
  wire                _zz_2421_;
  wire                _zz_2422_;
  wire                _zz_2423_;
  wire                _zz_2424_;
  wire                _zz_2425_;
  wire                _zz_2426_;
  wire                _zz_2427_;
  wire                _zz_2428_;
  wire       [31:0]   _zz_2429_;
  wire       [15:0]   _zz_2430_;
  wire       [15:0]   _zz_2431_;
  wire       [5:0]    _zz_2432_;
  wire       [63:0]   _zz_2433_;
  wire                _zz_2434_;
  wire                _zz_2435_;
  wire                _zz_2436_;
  wire                _zz_2437_;
  wire                _zz_2438_;
  wire                _zz_2439_;
  wire                _zz_2440_;
  wire                _zz_2441_;
  wire                _zz_2442_;
  wire                _zz_2443_;
  wire                _zz_2444_;
  wire                _zz_2445_;
  wire                _zz_2446_;
  wire                _zz_2447_;
  wire                _zz_2448_;
  wire                _zz_2449_;
  wire                _zz_2450_;
  wire                _zz_2451_;
  wire                _zz_2452_;
  wire                _zz_2453_;
  wire                _zz_2454_;
  wire                _zz_2455_;
  wire                _zz_2456_;
  wire                _zz_2457_;
  wire                _zz_2458_;
  wire                _zz_2459_;
  wire                _zz_2460_;
  wire                _zz_2461_;
  wire                _zz_2462_;
  wire                _zz_2463_;
  wire                _zz_2464_;
  wire                _zz_2465_;
  wire                _zz_2466_;
  wire                _zz_2467_;
  wire                _zz_2468_;
  wire                _zz_2469_;
  wire                _zz_2470_;
  wire                _zz_2471_;
  wire                _zz_2472_;
  wire                _zz_2473_;
  wire                _zz_2474_;
  wire                _zz_2475_;
  wire                _zz_2476_;
  wire                _zz_2477_;
  wire                _zz_2478_;
  wire                _zz_2479_;
  wire                _zz_2480_;
  wire                _zz_2481_;
  wire                _zz_2482_;
  wire                _zz_2483_;
  wire                _zz_2484_;
  wire                _zz_2485_;
  wire                _zz_2486_;
  wire                _zz_2487_;
  wire                _zz_2488_;
  wire                _zz_2489_;
  wire                _zz_2490_;
  wire                _zz_2491_;
  wire                _zz_2492_;
  wire                _zz_2493_;
  wire                _zz_2494_;
  wire                _zz_2495_;
  wire                _zz_2496_;
  wire                _zz_2497_;
  wire       [31:0]   _zz_2498_;
  wire       [15:0]   _zz_2499_;
  wire       [15:0]   _zz_2500_;
  wire       [5:0]    _zz_2501_;
  wire       [63:0]   _zz_2502_;
  wire                _zz_2503_;
  wire                _zz_2504_;
  wire                _zz_2505_;
  wire                _zz_2506_;
  wire                _zz_2507_;
  wire                _zz_2508_;
  wire                _zz_2509_;
  wire                _zz_2510_;
  wire                _zz_2511_;
  wire                _zz_2512_;
  wire                _zz_2513_;
  wire                _zz_2514_;
  wire                _zz_2515_;
  wire                _zz_2516_;
  wire                _zz_2517_;
  wire                _zz_2518_;
  wire                _zz_2519_;
  wire                _zz_2520_;
  wire                _zz_2521_;
  wire                _zz_2522_;
  wire                _zz_2523_;
  wire                _zz_2524_;
  wire                _zz_2525_;
  wire                _zz_2526_;
  wire                _zz_2527_;
  wire                _zz_2528_;
  wire                _zz_2529_;
  wire                _zz_2530_;
  wire                _zz_2531_;
  wire                _zz_2532_;
  wire                _zz_2533_;
  wire                _zz_2534_;
  wire                _zz_2535_;
  wire                _zz_2536_;
  wire                _zz_2537_;
  wire                _zz_2538_;
  wire                _zz_2539_;
  wire                _zz_2540_;
  wire                _zz_2541_;
  wire                _zz_2542_;
  wire                _zz_2543_;
  wire                _zz_2544_;
  wire                _zz_2545_;
  wire                _zz_2546_;
  wire                _zz_2547_;
  wire                _zz_2548_;
  wire                _zz_2549_;
  wire                _zz_2550_;
  wire                _zz_2551_;
  wire                _zz_2552_;
  wire                _zz_2553_;
  wire                _zz_2554_;
  wire                _zz_2555_;
  wire                _zz_2556_;
  wire                _zz_2557_;
  wire                _zz_2558_;
  wire                _zz_2559_;
  wire                _zz_2560_;
  wire                _zz_2561_;
  wire                _zz_2562_;
  wire                _zz_2563_;
  wire                _zz_2564_;
  wire                _zz_2565_;
  wire                _zz_2566_;
  wire       [31:0]   _zz_2567_;
  wire       [15:0]   _zz_2568_;
  wire       [15:0]   _zz_2569_;
  wire       [5:0]    _zz_2570_;
  wire       [63:0]   _zz_2571_;
  wire                _zz_2572_;
  wire                _zz_2573_;
  wire                _zz_2574_;
  wire                _zz_2575_;
  wire                _zz_2576_;
  wire                _zz_2577_;
  wire                _zz_2578_;
  wire                _zz_2579_;
  wire                _zz_2580_;
  wire                _zz_2581_;
  wire                _zz_2582_;
  wire                _zz_2583_;
  wire                _zz_2584_;
  wire                _zz_2585_;
  wire                _zz_2586_;
  wire                _zz_2587_;
  wire                _zz_2588_;
  wire                _zz_2589_;
  wire                _zz_2590_;
  wire                _zz_2591_;
  wire                _zz_2592_;
  wire                _zz_2593_;
  wire                _zz_2594_;
  wire                _zz_2595_;
  wire                _zz_2596_;
  wire                _zz_2597_;
  wire                _zz_2598_;
  wire                _zz_2599_;
  wire                _zz_2600_;
  wire                _zz_2601_;
  wire                _zz_2602_;
  wire                _zz_2603_;
  wire                _zz_2604_;
  wire                _zz_2605_;
  wire                _zz_2606_;
  wire                _zz_2607_;
  wire                _zz_2608_;
  wire                _zz_2609_;
  wire                _zz_2610_;
  wire                _zz_2611_;
  wire                _zz_2612_;
  wire                _zz_2613_;
  wire                _zz_2614_;
  wire                _zz_2615_;
  wire                _zz_2616_;
  wire                _zz_2617_;
  wire                _zz_2618_;
  wire                _zz_2619_;
  wire                _zz_2620_;
  wire                _zz_2621_;
  wire                _zz_2622_;
  wire                _zz_2623_;
  wire                _zz_2624_;
  wire                _zz_2625_;
  wire                _zz_2626_;
  wire                _zz_2627_;
  wire                _zz_2628_;
  wire                _zz_2629_;
  wire                _zz_2630_;
  wire                _zz_2631_;
  wire                _zz_2632_;
  wire                _zz_2633_;
  wire                _zz_2634_;
  wire                _zz_2635_;
  wire       [31:0]   _zz_2636_;
  wire       [15:0]   _zz_2637_;
  wire       [15:0]   _zz_2638_;
  wire       [5:0]    _zz_2639_;
  wire       [63:0]   _zz_2640_;
  wire                _zz_2641_;
  wire                _zz_2642_;
  wire                _zz_2643_;
  wire                _zz_2644_;
  wire                _zz_2645_;
  wire                _zz_2646_;
  wire                _zz_2647_;
  wire                _zz_2648_;
  wire                _zz_2649_;
  wire                _zz_2650_;
  wire                _zz_2651_;
  wire                _zz_2652_;
  wire                _zz_2653_;
  wire                _zz_2654_;
  wire                _zz_2655_;
  wire                _zz_2656_;
  wire                _zz_2657_;
  wire                _zz_2658_;
  wire                _zz_2659_;
  wire                _zz_2660_;
  wire                _zz_2661_;
  wire                _zz_2662_;
  wire                _zz_2663_;
  wire                _zz_2664_;
  wire                _zz_2665_;
  wire                _zz_2666_;
  wire                _zz_2667_;
  wire                _zz_2668_;
  wire                _zz_2669_;
  wire                _zz_2670_;
  wire                _zz_2671_;
  wire                _zz_2672_;
  wire                _zz_2673_;
  wire                _zz_2674_;
  wire                _zz_2675_;
  wire                _zz_2676_;
  wire                _zz_2677_;
  wire                _zz_2678_;
  wire                _zz_2679_;
  wire                _zz_2680_;
  wire                _zz_2681_;
  wire                _zz_2682_;
  wire                _zz_2683_;
  wire                _zz_2684_;
  wire                _zz_2685_;
  wire                _zz_2686_;
  wire                _zz_2687_;
  wire                _zz_2688_;
  wire                _zz_2689_;
  wire                _zz_2690_;
  wire                _zz_2691_;
  wire                _zz_2692_;
  wire                _zz_2693_;
  wire                _zz_2694_;
  wire                _zz_2695_;
  wire                _zz_2696_;
  wire                _zz_2697_;
  wire                _zz_2698_;
  wire                _zz_2699_;
  wire                _zz_2700_;
  wire                _zz_2701_;
  wire                _zz_2702_;
  wire                _zz_2703_;
  wire                _zz_2704_;
  wire       [31:0]   _zz_2705_;
  wire       [15:0]   _zz_2706_;
  wire       [15:0]   _zz_2707_;
  wire       [5:0]    _zz_2708_;
  wire       [63:0]   _zz_2709_;
  wire                _zz_2710_;
  wire                _zz_2711_;
  wire                _zz_2712_;
  wire                _zz_2713_;
  wire                _zz_2714_;
  wire                _zz_2715_;
  wire                _zz_2716_;
  wire                _zz_2717_;
  wire                _zz_2718_;
  wire                _zz_2719_;
  wire                _zz_2720_;
  wire                _zz_2721_;
  wire                _zz_2722_;
  wire                _zz_2723_;
  wire                _zz_2724_;
  wire                _zz_2725_;
  wire                _zz_2726_;
  wire                _zz_2727_;
  wire                _zz_2728_;
  wire                _zz_2729_;
  wire                _zz_2730_;
  wire                _zz_2731_;
  wire                _zz_2732_;
  wire                _zz_2733_;
  wire                _zz_2734_;
  wire                _zz_2735_;
  wire                _zz_2736_;
  wire                _zz_2737_;
  wire                _zz_2738_;
  wire                _zz_2739_;
  wire                _zz_2740_;
  wire                _zz_2741_;
  wire                _zz_2742_;
  wire                _zz_2743_;
  wire                _zz_2744_;
  wire                _zz_2745_;
  wire                _zz_2746_;
  wire                _zz_2747_;
  wire                _zz_2748_;
  wire                _zz_2749_;
  wire                _zz_2750_;
  wire                _zz_2751_;
  wire                _zz_2752_;
  wire                _zz_2753_;
  wire                _zz_2754_;
  wire                _zz_2755_;
  wire                _zz_2756_;
  wire                _zz_2757_;
  wire                _zz_2758_;
  wire                _zz_2759_;
  wire                _zz_2760_;
  wire                _zz_2761_;
  wire                _zz_2762_;
  wire                _zz_2763_;
  wire                _zz_2764_;
  wire                _zz_2765_;
  wire                _zz_2766_;
  wire                _zz_2767_;
  wire                _zz_2768_;
  wire                _zz_2769_;
  wire                _zz_2770_;
  wire                _zz_2771_;
  wire                _zz_2772_;
  wire                _zz_2773_;
  wire       [31:0]   _zz_2774_;
  wire       [15:0]   _zz_2775_;
  wire       [15:0]   _zz_2776_;
  wire       [5:0]    _zz_2777_;
  wire       [63:0]   _zz_2778_;
  wire                _zz_2779_;
  wire                _zz_2780_;
  wire                _zz_2781_;
  wire                _zz_2782_;
  wire                _zz_2783_;
  wire                _zz_2784_;
  wire                _zz_2785_;
  wire                _zz_2786_;
  wire                _zz_2787_;
  wire                _zz_2788_;
  wire                _zz_2789_;
  wire                _zz_2790_;
  wire                _zz_2791_;
  wire                _zz_2792_;
  wire                _zz_2793_;
  wire                _zz_2794_;
  wire                _zz_2795_;
  wire                _zz_2796_;
  wire                _zz_2797_;
  wire                _zz_2798_;
  wire                _zz_2799_;
  wire                _zz_2800_;
  wire                _zz_2801_;
  wire                _zz_2802_;
  wire                _zz_2803_;
  wire                _zz_2804_;
  wire                _zz_2805_;
  wire                _zz_2806_;
  wire                _zz_2807_;
  wire                _zz_2808_;
  wire                _zz_2809_;
  wire                _zz_2810_;
  wire                _zz_2811_;
  wire                _zz_2812_;
  wire                _zz_2813_;
  wire                _zz_2814_;
  wire                _zz_2815_;
  wire                _zz_2816_;
  wire                _zz_2817_;
  wire                _zz_2818_;
  wire                _zz_2819_;
  wire                _zz_2820_;
  wire                _zz_2821_;
  wire                _zz_2822_;
  wire                _zz_2823_;
  wire                _zz_2824_;
  wire                _zz_2825_;
  wire                _zz_2826_;
  wire                _zz_2827_;
  wire                _zz_2828_;
  wire                _zz_2829_;
  wire                _zz_2830_;
  wire                _zz_2831_;
  wire                _zz_2832_;
  wire                _zz_2833_;
  wire                _zz_2834_;
  wire                _zz_2835_;
  wire                _zz_2836_;
  wire                _zz_2837_;
  wire                _zz_2838_;
  wire                _zz_2839_;
  wire                _zz_2840_;
  wire                _zz_2841_;
  wire                _zz_2842_;
  wire       [31:0]   _zz_2843_;
  wire       [15:0]   _zz_2844_;
  wire       [15:0]   _zz_2845_;
  wire       [5:0]    _zz_2846_;
  wire       [63:0]   _zz_2847_;
  wire                _zz_2848_;
  wire                _zz_2849_;
  wire                _zz_2850_;
  wire                _zz_2851_;
  wire                _zz_2852_;
  wire                _zz_2853_;
  wire                _zz_2854_;
  wire                _zz_2855_;
  wire                _zz_2856_;
  wire                _zz_2857_;
  wire                _zz_2858_;
  wire                _zz_2859_;
  wire                _zz_2860_;
  wire                _zz_2861_;
  wire                _zz_2862_;
  wire                _zz_2863_;
  wire                _zz_2864_;
  wire                _zz_2865_;
  wire                _zz_2866_;
  wire                _zz_2867_;
  wire                _zz_2868_;
  wire                _zz_2869_;
  wire                _zz_2870_;
  wire                _zz_2871_;
  wire                _zz_2872_;
  wire                _zz_2873_;
  wire                _zz_2874_;
  wire                _zz_2875_;
  wire                _zz_2876_;
  wire                _zz_2877_;
  wire                _zz_2878_;
  wire                _zz_2879_;
  wire                _zz_2880_;
  wire                _zz_2881_;
  wire                _zz_2882_;
  wire                _zz_2883_;
  wire                _zz_2884_;
  wire                _zz_2885_;
  wire                _zz_2886_;
  wire                _zz_2887_;
  wire                _zz_2888_;
  wire                _zz_2889_;
  wire                _zz_2890_;
  wire                _zz_2891_;
  wire                _zz_2892_;
  wire                _zz_2893_;
  wire                _zz_2894_;
  wire                _zz_2895_;
  wire                _zz_2896_;
  wire                _zz_2897_;
  wire                _zz_2898_;
  wire                _zz_2899_;
  wire                _zz_2900_;
  wire                _zz_2901_;
  wire                _zz_2902_;
  wire                _zz_2903_;
  wire                _zz_2904_;
  wire                _zz_2905_;
  wire                _zz_2906_;
  wire                _zz_2907_;
  wire                _zz_2908_;
  wire                _zz_2909_;
  wire                _zz_2910_;
  wire                _zz_2911_;
  wire       [31:0]   _zz_2912_;
  wire       [15:0]   _zz_2913_;
  wire       [15:0]   _zz_2914_;
  wire       [5:0]    _zz_2915_;
  wire       [63:0]   _zz_2916_;
  wire                _zz_2917_;
  wire                _zz_2918_;
  wire                _zz_2919_;
  wire                _zz_2920_;
  wire                _zz_2921_;
  wire                _zz_2922_;
  wire                _zz_2923_;
  wire                _zz_2924_;
  wire                _zz_2925_;
  wire                _zz_2926_;
  wire                _zz_2927_;
  wire                _zz_2928_;
  wire                _zz_2929_;
  wire                _zz_2930_;
  wire                _zz_2931_;
  wire                _zz_2932_;
  wire                _zz_2933_;
  wire                _zz_2934_;
  wire                _zz_2935_;
  wire                _zz_2936_;
  wire                _zz_2937_;
  wire                _zz_2938_;
  wire                _zz_2939_;
  wire                _zz_2940_;
  wire                _zz_2941_;
  wire                _zz_2942_;
  wire                _zz_2943_;
  wire                _zz_2944_;
  wire                _zz_2945_;
  wire                _zz_2946_;
  wire                _zz_2947_;
  wire                _zz_2948_;
  wire                _zz_2949_;
  wire                _zz_2950_;
  wire                _zz_2951_;
  wire                _zz_2952_;
  wire                _zz_2953_;
  wire                _zz_2954_;
  wire                _zz_2955_;
  wire                _zz_2956_;
  wire                _zz_2957_;
  wire                _zz_2958_;
  wire                _zz_2959_;
  wire                _zz_2960_;
  wire                _zz_2961_;
  wire                _zz_2962_;
  wire                _zz_2963_;
  wire                _zz_2964_;
  wire                _zz_2965_;
  wire                _zz_2966_;
  wire                _zz_2967_;
  wire                _zz_2968_;
  wire                _zz_2969_;
  wire                _zz_2970_;
  wire                _zz_2971_;
  wire                _zz_2972_;
  wire                _zz_2973_;
  wire                _zz_2974_;
  wire                _zz_2975_;
  wire                _zz_2976_;
  wire                _zz_2977_;
  wire                _zz_2978_;
  wire                _zz_2979_;
  wire                _zz_2980_;
  wire       [31:0]   _zz_2981_;
  wire       [15:0]   _zz_2982_;
  wire       [15:0]   _zz_2983_;
  wire       [5:0]    _zz_2984_;
  wire       [63:0]   _zz_2985_;
  wire                _zz_2986_;
  wire                _zz_2987_;
  wire                _zz_2988_;
  wire                _zz_2989_;
  wire                _zz_2990_;
  wire                _zz_2991_;
  wire                _zz_2992_;
  wire                _zz_2993_;
  wire                _zz_2994_;
  wire                _zz_2995_;
  wire                _zz_2996_;
  wire                _zz_2997_;
  wire                _zz_2998_;
  wire                _zz_2999_;
  wire                _zz_3000_;
  wire                _zz_3001_;
  wire                _zz_3002_;
  wire                _zz_3003_;
  wire                _zz_3004_;
  wire                _zz_3005_;
  wire                _zz_3006_;
  wire                _zz_3007_;
  wire                _zz_3008_;
  wire                _zz_3009_;
  wire                _zz_3010_;
  wire                _zz_3011_;
  wire                _zz_3012_;
  wire                _zz_3013_;
  wire                _zz_3014_;
  wire                _zz_3015_;
  wire                _zz_3016_;
  wire                _zz_3017_;
  wire                _zz_3018_;
  wire                _zz_3019_;
  wire                _zz_3020_;
  wire                _zz_3021_;
  wire                _zz_3022_;
  wire                _zz_3023_;
  wire                _zz_3024_;
  wire                _zz_3025_;
  wire                _zz_3026_;
  wire                _zz_3027_;
  wire                _zz_3028_;
  wire                _zz_3029_;
  wire                _zz_3030_;
  wire                _zz_3031_;
  wire                _zz_3032_;
  wire                _zz_3033_;
  wire                _zz_3034_;
  wire                _zz_3035_;
  wire                _zz_3036_;
  wire                _zz_3037_;
  wire                _zz_3038_;
  wire                _zz_3039_;
  wire                _zz_3040_;
  wire                _zz_3041_;
  wire                _zz_3042_;
  wire                _zz_3043_;
  wire                _zz_3044_;
  wire                _zz_3045_;
  wire                _zz_3046_;
  wire                _zz_3047_;
  wire                _zz_3048_;
  wire                _zz_3049_;
  wire       [31:0]   _zz_3050_;
  wire       [15:0]   _zz_3051_;
  wire       [15:0]   _zz_3052_;
  wire       [5:0]    _zz_3053_;
  wire       [63:0]   _zz_3054_;
  wire                _zz_3055_;
  wire                _zz_3056_;
  wire                _zz_3057_;
  wire                _zz_3058_;
  wire                _zz_3059_;
  wire                _zz_3060_;
  wire                _zz_3061_;
  wire                _zz_3062_;
  wire                _zz_3063_;
  wire                _zz_3064_;
  wire                _zz_3065_;
  wire                _zz_3066_;
  wire                _zz_3067_;
  wire                _zz_3068_;
  wire                _zz_3069_;
  wire                _zz_3070_;
  wire                _zz_3071_;
  wire                _zz_3072_;
  wire                _zz_3073_;
  wire                _zz_3074_;
  wire                _zz_3075_;
  wire                _zz_3076_;
  wire                _zz_3077_;
  wire                _zz_3078_;
  wire                _zz_3079_;
  wire                _zz_3080_;
  wire                _zz_3081_;
  wire                _zz_3082_;
  wire                _zz_3083_;
  wire                _zz_3084_;
  wire                _zz_3085_;
  wire                _zz_3086_;
  wire                _zz_3087_;
  wire                _zz_3088_;
  wire                _zz_3089_;
  wire                _zz_3090_;
  wire                _zz_3091_;
  wire                _zz_3092_;
  wire                _zz_3093_;
  wire                _zz_3094_;
  wire                _zz_3095_;
  wire                _zz_3096_;
  wire                _zz_3097_;
  wire                _zz_3098_;
  wire                _zz_3099_;
  wire                _zz_3100_;
  wire                _zz_3101_;
  wire                _zz_3102_;
  wire                _zz_3103_;
  wire                _zz_3104_;
  wire                _zz_3105_;
  wire                _zz_3106_;
  wire                _zz_3107_;
  wire                _zz_3108_;
  wire                _zz_3109_;
  wire                _zz_3110_;
  wire                _zz_3111_;
  wire                _zz_3112_;
  wire                _zz_3113_;
  wire                _zz_3114_;
  wire                _zz_3115_;
  wire                _zz_3116_;
  wire                _zz_3117_;
  wire                _zz_3118_;
  wire       [31:0]   _zz_3119_;
  wire       [15:0]   _zz_3120_;
  wire       [15:0]   _zz_3121_;
  wire       [5:0]    _zz_3122_;
  wire       [63:0]   _zz_3123_;
  wire                _zz_3124_;
  wire                _zz_3125_;
  wire                _zz_3126_;
  wire                _zz_3127_;
  wire                _zz_3128_;
  wire                _zz_3129_;
  wire                _zz_3130_;
  wire                _zz_3131_;
  wire                _zz_3132_;
  wire                _zz_3133_;
  wire                _zz_3134_;
  wire                _zz_3135_;
  wire                _zz_3136_;
  wire                _zz_3137_;
  wire                _zz_3138_;
  wire                _zz_3139_;
  wire                _zz_3140_;
  wire                _zz_3141_;
  wire                _zz_3142_;
  wire                _zz_3143_;
  wire                _zz_3144_;
  wire                _zz_3145_;
  wire                _zz_3146_;
  wire                _zz_3147_;
  wire                _zz_3148_;
  wire                _zz_3149_;
  wire                _zz_3150_;
  wire                _zz_3151_;
  wire                _zz_3152_;
  wire                _zz_3153_;
  wire                _zz_3154_;
  wire                _zz_3155_;
  wire                _zz_3156_;
  wire                _zz_3157_;
  wire                _zz_3158_;
  wire                _zz_3159_;
  wire                _zz_3160_;
  wire                _zz_3161_;
  wire                _zz_3162_;
  wire                _zz_3163_;
  wire                _zz_3164_;
  wire                _zz_3165_;
  wire                _zz_3166_;
  wire                _zz_3167_;
  wire                _zz_3168_;
  wire                _zz_3169_;
  wire                _zz_3170_;
  wire                _zz_3171_;
  wire                _zz_3172_;
  wire                _zz_3173_;
  wire                _zz_3174_;
  wire                _zz_3175_;
  wire                _zz_3176_;
  wire                _zz_3177_;
  wire                _zz_3178_;
  wire                _zz_3179_;
  wire                _zz_3180_;
  wire                _zz_3181_;
  wire                _zz_3182_;
  wire                _zz_3183_;
  wire                _zz_3184_;
  wire                _zz_3185_;
  wire                _zz_3186_;
  wire                _zz_3187_;
  wire       [31:0]   _zz_3188_;
  wire       [15:0]   _zz_3189_;
  wire       [15:0]   _zz_3190_;
  wire       [5:0]    _zz_3191_;
  wire       [63:0]   _zz_3192_;
  wire                _zz_3193_;
  wire                _zz_3194_;
  wire                _zz_3195_;
  wire                _zz_3196_;
  wire                _zz_3197_;
  wire                _zz_3198_;
  wire                _zz_3199_;
  wire                _zz_3200_;
  wire                _zz_3201_;
  wire                _zz_3202_;
  wire                _zz_3203_;
  wire                _zz_3204_;
  wire                _zz_3205_;
  wire                _zz_3206_;
  wire                _zz_3207_;
  wire                _zz_3208_;
  wire                _zz_3209_;
  wire                _zz_3210_;
  wire                _zz_3211_;
  wire                _zz_3212_;
  wire                _zz_3213_;
  wire                _zz_3214_;
  wire                _zz_3215_;
  wire                _zz_3216_;
  wire                _zz_3217_;
  wire                _zz_3218_;
  wire                _zz_3219_;
  wire                _zz_3220_;
  wire                _zz_3221_;
  wire                _zz_3222_;
  wire                _zz_3223_;
  wire                _zz_3224_;
  wire                _zz_3225_;
  wire                _zz_3226_;
  wire                _zz_3227_;
  wire                _zz_3228_;
  wire                _zz_3229_;
  wire                _zz_3230_;
  wire                _zz_3231_;
  wire                _zz_3232_;
  wire                _zz_3233_;
  wire                _zz_3234_;
  wire                _zz_3235_;
  wire                _zz_3236_;
  wire                _zz_3237_;
  wire                _zz_3238_;
  wire                _zz_3239_;
  wire                _zz_3240_;
  wire                _zz_3241_;
  wire                _zz_3242_;
  wire                _zz_3243_;
  wire                _zz_3244_;
  wire                _zz_3245_;
  wire                _zz_3246_;
  wire                _zz_3247_;
  wire                _zz_3248_;
  wire                _zz_3249_;
  wire                _zz_3250_;
  wire                _zz_3251_;
  wire                _zz_3252_;
  wire                _zz_3253_;
  wire                _zz_3254_;
  wire                _zz_3255_;
  wire                _zz_3256_;
  wire       [31:0]   _zz_3257_;
  wire       [15:0]   _zz_3258_;
  wire       [15:0]   _zz_3259_;
  wire       [5:0]    _zz_3260_;
  wire       [63:0]   _zz_3261_;
  wire                _zz_3262_;
  wire                _zz_3263_;
  wire                _zz_3264_;
  wire                _zz_3265_;
  wire                _zz_3266_;
  wire                _zz_3267_;
  wire                _zz_3268_;
  wire                _zz_3269_;
  wire                _zz_3270_;
  wire                _zz_3271_;
  wire                _zz_3272_;
  wire                _zz_3273_;
  wire                _zz_3274_;
  wire                _zz_3275_;
  wire                _zz_3276_;
  wire                _zz_3277_;
  wire                _zz_3278_;
  wire                _zz_3279_;
  wire                _zz_3280_;
  wire                _zz_3281_;
  wire                _zz_3282_;
  wire                _zz_3283_;
  wire                _zz_3284_;
  wire                _zz_3285_;
  wire                _zz_3286_;
  wire                _zz_3287_;
  wire                _zz_3288_;
  wire                _zz_3289_;
  wire                _zz_3290_;
  wire                _zz_3291_;
  wire                _zz_3292_;
  wire                _zz_3293_;
  wire                _zz_3294_;
  wire                _zz_3295_;
  wire                _zz_3296_;
  wire                _zz_3297_;
  wire                _zz_3298_;
  wire                _zz_3299_;
  wire                _zz_3300_;
  wire                _zz_3301_;
  wire                _zz_3302_;
  wire                _zz_3303_;
  wire                _zz_3304_;
  wire                _zz_3305_;
  wire                _zz_3306_;
  wire                _zz_3307_;
  wire                _zz_3308_;
  wire                _zz_3309_;
  wire                _zz_3310_;
  wire                _zz_3311_;
  wire                _zz_3312_;
  wire                _zz_3313_;
  wire                _zz_3314_;
  wire                _zz_3315_;
  wire                _zz_3316_;
  wire                _zz_3317_;
  wire                _zz_3318_;
  wire                _zz_3319_;
  wire                _zz_3320_;
  wire                _zz_3321_;
  wire                _zz_3322_;
  wire                _zz_3323_;
  wire                _zz_3324_;
  wire                _zz_3325_;
  wire       [31:0]   _zz_3326_;
  wire       [15:0]   _zz_3327_;
  wire       [15:0]   _zz_3328_;
  wire       [5:0]    _zz_3329_;
  wire       [63:0]   _zz_3330_;
  wire                _zz_3331_;
  wire                _zz_3332_;
  wire                _zz_3333_;
  wire                _zz_3334_;
  wire                _zz_3335_;
  wire                _zz_3336_;
  wire                _zz_3337_;
  wire                _zz_3338_;
  wire                _zz_3339_;
  wire                _zz_3340_;
  wire                _zz_3341_;
  wire                _zz_3342_;
  wire                _zz_3343_;
  wire                _zz_3344_;
  wire                _zz_3345_;
  wire                _zz_3346_;
  wire                _zz_3347_;
  wire                _zz_3348_;
  wire                _zz_3349_;
  wire                _zz_3350_;
  wire                _zz_3351_;
  wire                _zz_3352_;
  wire                _zz_3353_;
  wire                _zz_3354_;
  wire                _zz_3355_;
  wire                _zz_3356_;
  wire                _zz_3357_;
  wire                _zz_3358_;
  wire                _zz_3359_;
  wire                _zz_3360_;
  wire                _zz_3361_;
  wire                _zz_3362_;
  wire                _zz_3363_;
  wire                _zz_3364_;
  wire                _zz_3365_;
  wire                _zz_3366_;
  wire                _zz_3367_;
  wire                _zz_3368_;
  wire                _zz_3369_;
  wire                _zz_3370_;
  wire                _zz_3371_;
  wire                _zz_3372_;
  wire                _zz_3373_;
  wire                _zz_3374_;
  wire                _zz_3375_;
  wire                _zz_3376_;
  wire                _zz_3377_;
  wire                _zz_3378_;
  wire                _zz_3379_;
  wire                _zz_3380_;
  wire                _zz_3381_;
  wire                _zz_3382_;
  wire                _zz_3383_;
  wire                _zz_3384_;
  wire                _zz_3385_;
  wire                _zz_3386_;
  wire                _zz_3387_;
  wire                _zz_3388_;
  wire                _zz_3389_;
  wire                _zz_3390_;
  wire                _zz_3391_;
  wire                _zz_3392_;
  wire                _zz_3393_;
  wire                _zz_3394_;
  wire       [31:0]   _zz_3395_;
  wire       [15:0]   _zz_3396_;
  wire       [15:0]   _zz_3397_;
  wire       [5:0]    _zz_3398_;
  wire       [63:0]   _zz_3399_;
  wire                _zz_3400_;
  wire                _zz_3401_;
  wire                _zz_3402_;
  wire                _zz_3403_;
  wire                _zz_3404_;
  wire                _zz_3405_;
  wire                _zz_3406_;
  wire                _zz_3407_;
  wire                _zz_3408_;
  wire                _zz_3409_;
  wire                _zz_3410_;
  wire                _zz_3411_;
  wire                _zz_3412_;
  wire                _zz_3413_;
  wire                _zz_3414_;
  wire                _zz_3415_;
  wire                _zz_3416_;
  wire                _zz_3417_;
  wire                _zz_3418_;
  wire                _zz_3419_;
  wire                _zz_3420_;
  wire                _zz_3421_;
  wire                _zz_3422_;
  wire                _zz_3423_;
  wire                _zz_3424_;
  wire                _zz_3425_;
  wire                _zz_3426_;
  wire                _zz_3427_;
  wire                _zz_3428_;
  wire                _zz_3429_;
  wire                _zz_3430_;
  wire                _zz_3431_;
  wire                _zz_3432_;
  wire                _zz_3433_;
  wire                _zz_3434_;
  wire                _zz_3435_;
  wire                _zz_3436_;
  wire                _zz_3437_;
  wire                _zz_3438_;
  wire                _zz_3439_;
  wire                _zz_3440_;
  wire                _zz_3441_;
  wire                _zz_3442_;
  wire                _zz_3443_;
  wire                _zz_3444_;
  wire                _zz_3445_;
  wire                _zz_3446_;
  wire                _zz_3447_;
  wire                _zz_3448_;
  wire                _zz_3449_;
  wire                _zz_3450_;
  wire                _zz_3451_;
  wire                _zz_3452_;
  wire                _zz_3453_;
  wire                _zz_3454_;
  wire                _zz_3455_;
  wire                _zz_3456_;
  wire                _zz_3457_;
  wire                _zz_3458_;
  wire                _zz_3459_;
  wire                _zz_3460_;
  wire                _zz_3461_;
  wire                _zz_3462_;
  wire                _zz_3463_;
  wire       [31:0]   _zz_3464_;
  wire       [15:0]   _zz_3465_;
  wire       [15:0]   _zz_3466_;
  wire       [5:0]    _zz_3467_;
  wire       [63:0]   _zz_3468_;
  wire                _zz_3469_;
  wire                _zz_3470_;
  wire                _zz_3471_;
  wire                _zz_3472_;
  wire                _zz_3473_;
  wire                _zz_3474_;
  wire                _zz_3475_;
  wire                _zz_3476_;
  wire                _zz_3477_;
  wire                _zz_3478_;
  wire                _zz_3479_;
  wire                _zz_3480_;
  wire                _zz_3481_;
  wire                _zz_3482_;
  wire                _zz_3483_;
  wire                _zz_3484_;
  wire                _zz_3485_;
  wire                _zz_3486_;
  wire                _zz_3487_;
  wire                _zz_3488_;
  wire                _zz_3489_;
  wire                _zz_3490_;
  wire                _zz_3491_;
  wire                _zz_3492_;
  wire                _zz_3493_;
  wire                _zz_3494_;
  wire                _zz_3495_;
  wire                _zz_3496_;
  wire                _zz_3497_;
  wire                _zz_3498_;
  wire                _zz_3499_;
  wire                _zz_3500_;
  wire                _zz_3501_;
  wire                _zz_3502_;
  wire                _zz_3503_;
  wire                _zz_3504_;
  wire                _zz_3505_;
  wire                _zz_3506_;
  wire                _zz_3507_;
  wire                _zz_3508_;
  wire                _zz_3509_;
  wire                _zz_3510_;
  wire                _zz_3511_;
  wire                _zz_3512_;
  wire                _zz_3513_;
  wire                _zz_3514_;
  wire                _zz_3515_;
  wire                _zz_3516_;
  wire                _zz_3517_;
  wire                _zz_3518_;
  wire                _zz_3519_;
  wire                _zz_3520_;
  wire                _zz_3521_;
  wire                _zz_3522_;
  wire                _zz_3523_;
  wire                _zz_3524_;
  wire                _zz_3525_;
  wire                _zz_3526_;
  wire                _zz_3527_;
  wire                _zz_3528_;
  wire                _zz_3529_;
  wire                _zz_3530_;
  wire                _zz_3531_;
  wire                _zz_3532_;
  wire       [31:0]   _zz_3533_;
  wire       [15:0]   _zz_3534_;
  wire       [15:0]   _zz_3535_;
  wire       [5:0]    _zz_3536_;
  wire       [63:0]   _zz_3537_;
  wire                _zz_3538_;
  wire                _zz_3539_;
  wire                _zz_3540_;
  wire                _zz_3541_;
  wire                _zz_3542_;
  wire                _zz_3543_;
  wire                _zz_3544_;
  wire                _zz_3545_;
  wire                _zz_3546_;
  wire                _zz_3547_;
  wire                _zz_3548_;
  wire                _zz_3549_;
  wire                _zz_3550_;
  wire                _zz_3551_;
  wire                _zz_3552_;
  wire                _zz_3553_;
  wire                _zz_3554_;
  wire                _zz_3555_;
  wire                _zz_3556_;
  wire                _zz_3557_;
  wire                _zz_3558_;
  wire                _zz_3559_;
  wire                _zz_3560_;
  wire                _zz_3561_;
  wire                _zz_3562_;
  wire                _zz_3563_;
  wire                _zz_3564_;
  wire                _zz_3565_;
  wire                _zz_3566_;
  wire                _zz_3567_;
  wire                _zz_3568_;
  wire                _zz_3569_;
  wire                _zz_3570_;
  wire                _zz_3571_;
  wire                _zz_3572_;
  wire                _zz_3573_;
  wire                _zz_3574_;
  wire                _zz_3575_;
  wire                _zz_3576_;
  wire                _zz_3577_;
  wire                _zz_3578_;
  wire                _zz_3579_;
  wire                _zz_3580_;
  wire                _zz_3581_;
  wire                _zz_3582_;
  wire                _zz_3583_;
  wire                _zz_3584_;
  wire                _zz_3585_;
  wire                _zz_3586_;
  wire                _zz_3587_;
  wire                _zz_3588_;
  wire                _zz_3589_;
  wire                _zz_3590_;
  wire                _zz_3591_;
  wire                _zz_3592_;
  wire                _zz_3593_;
  wire                _zz_3594_;
  wire                _zz_3595_;
  wire                _zz_3596_;
  wire                _zz_3597_;
  wire                _zz_3598_;
  wire                _zz_3599_;
  wire                _zz_3600_;
  wire                _zz_3601_;
  wire       [31:0]   _zz_3602_;
  wire       [15:0]   _zz_3603_;
  wire       [15:0]   _zz_3604_;
  wire       [5:0]    _zz_3605_;
  wire       [63:0]   _zz_3606_;
  wire                _zz_3607_;
  wire                _zz_3608_;
  wire                _zz_3609_;
  wire                _zz_3610_;
  wire                _zz_3611_;
  wire                _zz_3612_;
  wire                _zz_3613_;
  wire                _zz_3614_;
  wire                _zz_3615_;
  wire                _zz_3616_;
  wire                _zz_3617_;
  wire                _zz_3618_;
  wire                _zz_3619_;
  wire                _zz_3620_;
  wire                _zz_3621_;
  wire                _zz_3622_;
  wire                _zz_3623_;
  wire                _zz_3624_;
  wire                _zz_3625_;
  wire                _zz_3626_;
  wire                _zz_3627_;
  wire                _zz_3628_;
  wire                _zz_3629_;
  wire                _zz_3630_;
  wire                _zz_3631_;
  wire                _zz_3632_;
  wire                _zz_3633_;
  wire                _zz_3634_;
  wire                _zz_3635_;
  wire                _zz_3636_;
  wire                _zz_3637_;
  wire                _zz_3638_;
  wire                _zz_3639_;
  wire                _zz_3640_;
  wire                _zz_3641_;
  wire                _zz_3642_;
  wire                _zz_3643_;
  wire                _zz_3644_;
  wire                _zz_3645_;
  wire                _zz_3646_;
  wire                _zz_3647_;
  wire                _zz_3648_;
  wire                _zz_3649_;
  wire                _zz_3650_;
  wire                _zz_3651_;
  wire                _zz_3652_;
  wire                _zz_3653_;
  wire                _zz_3654_;
  wire                _zz_3655_;
  wire                _zz_3656_;
  wire                _zz_3657_;
  wire                _zz_3658_;
  wire                _zz_3659_;
  wire                _zz_3660_;
  wire                _zz_3661_;
  wire                _zz_3662_;
  wire                _zz_3663_;
  wire                _zz_3664_;
  wire                _zz_3665_;
  wire                _zz_3666_;
  wire                _zz_3667_;
  wire                _zz_3668_;
  wire                _zz_3669_;
  wire                _zz_3670_;
  wire       [31:0]   _zz_3671_;
  wire       [15:0]   _zz_3672_;
  wire       [15:0]   _zz_3673_;
  wire       [5:0]    _zz_3674_;
  wire       [63:0]   _zz_3675_;
  wire                _zz_3676_;
  wire                _zz_3677_;
  wire                _zz_3678_;
  wire                _zz_3679_;
  wire                _zz_3680_;
  wire                _zz_3681_;
  wire                _zz_3682_;
  wire                _zz_3683_;
  wire                _zz_3684_;
  wire                _zz_3685_;
  wire                _zz_3686_;
  wire                _zz_3687_;
  wire                _zz_3688_;
  wire                _zz_3689_;
  wire                _zz_3690_;
  wire                _zz_3691_;
  wire                _zz_3692_;
  wire                _zz_3693_;
  wire                _zz_3694_;
  wire                _zz_3695_;
  wire                _zz_3696_;
  wire                _zz_3697_;
  wire                _zz_3698_;
  wire                _zz_3699_;
  wire                _zz_3700_;
  wire                _zz_3701_;
  wire                _zz_3702_;
  wire                _zz_3703_;
  wire                _zz_3704_;
  wire                _zz_3705_;
  wire                _zz_3706_;
  wire                _zz_3707_;
  wire                _zz_3708_;
  wire                _zz_3709_;
  wire                _zz_3710_;
  wire                _zz_3711_;
  wire                _zz_3712_;
  wire                _zz_3713_;
  wire                _zz_3714_;
  wire                _zz_3715_;
  wire                _zz_3716_;
  wire                _zz_3717_;
  wire                _zz_3718_;
  wire                _zz_3719_;
  wire                _zz_3720_;
  wire                _zz_3721_;
  wire                _zz_3722_;
  wire                _zz_3723_;
  wire                _zz_3724_;
  wire                _zz_3725_;
  wire                _zz_3726_;
  wire                _zz_3727_;
  wire                _zz_3728_;
  wire                _zz_3729_;
  wire                _zz_3730_;
  wire                _zz_3731_;
  wire                _zz_3732_;
  wire                _zz_3733_;
  wire                _zz_3734_;
  wire                _zz_3735_;
  wire                _zz_3736_;
  wire                _zz_3737_;
  wire                _zz_3738_;
  wire                _zz_3739_;
  wire       [31:0]   _zz_3740_;
  wire       [15:0]   _zz_3741_;
  wire       [15:0]   _zz_3742_;
  wire       [5:0]    _zz_3743_;
  wire       [63:0]   _zz_3744_;
  wire                _zz_3745_;
  wire                _zz_3746_;
  wire                _zz_3747_;
  wire                _zz_3748_;
  wire                _zz_3749_;
  wire                _zz_3750_;
  wire                _zz_3751_;
  wire                _zz_3752_;
  wire                _zz_3753_;
  wire                _zz_3754_;
  wire                _zz_3755_;
  wire                _zz_3756_;
  wire                _zz_3757_;
  wire                _zz_3758_;
  wire                _zz_3759_;
  wire                _zz_3760_;
  wire                _zz_3761_;
  wire                _zz_3762_;
  wire                _zz_3763_;
  wire                _zz_3764_;
  wire                _zz_3765_;
  wire                _zz_3766_;
  wire                _zz_3767_;
  wire                _zz_3768_;
  wire                _zz_3769_;
  wire                _zz_3770_;
  wire                _zz_3771_;
  wire                _zz_3772_;
  wire                _zz_3773_;
  wire                _zz_3774_;
  wire                _zz_3775_;
  wire                _zz_3776_;
  wire                _zz_3777_;
  wire                _zz_3778_;
  wire                _zz_3779_;
  wire                _zz_3780_;
  wire                _zz_3781_;
  wire                _zz_3782_;
  wire                _zz_3783_;
  wire                _zz_3784_;
  wire                _zz_3785_;
  wire                _zz_3786_;
  wire                _zz_3787_;
  wire                _zz_3788_;
  wire                _zz_3789_;
  wire                _zz_3790_;
  wire                _zz_3791_;
  wire                _zz_3792_;
  wire                _zz_3793_;
  wire                _zz_3794_;
  wire                _zz_3795_;
  wire                _zz_3796_;
  wire                _zz_3797_;
  wire                _zz_3798_;
  wire                _zz_3799_;
  wire                _zz_3800_;
  wire                _zz_3801_;
  wire                _zz_3802_;
  wire                _zz_3803_;
  wire                _zz_3804_;
  wire                _zz_3805_;
  wire                _zz_3806_;
  wire                _zz_3807_;
  wire                _zz_3808_;
  wire       [31:0]   _zz_3809_;
  wire       [15:0]   _zz_3810_;
  wire       [15:0]   _zz_3811_;
  wire       [5:0]    _zz_3812_;
  wire       [63:0]   _zz_3813_;
  wire                _zz_3814_;
  wire                _zz_3815_;
  wire                _zz_3816_;
  wire                _zz_3817_;
  wire                _zz_3818_;
  wire                _zz_3819_;
  wire                _zz_3820_;
  wire                _zz_3821_;
  wire                _zz_3822_;
  wire                _zz_3823_;
  wire                _zz_3824_;
  wire                _zz_3825_;
  wire                _zz_3826_;
  wire                _zz_3827_;
  wire                _zz_3828_;
  wire                _zz_3829_;
  wire                _zz_3830_;
  wire                _zz_3831_;
  wire                _zz_3832_;
  wire                _zz_3833_;
  wire                _zz_3834_;
  wire                _zz_3835_;
  wire                _zz_3836_;
  wire                _zz_3837_;
  wire                _zz_3838_;
  wire                _zz_3839_;
  wire                _zz_3840_;
  wire                _zz_3841_;
  wire                _zz_3842_;
  wire                _zz_3843_;
  wire                _zz_3844_;
  wire                _zz_3845_;
  wire                _zz_3846_;
  wire                _zz_3847_;
  wire                _zz_3848_;
  wire                _zz_3849_;
  wire                _zz_3850_;
  wire                _zz_3851_;
  wire                _zz_3852_;
  wire                _zz_3853_;
  wire                _zz_3854_;
  wire                _zz_3855_;
  wire                _zz_3856_;
  wire                _zz_3857_;
  wire                _zz_3858_;
  wire                _zz_3859_;
  wire                _zz_3860_;
  wire                _zz_3861_;
  wire                _zz_3862_;
  wire                _zz_3863_;
  wire                _zz_3864_;
  wire                _zz_3865_;
  wire                _zz_3866_;
  wire                _zz_3867_;
  wire                _zz_3868_;
  wire                _zz_3869_;
  wire                _zz_3870_;
  wire                _zz_3871_;
  wire                _zz_3872_;
  wire                _zz_3873_;
  wire                _zz_3874_;
  wire                _zz_3875_;
  wire                _zz_3876_;
  wire                _zz_3877_;
  wire       [31:0]   _zz_3878_;
  wire       [15:0]   _zz_3879_;
  wire       [15:0]   _zz_3880_;
  wire       [5:0]    _zz_3881_;
  wire       [63:0]   _zz_3882_;
  wire                _zz_3883_;
  wire                _zz_3884_;
  wire                _zz_3885_;
  wire                _zz_3886_;
  wire                _zz_3887_;
  wire                _zz_3888_;
  wire                _zz_3889_;
  wire                _zz_3890_;
  wire                _zz_3891_;
  wire                _zz_3892_;
  wire                _zz_3893_;
  wire                _zz_3894_;
  wire                _zz_3895_;
  wire                _zz_3896_;
  wire                _zz_3897_;
  wire                _zz_3898_;
  wire                _zz_3899_;
  wire                _zz_3900_;
  wire                _zz_3901_;
  wire                _zz_3902_;
  wire                _zz_3903_;
  wire                _zz_3904_;
  wire                _zz_3905_;
  wire                _zz_3906_;
  wire                _zz_3907_;
  wire                _zz_3908_;
  wire                _zz_3909_;
  wire                _zz_3910_;
  wire                _zz_3911_;
  wire                _zz_3912_;
  wire                _zz_3913_;
  wire                _zz_3914_;
  wire                _zz_3915_;
  wire                _zz_3916_;
  wire                _zz_3917_;
  wire                _zz_3918_;
  wire                _zz_3919_;
  wire                _zz_3920_;
  wire                _zz_3921_;
  wire                _zz_3922_;
  wire                _zz_3923_;
  wire                _zz_3924_;
  wire                _zz_3925_;
  wire                _zz_3926_;
  wire                _zz_3927_;
  wire                _zz_3928_;
  wire                _zz_3929_;
  wire                _zz_3930_;
  wire                _zz_3931_;
  wire                _zz_3932_;
  wire                _zz_3933_;
  wire                _zz_3934_;
  wire                _zz_3935_;
  wire                _zz_3936_;
  wire                _zz_3937_;
  wire                _zz_3938_;
  wire                _zz_3939_;
  wire                _zz_3940_;
  wire                _zz_3941_;
  wire                _zz_3942_;
  wire                _zz_3943_;
  wire                _zz_3944_;
  wire                _zz_3945_;
  wire                _zz_3946_;
  wire       [31:0]   _zz_3947_;
  wire       [15:0]   _zz_3948_;
  wire       [15:0]   _zz_3949_;
  wire       [5:0]    _zz_3950_;
  wire       [63:0]   _zz_3951_;
  wire                _zz_3952_;
  wire                _zz_3953_;
  wire                _zz_3954_;
  wire                _zz_3955_;
  wire                _zz_3956_;
  wire                _zz_3957_;
  wire                _zz_3958_;
  wire                _zz_3959_;
  wire                _zz_3960_;
  wire                _zz_3961_;
  wire                _zz_3962_;
  wire                _zz_3963_;
  wire                _zz_3964_;
  wire                _zz_3965_;
  wire                _zz_3966_;
  wire                _zz_3967_;
  wire                _zz_3968_;
  wire                _zz_3969_;
  wire                _zz_3970_;
  wire                _zz_3971_;
  wire                _zz_3972_;
  wire                _zz_3973_;
  wire                _zz_3974_;
  wire                _zz_3975_;
  wire                _zz_3976_;
  wire                _zz_3977_;
  wire                _zz_3978_;
  wire                _zz_3979_;
  wire                _zz_3980_;
  wire                _zz_3981_;
  wire                _zz_3982_;
  wire                _zz_3983_;
  wire                _zz_3984_;
  wire                _zz_3985_;
  wire                _zz_3986_;
  wire                _zz_3987_;
  wire                _zz_3988_;
  wire                _zz_3989_;
  wire                _zz_3990_;
  wire                _zz_3991_;
  wire                _zz_3992_;
  wire                _zz_3993_;
  wire                _zz_3994_;
  wire                _zz_3995_;
  wire                _zz_3996_;
  wire                _zz_3997_;
  wire                _zz_3998_;
  wire                _zz_3999_;
  wire                _zz_4000_;
  wire                _zz_4001_;
  wire                _zz_4002_;
  wire                _zz_4003_;
  wire                _zz_4004_;
  wire                _zz_4005_;
  wire                _zz_4006_;
  wire                _zz_4007_;
  wire                _zz_4008_;
  wire                _zz_4009_;
  wire                _zz_4010_;
  wire                _zz_4011_;
  wire                _zz_4012_;
  wire                _zz_4013_;
  wire                _zz_4014_;
  wire                _zz_4015_;
  wire       [31:0]   _zz_4016_;
  wire       [15:0]   _zz_4017_;
  wire       [15:0]   _zz_4018_;
  wire       [5:0]    _zz_4019_;
  wire       [63:0]   _zz_4020_;
  wire                _zz_4021_;
  wire                _zz_4022_;
  wire                _zz_4023_;
  wire                _zz_4024_;
  wire                _zz_4025_;
  wire                _zz_4026_;
  wire                _zz_4027_;
  wire                _zz_4028_;
  wire                _zz_4029_;
  wire                _zz_4030_;
  wire                _zz_4031_;
  wire                _zz_4032_;
  wire                _zz_4033_;
  wire                _zz_4034_;
  wire                _zz_4035_;
  wire                _zz_4036_;
  wire                _zz_4037_;
  wire                _zz_4038_;
  wire                _zz_4039_;
  wire                _zz_4040_;
  wire                _zz_4041_;
  wire                _zz_4042_;
  wire                _zz_4043_;
  wire                _zz_4044_;
  wire                _zz_4045_;
  wire                _zz_4046_;
  wire                _zz_4047_;
  wire                _zz_4048_;
  wire                _zz_4049_;
  wire                _zz_4050_;
  wire                _zz_4051_;
  wire                _zz_4052_;
  wire                _zz_4053_;
  wire                _zz_4054_;
  wire                _zz_4055_;
  wire                _zz_4056_;
  wire                _zz_4057_;
  wire                _zz_4058_;
  wire                _zz_4059_;
  wire                _zz_4060_;
  wire                _zz_4061_;
  wire                _zz_4062_;
  wire                _zz_4063_;
  wire                _zz_4064_;
  wire                _zz_4065_;
  wire                _zz_4066_;
  wire                _zz_4067_;
  wire                _zz_4068_;
  wire                _zz_4069_;
  wire                _zz_4070_;
  wire                _zz_4071_;
  wire                _zz_4072_;
  wire                _zz_4073_;
  wire                _zz_4074_;
  wire                _zz_4075_;
  wire                _zz_4076_;
  wire                _zz_4077_;
  wire                _zz_4078_;
  wire                _zz_4079_;
  wire                _zz_4080_;
  wire                _zz_4081_;
  wire                _zz_4082_;
  wire                _zz_4083_;
  wire                _zz_4084_;
  wire       [31:0]   _zz_4085_;
  wire       [15:0]   _zz_4086_;
  wire       [15:0]   _zz_4087_;
  wire       [5:0]    _zz_4088_;
  wire       [63:0]   _zz_4089_;
  wire                _zz_4090_;
  wire                _zz_4091_;
  wire                _zz_4092_;
  wire                _zz_4093_;
  wire                _zz_4094_;
  wire                _zz_4095_;
  wire                _zz_4096_;
  wire                _zz_4097_;
  wire                _zz_4098_;
  wire                _zz_4099_;
  wire                _zz_4100_;
  wire                _zz_4101_;
  wire                _zz_4102_;
  wire                _zz_4103_;
  wire                _zz_4104_;
  wire                _zz_4105_;
  wire                _zz_4106_;
  wire                _zz_4107_;
  wire                _zz_4108_;
  wire                _zz_4109_;
  wire                _zz_4110_;
  wire                _zz_4111_;
  wire                _zz_4112_;
  wire                _zz_4113_;
  wire                _zz_4114_;
  wire                _zz_4115_;
  wire                _zz_4116_;
  wire                _zz_4117_;
  wire                _zz_4118_;
  wire                _zz_4119_;
  wire                _zz_4120_;
  wire                _zz_4121_;
  wire                _zz_4122_;
  wire                _zz_4123_;
  wire                _zz_4124_;
  wire                _zz_4125_;
  wire                _zz_4126_;
  wire                _zz_4127_;
  wire                _zz_4128_;
  wire                _zz_4129_;
  wire                _zz_4130_;
  wire                _zz_4131_;
  wire                _zz_4132_;
  wire                _zz_4133_;
  wire                _zz_4134_;
  wire                _zz_4135_;
  wire                _zz_4136_;
  wire                _zz_4137_;
  wire                _zz_4138_;
  wire                _zz_4139_;
  wire                _zz_4140_;
  wire                _zz_4141_;
  wire                _zz_4142_;
  wire                _zz_4143_;
  wire                _zz_4144_;
  wire                _zz_4145_;
  wire                _zz_4146_;
  wire                _zz_4147_;
  wire                _zz_4148_;
  wire                _zz_4149_;
  wire                _zz_4150_;
  wire                _zz_4151_;
  wire                _zz_4152_;
  wire                _zz_4153_;
  wire       [31:0]   _zz_4154_;
  wire       [15:0]   _zz_4155_;
  wire       [15:0]   _zz_4156_;
  wire       [5:0]    _zz_4157_;
  wire       [63:0]   _zz_4158_;
  wire                _zz_4159_;
  wire                _zz_4160_;
  wire                _zz_4161_;
  wire                _zz_4162_;
  wire                _zz_4163_;
  wire                _zz_4164_;
  wire                _zz_4165_;
  wire                _zz_4166_;
  wire                _zz_4167_;
  wire                _zz_4168_;
  wire                _zz_4169_;
  wire                _zz_4170_;
  wire                _zz_4171_;
  wire                _zz_4172_;
  wire                _zz_4173_;
  wire                _zz_4174_;
  wire                _zz_4175_;
  wire                _zz_4176_;
  wire                _zz_4177_;
  wire                _zz_4178_;
  wire                _zz_4179_;
  wire                _zz_4180_;
  wire                _zz_4181_;
  wire                _zz_4182_;
  wire                _zz_4183_;
  wire                _zz_4184_;
  wire                _zz_4185_;
  wire                _zz_4186_;
  wire                _zz_4187_;
  wire                _zz_4188_;
  wire                _zz_4189_;
  wire                _zz_4190_;
  wire                _zz_4191_;
  wire                _zz_4192_;
  wire                _zz_4193_;
  wire                _zz_4194_;
  wire                _zz_4195_;
  wire                _zz_4196_;
  wire                _zz_4197_;
  wire                _zz_4198_;
  wire                _zz_4199_;
  wire                _zz_4200_;
  wire                _zz_4201_;
  wire                _zz_4202_;
  wire                _zz_4203_;
  wire                _zz_4204_;
  wire                _zz_4205_;
  wire                _zz_4206_;
  wire                _zz_4207_;
  wire                _zz_4208_;
  wire                _zz_4209_;
  wire                _zz_4210_;
  wire                _zz_4211_;
  wire                _zz_4212_;
  wire                _zz_4213_;
  wire                _zz_4214_;
  wire                _zz_4215_;
  wire                _zz_4216_;
  wire                _zz_4217_;
  wire                _zz_4218_;
  wire                _zz_4219_;
  wire                _zz_4220_;
  wire                _zz_4221_;
  wire                _zz_4222_;
  wire       [31:0]   _zz_4223_;
  wire       [15:0]   _zz_4224_;
  wire       [15:0]   _zz_4225_;
  wire       [5:0]    _zz_4226_;
  wire       [63:0]   _zz_4227_;
  wire                _zz_4228_;
  wire                _zz_4229_;
  wire                _zz_4230_;
  wire                _zz_4231_;
  wire                _zz_4232_;
  wire                _zz_4233_;
  wire                _zz_4234_;
  wire                _zz_4235_;
  wire                _zz_4236_;
  wire                _zz_4237_;
  wire                _zz_4238_;
  wire                _zz_4239_;
  wire                _zz_4240_;
  wire                _zz_4241_;
  wire                _zz_4242_;
  wire                _zz_4243_;
  wire                _zz_4244_;
  wire                _zz_4245_;
  wire                _zz_4246_;
  wire                _zz_4247_;
  wire                _zz_4248_;
  wire                _zz_4249_;
  wire                _zz_4250_;
  wire                _zz_4251_;
  wire                _zz_4252_;
  wire                _zz_4253_;
  wire                _zz_4254_;
  wire                _zz_4255_;
  wire                _zz_4256_;
  wire                _zz_4257_;
  wire                _zz_4258_;
  wire                _zz_4259_;
  wire                _zz_4260_;
  wire                _zz_4261_;
  wire                _zz_4262_;
  wire                _zz_4263_;
  wire                _zz_4264_;
  wire                _zz_4265_;
  wire                _zz_4266_;
  wire                _zz_4267_;
  wire                _zz_4268_;
  wire                _zz_4269_;
  wire                _zz_4270_;
  wire                _zz_4271_;
  wire                _zz_4272_;
  wire                _zz_4273_;
  wire                _zz_4274_;
  wire                _zz_4275_;
  wire                _zz_4276_;
  wire                _zz_4277_;
  wire                _zz_4278_;
  wire                _zz_4279_;
  wire                _zz_4280_;
  wire                _zz_4281_;
  wire                _zz_4282_;
  wire                _zz_4283_;
  wire                _zz_4284_;
  wire                _zz_4285_;
  wire                _zz_4286_;
  wire                _zz_4287_;
  wire                _zz_4288_;
  wire                _zz_4289_;
  wire                _zz_4290_;
  wire                _zz_4291_;
  wire       [31:0]   _zz_4292_;
  wire       [15:0]   _zz_4293_;
  wire       [15:0]   _zz_4294_;
  wire       [5:0]    _zz_4295_;
  wire       [63:0]   _zz_4296_;
  wire                _zz_4297_;
  wire                _zz_4298_;
  wire                _zz_4299_;
  wire                _zz_4300_;
  wire                _zz_4301_;
  wire                _zz_4302_;
  wire                _zz_4303_;
  wire                _zz_4304_;
  wire                _zz_4305_;
  wire                _zz_4306_;
  wire                _zz_4307_;
  wire                _zz_4308_;
  wire                _zz_4309_;
  wire                _zz_4310_;
  wire                _zz_4311_;
  wire                _zz_4312_;
  wire                _zz_4313_;
  wire                _zz_4314_;
  wire                _zz_4315_;
  wire                _zz_4316_;
  wire                _zz_4317_;
  wire                _zz_4318_;
  wire                _zz_4319_;
  wire                _zz_4320_;
  wire                _zz_4321_;
  wire                _zz_4322_;
  wire                _zz_4323_;
  wire                _zz_4324_;
  wire                _zz_4325_;
  wire                _zz_4326_;
  wire                _zz_4327_;
  wire                _zz_4328_;
  wire                _zz_4329_;
  wire                _zz_4330_;
  wire                _zz_4331_;
  wire                _zz_4332_;
  wire                _zz_4333_;
  wire                _zz_4334_;
  wire                _zz_4335_;
  wire                _zz_4336_;
  wire                _zz_4337_;
  wire                _zz_4338_;
  wire                _zz_4339_;
  wire                _zz_4340_;
  wire                _zz_4341_;
  wire                _zz_4342_;
  wire                _zz_4343_;
  wire                _zz_4344_;
  wire                _zz_4345_;
  wire                _zz_4346_;
  wire                _zz_4347_;
  wire                _zz_4348_;
  wire                _zz_4349_;
  wire                _zz_4350_;
  wire                _zz_4351_;
  wire                _zz_4352_;
  wire                _zz_4353_;
  wire                _zz_4354_;
  wire                _zz_4355_;
  wire                _zz_4356_;
  wire                _zz_4357_;
  wire                _zz_4358_;
  wire                _zz_4359_;
  wire                _zz_4360_;
  wire       [31:0]   _zz_4361_;
  wire       [15:0]   _zz_4362_;
  wire       [15:0]   _zz_4363_;
  wire       [5:0]    _zz_4364_;
  wire       [63:0]   _zz_4365_;
  wire                _zz_4366_;
  wire                _zz_4367_;
  wire                _zz_4368_;
  wire                _zz_4369_;
  wire                _zz_4370_;
  wire                _zz_4371_;
  wire                _zz_4372_;
  wire                _zz_4373_;
  wire                _zz_4374_;
  wire                _zz_4375_;
  wire                _zz_4376_;
  wire                _zz_4377_;
  wire                _zz_4378_;
  wire                _zz_4379_;
  wire                _zz_4380_;
  wire                _zz_4381_;
  wire                _zz_4382_;
  wire                _zz_4383_;
  wire                _zz_4384_;
  wire                _zz_4385_;
  wire                _zz_4386_;
  wire                _zz_4387_;
  wire                _zz_4388_;
  wire                _zz_4389_;
  wire                _zz_4390_;
  wire                _zz_4391_;
  wire                _zz_4392_;
  wire                _zz_4393_;
  wire                _zz_4394_;
  wire                _zz_4395_;
  wire                _zz_4396_;
  wire                _zz_4397_;
  wire                _zz_4398_;
  wire                _zz_4399_;
  wire                _zz_4400_;
  wire                _zz_4401_;
  wire                _zz_4402_;
  wire                _zz_4403_;
  wire                _zz_4404_;
  wire                _zz_4405_;
  wire                _zz_4406_;
  wire                _zz_4407_;
  wire                _zz_4408_;
  wire                _zz_4409_;
  wire                _zz_4410_;
  wire                _zz_4411_;
  wire                _zz_4412_;
  wire                _zz_4413_;
  wire                _zz_4414_;
  wire                _zz_4415_;
  wire                _zz_4416_;
  wire                _zz_4417_;
  wire                _zz_4418_;
  wire                _zz_4419_;
  wire                _zz_4420_;
  wire                _zz_4421_;
  wire                _zz_4422_;
  wire                _zz_4423_;
  wire                _zz_4424_;
  wire                _zz_4425_;
  wire                _zz_4426_;
  wire                _zz_4427_;
  wire                _zz_4428_;
  wire                _zz_4429_;
  wire       [31:0]   _zz_4430_;
  wire       [15:0]   _zz_4431_;
  wire       [15:0]   _zz_4432_;

  assign _zz_4562_ = _zz_13_[11 : 0];
  assign _zz_4563_ = _zz_4562_;
  assign _zz_4564_ = {11'd0, Axi4Incr_sizeValue};
  assign _zz_4565_ = transfer_done;
  assign _zz_4566_ = (load_data_area_current_addr - 32'h0);
  assign _zz_4567_ = (load_data_area_current_addr - 32'h00000f00);
  assign _zz_4568_ = (load_data_area_current_addr - 32'h00000b80);
  assign _zz_4569_ = (load_data_area_current_addr - 32'h000009c0);
  assign _zz_4570_ = (load_data_area_current_addr - 32'h00000b00);
  assign _zz_4571_ = (load_data_area_current_addr - 32'h000005c0);
  assign _zz_4572_ = (load_data_area_current_addr - 32'h00000c80);
  assign _zz_4573_ = (load_data_area_current_addr - 32'h00000a40);
  assign _zz_4574_ = (load_data_area_current_addr - 32'h000002c0);
  assign _zz_4575_ = (load_data_area_current_addr - 32'h00000f80);
  assign _zz_4576_ = (load_data_area_current_addr - 32'h00000780);
  assign _zz_4577_ = (load_data_area_current_addr - 32'h00000580);
  assign _zz_4578_ = (load_data_area_current_addr - 32'h00000500);
  assign _zz_4579_ = (load_data_area_current_addr - 32'h00000880);
  assign _zz_4580_ = (load_data_area_current_addr - 32'h00000180);
  assign _zz_4581_ = (load_data_area_current_addr - 32'h00000200);
  assign _zz_4582_ = (load_data_area_current_addr - 32'h000006c0);
  assign _zz_4583_ = (load_data_area_current_addr - 32'h000004c0);
  assign _zz_4584_ = (load_data_area_current_addr - 32'h00000c40);
  assign _zz_4585_ = (load_data_area_current_addr - 32'h000001c0);
  assign _zz_4586_ = (load_data_area_current_addr - 32'h00000e80);
  assign _zz_4587_ = (load_data_area_current_addr - 32'h00000700);
  assign _zz_4588_ = (load_data_area_current_addr - 32'h00000d80);
  assign _zz_4589_ = (load_data_area_current_addr - 32'h00000ac0);
  assign _zz_4590_ = (load_data_area_current_addr - 32'h00000380);
  assign _zz_4591_ = (load_data_area_current_addr - 32'h00000800);
  assign _zz_4592_ = (load_data_area_current_addr - 32'h00000f40);
  assign _zz_4593_ = (load_data_area_current_addr - 32'h00000680);
  assign _zz_4594_ = (load_data_area_current_addr - 32'h00000400);
  assign _zz_4595_ = (load_data_area_current_addr - 32'h00000980);
  assign _zz_4596_ = (load_data_area_current_addr - 32'h00000e00);
  assign _zz_4597_ = (load_data_area_current_addr - 32'h00000e40);
  assign _zz_4598_ = (load_data_area_current_addr - 32'h00000600);
  assign _zz_4599_ = (load_data_area_current_addr - 32'h00000040);
  assign _zz_4600_ = (load_data_area_current_addr - 32'h00000d00);
  assign _zz_4601_ = (load_data_area_current_addr - 32'h00000240);
  assign _zz_4602_ = (load_data_area_current_addr - 32'h00000a00);
  assign _zz_4603_ = (load_data_area_current_addr - 32'h00000640);
  assign _zz_4604_ = (load_data_area_current_addr - 32'h00000080);
  assign _zz_4605_ = (load_data_area_current_addr - 32'h00000840);
  assign _zz_4606_ = (load_data_area_current_addr - 32'h00000140);
  assign _zz_4607_ = (load_data_area_current_addr - 32'h000000c0);
  assign _zz_4608_ = (load_data_area_current_addr - 32'h00000340);
  assign _zz_4609_ = (load_data_area_current_addr - 32'h00000dc0);
  assign _zz_4610_ = (load_data_area_current_addr - 32'h00000d40);
  assign _zz_4611_ = (load_data_area_current_addr - 32'h00000280);
  assign _zz_4612_ = (load_data_area_current_addr - 32'h00000740);
  assign _zz_4613_ = (load_data_area_current_addr - 32'h00000ec0);
  assign _zz_4614_ = (load_data_area_current_addr - 32'h00000b40);
  assign _zz_4615_ = (load_data_area_current_addr - 32'h00000100);
  assign _zz_4616_ = (load_data_area_current_addr - 32'h00000cc0);
  assign _zz_4617_ = (load_data_area_current_addr - 32'h00000440);
  assign _zz_4618_ = (load_data_area_current_addr - 32'h00000540);
  assign _zz_4619_ = (load_data_area_current_addr - 32'h000008c0);
  assign _zz_4620_ = (load_data_area_current_addr - 32'h00000a80);
  assign _zz_4621_ = (load_data_area_current_addr - 32'h000007c0);
  assign _zz_4622_ = (load_data_area_current_addr - 32'h00000c00);
  assign _zz_4623_ = (load_data_area_current_addr - 32'h00000940);
  assign _zz_4624_ = (load_data_area_current_addr - 32'h00000300);
  assign _zz_4625_ = (load_data_area_current_addr - 32'h00000900);
  assign _zz_4626_ = (load_data_area_current_addr - 32'h00000fc0);
  assign _zz_4627_ = (load_data_area_current_addr - 32'h000003c0);
  assign _zz_4628_ = (load_data_area_current_addr - 32'h00000bc0);
  assign _zz_4629_ = (load_data_area_current_addr - 32'h00000480);
  always @(*) begin
    case(Axi4Incr_wrapCase)
      2'b00 : begin
        _zz_4433_ = {Axi4Incr_base[11 : 1],Axi4Incr_baseIncr[0 : 0]};
      end
      2'b01 : begin
        _zz_4433_ = {Axi4Incr_base[11 : 2],Axi4Incr_baseIncr[1 : 0]};
      end
      2'b10 : begin
        _zz_4433_ = {Axi4Incr_base[11 : 3],Axi4Incr_baseIncr[2 : 0]};
      end
      default : begin
        _zz_4433_ = {Axi4Incr_base[11 : 4],Axi4Incr_baseIncr[3 : 0]};
      end
    endcase
  end

  always @(*) begin
    case(_zz_17_)
      6'b000000 : begin
        _zz_4434_ = int_reg_array_0_0_imag;
        _zz_4435_ = int_reg_array_0_0_real;
      end
      6'b000001 : begin
        _zz_4434_ = int_reg_array_0_1_imag;
        _zz_4435_ = int_reg_array_0_1_real;
      end
      6'b000010 : begin
        _zz_4434_ = int_reg_array_0_2_imag;
        _zz_4435_ = int_reg_array_0_2_real;
      end
      6'b000011 : begin
        _zz_4434_ = int_reg_array_0_3_imag;
        _zz_4435_ = int_reg_array_0_3_real;
      end
      6'b000100 : begin
        _zz_4434_ = int_reg_array_0_4_imag;
        _zz_4435_ = int_reg_array_0_4_real;
      end
      6'b000101 : begin
        _zz_4434_ = int_reg_array_0_5_imag;
        _zz_4435_ = int_reg_array_0_5_real;
      end
      6'b000110 : begin
        _zz_4434_ = int_reg_array_0_6_imag;
        _zz_4435_ = int_reg_array_0_6_real;
      end
      6'b000111 : begin
        _zz_4434_ = int_reg_array_0_7_imag;
        _zz_4435_ = int_reg_array_0_7_real;
      end
      6'b001000 : begin
        _zz_4434_ = int_reg_array_0_8_imag;
        _zz_4435_ = int_reg_array_0_8_real;
      end
      6'b001001 : begin
        _zz_4434_ = int_reg_array_0_9_imag;
        _zz_4435_ = int_reg_array_0_9_real;
      end
      6'b001010 : begin
        _zz_4434_ = int_reg_array_0_10_imag;
        _zz_4435_ = int_reg_array_0_10_real;
      end
      6'b001011 : begin
        _zz_4434_ = int_reg_array_0_11_imag;
        _zz_4435_ = int_reg_array_0_11_real;
      end
      6'b001100 : begin
        _zz_4434_ = int_reg_array_0_12_imag;
        _zz_4435_ = int_reg_array_0_12_real;
      end
      6'b001101 : begin
        _zz_4434_ = int_reg_array_0_13_imag;
        _zz_4435_ = int_reg_array_0_13_real;
      end
      6'b001110 : begin
        _zz_4434_ = int_reg_array_0_14_imag;
        _zz_4435_ = int_reg_array_0_14_real;
      end
      6'b001111 : begin
        _zz_4434_ = int_reg_array_0_15_imag;
        _zz_4435_ = int_reg_array_0_15_real;
      end
      6'b010000 : begin
        _zz_4434_ = int_reg_array_0_16_imag;
        _zz_4435_ = int_reg_array_0_16_real;
      end
      6'b010001 : begin
        _zz_4434_ = int_reg_array_0_17_imag;
        _zz_4435_ = int_reg_array_0_17_real;
      end
      6'b010010 : begin
        _zz_4434_ = int_reg_array_0_18_imag;
        _zz_4435_ = int_reg_array_0_18_real;
      end
      6'b010011 : begin
        _zz_4434_ = int_reg_array_0_19_imag;
        _zz_4435_ = int_reg_array_0_19_real;
      end
      6'b010100 : begin
        _zz_4434_ = int_reg_array_0_20_imag;
        _zz_4435_ = int_reg_array_0_20_real;
      end
      6'b010101 : begin
        _zz_4434_ = int_reg_array_0_21_imag;
        _zz_4435_ = int_reg_array_0_21_real;
      end
      6'b010110 : begin
        _zz_4434_ = int_reg_array_0_22_imag;
        _zz_4435_ = int_reg_array_0_22_real;
      end
      6'b010111 : begin
        _zz_4434_ = int_reg_array_0_23_imag;
        _zz_4435_ = int_reg_array_0_23_real;
      end
      6'b011000 : begin
        _zz_4434_ = int_reg_array_0_24_imag;
        _zz_4435_ = int_reg_array_0_24_real;
      end
      6'b011001 : begin
        _zz_4434_ = int_reg_array_0_25_imag;
        _zz_4435_ = int_reg_array_0_25_real;
      end
      6'b011010 : begin
        _zz_4434_ = int_reg_array_0_26_imag;
        _zz_4435_ = int_reg_array_0_26_real;
      end
      6'b011011 : begin
        _zz_4434_ = int_reg_array_0_27_imag;
        _zz_4435_ = int_reg_array_0_27_real;
      end
      6'b011100 : begin
        _zz_4434_ = int_reg_array_0_28_imag;
        _zz_4435_ = int_reg_array_0_28_real;
      end
      6'b011101 : begin
        _zz_4434_ = int_reg_array_0_29_imag;
        _zz_4435_ = int_reg_array_0_29_real;
      end
      6'b011110 : begin
        _zz_4434_ = int_reg_array_0_30_imag;
        _zz_4435_ = int_reg_array_0_30_real;
      end
      6'b011111 : begin
        _zz_4434_ = int_reg_array_0_31_imag;
        _zz_4435_ = int_reg_array_0_31_real;
      end
      6'b100000 : begin
        _zz_4434_ = int_reg_array_0_32_imag;
        _zz_4435_ = int_reg_array_0_32_real;
      end
      6'b100001 : begin
        _zz_4434_ = int_reg_array_0_33_imag;
        _zz_4435_ = int_reg_array_0_33_real;
      end
      6'b100010 : begin
        _zz_4434_ = int_reg_array_0_34_imag;
        _zz_4435_ = int_reg_array_0_34_real;
      end
      6'b100011 : begin
        _zz_4434_ = int_reg_array_0_35_imag;
        _zz_4435_ = int_reg_array_0_35_real;
      end
      6'b100100 : begin
        _zz_4434_ = int_reg_array_0_36_imag;
        _zz_4435_ = int_reg_array_0_36_real;
      end
      6'b100101 : begin
        _zz_4434_ = int_reg_array_0_37_imag;
        _zz_4435_ = int_reg_array_0_37_real;
      end
      6'b100110 : begin
        _zz_4434_ = int_reg_array_0_38_imag;
        _zz_4435_ = int_reg_array_0_38_real;
      end
      6'b100111 : begin
        _zz_4434_ = int_reg_array_0_39_imag;
        _zz_4435_ = int_reg_array_0_39_real;
      end
      6'b101000 : begin
        _zz_4434_ = int_reg_array_0_40_imag;
        _zz_4435_ = int_reg_array_0_40_real;
      end
      6'b101001 : begin
        _zz_4434_ = int_reg_array_0_41_imag;
        _zz_4435_ = int_reg_array_0_41_real;
      end
      6'b101010 : begin
        _zz_4434_ = int_reg_array_0_42_imag;
        _zz_4435_ = int_reg_array_0_42_real;
      end
      6'b101011 : begin
        _zz_4434_ = int_reg_array_0_43_imag;
        _zz_4435_ = int_reg_array_0_43_real;
      end
      6'b101100 : begin
        _zz_4434_ = int_reg_array_0_44_imag;
        _zz_4435_ = int_reg_array_0_44_real;
      end
      6'b101101 : begin
        _zz_4434_ = int_reg_array_0_45_imag;
        _zz_4435_ = int_reg_array_0_45_real;
      end
      6'b101110 : begin
        _zz_4434_ = int_reg_array_0_46_imag;
        _zz_4435_ = int_reg_array_0_46_real;
      end
      6'b101111 : begin
        _zz_4434_ = int_reg_array_0_47_imag;
        _zz_4435_ = int_reg_array_0_47_real;
      end
      6'b110000 : begin
        _zz_4434_ = int_reg_array_0_48_imag;
        _zz_4435_ = int_reg_array_0_48_real;
      end
      6'b110001 : begin
        _zz_4434_ = int_reg_array_0_49_imag;
        _zz_4435_ = int_reg_array_0_49_real;
      end
      6'b110010 : begin
        _zz_4434_ = int_reg_array_0_50_imag;
        _zz_4435_ = int_reg_array_0_50_real;
      end
      6'b110011 : begin
        _zz_4434_ = int_reg_array_0_51_imag;
        _zz_4435_ = int_reg_array_0_51_real;
      end
      6'b110100 : begin
        _zz_4434_ = int_reg_array_0_52_imag;
        _zz_4435_ = int_reg_array_0_52_real;
      end
      6'b110101 : begin
        _zz_4434_ = int_reg_array_0_53_imag;
        _zz_4435_ = int_reg_array_0_53_real;
      end
      6'b110110 : begin
        _zz_4434_ = int_reg_array_0_54_imag;
        _zz_4435_ = int_reg_array_0_54_real;
      end
      6'b110111 : begin
        _zz_4434_ = int_reg_array_0_55_imag;
        _zz_4435_ = int_reg_array_0_55_real;
      end
      6'b111000 : begin
        _zz_4434_ = int_reg_array_0_56_imag;
        _zz_4435_ = int_reg_array_0_56_real;
      end
      6'b111001 : begin
        _zz_4434_ = int_reg_array_0_57_imag;
        _zz_4435_ = int_reg_array_0_57_real;
      end
      6'b111010 : begin
        _zz_4434_ = int_reg_array_0_58_imag;
        _zz_4435_ = int_reg_array_0_58_real;
      end
      6'b111011 : begin
        _zz_4434_ = int_reg_array_0_59_imag;
        _zz_4435_ = int_reg_array_0_59_real;
      end
      6'b111100 : begin
        _zz_4434_ = int_reg_array_0_60_imag;
        _zz_4435_ = int_reg_array_0_60_real;
      end
      6'b111101 : begin
        _zz_4434_ = int_reg_array_0_61_imag;
        _zz_4435_ = int_reg_array_0_61_real;
      end
      6'b111110 : begin
        _zz_4434_ = int_reg_array_0_62_imag;
        _zz_4435_ = int_reg_array_0_62_real;
      end
      default : begin
        _zz_4434_ = int_reg_array_0_63_imag;
        _zz_4435_ = int_reg_array_0_63_real;
      end
    endcase
  end

  always @(*) begin
    case(_zz_86_)
      6'b000000 : begin
        _zz_4436_ = int_reg_array_1_0_imag;
        _zz_4437_ = int_reg_array_1_0_real;
      end
      6'b000001 : begin
        _zz_4436_ = int_reg_array_1_1_imag;
        _zz_4437_ = int_reg_array_1_1_real;
      end
      6'b000010 : begin
        _zz_4436_ = int_reg_array_1_2_imag;
        _zz_4437_ = int_reg_array_1_2_real;
      end
      6'b000011 : begin
        _zz_4436_ = int_reg_array_1_3_imag;
        _zz_4437_ = int_reg_array_1_3_real;
      end
      6'b000100 : begin
        _zz_4436_ = int_reg_array_1_4_imag;
        _zz_4437_ = int_reg_array_1_4_real;
      end
      6'b000101 : begin
        _zz_4436_ = int_reg_array_1_5_imag;
        _zz_4437_ = int_reg_array_1_5_real;
      end
      6'b000110 : begin
        _zz_4436_ = int_reg_array_1_6_imag;
        _zz_4437_ = int_reg_array_1_6_real;
      end
      6'b000111 : begin
        _zz_4436_ = int_reg_array_1_7_imag;
        _zz_4437_ = int_reg_array_1_7_real;
      end
      6'b001000 : begin
        _zz_4436_ = int_reg_array_1_8_imag;
        _zz_4437_ = int_reg_array_1_8_real;
      end
      6'b001001 : begin
        _zz_4436_ = int_reg_array_1_9_imag;
        _zz_4437_ = int_reg_array_1_9_real;
      end
      6'b001010 : begin
        _zz_4436_ = int_reg_array_1_10_imag;
        _zz_4437_ = int_reg_array_1_10_real;
      end
      6'b001011 : begin
        _zz_4436_ = int_reg_array_1_11_imag;
        _zz_4437_ = int_reg_array_1_11_real;
      end
      6'b001100 : begin
        _zz_4436_ = int_reg_array_1_12_imag;
        _zz_4437_ = int_reg_array_1_12_real;
      end
      6'b001101 : begin
        _zz_4436_ = int_reg_array_1_13_imag;
        _zz_4437_ = int_reg_array_1_13_real;
      end
      6'b001110 : begin
        _zz_4436_ = int_reg_array_1_14_imag;
        _zz_4437_ = int_reg_array_1_14_real;
      end
      6'b001111 : begin
        _zz_4436_ = int_reg_array_1_15_imag;
        _zz_4437_ = int_reg_array_1_15_real;
      end
      6'b010000 : begin
        _zz_4436_ = int_reg_array_1_16_imag;
        _zz_4437_ = int_reg_array_1_16_real;
      end
      6'b010001 : begin
        _zz_4436_ = int_reg_array_1_17_imag;
        _zz_4437_ = int_reg_array_1_17_real;
      end
      6'b010010 : begin
        _zz_4436_ = int_reg_array_1_18_imag;
        _zz_4437_ = int_reg_array_1_18_real;
      end
      6'b010011 : begin
        _zz_4436_ = int_reg_array_1_19_imag;
        _zz_4437_ = int_reg_array_1_19_real;
      end
      6'b010100 : begin
        _zz_4436_ = int_reg_array_1_20_imag;
        _zz_4437_ = int_reg_array_1_20_real;
      end
      6'b010101 : begin
        _zz_4436_ = int_reg_array_1_21_imag;
        _zz_4437_ = int_reg_array_1_21_real;
      end
      6'b010110 : begin
        _zz_4436_ = int_reg_array_1_22_imag;
        _zz_4437_ = int_reg_array_1_22_real;
      end
      6'b010111 : begin
        _zz_4436_ = int_reg_array_1_23_imag;
        _zz_4437_ = int_reg_array_1_23_real;
      end
      6'b011000 : begin
        _zz_4436_ = int_reg_array_1_24_imag;
        _zz_4437_ = int_reg_array_1_24_real;
      end
      6'b011001 : begin
        _zz_4436_ = int_reg_array_1_25_imag;
        _zz_4437_ = int_reg_array_1_25_real;
      end
      6'b011010 : begin
        _zz_4436_ = int_reg_array_1_26_imag;
        _zz_4437_ = int_reg_array_1_26_real;
      end
      6'b011011 : begin
        _zz_4436_ = int_reg_array_1_27_imag;
        _zz_4437_ = int_reg_array_1_27_real;
      end
      6'b011100 : begin
        _zz_4436_ = int_reg_array_1_28_imag;
        _zz_4437_ = int_reg_array_1_28_real;
      end
      6'b011101 : begin
        _zz_4436_ = int_reg_array_1_29_imag;
        _zz_4437_ = int_reg_array_1_29_real;
      end
      6'b011110 : begin
        _zz_4436_ = int_reg_array_1_30_imag;
        _zz_4437_ = int_reg_array_1_30_real;
      end
      6'b011111 : begin
        _zz_4436_ = int_reg_array_1_31_imag;
        _zz_4437_ = int_reg_array_1_31_real;
      end
      6'b100000 : begin
        _zz_4436_ = int_reg_array_1_32_imag;
        _zz_4437_ = int_reg_array_1_32_real;
      end
      6'b100001 : begin
        _zz_4436_ = int_reg_array_1_33_imag;
        _zz_4437_ = int_reg_array_1_33_real;
      end
      6'b100010 : begin
        _zz_4436_ = int_reg_array_1_34_imag;
        _zz_4437_ = int_reg_array_1_34_real;
      end
      6'b100011 : begin
        _zz_4436_ = int_reg_array_1_35_imag;
        _zz_4437_ = int_reg_array_1_35_real;
      end
      6'b100100 : begin
        _zz_4436_ = int_reg_array_1_36_imag;
        _zz_4437_ = int_reg_array_1_36_real;
      end
      6'b100101 : begin
        _zz_4436_ = int_reg_array_1_37_imag;
        _zz_4437_ = int_reg_array_1_37_real;
      end
      6'b100110 : begin
        _zz_4436_ = int_reg_array_1_38_imag;
        _zz_4437_ = int_reg_array_1_38_real;
      end
      6'b100111 : begin
        _zz_4436_ = int_reg_array_1_39_imag;
        _zz_4437_ = int_reg_array_1_39_real;
      end
      6'b101000 : begin
        _zz_4436_ = int_reg_array_1_40_imag;
        _zz_4437_ = int_reg_array_1_40_real;
      end
      6'b101001 : begin
        _zz_4436_ = int_reg_array_1_41_imag;
        _zz_4437_ = int_reg_array_1_41_real;
      end
      6'b101010 : begin
        _zz_4436_ = int_reg_array_1_42_imag;
        _zz_4437_ = int_reg_array_1_42_real;
      end
      6'b101011 : begin
        _zz_4436_ = int_reg_array_1_43_imag;
        _zz_4437_ = int_reg_array_1_43_real;
      end
      6'b101100 : begin
        _zz_4436_ = int_reg_array_1_44_imag;
        _zz_4437_ = int_reg_array_1_44_real;
      end
      6'b101101 : begin
        _zz_4436_ = int_reg_array_1_45_imag;
        _zz_4437_ = int_reg_array_1_45_real;
      end
      6'b101110 : begin
        _zz_4436_ = int_reg_array_1_46_imag;
        _zz_4437_ = int_reg_array_1_46_real;
      end
      6'b101111 : begin
        _zz_4436_ = int_reg_array_1_47_imag;
        _zz_4437_ = int_reg_array_1_47_real;
      end
      6'b110000 : begin
        _zz_4436_ = int_reg_array_1_48_imag;
        _zz_4437_ = int_reg_array_1_48_real;
      end
      6'b110001 : begin
        _zz_4436_ = int_reg_array_1_49_imag;
        _zz_4437_ = int_reg_array_1_49_real;
      end
      6'b110010 : begin
        _zz_4436_ = int_reg_array_1_50_imag;
        _zz_4437_ = int_reg_array_1_50_real;
      end
      6'b110011 : begin
        _zz_4436_ = int_reg_array_1_51_imag;
        _zz_4437_ = int_reg_array_1_51_real;
      end
      6'b110100 : begin
        _zz_4436_ = int_reg_array_1_52_imag;
        _zz_4437_ = int_reg_array_1_52_real;
      end
      6'b110101 : begin
        _zz_4436_ = int_reg_array_1_53_imag;
        _zz_4437_ = int_reg_array_1_53_real;
      end
      6'b110110 : begin
        _zz_4436_ = int_reg_array_1_54_imag;
        _zz_4437_ = int_reg_array_1_54_real;
      end
      6'b110111 : begin
        _zz_4436_ = int_reg_array_1_55_imag;
        _zz_4437_ = int_reg_array_1_55_real;
      end
      6'b111000 : begin
        _zz_4436_ = int_reg_array_1_56_imag;
        _zz_4437_ = int_reg_array_1_56_real;
      end
      6'b111001 : begin
        _zz_4436_ = int_reg_array_1_57_imag;
        _zz_4437_ = int_reg_array_1_57_real;
      end
      6'b111010 : begin
        _zz_4436_ = int_reg_array_1_58_imag;
        _zz_4437_ = int_reg_array_1_58_real;
      end
      6'b111011 : begin
        _zz_4436_ = int_reg_array_1_59_imag;
        _zz_4437_ = int_reg_array_1_59_real;
      end
      6'b111100 : begin
        _zz_4436_ = int_reg_array_1_60_imag;
        _zz_4437_ = int_reg_array_1_60_real;
      end
      6'b111101 : begin
        _zz_4436_ = int_reg_array_1_61_imag;
        _zz_4437_ = int_reg_array_1_61_real;
      end
      6'b111110 : begin
        _zz_4436_ = int_reg_array_1_62_imag;
        _zz_4437_ = int_reg_array_1_62_real;
      end
      default : begin
        _zz_4436_ = int_reg_array_1_63_imag;
        _zz_4437_ = int_reg_array_1_63_real;
      end
    endcase
  end

  always @(*) begin
    case(_zz_155_)
      6'b000000 : begin
        _zz_4438_ = int_reg_array_2_0_imag;
        _zz_4439_ = int_reg_array_2_0_real;
      end
      6'b000001 : begin
        _zz_4438_ = int_reg_array_2_1_imag;
        _zz_4439_ = int_reg_array_2_1_real;
      end
      6'b000010 : begin
        _zz_4438_ = int_reg_array_2_2_imag;
        _zz_4439_ = int_reg_array_2_2_real;
      end
      6'b000011 : begin
        _zz_4438_ = int_reg_array_2_3_imag;
        _zz_4439_ = int_reg_array_2_3_real;
      end
      6'b000100 : begin
        _zz_4438_ = int_reg_array_2_4_imag;
        _zz_4439_ = int_reg_array_2_4_real;
      end
      6'b000101 : begin
        _zz_4438_ = int_reg_array_2_5_imag;
        _zz_4439_ = int_reg_array_2_5_real;
      end
      6'b000110 : begin
        _zz_4438_ = int_reg_array_2_6_imag;
        _zz_4439_ = int_reg_array_2_6_real;
      end
      6'b000111 : begin
        _zz_4438_ = int_reg_array_2_7_imag;
        _zz_4439_ = int_reg_array_2_7_real;
      end
      6'b001000 : begin
        _zz_4438_ = int_reg_array_2_8_imag;
        _zz_4439_ = int_reg_array_2_8_real;
      end
      6'b001001 : begin
        _zz_4438_ = int_reg_array_2_9_imag;
        _zz_4439_ = int_reg_array_2_9_real;
      end
      6'b001010 : begin
        _zz_4438_ = int_reg_array_2_10_imag;
        _zz_4439_ = int_reg_array_2_10_real;
      end
      6'b001011 : begin
        _zz_4438_ = int_reg_array_2_11_imag;
        _zz_4439_ = int_reg_array_2_11_real;
      end
      6'b001100 : begin
        _zz_4438_ = int_reg_array_2_12_imag;
        _zz_4439_ = int_reg_array_2_12_real;
      end
      6'b001101 : begin
        _zz_4438_ = int_reg_array_2_13_imag;
        _zz_4439_ = int_reg_array_2_13_real;
      end
      6'b001110 : begin
        _zz_4438_ = int_reg_array_2_14_imag;
        _zz_4439_ = int_reg_array_2_14_real;
      end
      6'b001111 : begin
        _zz_4438_ = int_reg_array_2_15_imag;
        _zz_4439_ = int_reg_array_2_15_real;
      end
      6'b010000 : begin
        _zz_4438_ = int_reg_array_2_16_imag;
        _zz_4439_ = int_reg_array_2_16_real;
      end
      6'b010001 : begin
        _zz_4438_ = int_reg_array_2_17_imag;
        _zz_4439_ = int_reg_array_2_17_real;
      end
      6'b010010 : begin
        _zz_4438_ = int_reg_array_2_18_imag;
        _zz_4439_ = int_reg_array_2_18_real;
      end
      6'b010011 : begin
        _zz_4438_ = int_reg_array_2_19_imag;
        _zz_4439_ = int_reg_array_2_19_real;
      end
      6'b010100 : begin
        _zz_4438_ = int_reg_array_2_20_imag;
        _zz_4439_ = int_reg_array_2_20_real;
      end
      6'b010101 : begin
        _zz_4438_ = int_reg_array_2_21_imag;
        _zz_4439_ = int_reg_array_2_21_real;
      end
      6'b010110 : begin
        _zz_4438_ = int_reg_array_2_22_imag;
        _zz_4439_ = int_reg_array_2_22_real;
      end
      6'b010111 : begin
        _zz_4438_ = int_reg_array_2_23_imag;
        _zz_4439_ = int_reg_array_2_23_real;
      end
      6'b011000 : begin
        _zz_4438_ = int_reg_array_2_24_imag;
        _zz_4439_ = int_reg_array_2_24_real;
      end
      6'b011001 : begin
        _zz_4438_ = int_reg_array_2_25_imag;
        _zz_4439_ = int_reg_array_2_25_real;
      end
      6'b011010 : begin
        _zz_4438_ = int_reg_array_2_26_imag;
        _zz_4439_ = int_reg_array_2_26_real;
      end
      6'b011011 : begin
        _zz_4438_ = int_reg_array_2_27_imag;
        _zz_4439_ = int_reg_array_2_27_real;
      end
      6'b011100 : begin
        _zz_4438_ = int_reg_array_2_28_imag;
        _zz_4439_ = int_reg_array_2_28_real;
      end
      6'b011101 : begin
        _zz_4438_ = int_reg_array_2_29_imag;
        _zz_4439_ = int_reg_array_2_29_real;
      end
      6'b011110 : begin
        _zz_4438_ = int_reg_array_2_30_imag;
        _zz_4439_ = int_reg_array_2_30_real;
      end
      6'b011111 : begin
        _zz_4438_ = int_reg_array_2_31_imag;
        _zz_4439_ = int_reg_array_2_31_real;
      end
      6'b100000 : begin
        _zz_4438_ = int_reg_array_2_32_imag;
        _zz_4439_ = int_reg_array_2_32_real;
      end
      6'b100001 : begin
        _zz_4438_ = int_reg_array_2_33_imag;
        _zz_4439_ = int_reg_array_2_33_real;
      end
      6'b100010 : begin
        _zz_4438_ = int_reg_array_2_34_imag;
        _zz_4439_ = int_reg_array_2_34_real;
      end
      6'b100011 : begin
        _zz_4438_ = int_reg_array_2_35_imag;
        _zz_4439_ = int_reg_array_2_35_real;
      end
      6'b100100 : begin
        _zz_4438_ = int_reg_array_2_36_imag;
        _zz_4439_ = int_reg_array_2_36_real;
      end
      6'b100101 : begin
        _zz_4438_ = int_reg_array_2_37_imag;
        _zz_4439_ = int_reg_array_2_37_real;
      end
      6'b100110 : begin
        _zz_4438_ = int_reg_array_2_38_imag;
        _zz_4439_ = int_reg_array_2_38_real;
      end
      6'b100111 : begin
        _zz_4438_ = int_reg_array_2_39_imag;
        _zz_4439_ = int_reg_array_2_39_real;
      end
      6'b101000 : begin
        _zz_4438_ = int_reg_array_2_40_imag;
        _zz_4439_ = int_reg_array_2_40_real;
      end
      6'b101001 : begin
        _zz_4438_ = int_reg_array_2_41_imag;
        _zz_4439_ = int_reg_array_2_41_real;
      end
      6'b101010 : begin
        _zz_4438_ = int_reg_array_2_42_imag;
        _zz_4439_ = int_reg_array_2_42_real;
      end
      6'b101011 : begin
        _zz_4438_ = int_reg_array_2_43_imag;
        _zz_4439_ = int_reg_array_2_43_real;
      end
      6'b101100 : begin
        _zz_4438_ = int_reg_array_2_44_imag;
        _zz_4439_ = int_reg_array_2_44_real;
      end
      6'b101101 : begin
        _zz_4438_ = int_reg_array_2_45_imag;
        _zz_4439_ = int_reg_array_2_45_real;
      end
      6'b101110 : begin
        _zz_4438_ = int_reg_array_2_46_imag;
        _zz_4439_ = int_reg_array_2_46_real;
      end
      6'b101111 : begin
        _zz_4438_ = int_reg_array_2_47_imag;
        _zz_4439_ = int_reg_array_2_47_real;
      end
      6'b110000 : begin
        _zz_4438_ = int_reg_array_2_48_imag;
        _zz_4439_ = int_reg_array_2_48_real;
      end
      6'b110001 : begin
        _zz_4438_ = int_reg_array_2_49_imag;
        _zz_4439_ = int_reg_array_2_49_real;
      end
      6'b110010 : begin
        _zz_4438_ = int_reg_array_2_50_imag;
        _zz_4439_ = int_reg_array_2_50_real;
      end
      6'b110011 : begin
        _zz_4438_ = int_reg_array_2_51_imag;
        _zz_4439_ = int_reg_array_2_51_real;
      end
      6'b110100 : begin
        _zz_4438_ = int_reg_array_2_52_imag;
        _zz_4439_ = int_reg_array_2_52_real;
      end
      6'b110101 : begin
        _zz_4438_ = int_reg_array_2_53_imag;
        _zz_4439_ = int_reg_array_2_53_real;
      end
      6'b110110 : begin
        _zz_4438_ = int_reg_array_2_54_imag;
        _zz_4439_ = int_reg_array_2_54_real;
      end
      6'b110111 : begin
        _zz_4438_ = int_reg_array_2_55_imag;
        _zz_4439_ = int_reg_array_2_55_real;
      end
      6'b111000 : begin
        _zz_4438_ = int_reg_array_2_56_imag;
        _zz_4439_ = int_reg_array_2_56_real;
      end
      6'b111001 : begin
        _zz_4438_ = int_reg_array_2_57_imag;
        _zz_4439_ = int_reg_array_2_57_real;
      end
      6'b111010 : begin
        _zz_4438_ = int_reg_array_2_58_imag;
        _zz_4439_ = int_reg_array_2_58_real;
      end
      6'b111011 : begin
        _zz_4438_ = int_reg_array_2_59_imag;
        _zz_4439_ = int_reg_array_2_59_real;
      end
      6'b111100 : begin
        _zz_4438_ = int_reg_array_2_60_imag;
        _zz_4439_ = int_reg_array_2_60_real;
      end
      6'b111101 : begin
        _zz_4438_ = int_reg_array_2_61_imag;
        _zz_4439_ = int_reg_array_2_61_real;
      end
      6'b111110 : begin
        _zz_4438_ = int_reg_array_2_62_imag;
        _zz_4439_ = int_reg_array_2_62_real;
      end
      default : begin
        _zz_4438_ = int_reg_array_2_63_imag;
        _zz_4439_ = int_reg_array_2_63_real;
      end
    endcase
  end

  always @(*) begin
    case(_zz_224_)
      6'b000000 : begin
        _zz_4440_ = int_reg_array_3_0_imag;
        _zz_4441_ = int_reg_array_3_0_real;
      end
      6'b000001 : begin
        _zz_4440_ = int_reg_array_3_1_imag;
        _zz_4441_ = int_reg_array_3_1_real;
      end
      6'b000010 : begin
        _zz_4440_ = int_reg_array_3_2_imag;
        _zz_4441_ = int_reg_array_3_2_real;
      end
      6'b000011 : begin
        _zz_4440_ = int_reg_array_3_3_imag;
        _zz_4441_ = int_reg_array_3_3_real;
      end
      6'b000100 : begin
        _zz_4440_ = int_reg_array_3_4_imag;
        _zz_4441_ = int_reg_array_3_4_real;
      end
      6'b000101 : begin
        _zz_4440_ = int_reg_array_3_5_imag;
        _zz_4441_ = int_reg_array_3_5_real;
      end
      6'b000110 : begin
        _zz_4440_ = int_reg_array_3_6_imag;
        _zz_4441_ = int_reg_array_3_6_real;
      end
      6'b000111 : begin
        _zz_4440_ = int_reg_array_3_7_imag;
        _zz_4441_ = int_reg_array_3_7_real;
      end
      6'b001000 : begin
        _zz_4440_ = int_reg_array_3_8_imag;
        _zz_4441_ = int_reg_array_3_8_real;
      end
      6'b001001 : begin
        _zz_4440_ = int_reg_array_3_9_imag;
        _zz_4441_ = int_reg_array_3_9_real;
      end
      6'b001010 : begin
        _zz_4440_ = int_reg_array_3_10_imag;
        _zz_4441_ = int_reg_array_3_10_real;
      end
      6'b001011 : begin
        _zz_4440_ = int_reg_array_3_11_imag;
        _zz_4441_ = int_reg_array_3_11_real;
      end
      6'b001100 : begin
        _zz_4440_ = int_reg_array_3_12_imag;
        _zz_4441_ = int_reg_array_3_12_real;
      end
      6'b001101 : begin
        _zz_4440_ = int_reg_array_3_13_imag;
        _zz_4441_ = int_reg_array_3_13_real;
      end
      6'b001110 : begin
        _zz_4440_ = int_reg_array_3_14_imag;
        _zz_4441_ = int_reg_array_3_14_real;
      end
      6'b001111 : begin
        _zz_4440_ = int_reg_array_3_15_imag;
        _zz_4441_ = int_reg_array_3_15_real;
      end
      6'b010000 : begin
        _zz_4440_ = int_reg_array_3_16_imag;
        _zz_4441_ = int_reg_array_3_16_real;
      end
      6'b010001 : begin
        _zz_4440_ = int_reg_array_3_17_imag;
        _zz_4441_ = int_reg_array_3_17_real;
      end
      6'b010010 : begin
        _zz_4440_ = int_reg_array_3_18_imag;
        _zz_4441_ = int_reg_array_3_18_real;
      end
      6'b010011 : begin
        _zz_4440_ = int_reg_array_3_19_imag;
        _zz_4441_ = int_reg_array_3_19_real;
      end
      6'b010100 : begin
        _zz_4440_ = int_reg_array_3_20_imag;
        _zz_4441_ = int_reg_array_3_20_real;
      end
      6'b010101 : begin
        _zz_4440_ = int_reg_array_3_21_imag;
        _zz_4441_ = int_reg_array_3_21_real;
      end
      6'b010110 : begin
        _zz_4440_ = int_reg_array_3_22_imag;
        _zz_4441_ = int_reg_array_3_22_real;
      end
      6'b010111 : begin
        _zz_4440_ = int_reg_array_3_23_imag;
        _zz_4441_ = int_reg_array_3_23_real;
      end
      6'b011000 : begin
        _zz_4440_ = int_reg_array_3_24_imag;
        _zz_4441_ = int_reg_array_3_24_real;
      end
      6'b011001 : begin
        _zz_4440_ = int_reg_array_3_25_imag;
        _zz_4441_ = int_reg_array_3_25_real;
      end
      6'b011010 : begin
        _zz_4440_ = int_reg_array_3_26_imag;
        _zz_4441_ = int_reg_array_3_26_real;
      end
      6'b011011 : begin
        _zz_4440_ = int_reg_array_3_27_imag;
        _zz_4441_ = int_reg_array_3_27_real;
      end
      6'b011100 : begin
        _zz_4440_ = int_reg_array_3_28_imag;
        _zz_4441_ = int_reg_array_3_28_real;
      end
      6'b011101 : begin
        _zz_4440_ = int_reg_array_3_29_imag;
        _zz_4441_ = int_reg_array_3_29_real;
      end
      6'b011110 : begin
        _zz_4440_ = int_reg_array_3_30_imag;
        _zz_4441_ = int_reg_array_3_30_real;
      end
      6'b011111 : begin
        _zz_4440_ = int_reg_array_3_31_imag;
        _zz_4441_ = int_reg_array_3_31_real;
      end
      6'b100000 : begin
        _zz_4440_ = int_reg_array_3_32_imag;
        _zz_4441_ = int_reg_array_3_32_real;
      end
      6'b100001 : begin
        _zz_4440_ = int_reg_array_3_33_imag;
        _zz_4441_ = int_reg_array_3_33_real;
      end
      6'b100010 : begin
        _zz_4440_ = int_reg_array_3_34_imag;
        _zz_4441_ = int_reg_array_3_34_real;
      end
      6'b100011 : begin
        _zz_4440_ = int_reg_array_3_35_imag;
        _zz_4441_ = int_reg_array_3_35_real;
      end
      6'b100100 : begin
        _zz_4440_ = int_reg_array_3_36_imag;
        _zz_4441_ = int_reg_array_3_36_real;
      end
      6'b100101 : begin
        _zz_4440_ = int_reg_array_3_37_imag;
        _zz_4441_ = int_reg_array_3_37_real;
      end
      6'b100110 : begin
        _zz_4440_ = int_reg_array_3_38_imag;
        _zz_4441_ = int_reg_array_3_38_real;
      end
      6'b100111 : begin
        _zz_4440_ = int_reg_array_3_39_imag;
        _zz_4441_ = int_reg_array_3_39_real;
      end
      6'b101000 : begin
        _zz_4440_ = int_reg_array_3_40_imag;
        _zz_4441_ = int_reg_array_3_40_real;
      end
      6'b101001 : begin
        _zz_4440_ = int_reg_array_3_41_imag;
        _zz_4441_ = int_reg_array_3_41_real;
      end
      6'b101010 : begin
        _zz_4440_ = int_reg_array_3_42_imag;
        _zz_4441_ = int_reg_array_3_42_real;
      end
      6'b101011 : begin
        _zz_4440_ = int_reg_array_3_43_imag;
        _zz_4441_ = int_reg_array_3_43_real;
      end
      6'b101100 : begin
        _zz_4440_ = int_reg_array_3_44_imag;
        _zz_4441_ = int_reg_array_3_44_real;
      end
      6'b101101 : begin
        _zz_4440_ = int_reg_array_3_45_imag;
        _zz_4441_ = int_reg_array_3_45_real;
      end
      6'b101110 : begin
        _zz_4440_ = int_reg_array_3_46_imag;
        _zz_4441_ = int_reg_array_3_46_real;
      end
      6'b101111 : begin
        _zz_4440_ = int_reg_array_3_47_imag;
        _zz_4441_ = int_reg_array_3_47_real;
      end
      6'b110000 : begin
        _zz_4440_ = int_reg_array_3_48_imag;
        _zz_4441_ = int_reg_array_3_48_real;
      end
      6'b110001 : begin
        _zz_4440_ = int_reg_array_3_49_imag;
        _zz_4441_ = int_reg_array_3_49_real;
      end
      6'b110010 : begin
        _zz_4440_ = int_reg_array_3_50_imag;
        _zz_4441_ = int_reg_array_3_50_real;
      end
      6'b110011 : begin
        _zz_4440_ = int_reg_array_3_51_imag;
        _zz_4441_ = int_reg_array_3_51_real;
      end
      6'b110100 : begin
        _zz_4440_ = int_reg_array_3_52_imag;
        _zz_4441_ = int_reg_array_3_52_real;
      end
      6'b110101 : begin
        _zz_4440_ = int_reg_array_3_53_imag;
        _zz_4441_ = int_reg_array_3_53_real;
      end
      6'b110110 : begin
        _zz_4440_ = int_reg_array_3_54_imag;
        _zz_4441_ = int_reg_array_3_54_real;
      end
      6'b110111 : begin
        _zz_4440_ = int_reg_array_3_55_imag;
        _zz_4441_ = int_reg_array_3_55_real;
      end
      6'b111000 : begin
        _zz_4440_ = int_reg_array_3_56_imag;
        _zz_4441_ = int_reg_array_3_56_real;
      end
      6'b111001 : begin
        _zz_4440_ = int_reg_array_3_57_imag;
        _zz_4441_ = int_reg_array_3_57_real;
      end
      6'b111010 : begin
        _zz_4440_ = int_reg_array_3_58_imag;
        _zz_4441_ = int_reg_array_3_58_real;
      end
      6'b111011 : begin
        _zz_4440_ = int_reg_array_3_59_imag;
        _zz_4441_ = int_reg_array_3_59_real;
      end
      6'b111100 : begin
        _zz_4440_ = int_reg_array_3_60_imag;
        _zz_4441_ = int_reg_array_3_60_real;
      end
      6'b111101 : begin
        _zz_4440_ = int_reg_array_3_61_imag;
        _zz_4441_ = int_reg_array_3_61_real;
      end
      6'b111110 : begin
        _zz_4440_ = int_reg_array_3_62_imag;
        _zz_4441_ = int_reg_array_3_62_real;
      end
      default : begin
        _zz_4440_ = int_reg_array_3_63_imag;
        _zz_4441_ = int_reg_array_3_63_real;
      end
    endcase
  end

  always @(*) begin
    case(_zz_293_)
      6'b000000 : begin
        _zz_4442_ = int_reg_array_4_0_imag;
        _zz_4443_ = int_reg_array_4_0_real;
      end
      6'b000001 : begin
        _zz_4442_ = int_reg_array_4_1_imag;
        _zz_4443_ = int_reg_array_4_1_real;
      end
      6'b000010 : begin
        _zz_4442_ = int_reg_array_4_2_imag;
        _zz_4443_ = int_reg_array_4_2_real;
      end
      6'b000011 : begin
        _zz_4442_ = int_reg_array_4_3_imag;
        _zz_4443_ = int_reg_array_4_3_real;
      end
      6'b000100 : begin
        _zz_4442_ = int_reg_array_4_4_imag;
        _zz_4443_ = int_reg_array_4_4_real;
      end
      6'b000101 : begin
        _zz_4442_ = int_reg_array_4_5_imag;
        _zz_4443_ = int_reg_array_4_5_real;
      end
      6'b000110 : begin
        _zz_4442_ = int_reg_array_4_6_imag;
        _zz_4443_ = int_reg_array_4_6_real;
      end
      6'b000111 : begin
        _zz_4442_ = int_reg_array_4_7_imag;
        _zz_4443_ = int_reg_array_4_7_real;
      end
      6'b001000 : begin
        _zz_4442_ = int_reg_array_4_8_imag;
        _zz_4443_ = int_reg_array_4_8_real;
      end
      6'b001001 : begin
        _zz_4442_ = int_reg_array_4_9_imag;
        _zz_4443_ = int_reg_array_4_9_real;
      end
      6'b001010 : begin
        _zz_4442_ = int_reg_array_4_10_imag;
        _zz_4443_ = int_reg_array_4_10_real;
      end
      6'b001011 : begin
        _zz_4442_ = int_reg_array_4_11_imag;
        _zz_4443_ = int_reg_array_4_11_real;
      end
      6'b001100 : begin
        _zz_4442_ = int_reg_array_4_12_imag;
        _zz_4443_ = int_reg_array_4_12_real;
      end
      6'b001101 : begin
        _zz_4442_ = int_reg_array_4_13_imag;
        _zz_4443_ = int_reg_array_4_13_real;
      end
      6'b001110 : begin
        _zz_4442_ = int_reg_array_4_14_imag;
        _zz_4443_ = int_reg_array_4_14_real;
      end
      6'b001111 : begin
        _zz_4442_ = int_reg_array_4_15_imag;
        _zz_4443_ = int_reg_array_4_15_real;
      end
      6'b010000 : begin
        _zz_4442_ = int_reg_array_4_16_imag;
        _zz_4443_ = int_reg_array_4_16_real;
      end
      6'b010001 : begin
        _zz_4442_ = int_reg_array_4_17_imag;
        _zz_4443_ = int_reg_array_4_17_real;
      end
      6'b010010 : begin
        _zz_4442_ = int_reg_array_4_18_imag;
        _zz_4443_ = int_reg_array_4_18_real;
      end
      6'b010011 : begin
        _zz_4442_ = int_reg_array_4_19_imag;
        _zz_4443_ = int_reg_array_4_19_real;
      end
      6'b010100 : begin
        _zz_4442_ = int_reg_array_4_20_imag;
        _zz_4443_ = int_reg_array_4_20_real;
      end
      6'b010101 : begin
        _zz_4442_ = int_reg_array_4_21_imag;
        _zz_4443_ = int_reg_array_4_21_real;
      end
      6'b010110 : begin
        _zz_4442_ = int_reg_array_4_22_imag;
        _zz_4443_ = int_reg_array_4_22_real;
      end
      6'b010111 : begin
        _zz_4442_ = int_reg_array_4_23_imag;
        _zz_4443_ = int_reg_array_4_23_real;
      end
      6'b011000 : begin
        _zz_4442_ = int_reg_array_4_24_imag;
        _zz_4443_ = int_reg_array_4_24_real;
      end
      6'b011001 : begin
        _zz_4442_ = int_reg_array_4_25_imag;
        _zz_4443_ = int_reg_array_4_25_real;
      end
      6'b011010 : begin
        _zz_4442_ = int_reg_array_4_26_imag;
        _zz_4443_ = int_reg_array_4_26_real;
      end
      6'b011011 : begin
        _zz_4442_ = int_reg_array_4_27_imag;
        _zz_4443_ = int_reg_array_4_27_real;
      end
      6'b011100 : begin
        _zz_4442_ = int_reg_array_4_28_imag;
        _zz_4443_ = int_reg_array_4_28_real;
      end
      6'b011101 : begin
        _zz_4442_ = int_reg_array_4_29_imag;
        _zz_4443_ = int_reg_array_4_29_real;
      end
      6'b011110 : begin
        _zz_4442_ = int_reg_array_4_30_imag;
        _zz_4443_ = int_reg_array_4_30_real;
      end
      6'b011111 : begin
        _zz_4442_ = int_reg_array_4_31_imag;
        _zz_4443_ = int_reg_array_4_31_real;
      end
      6'b100000 : begin
        _zz_4442_ = int_reg_array_4_32_imag;
        _zz_4443_ = int_reg_array_4_32_real;
      end
      6'b100001 : begin
        _zz_4442_ = int_reg_array_4_33_imag;
        _zz_4443_ = int_reg_array_4_33_real;
      end
      6'b100010 : begin
        _zz_4442_ = int_reg_array_4_34_imag;
        _zz_4443_ = int_reg_array_4_34_real;
      end
      6'b100011 : begin
        _zz_4442_ = int_reg_array_4_35_imag;
        _zz_4443_ = int_reg_array_4_35_real;
      end
      6'b100100 : begin
        _zz_4442_ = int_reg_array_4_36_imag;
        _zz_4443_ = int_reg_array_4_36_real;
      end
      6'b100101 : begin
        _zz_4442_ = int_reg_array_4_37_imag;
        _zz_4443_ = int_reg_array_4_37_real;
      end
      6'b100110 : begin
        _zz_4442_ = int_reg_array_4_38_imag;
        _zz_4443_ = int_reg_array_4_38_real;
      end
      6'b100111 : begin
        _zz_4442_ = int_reg_array_4_39_imag;
        _zz_4443_ = int_reg_array_4_39_real;
      end
      6'b101000 : begin
        _zz_4442_ = int_reg_array_4_40_imag;
        _zz_4443_ = int_reg_array_4_40_real;
      end
      6'b101001 : begin
        _zz_4442_ = int_reg_array_4_41_imag;
        _zz_4443_ = int_reg_array_4_41_real;
      end
      6'b101010 : begin
        _zz_4442_ = int_reg_array_4_42_imag;
        _zz_4443_ = int_reg_array_4_42_real;
      end
      6'b101011 : begin
        _zz_4442_ = int_reg_array_4_43_imag;
        _zz_4443_ = int_reg_array_4_43_real;
      end
      6'b101100 : begin
        _zz_4442_ = int_reg_array_4_44_imag;
        _zz_4443_ = int_reg_array_4_44_real;
      end
      6'b101101 : begin
        _zz_4442_ = int_reg_array_4_45_imag;
        _zz_4443_ = int_reg_array_4_45_real;
      end
      6'b101110 : begin
        _zz_4442_ = int_reg_array_4_46_imag;
        _zz_4443_ = int_reg_array_4_46_real;
      end
      6'b101111 : begin
        _zz_4442_ = int_reg_array_4_47_imag;
        _zz_4443_ = int_reg_array_4_47_real;
      end
      6'b110000 : begin
        _zz_4442_ = int_reg_array_4_48_imag;
        _zz_4443_ = int_reg_array_4_48_real;
      end
      6'b110001 : begin
        _zz_4442_ = int_reg_array_4_49_imag;
        _zz_4443_ = int_reg_array_4_49_real;
      end
      6'b110010 : begin
        _zz_4442_ = int_reg_array_4_50_imag;
        _zz_4443_ = int_reg_array_4_50_real;
      end
      6'b110011 : begin
        _zz_4442_ = int_reg_array_4_51_imag;
        _zz_4443_ = int_reg_array_4_51_real;
      end
      6'b110100 : begin
        _zz_4442_ = int_reg_array_4_52_imag;
        _zz_4443_ = int_reg_array_4_52_real;
      end
      6'b110101 : begin
        _zz_4442_ = int_reg_array_4_53_imag;
        _zz_4443_ = int_reg_array_4_53_real;
      end
      6'b110110 : begin
        _zz_4442_ = int_reg_array_4_54_imag;
        _zz_4443_ = int_reg_array_4_54_real;
      end
      6'b110111 : begin
        _zz_4442_ = int_reg_array_4_55_imag;
        _zz_4443_ = int_reg_array_4_55_real;
      end
      6'b111000 : begin
        _zz_4442_ = int_reg_array_4_56_imag;
        _zz_4443_ = int_reg_array_4_56_real;
      end
      6'b111001 : begin
        _zz_4442_ = int_reg_array_4_57_imag;
        _zz_4443_ = int_reg_array_4_57_real;
      end
      6'b111010 : begin
        _zz_4442_ = int_reg_array_4_58_imag;
        _zz_4443_ = int_reg_array_4_58_real;
      end
      6'b111011 : begin
        _zz_4442_ = int_reg_array_4_59_imag;
        _zz_4443_ = int_reg_array_4_59_real;
      end
      6'b111100 : begin
        _zz_4442_ = int_reg_array_4_60_imag;
        _zz_4443_ = int_reg_array_4_60_real;
      end
      6'b111101 : begin
        _zz_4442_ = int_reg_array_4_61_imag;
        _zz_4443_ = int_reg_array_4_61_real;
      end
      6'b111110 : begin
        _zz_4442_ = int_reg_array_4_62_imag;
        _zz_4443_ = int_reg_array_4_62_real;
      end
      default : begin
        _zz_4442_ = int_reg_array_4_63_imag;
        _zz_4443_ = int_reg_array_4_63_real;
      end
    endcase
  end

  always @(*) begin
    case(_zz_362_)
      6'b000000 : begin
        _zz_4444_ = int_reg_array_5_0_imag;
        _zz_4445_ = int_reg_array_5_0_real;
      end
      6'b000001 : begin
        _zz_4444_ = int_reg_array_5_1_imag;
        _zz_4445_ = int_reg_array_5_1_real;
      end
      6'b000010 : begin
        _zz_4444_ = int_reg_array_5_2_imag;
        _zz_4445_ = int_reg_array_5_2_real;
      end
      6'b000011 : begin
        _zz_4444_ = int_reg_array_5_3_imag;
        _zz_4445_ = int_reg_array_5_3_real;
      end
      6'b000100 : begin
        _zz_4444_ = int_reg_array_5_4_imag;
        _zz_4445_ = int_reg_array_5_4_real;
      end
      6'b000101 : begin
        _zz_4444_ = int_reg_array_5_5_imag;
        _zz_4445_ = int_reg_array_5_5_real;
      end
      6'b000110 : begin
        _zz_4444_ = int_reg_array_5_6_imag;
        _zz_4445_ = int_reg_array_5_6_real;
      end
      6'b000111 : begin
        _zz_4444_ = int_reg_array_5_7_imag;
        _zz_4445_ = int_reg_array_5_7_real;
      end
      6'b001000 : begin
        _zz_4444_ = int_reg_array_5_8_imag;
        _zz_4445_ = int_reg_array_5_8_real;
      end
      6'b001001 : begin
        _zz_4444_ = int_reg_array_5_9_imag;
        _zz_4445_ = int_reg_array_5_9_real;
      end
      6'b001010 : begin
        _zz_4444_ = int_reg_array_5_10_imag;
        _zz_4445_ = int_reg_array_5_10_real;
      end
      6'b001011 : begin
        _zz_4444_ = int_reg_array_5_11_imag;
        _zz_4445_ = int_reg_array_5_11_real;
      end
      6'b001100 : begin
        _zz_4444_ = int_reg_array_5_12_imag;
        _zz_4445_ = int_reg_array_5_12_real;
      end
      6'b001101 : begin
        _zz_4444_ = int_reg_array_5_13_imag;
        _zz_4445_ = int_reg_array_5_13_real;
      end
      6'b001110 : begin
        _zz_4444_ = int_reg_array_5_14_imag;
        _zz_4445_ = int_reg_array_5_14_real;
      end
      6'b001111 : begin
        _zz_4444_ = int_reg_array_5_15_imag;
        _zz_4445_ = int_reg_array_5_15_real;
      end
      6'b010000 : begin
        _zz_4444_ = int_reg_array_5_16_imag;
        _zz_4445_ = int_reg_array_5_16_real;
      end
      6'b010001 : begin
        _zz_4444_ = int_reg_array_5_17_imag;
        _zz_4445_ = int_reg_array_5_17_real;
      end
      6'b010010 : begin
        _zz_4444_ = int_reg_array_5_18_imag;
        _zz_4445_ = int_reg_array_5_18_real;
      end
      6'b010011 : begin
        _zz_4444_ = int_reg_array_5_19_imag;
        _zz_4445_ = int_reg_array_5_19_real;
      end
      6'b010100 : begin
        _zz_4444_ = int_reg_array_5_20_imag;
        _zz_4445_ = int_reg_array_5_20_real;
      end
      6'b010101 : begin
        _zz_4444_ = int_reg_array_5_21_imag;
        _zz_4445_ = int_reg_array_5_21_real;
      end
      6'b010110 : begin
        _zz_4444_ = int_reg_array_5_22_imag;
        _zz_4445_ = int_reg_array_5_22_real;
      end
      6'b010111 : begin
        _zz_4444_ = int_reg_array_5_23_imag;
        _zz_4445_ = int_reg_array_5_23_real;
      end
      6'b011000 : begin
        _zz_4444_ = int_reg_array_5_24_imag;
        _zz_4445_ = int_reg_array_5_24_real;
      end
      6'b011001 : begin
        _zz_4444_ = int_reg_array_5_25_imag;
        _zz_4445_ = int_reg_array_5_25_real;
      end
      6'b011010 : begin
        _zz_4444_ = int_reg_array_5_26_imag;
        _zz_4445_ = int_reg_array_5_26_real;
      end
      6'b011011 : begin
        _zz_4444_ = int_reg_array_5_27_imag;
        _zz_4445_ = int_reg_array_5_27_real;
      end
      6'b011100 : begin
        _zz_4444_ = int_reg_array_5_28_imag;
        _zz_4445_ = int_reg_array_5_28_real;
      end
      6'b011101 : begin
        _zz_4444_ = int_reg_array_5_29_imag;
        _zz_4445_ = int_reg_array_5_29_real;
      end
      6'b011110 : begin
        _zz_4444_ = int_reg_array_5_30_imag;
        _zz_4445_ = int_reg_array_5_30_real;
      end
      6'b011111 : begin
        _zz_4444_ = int_reg_array_5_31_imag;
        _zz_4445_ = int_reg_array_5_31_real;
      end
      6'b100000 : begin
        _zz_4444_ = int_reg_array_5_32_imag;
        _zz_4445_ = int_reg_array_5_32_real;
      end
      6'b100001 : begin
        _zz_4444_ = int_reg_array_5_33_imag;
        _zz_4445_ = int_reg_array_5_33_real;
      end
      6'b100010 : begin
        _zz_4444_ = int_reg_array_5_34_imag;
        _zz_4445_ = int_reg_array_5_34_real;
      end
      6'b100011 : begin
        _zz_4444_ = int_reg_array_5_35_imag;
        _zz_4445_ = int_reg_array_5_35_real;
      end
      6'b100100 : begin
        _zz_4444_ = int_reg_array_5_36_imag;
        _zz_4445_ = int_reg_array_5_36_real;
      end
      6'b100101 : begin
        _zz_4444_ = int_reg_array_5_37_imag;
        _zz_4445_ = int_reg_array_5_37_real;
      end
      6'b100110 : begin
        _zz_4444_ = int_reg_array_5_38_imag;
        _zz_4445_ = int_reg_array_5_38_real;
      end
      6'b100111 : begin
        _zz_4444_ = int_reg_array_5_39_imag;
        _zz_4445_ = int_reg_array_5_39_real;
      end
      6'b101000 : begin
        _zz_4444_ = int_reg_array_5_40_imag;
        _zz_4445_ = int_reg_array_5_40_real;
      end
      6'b101001 : begin
        _zz_4444_ = int_reg_array_5_41_imag;
        _zz_4445_ = int_reg_array_5_41_real;
      end
      6'b101010 : begin
        _zz_4444_ = int_reg_array_5_42_imag;
        _zz_4445_ = int_reg_array_5_42_real;
      end
      6'b101011 : begin
        _zz_4444_ = int_reg_array_5_43_imag;
        _zz_4445_ = int_reg_array_5_43_real;
      end
      6'b101100 : begin
        _zz_4444_ = int_reg_array_5_44_imag;
        _zz_4445_ = int_reg_array_5_44_real;
      end
      6'b101101 : begin
        _zz_4444_ = int_reg_array_5_45_imag;
        _zz_4445_ = int_reg_array_5_45_real;
      end
      6'b101110 : begin
        _zz_4444_ = int_reg_array_5_46_imag;
        _zz_4445_ = int_reg_array_5_46_real;
      end
      6'b101111 : begin
        _zz_4444_ = int_reg_array_5_47_imag;
        _zz_4445_ = int_reg_array_5_47_real;
      end
      6'b110000 : begin
        _zz_4444_ = int_reg_array_5_48_imag;
        _zz_4445_ = int_reg_array_5_48_real;
      end
      6'b110001 : begin
        _zz_4444_ = int_reg_array_5_49_imag;
        _zz_4445_ = int_reg_array_5_49_real;
      end
      6'b110010 : begin
        _zz_4444_ = int_reg_array_5_50_imag;
        _zz_4445_ = int_reg_array_5_50_real;
      end
      6'b110011 : begin
        _zz_4444_ = int_reg_array_5_51_imag;
        _zz_4445_ = int_reg_array_5_51_real;
      end
      6'b110100 : begin
        _zz_4444_ = int_reg_array_5_52_imag;
        _zz_4445_ = int_reg_array_5_52_real;
      end
      6'b110101 : begin
        _zz_4444_ = int_reg_array_5_53_imag;
        _zz_4445_ = int_reg_array_5_53_real;
      end
      6'b110110 : begin
        _zz_4444_ = int_reg_array_5_54_imag;
        _zz_4445_ = int_reg_array_5_54_real;
      end
      6'b110111 : begin
        _zz_4444_ = int_reg_array_5_55_imag;
        _zz_4445_ = int_reg_array_5_55_real;
      end
      6'b111000 : begin
        _zz_4444_ = int_reg_array_5_56_imag;
        _zz_4445_ = int_reg_array_5_56_real;
      end
      6'b111001 : begin
        _zz_4444_ = int_reg_array_5_57_imag;
        _zz_4445_ = int_reg_array_5_57_real;
      end
      6'b111010 : begin
        _zz_4444_ = int_reg_array_5_58_imag;
        _zz_4445_ = int_reg_array_5_58_real;
      end
      6'b111011 : begin
        _zz_4444_ = int_reg_array_5_59_imag;
        _zz_4445_ = int_reg_array_5_59_real;
      end
      6'b111100 : begin
        _zz_4444_ = int_reg_array_5_60_imag;
        _zz_4445_ = int_reg_array_5_60_real;
      end
      6'b111101 : begin
        _zz_4444_ = int_reg_array_5_61_imag;
        _zz_4445_ = int_reg_array_5_61_real;
      end
      6'b111110 : begin
        _zz_4444_ = int_reg_array_5_62_imag;
        _zz_4445_ = int_reg_array_5_62_real;
      end
      default : begin
        _zz_4444_ = int_reg_array_5_63_imag;
        _zz_4445_ = int_reg_array_5_63_real;
      end
    endcase
  end

  always @(*) begin
    case(_zz_431_)
      6'b000000 : begin
        _zz_4446_ = int_reg_array_6_0_imag;
        _zz_4447_ = int_reg_array_6_0_real;
      end
      6'b000001 : begin
        _zz_4446_ = int_reg_array_6_1_imag;
        _zz_4447_ = int_reg_array_6_1_real;
      end
      6'b000010 : begin
        _zz_4446_ = int_reg_array_6_2_imag;
        _zz_4447_ = int_reg_array_6_2_real;
      end
      6'b000011 : begin
        _zz_4446_ = int_reg_array_6_3_imag;
        _zz_4447_ = int_reg_array_6_3_real;
      end
      6'b000100 : begin
        _zz_4446_ = int_reg_array_6_4_imag;
        _zz_4447_ = int_reg_array_6_4_real;
      end
      6'b000101 : begin
        _zz_4446_ = int_reg_array_6_5_imag;
        _zz_4447_ = int_reg_array_6_5_real;
      end
      6'b000110 : begin
        _zz_4446_ = int_reg_array_6_6_imag;
        _zz_4447_ = int_reg_array_6_6_real;
      end
      6'b000111 : begin
        _zz_4446_ = int_reg_array_6_7_imag;
        _zz_4447_ = int_reg_array_6_7_real;
      end
      6'b001000 : begin
        _zz_4446_ = int_reg_array_6_8_imag;
        _zz_4447_ = int_reg_array_6_8_real;
      end
      6'b001001 : begin
        _zz_4446_ = int_reg_array_6_9_imag;
        _zz_4447_ = int_reg_array_6_9_real;
      end
      6'b001010 : begin
        _zz_4446_ = int_reg_array_6_10_imag;
        _zz_4447_ = int_reg_array_6_10_real;
      end
      6'b001011 : begin
        _zz_4446_ = int_reg_array_6_11_imag;
        _zz_4447_ = int_reg_array_6_11_real;
      end
      6'b001100 : begin
        _zz_4446_ = int_reg_array_6_12_imag;
        _zz_4447_ = int_reg_array_6_12_real;
      end
      6'b001101 : begin
        _zz_4446_ = int_reg_array_6_13_imag;
        _zz_4447_ = int_reg_array_6_13_real;
      end
      6'b001110 : begin
        _zz_4446_ = int_reg_array_6_14_imag;
        _zz_4447_ = int_reg_array_6_14_real;
      end
      6'b001111 : begin
        _zz_4446_ = int_reg_array_6_15_imag;
        _zz_4447_ = int_reg_array_6_15_real;
      end
      6'b010000 : begin
        _zz_4446_ = int_reg_array_6_16_imag;
        _zz_4447_ = int_reg_array_6_16_real;
      end
      6'b010001 : begin
        _zz_4446_ = int_reg_array_6_17_imag;
        _zz_4447_ = int_reg_array_6_17_real;
      end
      6'b010010 : begin
        _zz_4446_ = int_reg_array_6_18_imag;
        _zz_4447_ = int_reg_array_6_18_real;
      end
      6'b010011 : begin
        _zz_4446_ = int_reg_array_6_19_imag;
        _zz_4447_ = int_reg_array_6_19_real;
      end
      6'b010100 : begin
        _zz_4446_ = int_reg_array_6_20_imag;
        _zz_4447_ = int_reg_array_6_20_real;
      end
      6'b010101 : begin
        _zz_4446_ = int_reg_array_6_21_imag;
        _zz_4447_ = int_reg_array_6_21_real;
      end
      6'b010110 : begin
        _zz_4446_ = int_reg_array_6_22_imag;
        _zz_4447_ = int_reg_array_6_22_real;
      end
      6'b010111 : begin
        _zz_4446_ = int_reg_array_6_23_imag;
        _zz_4447_ = int_reg_array_6_23_real;
      end
      6'b011000 : begin
        _zz_4446_ = int_reg_array_6_24_imag;
        _zz_4447_ = int_reg_array_6_24_real;
      end
      6'b011001 : begin
        _zz_4446_ = int_reg_array_6_25_imag;
        _zz_4447_ = int_reg_array_6_25_real;
      end
      6'b011010 : begin
        _zz_4446_ = int_reg_array_6_26_imag;
        _zz_4447_ = int_reg_array_6_26_real;
      end
      6'b011011 : begin
        _zz_4446_ = int_reg_array_6_27_imag;
        _zz_4447_ = int_reg_array_6_27_real;
      end
      6'b011100 : begin
        _zz_4446_ = int_reg_array_6_28_imag;
        _zz_4447_ = int_reg_array_6_28_real;
      end
      6'b011101 : begin
        _zz_4446_ = int_reg_array_6_29_imag;
        _zz_4447_ = int_reg_array_6_29_real;
      end
      6'b011110 : begin
        _zz_4446_ = int_reg_array_6_30_imag;
        _zz_4447_ = int_reg_array_6_30_real;
      end
      6'b011111 : begin
        _zz_4446_ = int_reg_array_6_31_imag;
        _zz_4447_ = int_reg_array_6_31_real;
      end
      6'b100000 : begin
        _zz_4446_ = int_reg_array_6_32_imag;
        _zz_4447_ = int_reg_array_6_32_real;
      end
      6'b100001 : begin
        _zz_4446_ = int_reg_array_6_33_imag;
        _zz_4447_ = int_reg_array_6_33_real;
      end
      6'b100010 : begin
        _zz_4446_ = int_reg_array_6_34_imag;
        _zz_4447_ = int_reg_array_6_34_real;
      end
      6'b100011 : begin
        _zz_4446_ = int_reg_array_6_35_imag;
        _zz_4447_ = int_reg_array_6_35_real;
      end
      6'b100100 : begin
        _zz_4446_ = int_reg_array_6_36_imag;
        _zz_4447_ = int_reg_array_6_36_real;
      end
      6'b100101 : begin
        _zz_4446_ = int_reg_array_6_37_imag;
        _zz_4447_ = int_reg_array_6_37_real;
      end
      6'b100110 : begin
        _zz_4446_ = int_reg_array_6_38_imag;
        _zz_4447_ = int_reg_array_6_38_real;
      end
      6'b100111 : begin
        _zz_4446_ = int_reg_array_6_39_imag;
        _zz_4447_ = int_reg_array_6_39_real;
      end
      6'b101000 : begin
        _zz_4446_ = int_reg_array_6_40_imag;
        _zz_4447_ = int_reg_array_6_40_real;
      end
      6'b101001 : begin
        _zz_4446_ = int_reg_array_6_41_imag;
        _zz_4447_ = int_reg_array_6_41_real;
      end
      6'b101010 : begin
        _zz_4446_ = int_reg_array_6_42_imag;
        _zz_4447_ = int_reg_array_6_42_real;
      end
      6'b101011 : begin
        _zz_4446_ = int_reg_array_6_43_imag;
        _zz_4447_ = int_reg_array_6_43_real;
      end
      6'b101100 : begin
        _zz_4446_ = int_reg_array_6_44_imag;
        _zz_4447_ = int_reg_array_6_44_real;
      end
      6'b101101 : begin
        _zz_4446_ = int_reg_array_6_45_imag;
        _zz_4447_ = int_reg_array_6_45_real;
      end
      6'b101110 : begin
        _zz_4446_ = int_reg_array_6_46_imag;
        _zz_4447_ = int_reg_array_6_46_real;
      end
      6'b101111 : begin
        _zz_4446_ = int_reg_array_6_47_imag;
        _zz_4447_ = int_reg_array_6_47_real;
      end
      6'b110000 : begin
        _zz_4446_ = int_reg_array_6_48_imag;
        _zz_4447_ = int_reg_array_6_48_real;
      end
      6'b110001 : begin
        _zz_4446_ = int_reg_array_6_49_imag;
        _zz_4447_ = int_reg_array_6_49_real;
      end
      6'b110010 : begin
        _zz_4446_ = int_reg_array_6_50_imag;
        _zz_4447_ = int_reg_array_6_50_real;
      end
      6'b110011 : begin
        _zz_4446_ = int_reg_array_6_51_imag;
        _zz_4447_ = int_reg_array_6_51_real;
      end
      6'b110100 : begin
        _zz_4446_ = int_reg_array_6_52_imag;
        _zz_4447_ = int_reg_array_6_52_real;
      end
      6'b110101 : begin
        _zz_4446_ = int_reg_array_6_53_imag;
        _zz_4447_ = int_reg_array_6_53_real;
      end
      6'b110110 : begin
        _zz_4446_ = int_reg_array_6_54_imag;
        _zz_4447_ = int_reg_array_6_54_real;
      end
      6'b110111 : begin
        _zz_4446_ = int_reg_array_6_55_imag;
        _zz_4447_ = int_reg_array_6_55_real;
      end
      6'b111000 : begin
        _zz_4446_ = int_reg_array_6_56_imag;
        _zz_4447_ = int_reg_array_6_56_real;
      end
      6'b111001 : begin
        _zz_4446_ = int_reg_array_6_57_imag;
        _zz_4447_ = int_reg_array_6_57_real;
      end
      6'b111010 : begin
        _zz_4446_ = int_reg_array_6_58_imag;
        _zz_4447_ = int_reg_array_6_58_real;
      end
      6'b111011 : begin
        _zz_4446_ = int_reg_array_6_59_imag;
        _zz_4447_ = int_reg_array_6_59_real;
      end
      6'b111100 : begin
        _zz_4446_ = int_reg_array_6_60_imag;
        _zz_4447_ = int_reg_array_6_60_real;
      end
      6'b111101 : begin
        _zz_4446_ = int_reg_array_6_61_imag;
        _zz_4447_ = int_reg_array_6_61_real;
      end
      6'b111110 : begin
        _zz_4446_ = int_reg_array_6_62_imag;
        _zz_4447_ = int_reg_array_6_62_real;
      end
      default : begin
        _zz_4446_ = int_reg_array_6_63_imag;
        _zz_4447_ = int_reg_array_6_63_real;
      end
    endcase
  end

  always @(*) begin
    case(_zz_500_)
      6'b000000 : begin
        _zz_4448_ = int_reg_array_7_0_imag;
        _zz_4449_ = int_reg_array_7_0_real;
      end
      6'b000001 : begin
        _zz_4448_ = int_reg_array_7_1_imag;
        _zz_4449_ = int_reg_array_7_1_real;
      end
      6'b000010 : begin
        _zz_4448_ = int_reg_array_7_2_imag;
        _zz_4449_ = int_reg_array_7_2_real;
      end
      6'b000011 : begin
        _zz_4448_ = int_reg_array_7_3_imag;
        _zz_4449_ = int_reg_array_7_3_real;
      end
      6'b000100 : begin
        _zz_4448_ = int_reg_array_7_4_imag;
        _zz_4449_ = int_reg_array_7_4_real;
      end
      6'b000101 : begin
        _zz_4448_ = int_reg_array_7_5_imag;
        _zz_4449_ = int_reg_array_7_5_real;
      end
      6'b000110 : begin
        _zz_4448_ = int_reg_array_7_6_imag;
        _zz_4449_ = int_reg_array_7_6_real;
      end
      6'b000111 : begin
        _zz_4448_ = int_reg_array_7_7_imag;
        _zz_4449_ = int_reg_array_7_7_real;
      end
      6'b001000 : begin
        _zz_4448_ = int_reg_array_7_8_imag;
        _zz_4449_ = int_reg_array_7_8_real;
      end
      6'b001001 : begin
        _zz_4448_ = int_reg_array_7_9_imag;
        _zz_4449_ = int_reg_array_7_9_real;
      end
      6'b001010 : begin
        _zz_4448_ = int_reg_array_7_10_imag;
        _zz_4449_ = int_reg_array_7_10_real;
      end
      6'b001011 : begin
        _zz_4448_ = int_reg_array_7_11_imag;
        _zz_4449_ = int_reg_array_7_11_real;
      end
      6'b001100 : begin
        _zz_4448_ = int_reg_array_7_12_imag;
        _zz_4449_ = int_reg_array_7_12_real;
      end
      6'b001101 : begin
        _zz_4448_ = int_reg_array_7_13_imag;
        _zz_4449_ = int_reg_array_7_13_real;
      end
      6'b001110 : begin
        _zz_4448_ = int_reg_array_7_14_imag;
        _zz_4449_ = int_reg_array_7_14_real;
      end
      6'b001111 : begin
        _zz_4448_ = int_reg_array_7_15_imag;
        _zz_4449_ = int_reg_array_7_15_real;
      end
      6'b010000 : begin
        _zz_4448_ = int_reg_array_7_16_imag;
        _zz_4449_ = int_reg_array_7_16_real;
      end
      6'b010001 : begin
        _zz_4448_ = int_reg_array_7_17_imag;
        _zz_4449_ = int_reg_array_7_17_real;
      end
      6'b010010 : begin
        _zz_4448_ = int_reg_array_7_18_imag;
        _zz_4449_ = int_reg_array_7_18_real;
      end
      6'b010011 : begin
        _zz_4448_ = int_reg_array_7_19_imag;
        _zz_4449_ = int_reg_array_7_19_real;
      end
      6'b010100 : begin
        _zz_4448_ = int_reg_array_7_20_imag;
        _zz_4449_ = int_reg_array_7_20_real;
      end
      6'b010101 : begin
        _zz_4448_ = int_reg_array_7_21_imag;
        _zz_4449_ = int_reg_array_7_21_real;
      end
      6'b010110 : begin
        _zz_4448_ = int_reg_array_7_22_imag;
        _zz_4449_ = int_reg_array_7_22_real;
      end
      6'b010111 : begin
        _zz_4448_ = int_reg_array_7_23_imag;
        _zz_4449_ = int_reg_array_7_23_real;
      end
      6'b011000 : begin
        _zz_4448_ = int_reg_array_7_24_imag;
        _zz_4449_ = int_reg_array_7_24_real;
      end
      6'b011001 : begin
        _zz_4448_ = int_reg_array_7_25_imag;
        _zz_4449_ = int_reg_array_7_25_real;
      end
      6'b011010 : begin
        _zz_4448_ = int_reg_array_7_26_imag;
        _zz_4449_ = int_reg_array_7_26_real;
      end
      6'b011011 : begin
        _zz_4448_ = int_reg_array_7_27_imag;
        _zz_4449_ = int_reg_array_7_27_real;
      end
      6'b011100 : begin
        _zz_4448_ = int_reg_array_7_28_imag;
        _zz_4449_ = int_reg_array_7_28_real;
      end
      6'b011101 : begin
        _zz_4448_ = int_reg_array_7_29_imag;
        _zz_4449_ = int_reg_array_7_29_real;
      end
      6'b011110 : begin
        _zz_4448_ = int_reg_array_7_30_imag;
        _zz_4449_ = int_reg_array_7_30_real;
      end
      6'b011111 : begin
        _zz_4448_ = int_reg_array_7_31_imag;
        _zz_4449_ = int_reg_array_7_31_real;
      end
      6'b100000 : begin
        _zz_4448_ = int_reg_array_7_32_imag;
        _zz_4449_ = int_reg_array_7_32_real;
      end
      6'b100001 : begin
        _zz_4448_ = int_reg_array_7_33_imag;
        _zz_4449_ = int_reg_array_7_33_real;
      end
      6'b100010 : begin
        _zz_4448_ = int_reg_array_7_34_imag;
        _zz_4449_ = int_reg_array_7_34_real;
      end
      6'b100011 : begin
        _zz_4448_ = int_reg_array_7_35_imag;
        _zz_4449_ = int_reg_array_7_35_real;
      end
      6'b100100 : begin
        _zz_4448_ = int_reg_array_7_36_imag;
        _zz_4449_ = int_reg_array_7_36_real;
      end
      6'b100101 : begin
        _zz_4448_ = int_reg_array_7_37_imag;
        _zz_4449_ = int_reg_array_7_37_real;
      end
      6'b100110 : begin
        _zz_4448_ = int_reg_array_7_38_imag;
        _zz_4449_ = int_reg_array_7_38_real;
      end
      6'b100111 : begin
        _zz_4448_ = int_reg_array_7_39_imag;
        _zz_4449_ = int_reg_array_7_39_real;
      end
      6'b101000 : begin
        _zz_4448_ = int_reg_array_7_40_imag;
        _zz_4449_ = int_reg_array_7_40_real;
      end
      6'b101001 : begin
        _zz_4448_ = int_reg_array_7_41_imag;
        _zz_4449_ = int_reg_array_7_41_real;
      end
      6'b101010 : begin
        _zz_4448_ = int_reg_array_7_42_imag;
        _zz_4449_ = int_reg_array_7_42_real;
      end
      6'b101011 : begin
        _zz_4448_ = int_reg_array_7_43_imag;
        _zz_4449_ = int_reg_array_7_43_real;
      end
      6'b101100 : begin
        _zz_4448_ = int_reg_array_7_44_imag;
        _zz_4449_ = int_reg_array_7_44_real;
      end
      6'b101101 : begin
        _zz_4448_ = int_reg_array_7_45_imag;
        _zz_4449_ = int_reg_array_7_45_real;
      end
      6'b101110 : begin
        _zz_4448_ = int_reg_array_7_46_imag;
        _zz_4449_ = int_reg_array_7_46_real;
      end
      6'b101111 : begin
        _zz_4448_ = int_reg_array_7_47_imag;
        _zz_4449_ = int_reg_array_7_47_real;
      end
      6'b110000 : begin
        _zz_4448_ = int_reg_array_7_48_imag;
        _zz_4449_ = int_reg_array_7_48_real;
      end
      6'b110001 : begin
        _zz_4448_ = int_reg_array_7_49_imag;
        _zz_4449_ = int_reg_array_7_49_real;
      end
      6'b110010 : begin
        _zz_4448_ = int_reg_array_7_50_imag;
        _zz_4449_ = int_reg_array_7_50_real;
      end
      6'b110011 : begin
        _zz_4448_ = int_reg_array_7_51_imag;
        _zz_4449_ = int_reg_array_7_51_real;
      end
      6'b110100 : begin
        _zz_4448_ = int_reg_array_7_52_imag;
        _zz_4449_ = int_reg_array_7_52_real;
      end
      6'b110101 : begin
        _zz_4448_ = int_reg_array_7_53_imag;
        _zz_4449_ = int_reg_array_7_53_real;
      end
      6'b110110 : begin
        _zz_4448_ = int_reg_array_7_54_imag;
        _zz_4449_ = int_reg_array_7_54_real;
      end
      6'b110111 : begin
        _zz_4448_ = int_reg_array_7_55_imag;
        _zz_4449_ = int_reg_array_7_55_real;
      end
      6'b111000 : begin
        _zz_4448_ = int_reg_array_7_56_imag;
        _zz_4449_ = int_reg_array_7_56_real;
      end
      6'b111001 : begin
        _zz_4448_ = int_reg_array_7_57_imag;
        _zz_4449_ = int_reg_array_7_57_real;
      end
      6'b111010 : begin
        _zz_4448_ = int_reg_array_7_58_imag;
        _zz_4449_ = int_reg_array_7_58_real;
      end
      6'b111011 : begin
        _zz_4448_ = int_reg_array_7_59_imag;
        _zz_4449_ = int_reg_array_7_59_real;
      end
      6'b111100 : begin
        _zz_4448_ = int_reg_array_7_60_imag;
        _zz_4449_ = int_reg_array_7_60_real;
      end
      6'b111101 : begin
        _zz_4448_ = int_reg_array_7_61_imag;
        _zz_4449_ = int_reg_array_7_61_real;
      end
      6'b111110 : begin
        _zz_4448_ = int_reg_array_7_62_imag;
        _zz_4449_ = int_reg_array_7_62_real;
      end
      default : begin
        _zz_4448_ = int_reg_array_7_63_imag;
        _zz_4449_ = int_reg_array_7_63_real;
      end
    endcase
  end

  always @(*) begin
    case(_zz_569_)
      6'b000000 : begin
        _zz_4450_ = int_reg_array_8_0_imag;
        _zz_4451_ = int_reg_array_8_0_real;
      end
      6'b000001 : begin
        _zz_4450_ = int_reg_array_8_1_imag;
        _zz_4451_ = int_reg_array_8_1_real;
      end
      6'b000010 : begin
        _zz_4450_ = int_reg_array_8_2_imag;
        _zz_4451_ = int_reg_array_8_2_real;
      end
      6'b000011 : begin
        _zz_4450_ = int_reg_array_8_3_imag;
        _zz_4451_ = int_reg_array_8_3_real;
      end
      6'b000100 : begin
        _zz_4450_ = int_reg_array_8_4_imag;
        _zz_4451_ = int_reg_array_8_4_real;
      end
      6'b000101 : begin
        _zz_4450_ = int_reg_array_8_5_imag;
        _zz_4451_ = int_reg_array_8_5_real;
      end
      6'b000110 : begin
        _zz_4450_ = int_reg_array_8_6_imag;
        _zz_4451_ = int_reg_array_8_6_real;
      end
      6'b000111 : begin
        _zz_4450_ = int_reg_array_8_7_imag;
        _zz_4451_ = int_reg_array_8_7_real;
      end
      6'b001000 : begin
        _zz_4450_ = int_reg_array_8_8_imag;
        _zz_4451_ = int_reg_array_8_8_real;
      end
      6'b001001 : begin
        _zz_4450_ = int_reg_array_8_9_imag;
        _zz_4451_ = int_reg_array_8_9_real;
      end
      6'b001010 : begin
        _zz_4450_ = int_reg_array_8_10_imag;
        _zz_4451_ = int_reg_array_8_10_real;
      end
      6'b001011 : begin
        _zz_4450_ = int_reg_array_8_11_imag;
        _zz_4451_ = int_reg_array_8_11_real;
      end
      6'b001100 : begin
        _zz_4450_ = int_reg_array_8_12_imag;
        _zz_4451_ = int_reg_array_8_12_real;
      end
      6'b001101 : begin
        _zz_4450_ = int_reg_array_8_13_imag;
        _zz_4451_ = int_reg_array_8_13_real;
      end
      6'b001110 : begin
        _zz_4450_ = int_reg_array_8_14_imag;
        _zz_4451_ = int_reg_array_8_14_real;
      end
      6'b001111 : begin
        _zz_4450_ = int_reg_array_8_15_imag;
        _zz_4451_ = int_reg_array_8_15_real;
      end
      6'b010000 : begin
        _zz_4450_ = int_reg_array_8_16_imag;
        _zz_4451_ = int_reg_array_8_16_real;
      end
      6'b010001 : begin
        _zz_4450_ = int_reg_array_8_17_imag;
        _zz_4451_ = int_reg_array_8_17_real;
      end
      6'b010010 : begin
        _zz_4450_ = int_reg_array_8_18_imag;
        _zz_4451_ = int_reg_array_8_18_real;
      end
      6'b010011 : begin
        _zz_4450_ = int_reg_array_8_19_imag;
        _zz_4451_ = int_reg_array_8_19_real;
      end
      6'b010100 : begin
        _zz_4450_ = int_reg_array_8_20_imag;
        _zz_4451_ = int_reg_array_8_20_real;
      end
      6'b010101 : begin
        _zz_4450_ = int_reg_array_8_21_imag;
        _zz_4451_ = int_reg_array_8_21_real;
      end
      6'b010110 : begin
        _zz_4450_ = int_reg_array_8_22_imag;
        _zz_4451_ = int_reg_array_8_22_real;
      end
      6'b010111 : begin
        _zz_4450_ = int_reg_array_8_23_imag;
        _zz_4451_ = int_reg_array_8_23_real;
      end
      6'b011000 : begin
        _zz_4450_ = int_reg_array_8_24_imag;
        _zz_4451_ = int_reg_array_8_24_real;
      end
      6'b011001 : begin
        _zz_4450_ = int_reg_array_8_25_imag;
        _zz_4451_ = int_reg_array_8_25_real;
      end
      6'b011010 : begin
        _zz_4450_ = int_reg_array_8_26_imag;
        _zz_4451_ = int_reg_array_8_26_real;
      end
      6'b011011 : begin
        _zz_4450_ = int_reg_array_8_27_imag;
        _zz_4451_ = int_reg_array_8_27_real;
      end
      6'b011100 : begin
        _zz_4450_ = int_reg_array_8_28_imag;
        _zz_4451_ = int_reg_array_8_28_real;
      end
      6'b011101 : begin
        _zz_4450_ = int_reg_array_8_29_imag;
        _zz_4451_ = int_reg_array_8_29_real;
      end
      6'b011110 : begin
        _zz_4450_ = int_reg_array_8_30_imag;
        _zz_4451_ = int_reg_array_8_30_real;
      end
      6'b011111 : begin
        _zz_4450_ = int_reg_array_8_31_imag;
        _zz_4451_ = int_reg_array_8_31_real;
      end
      6'b100000 : begin
        _zz_4450_ = int_reg_array_8_32_imag;
        _zz_4451_ = int_reg_array_8_32_real;
      end
      6'b100001 : begin
        _zz_4450_ = int_reg_array_8_33_imag;
        _zz_4451_ = int_reg_array_8_33_real;
      end
      6'b100010 : begin
        _zz_4450_ = int_reg_array_8_34_imag;
        _zz_4451_ = int_reg_array_8_34_real;
      end
      6'b100011 : begin
        _zz_4450_ = int_reg_array_8_35_imag;
        _zz_4451_ = int_reg_array_8_35_real;
      end
      6'b100100 : begin
        _zz_4450_ = int_reg_array_8_36_imag;
        _zz_4451_ = int_reg_array_8_36_real;
      end
      6'b100101 : begin
        _zz_4450_ = int_reg_array_8_37_imag;
        _zz_4451_ = int_reg_array_8_37_real;
      end
      6'b100110 : begin
        _zz_4450_ = int_reg_array_8_38_imag;
        _zz_4451_ = int_reg_array_8_38_real;
      end
      6'b100111 : begin
        _zz_4450_ = int_reg_array_8_39_imag;
        _zz_4451_ = int_reg_array_8_39_real;
      end
      6'b101000 : begin
        _zz_4450_ = int_reg_array_8_40_imag;
        _zz_4451_ = int_reg_array_8_40_real;
      end
      6'b101001 : begin
        _zz_4450_ = int_reg_array_8_41_imag;
        _zz_4451_ = int_reg_array_8_41_real;
      end
      6'b101010 : begin
        _zz_4450_ = int_reg_array_8_42_imag;
        _zz_4451_ = int_reg_array_8_42_real;
      end
      6'b101011 : begin
        _zz_4450_ = int_reg_array_8_43_imag;
        _zz_4451_ = int_reg_array_8_43_real;
      end
      6'b101100 : begin
        _zz_4450_ = int_reg_array_8_44_imag;
        _zz_4451_ = int_reg_array_8_44_real;
      end
      6'b101101 : begin
        _zz_4450_ = int_reg_array_8_45_imag;
        _zz_4451_ = int_reg_array_8_45_real;
      end
      6'b101110 : begin
        _zz_4450_ = int_reg_array_8_46_imag;
        _zz_4451_ = int_reg_array_8_46_real;
      end
      6'b101111 : begin
        _zz_4450_ = int_reg_array_8_47_imag;
        _zz_4451_ = int_reg_array_8_47_real;
      end
      6'b110000 : begin
        _zz_4450_ = int_reg_array_8_48_imag;
        _zz_4451_ = int_reg_array_8_48_real;
      end
      6'b110001 : begin
        _zz_4450_ = int_reg_array_8_49_imag;
        _zz_4451_ = int_reg_array_8_49_real;
      end
      6'b110010 : begin
        _zz_4450_ = int_reg_array_8_50_imag;
        _zz_4451_ = int_reg_array_8_50_real;
      end
      6'b110011 : begin
        _zz_4450_ = int_reg_array_8_51_imag;
        _zz_4451_ = int_reg_array_8_51_real;
      end
      6'b110100 : begin
        _zz_4450_ = int_reg_array_8_52_imag;
        _zz_4451_ = int_reg_array_8_52_real;
      end
      6'b110101 : begin
        _zz_4450_ = int_reg_array_8_53_imag;
        _zz_4451_ = int_reg_array_8_53_real;
      end
      6'b110110 : begin
        _zz_4450_ = int_reg_array_8_54_imag;
        _zz_4451_ = int_reg_array_8_54_real;
      end
      6'b110111 : begin
        _zz_4450_ = int_reg_array_8_55_imag;
        _zz_4451_ = int_reg_array_8_55_real;
      end
      6'b111000 : begin
        _zz_4450_ = int_reg_array_8_56_imag;
        _zz_4451_ = int_reg_array_8_56_real;
      end
      6'b111001 : begin
        _zz_4450_ = int_reg_array_8_57_imag;
        _zz_4451_ = int_reg_array_8_57_real;
      end
      6'b111010 : begin
        _zz_4450_ = int_reg_array_8_58_imag;
        _zz_4451_ = int_reg_array_8_58_real;
      end
      6'b111011 : begin
        _zz_4450_ = int_reg_array_8_59_imag;
        _zz_4451_ = int_reg_array_8_59_real;
      end
      6'b111100 : begin
        _zz_4450_ = int_reg_array_8_60_imag;
        _zz_4451_ = int_reg_array_8_60_real;
      end
      6'b111101 : begin
        _zz_4450_ = int_reg_array_8_61_imag;
        _zz_4451_ = int_reg_array_8_61_real;
      end
      6'b111110 : begin
        _zz_4450_ = int_reg_array_8_62_imag;
        _zz_4451_ = int_reg_array_8_62_real;
      end
      default : begin
        _zz_4450_ = int_reg_array_8_63_imag;
        _zz_4451_ = int_reg_array_8_63_real;
      end
    endcase
  end

  always @(*) begin
    case(_zz_638_)
      6'b000000 : begin
        _zz_4452_ = int_reg_array_9_0_imag;
        _zz_4453_ = int_reg_array_9_0_real;
      end
      6'b000001 : begin
        _zz_4452_ = int_reg_array_9_1_imag;
        _zz_4453_ = int_reg_array_9_1_real;
      end
      6'b000010 : begin
        _zz_4452_ = int_reg_array_9_2_imag;
        _zz_4453_ = int_reg_array_9_2_real;
      end
      6'b000011 : begin
        _zz_4452_ = int_reg_array_9_3_imag;
        _zz_4453_ = int_reg_array_9_3_real;
      end
      6'b000100 : begin
        _zz_4452_ = int_reg_array_9_4_imag;
        _zz_4453_ = int_reg_array_9_4_real;
      end
      6'b000101 : begin
        _zz_4452_ = int_reg_array_9_5_imag;
        _zz_4453_ = int_reg_array_9_5_real;
      end
      6'b000110 : begin
        _zz_4452_ = int_reg_array_9_6_imag;
        _zz_4453_ = int_reg_array_9_6_real;
      end
      6'b000111 : begin
        _zz_4452_ = int_reg_array_9_7_imag;
        _zz_4453_ = int_reg_array_9_7_real;
      end
      6'b001000 : begin
        _zz_4452_ = int_reg_array_9_8_imag;
        _zz_4453_ = int_reg_array_9_8_real;
      end
      6'b001001 : begin
        _zz_4452_ = int_reg_array_9_9_imag;
        _zz_4453_ = int_reg_array_9_9_real;
      end
      6'b001010 : begin
        _zz_4452_ = int_reg_array_9_10_imag;
        _zz_4453_ = int_reg_array_9_10_real;
      end
      6'b001011 : begin
        _zz_4452_ = int_reg_array_9_11_imag;
        _zz_4453_ = int_reg_array_9_11_real;
      end
      6'b001100 : begin
        _zz_4452_ = int_reg_array_9_12_imag;
        _zz_4453_ = int_reg_array_9_12_real;
      end
      6'b001101 : begin
        _zz_4452_ = int_reg_array_9_13_imag;
        _zz_4453_ = int_reg_array_9_13_real;
      end
      6'b001110 : begin
        _zz_4452_ = int_reg_array_9_14_imag;
        _zz_4453_ = int_reg_array_9_14_real;
      end
      6'b001111 : begin
        _zz_4452_ = int_reg_array_9_15_imag;
        _zz_4453_ = int_reg_array_9_15_real;
      end
      6'b010000 : begin
        _zz_4452_ = int_reg_array_9_16_imag;
        _zz_4453_ = int_reg_array_9_16_real;
      end
      6'b010001 : begin
        _zz_4452_ = int_reg_array_9_17_imag;
        _zz_4453_ = int_reg_array_9_17_real;
      end
      6'b010010 : begin
        _zz_4452_ = int_reg_array_9_18_imag;
        _zz_4453_ = int_reg_array_9_18_real;
      end
      6'b010011 : begin
        _zz_4452_ = int_reg_array_9_19_imag;
        _zz_4453_ = int_reg_array_9_19_real;
      end
      6'b010100 : begin
        _zz_4452_ = int_reg_array_9_20_imag;
        _zz_4453_ = int_reg_array_9_20_real;
      end
      6'b010101 : begin
        _zz_4452_ = int_reg_array_9_21_imag;
        _zz_4453_ = int_reg_array_9_21_real;
      end
      6'b010110 : begin
        _zz_4452_ = int_reg_array_9_22_imag;
        _zz_4453_ = int_reg_array_9_22_real;
      end
      6'b010111 : begin
        _zz_4452_ = int_reg_array_9_23_imag;
        _zz_4453_ = int_reg_array_9_23_real;
      end
      6'b011000 : begin
        _zz_4452_ = int_reg_array_9_24_imag;
        _zz_4453_ = int_reg_array_9_24_real;
      end
      6'b011001 : begin
        _zz_4452_ = int_reg_array_9_25_imag;
        _zz_4453_ = int_reg_array_9_25_real;
      end
      6'b011010 : begin
        _zz_4452_ = int_reg_array_9_26_imag;
        _zz_4453_ = int_reg_array_9_26_real;
      end
      6'b011011 : begin
        _zz_4452_ = int_reg_array_9_27_imag;
        _zz_4453_ = int_reg_array_9_27_real;
      end
      6'b011100 : begin
        _zz_4452_ = int_reg_array_9_28_imag;
        _zz_4453_ = int_reg_array_9_28_real;
      end
      6'b011101 : begin
        _zz_4452_ = int_reg_array_9_29_imag;
        _zz_4453_ = int_reg_array_9_29_real;
      end
      6'b011110 : begin
        _zz_4452_ = int_reg_array_9_30_imag;
        _zz_4453_ = int_reg_array_9_30_real;
      end
      6'b011111 : begin
        _zz_4452_ = int_reg_array_9_31_imag;
        _zz_4453_ = int_reg_array_9_31_real;
      end
      6'b100000 : begin
        _zz_4452_ = int_reg_array_9_32_imag;
        _zz_4453_ = int_reg_array_9_32_real;
      end
      6'b100001 : begin
        _zz_4452_ = int_reg_array_9_33_imag;
        _zz_4453_ = int_reg_array_9_33_real;
      end
      6'b100010 : begin
        _zz_4452_ = int_reg_array_9_34_imag;
        _zz_4453_ = int_reg_array_9_34_real;
      end
      6'b100011 : begin
        _zz_4452_ = int_reg_array_9_35_imag;
        _zz_4453_ = int_reg_array_9_35_real;
      end
      6'b100100 : begin
        _zz_4452_ = int_reg_array_9_36_imag;
        _zz_4453_ = int_reg_array_9_36_real;
      end
      6'b100101 : begin
        _zz_4452_ = int_reg_array_9_37_imag;
        _zz_4453_ = int_reg_array_9_37_real;
      end
      6'b100110 : begin
        _zz_4452_ = int_reg_array_9_38_imag;
        _zz_4453_ = int_reg_array_9_38_real;
      end
      6'b100111 : begin
        _zz_4452_ = int_reg_array_9_39_imag;
        _zz_4453_ = int_reg_array_9_39_real;
      end
      6'b101000 : begin
        _zz_4452_ = int_reg_array_9_40_imag;
        _zz_4453_ = int_reg_array_9_40_real;
      end
      6'b101001 : begin
        _zz_4452_ = int_reg_array_9_41_imag;
        _zz_4453_ = int_reg_array_9_41_real;
      end
      6'b101010 : begin
        _zz_4452_ = int_reg_array_9_42_imag;
        _zz_4453_ = int_reg_array_9_42_real;
      end
      6'b101011 : begin
        _zz_4452_ = int_reg_array_9_43_imag;
        _zz_4453_ = int_reg_array_9_43_real;
      end
      6'b101100 : begin
        _zz_4452_ = int_reg_array_9_44_imag;
        _zz_4453_ = int_reg_array_9_44_real;
      end
      6'b101101 : begin
        _zz_4452_ = int_reg_array_9_45_imag;
        _zz_4453_ = int_reg_array_9_45_real;
      end
      6'b101110 : begin
        _zz_4452_ = int_reg_array_9_46_imag;
        _zz_4453_ = int_reg_array_9_46_real;
      end
      6'b101111 : begin
        _zz_4452_ = int_reg_array_9_47_imag;
        _zz_4453_ = int_reg_array_9_47_real;
      end
      6'b110000 : begin
        _zz_4452_ = int_reg_array_9_48_imag;
        _zz_4453_ = int_reg_array_9_48_real;
      end
      6'b110001 : begin
        _zz_4452_ = int_reg_array_9_49_imag;
        _zz_4453_ = int_reg_array_9_49_real;
      end
      6'b110010 : begin
        _zz_4452_ = int_reg_array_9_50_imag;
        _zz_4453_ = int_reg_array_9_50_real;
      end
      6'b110011 : begin
        _zz_4452_ = int_reg_array_9_51_imag;
        _zz_4453_ = int_reg_array_9_51_real;
      end
      6'b110100 : begin
        _zz_4452_ = int_reg_array_9_52_imag;
        _zz_4453_ = int_reg_array_9_52_real;
      end
      6'b110101 : begin
        _zz_4452_ = int_reg_array_9_53_imag;
        _zz_4453_ = int_reg_array_9_53_real;
      end
      6'b110110 : begin
        _zz_4452_ = int_reg_array_9_54_imag;
        _zz_4453_ = int_reg_array_9_54_real;
      end
      6'b110111 : begin
        _zz_4452_ = int_reg_array_9_55_imag;
        _zz_4453_ = int_reg_array_9_55_real;
      end
      6'b111000 : begin
        _zz_4452_ = int_reg_array_9_56_imag;
        _zz_4453_ = int_reg_array_9_56_real;
      end
      6'b111001 : begin
        _zz_4452_ = int_reg_array_9_57_imag;
        _zz_4453_ = int_reg_array_9_57_real;
      end
      6'b111010 : begin
        _zz_4452_ = int_reg_array_9_58_imag;
        _zz_4453_ = int_reg_array_9_58_real;
      end
      6'b111011 : begin
        _zz_4452_ = int_reg_array_9_59_imag;
        _zz_4453_ = int_reg_array_9_59_real;
      end
      6'b111100 : begin
        _zz_4452_ = int_reg_array_9_60_imag;
        _zz_4453_ = int_reg_array_9_60_real;
      end
      6'b111101 : begin
        _zz_4452_ = int_reg_array_9_61_imag;
        _zz_4453_ = int_reg_array_9_61_real;
      end
      6'b111110 : begin
        _zz_4452_ = int_reg_array_9_62_imag;
        _zz_4453_ = int_reg_array_9_62_real;
      end
      default : begin
        _zz_4452_ = int_reg_array_9_63_imag;
        _zz_4453_ = int_reg_array_9_63_real;
      end
    endcase
  end

  always @(*) begin
    case(_zz_707_)
      6'b000000 : begin
        _zz_4454_ = int_reg_array_10_0_imag;
        _zz_4455_ = int_reg_array_10_0_real;
      end
      6'b000001 : begin
        _zz_4454_ = int_reg_array_10_1_imag;
        _zz_4455_ = int_reg_array_10_1_real;
      end
      6'b000010 : begin
        _zz_4454_ = int_reg_array_10_2_imag;
        _zz_4455_ = int_reg_array_10_2_real;
      end
      6'b000011 : begin
        _zz_4454_ = int_reg_array_10_3_imag;
        _zz_4455_ = int_reg_array_10_3_real;
      end
      6'b000100 : begin
        _zz_4454_ = int_reg_array_10_4_imag;
        _zz_4455_ = int_reg_array_10_4_real;
      end
      6'b000101 : begin
        _zz_4454_ = int_reg_array_10_5_imag;
        _zz_4455_ = int_reg_array_10_5_real;
      end
      6'b000110 : begin
        _zz_4454_ = int_reg_array_10_6_imag;
        _zz_4455_ = int_reg_array_10_6_real;
      end
      6'b000111 : begin
        _zz_4454_ = int_reg_array_10_7_imag;
        _zz_4455_ = int_reg_array_10_7_real;
      end
      6'b001000 : begin
        _zz_4454_ = int_reg_array_10_8_imag;
        _zz_4455_ = int_reg_array_10_8_real;
      end
      6'b001001 : begin
        _zz_4454_ = int_reg_array_10_9_imag;
        _zz_4455_ = int_reg_array_10_9_real;
      end
      6'b001010 : begin
        _zz_4454_ = int_reg_array_10_10_imag;
        _zz_4455_ = int_reg_array_10_10_real;
      end
      6'b001011 : begin
        _zz_4454_ = int_reg_array_10_11_imag;
        _zz_4455_ = int_reg_array_10_11_real;
      end
      6'b001100 : begin
        _zz_4454_ = int_reg_array_10_12_imag;
        _zz_4455_ = int_reg_array_10_12_real;
      end
      6'b001101 : begin
        _zz_4454_ = int_reg_array_10_13_imag;
        _zz_4455_ = int_reg_array_10_13_real;
      end
      6'b001110 : begin
        _zz_4454_ = int_reg_array_10_14_imag;
        _zz_4455_ = int_reg_array_10_14_real;
      end
      6'b001111 : begin
        _zz_4454_ = int_reg_array_10_15_imag;
        _zz_4455_ = int_reg_array_10_15_real;
      end
      6'b010000 : begin
        _zz_4454_ = int_reg_array_10_16_imag;
        _zz_4455_ = int_reg_array_10_16_real;
      end
      6'b010001 : begin
        _zz_4454_ = int_reg_array_10_17_imag;
        _zz_4455_ = int_reg_array_10_17_real;
      end
      6'b010010 : begin
        _zz_4454_ = int_reg_array_10_18_imag;
        _zz_4455_ = int_reg_array_10_18_real;
      end
      6'b010011 : begin
        _zz_4454_ = int_reg_array_10_19_imag;
        _zz_4455_ = int_reg_array_10_19_real;
      end
      6'b010100 : begin
        _zz_4454_ = int_reg_array_10_20_imag;
        _zz_4455_ = int_reg_array_10_20_real;
      end
      6'b010101 : begin
        _zz_4454_ = int_reg_array_10_21_imag;
        _zz_4455_ = int_reg_array_10_21_real;
      end
      6'b010110 : begin
        _zz_4454_ = int_reg_array_10_22_imag;
        _zz_4455_ = int_reg_array_10_22_real;
      end
      6'b010111 : begin
        _zz_4454_ = int_reg_array_10_23_imag;
        _zz_4455_ = int_reg_array_10_23_real;
      end
      6'b011000 : begin
        _zz_4454_ = int_reg_array_10_24_imag;
        _zz_4455_ = int_reg_array_10_24_real;
      end
      6'b011001 : begin
        _zz_4454_ = int_reg_array_10_25_imag;
        _zz_4455_ = int_reg_array_10_25_real;
      end
      6'b011010 : begin
        _zz_4454_ = int_reg_array_10_26_imag;
        _zz_4455_ = int_reg_array_10_26_real;
      end
      6'b011011 : begin
        _zz_4454_ = int_reg_array_10_27_imag;
        _zz_4455_ = int_reg_array_10_27_real;
      end
      6'b011100 : begin
        _zz_4454_ = int_reg_array_10_28_imag;
        _zz_4455_ = int_reg_array_10_28_real;
      end
      6'b011101 : begin
        _zz_4454_ = int_reg_array_10_29_imag;
        _zz_4455_ = int_reg_array_10_29_real;
      end
      6'b011110 : begin
        _zz_4454_ = int_reg_array_10_30_imag;
        _zz_4455_ = int_reg_array_10_30_real;
      end
      6'b011111 : begin
        _zz_4454_ = int_reg_array_10_31_imag;
        _zz_4455_ = int_reg_array_10_31_real;
      end
      6'b100000 : begin
        _zz_4454_ = int_reg_array_10_32_imag;
        _zz_4455_ = int_reg_array_10_32_real;
      end
      6'b100001 : begin
        _zz_4454_ = int_reg_array_10_33_imag;
        _zz_4455_ = int_reg_array_10_33_real;
      end
      6'b100010 : begin
        _zz_4454_ = int_reg_array_10_34_imag;
        _zz_4455_ = int_reg_array_10_34_real;
      end
      6'b100011 : begin
        _zz_4454_ = int_reg_array_10_35_imag;
        _zz_4455_ = int_reg_array_10_35_real;
      end
      6'b100100 : begin
        _zz_4454_ = int_reg_array_10_36_imag;
        _zz_4455_ = int_reg_array_10_36_real;
      end
      6'b100101 : begin
        _zz_4454_ = int_reg_array_10_37_imag;
        _zz_4455_ = int_reg_array_10_37_real;
      end
      6'b100110 : begin
        _zz_4454_ = int_reg_array_10_38_imag;
        _zz_4455_ = int_reg_array_10_38_real;
      end
      6'b100111 : begin
        _zz_4454_ = int_reg_array_10_39_imag;
        _zz_4455_ = int_reg_array_10_39_real;
      end
      6'b101000 : begin
        _zz_4454_ = int_reg_array_10_40_imag;
        _zz_4455_ = int_reg_array_10_40_real;
      end
      6'b101001 : begin
        _zz_4454_ = int_reg_array_10_41_imag;
        _zz_4455_ = int_reg_array_10_41_real;
      end
      6'b101010 : begin
        _zz_4454_ = int_reg_array_10_42_imag;
        _zz_4455_ = int_reg_array_10_42_real;
      end
      6'b101011 : begin
        _zz_4454_ = int_reg_array_10_43_imag;
        _zz_4455_ = int_reg_array_10_43_real;
      end
      6'b101100 : begin
        _zz_4454_ = int_reg_array_10_44_imag;
        _zz_4455_ = int_reg_array_10_44_real;
      end
      6'b101101 : begin
        _zz_4454_ = int_reg_array_10_45_imag;
        _zz_4455_ = int_reg_array_10_45_real;
      end
      6'b101110 : begin
        _zz_4454_ = int_reg_array_10_46_imag;
        _zz_4455_ = int_reg_array_10_46_real;
      end
      6'b101111 : begin
        _zz_4454_ = int_reg_array_10_47_imag;
        _zz_4455_ = int_reg_array_10_47_real;
      end
      6'b110000 : begin
        _zz_4454_ = int_reg_array_10_48_imag;
        _zz_4455_ = int_reg_array_10_48_real;
      end
      6'b110001 : begin
        _zz_4454_ = int_reg_array_10_49_imag;
        _zz_4455_ = int_reg_array_10_49_real;
      end
      6'b110010 : begin
        _zz_4454_ = int_reg_array_10_50_imag;
        _zz_4455_ = int_reg_array_10_50_real;
      end
      6'b110011 : begin
        _zz_4454_ = int_reg_array_10_51_imag;
        _zz_4455_ = int_reg_array_10_51_real;
      end
      6'b110100 : begin
        _zz_4454_ = int_reg_array_10_52_imag;
        _zz_4455_ = int_reg_array_10_52_real;
      end
      6'b110101 : begin
        _zz_4454_ = int_reg_array_10_53_imag;
        _zz_4455_ = int_reg_array_10_53_real;
      end
      6'b110110 : begin
        _zz_4454_ = int_reg_array_10_54_imag;
        _zz_4455_ = int_reg_array_10_54_real;
      end
      6'b110111 : begin
        _zz_4454_ = int_reg_array_10_55_imag;
        _zz_4455_ = int_reg_array_10_55_real;
      end
      6'b111000 : begin
        _zz_4454_ = int_reg_array_10_56_imag;
        _zz_4455_ = int_reg_array_10_56_real;
      end
      6'b111001 : begin
        _zz_4454_ = int_reg_array_10_57_imag;
        _zz_4455_ = int_reg_array_10_57_real;
      end
      6'b111010 : begin
        _zz_4454_ = int_reg_array_10_58_imag;
        _zz_4455_ = int_reg_array_10_58_real;
      end
      6'b111011 : begin
        _zz_4454_ = int_reg_array_10_59_imag;
        _zz_4455_ = int_reg_array_10_59_real;
      end
      6'b111100 : begin
        _zz_4454_ = int_reg_array_10_60_imag;
        _zz_4455_ = int_reg_array_10_60_real;
      end
      6'b111101 : begin
        _zz_4454_ = int_reg_array_10_61_imag;
        _zz_4455_ = int_reg_array_10_61_real;
      end
      6'b111110 : begin
        _zz_4454_ = int_reg_array_10_62_imag;
        _zz_4455_ = int_reg_array_10_62_real;
      end
      default : begin
        _zz_4454_ = int_reg_array_10_63_imag;
        _zz_4455_ = int_reg_array_10_63_real;
      end
    endcase
  end

  always @(*) begin
    case(_zz_776_)
      6'b000000 : begin
        _zz_4456_ = int_reg_array_11_0_imag;
        _zz_4457_ = int_reg_array_11_0_real;
      end
      6'b000001 : begin
        _zz_4456_ = int_reg_array_11_1_imag;
        _zz_4457_ = int_reg_array_11_1_real;
      end
      6'b000010 : begin
        _zz_4456_ = int_reg_array_11_2_imag;
        _zz_4457_ = int_reg_array_11_2_real;
      end
      6'b000011 : begin
        _zz_4456_ = int_reg_array_11_3_imag;
        _zz_4457_ = int_reg_array_11_3_real;
      end
      6'b000100 : begin
        _zz_4456_ = int_reg_array_11_4_imag;
        _zz_4457_ = int_reg_array_11_4_real;
      end
      6'b000101 : begin
        _zz_4456_ = int_reg_array_11_5_imag;
        _zz_4457_ = int_reg_array_11_5_real;
      end
      6'b000110 : begin
        _zz_4456_ = int_reg_array_11_6_imag;
        _zz_4457_ = int_reg_array_11_6_real;
      end
      6'b000111 : begin
        _zz_4456_ = int_reg_array_11_7_imag;
        _zz_4457_ = int_reg_array_11_7_real;
      end
      6'b001000 : begin
        _zz_4456_ = int_reg_array_11_8_imag;
        _zz_4457_ = int_reg_array_11_8_real;
      end
      6'b001001 : begin
        _zz_4456_ = int_reg_array_11_9_imag;
        _zz_4457_ = int_reg_array_11_9_real;
      end
      6'b001010 : begin
        _zz_4456_ = int_reg_array_11_10_imag;
        _zz_4457_ = int_reg_array_11_10_real;
      end
      6'b001011 : begin
        _zz_4456_ = int_reg_array_11_11_imag;
        _zz_4457_ = int_reg_array_11_11_real;
      end
      6'b001100 : begin
        _zz_4456_ = int_reg_array_11_12_imag;
        _zz_4457_ = int_reg_array_11_12_real;
      end
      6'b001101 : begin
        _zz_4456_ = int_reg_array_11_13_imag;
        _zz_4457_ = int_reg_array_11_13_real;
      end
      6'b001110 : begin
        _zz_4456_ = int_reg_array_11_14_imag;
        _zz_4457_ = int_reg_array_11_14_real;
      end
      6'b001111 : begin
        _zz_4456_ = int_reg_array_11_15_imag;
        _zz_4457_ = int_reg_array_11_15_real;
      end
      6'b010000 : begin
        _zz_4456_ = int_reg_array_11_16_imag;
        _zz_4457_ = int_reg_array_11_16_real;
      end
      6'b010001 : begin
        _zz_4456_ = int_reg_array_11_17_imag;
        _zz_4457_ = int_reg_array_11_17_real;
      end
      6'b010010 : begin
        _zz_4456_ = int_reg_array_11_18_imag;
        _zz_4457_ = int_reg_array_11_18_real;
      end
      6'b010011 : begin
        _zz_4456_ = int_reg_array_11_19_imag;
        _zz_4457_ = int_reg_array_11_19_real;
      end
      6'b010100 : begin
        _zz_4456_ = int_reg_array_11_20_imag;
        _zz_4457_ = int_reg_array_11_20_real;
      end
      6'b010101 : begin
        _zz_4456_ = int_reg_array_11_21_imag;
        _zz_4457_ = int_reg_array_11_21_real;
      end
      6'b010110 : begin
        _zz_4456_ = int_reg_array_11_22_imag;
        _zz_4457_ = int_reg_array_11_22_real;
      end
      6'b010111 : begin
        _zz_4456_ = int_reg_array_11_23_imag;
        _zz_4457_ = int_reg_array_11_23_real;
      end
      6'b011000 : begin
        _zz_4456_ = int_reg_array_11_24_imag;
        _zz_4457_ = int_reg_array_11_24_real;
      end
      6'b011001 : begin
        _zz_4456_ = int_reg_array_11_25_imag;
        _zz_4457_ = int_reg_array_11_25_real;
      end
      6'b011010 : begin
        _zz_4456_ = int_reg_array_11_26_imag;
        _zz_4457_ = int_reg_array_11_26_real;
      end
      6'b011011 : begin
        _zz_4456_ = int_reg_array_11_27_imag;
        _zz_4457_ = int_reg_array_11_27_real;
      end
      6'b011100 : begin
        _zz_4456_ = int_reg_array_11_28_imag;
        _zz_4457_ = int_reg_array_11_28_real;
      end
      6'b011101 : begin
        _zz_4456_ = int_reg_array_11_29_imag;
        _zz_4457_ = int_reg_array_11_29_real;
      end
      6'b011110 : begin
        _zz_4456_ = int_reg_array_11_30_imag;
        _zz_4457_ = int_reg_array_11_30_real;
      end
      6'b011111 : begin
        _zz_4456_ = int_reg_array_11_31_imag;
        _zz_4457_ = int_reg_array_11_31_real;
      end
      6'b100000 : begin
        _zz_4456_ = int_reg_array_11_32_imag;
        _zz_4457_ = int_reg_array_11_32_real;
      end
      6'b100001 : begin
        _zz_4456_ = int_reg_array_11_33_imag;
        _zz_4457_ = int_reg_array_11_33_real;
      end
      6'b100010 : begin
        _zz_4456_ = int_reg_array_11_34_imag;
        _zz_4457_ = int_reg_array_11_34_real;
      end
      6'b100011 : begin
        _zz_4456_ = int_reg_array_11_35_imag;
        _zz_4457_ = int_reg_array_11_35_real;
      end
      6'b100100 : begin
        _zz_4456_ = int_reg_array_11_36_imag;
        _zz_4457_ = int_reg_array_11_36_real;
      end
      6'b100101 : begin
        _zz_4456_ = int_reg_array_11_37_imag;
        _zz_4457_ = int_reg_array_11_37_real;
      end
      6'b100110 : begin
        _zz_4456_ = int_reg_array_11_38_imag;
        _zz_4457_ = int_reg_array_11_38_real;
      end
      6'b100111 : begin
        _zz_4456_ = int_reg_array_11_39_imag;
        _zz_4457_ = int_reg_array_11_39_real;
      end
      6'b101000 : begin
        _zz_4456_ = int_reg_array_11_40_imag;
        _zz_4457_ = int_reg_array_11_40_real;
      end
      6'b101001 : begin
        _zz_4456_ = int_reg_array_11_41_imag;
        _zz_4457_ = int_reg_array_11_41_real;
      end
      6'b101010 : begin
        _zz_4456_ = int_reg_array_11_42_imag;
        _zz_4457_ = int_reg_array_11_42_real;
      end
      6'b101011 : begin
        _zz_4456_ = int_reg_array_11_43_imag;
        _zz_4457_ = int_reg_array_11_43_real;
      end
      6'b101100 : begin
        _zz_4456_ = int_reg_array_11_44_imag;
        _zz_4457_ = int_reg_array_11_44_real;
      end
      6'b101101 : begin
        _zz_4456_ = int_reg_array_11_45_imag;
        _zz_4457_ = int_reg_array_11_45_real;
      end
      6'b101110 : begin
        _zz_4456_ = int_reg_array_11_46_imag;
        _zz_4457_ = int_reg_array_11_46_real;
      end
      6'b101111 : begin
        _zz_4456_ = int_reg_array_11_47_imag;
        _zz_4457_ = int_reg_array_11_47_real;
      end
      6'b110000 : begin
        _zz_4456_ = int_reg_array_11_48_imag;
        _zz_4457_ = int_reg_array_11_48_real;
      end
      6'b110001 : begin
        _zz_4456_ = int_reg_array_11_49_imag;
        _zz_4457_ = int_reg_array_11_49_real;
      end
      6'b110010 : begin
        _zz_4456_ = int_reg_array_11_50_imag;
        _zz_4457_ = int_reg_array_11_50_real;
      end
      6'b110011 : begin
        _zz_4456_ = int_reg_array_11_51_imag;
        _zz_4457_ = int_reg_array_11_51_real;
      end
      6'b110100 : begin
        _zz_4456_ = int_reg_array_11_52_imag;
        _zz_4457_ = int_reg_array_11_52_real;
      end
      6'b110101 : begin
        _zz_4456_ = int_reg_array_11_53_imag;
        _zz_4457_ = int_reg_array_11_53_real;
      end
      6'b110110 : begin
        _zz_4456_ = int_reg_array_11_54_imag;
        _zz_4457_ = int_reg_array_11_54_real;
      end
      6'b110111 : begin
        _zz_4456_ = int_reg_array_11_55_imag;
        _zz_4457_ = int_reg_array_11_55_real;
      end
      6'b111000 : begin
        _zz_4456_ = int_reg_array_11_56_imag;
        _zz_4457_ = int_reg_array_11_56_real;
      end
      6'b111001 : begin
        _zz_4456_ = int_reg_array_11_57_imag;
        _zz_4457_ = int_reg_array_11_57_real;
      end
      6'b111010 : begin
        _zz_4456_ = int_reg_array_11_58_imag;
        _zz_4457_ = int_reg_array_11_58_real;
      end
      6'b111011 : begin
        _zz_4456_ = int_reg_array_11_59_imag;
        _zz_4457_ = int_reg_array_11_59_real;
      end
      6'b111100 : begin
        _zz_4456_ = int_reg_array_11_60_imag;
        _zz_4457_ = int_reg_array_11_60_real;
      end
      6'b111101 : begin
        _zz_4456_ = int_reg_array_11_61_imag;
        _zz_4457_ = int_reg_array_11_61_real;
      end
      6'b111110 : begin
        _zz_4456_ = int_reg_array_11_62_imag;
        _zz_4457_ = int_reg_array_11_62_real;
      end
      default : begin
        _zz_4456_ = int_reg_array_11_63_imag;
        _zz_4457_ = int_reg_array_11_63_real;
      end
    endcase
  end

  always @(*) begin
    case(_zz_845_)
      6'b000000 : begin
        _zz_4458_ = int_reg_array_12_0_imag;
        _zz_4459_ = int_reg_array_12_0_real;
      end
      6'b000001 : begin
        _zz_4458_ = int_reg_array_12_1_imag;
        _zz_4459_ = int_reg_array_12_1_real;
      end
      6'b000010 : begin
        _zz_4458_ = int_reg_array_12_2_imag;
        _zz_4459_ = int_reg_array_12_2_real;
      end
      6'b000011 : begin
        _zz_4458_ = int_reg_array_12_3_imag;
        _zz_4459_ = int_reg_array_12_3_real;
      end
      6'b000100 : begin
        _zz_4458_ = int_reg_array_12_4_imag;
        _zz_4459_ = int_reg_array_12_4_real;
      end
      6'b000101 : begin
        _zz_4458_ = int_reg_array_12_5_imag;
        _zz_4459_ = int_reg_array_12_5_real;
      end
      6'b000110 : begin
        _zz_4458_ = int_reg_array_12_6_imag;
        _zz_4459_ = int_reg_array_12_6_real;
      end
      6'b000111 : begin
        _zz_4458_ = int_reg_array_12_7_imag;
        _zz_4459_ = int_reg_array_12_7_real;
      end
      6'b001000 : begin
        _zz_4458_ = int_reg_array_12_8_imag;
        _zz_4459_ = int_reg_array_12_8_real;
      end
      6'b001001 : begin
        _zz_4458_ = int_reg_array_12_9_imag;
        _zz_4459_ = int_reg_array_12_9_real;
      end
      6'b001010 : begin
        _zz_4458_ = int_reg_array_12_10_imag;
        _zz_4459_ = int_reg_array_12_10_real;
      end
      6'b001011 : begin
        _zz_4458_ = int_reg_array_12_11_imag;
        _zz_4459_ = int_reg_array_12_11_real;
      end
      6'b001100 : begin
        _zz_4458_ = int_reg_array_12_12_imag;
        _zz_4459_ = int_reg_array_12_12_real;
      end
      6'b001101 : begin
        _zz_4458_ = int_reg_array_12_13_imag;
        _zz_4459_ = int_reg_array_12_13_real;
      end
      6'b001110 : begin
        _zz_4458_ = int_reg_array_12_14_imag;
        _zz_4459_ = int_reg_array_12_14_real;
      end
      6'b001111 : begin
        _zz_4458_ = int_reg_array_12_15_imag;
        _zz_4459_ = int_reg_array_12_15_real;
      end
      6'b010000 : begin
        _zz_4458_ = int_reg_array_12_16_imag;
        _zz_4459_ = int_reg_array_12_16_real;
      end
      6'b010001 : begin
        _zz_4458_ = int_reg_array_12_17_imag;
        _zz_4459_ = int_reg_array_12_17_real;
      end
      6'b010010 : begin
        _zz_4458_ = int_reg_array_12_18_imag;
        _zz_4459_ = int_reg_array_12_18_real;
      end
      6'b010011 : begin
        _zz_4458_ = int_reg_array_12_19_imag;
        _zz_4459_ = int_reg_array_12_19_real;
      end
      6'b010100 : begin
        _zz_4458_ = int_reg_array_12_20_imag;
        _zz_4459_ = int_reg_array_12_20_real;
      end
      6'b010101 : begin
        _zz_4458_ = int_reg_array_12_21_imag;
        _zz_4459_ = int_reg_array_12_21_real;
      end
      6'b010110 : begin
        _zz_4458_ = int_reg_array_12_22_imag;
        _zz_4459_ = int_reg_array_12_22_real;
      end
      6'b010111 : begin
        _zz_4458_ = int_reg_array_12_23_imag;
        _zz_4459_ = int_reg_array_12_23_real;
      end
      6'b011000 : begin
        _zz_4458_ = int_reg_array_12_24_imag;
        _zz_4459_ = int_reg_array_12_24_real;
      end
      6'b011001 : begin
        _zz_4458_ = int_reg_array_12_25_imag;
        _zz_4459_ = int_reg_array_12_25_real;
      end
      6'b011010 : begin
        _zz_4458_ = int_reg_array_12_26_imag;
        _zz_4459_ = int_reg_array_12_26_real;
      end
      6'b011011 : begin
        _zz_4458_ = int_reg_array_12_27_imag;
        _zz_4459_ = int_reg_array_12_27_real;
      end
      6'b011100 : begin
        _zz_4458_ = int_reg_array_12_28_imag;
        _zz_4459_ = int_reg_array_12_28_real;
      end
      6'b011101 : begin
        _zz_4458_ = int_reg_array_12_29_imag;
        _zz_4459_ = int_reg_array_12_29_real;
      end
      6'b011110 : begin
        _zz_4458_ = int_reg_array_12_30_imag;
        _zz_4459_ = int_reg_array_12_30_real;
      end
      6'b011111 : begin
        _zz_4458_ = int_reg_array_12_31_imag;
        _zz_4459_ = int_reg_array_12_31_real;
      end
      6'b100000 : begin
        _zz_4458_ = int_reg_array_12_32_imag;
        _zz_4459_ = int_reg_array_12_32_real;
      end
      6'b100001 : begin
        _zz_4458_ = int_reg_array_12_33_imag;
        _zz_4459_ = int_reg_array_12_33_real;
      end
      6'b100010 : begin
        _zz_4458_ = int_reg_array_12_34_imag;
        _zz_4459_ = int_reg_array_12_34_real;
      end
      6'b100011 : begin
        _zz_4458_ = int_reg_array_12_35_imag;
        _zz_4459_ = int_reg_array_12_35_real;
      end
      6'b100100 : begin
        _zz_4458_ = int_reg_array_12_36_imag;
        _zz_4459_ = int_reg_array_12_36_real;
      end
      6'b100101 : begin
        _zz_4458_ = int_reg_array_12_37_imag;
        _zz_4459_ = int_reg_array_12_37_real;
      end
      6'b100110 : begin
        _zz_4458_ = int_reg_array_12_38_imag;
        _zz_4459_ = int_reg_array_12_38_real;
      end
      6'b100111 : begin
        _zz_4458_ = int_reg_array_12_39_imag;
        _zz_4459_ = int_reg_array_12_39_real;
      end
      6'b101000 : begin
        _zz_4458_ = int_reg_array_12_40_imag;
        _zz_4459_ = int_reg_array_12_40_real;
      end
      6'b101001 : begin
        _zz_4458_ = int_reg_array_12_41_imag;
        _zz_4459_ = int_reg_array_12_41_real;
      end
      6'b101010 : begin
        _zz_4458_ = int_reg_array_12_42_imag;
        _zz_4459_ = int_reg_array_12_42_real;
      end
      6'b101011 : begin
        _zz_4458_ = int_reg_array_12_43_imag;
        _zz_4459_ = int_reg_array_12_43_real;
      end
      6'b101100 : begin
        _zz_4458_ = int_reg_array_12_44_imag;
        _zz_4459_ = int_reg_array_12_44_real;
      end
      6'b101101 : begin
        _zz_4458_ = int_reg_array_12_45_imag;
        _zz_4459_ = int_reg_array_12_45_real;
      end
      6'b101110 : begin
        _zz_4458_ = int_reg_array_12_46_imag;
        _zz_4459_ = int_reg_array_12_46_real;
      end
      6'b101111 : begin
        _zz_4458_ = int_reg_array_12_47_imag;
        _zz_4459_ = int_reg_array_12_47_real;
      end
      6'b110000 : begin
        _zz_4458_ = int_reg_array_12_48_imag;
        _zz_4459_ = int_reg_array_12_48_real;
      end
      6'b110001 : begin
        _zz_4458_ = int_reg_array_12_49_imag;
        _zz_4459_ = int_reg_array_12_49_real;
      end
      6'b110010 : begin
        _zz_4458_ = int_reg_array_12_50_imag;
        _zz_4459_ = int_reg_array_12_50_real;
      end
      6'b110011 : begin
        _zz_4458_ = int_reg_array_12_51_imag;
        _zz_4459_ = int_reg_array_12_51_real;
      end
      6'b110100 : begin
        _zz_4458_ = int_reg_array_12_52_imag;
        _zz_4459_ = int_reg_array_12_52_real;
      end
      6'b110101 : begin
        _zz_4458_ = int_reg_array_12_53_imag;
        _zz_4459_ = int_reg_array_12_53_real;
      end
      6'b110110 : begin
        _zz_4458_ = int_reg_array_12_54_imag;
        _zz_4459_ = int_reg_array_12_54_real;
      end
      6'b110111 : begin
        _zz_4458_ = int_reg_array_12_55_imag;
        _zz_4459_ = int_reg_array_12_55_real;
      end
      6'b111000 : begin
        _zz_4458_ = int_reg_array_12_56_imag;
        _zz_4459_ = int_reg_array_12_56_real;
      end
      6'b111001 : begin
        _zz_4458_ = int_reg_array_12_57_imag;
        _zz_4459_ = int_reg_array_12_57_real;
      end
      6'b111010 : begin
        _zz_4458_ = int_reg_array_12_58_imag;
        _zz_4459_ = int_reg_array_12_58_real;
      end
      6'b111011 : begin
        _zz_4458_ = int_reg_array_12_59_imag;
        _zz_4459_ = int_reg_array_12_59_real;
      end
      6'b111100 : begin
        _zz_4458_ = int_reg_array_12_60_imag;
        _zz_4459_ = int_reg_array_12_60_real;
      end
      6'b111101 : begin
        _zz_4458_ = int_reg_array_12_61_imag;
        _zz_4459_ = int_reg_array_12_61_real;
      end
      6'b111110 : begin
        _zz_4458_ = int_reg_array_12_62_imag;
        _zz_4459_ = int_reg_array_12_62_real;
      end
      default : begin
        _zz_4458_ = int_reg_array_12_63_imag;
        _zz_4459_ = int_reg_array_12_63_real;
      end
    endcase
  end

  always @(*) begin
    case(_zz_914_)
      6'b000000 : begin
        _zz_4460_ = int_reg_array_13_0_imag;
        _zz_4461_ = int_reg_array_13_0_real;
      end
      6'b000001 : begin
        _zz_4460_ = int_reg_array_13_1_imag;
        _zz_4461_ = int_reg_array_13_1_real;
      end
      6'b000010 : begin
        _zz_4460_ = int_reg_array_13_2_imag;
        _zz_4461_ = int_reg_array_13_2_real;
      end
      6'b000011 : begin
        _zz_4460_ = int_reg_array_13_3_imag;
        _zz_4461_ = int_reg_array_13_3_real;
      end
      6'b000100 : begin
        _zz_4460_ = int_reg_array_13_4_imag;
        _zz_4461_ = int_reg_array_13_4_real;
      end
      6'b000101 : begin
        _zz_4460_ = int_reg_array_13_5_imag;
        _zz_4461_ = int_reg_array_13_5_real;
      end
      6'b000110 : begin
        _zz_4460_ = int_reg_array_13_6_imag;
        _zz_4461_ = int_reg_array_13_6_real;
      end
      6'b000111 : begin
        _zz_4460_ = int_reg_array_13_7_imag;
        _zz_4461_ = int_reg_array_13_7_real;
      end
      6'b001000 : begin
        _zz_4460_ = int_reg_array_13_8_imag;
        _zz_4461_ = int_reg_array_13_8_real;
      end
      6'b001001 : begin
        _zz_4460_ = int_reg_array_13_9_imag;
        _zz_4461_ = int_reg_array_13_9_real;
      end
      6'b001010 : begin
        _zz_4460_ = int_reg_array_13_10_imag;
        _zz_4461_ = int_reg_array_13_10_real;
      end
      6'b001011 : begin
        _zz_4460_ = int_reg_array_13_11_imag;
        _zz_4461_ = int_reg_array_13_11_real;
      end
      6'b001100 : begin
        _zz_4460_ = int_reg_array_13_12_imag;
        _zz_4461_ = int_reg_array_13_12_real;
      end
      6'b001101 : begin
        _zz_4460_ = int_reg_array_13_13_imag;
        _zz_4461_ = int_reg_array_13_13_real;
      end
      6'b001110 : begin
        _zz_4460_ = int_reg_array_13_14_imag;
        _zz_4461_ = int_reg_array_13_14_real;
      end
      6'b001111 : begin
        _zz_4460_ = int_reg_array_13_15_imag;
        _zz_4461_ = int_reg_array_13_15_real;
      end
      6'b010000 : begin
        _zz_4460_ = int_reg_array_13_16_imag;
        _zz_4461_ = int_reg_array_13_16_real;
      end
      6'b010001 : begin
        _zz_4460_ = int_reg_array_13_17_imag;
        _zz_4461_ = int_reg_array_13_17_real;
      end
      6'b010010 : begin
        _zz_4460_ = int_reg_array_13_18_imag;
        _zz_4461_ = int_reg_array_13_18_real;
      end
      6'b010011 : begin
        _zz_4460_ = int_reg_array_13_19_imag;
        _zz_4461_ = int_reg_array_13_19_real;
      end
      6'b010100 : begin
        _zz_4460_ = int_reg_array_13_20_imag;
        _zz_4461_ = int_reg_array_13_20_real;
      end
      6'b010101 : begin
        _zz_4460_ = int_reg_array_13_21_imag;
        _zz_4461_ = int_reg_array_13_21_real;
      end
      6'b010110 : begin
        _zz_4460_ = int_reg_array_13_22_imag;
        _zz_4461_ = int_reg_array_13_22_real;
      end
      6'b010111 : begin
        _zz_4460_ = int_reg_array_13_23_imag;
        _zz_4461_ = int_reg_array_13_23_real;
      end
      6'b011000 : begin
        _zz_4460_ = int_reg_array_13_24_imag;
        _zz_4461_ = int_reg_array_13_24_real;
      end
      6'b011001 : begin
        _zz_4460_ = int_reg_array_13_25_imag;
        _zz_4461_ = int_reg_array_13_25_real;
      end
      6'b011010 : begin
        _zz_4460_ = int_reg_array_13_26_imag;
        _zz_4461_ = int_reg_array_13_26_real;
      end
      6'b011011 : begin
        _zz_4460_ = int_reg_array_13_27_imag;
        _zz_4461_ = int_reg_array_13_27_real;
      end
      6'b011100 : begin
        _zz_4460_ = int_reg_array_13_28_imag;
        _zz_4461_ = int_reg_array_13_28_real;
      end
      6'b011101 : begin
        _zz_4460_ = int_reg_array_13_29_imag;
        _zz_4461_ = int_reg_array_13_29_real;
      end
      6'b011110 : begin
        _zz_4460_ = int_reg_array_13_30_imag;
        _zz_4461_ = int_reg_array_13_30_real;
      end
      6'b011111 : begin
        _zz_4460_ = int_reg_array_13_31_imag;
        _zz_4461_ = int_reg_array_13_31_real;
      end
      6'b100000 : begin
        _zz_4460_ = int_reg_array_13_32_imag;
        _zz_4461_ = int_reg_array_13_32_real;
      end
      6'b100001 : begin
        _zz_4460_ = int_reg_array_13_33_imag;
        _zz_4461_ = int_reg_array_13_33_real;
      end
      6'b100010 : begin
        _zz_4460_ = int_reg_array_13_34_imag;
        _zz_4461_ = int_reg_array_13_34_real;
      end
      6'b100011 : begin
        _zz_4460_ = int_reg_array_13_35_imag;
        _zz_4461_ = int_reg_array_13_35_real;
      end
      6'b100100 : begin
        _zz_4460_ = int_reg_array_13_36_imag;
        _zz_4461_ = int_reg_array_13_36_real;
      end
      6'b100101 : begin
        _zz_4460_ = int_reg_array_13_37_imag;
        _zz_4461_ = int_reg_array_13_37_real;
      end
      6'b100110 : begin
        _zz_4460_ = int_reg_array_13_38_imag;
        _zz_4461_ = int_reg_array_13_38_real;
      end
      6'b100111 : begin
        _zz_4460_ = int_reg_array_13_39_imag;
        _zz_4461_ = int_reg_array_13_39_real;
      end
      6'b101000 : begin
        _zz_4460_ = int_reg_array_13_40_imag;
        _zz_4461_ = int_reg_array_13_40_real;
      end
      6'b101001 : begin
        _zz_4460_ = int_reg_array_13_41_imag;
        _zz_4461_ = int_reg_array_13_41_real;
      end
      6'b101010 : begin
        _zz_4460_ = int_reg_array_13_42_imag;
        _zz_4461_ = int_reg_array_13_42_real;
      end
      6'b101011 : begin
        _zz_4460_ = int_reg_array_13_43_imag;
        _zz_4461_ = int_reg_array_13_43_real;
      end
      6'b101100 : begin
        _zz_4460_ = int_reg_array_13_44_imag;
        _zz_4461_ = int_reg_array_13_44_real;
      end
      6'b101101 : begin
        _zz_4460_ = int_reg_array_13_45_imag;
        _zz_4461_ = int_reg_array_13_45_real;
      end
      6'b101110 : begin
        _zz_4460_ = int_reg_array_13_46_imag;
        _zz_4461_ = int_reg_array_13_46_real;
      end
      6'b101111 : begin
        _zz_4460_ = int_reg_array_13_47_imag;
        _zz_4461_ = int_reg_array_13_47_real;
      end
      6'b110000 : begin
        _zz_4460_ = int_reg_array_13_48_imag;
        _zz_4461_ = int_reg_array_13_48_real;
      end
      6'b110001 : begin
        _zz_4460_ = int_reg_array_13_49_imag;
        _zz_4461_ = int_reg_array_13_49_real;
      end
      6'b110010 : begin
        _zz_4460_ = int_reg_array_13_50_imag;
        _zz_4461_ = int_reg_array_13_50_real;
      end
      6'b110011 : begin
        _zz_4460_ = int_reg_array_13_51_imag;
        _zz_4461_ = int_reg_array_13_51_real;
      end
      6'b110100 : begin
        _zz_4460_ = int_reg_array_13_52_imag;
        _zz_4461_ = int_reg_array_13_52_real;
      end
      6'b110101 : begin
        _zz_4460_ = int_reg_array_13_53_imag;
        _zz_4461_ = int_reg_array_13_53_real;
      end
      6'b110110 : begin
        _zz_4460_ = int_reg_array_13_54_imag;
        _zz_4461_ = int_reg_array_13_54_real;
      end
      6'b110111 : begin
        _zz_4460_ = int_reg_array_13_55_imag;
        _zz_4461_ = int_reg_array_13_55_real;
      end
      6'b111000 : begin
        _zz_4460_ = int_reg_array_13_56_imag;
        _zz_4461_ = int_reg_array_13_56_real;
      end
      6'b111001 : begin
        _zz_4460_ = int_reg_array_13_57_imag;
        _zz_4461_ = int_reg_array_13_57_real;
      end
      6'b111010 : begin
        _zz_4460_ = int_reg_array_13_58_imag;
        _zz_4461_ = int_reg_array_13_58_real;
      end
      6'b111011 : begin
        _zz_4460_ = int_reg_array_13_59_imag;
        _zz_4461_ = int_reg_array_13_59_real;
      end
      6'b111100 : begin
        _zz_4460_ = int_reg_array_13_60_imag;
        _zz_4461_ = int_reg_array_13_60_real;
      end
      6'b111101 : begin
        _zz_4460_ = int_reg_array_13_61_imag;
        _zz_4461_ = int_reg_array_13_61_real;
      end
      6'b111110 : begin
        _zz_4460_ = int_reg_array_13_62_imag;
        _zz_4461_ = int_reg_array_13_62_real;
      end
      default : begin
        _zz_4460_ = int_reg_array_13_63_imag;
        _zz_4461_ = int_reg_array_13_63_real;
      end
    endcase
  end

  always @(*) begin
    case(_zz_983_)
      6'b000000 : begin
        _zz_4462_ = int_reg_array_14_0_imag;
        _zz_4463_ = int_reg_array_14_0_real;
      end
      6'b000001 : begin
        _zz_4462_ = int_reg_array_14_1_imag;
        _zz_4463_ = int_reg_array_14_1_real;
      end
      6'b000010 : begin
        _zz_4462_ = int_reg_array_14_2_imag;
        _zz_4463_ = int_reg_array_14_2_real;
      end
      6'b000011 : begin
        _zz_4462_ = int_reg_array_14_3_imag;
        _zz_4463_ = int_reg_array_14_3_real;
      end
      6'b000100 : begin
        _zz_4462_ = int_reg_array_14_4_imag;
        _zz_4463_ = int_reg_array_14_4_real;
      end
      6'b000101 : begin
        _zz_4462_ = int_reg_array_14_5_imag;
        _zz_4463_ = int_reg_array_14_5_real;
      end
      6'b000110 : begin
        _zz_4462_ = int_reg_array_14_6_imag;
        _zz_4463_ = int_reg_array_14_6_real;
      end
      6'b000111 : begin
        _zz_4462_ = int_reg_array_14_7_imag;
        _zz_4463_ = int_reg_array_14_7_real;
      end
      6'b001000 : begin
        _zz_4462_ = int_reg_array_14_8_imag;
        _zz_4463_ = int_reg_array_14_8_real;
      end
      6'b001001 : begin
        _zz_4462_ = int_reg_array_14_9_imag;
        _zz_4463_ = int_reg_array_14_9_real;
      end
      6'b001010 : begin
        _zz_4462_ = int_reg_array_14_10_imag;
        _zz_4463_ = int_reg_array_14_10_real;
      end
      6'b001011 : begin
        _zz_4462_ = int_reg_array_14_11_imag;
        _zz_4463_ = int_reg_array_14_11_real;
      end
      6'b001100 : begin
        _zz_4462_ = int_reg_array_14_12_imag;
        _zz_4463_ = int_reg_array_14_12_real;
      end
      6'b001101 : begin
        _zz_4462_ = int_reg_array_14_13_imag;
        _zz_4463_ = int_reg_array_14_13_real;
      end
      6'b001110 : begin
        _zz_4462_ = int_reg_array_14_14_imag;
        _zz_4463_ = int_reg_array_14_14_real;
      end
      6'b001111 : begin
        _zz_4462_ = int_reg_array_14_15_imag;
        _zz_4463_ = int_reg_array_14_15_real;
      end
      6'b010000 : begin
        _zz_4462_ = int_reg_array_14_16_imag;
        _zz_4463_ = int_reg_array_14_16_real;
      end
      6'b010001 : begin
        _zz_4462_ = int_reg_array_14_17_imag;
        _zz_4463_ = int_reg_array_14_17_real;
      end
      6'b010010 : begin
        _zz_4462_ = int_reg_array_14_18_imag;
        _zz_4463_ = int_reg_array_14_18_real;
      end
      6'b010011 : begin
        _zz_4462_ = int_reg_array_14_19_imag;
        _zz_4463_ = int_reg_array_14_19_real;
      end
      6'b010100 : begin
        _zz_4462_ = int_reg_array_14_20_imag;
        _zz_4463_ = int_reg_array_14_20_real;
      end
      6'b010101 : begin
        _zz_4462_ = int_reg_array_14_21_imag;
        _zz_4463_ = int_reg_array_14_21_real;
      end
      6'b010110 : begin
        _zz_4462_ = int_reg_array_14_22_imag;
        _zz_4463_ = int_reg_array_14_22_real;
      end
      6'b010111 : begin
        _zz_4462_ = int_reg_array_14_23_imag;
        _zz_4463_ = int_reg_array_14_23_real;
      end
      6'b011000 : begin
        _zz_4462_ = int_reg_array_14_24_imag;
        _zz_4463_ = int_reg_array_14_24_real;
      end
      6'b011001 : begin
        _zz_4462_ = int_reg_array_14_25_imag;
        _zz_4463_ = int_reg_array_14_25_real;
      end
      6'b011010 : begin
        _zz_4462_ = int_reg_array_14_26_imag;
        _zz_4463_ = int_reg_array_14_26_real;
      end
      6'b011011 : begin
        _zz_4462_ = int_reg_array_14_27_imag;
        _zz_4463_ = int_reg_array_14_27_real;
      end
      6'b011100 : begin
        _zz_4462_ = int_reg_array_14_28_imag;
        _zz_4463_ = int_reg_array_14_28_real;
      end
      6'b011101 : begin
        _zz_4462_ = int_reg_array_14_29_imag;
        _zz_4463_ = int_reg_array_14_29_real;
      end
      6'b011110 : begin
        _zz_4462_ = int_reg_array_14_30_imag;
        _zz_4463_ = int_reg_array_14_30_real;
      end
      6'b011111 : begin
        _zz_4462_ = int_reg_array_14_31_imag;
        _zz_4463_ = int_reg_array_14_31_real;
      end
      6'b100000 : begin
        _zz_4462_ = int_reg_array_14_32_imag;
        _zz_4463_ = int_reg_array_14_32_real;
      end
      6'b100001 : begin
        _zz_4462_ = int_reg_array_14_33_imag;
        _zz_4463_ = int_reg_array_14_33_real;
      end
      6'b100010 : begin
        _zz_4462_ = int_reg_array_14_34_imag;
        _zz_4463_ = int_reg_array_14_34_real;
      end
      6'b100011 : begin
        _zz_4462_ = int_reg_array_14_35_imag;
        _zz_4463_ = int_reg_array_14_35_real;
      end
      6'b100100 : begin
        _zz_4462_ = int_reg_array_14_36_imag;
        _zz_4463_ = int_reg_array_14_36_real;
      end
      6'b100101 : begin
        _zz_4462_ = int_reg_array_14_37_imag;
        _zz_4463_ = int_reg_array_14_37_real;
      end
      6'b100110 : begin
        _zz_4462_ = int_reg_array_14_38_imag;
        _zz_4463_ = int_reg_array_14_38_real;
      end
      6'b100111 : begin
        _zz_4462_ = int_reg_array_14_39_imag;
        _zz_4463_ = int_reg_array_14_39_real;
      end
      6'b101000 : begin
        _zz_4462_ = int_reg_array_14_40_imag;
        _zz_4463_ = int_reg_array_14_40_real;
      end
      6'b101001 : begin
        _zz_4462_ = int_reg_array_14_41_imag;
        _zz_4463_ = int_reg_array_14_41_real;
      end
      6'b101010 : begin
        _zz_4462_ = int_reg_array_14_42_imag;
        _zz_4463_ = int_reg_array_14_42_real;
      end
      6'b101011 : begin
        _zz_4462_ = int_reg_array_14_43_imag;
        _zz_4463_ = int_reg_array_14_43_real;
      end
      6'b101100 : begin
        _zz_4462_ = int_reg_array_14_44_imag;
        _zz_4463_ = int_reg_array_14_44_real;
      end
      6'b101101 : begin
        _zz_4462_ = int_reg_array_14_45_imag;
        _zz_4463_ = int_reg_array_14_45_real;
      end
      6'b101110 : begin
        _zz_4462_ = int_reg_array_14_46_imag;
        _zz_4463_ = int_reg_array_14_46_real;
      end
      6'b101111 : begin
        _zz_4462_ = int_reg_array_14_47_imag;
        _zz_4463_ = int_reg_array_14_47_real;
      end
      6'b110000 : begin
        _zz_4462_ = int_reg_array_14_48_imag;
        _zz_4463_ = int_reg_array_14_48_real;
      end
      6'b110001 : begin
        _zz_4462_ = int_reg_array_14_49_imag;
        _zz_4463_ = int_reg_array_14_49_real;
      end
      6'b110010 : begin
        _zz_4462_ = int_reg_array_14_50_imag;
        _zz_4463_ = int_reg_array_14_50_real;
      end
      6'b110011 : begin
        _zz_4462_ = int_reg_array_14_51_imag;
        _zz_4463_ = int_reg_array_14_51_real;
      end
      6'b110100 : begin
        _zz_4462_ = int_reg_array_14_52_imag;
        _zz_4463_ = int_reg_array_14_52_real;
      end
      6'b110101 : begin
        _zz_4462_ = int_reg_array_14_53_imag;
        _zz_4463_ = int_reg_array_14_53_real;
      end
      6'b110110 : begin
        _zz_4462_ = int_reg_array_14_54_imag;
        _zz_4463_ = int_reg_array_14_54_real;
      end
      6'b110111 : begin
        _zz_4462_ = int_reg_array_14_55_imag;
        _zz_4463_ = int_reg_array_14_55_real;
      end
      6'b111000 : begin
        _zz_4462_ = int_reg_array_14_56_imag;
        _zz_4463_ = int_reg_array_14_56_real;
      end
      6'b111001 : begin
        _zz_4462_ = int_reg_array_14_57_imag;
        _zz_4463_ = int_reg_array_14_57_real;
      end
      6'b111010 : begin
        _zz_4462_ = int_reg_array_14_58_imag;
        _zz_4463_ = int_reg_array_14_58_real;
      end
      6'b111011 : begin
        _zz_4462_ = int_reg_array_14_59_imag;
        _zz_4463_ = int_reg_array_14_59_real;
      end
      6'b111100 : begin
        _zz_4462_ = int_reg_array_14_60_imag;
        _zz_4463_ = int_reg_array_14_60_real;
      end
      6'b111101 : begin
        _zz_4462_ = int_reg_array_14_61_imag;
        _zz_4463_ = int_reg_array_14_61_real;
      end
      6'b111110 : begin
        _zz_4462_ = int_reg_array_14_62_imag;
        _zz_4463_ = int_reg_array_14_62_real;
      end
      default : begin
        _zz_4462_ = int_reg_array_14_63_imag;
        _zz_4463_ = int_reg_array_14_63_real;
      end
    endcase
  end

  always @(*) begin
    case(_zz_1052_)
      6'b000000 : begin
        _zz_4464_ = int_reg_array_15_0_imag;
        _zz_4465_ = int_reg_array_15_0_real;
      end
      6'b000001 : begin
        _zz_4464_ = int_reg_array_15_1_imag;
        _zz_4465_ = int_reg_array_15_1_real;
      end
      6'b000010 : begin
        _zz_4464_ = int_reg_array_15_2_imag;
        _zz_4465_ = int_reg_array_15_2_real;
      end
      6'b000011 : begin
        _zz_4464_ = int_reg_array_15_3_imag;
        _zz_4465_ = int_reg_array_15_3_real;
      end
      6'b000100 : begin
        _zz_4464_ = int_reg_array_15_4_imag;
        _zz_4465_ = int_reg_array_15_4_real;
      end
      6'b000101 : begin
        _zz_4464_ = int_reg_array_15_5_imag;
        _zz_4465_ = int_reg_array_15_5_real;
      end
      6'b000110 : begin
        _zz_4464_ = int_reg_array_15_6_imag;
        _zz_4465_ = int_reg_array_15_6_real;
      end
      6'b000111 : begin
        _zz_4464_ = int_reg_array_15_7_imag;
        _zz_4465_ = int_reg_array_15_7_real;
      end
      6'b001000 : begin
        _zz_4464_ = int_reg_array_15_8_imag;
        _zz_4465_ = int_reg_array_15_8_real;
      end
      6'b001001 : begin
        _zz_4464_ = int_reg_array_15_9_imag;
        _zz_4465_ = int_reg_array_15_9_real;
      end
      6'b001010 : begin
        _zz_4464_ = int_reg_array_15_10_imag;
        _zz_4465_ = int_reg_array_15_10_real;
      end
      6'b001011 : begin
        _zz_4464_ = int_reg_array_15_11_imag;
        _zz_4465_ = int_reg_array_15_11_real;
      end
      6'b001100 : begin
        _zz_4464_ = int_reg_array_15_12_imag;
        _zz_4465_ = int_reg_array_15_12_real;
      end
      6'b001101 : begin
        _zz_4464_ = int_reg_array_15_13_imag;
        _zz_4465_ = int_reg_array_15_13_real;
      end
      6'b001110 : begin
        _zz_4464_ = int_reg_array_15_14_imag;
        _zz_4465_ = int_reg_array_15_14_real;
      end
      6'b001111 : begin
        _zz_4464_ = int_reg_array_15_15_imag;
        _zz_4465_ = int_reg_array_15_15_real;
      end
      6'b010000 : begin
        _zz_4464_ = int_reg_array_15_16_imag;
        _zz_4465_ = int_reg_array_15_16_real;
      end
      6'b010001 : begin
        _zz_4464_ = int_reg_array_15_17_imag;
        _zz_4465_ = int_reg_array_15_17_real;
      end
      6'b010010 : begin
        _zz_4464_ = int_reg_array_15_18_imag;
        _zz_4465_ = int_reg_array_15_18_real;
      end
      6'b010011 : begin
        _zz_4464_ = int_reg_array_15_19_imag;
        _zz_4465_ = int_reg_array_15_19_real;
      end
      6'b010100 : begin
        _zz_4464_ = int_reg_array_15_20_imag;
        _zz_4465_ = int_reg_array_15_20_real;
      end
      6'b010101 : begin
        _zz_4464_ = int_reg_array_15_21_imag;
        _zz_4465_ = int_reg_array_15_21_real;
      end
      6'b010110 : begin
        _zz_4464_ = int_reg_array_15_22_imag;
        _zz_4465_ = int_reg_array_15_22_real;
      end
      6'b010111 : begin
        _zz_4464_ = int_reg_array_15_23_imag;
        _zz_4465_ = int_reg_array_15_23_real;
      end
      6'b011000 : begin
        _zz_4464_ = int_reg_array_15_24_imag;
        _zz_4465_ = int_reg_array_15_24_real;
      end
      6'b011001 : begin
        _zz_4464_ = int_reg_array_15_25_imag;
        _zz_4465_ = int_reg_array_15_25_real;
      end
      6'b011010 : begin
        _zz_4464_ = int_reg_array_15_26_imag;
        _zz_4465_ = int_reg_array_15_26_real;
      end
      6'b011011 : begin
        _zz_4464_ = int_reg_array_15_27_imag;
        _zz_4465_ = int_reg_array_15_27_real;
      end
      6'b011100 : begin
        _zz_4464_ = int_reg_array_15_28_imag;
        _zz_4465_ = int_reg_array_15_28_real;
      end
      6'b011101 : begin
        _zz_4464_ = int_reg_array_15_29_imag;
        _zz_4465_ = int_reg_array_15_29_real;
      end
      6'b011110 : begin
        _zz_4464_ = int_reg_array_15_30_imag;
        _zz_4465_ = int_reg_array_15_30_real;
      end
      6'b011111 : begin
        _zz_4464_ = int_reg_array_15_31_imag;
        _zz_4465_ = int_reg_array_15_31_real;
      end
      6'b100000 : begin
        _zz_4464_ = int_reg_array_15_32_imag;
        _zz_4465_ = int_reg_array_15_32_real;
      end
      6'b100001 : begin
        _zz_4464_ = int_reg_array_15_33_imag;
        _zz_4465_ = int_reg_array_15_33_real;
      end
      6'b100010 : begin
        _zz_4464_ = int_reg_array_15_34_imag;
        _zz_4465_ = int_reg_array_15_34_real;
      end
      6'b100011 : begin
        _zz_4464_ = int_reg_array_15_35_imag;
        _zz_4465_ = int_reg_array_15_35_real;
      end
      6'b100100 : begin
        _zz_4464_ = int_reg_array_15_36_imag;
        _zz_4465_ = int_reg_array_15_36_real;
      end
      6'b100101 : begin
        _zz_4464_ = int_reg_array_15_37_imag;
        _zz_4465_ = int_reg_array_15_37_real;
      end
      6'b100110 : begin
        _zz_4464_ = int_reg_array_15_38_imag;
        _zz_4465_ = int_reg_array_15_38_real;
      end
      6'b100111 : begin
        _zz_4464_ = int_reg_array_15_39_imag;
        _zz_4465_ = int_reg_array_15_39_real;
      end
      6'b101000 : begin
        _zz_4464_ = int_reg_array_15_40_imag;
        _zz_4465_ = int_reg_array_15_40_real;
      end
      6'b101001 : begin
        _zz_4464_ = int_reg_array_15_41_imag;
        _zz_4465_ = int_reg_array_15_41_real;
      end
      6'b101010 : begin
        _zz_4464_ = int_reg_array_15_42_imag;
        _zz_4465_ = int_reg_array_15_42_real;
      end
      6'b101011 : begin
        _zz_4464_ = int_reg_array_15_43_imag;
        _zz_4465_ = int_reg_array_15_43_real;
      end
      6'b101100 : begin
        _zz_4464_ = int_reg_array_15_44_imag;
        _zz_4465_ = int_reg_array_15_44_real;
      end
      6'b101101 : begin
        _zz_4464_ = int_reg_array_15_45_imag;
        _zz_4465_ = int_reg_array_15_45_real;
      end
      6'b101110 : begin
        _zz_4464_ = int_reg_array_15_46_imag;
        _zz_4465_ = int_reg_array_15_46_real;
      end
      6'b101111 : begin
        _zz_4464_ = int_reg_array_15_47_imag;
        _zz_4465_ = int_reg_array_15_47_real;
      end
      6'b110000 : begin
        _zz_4464_ = int_reg_array_15_48_imag;
        _zz_4465_ = int_reg_array_15_48_real;
      end
      6'b110001 : begin
        _zz_4464_ = int_reg_array_15_49_imag;
        _zz_4465_ = int_reg_array_15_49_real;
      end
      6'b110010 : begin
        _zz_4464_ = int_reg_array_15_50_imag;
        _zz_4465_ = int_reg_array_15_50_real;
      end
      6'b110011 : begin
        _zz_4464_ = int_reg_array_15_51_imag;
        _zz_4465_ = int_reg_array_15_51_real;
      end
      6'b110100 : begin
        _zz_4464_ = int_reg_array_15_52_imag;
        _zz_4465_ = int_reg_array_15_52_real;
      end
      6'b110101 : begin
        _zz_4464_ = int_reg_array_15_53_imag;
        _zz_4465_ = int_reg_array_15_53_real;
      end
      6'b110110 : begin
        _zz_4464_ = int_reg_array_15_54_imag;
        _zz_4465_ = int_reg_array_15_54_real;
      end
      6'b110111 : begin
        _zz_4464_ = int_reg_array_15_55_imag;
        _zz_4465_ = int_reg_array_15_55_real;
      end
      6'b111000 : begin
        _zz_4464_ = int_reg_array_15_56_imag;
        _zz_4465_ = int_reg_array_15_56_real;
      end
      6'b111001 : begin
        _zz_4464_ = int_reg_array_15_57_imag;
        _zz_4465_ = int_reg_array_15_57_real;
      end
      6'b111010 : begin
        _zz_4464_ = int_reg_array_15_58_imag;
        _zz_4465_ = int_reg_array_15_58_real;
      end
      6'b111011 : begin
        _zz_4464_ = int_reg_array_15_59_imag;
        _zz_4465_ = int_reg_array_15_59_real;
      end
      6'b111100 : begin
        _zz_4464_ = int_reg_array_15_60_imag;
        _zz_4465_ = int_reg_array_15_60_real;
      end
      6'b111101 : begin
        _zz_4464_ = int_reg_array_15_61_imag;
        _zz_4465_ = int_reg_array_15_61_real;
      end
      6'b111110 : begin
        _zz_4464_ = int_reg_array_15_62_imag;
        _zz_4465_ = int_reg_array_15_62_real;
      end
      default : begin
        _zz_4464_ = int_reg_array_15_63_imag;
        _zz_4465_ = int_reg_array_15_63_real;
      end
    endcase
  end

  always @(*) begin
    case(_zz_1121_)
      6'b000000 : begin
        _zz_4466_ = int_reg_array_16_0_imag;
        _zz_4467_ = int_reg_array_16_0_real;
      end
      6'b000001 : begin
        _zz_4466_ = int_reg_array_16_1_imag;
        _zz_4467_ = int_reg_array_16_1_real;
      end
      6'b000010 : begin
        _zz_4466_ = int_reg_array_16_2_imag;
        _zz_4467_ = int_reg_array_16_2_real;
      end
      6'b000011 : begin
        _zz_4466_ = int_reg_array_16_3_imag;
        _zz_4467_ = int_reg_array_16_3_real;
      end
      6'b000100 : begin
        _zz_4466_ = int_reg_array_16_4_imag;
        _zz_4467_ = int_reg_array_16_4_real;
      end
      6'b000101 : begin
        _zz_4466_ = int_reg_array_16_5_imag;
        _zz_4467_ = int_reg_array_16_5_real;
      end
      6'b000110 : begin
        _zz_4466_ = int_reg_array_16_6_imag;
        _zz_4467_ = int_reg_array_16_6_real;
      end
      6'b000111 : begin
        _zz_4466_ = int_reg_array_16_7_imag;
        _zz_4467_ = int_reg_array_16_7_real;
      end
      6'b001000 : begin
        _zz_4466_ = int_reg_array_16_8_imag;
        _zz_4467_ = int_reg_array_16_8_real;
      end
      6'b001001 : begin
        _zz_4466_ = int_reg_array_16_9_imag;
        _zz_4467_ = int_reg_array_16_9_real;
      end
      6'b001010 : begin
        _zz_4466_ = int_reg_array_16_10_imag;
        _zz_4467_ = int_reg_array_16_10_real;
      end
      6'b001011 : begin
        _zz_4466_ = int_reg_array_16_11_imag;
        _zz_4467_ = int_reg_array_16_11_real;
      end
      6'b001100 : begin
        _zz_4466_ = int_reg_array_16_12_imag;
        _zz_4467_ = int_reg_array_16_12_real;
      end
      6'b001101 : begin
        _zz_4466_ = int_reg_array_16_13_imag;
        _zz_4467_ = int_reg_array_16_13_real;
      end
      6'b001110 : begin
        _zz_4466_ = int_reg_array_16_14_imag;
        _zz_4467_ = int_reg_array_16_14_real;
      end
      6'b001111 : begin
        _zz_4466_ = int_reg_array_16_15_imag;
        _zz_4467_ = int_reg_array_16_15_real;
      end
      6'b010000 : begin
        _zz_4466_ = int_reg_array_16_16_imag;
        _zz_4467_ = int_reg_array_16_16_real;
      end
      6'b010001 : begin
        _zz_4466_ = int_reg_array_16_17_imag;
        _zz_4467_ = int_reg_array_16_17_real;
      end
      6'b010010 : begin
        _zz_4466_ = int_reg_array_16_18_imag;
        _zz_4467_ = int_reg_array_16_18_real;
      end
      6'b010011 : begin
        _zz_4466_ = int_reg_array_16_19_imag;
        _zz_4467_ = int_reg_array_16_19_real;
      end
      6'b010100 : begin
        _zz_4466_ = int_reg_array_16_20_imag;
        _zz_4467_ = int_reg_array_16_20_real;
      end
      6'b010101 : begin
        _zz_4466_ = int_reg_array_16_21_imag;
        _zz_4467_ = int_reg_array_16_21_real;
      end
      6'b010110 : begin
        _zz_4466_ = int_reg_array_16_22_imag;
        _zz_4467_ = int_reg_array_16_22_real;
      end
      6'b010111 : begin
        _zz_4466_ = int_reg_array_16_23_imag;
        _zz_4467_ = int_reg_array_16_23_real;
      end
      6'b011000 : begin
        _zz_4466_ = int_reg_array_16_24_imag;
        _zz_4467_ = int_reg_array_16_24_real;
      end
      6'b011001 : begin
        _zz_4466_ = int_reg_array_16_25_imag;
        _zz_4467_ = int_reg_array_16_25_real;
      end
      6'b011010 : begin
        _zz_4466_ = int_reg_array_16_26_imag;
        _zz_4467_ = int_reg_array_16_26_real;
      end
      6'b011011 : begin
        _zz_4466_ = int_reg_array_16_27_imag;
        _zz_4467_ = int_reg_array_16_27_real;
      end
      6'b011100 : begin
        _zz_4466_ = int_reg_array_16_28_imag;
        _zz_4467_ = int_reg_array_16_28_real;
      end
      6'b011101 : begin
        _zz_4466_ = int_reg_array_16_29_imag;
        _zz_4467_ = int_reg_array_16_29_real;
      end
      6'b011110 : begin
        _zz_4466_ = int_reg_array_16_30_imag;
        _zz_4467_ = int_reg_array_16_30_real;
      end
      6'b011111 : begin
        _zz_4466_ = int_reg_array_16_31_imag;
        _zz_4467_ = int_reg_array_16_31_real;
      end
      6'b100000 : begin
        _zz_4466_ = int_reg_array_16_32_imag;
        _zz_4467_ = int_reg_array_16_32_real;
      end
      6'b100001 : begin
        _zz_4466_ = int_reg_array_16_33_imag;
        _zz_4467_ = int_reg_array_16_33_real;
      end
      6'b100010 : begin
        _zz_4466_ = int_reg_array_16_34_imag;
        _zz_4467_ = int_reg_array_16_34_real;
      end
      6'b100011 : begin
        _zz_4466_ = int_reg_array_16_35_imag;
        _zz_4467_ = int_reg_array_16_35_real;
      end
      6'b100100 : begin
        _zz_4466_ = int_reg_array_16_36_imag;
        _zz_4467_ = int_reg_array_16_36_real;
      end
      6'b100101 : begin
        _zz_4466_ = int_reg_array_16_37_imag;
        _zz_4467_ = int_reg_array_16_37_real;
      end
      6'b100110 : begin
        _zz_4466_ = int_reg_array_16_38_imag;
        _zz_4467_ = int_reg_array_16_38_real;
      end
      6'b100111 : begin
        _zz_4466_ = int_reg_array_16_39_imag;
        _zz_4467_ = int_reg_array_16_39_real;
      end
      6'b101000 : begin
        _zz_4466_ = int_reg_array_16_40_imag;
        _zz_4467_ = int_reg_array_16_40_real;
      end
      6'b101001 : begin
        _zz_4466_ = int_reg_array_16_41_imag;
        _zz_4467_ = int_reg_array_16_41_real;
      end
      6'b101010 : begin
        _zz_4466_ = int_reg_array_16_42_imag;
        _zz_4467_ = int_reg_array_16_42_real;
      end
      6'b101011 : begin
        _zz_4466_ = int_reg_array_16_43_imag;
        _zz_4467_ = int_reg_array_16_43_real;
      end
      6'b101100 : begin
        _zz_4466_ = int_reg_array_16_44_imag;
        _zz_4467_ = int_reg_array_16_44_real;
      end
      6'b101101 : begin
        _zz_4466_ = int_reg_array_16_45_imag;
        _zz_4467_ = int_reg_array_16_45_real;
      end
      6'b101110 : begin
        _zz_4466_ = int_reg_array_16_46_imag;
        _zz_4467_ = int_reg_array_16_46_real;
      end
      6'b101111 : begin
        _zz_4466_ = int_reg_array_16_47_imag;
        _zz_4467_ = int_reg_array_16_47_real;
      end
      6'b110000 : begin
        _zz_4466_ = int_reg_array_16_48_imag;
        _zz_4467_ = int_reg_array_16_48_real;
      end
      6'b110001 : begin
        _zz_4466_ = int_reg_array_16_49_imag;
        _zz_4467_ = int_reg_array_16_49_real;
      end
      6'b110010 : begin
        _zz_4466_ = int_reg_array_16_50_imag;
        _zz_4467_ = int_reg_array_16_50_real;
      end
      6'b110011 : begin
        _zz_4466_ = int_reg_array_16_51_imag;
        _zz_4467_ = int_reg_array_16_51_real;
      end
      6'b110100 : begin
        _zz_4466_ = int_reg_array_16_52_imag;
        _zz_4467_ = int_reg_array_16_52_real;
      end
      6'b110101 : begin
        _zz_4466_ = int_reg_array_16_53_imag;
        _zz_4467_ = int_reg_array_16_53_real;
      end
      6'b110110 : begin
        _zz_4466_ = int_reg_array_16_54_imag;
        _zz_4467_ = int_reg_array_16_54_real;
      end
      6'b110111 : begin
        _zz_4466_ = int_reg_array_16_55_imag;
        _zz_4467_ = int_reg_array_16_55_real;
      end
      6'b111000 : begin
        _zz_4466_ = int_reg_array_16_56_imag;
        _zz_4467_ = int_reg_array_16_56_real;
      end
      6'b111001 : begin
        _zz_4466_ = int_reg_array_16_57_imag;
        _zz_4467_ = int_reg_array_16_57_real;
      end
      6'b111010 : begin
        _zz_4466_ = int_reg_array_16_58_imag;
        _zz_4467_ = int_reg_array_16_58_real;
      end
      6'b111011 : begin
        _zz_4466_ = int_reg_array_16_59_imag;
        _zz_4467_ = int_reg_array_16_59_real;
      end
      6'b111100 : begin
        _zz_4466_ = int_reg_array_16_60_imag;
        _zz_4467_ = int_reg_array_16_60_real;
      end
      6'b111101 : begin
        _zz_4466_ = int_reg_array_16_61_imag;
        _zz_4467_ = int_reg_array_16_61_real;
      end
      6'b111110 : begin
        _zz_4466_ = int_reg_array_16_62_imag;
        _zz_4467_ = int_reg_array_16_62_real;
      end
      default : begin
        _zz_4466_ = int_reg_array_16_63_imag;
        _zz_4467_ = int_reg_array_16_63_real;
      end
    endcase
  end

  always @(*) begin
    case(_zz_1190_)
      6'b000000 : begin
        _zz_4468_ = int_reg_array_17_0_imag;
        _zz_4469_ = int_reg_array_17_0_real;
      end
      6'b000001 : begin
        _zz_4468_ = int_reg_array_17_1_imag;
        _zz_4469_ = int_reg_array_17_1_real;
      end
      6'b000010 : begin
        _zz_4468_ = int_reg_array_17_2_imag;
        _zz_4469_ = int_reg_array_17_2_real;
      end
      6'b000011 : begin
        _zz_4468_ = int_reg_array_17_3_imag;
        _zz_4469_ = int_reg_array_17_3_real;
      end
      6'b000100 : begin
        _zz_4468_ = int_reg_array_17_4_imag;
        _zz_4469_ = int_reg_array_17_4_real;
      end
      6'b000101 : begin
        _zz_4468_ = int_reg_array_17_5_imag;
        _zz_4469_ = int_reg_array_17_5_real;
      end
      6'b000110 : begin
        _zz_4468_ = int_reg_array_17_6_imag;
        _zz_4469_ = int_reg_array_17_6_real;
      end
      6'b000111 : begin
        _zz_4468_ = int_reg_array_17_7_imag;
        _zz_4469_ = int_reg_array_17_7_real;
      end
      6'b001000 : begin
        _zz_4468_ = int_reg_array_17_8_imag;
        _zz_4469_ = int_reg_array_17_8_real;
      end
      6'b001001 : begin
        _zz_4468_ = int_reg_array_17_9_imag;
        _zz_4469_ = int_reg_array_17_9_real;
      end
      6'b001010 : begin
        _zz_4468_ = int_reg_array_17_10_imag;
        _zz_4469_ = int_reg_array_17_10_real;
      end
      6'b001011 : begin
        _zz_4468_ = int_reg_array_17_11_imag;
        _zz_4469_ = int_reg_array_17_11_real;
      end
      6'b001100 : begin
        _zz_4468_ = int_reg_array_17_12_imag;
        _zz_4469_ = int_reg_array_17_12_real;
      end
      6'b001101 : begin
        _zz_4468_ = int_reg_array_17_13_imag;
        _zz_4469_ = int_reg_array_17_13_real;
      end
      6'b001110 : begin
        _zz_4468_ = int_reg_array_17_14_imag;
        _zz_4469_ = int_reg_array_17_14_real;
      end
      6'b001111 : begin
        _zz_4468_ = int_reg_array_17_15_imag;
        _zz_4469_ = int_reg_array_17_15_real;
      end
      6'b010000 : begin
        _zz_4468_ = int_reg_array_17_16_imag;
        _zz_4469_ = int_reg_array_17_16_real;
      end
      6'b010001 : begin
        _zz_4468_ = int_reg_array_17_17_imag;
        _zz_4469_ = int_reg_array_17_17_real;
      end
      6'b010010 : begin
        _zz_4468_ = int_reg_array_17_18_imag;
        _zz_4469_ = int_reg_array_17_18_real;
      end
      6'b010011 : begin
        _zz_4468_ = int_reg_array_17_19_imag;
        _zz_4469_ = int_reg_array_17_19_real;
      end
      6'b010100 : begin
        _zz_4468_ = int_reg_array_17_20_imag;
        _zz_4469_ = int_reg_array_17_20_real;
      end
      6'b010101 : begin
        _zz_4468_ = int_reg_array_17_21_imag;
        _zz_4469_ = int_reg_array_17_21_real;
      end
      6'b010110 : begin
        _zz_4468_ = int_reg_array_17_22_imag;
        _zz_4469_ = int_reg_array_17_22_real;
      end
      6'b010111 : begin
        _zz_4468_ = int_reg_array_17_23_imag;
        _zz_4469_ = int_reg_array_17_23_real;
      end
      6'b011000 : begin
        _zz_4468_ = int_reg_array_17_24_imag;
        _zz_4469_ = int_reg_array_17_24_real;
      end
      6'b011001 : begin
        _zz_4468_ = int_reg_array_17_25_imag;
        _zz_4469_ = int_reg_array_17_25_real;
      end
      6'b011010 : begin
        _zz_4468_ = int_reg_array_17_26_imag;
        _zz_4469_ = int_reg_array_17_26_real;
      end
      6'b011011 : begin
        _zz_4468_ = int_reg_array_17_27_imag;
        _zz_4469_ = int_reg_array_17_27_real;
      end
      6'b011100 : begin
        _zz_4468_ = int_reg_array_17_28_imag;
        _zz_4469_ = int_reg_array_17_28_real;
      end
      6'b011101 : begin
        _zz_4468_ = int_reg_array_17_29_imag;
        _zz_4469_ = int_reg_array_17_29_real;
      end
      6'b011110 : begin
        _zz_4468_ = int_reg_array_17_30_imag;
        _zz_4469_ = int_reg_array_17_30_real;
      end
      6'b011111 : begin
        _zz_4468_ = int_reg_array_17_31_imag;
        _zz_4469_ = int_reg_array_17_31_real;
      end
      6'b100000 : begin
        _zz_4468_ = int_reg_array_17_32_imag;
        _zz_4469_ = int_reg_array_17_32_real;
      end
      6'b100001 : begin
        _zz_4468_ = int_reg_array_17_33_imag;
        _zz_4469_ = int_reg_array_17_33_real;
      end
      6'b100010 : begin
        _zz_4468_ = int_reg_array_17_34_imag;
        _zz_4469_ = int_reg_array_17_34_real;
      end
      6'b100011 : begin
        _zz_4468_ = int_reg_array_17_35_imag;
        _zz_4469_ = int_reg_array_17_35_real;
      end
      6'b100100 : begin
        _zz_4468_ = int_reg_array_17_36_imag;
        _zz_4469_ = int_reg_array_17_36_real;
      end
      6'b100101 : begin
        _zz_4468_ = int_reg_array_17_37_imag;
        _zz_4469_ = int_reg_array_17_37_real;
      end
      6'b100110 : begin
        _zz_4468_ = int_reg_array_17_38_imag;
        _zz_4469_ = int_reg_array_17_38_real;
      end
      6'b100111 : begin
        _zz_4468_ = int_reg_array_17_39_imag;
        _zz_4469_ = int_reg_array_17_39_real;
      end
      6'b101000 : begin
        _zz_4468_ = int_reg_array_17_40_imag;
        _zz_4469_ = int_reg_array_17_40_real;
      end
      6'b101001 : begin
        _zz_4468_ = int_reg_array_17_41_imag;
        _zz_4469_ = int_reg_array_17_41_real;
      end
      6'b101010 : begin
        _zz_4468_ = int_reg_array_17_42_imag;
        _zz_4469_ = int_reg_array_17_42_real;
      end
      6'b101011 : begin
        _zz_4468_ = int_reg_array_17_43_imag;
        _zz_4469_ = int_reg_array_17_43_real;
      end
      6'b101100 : begin
        _zz_4468_ = int_reg_array_17_44_imag;
        _zz_4469_ = int_reg_array_17_44_real;
      end
      6'b101101 : begin
        _zz_4468_ = int_reg_array_17_45_imag;
        _zz_4469_ = int_reg_array_17_45_real;
      end
      6'b101110 : begin
        _zz_4468_ = int_reg_array_17_46_imag;
        _zz_4469_ = int_reg_array_17_46_real;
      end
      6'b101111 : begin
        _zz_4468_ = int_reg_array_17_47_imag;
        _zz_4469_ = int_reg_array_17_47_real;
      end
      6'b110000 : begin
        _zz_4468_ = int_reg_array_17_48_imag;
        _zz_4469_ = int_reg_array_17_48_real;
      end
      6'b110001 : begin
        _zz_4468_ = int_reg_array_17_49_imag;
        _zz_4469_ = int_reg_array_17_49_real;
      end
      6'b110010 : begin
        _zz_4468_ = int_reg_array_17_50_imag;
        _zz_4469_ = int_reg_array_17_50_real;
      end
      6'b110011 : begin
        _zz_4468_ = int_reg_array_17_51_imag;
        _zz_4469_ = int_reg_array_17_51_real;
      end
      6'b110100 : begin
        _zz_4468_ = int_reg_array_17_52_imag;
        _zz_4469_ = int_reg_array_17_52_real;
      end
      6'b110101 : begin
        _zz_4468_ = int_reg_array_17_53_imag;
        _zz_4469_ = int_reg_array_17_53_real;
      end
      6'b110110 : begin
        _zz_4468_ = int_reg_array_17_54_imag;
        _zz_4469_ = int_reg_array_17_54_real;
      end
      6'b110111 : begin
        _zz_4468_ = int_reg_array_17_55_imag;
        _zz_4469_ = int_reg_array_17_55_real;
      end
      6'b111000 : begin
        _zz_4468_ = int_reg_array_17_56_imag;
        _zz_4469_ = int_reg_array_17_56_real;
      end
      6'b111001 : begin
        _zz_4468_ = int_reg_array_17_57_imag;
        _zz_4469_ = int_reg_array_17_57_real;
      end
      6'b111010 : begin
        _zz_4468_ = int_reg_array_17_58_imag;
        _zz_4469_ = int_reg_array_17_58_real;
      end
      6'b111011 : begin
        _zz_4468_ = int_reg_array_17_59_imag;
        _zz_4469_ = int_reg_array_17_59_real;
      end
      6'b111100 : begin
        _zz_4468_ = int_reg_array_17_60_imag;
        _zz_4469_ = int_reg_array_17_60_real;
      end
      6'b111101 : begin
        _zz_4468_ = int_reg_array_17_61_imag;
        _zz_4469_ = int_reg_array_17_61_real;
      end
      6'b111110 : begin
        _zz_4468_ = int_reg_array_17_62_imag;
        _zz_4469_ = int_reg_array_17_62_real;
      end
      default : begin
        _zz_4468_ = int_reg_array_17_63_imag;
        _zz_4469_ = int_reg_array_17_63_real;
      end
    endcase
  end

  always @(*) begin
    case(_zz_1259_)
      6'b000000 : begin
        _zz_4470_ = int_reg_array_18_0_imag;
        _zz_4471_ = int_reg_array_18_0_real;
      end
      6'b000001 : begin
        _zz_4470_ = int_reg_array_18_1_imag;
        _zz_4471_ = int_reg_array_18_1_real;
      end
      6'b000010 : begin
        _zz_4470_ = int_reg_array_18_2_imag;
        _zz_4471_ = int_reg_array_18_2_real;
      end
      6'b000011 : begin
        _zz_4470_ = int_reg_array_18_3_imag;
        _zz_4471_ = int_reg_array_18_3_real;
      end
      6'b000100 : begin
        _zz_4470_ = int_reg_array_18_4_imag;
        _zz_4471_ = int_reg_array_18_4_real;
      end
      6'b000101 : begin
        _zz_4470_ = int_reg_array_18_5_imag;
        _zz_4471_ = int_reg_array_18_5_real;
      end
      6'b000110 : begin
        _zz_4470_ = int_reg_array_18_6_imag;
        _zz_4471_ = int_reg_array_18_6_real;
      end
      6'b000111 : begin
        _zz_4470_ = int_reg_array_18_7_imag;
        _zz_4471_ = int_reg_array_18_7_real;
      end
      6'b001000 : begin
        _zz_4470_ = int_reg_array_18_8_imag;
        _zz_4471_ = int_reg_array_18_8_real;
      end
      6'b001001 : begin
        _zz_4470_ = int_reg_array_18_9_imag;
        _zz_4471_ = int_reg_array_18_9_real;
      end
      6'b001010 : begin
        _zz_4470_ = int_reg_array_18_10_imag;
        _zz_4471_ = int_reg_array_18_10_real;
      end
      6'b001011 : begin
        _zz_4470_ = int_reg_array_18_11_imag;
        _zz_4471_ = int_reg_array_18_11_real;
      end
      6'b001100 : begin
        _zz_4470_ = int_reg_array_18_12_imag;
        _zz_4471_ = int_reg_array_18_12_real;
      end
      6'b001101 : begin
        _zz_4470_ = int_reg_array_18_13_imag;
        _zz_4471_ = int_reg_array_18_13_real;
      end
      6'b001110 : begin
        _zz_4470_ = int_reg_array_18_14_imag;
        _zz_4471_ = int_reg_array_18_14_real;
      end
      6'b001111 : begin
        _zz_4470_ = int_reg_array_18_15_imag;
        _zz_4471_ = int_reg_array_18_15_real;
      end
      6'b010000 : begin
        _zz_4470_ = int_reg_array_18_16_imag;
        _zz_4471_ = int_reg_array_18_16_real;
      end
      6'b010001 : begin
        _zz_4470_ = int_reg_array_18_17_imag;
        _zz_4471_ = int_reg_array_18_17_real;
      end
      6'b010010 : begin
        _zz_4470_ = int_reg_array_18_18_imag;
        _zz_4471_ = int_reg_array_18_18_real;
      end
      6'b010011 : begin
        _zz_4470_ = int_reg_array_18_19_imag;
        _zz_4471_ = int_reg_array_18_19_real;
      end
      6'b010100 : begin
        _zz_4470_ = int_reg_array_18_20_imag;
        _zz_4471_ = int_reg_array_18_20_real;
      end
      6'b010101 : begin
        _zz_4470_ = int_reg_array_18_21_imag;
        _zz_4471_ = int_reg_array_18_21_real;
      end
      6'b010110 : begin
        _zz_4470_ = int_reg_array_18_22_imag;
        _zz_4471_ = int_reg_array_18_22_real;
      end
      6'b010111 : begin
        _zz_4470_ = int_reg_array_18_23_imag;
        _zz_4471_ = int_reg_array_18_23_real;
      end
      6'b011000 : begin
        _zz_4470_ = int_reg_array_18_24_imag;
        _zz_4471_ = int_reg_array_18_24_real;
      end
      6'b011001 : begin
        _zz_4470_ = int_reg_array_18_25_imag;
        _zz_4471_ = int_reg_array_18_25_real;
      end
      6'b011010 : begin
        _zz_4470_ = int_reg_array_18_26_imag;
        _zz_4471_ = int_reg_array_18_26_real;
      end
      6'b011011 : begin
        _zz_4470_ = int_reg_array_18_27_imag;
        _zz_4471_ = int_reg_array_18_27_real;
      end
      6'b011100 : begin
        _zz_4470_ = int_reg_array_18_28_imag;
        _zz_4471_ = int_reg_array_18_28_real;
      end
      6'b011101 : begin
        _zz_4470_ = int_reg_array_18_29_imag;
        _zz_4471_ = int_reg_array_18_29_real;
      end
      6'b011110 : begin
        _zz_4470_ = int_reg_array_18_30_imag;
        _zz_4471_ = int_reg_array_18_30_real;
      end
      6'b011111 : begin
        _zz_4470_ = int_reg_array_18_31_imag;
        _zz_4471_ = int_reg_array_18_31_real;
      end
      6'b100000 : begin
        _zz_4470_ = int_reg_array_18_32_imag;
        _zz_4471_ = int_reg_array_18_32_real;
      end
      6'b100001 : begin
        _zz_4470_ = int_reg_array_18_33_imag;
        _zz_4471_ = int_reg_array_18_33_real;
      end
      6'b100010 : begin
        _zz_4470_ = int_reg_array_18_34_imag;
        _zz_4471_ = int_reg_array_18_34_real;
      end
      6'b100011 : begin
        _zz_4470_ = int_reg_array_18_35_imag;
        _zz_4471_ = int_reg_array_18_35_real;
      end
      6'b100100 : begin
        _zz_4470_ = int_reg_array_18_36_imag;
        _zz_4471_ = int_reg_array_18_36_real;
      end
      6'b100101 : begin
        _zz_4470_ = int_reg_array_18_37_imag;
        _zz_4471_ = int_reg_array_18_37_real;
      end
      6'b100110 : begin
        _zz_4470_ = int_reg_array_18_38_imag;
        _zz_4471_ = int_reg_array_18_38_real;
      end
      6'b100111 : begin
        _zz_4470_ = int_reg_array_18_39_imag;
        _zz_4471_ = int_reg_array_18_39_real;
      end
      6'b101000 : begin
        _zz_4470_ = int_reg_array_18_40_imag;
        _zz_4471_ = int_reg_array_18_40_real;
      end
      6'b101001 : begin
        _zz_4470_ = int_reg_array_18_41_imag;
        _zz_4471_ = int_reg_array_18_41_real;
      end
      6'b101010 : begin
        _zz_4470_ = int_reg_array_18_42_imag;
        _zz_4471_ = int_reg_array_18_42_real;
      end
      6'b101011 : begin
        _zz_4470_ = int_reg_array_18_43_imag;
        _zz_4471_ = int_reg_array_18_43_real;
      end
      6'b101100 : begin
        _zz_4470_ = int_reg_array_18_44_imag;
        _zz_4471_ = int_reg_array_18_44_real;
      end
      6'b101101 : begin
        _zz_4470_ = int_reg_array_18_45_imag;
        _zz_4471_ = int_reg_array_18_45_real;
      end
      6'b101110 : begin
        _zz_4470_ = int_reg_array_18_46_imag;
        _zz_4471_ = int_reg_array_18_46_real;
      end
      6'b101111 : begin
        _zz_4470_ = int_reg_array_18_47_imag;
        _zz_4471_ = int_reg_array_18_47_real;
      end
      6'b110000 : begin
        _zz_4470_ = int_reg_array_18_48_imag;
        _zz_4471_ = int_reg_array_18_48_real;
      end
      6'b110001 : begin
        _zz_4470_ = int_reg_array_18_49_imag;
        _zz_4471_ = int_reg_array_18_49_real;
      end
      6'b110010 : begin
        _zz_4470_ = int_reg_array_18_50_imag;
        _zz_4471_ = int_reg_array_18_50_real;
      end
      6'b110011 : begin
        _zz_4470_ = int_reg_array_18_51_imag;
        _zz_4471_ = int_reg_array_18_51_real;
      end
      6'b110100 : begin
        _zz_4470_ = int_reg_array_18_52_imag;
        _zz_4471_ = int_reg_array_18_52_real;
      end
      6'b110101 : begin
        _zz_4470_ = int_reg_array_18_53_imag;
        _zz_4471_ = int_reg_array_18_53_real;
      end
      6'b110110 : begin
        _zz_4470_ = int_reg_array_18_54_imag;
        _zz_4471_ = int_reg_array_18_54_real;
      end
      6'b110111 : begin
        _zz_4470_ = int_reg_array_18_55_imag;
        _zz_4471_ = int_reg_array_18_55_real;
      end
      6'b111000 : begin
        _zz_4470_ = int_reg_array_18_56_imag;
        _zz_4471_ = int_reg_array_18_56_real;
      end
      6'b111001 : begin
        _zz_4470_ = int_reg_array_18_57_imag;
        _zz_4471_ = int_reg_array_18_57_real;
      end
      6'b111010 : begin
        _zz_4470_ = int_reg_array_18_58_imag;
        _zz_4471_ = int_reg_array_18_58_real;
      end
      6'b111011 : begin
        _zz_4470_ = int_reg_array_18_59_imag;
        _zz_4471_ = int_reg_array_18_59_real;
      end
      6'b111100 : begin
        _zz_4470_ = int_reg_array_18_60_imag;
        _zz_4471_ = int_reg_array_18_60_real;
      end
      6'b111101 : begin
        _zz_4470_ = int_reg_array_18_61_imag;
        _zz_4471_ = int_reg_array_18_61_real;
      end
      6'b111110 : begin
        _zz_4470_ = int_reg_array_18_62_imag;
        _zz_4471_ = int_reg_array_18_62_real;
      end
      default : begin
        _zz_4470_ = int_reg_array_18_63_imag;
        _zz_4471_ = int_reg_array_18_63_real;
      end
    endcase
  end

  always @(*) begin
    case(_zz_1328_)
      6'b000000 : begin
        _zz_4472_ = int_reg_array_19_0_imag;
        _zz_4473_ = int_reg_array_19_0_real;
      end
      6'b000001 : begin
        _zz_4472_ = int_reg_array_19_1_imag;
        _zz_4473_ = int_reg_array_19_1_real;
      end
      6'b000010 : begin
        _zz_4472_ = int_reg_array_19_2_imag;
        _zz_4473_ = int_reg_array_19_2_real;
      end
      6'b000011 : begin
        _zz_4472_ = int_reg_array_19_3_imag;
        _zz_4473_ = int_reg_array_19_3_real;
      end
      6'b000100 : begin
        _zz_4472_ = int_reg_array_19_4_imag;
        _zz_4473_ = int_reg_array_19_4_real;
      end
      6'b000101 : begin
        _zz_4472_ = int_reg_array_19_5_imag;
        _zz_4473_ = int_reg_array_19_5_real;
      end
      6'b000110 : begin
        _zz_4472_ = int_reg_array_19_6_imag;
        _zz_4473_ = int_reg_array_19_6_real;
      end
      6'b000111 : begin
        _zz_4472_ = int_reg_array_19_7_imag;
        _zz_4473_ = int_reg_array_19_7_real;
      end
      6'b001000 : begin
        _zz_4472_ = int_reg_array_19_8_imag;
        _zz_4473_ = int_reg_array_19_8_real;
      end
      6'b001001 : begin
        _zz_4472_ = int_reg_array_19_9_imag;
        _zz_4473_ = int_reg_array_19_9_real;
      end
      6'b001010 : begin
        _zz_4472_ = int_reg_array_19_10_imag;
        _zz_4473_ = int_reg_array_19_10_real;
      end
      6'b001011 : begin
        _zz_4472_ = int_reg_array_19_11_imag;
        _zz_4473_ = int_reg_array_19_11_real;
      end
      6'b001100 : begin
        _zz_4472_ = int_reg_array_19_12_imag;
        _zz_4473_ = int_reg_array_19_12_real;
      end
      6'b001101 : begin
        _zz_4472_ = int_reg_array_19_13_imag;
        _zz_4473_ = int_reg_array_19_13_real;
      end
      6'b001110 : begin
        _zz_4472_ = int_reg_array_19_14_imag;
        _zz_4473_ = int_reg_array_19_14_real;
      end
      6'b001111 : begin
        _zz_4472_ = int_reg_array_19_15_imag;
        _zz_4473_ = int_reg_array_19_15_real;
      end
      6'b010000 : begin
        _zz_4472_ = int_reg_array_19_16_imag;
        _zz_4473_ = int_reg_array_19_16_real;
      end
      6'b010001 : begin
        _zz_4472_ = int_reg_array_19_17_imag;
        _zz_4473_ = int_reg_array_19_17_real;
      end
      6'b010010 : begin
        _zz_4472_ = int_reg_array_19_18_imag;
        _zz_4473_ = int_reg_array_19_18_real;
      end
      6'b010011 : begin
        _zz_4472_ = int_reg_array_19_19_imag;
        _zz_4473_ = int_reg_array_19_19_real;
      end
      6'b010100 : begin
        _zz_4472_ = int_reg_array_19_20_imag;
        _zz_4473_ = int_reg_array_19_20_real;
      end
      6'b010101 : begin
        _zz_4472_ = int_reg_array_19_21_imag;
        _zz_4473_ = int_reg_array_19_21_real;
      end
      6'b010110 : begin
        _zz_4472_ = int_reg_array_19_22_imag;
        _zz_4473_ = int_reg_array_19_22_real;
      end
      6'b010111 : begin
        _zz_4472_ = int_reg_array_19_23_imag;
        _zz_4473_ = int_reg_array_19_23_real;
      end
      6'b011000 : begin
        _zz_4472_ = int_reg_array_19_24_imag;
        _zz_4473_ = int_reg_array_19_24_real;
      end
      6'b011001 : begin
        _zz_4472_ = int_reg_array_19_25_imag;
        _zz_4473_ = int_reg_array_19_25_real;
      end
      6'b011010 : begin
        _zz_4472_ = int_reg_array_19_26_imag;
        _zz_4473_ = int_reg_array_19_26_real;
      end
      6'b011011 : begin
        _zz_4472_ = int_reg_array_19_27_imag;
        _zz_4473_ = int_reg_array_19_27_real;
      end
      6'b011100 : begin
        _zz_4472_ = int_reg_array_19_28_imag;
        _zz_4473_ = int_reg_array_19_28_real;
      end
      6'b011101 : begin
        _zz_4472_ = int_reg_array_19_29_imag;
        _zz_4473_ = int_reg_array_19_29_real;
      end
      6'b011110 : begin
        _zz_4472_ = int_reg_array_19_30_imag;
        _zz_4473_ = int_reg_array_19_30_real;
      end
      6'b011111 : begin
        _zz_4472_ = int_reg_array_19_31_imag;
        _zz_4473_ = int_reg_array_19_31_real;
      end
      6'b100000 : begin
        _zz_4472_ = int_reg_array_19_32_imag;
        _zz_4473_ = int_reg_array_19_32_real;
      end
      6'b100001 : begin
        _zz_4472_ = int_reg_array_19_33_imag;
        _zz_4473_ = int_reg_array_19_33_real;
      end
      6'b100010 : begin
        _zz_4472_ = int_reg_array_19_34_imag;
        _zz_4473_ = int_reg_array_19_34_real;
      end
      6'b100011 : begin
        _zz_4472_ = int_reg_array_19_35_imag;
        _zz_4473_ = int_reg_array_19_35_real;
      end
      6'b100100 : begin
        _zz_4472_ = int_reg_array_19_36_imag;
        _zz_4473_ = int_reg_array_19_36_real;
      end
      6'b100101 : begin
        _zz_4472_ = int_reg_array_19_37_imag;
        _zz_4473_ = int_reg_array_19_37_real;
      end
      6'b100110 : begin
        _zz_4472_ = int_reg_array_19_38_imag;
        _zz_4473_ = int_reg_array_19_38_real;
      end
      6'b100111 : begin
        _zz_4472_ = int_reg_array_19_39_imag;
        _zz_4473_ = int_reg_array_19_39_real;
      end
      6'b101000 : begin
        _zz_4472_ = int_reg_array_19_40_imag;
        _zz_4473_ = int_reg_array_19_40_real;
      end
      6'b101001 : begin
        _zz_4472_ = int_reg_array_19_41_imag;
        _zz_4473_ = int_reg_array_19_41_real;
      end
      6'b101010 : begin
        _zz_4472_ = int_reg_array_19_42_imag;
        _zz_4473_ = int_reg_array_19_42_real;
      end
      6'b101011 : begin
        _zz_4472_ = int_reg_array_19_43_imag;
        _zz_4473_ = int_reg_array_19_43_real;
      end
      6'b101100 : begin
        _zz_4472_ = int_reg_array_19_44_imag;
        _zz_4473_ = int_reg_array_19_44_real;
      end
      6'b101101 : begin
        _zz_4472_ = int_reg_array_19_45_imag;
        _zz_4473_ = int_reg_array_19_45_real;
      end
      6'b101110 : begin
        _zz_4472_ = int_reg_array_19_46_imag;
        _zz_4473_ = int_reg_array_19_46_real;
      end
      6'b101111 : begin
        _zz_4472_ = int_reg_array_19_47_imag;
        _zz_4473_ = int_reg_array_19_47_real;
      end
      6'b110000 : begin
        _zz_4472_ = int_reg_array_19_48_imag;
        _zz_4473_ = int_reg_array_19_48_real;
      end
      6'b110001 : begin
        _zz_4472_ = int_reg_array_19_49_imag;
        _zz_4473_ = int_reg_array_19_49_real;
      end
      6'b110010 : begin
        _zz_4472_ = int_reg_array_19_50_imag;
        _zz_4473_ = int_reg_array_19_50_real;
      end
      6'b110011 : begin
        _zz_4472_ = int_reg_array_19_51_imag;
        _zz_4473_ = int_reg_array_19_51_real;
      end
      6'b110100 : begin
        _zz_4472_ = int_reg_array_19_52_imag;
        _zz_4473_ = int_reg_array_19_52_real;
      end
      6'b110101 : begin
        _zz_4472_ = int_reg_array_19_53_imag;
        _zz_4473_ = int_reg_array_19_53_real;
      end
      6'b110110 : begin
        _zz_4472_ = int_reg_array_19_54_imag;
        _zz_4473_ = int_reg_array_19_54_real;
      end
      6'b110111 : begin
        _zz_4472_ = int_reg_array_19_55_imag;
        _zz_4473_ = int_reg_array_19_55_real;
      end
      6'b111000 : begin
        _zz_4472_ = int_reg_array_19_56_imag;
        _zz_4473_ = int_reg_array_19_56_real;
      end
      6'b111001 : begin
        _zz_4472_ = int_reg_array_19_57_imag;
        _zz_4473_ = int_reg_array_19_57_real;
      end
      6'b111010 : begin
        _zz_4472_ = int_reg_array_19_58_imag;
        _zz_4473_ = int_reg_array_19_58_real;
      end
      6'b111011 : begin
        _zz_4472_ = int_reg_array_19_59_imag;
        _zz_4473_ = int_reg_array_19_59_real;
      end
      6'b111100 : begin
        _zz_4472_ = int_reg_array_19_60_imag;
        _zz_4473_ = int_reg_array_19_60_real;
      end
      6'b111101 : begin
        _zz_4472_ = int_reg_array_19_61_imag;
        _zz_4473_ = int_reg_array_19_61_real;
      end
      6'b111110 : begin
        _zz_4472_ = int_reg_array_19_62_imag;
        _zz_4473_ = int_reg_array_19_62_real;
      end
      default : begin
        _zz_4472_ = int_reg_array_19_63_imag;
        _zz_4473_ = int_reg_array_19_63_real;
      end
    endcase
  end

  always @(*) begin
    case(_zz_1397_)
      6'b000000 : begin
        _zz_4474_ = int_reg_array_20_0_imag;
        _zz_4475_ = int_reg_array_20_0_real;
      end
      6'b000001 : begin
        _zz_4474_ = int_reg_array_20_1_imag;
        _zz_4475_ = int_reg_array_20_1_real;
      end
      6'b000010 : begin
        _zz_4474_ = int_reg_array_20_2_imag;
        _zz_4475_ = int_reg_array_20_2_real;
      end
      6'b000011 : begin
        _zz_4474_ = int_reg_array_20_3_imag;
        _zz_4475_ = int_reg_array_20_3_real;
      end
      6'b000100 : begin
        _zz_4474_ = int_reg_array_20_4_imag;
        _zz_4475_ = int_reg_array_20_4_real;
      end
      6'b000101 : begin
        _zz_4474_ = int_reg_array_20_5_imag;
        _zz_4475_ = int_reg_array_20_5_real;
      end
      6'b000110 : begin
        _zz_4474_ = int_reg_array_20_6_imag;
        _zz_4475_ = int_reg_array_20_6_real;
      end
      6'b000111 : begin
        _zz_4474_ = int_reg_array_20_7_imag;
        _zz_4475_ = int_reg_array_20_7_real;
      end
      6'b001000 : begin
        _zz_4474_ = int_reg_array_20_8_imag;
        _zz_4475_ = int_reg_array_20_8_real;
      end
      6'b001001 : begin
        _zz_4474_ = int_reg_array_20_9_imag;
        _zz_4475_ = int_reg_array_20_9_real;
      end
      6'b001010 : begin
        _zz_4474_ = int_reg_array_20_10_imag;
        _zz_4475_ = int_reg_array_20_10_real;
      end
      6'b001011 : begin
        _zz_4474_ = int_reg_array_20_11_imag;
        _zz_4475_ = int_reg_array_20_11_real;
      end
      6'b001100 : begin
        _zz_4474_ = int_reg_array_20_12_imag;
        _zz_4475_ = int_reg_array_20_12_real;
      end
      6'b001101 : begin
        _zz_4474_ = int_reg_array_20_13_imag;
        _zz_4475_ = int_reg_array_20_13_real;
      end
      6'b001110 : begin
        _zz_4474_ = int_reg_array_20_14_imag;
        _zz_4475_ = int_reg_array_20_14_real;
      end
      6'b001111 : begin
        _zz_4474_ = int_reg_array_20_15_imag;
        _zz_4475_ = int_reg_array_20_15_real;
      end
      6'b010000 : begin
        _zz_4474_ = int_reg_array_20_16_imag;
        _zz_4475_ = int_reg_array_20_16_real;
      end
      6'b010001 : begin
        _zz_4474_ = int_reg_array_20_17_imag;
        _zz_4475_ = int_reg_array_20_17_real;
      end
      6'b010010 : begin
        _zz_4474_ = int_reg_array_20_18_imag;
        _zz_4475_ = int_reg_array_20_18_real;
      end
      6'b010011 : begin
        _zz_4474_ = int_reg_array_20_19_imag;
        _zz_4475_ = int_reg_array_20_19_real;
      end
      6'b010100 : begin
        _zz_4474_ = int_reg_array_20_20_imag;
        _zz_4475_ = int_reg_array_20_20_real;
      end
      6'b010101 : begin
        _zz_4474_ = int_reg_array_20_21_imag;
        _zz_4475_ = int_reg_array_20_21_real;
      end
      6'b010110 : begin
        _zz_4474_ = int_reg_array_20_22_imag;
        _zz_4475_ = int_reg_array_20_22_real;
      end
      6'b010111 : begin
        _zz_4474_ = int_reg_array_20_23_imag;
        _zz_4475_ = int_reg_array_20_23_real;
      end
      6'b011000 : begin
        _zz_4474_ = int_reg_array_20_24_imag;
        _zz_4475_ = int_reg_array_20_24_real;
      end
      6'b011001 : begin
        _zz_4474_ = int_reg_array_20_25_imag;
        _zz_4475_ = int_reg_array_20_25_real;
      end
      6'b011010 : begin
        _zz_4474_ = int_reg_array_20_26_imag;
        _zz_4475_ = int_reg_array_20_26_real;
      end
      6'b011011 : begin
        _zz_4474_ = int_reg_array_20_27_imag;
        _zz_4475_ = int_reg_array_20_27_real;
      end
      6'b011100 : begin
        _zz_4474_ = int_reg_array_20_28_imag;
        _zz_4475_ = int_reg_array_20_28_real;
      end
      6'b011101 : begin
        _zz_4474_ = int_reg_array_20_29_imag;
        _zz_4475_ = int_reg_array_20_29_real;
      end
      6'b011110 : begin
        _zz_4474_ = int_reg_array_20_30_imag;
        _zz_4475_ = int_reg_array_20_30_real;
      end
      6'b011111 : begin
        _zz_4474_ = int_reg_array_20_31_imag;
        _zz_4475_ = int_reg_array_20_31_real;
      end
      6'b100000 : begin
        _zz_4474_ = int_reg_array_20_32_imag;
        _zz_4475_ = int_reg_array_20_32_real;
      end
      6'b100001 : begin
        _zz_4474_ = int_reg_array_20_33_imag;
        _zz_4475_ = int_reg_array_20_33_real;
      end
      6'b100010 : begin
        _zz_4474_ = int_reg_array_20_34_imag;
        _zz_4475_ = int_reg_array_20_34_real;
      end
      6'b100011 : begin
        _zz_4474_ = int_reg_array_20_35_imag;
        _zz_4475_ = int_reg_array_20_35_real;
      end
      6'b100100 : begin
        _zz_4474_ = int_reg_array_20_36_imag;
        _zz_4475_ = int_reg_array_20_36_real;
      end
      6'b100101 : begin
        _zz_4474_ = int_reg_array_20_37_imag;
        _zz_4475_ = int_reg_array_20_37_real;
      end
      6'b100110 : begin
        _zz_4474_ = int_reg_array_20_38_imag;
        _zz_4475_ = int_reg_array_20_38_real;
      end
      6'b100111 : begin
        _zz_4474_ = int_reg_array_20_39_imag;
        _zz_4475_ = int_reg_array_20_39_real;
      end
      6'b101000 : begin
        _zz_4474_ = int_reg_array_20_40_imag;
        _zz_4475_ = int_reg_array_20_40_real;
      end
      6'b101001 : begin
        _zz_4474_ = int_reg_array_20_41_imag;
        _zz_4475_ = int_reg_array_20_41_real;
      end
      6'b101010 : begin
        _zz_4474_ = int_reg_array_20_42_imag;
        _zz_4475_ = int_reg_array_20_42_real;
      end
      6'b101011 : begin
        _zz_4474_ = int_reg_array_20_43_imag;
        _zz_4475_ = int_reg_array_20_43_real;
      end
      6'b101100 : begin
        _zz_4474_ = int_reg_array_20_44_imag;
        _zz_4475_ = int_reg_array_20_44_real;
      end
      6'b101101 : begin
        _zz_4474_ = int_reg_array_20_45_imag;
        _zz_4475_ = int_reg_array_20_45_real;
      end
      6'b101110 : begin
        _zz_4474_ = int_reg_array_20_46_imag;
        _zz_4475_ = int_reg_array_20_46_real;
      end
      6'b101111 : begin
        _zz_4474_ = int_reg_array_20_47_imag;
        _zz_4475_ = int_reg_array_20_47_real;
      end
      6'b110000 : begin
        _zz_4474_ = int_reg_array_20_48_imag;
        _zz_4475_ = int_reg_array_20_48_real;
      end
      6'b110001 : begin
        _zz_4474_ = int_reg_array_20_49_imag;
        _zz_4475_ = int_reg_array_20_49_real;
      end
      6'b110010 : begin
        _zz_4474_ = int_reg_array_20_50_imag;
        _zz_4475_ = int_reg_array_20_50_real;
      end
      6'b110011 : begin
        _zz_4474_ = int_reg_array_20_51_imag;
        _zz_4475_ = int_reg_array_20_51_real;
      end
      6'b110100 : begin
        _zz_4474_ = int_reg_array_20_52_imag;
        _zz_4475_ = int_reg_array_20_52_real;
      end
      6'b110101 : begin
        _zz_4474_ = int_reg_array_20_53_imag;
        _zz_4475_ = int_reg_array_20_53_real;
      end
      6'b110110 : begin
        _zz_4474_ = int_reg_array_20_54_imag;
        _zz_4475_ = int_reg_array_20_54_real;
      end
      6'b110111 : begin
        _zz_4474_ = int_reg_array_20_55_imag;
        _zz_4475_ = int_reg_array_20_55_real;
      end
      6'b111000 : begin
        _zz_4474_ = int_reg_array_20_56_imag;
        _zz_4475_ = int_reg_array_20_56_real;
      end
      6'b111001 : begin
        _zz_4474_ = int_reg_array_20_57_imag;
        _zz_4475_ = int_reg_array_20_57_real;
      end
      6'b111010 : begin
        _zz_4474_ = int_reg_array_20_58_imag;
        _zz_4475_ = int_reg_array_20_58_real;
      end
      6'b111011 : begin
        _zz_4474_ = int_reg_array_20_59_imag;
        _zz_4475_ = int_reg_array_20_59_real;
      end
      6'b111100 : begin
        _zz_4474_ = int_reg_array_20_60_imag;
        _zz_4475_ = int_reg_array_20_60_real;
      end
      6'b111101 : begin
        _zz_4474_ = int_reg_array_20_61_imag;
        _zz_4475_ = int_reg_array_20_61_real;
      end
      6'b111110 : begin
        _zz_4474_ = int_reg_array_20_62_imag;
        _zz_4475_ = int_reg_array_20_62_real;
      end
      default : begin
        _zz_4474_ = int_reg_array_20_63_imag;
        _zz_4475_ = int_reg_array_20_63_real;
      end
    endcase
  end

  always @(*) begin
    case(_zz_1466_)
      6'b000000 : begin
        _zz_4476_ = int_reg_array_21_0_imag;
        _zz_4477_ = int_reg_array_21_0_real;
      end
      6'b000001 : begin
        _zz_4476_ = int_reg_array_21_1_imag;
        _zz_4477_ = int_reg_array_21_1_real;
      end
      6'b000010 : begin
        _zz_4476_ = int_reg_array_21_2_imag;
        _zz_4477_ = int_reg_array_21_2_real;
      end
      6'b000011 : begin
        _zz_4476_ = int_reg_array_21_3_imag;
        _zz_4477_ = int_reg_array_21_3_real;
      end
      6'b000100 : begin
        _zz_4476_ = int_reg_array_21_4_imag;
        _zz_4477_ = int_reg_array_21_4_real;
      end
      6'b000101 : begin
        _zz_4476_ = int_reg_array_21_5_imag;
        _zz_4477_ = int_reg_array_21_5_real;
      end
      6'b000110 : begin
        _zz_4476_ = int_reg_array_21_6_imag;
        _zz_4477_ = int_reg_array_21_6_real;
      end
      6'b000111 : begin
        _zz_4476_ = int_reg_array_21_7_imag;
        _zz_4477_ = int_reg_array_21_7_real;
      end
      6'b001000 : begin
        _zz_4476_ = int_reg_array_21_8_imag;
        _zz_4477_ = int_reg_array_21_8_real;
      end
      6'b001001 : begin
        _zz_4476_ = int_reg_array_21_9_imag;
        _zz_4477_ = int_reg_array_21_9_real;
      end
      6'b001010 : begin
        _zz_4476_ = int_reg_array_21_10_imag;
        _zz_4477_ = int_reg_array_21_10_real;
      end
      6'b001011 : begin
        _zz_4476_ = int_reg_array_21_11_imag;
        _zz_4477_ = int_reg_array_21_11_real;
      end
      6'b001100 : begin
        _zz_4476_ = int_reg_array_21_12_imag;
        _zz_4477_ = int_reg_array_21_12_real;
      end
      6'b001101 : begin
        _zz_4476_ = int_reg_array_21_13_imag;
        _zz_4477_ = int_reg_array_21_13_real;
      end
      6'b001110 : begin
        _zz_4476_ = int_reg_array_21_14_imag;
        _zz_4477_ = int_reg_array_21_14_real;
      end
      6'b001111 : begin
        _zz_4476_ = int_reg_array_21_15_imag;
        _zz_4477_ = int_reg_array_21_15_real;
      end
      6'b010000 : begin
        _zz_4476_ = int_reg_array_21_16_imag;
        _zz_4477_ = int_reg_array_21_16_real;
      end
      6'b010001 : begin
        _zz_4476_ = int_reg_array_21_17_imag;
        _zz_4477_ = int_reg_array_21_17_real;
      end
      6'b010010 : begin
        _zz_4476_ = int_reg_array_21_18_imag;
        _zz_4477_ = int_reg_array_21_18_real;
      end
      6'b010011 : begin
        _zz_4476_ = int_reg_array_21_19_imag;
        _zz_4477_ = int_reg_array_21_19_real;
      end
      6'b010100 : begin
        _zz_4476_ = int_reg_array_21_20_imag;
        _zz_4477_ = int_reg_array_21_20_real;
      end
      6'b010101 : begin
        _zz_4476_ = int_reg_array_21_21_imag;
        _zz_4477_ = int_reg_array_21_21_real;
      end
      6'b010110 : begin
        _zz_4476_ = int_reg_array_21_22_imag;
        _zz_4477_ = int_reg_array_21_22_real;
      end
      6'b010111 : begin
        _zz_4476_ = int_reg_array_21_23_imag;
        _zz_4477_ = int_reg_array_21_23_real;
      end
      6'b011000 : begin
        _zz_4476_ = int_reg_array_21_24_imag;
        _zz_4477_ = int_reg_array_21_24_real;
      end
      6'b011001 : begin
        _zz_4476_ = int_reg_array_21_25_imag;
        _zz_4477_ = int_reg_array_21_25_real;
      end
      6'b011010 : begin
        _zz_4476_ = int_reg_array_21_26_imag;
        _zz_4477_ = int_reg_array_21_26_real;
      end
      6'b011011 : begin
        _zz_4476_ = int_reg_array_21_27_imag;
        _zz_4477_ = int_reg_array_21_27_real;
      end
      6'b011100 : begin
        _zz_4476_ = int_reg_array_21_28_imag;
        _zz_4477_ = int_reg_array_21_28_real;
      end
      6'b011101 : begin
        _zz_4476_ = int_reg_array_21_29_imag;
        _zz_4477_ = int_reg_array_21_29_real;
      end
      6'b011110 : begin
        _zz_4476_ = int_reg_array_21_30_imag;
        _zz_4477_ = int_reg_array_21_30_real;
      end
      6'b011111 : begin
        _zz_4476_ = int_reg_array_21_31_imag;
        _zz_4477_ = int_reg_array_21_31_real;
      end
      6'b100000 : begin
        _zz_4476_ = int_reg_array_21_32_imag;
        _zz_4477_ = int_reg_array_21_32_real;
      end
      6'b100001 : begin
        _zz_4476_ = int_reg_array_21_33_imag;
        _zz_4477_ = int_reg_array_21_33_real;
      end
      6'b100010 : begin
        _zz_4476_ = int_reg_array_21_34_imag;
        _zz_4477_ = int_reg_array_21_34_real;
      end
      6'b100011 : begin
        _zz_4476_ = int_reg_array_21_35_imag;
        _zz_4477_ = int_reg_array_21_35_real;
      end
      6'b100100 : begin
        _zz_4476_ = int_reg_array_21_36_imag;
        _zz_4477_ = int_reg_array_21_36_real;
      end
      6'b100101 : begin
        _zz_4476_ = int_reg_array_21_37_imag;
        _zz_4477_ = int_reg_array_21_37_real;
      end
      6'b100110 : begin
        _zz_4476_ = int_reg_array_21_38_imag;
        _zz_4477_ = int_reg_array_21_38_real;
      end
      6'b100111 : begin
        _zz_4476_ = int_reg_array_21_39_imag;
        _zz_4477_ = int_reg_array_21_39_real;
      end
      6'b101000 : begin
        _zz_4476_ = int_reg_array_21_40_imag;
        _zz_4477_ = int_reg_array_21_40_real;
      end
      6'b101001 : begin
        _zz_4476_ = int_reg_array_21_41_imag;
        _zz_4477_ = int_reg_array_21_41_real;
      end
      6'b101010 : begin
        _zz_4476_ = int_reg_array_21_42_imag;
        _zz_4477_ = int_reg_array_21_42_real;
      end
      6'b101011 : begin
        _zz_4476_ = int_reg_array_21_43_imag;
        _zz_4477_ = int_reg_array_21_43_real;
      end
      6'b101100 : begin
        _zz_4476_ = int_reg_array_21_44_imag;
        _zz_4477_ = int_reg_array_21_44_real;
      end
      6'b101101 : begin
        _zz_4476_ = int_reg_array_21_45_imag;
        _zz_4477_ = int_reg_array_21_45_real;
      end
      6'b101110 : begin
        _zz_4476_ = int_reg_array_21_46_imag;
        _zz_4477_ = int_reg_array_21_46_real;
      end
      6'b101111 : begin
        _zz_4476_ = int_reg_array_21_47_imag;
        _zz_4477_ = int_reg_array_21_47_real;
      end
      6'b110000 : begin
        _zz_4476_ = int_reg_array_21_48_imag;
        _zz_4477_ = int_reg_array_21_48_real;
      end
      6'b110001 : begin
        _zz_4476_ = int_reg_array_21_49_imag;
        _zz_4477_ = int_reg_array_21_49_real;
      end
      6'b110010 : begin
        _zz_4476_ = int_reg_array_21_50_imag;
        _zz_4477_ = int_reg_array_21_50_real;
      end
      6'b110011 : begin
        _zz_4476_ = int_reg_array_21_51_imag;
        _zz_4477_ = int_reg_array_21_51_real;
      end
      6'b110100 : begin
        _zz_4476_ = int_reg_array_21_52_imag;
        _zz_4477_ = int_reg_array_21_52_real;
      end
      6'b110101 : begin
        _zz_4476_ = int_reg_array_21_53_imag;
        _zz_4477_ = int_reg_array_21_53_real;
      end
      6'b110110 : begin
        _zz_4476_ = int_reg_array_21_54_imag;
        _zz_4477_ = int_reg_array_21_54_real;
      end
      6'b110111 : begin
        _zz_4476_ = int_reg_array_21_55_imag;
        _zz_4477_ = int_reg_array_21_55_real;
      end
      6'b111000 : begin
        _zz_4476_ = int_reg_array_21_56_imag;
        _zz_4477_ = int_reg_array_21_56_real;
      end
      6'b111001 : begin
        _zz_4476_ = int_reg_array_21_57_imag;
        _zz_4477_ = int_reg_array_21_57_real;
      end
      6'b111010 : begin
        _zz_4476_ = int_reg_array_21_58_imag;
        _zz_4477_ = int_reg_array_21_58_real;
      end
      6'b111011 : begin
        _zz_4476_ = int_reg_array_21_59_imag;
        _zz_4477_ = int_reg_array_21_59_real;
      end
      6'b111100 : begin
        _zz_4476_ = int_reg_array_21_60_imag;
        _zz_4477_ = int_reg_array_21_60_real;
      end
      6'b111101 : begin
        _zz_4476_ = int_reg_array_21_61_imag;
        _zz_4477_ = int_reg_array_21_61_real;
      end
      6'b111110 : begin
        _zz_4476_ = int_reg_array_21_62_imag;
        _zz_4477_ = int_reg_array_21_62_real;
      end
      default : begin
        _zz_4476_ = int_reg_array_21_63_imag;
        _zz_4477_ = int_reg_array_21_63_real;
      end
    endcase
  end

  always @(*) begin
    case(_zz_1535_)
      6'b000000 : begin
        _zz_4478_ = int_reg_array_22_0_imag;
        _zz_4479_ = int_reg_array_22_0_real;
      end
      6'b000001 : begin
        _zz_4478_ = int_reg_array_22_1_imag;
        _zz_4479_ = int_reg_array_22_1_real;
      end
      6'b000010 : begin
        _zz_4478_ = int_reg_array_22_2_imag;
        _zz_4479_ = int_reg_array_22_2_real;
      end
      6'b000011 : begin
        _zz_4478_ = int_reg_array_22_3_imag;
        _zz_4479_ = int_reg_array_22_3_real;
      end
      6'b000100 : begin
        _zz_4478_ = int_reg_array_22_4_imag;
        _zz_4479_ = int_reg_array_22_4_real;
      end
      6'b000101 : begin
        _zz_4478_ = int_reg_array_22_5_imag;
        _zz_4479_ = int_reg_array_22_5_real;
      end
      6'b000110 : begin
        _zz_4478_ = int_reg_array_22_6_imag;
        _zz_4479_ = int_reg_array_22_6_real;
      end
      6'b000111 : begin
        _zz_4478_ = int_reg_array_22_7_imag;
        _zz_4479_ = int_reg_array_22_7_real;
      end
      6'b001000 : begin
        _zz_4478_ = int_reg_array_22_8_imag;
        _zz_4479_ = int_reg_array_22_8_real;
      end
      6'b001001 : begin
        _zz_4478_ = int_reg_array_22_9_imag;
        _zz_4479_ = int_reg_array_22_9_real;
      end
      6'b001010 : begin
        _zz_4478_ = int_reg_array_22_10_imag;
        _zz_4479_ = int_reg_array_22_10_real;
      end
      6'b001011 : begin
        _zz_4478_ = int_reg_array_22_11_imag;
        _zz_4479_ = int_reg_array_22_11_real;
      end
      6'b001100 : begin
        _zz_4478_ = int_reg_array_22_12_imag;
        _zz_4479_ = int_reg_array_22_12_real;
      end
      6'b001101 : begin
        _zz_4478_ = int_reg_array_22_13_imag;
        _zz_4479_ = int_reg_array_22_13_real;
      end
      6'b001110 : begin
        _zz_4478_ = int_reg_array_22_14_imag;
        _zz_4479_ = int_reg_array_22_14_real;
      end
      6'b001111 : begin
        _zz_4478_ = int_reg_array_22_15_imag;
        _zz_4479_ = int_reg_array_22_15_real;
      end
      6'b010000 : begin
        _zz_4478_ = int_reg_array_22_16_imag;
        _zz_4479_ = int_reg_array_22_16_real;
      end
      6'b010001 : begin
        _zz_4478_ = int_reg_array_22_17_imag;
        _zz_4479_ = int_reg_array_22_17_real;
      end
      6'b010010 : begin
        _zz_4478_ = int_reg_array_22_18_imag;
        _zz_4479_ = int_reg_array_22_18_real;
      end
      6'b010011 : begin
        _zz_4478_ = int_reg_array_22_19_imag;
        _zz_4479_ = int_reg_array_22_19_real;
      end
      6'b010100 : begin
        _zz_4478_ = int_reg_array_22_20_imag;
        _zz_4479_ = int_reg_array_22_20_real;
      end
      6'b010101 : begin
        _zz_4478_ = int_reg_array_22_21_imag;
        _zz_4479_ = int_reg_array_22_21_real;
      end
      6'b010110 : begin
        _zz_4478_ = int_reg_array_22_22_imag;
        _zz_4479_ = int_reg_array_22_22_real;
      end
      6'b010111 : begin
        _zz_4478_ = int_reg_array_22_23_imag;
        _zz_4479_ = int_reg_array_22_23_real;
      end
      6'b011000 : begin
        _zz_4478_ = int_reg_array_22_24_imag;
        _zz_4479_ = int_reg_array_22_24_real;
      end
      6'b011001 : begin
        _zz_4478_ = int_reg_array_22_25_imag;
        _zz_4479_ = int_reg_array_22_25_real;
      end
      6'b011010 : begin
        _zz_4478_ = int_reg_array_22_26_imag;
        _zz_4479_ = int_reg_array_22_26_real;
      end
      6'b011011 : begin
        _zz_4478_ = int_reg_array_22_27_imag;
        _zz_4479_ = int_reg_array_22_27_real;
      end
      6'b011100 : begin
        _zz_4478_ = int_reg_array_22_28_imag;
        _zz_4479_ = int_reg_array_22_28_real;
      end
      6'b011101 : begin
        _zz_4478_ = int_reg_array_22_29_imag;
        _zz_4479_ = int_reg_array_22_29_real;
      end
      6'b011110 : begin
        _zz_4478_ = int_reg_array_22_30_imag;
        _zz_4479_ = int_reg_array_22_30_real;
      end
      6'b011111 : begin
        _zz_4478_ = int_reg_array_22_31_imag;
        _zz_4479_ = int_reg_array_22_31_real;
      end
      6'b100000 : begin
        _zz_4478_ = int_reg_array_22_32_imag;
        _zz_4479_ = int_reg_array_22_32_real;
      end
      6'b100001 : begin
        _zz_4478_ = int_reg_array_22_33_imag;
        _zz_4479_ = int_reg_array_22_33_real;
      end
      6'b100010 : begin
        _zz_4478_ = int_reg_array_22_34_imag;
        _zz_4479_ = int_reg_array_22_34_real;
      end
      6'b100011 : begin
        _zz_4478_ = int_reg_array_22_35_imag;
        _zz_4479_ = int_reg_array_22_35_real;
      end
      6'b100100 : begin
        _zz_4478_ = int_reg_array_22_36_imag;
        _zz_4479_ = int_reg_array_22_36_real;
      end
      6'b100101 : begin
        _zz_4478_ = int_reg_array_22_37_imag;
        _zz_4479_ = int_reg_array_22_37_real;
      end
      6'b100110 : begin
        _zz_4478_ = int_reg_array_22_38_imag;
        _zz_4479_ = int_reg_array_22_38_real;
      end
      6'b100111 : begin
        _zz_4478_ = int_reg_array_22_39_imag;
        _zz_4479_ = int_reg_array_22_39_real;
      end
      6'b101000 : begin
        _zz_4478_ = int_reg_array_22_40_imag;
        _zz_4479_ = int_reg_array_22_40_real;
      end
      6'b101001 : begin
        _zz_4478_ = int_reg_array_22_41_imag;
        _zz_4479_ = int_reg_array_22_41_real;
      end
      6'b101010 : begin
        _zz_4478_ = int_reg_array_22_42_imag;
        _zz_4479_ = int_reg_array_22_42_real;
      end
      6'b101011 : begin
        _zz_4478_ = int_reg_array_22_43_imag;
        _zz_4479_ = int_reg_array_22_43_real;
      end
      6'b101100 : begin
        _zz_4478_ = int_reg_array_22_44_imag;
        _zz_4479_ = int_reg_array_22_44_real;
      end
      6'b101101 : begin
        _zz_4478_ = int_reg_array_22_45_imag;
        _zz_4479_ = int_reg_array_22_45_real;
      end
      6'b101110 : begin
        _zz_4478_ = int_reg_array_22_46_imag;
        _zz_4479_ = int_reg_array_22_46_real;
      end
      6'b101111 : begin
        _zz_4478_ = int_reg_array_22_47_imag;
        _zz_4479_ = int_reg_array_22_47_real;
      end
      6'b110000 : begin
        _zz_4478_ = int_reg_array_22_48_imag;
        _zz_4479_ = int_reg_array_22_48_real;
      end
      6'b110001 : begin
        _zz_4478_ = int_reg_array_22_49_imag;
        _zz_4479_ = int_reg_array_22_49_real;
      end
      6'b110010 : begin
        _zz_4478_ = int_reg_array_22_50_imag;
        _zz_4479_ = int_reg_array_22_50_real;
      end
      6'b110011 : begin
        _zz_4478_ = int_reg_array_22_51_imag;
        _zz_4479_ = int_reg_array_22_51_real;
      end
      6'b110100 : begin
        _zz_4478_ = int_reg_array_22_52_imag;
        _zz_4479_ = int_reg_array_22_52_real;
      end
      6'b110101 : begin
        _zz_4478_ = int_reg_array_22_53_imag;
        _zz_4479_ = int_reg_array_22_53_real;
      end
      6'b110110 : begin
        _zz_4478_ = int_reg_array_22_54_imag;
        _zz_4479_ = int_reg_array_22_54_real;
      end
      6'b110111 : begin
        _zz_4478_ = int_reg_array_22_55_imag;
        _zz_4479_ = int_reg_array_22_55_real;
      end
      6'b111000 : begin
        _zz_4478_ = int_reg_array_22_56_imag;
        _zz_4479_ = int_reg_array_22_56_real;
      end
      6'b111001 : begin
        _zz_4478_ = int_reg_array_22_57_imag;
        _zz_4479_ = int_reg_array_22_57_real;
      end
      6'b111010 : begin
        _zz_4478_ = int_reg_array_22_58_imag;
        _zz_4479_ = int_reg_array_22_58_real;
      end
      6'b111011 : begin
        _zz_4478_ = int_reg_array_22_59_imag;
        _zz_4479_ = int_reg_array_22_59_real;
      end
      6'b111100 : begin
        _zz_4478_ = int_reg_array_22_60_imag;
        _zz_4479_ = int_reg_array_22_60_real;
      end
      6'b111101 : begin
        _zz_4478_ = int_reg_array_22_61_imag;
        _zz_4479_ = int_reg_array_22_61_real;
      end
      6'b111110 : begin
        _zz_4478_ = int_reg_array_22_62_imag;
        _zz_4479_ = int_reg_array_22_62_real;
      end
      default : begin
        _zz_4478_ = int_reg_array_22_63_imag;
        _zz_4479_ = int_reg_array_22_63_real;
      end
    endcase
  end

  always @(*) begin
    case(_zz_1604_)
      6'b000000 : begin
        _zz_4480_ = int_reg_array_23_0_imag;
        _zz_4481_ = int_reg_array_23_0_real;
      end
      6'b000001 : begin
        _zz_4480_ = int_reg_array_23_1_imag;
        _zz_4481_ = int_reg_array_23_1_real;
      end
      6'b000010 : begin
        _zz_4480_ = int_reg_array_23_2_imag;
        _zz_4481_ = int_reg_array_23_2_real;
      end
      6'b000011 : begin
        _zz_4480_ = int_reg_array_23_3_imag;
        _zz_4481_ = int_reg_array_23_3_real;
      end
      6'b000100 : begin
        _zz_4480_ = int_reg_array_23_4_imag;
        _zz_4481_ = int_reg_array_23_4_real;
      end
      6'b000101 : begin
        _zz_4480_ = int_reg_array_23_5_imag;
        _zz_4481_ = int_reg_array_23_5_real;
      end
      6'b000110 : begin
        _zz_4480_ = int_reg_array_23_6_imag;
        _zz_4481_ = int_reg_array_23_6_real;
      end
      6'b000111 : begin
        _zz_4480_ = int_reg_array_23_7_imag;
        _zz_4481_ = int_reg_array_23_7_real;
      end
      6'b001000 : begin
        _zz_4480_ = int_reg_array_23_8_imag;
        _zz_4481_ = int_reg_array_23_8_real;
      end
      6'b001001 : begin
        _zz_4480_ = int_reg_array_23_9_imag;
        _zz_4481_ = int_reg_array_23_9_real;
      end
      6'b001010 : begin
        _zz_4480_ = int_reg_array_23_10_imag;
        _zz_4481_ = int_reg_array_23_10_real;
      end
      6'b001011 : begin
        _zz_4480_ = int_reg_array_23_11_imag;
        _zz_4481_ = int_reg_array_23_11_real;
      end
      6'b001100 : begin
        _zz_4480_ = int_reg_array_23_12_imag;
        _zz_4481_ = int_reg_array_23_12_real;
      end
      6'b001101 : begin
        _zz_4480_ = int_reg_array_23_13_imag;
        _zz_4481_ = int_reg_array_23_13_real;
      end
      6'b001110 : begin
        _zz_4480_ = int_reg_array_23_14_imag;
        _zz_4481_ = int_reg_array_23_14_real;
      end
      6'b001111 : begin
        _zz_4480_ = int_reg_array_23_15_imag;
        _zz_4481_ = int_reg_array_23_15_real;
      end
      6'b010000 : begin
        _zz_4480_ = int_reg_array_23_16_imag;
        _zz_4481_ = int_reg_array_23_16_real;
      end
      6'b010001 : begin
        _zz_4480_ = int_reg_array_23_17_imag;
        _zz_4481_ = int_reg_array_23_17_real;
      end
      6'b010010 : begin
        _zz_4480_ = int_reg_array_23_18_imag;
        _zz_4481_ = int_reg_array_23_18_real;
      end
      6'b010011 : begin
        _zz_4480_ = int_reg_array_23_19_imag;
        _zz_4481_ = int_reg_array_23_19_real;
      end
      6'b010100 : begin
        _zz_4480_ = int_reg_array_23_20_imag;
        _zz_4481_ = int_reg_array_23_20_real;
      end
      6'b010101 : begin
        _zz_4480_ = int_reg_array_23_21_imag;
        _zz_4481_ = int_reg_array_23_21_real;
      end
      6'b010110 : begin
        _zz_4480_ = int_reg_array_23_22_imag;
        _zz_4481_ = int_reg_array_23_22_real;
      end
      6'b010111 : begin
        _zz_4480_ = int_reg_array_23_23_imag;
        _zz_4481_ = int_reg_array_23_23_real;
      end
      6'b011000 : begin
        _zz_4480_ = int_reg_array_23_24_imag;
        _zz_4481_ = int_reg_array_23_24_real;
      end
      6'b011001 : begin
        _zz_4480_ = int_reg_array_23_25_imag;
        _zz_4481_ = int_reg_array_23_25_real;
      end
      6'b011010 : begin
        _zz_4480_ = int_reg_array_23_26_imag;
        _zz_4481_ = int_reg_array_23_26_real;
      end
      6'b011011 : begin
        _zz_4480_ = int_reg_array_23_27_imag;
        _zz_4481_ = int_reg_array_23_27_real;
      end
      6'b011100 : begin
        _zz_4480_ = int_reg_array_23_28_imag;
        _zz_4481_ = int_reg_array_23_28_real;
      end
      6'b011101 : begin
        _zz_4480_ = int_reg_array_23_29_imag;
        _zz_4481_ = int_reg_array_23_29_real;
      end
      6'b011110 : begin
        _zz_4480_ = int_reg_array_23_30_imag;
        _zz_4481_ = int_reg_array_23_30_real;
      end
      6'b011111 : begin
        _zz_4480_ = int_reg_array_23_31_imag;
        _zz_4481_ = int_reg_array_23_31_real;
      end
      6'b100000 : begin
        _zz_4480_ = int_reg_array_23_32_imag;
        _zz_4481_ = int_reg_array_23_32_real;
      end
      6'b100001 : begin
        _zz_4480_ = int_reg_array_23_33_imag;
        _zz_4481_ = int_reg_array_23_33_real;
      end
      6'b100010 : begin
        _zz_4480_ = int_reg_array_23_34_imag;
        _zz_4481_ = int_reg_array_23_34_real;
      end
      6'b100011 : begin
        _zz_4480_ = int_reg_array_23_35_imag;
        _zz_4481_ = int_reg_array_23_35_real;
      end
      6'b100100 : begin
        _zz_4480_ = int_reg_array_23_36_imag;
        _zz_4481_ = int_reg_array_23_36_real;
      end
      6'b100101 : begin
        _zz_4480_ = int_reg_array_23_37_imag;
        _zz_4481_ = int_reg_array_23_37_real;
      end
      6'b100110 : begin
        _zz_4480_ = int_reg_array_23_38_imag;
        _zz_4481_ = int_reg_array_23_38_real;
      end
      6'b100111 : begin
        _zz_4480_ = int_reg_array_23_39_imag;
        _zz_4481_ = int_reg_array_23_39_real;
      end
      6'b101000 : begin
        _zz_4480_ = int_reg_array_23_40_imag;
        _zz_4481_ = int_reg_array_23_40_real;
      end
      6'b101001 : begin
        _zz_4480_ = int_reg_array_23_41_imag;
        _zz_4481_ = int_reg_array_23_41_real;
      end
      6'b101010 : begin
        _zz_4480_ = int_reg_array_23_42_imag;
        _zz_4481_ = int_reg_array_23_42_real;
      end
      6'b101011 : begin
        _zz_4480_ = int_reg_array_23_43_imag;
        _zz_4481_ = int_reg_array_23_43_real;
      end
      6'b101100 : begin
        _zz_4480_ = int_reg_array_23_44_imag;
        _zz_4481_ = int_reg_array_23_44_real;
      end
      6'b101101 : begin
        _zz_4480_ = int_reg_array_23_45_imag;
        _zz_4481_ = int_reg_array_23_45_real;
      end
      6'b101110 : begin
        _zz_4480_ = int_reg_array_23_46_imag;
        _zz_4481_ = int_reg_array_23_46_real;
      end
      6'b101111 : begin
        _zz_4480_ = int_reg_array_23_47_imag;
        _zz_4481_ = int_reg_array_23_47_real;
      end
      6'b110000 : begin
        _zz_4480_ = int_reg_array_23_48_imag;
        _zz_4481_ = int_reg_array_23_48_real;
      end
      6'b110001 : begin
        _zz_4480_ = int_reg_array_23_49_imag;
        _zz_4481_ = int_reg_array_23_49_real;
      end
      6'b110010 : begin
        _zz_4480_ = int_reg_array_23_50_imag;
        _zz_4481_ = int_reg_array_23_50_real;
      end
      6'b110011 : begin
        _zz_4480_ = int_reg_array_23_51_imag;
        _zz_4481_ = int_reg_array_23_51_real;
      end
      6'b110100 : begin
        _zz_4480_ = int_reg_array_23_52_imag;
        _zz_4481_ = int_reg_array_23_52_real;
      end
      6'b110101 : begin
        _zz_4480_ = int_reg_array_23_53_imag;
        _zz_4481_ = int_reg_array_23_53_real;
      end
      6'b110110 : begin
        _zz_4480_ = int_reg_array_23_54_imag;
        _zz_4481_ = int_reg_array_23_54_real;
      end
      6'b110111 : begin
        _zz_4480_ = int_reg_array_23_55_imag;
        _zz_4481_ = int_reg_array_23_55_real;
      end
      6'b111000 : begin
        _zz_4480_ = int_reg_array_23_56_imag;
        _zz_4481_ = int_reg_array_23_56_real;
      end
      6'b111001 : begin
        _zz_4480_ = int_reg_array_23_57_imag;
        _zz_4481_ = int_reg_array_23_57_real;
      end
      6'b111010 : begin
        _zz_4480_ = int_reg_array_23_58_imag;
        _zz_4481_ = int_reg_array_23_58_real;
      end
      6'b111011 : begin
        _zz_4480_ = int_reg_array_23_59_imag;
        _zz_4481_ = int_reg_array_23_59_real;
      end
      6'b111100 : begin
        _zz_4480_ = int_reg_array_23_60_imag;
        _zz_4481_ = int_reg_array_23_60_real;
      end
      6'b111101 : begin
        _zz_4480_ = int_reg_array_23_61_imag;
        _zz_4481_ = int_reg_array_23_61_real;
      end
      6'b111110 : begin
        _zz_4480_ = int_reg_array_23_62_imag;
        _zz_4481_ = int_reg_array_23_62_real;
      end
      default : begin
        _zz_4480_ = int_reg_array_23_63_imag;
        _zz_4481_ = int_reg_array_23_63_real;
      end
    endcase
  end

  always @(*) begin
    case(_zz_1673_)
      6'b000000 : begin
        _zz_4482_ = int_reg_array_24_0_imag;
        _zz_4483_ = int_reg_array_24_0_real;
      end
      6'b000001 : begin
        _zz_4482_ = int_reg_array_24_1_imag;
        _zz_4483_ = int_reg_array_24_1_real;
      end
      6'b000010 : begin
        _zz_4482_ = int_reg_array_24_2_imag;
        _zz_4483_ = int_reg_array_24_2_real;
      end
      6'b000011 : begin
        _zz_4482_ = int_reg_array_24_3_imag;
        _zz_4483_ = int_reg_array_24_3_real;
      end
      6'b000100 : begin
        _zz_4482_ = int_reg_array_24_4_imag;
        _zz_4483_ = int_reg_array_24_4_real;
      end
      6'b000101 : begin
        _zz_4482_ = int_reg_array_24_5_imag;
        _zz_4483_ = int_reg_array_24_5_real;
      end
      6'b000110 : begin
        _zz_4482_ = int_reg_array_24_6_imag;
        _zz_4483_ = int_reg_array_24_6_real;
      end
      6'b000111 : begin
        _zz_4482_ = int_reg_array_24_7_imag;
        _zz_4483_ = int_reg_array_24_7_real;
      end
      6'b001000 : begin
        _zz_4482_ = int_reg_array_24_8_imag;
        _zz_4483_ = int_reg_array_24_8_real;
      end
      6'b001001 : begin
        _zz_4482_ = int_reg_array_24_9_imag;
        _zz_4483_ = int_reg_array_24_9_real;
      end
      6'b001010 : begin
        _zz_4482_ = int_reg_array_24_10_imag;
        _zz_4483_ = int_reg_array_24_10_real;
      end
      6'b001011 : begin
        _zz_4482_ = int_reg_array_24_11_imag;
        _zz_4483_ = int_reg_array_24_11_real;
      end
      6'b001100 : begin
        _zz_4482_ = int_reg_array_24_12_imag;
        _zz_4483_ = int_reg_array_24_12_real;
      end
      6'b001101 : begin
        _zz_4482_ = int_reg_array_24_13_imag;
        _zz_4483_ = int_reg_array_24_13_real;
      end
      6'b001110 : begin
        _zz_4482_ = int_reg_array_24_14_imag;
        _zz_4483_ = int_reg_array_24_14_real;
      end
      6'b001111 : begin
        _zz_4482_ = int_reg_array_24_15_imag;
        _zz_4483_ = int_reg_array_24_15_real;
      end
      6'b010000 : begin
        _zz_4482_ = int_reg_array_24_16_imag;
        _zz_4483_ = int_reg_array_24_16_real;
      end
      6'b010001 : begin
        _zz_4482_ = int_reg_array_24_17_imag;
        _zz_4483_ = int_reg_array_24_17_real;
      end
      6'b010010 : begin
        _zz_4482_ = int_reg_array_24_18_imag;
        _zz_4483_ = int_reg_array_24_18_real;
      end
      6'b010011 : begin
        _zz_4482_ = int_reg_array_24_19_imag;
        _zz_4483_ = int_reg_array_24_19_real;
      end
      6'b010100 : begin
        _zz_4482_ = int_reg_array_24_20_imag;
        _zz_4483_ = int_reg_array_24_20_real;
      end
      6'b010101 : begin
        _zz_4482_ = int_reg_array_24_21_imag;
        _zz_4483_ = int_reg_array_24_21_real;
      end
      6'b010110 : begin
        _zz_4482_ = int_reg_array_24_22_imag;
        _zz_4483_ = int_reg_array_24_22_real;
      end
      6'b010111 : begin
        _zz_4482_ = int_reg_array_24_23_imag;
        _zz_4483_ = int_reg_array_24_23_real;
      end
      6'b011000 : begin
        _zz_4482_ = int_reg_array_24_24_imag;
        _zz_4483_ = int_reg_array_24_24_real;
      end
      6'b011001 : begin
        _zz_4482_ = int_reg_array_24_25_imag;
        _zz_4483_ = int_reg_array_24_25_real;
      end
      6'b011010 : begin
        _zz_4482_ = int_reg_array_24_26_imag;
        _zz_4483_ = int_reg_array_24_26_real;
      end
      6'b011011 : begin
        _zz_4482_ = int_reg_array_24_27_imag;
        _zz_4483_ = int_reg_array_24_27_real;
      end
      6'b011100 : begin
        _zz_4482_ = int_reg_array_24_28_imag;
        _zz_4483_ = int_reg_array_24_28_real;
      end
      6'b011101 : begin
        _zz_4482_ = int_reg_array_24_29_imag;
        _zz_4483_ = int_reg_array_24_29_real;
      end
      6'b011110 : begin
        _zz_4482_ = int_reg_array_24_30_imag;
        _zz_4483_ = int_reg_array_24_30_real;
      end
      6'b011111 : begin
        _zz_4482_ = int_reg_array_24_31_imag;
        _zz_4483_ = int_reg_array_24_31_real;
      end
      6'b100000 : begin
        _zz_4482_ = int_reg_array_24_32_imag;
        _zz_4483_ = int_reg_array_24_32_real;
      end
      6'b100001 : begin
        _zz_4482_ = int_reg_array_24_33_imag;
        _zz_4483_ = int_reg_array_24_33_real;
      end
      6'b100010 : begin
        _zz_4482_ = int_reg_array_24_34_imag;
        _zz_4483_ = int_reg_array_24_34_real;
      end
      6'b100011 : begin
        _zz_4482_ = int_reg_array_24_35_imag;
        _zz_4483_ = int_reg_array_24_35_real;
      end
      6'b100100 : begin
        _zz_4482_ = int_reg_array_24_36_imag;
        _zz_4483_ = int_reg_array_24_36_real;
      end
      6'b100101 : begin
        _zz_4482_ = int_reg_array_24_37_imag;
        _zz_4483_ = int_reg_array_24_37_real;
      end
      6'b100110 : begin
        _zz_4482_ = int_reg_array_24_38_imag;
        _zz_4483_ = int_reg_array_24_38_real;
      end
      6'b100111 : begin
        _zz_4482_ = int_reg_array_24_39_imag;
        _zz_4483_ = int_reg_array_24_39_real;
      end
      6'b101000 : begin
        _zz_4482_ = int_reg_array_24_40_imag;
        _zz_4483_ = int_reg_array_24_40_real;
      end
      6'b101001 : begin
        _zz_4482_ = int_reg_array_24_41_imag;
        _zz_4483_ = int_reg_array_24_41_real;
      end
      6'b101010 : begin
        _zz_4482_ = int_reg_array_24_42_imag;
        _zz_4483_ = int_reg_array_24_42_real;
      end
      6'b101011 : begin
        _zz_4482_ = int_reg_array_24_43_imag;
        _zz_4483_ = int_reg_array_24_43_real;
      end
      6'b101100 : begin
        _zz_4482_ = int_reg_array_24_44_imag;
        _zz_4483_ = int_reg_array_24_44_real;
      end
      6'b101101 : begin
        _zz_4482_ = int_reg_array_24_45_imag;
        _zz_4483_ = int_reg_array_24_45_real;
      end
      6'b101110 : begin
        _zz_4482_ = int_reg_array_24_46_imag;
        _zz_4483_ = int_reg_array_24_46_real;
      end
      6'b101111 : begin
        _zz_4482_ = int_reg_array_24_47_imag;
        _zz_4483_ = int_reg_array_24_47_real;
      end
      6'b110000 : begin
        _zz_4482_ = int_reg_array_24_48_imag;
        _zz_4483_ = int_reg_array_24_48_real;
      end
      6'b110001 : begin
        _zz_4482_ = int_reg_array_24_49_imag;
        _zz_4483_ = int_reg_array_24_49_real;
      end
      6'b110010 : begin
        _zz_4482_ = int_reg_array_24_50_imag;
        _zz_4483_ = int_reg_array_24_50_real;
      end
      6'b110011 : begin
        _zz_4482_ = int_reg_array_24_51_imag;
        _zz_4483_ = int_reg_array_24_51_real;
      end
      6'b110100 : begin
        _zz_4482_ = int_reg_array_24_52_imag;
        _zz_4483_ = int_reg_array_24_52_real;
      end
      6'b110101 : begin
        _zz_4482_ = int_reg_array_24_53_imag;
        _zz_4483_ = int_reg_array_24_53_real;
      end
      6'b110110 : begin
        _zz_4482_ = int_reg_array_24_54_imag;
        _zz_4483_ = int_reg_array_24_54_real;
      end
      6'b110111 : begin
        _zz_4482_ = int_reg_array_24_55_imag;
        _zz_4483_ = int_reg_array_24_55_real;
      end
      6'b111000 : begin
        _zz_4482_ = int_reg_array_24_56_imag;
        _zz_4483_ = int_reg_array_24_56_real;
      end
      6'b111001 : begin
        _zz_4482_ = int_reg_array_24_57_imag;
        _zz_4483_ = int_reg_array_24_57_real;
      end
      6'b111010 : begin
        _zz_4482_ = int_reg_array_24_58_imag;
        _zz_4483_ = int_reg_array_24_58_real;
      end
      6'b111011 : begin
        _zz_4482_ = int_reg_array_24_59_imag;
        _zz_4483_ = int_reg_array_24_59_real;
      end
      6'b111100 : begin
        _zz_4482_ = int_reg_array_24_60_imag;
        _zz_4483_ = int_reg_array_24_60_real;
      end
      6'b111101 : begin
        _zz_4482_ = int_reg_array_24_61_imag;
        _zz_4483_ = int_reg_array_24_61_real;
      end
      6'b111110 : begin
        _zz_4482_ = int_reg_array_24_62_imag;
        _zz_4483_ = int_reg_array_24_62_real;
      end
      default : begin
        _zz_4482_ = int_reg_array_24_63_imag;
        _zz_4483_ = int_reg_array_24_63_real;
      end
    endcase
  end

  always @(*) begin
    case(_zz_1742_)
      6'b000000 : begin
        _zz_4484_ = int_reg_array_25_0_imag;
        _zz_4485_ = int_reg_array_25_0_real;
      end
      6'b000001 : begin
        _zz_4484_ = int_reg_array_25_1_imag;
        _zz_4485_ = int_reg_array_25_1_real;
      end
      6'b000010 : begin
        _zz_4484_ = int_reg_array_25_2_imag;
        _zz_4485_ = int_reg_array_25_2_real;
      end
      6'b000011 : begin
        _zz_4484_ = int_reg_array_25_3_imag;
        _zz_4485_ = int_reg_array_25_3_real;
      end
      6'b000100 : begin
        _zz_4484_ = int_reg_array_25_4_imag;
        _zz_4485_ = int_reg_array_25_4_real;
      end
      6'b000101 : begin
        _zz_4484_ = int_reg_array_25_5_imag;
        _zz_4485_ = int_reg_array_25_5_real;
      end
      6'b000110 : begin
        _zz_4484_ = int_reg_array_25_6_imag;
        _zz_4485_ = int_reg_array_25_6_real;
      end
      6'b000111 : begin
        _zz_4484_ = int_reg_array_25_7_imag;
        _zz_4485_ = int_reg_array_25_7_real;
      end
      6'b001000 : begin
        _zz_4484_ = int_reg_array_25_8_imag;
        _zz_4485_ = int_reg_array_25_8_real;
      end
      6'b001001 : begin
        _zz_4484_ = int_reg_array_25_9_imag;
        _zz_4485_ = int_reg_array_25_9_real;
      end
      6'b001010 : begin
        _zz_4484_ = int_reg_array_25_10_imag;
        _zz_4485_ = int_reg_array_25_10_real;
      end
      6'b001011 : begin
        _zz_4484_ = int_reg_array_25_11_imag;
        _zz_4485_ = int_reg_array_25_11_real;
      end
      6'b001100 : begin
        _zz_4484_ = int_reg_array_25_12_imag;
        _zz_4485_ = int_reg_array_25_12_real;
      end
      6'b001101 : begin
        _zz_4484_ = int_reg_array_25_13_imag;
        _zz_4485_ = int_reg_array_25_13_real;
      end
      6'b001110 : begin
        _zz_4484_ = int_reg_array_25_14_imag;
        _zz_4485_ = int_reg_array_25_14_real;
      end
      6'b001111 : begin
        _zz_4484_ = int_reg_array_25_15_imag;
        _zz_4485_ = int_reg_array_25_15_real;
      end
      6'b010000 : begin
        _zz_4484_ = int_reg_array_25_16_imag;
        _zz_4485_ = int_reg_array_25_16_real;
      end
      6'b010001 : begin
        _zz_4484_ = int_reg_array_25_17_imag;
        _zz_4485_ = int_reg_array_25_17_real;
      end
      6'b010010 : begin
        _zz_4484_ = int_reg_array_25_18_imag;
        _zz_4485_ = int_reg_array_25_18_real;
      end
      6'b010011 : begin
        _zz_4484_ = int_reg_array_25_19_imag;
        _zz_4485_ = int_reg_array_25_19_real;
      end
      6'b010100 : begin
        _zz_4484_ = int_reg_array_25_20_imag;
        _zz_4485_ = int_reg_array_25_20_real;
      end
      6'b010101 : begin
        _zz_4484_ = int_reg_array_25_21_imag;
        _zz_4485_ = int_reg_array_25_21_real;
      end
      6'b010110 : begin
        _zz_4484_ = int_reg_array_25_22_imag;
        _zz_4485_ = int_reg_array_25_22_real;
      end
      6'b010111 : begin
        _zz_4484_ = int_reg_array_25_23_imag;
        _zz_4485_ = int_reg_array_25_23_real;
      end
      6'b011000 : begin
        _zz_4484_ = int_reg_array_25_24_imag;
        _zz_4485_ = int_reg_array_25_24_real;
      end
      6'b011001 : begin
        _zz_4484_ = int_reg_array_25_25_imag;
        _zz_4485_ = int_reg_array_25_25_real;
      end
      6'b011010 : begin
        _zz_4484_ = int_reg_array_25_26_imag;
        _zz_4485_ = int_reg_array_25_26_real;
      end
      6'b011011 : begin
        _zz_4484_ = int_reg_array_25_27_imag;
        _zz_4485_ = int_reg_array_25_27_real;
      end
      6'b011100 : begin
        _zz_4484_ = int_reg_array_25_28_imag;
        _zz_4485_ = int_reg_array_25_28_real;
      end
      6'b011101 : begin
        _zz_4484_ = int_reg_array_25_29_imag;
        _zz_4485_ = int_reg_array_25_29_real;
      end
      6'b011110 : begin
        _zz_4484_ = int_reg_array_25_30_imag;
        _zz_4485_ = int_reg_array_25_30_real;
      end
      6'b011111 : begin
        _zz_4484_ = int_reg_array_25_31_imag;
        _zz_4485_ = int_reg_array_25_31_real;
      end
      6'b100000 : begin
        _zz_4484_ = int_reg_array_25_32_imag;
        _zz_4485_ = int_reg_array_25_32_real;
      end
      6'b100001 : begin
        _zz_4484_ = int_reg_array_25_33_imag;
        _zz_4485_ = int_reg_array_25_33_real;
      end
      6'b100010 : begin
        _zz_4484_ = int_reg_array_25_34_imag;
        _zz_4485_ = int_reg_array_25_34_real;
      end
      6'b100011 : begin
        _zz_4484_ = int_reg_array_25_35_imag;
        _zz_4485_ = int_reg_array_25_35_real;
      end
      6'b100100 : begin
        _zz_4484_ = int_reg_array_25_36_imag;
        _zz_4485_ = int_reg_array_25_36_real;
      end
      6'b100101 : begin
        _zz_4484_ = int_reg_array_25_37_imag;
        _zz_4485_ = int_reg_array_25_37_real;
      end
      6'b100110 : begin
        _zz_4484_ = int_reg_array_25_38_imag;
        _zz_4485_ = int_reg_array_25_38_real;
      end
      6'b100111 : begin
        _zz_4484_ = int_reg_array_25_39_imag;
        _zz_4485_ = int_reg_array_25_39_real;
      end
      6'b101000 : begin
        _zz_4484_ = int_reg_array_25_40_imag;
        _zz_4485_ = int_reg_array_25_40_real;
      end
      6'b101001 : begin
        _zz_4484_ = int_reg_array_25_41_imag;
        _zz_4485_ = int_reg_array_25_41_real;
      end
      6'b101010 : begin
        _zz_4484_ = int_reg_array_25_42_imag;
        _zz_4485_ = int_reg_array_25_42_real;
      end
      6'b101011 : begin
        _zz_4484_ = int_reg_array_25_43_imag;
        _zz_4485_ = int_reg_array_25_43_real;
      end
      6'b101100 : begin
        _zz_4484_ = int_reg_array_25_44_imag;
        _zz_4485_ = int_reg_array_25_44_real;
      end
      6'b101101 : begin
        _zz_4484_ = int_reg_array_25_45_imag;
        _zz_4485_ = int_reg_array_25_45_real;
      end
      6'b101110 : begin
        _zz_4484_ = int_reg_array_25_46_imag;
        _zz_4485_ = int_reg_array_25_46_real;
      end
      6'b101111 : begin
        _zz_4484_ = int_reg_array_25_47_imag;
        _zz_4485_ = int_reg_array_25_47_real;
      end
      6'b110000 : begin
        _zz_4484_ = int_reg_array_25_48_imag;
        _zz_4485_ = int_reg_array_25_48_real;
      end
      6'b110001 : begin
        _zz_4484_ = int_reg_array_25_49_imag;
        _zz_4485_ = int_reg_array_25_49_real;
      end
      6'b110010 : begin
        _zz_4484_ = int_reg_array_25_50_imag;
        _zz_4485_ = int_reg_array_25_50_real;
      end
      6'b110011 : begin
        _zz_4484_ = int_reg_array_25_51_imag;
        _zz_4485_ = int_reg_array_25_51_real;
      end
      6'b110100 : begin
        _zz_4484_ = int_reg_array_25_52_imag;
        _zz_4485_ = int_reg_array_25_52_real;
      end
      6'b110101 : begin
        _zz_4484_ = int_reg_array_25_53_imag;
        _zz_4485_ = int_reg_array_25_53_real;
      end
      6'b110110 : begin
        _zz_4484_ = int_reg_array_25_54_imag;
        _zz_4485_ = int_reg_array_25_54_real;
      end
      6'b110111 : begin
        _zz_4484_ = int_reg_array_25_55_imag;
        _zz_4485_ = int_reg_array_25_55_real;
      end
      6'b111000 : begin
        _zz_4484_ = int_reg_array_25_56_imag;
        _zz_4485_ = int_reg_array_25_56_real;
      end
      6'b111001 : begin
        _zz_4484_ = int_reg_array_25_57_imag;
        _zz_4485_ = int_reg_array_25_57_real;
      end
      6'b111010 : begin
        _zz_4484_ = int_reg_array_25_58_imag;
        _zz_4485_ = int_reg_array_25_58_real;
      end
      6'b111011 : begin
        _zz_4484_ = int_reg_array_25_59_imag;
        _zz_4485_ = int_reg_array_25_59_real;
      end
      6'b111100 : begin
        _zz_4484_ = int_reg_array_25_60_imag;
        _zz_4485_ = int_reg_array_25_60_real;
      end
      6'b111101 : begin
        _zz_4484_ = int_reg_array_25_61_imag;
        _zz_4485_ = int_reg_array_25_61_real;
      end
      6'b111110 : begin
        _zz_4484_ = int_reg_array_25_62_imag;
        _zz_4485_ = int_reg_array_25_62_real;
      end
      default : begin
        _zz_4484_ = int_reg_array_25_63_imag;
        _zz_4485_ = int_reg_array_25_63_real;
      end
    endcase
  end

  always @(*) begin
    case(_zz_1811_)
      6'b000000 : begin
        _zz_4486_ = int_reg_array_26_0_imag;
        _zz_4487_ = int_reg_array_26_0_real;
      end
      6'b000001 : begin
        _zz_4486_ = int_reg_array_26_1_imag;
        _zz_4487_ = int_reg_array_26_1_real;
      end
      6'b000010 : begin
        _zz_4486_ = int_reg_array_26_2_imag;
        _zz_4487_ = int_reg_array_26_2_real;
      end
      6'b000011 : begin
        _zz_4486_ = int_reg_array_26_3_imag;
        _zz_4487_ = int_reg_array_26_3_real;
      end
      6'b000100 : begin
        _zz_4486_ = int_reg_array_26_4_imag;
        _zz_4487_ = int_reg_array_26_4_real;
      end
      6'b000101 : begin
        _zz_4486_ = int_reg_array_26_5_imag;
        _zz_4487_ = int_reg_array_26_5_real;
      end
      6'b000110 : begin
        _zz_4486_ = int_reg_array_26_6_imag;
        _zz_4487_ = int_reg_array_26_6_real;
      end
      6'b000111 : begin
        _zz_4486_ = int_reg_array_26_7_imag;
        _zz_4487_ = int_reg_array_26_7_real;
      end
      6'b001000 : begin
        _zz_4486_ = int_reg_array_26_8_imag;
        _zz_4487_ = int_reg_array_26_8_real;
      end
      6'b001001 : begin
        _zz_4486_ = int_reg_array_26_9_imag;
        _zz_4487_ = int_reg_array_26_9_real;
      end
      6'b001010 : begin
        _zz_4486_ = int_reg_array_26_10_imag;
        _zz_4487_ = int_reg_array_26_10_real;
      end
      6'b001011 : begin
        _zz_4486_ = int_reg_array_26_11_imag;
        _zz_4487_ = int_reg_array_26_11_real;
      end
      6'b001100 : begin
        _zz_4486_ = int_reg_array_26_12_imag;
        _zz_4487_ = int_reg_array_26_12_real;
      end
      6'b001101 : begin
        _zz_4486_ = int_reg_array_26_13_imag;
        _zz_4487_ = int_reg_array_26_13_real;
      end
      6'b001110 : begin
        _zz_4486_ = int_reg_array_26_14_imag;
        _zz_4487_ = int_reg_array_26_14_real;
      end
      6'b001111 : begin
        _zz_4486_ = int_reg_array_26_15_imag;
        _zz_4487_ = int_reg_array_26_15_real;
      end
      6'b010000 : begin
        _zz_4486_ = int_reg_array_26_16_imag;
        _zz_4487_ = int_reg_array_26_16_real;
      end
      6'b010001 : begin
        _zz_4486_ = int_reg_array_26_17_imag;
        _zz_4487_ = int_reg_array_26_17_real;
      end
      6'b010010 : begin
        _zz_4486_ = int_reg_array_26_18_imag;
        _zz_4487_ = int_reg_array_26_18_real;
      end
      6'b010011 : begin
        _zz_4486_ = int_reg_array_26_19_imag;
        _zz_4487_ = int_reg_array_26_19_real;
      end
      6'b010100 : begin
        _zz_4486_ = int_reg_array_26_20_imag;
        _zz_4487_ = int_reg_array_26_20_real;
      end
      6'b010101 : begin
        _zz_4486_ = int_reg_array_26_21_imag;
        _zz_4487_ = int_reg_array_26_21_real;
      end
      6'b010110 : begin
        _zz_4486_ = int_reg_array_26_22_imag;
        _zz_4487_ = int_reg_array_26_22_real;
      end
      6'b010111 : begin
        _zz_4486_ = int_reg_array_26_23_imag;
        _zz_4487_ = int_reg_array_26_23_real;
      end
      6'b011000 : begin
        _zz_4486_ = int_reg_array_26_24_imag;
        _zz_4487_ = int_reg_array_26_24_real;
      end
      6'b011001 : begin
        _zz_4486_ = int_reg_array_26_25_imag;
        _zz_4487_ = int_reg_array_26_25_real;
      end
      6'b011010 : begin
        _zz_4486_ = int_reg_array_26_26_imag;
        _zz_4487_ = int_reg_array_26_26_real;
      end
      6'b011011 : begin
        _zz_4486_ = int_reg_array_26_27_imag;
        _zz_4487_ = int_reg_array_26_27_real;
      end
      6'b011100 : begin
        _zz_4486_ = int_reg_array_26_28_imag;
        _zz_4487_ = int_reg_array_26_28_real;
      end
      6'b011101 : begin
        _zz_4486_ = int_reg_array_26_29_imag;
        _zz_4487_ = int_reg_array_26_29_real;
      end
      6'b011110 : begin
        _zz_4486_ = int_reg_array_26_30_imag;
        _zz_4487_ = int_reg_array_26_30_real;
      end
      6'b011111 : begin
        _zz_4486_ = int_reg_array_26_31_imag;
        _zz_4487_ = int_reg_array_26_31_real;
      end
      6'b100000 : begin
        _zz_4486_ = int_reg_array_26_32_imag;
        _zz_4487_ = int_reg_array_26_32_real;
      end
      6'b100001 : begin
        _zz_4486_ = int_reg_array_26_33_imag;
        _zz_4487_ = int_reg_array_26_33_real;
      end
      6'b100010 : begin
        _zz_4486_ = int_reg_array_26_34_imag;
        _zz_4487_ = int_reg_array_26_34_real;
      end
      6'b100011 : begin
        _zz_4486_ = int_reg_array_26_35_imag;
        _zz_4487_ = int_reg_array_26_35_real;
      end
      6'b100100 : begin
        _zz_4486_ = int_reg_array_26_36_imag;
        _zz_4487_ = int_reg_array_26_36_real;
      end
      6'b100101 : begin
        _zz_4486_ = int_reg_array_26_37_imag;
        _zz_4487_ = int_reg_array_26_37_real;
      end
      6'b100110 : begin
        _zz_4486_ = int_reg_array_26_38_imag;
        _zz_4487_ = int_reg_array_26_38_real;
      end
      6'b100111 : begin
        _zz_4486_ = int_reg_array_26_39_imag;
        _zz_4487_ = int_reg_array_26_39_real;
      end
      6'b101000 : begin
        _zz_4486_ = int_reg_array_26_40_imag;
        _zz_4487_ = int_reg_array_26_40_real;
      end
      6'b101001 : begin
        _zz_4486_ = int_reg_array_26_41_imag;
        _zz_4487_ = int_reg_array_26_41_real;
      end
      6'b101010 : begin
        _zz_4486_ = int_reg_array_26_42_imag;
        _zz_4487_ = int_reg_array_26_42_real;
      end
      6'b101011 : begin
        _zz_4486_ = int_reg_array_26_43_imag;
        _zz_4487_ = int_reg_array_26_43_real;
      end
      6'b101100 : begin
        _zz_4486_ = int_reg_array_26_44_imag;
        _zz_4487_ = int_reg_array_26_44_real;
      end
      6'b101101 : begin
        _zz_4486_ = int_reg_array_26_45_imag;
        _zz_4487_ = int_reg_array_26_45_real;
      end
      6'b101110 : begin
        _zz_4486_ = int_reg_array_26_46_imag;
        _zz_4487_ = int_reg_array_26_46_real;
      end
      6'b101111 : begin
        _zz_4486_ = int_reg_array_26_47_imag;
        _zz_4487_ = int_reg_array_26_47_real;
      end
      6'b110000 : begin
        _zz_4486_ = int_reg_array_26_48_imag;
        _zz_4487_ = int_reg_array_26_48_real;
      end
      6'b110001 : begin
        _zz_4486_ = int_reg_array_26_49_imag;
        _zz_4487_ = int_reg_array_26_49_real;
      end
      6'b110010 : begin
        _zz_4486_ = int_reg_array_26_50_imag;
        _zz_4487_ = int_reg_array_26_50_real;
      end
      6'b110011 : begin
        _zz_4486_ = int_reg_array_26_51_imag;
        _zz_4487_ = int_reg_array_26_51_real;
      end
      6'b110100 : begin
        _zz_4486_ = int_reg_array_26_52_imag;
        _zz_4487_ = int_reg_array_26_52_real;
      end
      6'b110101 : begin
        _zz_4486_ = int_reg_array_26_53_imag;
        _zz_4487_ = int_reg_array_26_53_real;
      end
      6'b110110 : begin
        _zz_4486_ = int_reg_array_26_54_imag;
        _zz_4487_ = int_reg_array_26_54_real;
      end
      6'b110111 : begin
        _zz_4486_ = int_reg_array_26_55_imag;
        _zz_4487_ = int_reg_array_26_55_real;
      end
      6'b111000 : begin
        _zz_4486_ = int_reg_array_26_56_imag;
        _zz_4487_ = int_reg_array_26_56_real;
      end
      6'b111001 : begin
        _zz_4486_ = int_reg_array_26_57_imag;
        _zz_4487_ = int_reg_array_26_57_real;
      end
      6'b111010 : begin
        _zz_4486_ = int_reg_array_26_58_imag;
        _zz_4487_ = int_reg_array_26_58_real;
      end
      6'b111011 : begin
        _zz_4486_ = int_reg_array_26_59_imag;
        _zz_4487_ = int_reg_array_26_59_real;
      end
      6'b111100 : begin
        _zz_4486_ = int_reg_array_26_60_imag;
        _zz_4487_ = int_reg_array_26_60_real;
      end
      6'b111101 : begin
        _zz_4486_ = int_reg_array_26_61_imag;
        _zz_4487_ = int_reg_array_26_61_real;
      end
      6'b111110 : begin
        _zz_4486_ = int_reg_array_26_62_imag;
        _zz_4487_ = int_reg_array_26_62_real;
      end
      default : begin
        _zz_4486_ = int_reg_array_26_63_imag;
        _zz_4487_ = int_reg_array_26_63_real;
      end
    endcase
  end

  always @(*) begin
    case(_zz_1880_)
      6'b000000 : begin
        _zz_4488_ = int_reg_array_27_0_imag;
        _zz_4489_ = int_reg_array_27_0_real;
      end
      6'b000001 : begin
        _zz_4488_ = int_reg_array_27_1_imag;
        _zz_4489_ = int_reg_array_27_1_real;
      end
      6'b000010 : begin
        _zz_4488_ = int_reg_array_27_2_imag;
        _zz_4489_ = int_reg_array_27_2_real;
      end
      6'b000011 : begin
        _zz_4488_ = int_reg_array_27_3_imag;
        _zz_4489_ = int_reg_array_27_3_real;
      end
      6'b000100 : begin
        _zz_4488_ = int_reg_array_27_4_imag;
        _zz_4489_ = int_reg_array_27_4_real;
      end
      6'b000101 : begin
        _zz_4488_ = int_reg_array_27_5_imag;
        _zz_4489_ = int_reg_array_27_5_real;
      end
      6'b000110 : begin
        _zz_4488_ = int_reg_array_27_6_imag;
        _zz_4489_ = int_reg_array_27_6_real;
      end
      6'b000111 : begin
        _zz_4488_ = int_reg_array_27_7_imag;
        _zz_4489_ = int_reg_array_27_7_real;
      end
      6'b001000 : begin
        _zz_4488_ = int_reg_array_27_8_imag;
        _zz_4489_ = int_reg_array_27_8_real;
      end
      6'b001001 : begin
        _zz_4488_ = int_reg_array_27_9_imag;
        _zz_4489_ = int_reg_array_27_9_real;
      end
      6'b001010 : begin
        _zz_4488_ = int_reg_array_27_10_imag;
        _zz_4489_ = int_reg_array_27_10_real;
      end
      6'b001011 : begin
        _zz_4488_ = int_reg_array_27_11_imag;
        _zz_4489_ = int_reg_array_27_11_real;
      end
      6'b001100 : begin
        _zz_4488_ = int_reg_array_27_12_imag;
        _zz_4489_ = int_reg_array_27_12_real;
      end
      6'b001101 : begin
        _zz_4488_ = int_reg_array_27_13_imag;
        _zz_4489_ = int_reg_array_27_13_real;
      end
      6'b001110 : begin
        _zz_4488_ = int_reg_array_27_14_imag;
        _zz_4489_ = int_reg_array_27_14_real;
      end
      6'b001111 : begin
        _zz_4488_ = int_reg_array_27_15_imag;
        _zz_4489_ = int_reg_array_27_15_real;
      end
      6'b010000 : begin
        _zz_4488_ = int_reg_array_27_16_imag;
        _zz_4489_ = int_reg_array_27_16_real;
      end
      6'b010001 : begin
        _zz_4488_ = int_reg_array_27_17_imag;
        _zz_4489_ = int_reg_array_27_17_real;
      end
      6'b010010 : begin
        _zz_4488_ = int_reg_array_27_18_imag;
        _zz_4489_ = int_reg_array_27_18_real;
      end
      6'b010011 : begin
        _zz_4488_ = int_reg_array_27_19_imag;
        _zz_4489_ = int_reg_array_27_19_real;
      end
      6'b010100 : begin
        _zz_4488_ = int_reg_array_27_20_imag;
        _zz_4489_ = int_reg_array_27_20_real;
      end
      6'b010101 : begin
        _zz_4488_ = int_reg_array_27_21_imag;
        _zz_4489_ = int_reg_array_27_21_real;
      end
      6'b010110 : begin
        _zz_4488_ = int_reg_array_27_22_imag;
        _zz_4489_ = int_reg_array_27_22_real;
      end
      6'b010111 : begin
        _zz_4488_ = int_reg_array_27_23_imag;
        _zz_4489_ = int_reg_array_27_23_real;
      end
      6'b011000 : begin
        _zz_4488_ = int_reg_array_27_24_imag;
        _zz_4489_ = int_reg_array_27_24_real;
      end
      6'b011001 : begin
        _zz_4488_ = int_reg_array_27_25_imag;
        _zz_4489_ = int_reg_array_27_25_real;
      end
      6'b011010 : begin
        _zz_4488_ = int_reg_array_27_26_imag;
        _zz_4489_ = int_reg_array_27_26_real;
      end
      6'b011011 : begin
        _zz_4488_ = int_reg_array_27_27_imag;
        _zz_4489_ = int_reg_array_27_27_real;
      end
      6'b011100 : begin
        _zz_4488_ = int_reg_array_27_28_imag;
        _zz_4489_ = int_reg_array_27_28_real;
      end
      6'b011101 : begin
        _zz_4488_ = int_reg_array_27_29_imag;
        _zz_4489_ = int_reg_array_27_29_real;
      end
      6'b011110 : begin
        _zz_4488_ = int_reg_array_27_30_imag;
        _zz_4489_ = int_reg_array_27_30_real;
      end
      6'b011111 : begin
        _zz_4488_ = int_reg_array_27_31_imag;
        _zz_4489_ = int_reg_array_27_31_real;
      end
      6'b100000 : begin
        _zz_4488_ = int_reg_array_27_32_imag;
        _zz_4489_ = int_reg_array_27_32_real;
      end
      6'b100001 : begin
        _zz_4488_ = int_reg_array_27_33_imag;
        _zz_4489_ = int_reg_array_27_33_real;
      end
      6'b100010 : begin
        _zz_4488_ = int_reg_array_27_34_imag;
        _zz_4489_ = int_reg_array_27_34_real;
      end
      6'b100011 : begin
        _zz_4488_ = int_reg_array_27_35_imag;
        _zz_4489_ = int_reg_array_27_35_real;
      end
      6'b100100 : begin
        _zz_4488_ = int_reg_array_27_36_imag;
        _zz_4489_ = int_reg_array_27_36_real;
      end
      6'b100101 : begin
        _zz_4488_ = int_reg_array_27_37_imag;
        _zz_4489_ = int_reg_array_27_37_real;
      end
      6'b100110 : begin
        _zz_4488_ = int_reg_array_27_38_imag;
        _zz_4489_ = int_reg_array_27_38_real;
      end
      6'b100111 : begin
        _zz_4488_ = int_reg_array_27_39_imag;
        _zz_4489_ = int_reg_array_27_39_real;
      end
      6'b101000 : begin
        _zz_4488_ = int_reg_array_27_40_imag;
        _zz_4489_ = int_reg_array_27_40_real;
      end
      6'b101001 : begin
        _zz_4488_ = int_reg_array_27_41_imag;
        _zz_4489_ = int_reg_array_27_41_real;
      end
      6'b101010 : begin
        _zz_4488_ = int_reg_array_27_42_imag;
        _zz_4489_ = int_reg_array_27_42_real;
      end
      6'b101011 : begin
        _zz_4488_ = int_reg_array_27_43_imag;
        _zz_4489_ = int_reg_array_27_43_real;
      end
      6'b101100 : begin
        _zz_4488_ = int_reg_array_27_44_imag;
        _zz_4489_ = int_reg_array_27_44_real;
      end
      6'b101101 : begin
        _zz_4488_ = int_reg_array_27_45_imag;
        _zz_4489_ = int_reg_array_27_45_real;
      end
      6'b101110 : begin
        _zz_4488_ = int_reg_array_27_46_imag;
        _zz_4489_ = int_reg_array_27_46_real;
      end
      6'b101111 : begin
        _zz_4488_ = int_reg_array_27_47_imag;
        _zz_4489_ = int_reg_array_27_47_real;
      end
      6'b110000 : begin
        _zz_4488_ = int_reg_array_27_48_imag;
        _zz_4489_ = int_reg_array_27_48_real;
      end
      6'b110001 : begin
        _zz_4488_ = int_reg_array_27_49_imag;
        _zz_4489_ = int_reg_array_27_49_real;
      end
      6'b110010 : begin
        _zz_4488_ = int_reg_array_27_50_imag;
        _zz_4489_ = int_reg_array_27_50_real;
      end
      6'b110011 : begin
        _zz_4488_ = int_reg_array_27_51_imag;
        _zz_4489_ = int_reg_array_27_51_real;
      end
      6'b110100 : begin
        _zz_4488_ = int_reg_array_27_52_imag;
        _zz_4489_ = int_reg_array_27_52_real;
      end
      6'b110101 : begin
        _zz_4488_ = int_reg_array_27_53_imag;
        _zz_4489_ = int_reg_array_27_53_real;
      end
      6'b110110 : begin
        _zz_4488_ = int_reg_array_27_54_imag;
        _zz_4489_ = int_reg_array_27_54_real;
      end
      6'b110111 : begin
        _zz_4488_ = int_reg_array_27_55_imag;
        _zz_4489_ = int_reg_array_27_55_real;
      end
      6'b111000 : begin
        _zz_4488_ = int_reg_array_27_56_imag;
        _zz_4489_ = int_reg_array_27_56_real;
      end
      6'b111001 : begin
        _zz_4488_ = int_reg_array_27_57_imag;
        _zz_4489_ = int_reg_array_27_57_real;
      end
      6'b111010 : begin
        _zz_4488_ = int_reg_array_27_58_imag;
        _zz_4489_ = int_reg_array_27_58_real;
      end
      6'b111011 : begin
        _zz_4488_ = int_reg_array_27_59_imag;
        _zz_4489_ = int_reg_array_27_59_real;
      end
      6'b111100 : begin
        _zz_4488_ = int_reg_array_27_60_imag;
        _zz_4489_ = int_reg_array_27_60_real;
      end
      6'b111101 : begin
        _zz_4488_ = int_reg_array_27_61_imag;
        _zz_4489_ = int_reg_array_27_61_real;
      end
      6'b111110 : begin
        _zz_4488_ = int_reg_array_27_62_imag;
        _zz_4489_ = int_reg_array_27_62_real;
      end
      default : begin
        _zz_4488_ = int_reg_array_27_63_imag;
        _zz_4489_ = int_reg_array_27_63_real;
      end
    endcase
  end

  always @(*) begin
    case(_zz_1949_)
      6'b000000 : begin
        _zz_4490_ = int_reg_array_28_0_imag;
        _zz_4491_ = int_reg_array_28_0_real;
      end
      6'b000001 : begin
        _zz_4490_ = int_reg_array_28_1_imag;
        _zz_4491_ = int_reg_array_28_1_real;
      end
      6'b000010 : begin
        _zz_4490_ = int_reg_array_28_2_imag;
        _zz_4491_ = int_reg_array_28_2_real;
      end
      6'b000011 : begin
        _zz_4490_ = int_reg_array_28_3_imag;
        _zz_4491_ = int_reg_array_28_3_real;
      end
      6'b000100 : begin
        _zz_4490_ = int_reg_array_28_4_imag;
        _zz_4491_ = int_reg_array_28_4_real;
      end
      6'b000101 : begin
        _zz_4490_ = int_reg_array_28_5_imag;
        _zz_4491_ = int_reg_array_28_5_real;
      end
      6'b000110 : begin
        _zz_4490_ = int_reg_array_28_6_imag;
        _zz_4491_ = int_reg_array_28_6_real;
      end
      6'b000111 : begin
        _zz_4490_ = int_reg_array_28_7_imag;
        _zz_4491_ = int_reg_array_28_7_real;
      end
      6'b001000 : begin
        _zz_4490_ = int_reg_array_28_8_imag;
        _zz_4491_ = int_reg_array_28_8_real;
      end
      6'b001001 : begin
        _zz_4490_ = int_reg_array_28_9_imag;
        _zz_4491_ = int_reg_array_28_9_real;
      end
      6'b001010 : begin
        _zz_4490_ = int_reg_array_28_10_imag;
        _zz_4491_ = int_reg_array_28_10_real;
      end
      6'b001011 : begin
        _zz_4490_ = int_reg_array_28_11_imag;
        _zz_4491_ = int_reg_array_28_11_real;
      end
      6'b001100 : begin
        _zz_4490_ = int_reg_array_28_12_imag;
        _zz_4491_ = int_reg_array_28_12_real;
      end
      6'b001101 : begin
        _zz_4490_ = int_reg_array_28_13_imag;
        _zz_4491_ = int_reg_array_28_13_real;
      end
      6'b001110 : begin
        _zz_4490_ = int_reg_array_28_14_imag;
        _zz_4491_ = int_reg_array_28_14_real;
      end
      6'b001111 : begin
        _zz_4490_ = int_reg_array_28_15_imag;
        _zz_4491_ = int_reg_array_28_15_real;
      end
      6'b010000 : begin
        _zz_4490_ = int_reg_array_28_16_imag;
        _zz_4491_ = int_reg_array_28_16_real;
      end
      6'b010001 : begin
        _zz_4490_ = int_reg_array_28_17_imag;
        _zz_4491_ = int_reg_array_28_17_real;
      end
      6'b010010 : begin
        _zz_4490_ = int_reg_array_28_18_imag;
        _zz_4491_ = int_reg_array_28_18_real;
      end
      6'b010011 : begin
        _zz_4490_ = int_reg_array_28_19_imag;
        _zz_4491_ = int_reg_array_28_19_real;
      end
      6'b010100 : begin
        _zz_4490_ = int_reg_array_28_20_imag;
        _zz_4491_ = int_reg_array_28_20_real;
      end
      6'b010101 : begin
        _zz_4490_ = int_reg_array_28_21_imag;
        _zz_4491_ = int_reg_array_28_21_real;
      end
      6'b010110 : begin
        _zz_4490_ = int_reg_array_28_22_imag;
        _zz_4491_ = int_reg_array_28_22_real;
      end
      6'b010111 : begin
        _zz_4490_ = int_reg_array_28_23_imag;
        _zz_4491_ = int_reg_array_28_23_real;
      end
      6'b011000 : begin
        _zz_4490_ = int_reg_array_28_24_imag;
        _zz_4491_ = int_reg_array_28_24_real;
      end
      6'b011001 : begin
        _zz_4490_ = int_reg_array_28_25_imag;
        _zz_4491_ = int_reg_array_28_25_real;
      end
      6'b011010 : begin
        _zz_4490_ = int_reg_array_28_26_imag;
        _zz_4491_ = int_reg_array_28_26_real;
      end
      6'b011011 : begin
        _zz_4490_ = int_reg_array_28_27_imag;
        _zz_4491_ = int_reg_array_28_27_real;
      end
      6'b011100 : begin
        _zz_4490_ = int_reg_array_28_28_imag;
        _zz_4491_ = int_reg_array_28_28_real;
      end
      6'b011101 : begin
        _zz_4490_ = int_reg_array_28_29_imag;
        _zz_4491_ = int_reg_array_28_29_real;
      end
      6'b011110 : begin
        _zz_4490_ = int_reg_array_28_30_imag;
        _zz_4491_ = int_reg_array_28_30_real;
      end
      6'b011111 : begin
        _zz_4490_ = int_reg_array_28_31_imag;
        _zz_4491_ = int_reg_array_28_31_real;
      end
      6'b100000 : begin
        _zz_4490_ = int_reg_array_28_32_imag;
        _zz_4491_ = int_reg_array_28_32_real;
      end
      6'b100001 : begin
        _zz_4490_ = int_reg_array_28_33_imag;
        _zz_4491_ = int_reg_array_28_33_real;
      end
      6'b100010 : begin
        _zz_4490_ = int_reg_array_28_34_imag;
        _zz_4491_ = int_reg_array_28_34_real;
      end
      6'b100011 : begin
        _zz_4490_ = int_reg_array_28_35_imag;
        _zz_4491_ = int_reg_array_28_35_real;
      end
      6'b100100 : begin
        _zz_4490_ = int_reg_array_28_36_imag;
        _zz_4491_ = int_reg_array_28_36_real;
      end
      6'b100101 : begin
        _zz_4490_ = int_reg_array_28_37_imag;
        _zz_4491_ = int_reg_array_28_37_real;
      end
      6'b100110 : begin
        _zz_4490_ = int_reg_array_28_38_imag;
        _zz_4491_ = int_reg_array_28_38_real;
      end
      6'b100111 : begin
        _zz_4490_ = int_reg_array_28_39_imag;
        _zz_4491_ = int_reg_array_28_39_real;
      end
      6'b101000 : begin
        _zz_4490_ = int_reg_array_28_40_imag;
        _zz_4491_ = int_reg_array_28_40_real;
      end
      6'b101001 : begin
        _zz_4490_ = int_reg_array_28_41_imag;
        _zz_4491_ = int_reg_array_28_41_real;
      end
      6'b101010 : begin
        _zz_4490_ = int_reg_array_28_42_imag;
        _zz_4491_ = int_reg_array_28_42_real;
      end
      6'b101011 : begin
        _zz_4490_ = int_reg_array_28_43_imag;
        _zz_4491_ = int_reg_array_28_43_real;
      end
      6'b101100 : begin
        _zz_4490_ = int_reg_array_28_44_imag;
        _zz_4491_ = int_reg_array_28_44_real;
      end
      6'b101101 : begin
        _zz_4490_ = int_reg_array_28_45_imag;
        _zz_4491_ = int_reg_array_28_45_real;
      end
      6'b101110 : begin
        _zz_4490_ = int_reg_array_28_46_imag;
        _zz_4491_ = int_reg_array_28_46_real;
      end
      6'b101111 : begin
        _zz_4490_ = int_reg_array_28_47_imag;
        _zz_4491_ = int_reg_array_28_47_real;
      end
      6'b110000 : begin
        _zz_4490_ = int_reg_array_28_48_imag;
        _zz_4491_ = int_reg_array_28_48_real;
      end
      6'b110001 : begin
        _zz_4490_ = int_reg_array_28_49_imag;
        _zz_4491_ = int_reg_array_28_49_real;
      end
      6'b110010 : begin
        _zz_4490_ = int_reg_array_28_50_imag;
        _zz_4491_ = int_reg_array_28_50_real;
      end
      6'b110011 : begin
        _zz_4490_ = int_reg_array_28_51_imag;
        _zz_4491_ = int_reg_array_28_51_real;
      end
      6'b110100 : begin
        _zz_4490_ = int_reg_array_28_52_imag;
        _zz_4491_ = int_reg_array_28_52_real;
      end
      6'b110101 : begin
        _zz_4490_ = int_reg_array_28_53_imag;
        _zz_4491_ = int_reg_array_28_53_real;
      end
      6'b110110 : begin
        _zz_4490_ = int_reg_array_28_54_imag;
        _zz_4491_ = int_reg_array_28_54_real;
      end
      6'b110111 : begin
        _zz_4490_ = int_reg_array_28_55_imag;
        _zz_4491_ = int_reg_array_28_55_real;
      end
      6'b111000 : begin
        _zz_4490_ = int_reg_array_28_56_imag;
        _zz_4491_ = int_reg_array_28_56_real;
      end
      6'b111001 : begin
        _zz_4490_ = int_reg_array_28_57_imag;
        _zz_4491_ = int_reg_array_28_57_real;
      end
      6'b111010 : begin
        _zz_4490_ = int_reg_array_28_58_imag;
        _zz_4491_ = int_reg_array_28_58_real;
      end
      6'b111011 : begin
        _zz_4490_ = int_reg_array_28_59_imag;
        _zz_4491_ = int_reg_array_28_59_real;
      end
      6'b111100 : begin
        _zz_4490_ = int_reg_array_28_60_imag;
        _zz_4491_ = int_reg_array_28_60_real;
      end
      6'b111101 : begin
        _zz_4490_ = int_reg_array_28_61_imag;
        _zz_4491_ = int_reg_array_28_61_real;
      end
      6'b111110 : begin
        _zz_4490_ = int_reg_array_28_62_imag;
        _zz_4491_ = int_reg_array_28_62_real;
      end
      default : begin
        _zz_4490_ = int_reg_array_28_63_imag;
        _zz_4491_ = int_reg_array_28_63_real;
      end
    endcase
  end

  always @(*) begin
    case(_zz_2018_)
      6'b000000 : begin
        _zz_4492_ = int_reg_array_29_0_imag;
        _zz_4493_ = int_reg_array_29_0_real;
      end
      6'b000001 : begin
        _zz_4492_ = int_reg_array_29_1_imag;
        _zz_4493_ = int_reg_array_29_1_real;
      end
      6'b000010 : begin
        _zz_4492_ = int_reg_array_29_2_imag;
        _zz_4493_ = int_reg_array_29_2_real;
      end
      6'b000011 : begin
        _zz_4492_ = int_reg_array_29_3_imag;
        _zz_4493_ = int_reg_array_29_3_real;
      end
      6'b000100 : begin
        _zz_4492_ = int_reg_array_29_4_imag;
        _zz_4493_ = int_reg_array_29_4_real;
      end
      6'b000101 : begin
        _zz_4492_ = int_reg_array_29_5_imag;
        _zz_4493_ = int_reg_array_29_5_real;
      end
      6'b000110 : begin
        _zz_4492_ = int_reg_array_29_6_imag;
        _zz_4493_ = int_reg_array_29_6_real;
      end
      6'b000111 : begin
        _zz_4492_ = int_reg_array_29_7_imag;
        _zz_4493_ = int_reg_array_29_7_real;
      end
      6'b001000 : begin
        _zz_4492_ = int_reg_array_29_8_imag;
        _zz_4493_ = int_reg_array_29_8_real;
      end
      6'b001001 : begin
        _zz_4492_ = int_reg_array_29_9_imag;
        _zz_4493_ = int_reg_array_29_9_real;
      end
      6'b001010 : begin
        _zz_4492_ = int_reg_array_29_10_imag;
        _zz_4493_ = int_reg_array_29_10_real;
      end
      6'b001011 : begin
        _zz_4492_ = int_reg_array_29_11_imag;
        _zz_4493_ = int_reg_array_29_11_real;
      end
      6'b001100 : begin
        _zz_4492_ = int_reg_array_29_12_imag;
        _zz_4493_ = int_reg_array_29_12_real;
      end
      6'b001101 : begin
        _zz_4492_ = int_reg_array_29_13_imag;
        _zz_4493_ = int_reg_array_29_13_real;
      end
      6'b001110 : begin
        _zz_4492_ = int_reg_array_29_14_imag;
        _zz_4493_ = int_reg_array_29_14_real;
      end
      6'b001111 : begin
        _zz_4492_ = int_reg_array_29_15_imag;
        _zz_4493_ = int_reg_array_29_15_real;
      end
      6'b010000 : begin
        _zz_4492_ = int_reg_array_29_16_imag;
        _zz_4493_ = int_reg_array_29_16_real;
      end
      6'b010001 : begin
        _zz_4492_ = int_reg_array_29_17_imag;
        _zz_4493_ = int_reg_array_29_17_real;
      end
      6'b010010 : begin
        _zz_4492_ = int_reg_array_29_18_imag;
        _zz_4493_ = int_reg_array_29_18_real;
      end
      6'b010011 : begin
        _zz_4492_ = int_reg_array_29_19_imag;
        _zz_4493_ = int_reg_array_29_19_real;
      end
      6'b010100 : begin
        _zz_4492_ = int_reg_array_29_20_imag;
        _zz_4493_ = int_reg_array_29_20_real;
      end
      6'b010101 : begin
        _zz_4492_ = int_reg_array_29_21_imag;
        _zz_4493_ = int_reg_array_29_21_real;
      end
      6'b010110 : begin
        _zz_4492_ = int_reg_array_29_22_imag;
        _zz_4493_ = int_reg_array_29_22_real;
      end
      6'b010111 : begin
        _zz_4492_ = int_reg_array_29_23_imag;
        _zz_4493_ = int_reg_array_29_23_real;
      end
      6'b011000 : begin
        _zz_4492_ = int_reg_array_29_24_imag;
        _zz_4493_ = int_reg_array_29_24_real;
      end
      6'b011001 : begin
        _zz_4492_ = int_reg_array_29_25_imag;
        _zz_4493_ = int_reg_array_29_25_real;
      end
      6'b011010 : begin
        _zz_4492_ = int_reg_array_29_26_imag;
        _zz_4493_ = int_reg_array_29_26_real;
      end
      6'b011011 : begin
        _zz_4492_ = int_reg_array_29_27_imag;
        _zz_4493_ = int_reg_array_29_27_real;
      end
      6'b011100 : begin
        _zz_4492_ = int_reg_array_29_28_imag;
        _zz_4493_ = int_reg_array_29_28_real;
      end
      6'b011101 : begin
        _zz_4492_ = int_reg_array_29_29_imag;
        _zz_4493_ = int_reg_array_29_29_real;
      end
      6'b011110 : begin
        _zz_4492_ = int_reg_array_29_30_imag;
        _zz_4493_ = int_reg_array_29_30_real;
      end
      6'b011111 : begin
        _zz_4492_ = int_reg_array_29_31_imag;
        _zz_4493_ = int_reg_array_29_31_real;
      end
      6'b100000 : begin
        _zz_4492_ = int_reg_array_29_32_imag;
        _zz_4493_ = int_reg_array_29_32_real;
      end
      6'b100001 : begin
        _zz_4492_ = int_reg_array_29_33_imag;
        _zz_4493_ = int_reg_array_29_33_real;
      end
      6'b100010 : begin
        _zz_4492_ = int_reg_array_29_34_imag;
        _zz_4493_ = int_reg_array_29_34_real;
      end
      6'b100011 : begin
        _zz_4492_ = int_reg_array_29_35_imag;
        _zz_4493_ = int_reg_array_29_35_real;
      end
      6'b100100 : begin
        _zz_4492_ = int_reg_array_29_36_imag;
        _zz_4493_ = int_reg_array_29_36_real;
      end
      6'b100101 : begin
        _zz_4492_ = int_reg_array_29_37_imag;
        _zz_4493_ = int_reg_array_29_37_real;
      end
      6'b100110 : begin
        _zz_4492_ = int_reg_array_29_38_imag;
        _zz_4493_ = int_reg_array_29_38_real;
      end
      6'b100111 : begin
        _zz_4492_ = int_reg_array_29_39_imag;
        _zz_4493_ = int_reg_array_29_39_real;
      end
      6'b101000 : begin
        _zz_4492_ = int_reg_array_29_40_imag;
        _zz_4493_ = int_reg_array_29_40_real;
      end
      6'b101001 : begin
        _zz_4492_ = int_reg_array_29_41_imag;
        _zz_4493_ = int_reg_array_29_41_real;
      end
      6'b101010 : begin
        _zz_4492_ = int_reg_array_29_42_imag;
        _zz_4493_ = int_reg_array_29_42_real;
      end
      6'b101011 : begin
        _zz_4492_ = int_reg_array_29_43_imag;
        _zz_4493_ = int_reg_array_29_43_real;
      end
      6'b101100 : begin
        _zz_4492_ = int_reg_array_29_44_imag;
        _zz_4493_ = int_reg_array_29_44_real;
      end
      6'b101101 : begin
        _zz_4492_ = int_reg_array_29_45_imag;
        _zz_4493_ = int_reg_array_29_45_real;
      end
      6'b101110 : begin
        _zz_4492_ = int_reg_array_29_46_imag;
        _zz_4493_ = int_reg_array_29_46_real;
      end
      6'b101111 : begin
        _zz_4492_ = int_reg_array_29_47_imag;
        _zz_4493_ = int_reg_array_29_47_real;
      end
      6'b110000 : begin
        _zz_4492_ = int_reg_array_29_48_imag;
        _zz_4493_ = int_reg_array_29_48_real;
      end
      6'b110001 : begin
        _zz_4492_ = int_reg_array_29_49_imag;
        _zz_4493_ = int_reg_array_29_49_real;
      end
      6'b110010 : begin
        _zz_4492_ = int_reg_array_29_50_imag;
        _zz_4493_ = int_reg_array_29_50_real;
      end
      6'b110011 : begin
        _zz_4492_ = int_reg_array_29_51_imag;
        _zz_4493_ = int_reg_array_29_51_real;
      end
      6'b110100 : begin
        _zz_4492_ = int_reg_array_29_52_imag;
        _zz_4493_ = int_reg_array_29_52_real;
      end
      6'b110101 : begin
        _zz_4492_ = int_reg_array_29_53_imag;
        _zz_4493_ = int_reg_array_29_53_real;
      end
      6'b110110 : begin
        _zz_4492_ = int_reg_array_29_54_imag;
        _zz_4493_ = int_reg_array_29_54_real;
      end
      6'b110111 : begin
        _zz_4492_ = int_reg_array_29_55_imag;
        _zz_4493_ = int_reg_array_29_55_real;
      end
      6'b111000 : begin
        _zz_4492_ = int_reg_array_29_56_imag;
        _zz_4493_ = int_reg_array_29_56_real;
      end
      6'b111001 : begin
        _zz_4492_ = int_reg_array_29_57_imag;
        _zz_4493_ = int_reg_array_29_57_real;
      end
      6'b111010 : begin
        _zz_4492_ = int_reg_array_29_58_imag;
        _zz_4493_ = int_reg_array_29_58_real;
      end
      6'b111011 : begin
        _zz_4492_ = int_reg_array_29_59_imag;
        _zz_4493_ = int_reg_array_29_59_real;
      end
      6'b111100 : begin
        _zz_4492_ = int_reg_array_29_60_imag;
        _zz_4493_ = int_reg_array_29_60_real;
      end
      6'b111101 : begin
        _zz_4492_ = int_reg_array_29_61_imag;
        _zz_4493_ = int_reg_array_29_61_real;
      end
      6'b111110 : begin
        _zz_4492_ = int_reg_array_29_62_imag;
        _zz_4493_ = int_reg_array_29_62_real;
      end
      default : begin
        _zz_4492_ = int_reg_array_29_63_imag;
        _zz_4493_ = int_reg_array_29_63_real;
      end
    endcase
  end

  always @(*) begin
    case(_zz_2087_)
      6'b000000 : begin
        _zz_4494_ = int_reg_array_30_0_imag;
        _zz_4495_ = int_reg_array_30_0_real;
      end
      6'b000001 : begin
        _zz_4494_ = int_reg_array_30_1_imag;
        _zz_4495_ = int_reg_array_30_1_real;
      end
      6'b000010 : begin
        _zz_4494_ = int_reg_array_30_2_imag;
        _zz_4495_ = int_reg_array_30_2_real;
      end
      6'b000011 : begin
        _zz_4494_ = int_reg_array_30_3_imag;
        _zz_4495_ = int_reg_array_30_3_real;
      end
      6'b000100 : begin
        _zz_4494_ = int_reg_array_30_4_imag;
        _zz_4495_ = int_reg_array_30_4_real;
      end
      6'b000101 : begin
        _zz_4494_ = int_reg_array_30_5_imag;
        _zz_4495_ = int_reg_array_30_5_real;
      end
      6'b000110 : begin
        _zz_4494_ = int_reg_array_30_6_imag;
        _zz_4495_ = int_reg_array_30_6_real;
      end
      6'b000111 : begin
        _zz_4494_ = int_reg_array_30_7_imag;
        _zz_4495_ = int_reg_array_30_7_real;
      end
      6'b001000 : begin
        _zz_4494_ = int_reg_array_30_8_imag;
        _zz_4495_ = int_reg_array_30_8_real;
      end
      6'b001001 : begin
        _zz_4494_ = int_reg_array_30_9_imag;
        _zz_4495_ = int_reg_array_30_9_real;
      end
      6'b001010 : begin
        _zz_4494_ = int_reg_array_30_10_imag;
        _zz_4495_ = int_reg_array_30_10_real;
      end
      6'b001011 : begin
        _zz_4494_ = int_reg_array_30_11_imag;
        _zz_4495_ = int_reg_array_30_11_real;
      end
      6'b001100 : begin
        _zz_4494_ = int_reg_array_30_12_imag;
        _zz_4495_ = int_reg_array_30_12_real;
      end
      6'b001101 : begin
        _zz_4494_ = int_reg_array_30_13_imag;
        _zz_4495_ = int_reg_array_30_13_real;
      end
      6'b001110 : begin
        _zz_4494_ = int_reg_array_30_14_imag;
        _zz_4495_ = int_reg_array_30_14_real;
      end
      6'b001111 : begin
        _zz_4494_ = int_reg_array_30_15_imag;
        _zz_4495_ = int_reg_array_30_15_real;
      end
      6'b010000 : begin
        _zz_4494_ = int_reg_array_30_16_imag;
        _zz_4495_ = int_reg_array_30_16_real;
      end
      6'b010001 : begin
        _zz_4494_ = int_reg_array_30_17_imag;
        _zz_4495_ = int_reg_array_30_17_real;
      end
      6'b010010 : begin
        _zz_4494_ = int_reg_array_30_18_imag;
        _zz_4495_ = int_reg_array_30_18_real;
      end
      6'b010011 : begin
        _zz_4494_ = int_reg_array_30_19_imag;
        _zz_4495_ = int_reg_array_30_19_real;
      end
      6'b010100 : begin
        _zz_4494_ = int_reg_array_30_20_imag;
        _zz_4495_ = int_reg_array_30_20_real;
      end
      6'b010101 : begin
        _zz_4494_ = int_reg_array_30_21_imag;
        _zz_4495_ = int_reg_array_30_21_real;
      end
      6'b010110 : begin
        _zz_4494_ = int_reg_array_30_22_imag;
        _zz_4495_ = int_reg_array_30_22_real;
      end
      6'b010111 : begin
        _zz_4494_ = int_reg_array_30_23_imag;
        _zz_4495_ = int_reg_array_30_23_real;
      end
      6'b011000 : begin
        _zz_4494_ = int_reg_array_30_24_imag;
        _zz_4495_ = int_reg_array_30_24_real;
      end
      6'b011001 : begin
        _zz_4494_ = int_reg_array_30_25_imag;
        _zz_4495_ = int_reg_array_30_25_real;
      end
      6'b011010 : begin
        _zz_4494_ = int_reg_array_30_26_imag;
        _zz_4495_ = int_reg_array_30_26_real;
      end
      6'b011011 : begin
        _zz_4494_ = int_reg_array_30_27_imag;
        _zz_4495_ = int_reg_array_30_27_real;
      end
      6'b011100 : begin
        _zz_4494_ = int_reg_array_30_28_imag;
        _zz_4495_ = int_reg_array_30_28_real;
      end
      6'b011101 : begin
        _zz_4494_ = int_reg_array_30_29_imag;
        _zz_4495_ = int_reg_array_30_29_real;
      end
      6'b011110 : begin
        _zz_4494_ = int_reg_array_30_30_imag;
        _zz_4495_ = int_reg_array_30_30_real;
      end
      6'b011111 : begin
        _zz_4494_ = int_reg_array_30_31_imag;
        _zz_4495_ = int_reg_array_30_31_real;
      end
      6'b100000 : begin
        _zz_4494_ = int_reg_array_30_32_imag;
        _zz_4495_ = int_reg_array_30_32_real;
      end
      6'b100001 : begin
        _zz_4494_ = int_reg_array_30_33_imag;
        _zz_4495_ = int_reg_array_30_33_real;
      end
      6'b100010 : begin
        _zz_4494_ = int_reg_array_30_34_imag;
        _zz_4495_ = int_reg_array_30_34_real;
      end
      6'b100011 : begin
        _zz_4494_ = int_reg_array_30_35_imag;
        _zz_4495_ = int_reg_array_30_35_real;
      end
      6'b100100 : begin
        _zz_4494_ = int_reg_array_30_36_imag;
        _zz_4495_ = int_reg_array_30_36_real;
      end
      6'b100101 : begin
        _zz_4494_ = int_reg_array_30_37_imag;
        _zz_4495_ = int_reg_array_30_37_real;
      end
      6'b100110 : begin
        _zz_4494_ = int_reg_array_30_38_imag;
        _zz_4495_ = int_reg_array_30_38_real;
      end
      6'b100111 : begin
        _zz_4494_ = int_reg_array_30_39_imag;
        _zz_4495_ = int_reg_array_30_39_real;
      end
      6'b101000 : begin
        _zz_4494_ = int_reg_array_30_40_imag;
        _zz_4495_ = int_reg_array_30_40_real;
      end
      6'b101001 : begin
        _zz_4494_ = int_reg_array_30_41_imag;
        _zz_4495_ = int_reg_array_30_41_real;
      end
      6'b101010 : begin
        _zz_4494_ = int_reg_array_30_42_imag;
        _zz_4495_ = int_reg_array_30_42_real;
      end
      6'b101011 : begin
        _zz_4494_ = int_reg_array_30_43_imag;
        _zz_4495_ = int_reg_array_30_43_real;
      end
      6'b101100 : begin
        _zz_4494_ = int_reg_array_30_44_imag;
        _zz_4495_ = int_reg_array_30_44_real;
      end
      6'b101101 : begin
        _zz_4494_ = int_reg_array_30_45_imag;
        _zz_4495_ = int_reg_array_30_45_real;
      end
      6'b101110 : begin
        _zz_4494_ = int_reg_array_30_46_imag;
        _zz_4495_ = int_reg_array_30_46_real;
      end
      6'b101111 : begin
        _zz_4494_ = int_reg_array_30_47_imag;
        _zz_4495_ = int_reg_array_30_47_real;
      end
      6'b110000 : begin
        _zz_4494_ = int_reg_array_30_48_imag;
        _zz_4495_ = int_reg_array_30_48_real;
      end
      6'b110001 : begin
        _zz_4494_ = int_reg_array_30_49_imag;
        _zz_4495_ = int_reg_array_30_49_real;
      end
      6'b110010 : begin
        _zz_4494_ = int_reg_array_30_50_imag;
        _zz_4495_ = int_reg_array_30_50_real;
      end
      6'b110011 : begin
        _zz_4494_ = int_reg_array_30_51_imag;
        _zz_4495_ = int_reg_array_30_51_real;
      end
      6'b110100 : begin
        _zz_4494_ = int_reg_array_30_52_imag;
        _zz_4495_ = int_reg_array_30_52_real;
      end
      6'b110101 : begin
        _zz_4494_ = int_reg_array_30_53_imag;
        _zz_4495_ = int_reg_array_30_53_real;
      end
      6'b110110 : begin
        _zz_4494_ = int_reg_array_30_54_imag;
        _zz_4495_ = int_reg_array_30_54_real;
      end
      6'b110111 : begin
        _zz_4494_ = int_reg_array_30_55_imag;
        _zz_4495_ = int_reg_array_30_55_real;
      end
      6'b111000 : begin
        _zz_4494_ = int_reg_array_30_56_imag;
        _zz_4495_ = int_reg_array_30_56_real;
      end
      6'b111001 : begin
        _zz_4494_ = int_reg_array_30_57_imag;
        _zz_4495_ = int_reg_array_30_57_real;
      end
      6'b111010 : begin
        _zz_4494_ = int_reg_array_30_58_imag;
        _zz_4495_ = int_reg_array_30_58_real;
      end
      6'b111011 : begin
        _zz_4494_ = int_reg_array_30_59_imag;
        _zz_4495_ = int_reg_array_30_59_real;
      end
      6'b111100 : begin
        _zz_4494_ = int_reg_array_30_60_imag;
        _zz_4495_ = int_reg_array_30_60_real;
      end
      6'b111101 : begin
        _zz_4494_ = int_reg_array_30_61_imag;
        _zz_4495_ = int_reg_array_30_61_real;
      end
      6'b111110 : begin
        _zz_4494_ = int_reg_array_30_62_imag;
        _zz_4495_ = int_reg_array_30_62_real;
      end
      default : begin
        _zz_4494_ = int_reg_array_30_63_imag;
        _zz_4495_ = int_reg_array_30_63_real;
      end
    endcase
  end

  always @(*) begin
    case(_zz_2156_)
      6'b000000 : begin
        _zz_4496_ = int_reg_array_31_0_imag;
        _zz_4497_ = int_reg_array_31_0_real;
      end
      6'b000001 : begin
        _zz_4496_ = int_reg_array_31_1_imag;
        _zz_4497_ = int_reg_array_31_1_real;
      end
      6'b000010 : begin
        _zz_4496_ = int_reg_array_31_2_imag;
        _zz_4497_ = int_reg_array_31_2_real;
      end
      6'b000011 : begin
        _zz_4496_ = int_reg_array_31_3_imag;
        _zz_4497_ = int_reg_array_31_3_real;
      end
      6'b000100 : begin
        _zz_4496_ = int_reg_array_31_4_imag;
        _zz_4497_ = int_reg_array_31_4_real;
      end
      6'b000101 : begin
        _zz_4496_ = int_reg_array_31_5_imag;
        _zz_4497_ = int_reg_array_31_5_real;
      end
      6'b000110 : begin
        _zz_4496_ = int_reg_array_31_6_imag;
        _zz_4497_ = int_reg_array_31_6_real;
      end
      6'b000111 : begin
        _zz_4496_ = int_reg_array_31_7_imag;
        _zz_4497_ = int_reg_array_31_7_real;
      end
      6'b001000 : begin
        _zz_4496_ = int_reg_array_31_8_imag;
        _zz_4497_ = int_reg_array_31_8_real;
      end
      6'b001001 : begin
        _zz_4496_ = int_reg_array_31_9_imag;
        _zz_4497_ = int_reg_array_31_9_real;
      end
      6'b001010 : begin
        _zz_4496_ = int_reg_array_31_10_imag;
        _zz_4497_ = int_reg_array_31_10_real;
      end
      6'b001011 : begin
        _zz_4496_ = int_reg_array_31_11_imag;
        _zz_4497_ = int_reg_array_31_11_real;
      end
      6'b001100 : begin
        _zz_4496_ = int_reg_array_31_12_imag;
        _zz_4497_ = int_reg_array_31_12_real;
      end
      6'b001101 : begin
        _zz_4496_ = int_reg_array_31_13_imag;
        _zz_4497_ = int_reg_array_31_13_real;
      end
      6'b001110 : begin
        _zz_4496_ = int_reg_array_31_14_imag;
        _zz_4497_ = int_reg_array_31_14_real;
      end
      6'b001111 : begin
        _zz_4496_ = int_reg_array_31_15_imag;
        _zz_4497_ = int_reg_array_31_15_real;
      end
      6'b010000 : begin
        _zz_4496_ = int_reg_array_31_16_imag;
        _zz_4497_ = int_reg_array_31_16_real;
      end
      6'b010001 : begin
        _zz_4496_ = int_reg_array_31_17_imag;
        _zz_4497_ = int_reg_array_31_17_real;
      end
      6'b010010 : begin
        _zz_4496_ = int_reg_array_31_18_imag;
        _zz_4497_ = int_reg_array_31_18_real;
      end
      6'b010011 : begin
        _zz_4496_ = int_reg_array_31_19_imag;
        _zz_4497_ = int_reg_array_31_19_real;
      end
      6'b010100 : begin
        _zz_4496_ = int_reg_array_31_20_imag;
        _zz_4497_ = int_reg_array_31_20_real;
      end
      6'b010101 : begin
        _zz_4496_ = int_reg_array_31_21_imag;
        _zz_4497_ = int_reg_array_31_21_real;
      end
      6'b010110 : begin
        _zz_4496_ = int_reg_array_31_22_imag;
        _zz_4497_ = int_reg_array_31_22_real;
      end
      6'b010111 : begin
        _zz_4496_ = int_reg_array_31_23_imag;
        _zz_4497_ = int_reg_array_31_23_real;
      end
      6'b011000 : begin
        _zz_4496_ = int_reg_array_31_24_imag;
        _zz_4497_ = int_reg_array_31_24_real;
      end
      6'b011001 : begin
        _zz_4496_ = int_reg_array_31_25_imag;
        _zz_4497_ = int_reg_array_31_25_real;
      end
      6'b011010 : begin
        _zz_4496_ = int_reg_array_31_26_imag;
        _zz_4497_ = int_reg_array_31_26_real;
      end
      6'b011011 : begin
        _zz_4496_ = int_reg_array_31_27_imag;
        _zz_4497_ = int_reg_array_31_27_real;
      end
      6'b011100 : begin
        _zz_4496_ = int_reg_array_31_28_imag;
        _zz_4497_ = int_reg_array_31_28_real;
      end
      6'b011101 : begin
        _zz_4496_ = int_reg_array_31_29_imag;
        _zz_4497_ = int_reg_array_31_29_real;
      end
      6'b011110 : begin
        _zz_4496_ = int_reg_array_31_30_imag;
        _zz_4497_ = int_reg_array_31_30_real;
      end
      6'b011111 : begin
        _zz_4496_ = int_reg_array_31_31_imag;
        _zz_4497_ = int_reg_array_31_31_real;
      end
      6'b100000 : begin
        _zz_4496_ = int_reg_array_31_32_imag;
        _zz_4497_ = int_reg_array_31_32_real;
      end
      6'b100001 : begin
        _zz_4496_ = int_reg_array_31_33_imag;
        _zz_4497_ = int_reg_array_31_33_real;
      end
      6'b100010 : begin
        _zz_4496_ = int_reg_array_31_34_imag;
        _zz_4497_ = int_reg_array_31_34_real;
      end
      6'b100011 : begin
        _zz_4496_ = int_reg_array_31_35_imag;
        _zz_4497_ = int_reg_array_31_35_real;
      end
      6'b100100 : begin
        _zz_4496_ = int_reg_array_31_36_imag;
        _zz_4497_ = int_reg_array_31_36_real;
      end
      6'b100101 : begin
        _zz_4496_ = int_reg_array_31_37_imag;
        _zz_4497_ = int_reg_array_31_37_real;
      end
      6'b100110 : begin
        _zz_4496_ = int_reg_array_31_38_imag;
        _zz_4497_ = int_reg_array_31_38_real;
      end
      6'b100111 : begin
        _zz_4496_ = int_reg_array_31_39_imag;
        _zz_4497_ = int_reg_array_31_39_real;
      end
      6'b101000 : begin
        _zz_4496_ = int_reg_array_31_40_imag;
        _zz_4497_ = int_reg_array_31_40_real;
      end
      6'b101001 : begin
        _zz_4496_ = int_reg_array_31_41_imag;
        _zz_4497_ = int_reg_array_31_41_real;
      end
      6'b101010 : begin
        _zz_4496_ = int_reg_array_31_42_imag;
        _zz_4497_ = int_reg_array_31_42_real;
      end
      6'b101011 : begin
        _zz_4496_ = int_reg_array_31_43_imag;
        _zz_4497_ = int_reg_array_31_43_real;
      end
      6'b101100 : begin
        _zz_4496_ = int_reg_array_31_44_imag;
        _zz_4497_ = int_reg_array_31_44_real;
      end
      6'b101101 : begin
        _zz_4496_ = int_reg_array_31_45_imag;
        _zz_4497_ = int_reg_array_31_45_real;
      end
      6'b101110 : begin
        _zz_4496_ = int_reg_array_31_46_imag;
        _zz_4497_ = int_reg_array_31_46_real;
      end
      6'b101111 : begin
        _zz_4496_ = int_reg_array_31_47_imag;
        _zz_4497_ = int_reg_array_31_47_real;
      end
      6'b110000 : begin
        _zz_4496_ = int_reg_array_31_48_imag;
        _zz_4497_ = int_reg_array_31_48_real;
      end
      6'b110001 : begin
        _zz_4496_ = int_reg_array_31_49_imag;
        _zz_4497_ = int_reg_array_31_49_real;
      end
      6'b110010 : begin
        _zz_4496_ = int_reg_array_31_50_imag;
        _zz_4497_ = int_reg_array_31_50_real;
      end
      6'b110011 : begin
        _zz_4496_ = int_reg_array_31_51_imag;
        _zz_4497_ = int_reg_array_31_51_real;
      end
      6'b110100 : begin
        _zz_4496_ = int_reg_array_31_52_imag;
        _zz_4497_ = int_reg_array_31_52_real;
      end
      6'b110101 : begin
        _zz_4496_ = int_reg_array_31_53_imag;
        _zz_4497_ = int_reg_array_31_53_real;
      end
      6'b110110 : begin
        _zz_4496_ = int_reg_array_31_54_imag;
        _zz_4497_ = int_reg_array_31_54_real;
      end
      6'b110111 : begin
        _zz_4496_ = int_reg_array_31_55_imag;
        _zz_4497_ = int_reg_array_31_55_real;
      end
      6'b111000 : begin
        _zz_4496_ = int_reg_array_31_56_imag;
        _zz_4497_ = int_reg_array_31_56_real;
      end
      6'b111001 : begin
        _zz_4496_ = int_reg_array_31_57_imag;
        _zz_4497_ = int_reg_array_31_57_real;
      end
      6'b111010 : begin
        _zz_4496_ = int_reg_array_31_58_imag;
        _zz_4497_ = int_reg_array_31_58_real;
      end
      6'b111011 : begin
        _zz_4496_ = int_reg_array_31_59_imag;
        _zz_4497_ = int_reg_array_31_59_real;
      end
      6'b111100 : begin
        _zz_4496_ = int_reg_array_31_60_imag;
        _zz_4497_ = int_reg_array_31_60_real;
      end
      6'b111101 : begin
        _zz_4496_ = int_reg_array_31_61_imag;
        _zz_4497_ = int_reg_array_31_61_real;
      end
      6'b111110 : begin
        _zz_4496_ = int_reg_array_31_62_imag;
        _zz_4497_ = int_reg_array_31_62_real;
      end
      default : begin
        _zz_4496_ = int_reg_array_31_63_imag;
        _zz_4497_ = int_reg_array_31_63_real;
      end
    endcase
  end

  always @(*) begin
    case(_zz_2225_)
      6'b000000 : begin
        _zz_4498_ = int_reg_array_32_0_imag;
        _zz_4499_ = int_reg_array_32_0_real;
      end
      6'b000001 : begin
        _zz_4498_ = int_reg_array_32_1_imag;
        _zz_4499_ = int_reg_array_32_1_real;
      end
      6'b000010 : begin
        _zz_4498_ = int_reg_array_32_2_imag;
        _zz_4499_ = int_reg_array_32_2_real;
      end
      6'b000011 : begin
        _zz_4498_ = int_reg_array_32_3_imag;
        _zz_4499_ = int_reg_array_32_3_real;
      end
      6'b000100 : begin
        _zz_4498_ = int_reg_array_32_4_imag;
        _zz_4499_ = int_reg_array_32_4_real;
      end
      6'b000101 : begin
        _zz_4498_ = int_reg_array_32_5_imag;
        _zz_4499_ = int_reg_array_32_5_real;
      end
      6'b000110 : begin
        _zz_4498_ = int_reg_array_32_6_imag;
        _zz_4499_ = int_reg_array_32_6_real;
      end
      6'b000111 : begin
        _zz_4498_ = int_reg_array_32_7_imag;
        _zz_4499_ = int_reg_array_32_7_real;
      end
      6'b001000 : begin
        _zz_4498_ = int_reg_array_32_8_imag;
        _zz_4499_ = int_reg_array_32_8_real;
      end
      6'b001001 : begin
        _zz_4498_ = int_reg_array_32_9_imag;
        _zz_4499_ = int_reg_array_32_9_real;
      end
      6'b001010 : begin
        _zz_4498_ = int_reg_array_32_10_imag;
        _zz_4499_ = int_reg_array_32_10_real;
      end
      6'b001011 : begin
        _zz_4498_ = int_reg_array_32_11_imag;
        _zz_4499_ = int_reg_array_32_11_real;
      end
      6'b001100 : begin
        _zz_4498_ = int_reg_array_32_12_imag;
        _zz_4499_ = int_reg_array_32_12_real;
      end
      6'b001101 : begin
        _zz_4498_ = int_reg_array_32_13_imag;
        _zz_4499_ = int_reg_array_32_13_real;
      end
      6'b001110 : begin
        _zz_4498_ = int_reg_array_32_14_imag;
        _zz_4499_ = int_reg_array_32_14_real;
      end
      6'b001111 : begin
        _zz_4498_ = int_reg_array_32_15_imag;
        _zz_4499_ = int_reg_array_32_15_real;
      end
      6'b010000 : begin
        _zz_4498_ = int_reg_array_32_16_imag;
        _zz_4499_ = int_reg_array_32_16_real;
      end
      6'b010001 : begin
        _zz_4498_ = int_reg_array_32_17_imag;
        _zz_4499_ = int_reg_array_32_17_real;
      end
      6'b010010 : begin
        _zz_4498_ = int_reg_array_32_18_imag;
        _zz_4499_ = int_reg_array_32_18_real;
      end
      6'b010011 : begin
        _zz_4498_ = int_reg_array_32_19_imag;
        _zz_4499_ = int_reg_array_32_19_real;
      end
      6'b010100 : begin
        _zz_4498_ = int_reg_array_32_20_imag;
        _zz_4499_ = int_reg_array_32_20_real;
      end
      6'b010101 : begin
        _zz_4498_ = int_reg_array_32_21_imag;
        _zz_4499_ = int_reg_array_32_21_real;
      end
      6'b010110 : begin
        _zz_4498_ = int_reg_array_32_22_imag;
        _zz_4499_ = int_reg_array_32_22_real;
      end
      6'b010111 : begin
        _zz_4498_ = int_reg_array_32_23_imag;
        _zz_4499_ = int_reg_array_32_23_real;
      end
      6'b011000 : begin
        _zz_4498_ = int_reg_array_32_24_imag;
        _zz_4499_ = int_reg_array_32_24_real;
      end
      6'b011001 : begin
        _zz_4498_ = int_reg_array_32_25_imag;
        _zz_4499_ = int_reg_array_32_25_real;
      end
      6'b011010 : begin
        _zz_4498_ = int_reg_array_32_26_imag;
        _zz_4499_ = int_reg_array_32_26_real;
      end
      6'b011011 : begin
        _zz_4498_ = int_reg_array_32_27_imag;
        _zz_4499_ = int_reg_array_32_27_real;
      end
      6'b011100 : begin
        _zz_4498_ = int_reg_array_32_28_imag;
        _zz_4499_ = int_reg_array_32_28_real;
      end
      6'b011101 : begin
        _zz_4498_ = int_reg_array_32_29_imag;
        _zz_4499_ = int_reg_array_32_29_real;
      end
      6'b011110 : begin
        _zz_4498_ = int_reg_array_32_30_imag;
        _zz_4499_ = int_reg_array_32_30_real;
      end
      6'b011111 : begin
        _zz_4498_ = int_reg_array_32_31_imag;
        _zz_4499_ = int_reg_array_32_31_real;
      end
      6'b100000 : begin
        _zz_4498_ = int_reg_array_32_32_imag;
        _zz_4499_ = int_reg_array_32_32_real;
      end
      6'b100001 : begin
        _zz_4498_ = int_reg_array_32_33_imag;
        _zz_4499_ = int_reg_array_32_33_real;
      end
      6'b100010 : begin
        _zz_4498_ = int_reg_array_32_34_imag;
        _zz_4499_ = int_reg_array_32_34_real;
      end
      6'b100011 : begin
        _zz_4498_ = int_reg_array_32_35_imag;
        _zz_4499_ = int_reg_array_32_35_real;
      end
      6'b100100 : begin
        _zz_4498_ = int_reg_array_32_36_imag;
        _zz_4499_ = int_reg_array_32_36_real;
      end
      6'b100101 : begin
        _zz_4498_ = int_reg_array_32_37_imag;
        _zz_4499_ = int_reg_array_32_37_real;
      end
      6'b100110 : begin
        _zz_4498_ = int_reg_array_32_38_imag;
        _zz_4499_ = int_reg_array_32_38_real;
      end
      6'b100111 : begin
        _zz_4498_ = int_reg_array_32_39_imag;
        _zz_4499_ = int_reg_array_32_39_real;
      end
      6'b101000 : begin
        _zz_4498_ = int_reg_array_32_40_imag;
        _zz_4499_ = int_reg_array_32_40_real;
      end
      6'b101001 : begin
        _zz_4498_ = int_reg_array_32_41_imag;
        _zz_4499_ = int_reg_array_32_41_real;
      end
      6'b101010 : begin
        _zz_4498_ = int_reg_array_32_42_imag;
        _zz_4499_ = int_reg_array_32_42_real;
      end
      6'b101011 : begin
        _zz_4498_ = int_reg_array_32_43_imag;
        _zz_4499_ = int_reg_array_32_43_real;
      end
      6'b101100 : begin
        _zz_4498_ = int_reg_array_32_44_imag;
        _zz_4499_ = int_reg_array_32_44_real;
      end
      6'b101101 : begin
        _zz_4498_ = int_reg_array_32_45_imag;
        _zz_4499_ = int_reg_array_32_45_real;
      end
      6'b101110 : begin
        _zz_4498_ = int_reg_array_32_46_imag;
        _zz_4499_ = int_reg_array_32_46_real;
      end
      6'b101111 : begin
        _zz_4498_ = int_reg_array_32_47_imag;
        _zz_4499_ = int_reg_array_32_47_real;
      end
      6'b110000 : begin
        _zz_4498_ = int_reg_array_32_48_imag;
        _zz_4499_ = int_reg_array_32_48_real;
      end
      6'b110001 : begin
        _zz_4498_ = int_reg_array_32_49_imag;
        _zz_4499_ = int_reg_array_32_49_real;
      end
      6'b110010 : begin
        _zz_4498_ = int_reg_array_32_50_imag;
        _zz_4499_ = int_reg_array_32_50_real;
      end
      6'b110011 : begin
        _zz_4498_ = int_reg_array_32_51_imag;
        _zz_4499_ = int_reg_array_32_51_real;
      end
      6'b110100 : begin
        _zz_4498_ = int_reg_array_32_52_imag;
        _zz_4499_ = int_reg_array_32_52_real;
      end
      6'b110101 : begin
        _zz_4498_ = int_reg_array_32_53_imag;
        _zz_4499_ = int_reg_array_32_53_real;
      end
      6'b110110 : begin
        _zz_4498_ = int_reg_array_32_54_imag;
        _zz_4499_ = int_reg_array_32_54_real;
      end
      6'b110111 : begin
        _zz_4498_ = int_reg_array_32_55_imag;
        _zz_4499_ = int_reg_array_32_55_real;
      end
      6'b111000 : begin
        _zz_4498_ = int_reg_array_32_56_imag;
        _zz_4499_ = int_reg_array_32_56_real;
      end
      6'b111001 : begin
        _zz_4498_ = int_reg_array_32_57_imag;
        _zz_4499_ = int_reg_array_32_57_real;
      end
      6'b111010 : begin
        _zz_4498_ = int_reg_array_32_58_imag;
        _zz_4499_ = int_reg_array_32_58_real;
      end
      6'b111011 : begin
        _zz_4498_ = int_reg_array_32_59_imag;
        _zz_4499_ = int_reg_array_32_59_real;
      end
      6'b111100 : begin
        _zz_4498_ = int_reg_array_32_60_imag;
        _zz_4499_ = int_reg_array_32_60_real;
      end
      6'b111101 : begin
        _zz_4498_ = int_reg_array_32_61_imag;
        _zz_4499_ = int_reg_array_32_61_real;
      end
      6'b111110 : begin
        _zz_4498_ = int_reg_array_32_62_imag;
        _zz_4499_ = int_reg_array_32_62_real;
      end
      default : begin
        _zz_4498_ = int_reg_array_32_63_imag;
        _zz_4499_ = int_reg_array_32_63_real;
      end
    endcase
  end

  always @(*) begin
    case(_zz_2294_)
      6'b000000 : begin
        _zz_4500_ = int_reg_array_33_0_imag;
        _zz_4501_ = int_reg_array_33_0_real;
      end
      6'b000001 : begin
        _zz_4500_ = int_reg_array_33_1_imag;
        _zz_4501_ = int_reg_array_33_1_real;
      end
      6'b000010 : begin
        _zz_4500_ = int_reg_array_33_2_imag;
        _zz_4501_ = int_reg_array_33_2_real;
      end
      6'b000011 : begin
        _zz_4500_ = int_reg_array_33_3_imag;
        _zz_4501_ = int_reg_array_33_3_real;
      end
      6'b000100 : begin
        _zz_4500_ = int_reg_array_33_4_imag;
        _zz_4501_ = int_reg_array_33_4_real;
      end
      6'b000101 : begin
        _zz_4500_ = int_reg_array_33_5_imag;
        _zz_4501_ = int_reg_array_33_5_real;
      end
      6'b000110 : begin
        _zz_4500_ = int_reg_array_33_6_imag;
        _zz_4501_ = int_reg_array_33_6_real;
      end
      6'b000111 : begin
        _zz_4500_ = int_reg_array_33_7_imag;
        _zz_4501_ = int_reg_array_33_7_real;
      end
      6'b001000 : begin
        _zz_4500_ = int_reg_array_33_8_imag;
        _zz_4501_ = int_reg_array_33_8_real;
      end
      6'b001001 : begin
        _zz_4500_ = int_reg_array_33_9_imag;
        _zz_4501_ = int_reg_array_33_9_real;
      end
      6'b001010 : begin
        _zz_4500_ = int_reg_array_33_10_imag;
        _zz_4501_ = int_reg_array_33_10_real;
      end
      6'b001011 : begin
        _zz_4500_ = int_reg_array_33_11_imag;
        _zz_4501_ = int_reg_array_33_11_real;
      end
      6'b001100 : begin
        _zz_4500_ = int_reg_array_33_12_imag;
        _zz_4501_ = int_reg_array_33_12_real;
      end
      6'b001101 : begin
        _zz_4500_ = int_reg_array_33_13_imag;
        _zz_4501_ = int_reg_array_33_13_real;
      end
      6'b001110 : begin
        _zz_4500_ = int_reg_array_33_14_imag;
        _zz_4501_ = int_reg_array_33_14_real;
      end
      6'b001111 : begin
        _zz_4500_ = int_reg_array_33_15_imag;
        _zz_4501_ = int_reg_array_33_15_real;
      end
      6'b010000 : begin
        _zz_4500_ = int_reg_array_33_16_imag;
        _zz_4501_ = int_reg_array_33_16_real;
      end
      6'b010001 : begin
        _zz_4500_ = int_reg_array_33_17_imag;
        _zz_4501_ = int_reg_array_33_17_real;
      end
      6'b010010 : begin
        _zz_4500_ = int_reg_array_33_18_imag;
        _zz_4501_ = int_reg_array_33_18_real;
      end
      6'b010011 : begin
        _zz_4500_ = int_reg_array_33_19_imag;
        _zz_4501_ = int_reg_array_33_19_real;
      end
      6'b010100 : begin
        _zz_4500_ = int_reg_array_33_20_imag;
        _zz_4501_ = int_reg_array_33_20_real;
      end
      6'b010101 : begin
        _zz_4500_ = int_reg_array_33_21_imag;
        _zz_4501_ = int_reg_array_33_21_real;
      end
      6'b010110 : begin
        _zz_4500_ = int_reg_array_33_22_imag;
        _zz_4501_ = int_reg_array_33_22_real;
      end
      6'b010111 : begin
        _zz_4500_ = int_reg_array_33_23_imag;
        _zz_4501_ = int_reg_array_33_23_real;
      end
      6'b011000 : begin
        _zz_4500_ = int_reg_array_33_24_imag;
        _zz_4501_ = int_reg_array_33_24_real;
      end
      6'b011001 : begin
        _zz_4500_ = int_reg_array_33_25_imag;
        _zz_4501_ = int_reg_array_33_25_real;
      end
      6'b011010 : begin
        _zz_4500_ = int_reg_array_33_26_imag;
        _zz_4501_ = int_reg_array_33_26_real;
      end
      6'b011011 : begin
        _zz_4500_ = int_reg_array_33_27_imag;
        _zz_4501_ = int_reg_array_33_27_real;
      end
      6'b011100 : begin
        _zz_4500_ = int_reg_array_33_28_imag;
        _zz_4501_ = int_reg_array_33_28_real;
      end
      6'b011101 : begin
        _zz_4500_ = int_reg_array_33_29_imag;
        _zz_4501_ = int_reg_array_33_29_real;
      end
      6'b011110 : begin
        _zz_4500_ = int_reg_array_33_30_imag;
        _zz_4501_ = int_reg_array_33_30_real;
      end
      6'b011111 : begin
        _zz_4500_ = int_reg_array_33_31_imag;
        _zz_4501_ = int_reg_array_33_31_real;
      end
      6'b100000 : begin
        _zz_4500_ = int_reg_array_33_32_imag;
        _zz_4501_ = int_reg_array_33_32_real;
      end
      6'b100001 : begin
        _zz_4500_ = int_reg_array_33_33_imag;
        _zz_4501_ = int_reg_array_33_33_real;
      end
      6'b100010 : begin
        _zz_4500_ = int_reg_array_33_34_imag;
        _zz_4501_ = int_reg_array_33_34_real;
      end
      6'b100011 : begin
        _zz_4500_ = int_reg_array_33_35_imag;
        _zz_4501_ = int_reg_array_33_35_real;
      end
      6'b100100 : begin
        _zz_4500_ = int_reg_array_33_36_imag;
        _zz_4501_ = int_reg_array_33_36_real;
      end
      6'b100101 : begin
        _zz_4500_ = int_reg_array_33_37_imag;
        _zz_4501_ = int_reg_array_33_37_real;
      end
      6'b100110 : begin
        _zz_4500_ = int_reg_array_33_38_imag;
        _zz_4501_ = int_reg_array_33_38_real;
      end
      6'b100111 : begin
        _zz_4500_ = int_reg_array_33_39_imag;
        _zz_4501_ = int_reg_array_33_39_real;
      end
      6'b101000 : begin
        _zz_4500_ = int_reg_array_33_40_imag;
        _zz_4501_ = int_reg_array_33_40_real;
      end
      6'b101001 : begin
        _zz_4500_ = int_reg_array_33_41_imag;
        _zz_4501_ = int_reg_array_33_41_real;
      end
      6'b101010 : begin
        _zz_4500_ = int_reg_array_33_42_imag;
        _zz_4501_ = int_reg_array_33_42_real;
      end
      6'b101011 : begin
        _zz_4500_ = int_reg_array_33_43_imag;
        _zz_4501_ = int_reg_array_33_43_real;
      end
      6'b101100 : begin
        _zz_4500_ = int_reg_array_33_44_imag;
        _zz_4501_ = int_reg_array_33_44_real;
      end
      6'b101101 : begin
        _zz_4500_ = int_reg_array_33_45_imag;
        _zz_4501_ = int_reg_array_33_45_real;
      end
      6'b101110 : begin
        _zz_4500_ = int_reg_array_33_46_imag;
        _zz_4501_ = int_reg_array_33_46_real;
      end
      6'b101111 : begin
        _zz_4500_ = int_reg_array_33_47_imag;
        _zz_4501_ = int_reg_array_33_47_real;
      end
      6'b110000 : begin
        _zz_4500_ = int_reg_array_33_48_imag;
        _zz_4501_ = int_reg_array_33_48_real;
      end
      6'b110001 : begin
        _zz_4500_ = int_reg_array_33_49_imag;
        _zz_4501_ = int_reg_array_33_49_real;
      end
      6'b110010 : begin
        _zz_4500_ = int_reg_array_33_50_imag;
        _zz_4501_ = int_reg_array_33_50_real;
      end
      6'b110011 : begin
        _zz_4500_ = int_reg_array_33_51_imag;
        _zz_4501_ = int_reg_array_33_51_real;
      end
      6'b110100 : begin
        _zz_4500_ = int_reg_array_33_52_imag;
        _zz_4501_ = int_reg_array_33_52_real;
      end
      6'b110101 : begin
        _zz_4500_ = int_reg_array_33_53_imag;
        _zz_4501_ = int_reg_array_33_53_real;
      end
      6'b110110 : begin
        _zz_4500_ = int_reg_array_33_54_imag;
        _zz_4501_ = int_reg_array_33_54_real;
      end
      6'b110111 : begin
        _zz_4500_ = int_reg_array_33_55_imag;
        _zz_4501_ = int_reg_array_33_55_real;
      end
      6'b111000 : begin
        _zz_4500_ = int_reg_array_33_56_imag;
        _zz_4501_ = int_reg_array_33_56_real;
      end
      6'b111001 : begin
        _zz_4500_ = int_reg_array_33_57_imag;
        _zz_4501_ = int_reg_array_33_57_real;
      end
      6'b111010 : begin
        _zz_4500_ = int_reg_array_33_58_imag;
        _zz_4501_ = int_reg_array_33_58_real;
      end
      6'b111011 : begin
        _zz_4500_ = int_reg_array_33_59_imag;
        _zz_4501_ = int_reg_array_33_59_real;
      end
      6'b111100 : begin
        _zz_4500_ = int_reg_array_33_60_imag;
        _zz_4501_ = int_reg_array_33_60_real;
      end
      6'b111101 : begin
        _zz_4500_ = int_reg_array_33_61_imag;
        _zz_4501_ = int_reg_array_33_61_real;
      end
      6'b111110 : begin
        _zz_4500_ = int_reg_array_33_62_imag;
        _zz_4501_ = int_reg_array_33_62_real;
      end
      default : begin
        _zz_4500_ = int_reg_array_33_63_imag;
        _zz_4501_ = int_reg_array_33_63_real;
      end
    endcase
  end

  always @(*) begin
    case(_zz_2363_)
      6'b000000 : begin
        _zz_4502_ = int_reg_array_34_0_imag;
        _zz_4503_ = int_reg_array_34_0_real;
      end
      6'b000001 : begin
        _zz_4502_ = int_reg_array_34_1_imag;
        _zz_4503_ = int_reg_array_34_1_real;
      end
      6'b000010 : begin
        _zz_4502_ = int_reg_array_34_2_imag;
        _zz_4503_ = int_reg_array_34_2_real;
      end
      6'b000011 : begin
        _zz_4502_ = int_reg_array_34_3_imag;
        _zz_4503_ = int_reg_array_34_3_real;
      end
      6'b000100 : begin
        _zz_4502_ = int_reg_array_34_4_imag;
        _zz_4503_ = int_reg_array_34_4_real;
      end
      6'b000101 : begin
        _zz_4502_ = int_reg_array_34_5_imag;
        _zz_4503_ = int_reg_array_34_5_real;
      end
      6'b000110 : begin
        _zz_4502_ = int_reg_array_34_6_imag;
        _zz_4503_ = int_reg_array_34_6_real;
      end
      6'b000111 : begin
        _zz_4502_ = int_reg_array_34_7_imag;
        _zz_4503_ = int_reg_array_34_7_real;
      end
      6'b001000 : begin
        _zz_4502_ = int_reg_array_34_8_imag;
        _zz_4503_ = int_reg_array_34_8_real;
      end
      6'b001001 : begin
        _zz_4502_ = int_reg_array_34_9_imag;
        _zz_4503_ = int_reg_array_34_9_real;
      end
      6'b001010 : begin
        _zz_4502_ = int_reg_array_34_10_imag;
        _zz_4503_ = int_reg_array_34_10_real;
      end
      6'b001011 : begin
        _zz_4502_ = int_reg_array_34_11_imag;
        _zz_4503_ = int_reg_array_34_11_real;
      end
      6'b001100 : begin
        _zz_4502_ = int_reg_array_34_12_imag;
        _zz_4503_ = int_reg_array_34_12_real;
      end
      6'b001101 : begin
        _zz_4502_ = int_reg_array_34_13_imag;
        _zz_4503_ = int_reg_array_34_13_real;
      end
      6'b001110 : begin
        _zz_4502_ = int_reg_array_34_14_imag;
        _zz_4503_ = int_reg_array_34_14_real;
      end
      6'b001111 : begin
        _zz_4502_ = int_reg_array_34_15_imag;
        _zz_4503_ = int_reg_array_34_15_real;
      end
      6'b010000 : begin
        _zz_4502_ = int_reg_array_34_16_imag;
        _zz_4503_ = int_reg_array_34_16_real;
      end
      6'b010001 : begin
        _zz_4502_ = int_reg_array_34_17_imag;
        _zz_4503_ = int_reg_array_34_17_real;
      end
      6'b010010 : begin
        _zz_4502_ = int_reg_array_34_18_imag;
        _zz_4503_ = int_reg_array_34_18_real;
      end
      6'b010011 : begin
        _zz_4502_ = int_reg_array_34_19_imag;
        _zz_4503_ = int_reg_array_34_19_real;
      end
      6'b010100 : begin
        _zz_4502_ = int_reg_array_34_20_imag;
        _zz_4503_ = int_reg_array_34_20_real;
      end
      6'b010101 : begin
        _zz_4502_ = int_reg_array_34_21_imag;
        _zz_4503_ = int_reg_array_34_21_real;
      end
      6'b010110 : begin
        _zz_4502_ = int_reg_array_34_22_imag;
        _zz_4503_ = int_reg_array_34_22_real;
      end
      6'b010111 : begin
        _zz_4502_ = int_reg_array_34_23_imag;
        _zz_4503_ = int_reg_array_34_23_real;
      end
      6'b011000 : begin
        _zz_4502_ = int_reg_array_34_24_imag;
        _zz_4503_ = int_reg_array_34_24_real;
      end
      6'b011001 : begin
        _zz_4502_ = int_reg_array_34_25_imag;
        _zz_4503_ = int_reg_array_34_25_real;
      end
      6'b011010 : begin
        _zz_4502_ = int_reg_array_34_26_imag;
        _zz_4503_ = int_reg_array_34_26_real;
      end
      6'b011011 : begin
        _zz_4502_ = int_reg_array_34_27_imag;
        _zz_4503_ = int_reg_array_34_27_real;
      end
      6'b011100 : begin
        _zz_4502_ = int_reg_array_34_28_imag;
        _zz_4503_ = int_reg_array_34_28_real;
      end
      6'b011101 : begin
        _zz_4502_ = int_reg_array_34_29_imag;
        _zz_4503_ = int_reg_array_34_29_real;
      end
      6'b011110 : begin
        _zz_4502_ = int_reg_array_34_30_imag;
        _zz_4503_ = int_reg_array_34_30_real;
      end
      6'b011111 : begin
        _zz_4502_ = int_reg_array_34_31_imag;
        _zz_4503_ = int_reg_array_34_31_real;
      end
      6'b100000 : begin
        _zz_4502_ = int_reg_array_34_32_imag;
        _zz_4503_ = int_reg_array_34_32_real;
      end
      6'b100001 : begin
        _zz_4502_ = int_reg_array_34_33_imag;
        _zz_4503_ = int_reg_array_34_33_real;
      end
      6'b100010 : begin
        _zz_4502_ = int_reg_array_34_34_imag;
        _zz_4503_ = int_reg_array_34_34_real;
      end
      6'b100011 : begin
        _zz_4502_ = int_reg_array_34_35_imag;
        _zz_4503_ = int_reg_array_34_35_real;
      end
      6'b100100 : begin
        _zz_4502_ = int_reg_array_34_36_imag;
        _zz_4503_ = int_reg_array_34_36_real;
      end
      6'b100101 : begin
        _zz_4502_ = int_reg_array_34_37_imag;
        _zz_4503_ = int_reg_array_34_37_real;
      end
      6'b100110 : begin
        _zz_4502_ = int_reg_array_34_38_imag;
        _zz_4503_ = int_reg_array_34_38_real;
      end
      6'b100111 : begin
        _zz_4502_ = int_reg_array_34_39_imag;
        _zz_4503_ = int_reg_array_34_39_real;
      end
      6'b101000 : begin
        _zz_4502_ = int_reg_array_34_40_imag;
        _zz_4503_ = int_reg_array_34_40_real;
      end
      6'b101001 : begin
        _zz_4502_ = int_reg_array_34_41_imag;
        _zz_4503_ = int_reg_array_34_41_real;
      end
      6'b101010 : begin
        _zz_4502_ = int_reg_array_34_42_imag;
        _zz_4503_ = int_reg_array_34_42_real;
      end
      6'b101011 : begin
        _zz_4502_ = int_reg_array_34_43_imag;
        _zz_4503_ = int_reg_array_34_43_real;
      end
      6'b101100 : begin
        _zz_4502_ = int_reg_array_34_44_imag;
        _zz_4503_ = int_reg_array_34_44_real;
      end
      6'b101101 : begin
        _zz_4502_ = int_reg_array_34_45_imag;
        _zz_4503_ = int_reg_array_34_45_real;
      end
      6'b101110 : begin
        _zz_4502_ = int_reg_array_34_46_imag;
        _zz_4503_ = int_reg_array_34_46_real;
      end
      6'b101111 : begin
        _zz_4502_ = int_reg_array_34_47_imag;
        _zz_4503_ = int_reg_array_34_47_real;
      end
      6'b110000 : begin
        _zz_4502_ = int_reg_array_34_48_imag;
        _zz_4503_ = int_reg_array_34_48_real;
      end
      6'b110001 : begin
        _zz_4502_ = int_reg_array_34_49_imag;
        _zz_4503_ = int_reg_array_34_49_real;
      end
      6'b110010 : begin
        _zz_4502_ = int_reg_array_34_50_imag;
        _zz_4503_ = int_reg_array_34_50_real;
      end
      6'b110011 : begin
        _zz_4502_ = int_reg_array_34_51_imag;
        _zz_4503_ = int_reg_array_34_51_real;
      end
      6'b110100 : begin
        _zz_4502_ = int_reg_array_34_52_imag;
        _zz_4503_ = int_reg_array_34_52_real;
      end
      6'b110101 : begin
        _zz_4502_ = int_reg_array_34_53_imag;
        _zz_4503_ = int_reg_array_34_53_real;
      end
      6'b110110 : begin
        _zz_4502_ = int_reg_array_34_54_imag;
        _zz_4503_ = int_reg_array_34_54_real;
      end
      6'b110111 : begin
        _zz_4502_ = int_reg_array_34_55_imag;
        _zz_4503_ = int_reg_array_34_55_real;
      end
      6'b111000 : begin
        _zz_4502_ = int_reg_array_34_56_imag;
        _zz_4503_ = int_reg_array_34_56_real;
      end
      6'b111001 : begin
        _zz_4502_ = int_reg_array_34_57_imag;
        _zz_4503_ = int_reg_array_34_57_real;
      end
      6'b111010 : begin
        _zz_4502_ = int_reg_array_34_58_imag;
        _zz_4503_ = int_reg_array_34_58_real;
      end
      6'b111011 : begin
        _zz_4502_ = int_reg_array_34_59_imag;
        _zz_4503_ = int_reg_array_34_59_real;
      end
      6'b111100 : begin
        _zz_4502_ = int_reg_array_34_60_imag;
        _zz_4503_ = int_reg_array_34_60_real;
      end
      6'b111101 : begin
        _zz_4502_ = int_reg_array_34_61_imag;
        _zz_4503_ = int_reg_array_34_61_real;
      end
      6'b111110 : begin
        _zz_4502_ = int_reg_array_34_62_imag;
        _zz_4503_ = int_reg_array_34_62_real;
      end
      default : begin
        _zz_4502_ = int_reg_array_34_63_imag;
        _zz_4503_ = int_reg_array_34_63_real;
      end
    endcase
  end

  always @(*) begin
    case(_zz_2432_)
      6'b000000 : begin
        _zz_4504_ = int_reg_array_35_0_imag;
        _zz_4505_ = int_reg_array_35_0_real;
      end
      6'b000001 : begin
        _zz_4504_ = int_reg_array_35_1_imag;
        _zz_4505_ = int_reg_array_35_1_real;
      end
      6'b000010 : begin
        _zz_4504_ = int_reg_array_35_2_imag;
        _zz_4505_ = int_reg_array_35_2_real;
      end
      6'b000011 : begin
        _zz_4504_ = int_reg_array_35_3_imag;
        _zz_4505_ = int_reg_array_35_3_real;
      end
      6'b000100 : begin
        _zz_4504_ = int_reg_array_35_4_imag;
        _zz_4505_ = int_reg_array_35_4_real;
      end
      6'b000101 : begin
        _zz_4504_ = int_reg_array_35_5_imag;
        _zz_4505_ = int_reg_array_35_5_real;
      end
      6'b000110 : begin
        _zz_4504_ = int_reg_array_35_6_imag;
        _zz_4505_ = int_reg_array_35_6_real;
      end
      6'b000111 : begin
        _zz_4504_ = int_reg_array_35_7_imag;
        _zz_4505_ = int_reg_array_35_7_real;
      end
      6'b001000 : begin
        _zz_4504_ = int_reg_array_35_8_imag;
        _zz_4505_ = int_reg_array_35_8_real;
      end
      6'b001001 : begin
        _zz_4504_ = int_reg_array_35_9_imag;
        _zz_4505_ = int_reg_array_35_9_real;
      end
      6'b001010 : begin
        _zz_4504_ = int_reg_array_35_10_imag;
        _zz_4505_ = int_reg_array_35_10_real;
      end
      6'b001011 : begin
        _zz_4504_ = int_reg_array_35_11_imag;
        _zz_4505_ = int_reg_array_35_11_real;
      end
      6'b001100 : begin
        _zz_4504_ = int_reg_array_35_12_imag;
        _zz_4505_ = int_reg_array_35_12_real;
      end
      6'b001101 : begin
        _zz_4504_ = int_reg_array_35_13_imag;
        _zz_4505_ = int_reg_array_35_13_real;
      end
      6'b001110 : begin
        _zz_4504_ = int_reg_array_35_14_imag;
        _zz_4505_ = int_reg_array_35_14_real;
      end
      6'b001111 : begin
        _zz_4504_ = int_reg_array_35_15_imag;
        _zz_4505_ = int_reg_array_35_15_real;
      end
      6'b010000 : begin
        _zz_4504_ = int_reg_array_35_16_imag;
        _zz_4505_ = int_reg_array_35_16_real;
      end
      6'b010001 : begin
        _zz_4504_ = int_reg_array_35_17_imag;
        _zz_4505_ = int_reg_array_35_17_real;
      end
      6'b010010 : begin
        _zz_4504_ = int_reg_array_35_18_imag;
        _zz_4505_ = int_reg_array_35_18_real;
      end
      6'b010011 : begin
        _zz_4504_ = int_reg_array_35_19_imag;
        _zz_4505_ = int_reg_array_35_19_real;
      end
      6'b010100 : begin
        _zz_4504_ = int_reg_array_35_20_imag;
        _zz_4505_ = int_reg_array_35_20_real;
      end
      6'b010101 : begin
        _zz_4504_ = int_reg_array_35_21_imag;
        _zz_4505_ = int_reg_array_35_21_real;
      end
      6'b010110 : begin
        _zz_4504_ = int_reg_array_35_22_imag;
        _zz_4505_ = int_reg_array_35_22_real;
      end
      6'b010111 : begin
        _zz_4504_ = int_reg_array_35_23_imag;
        _zz_4505_ = int_reg_array_35_23_real;
      end
      6'b011000 : begin
        _zz_4504_ = int_reg_array_35_24_imag;
        _zz_4505_ = int_reg_array_35_24_real;
      end
      6'b011001 : begin
        _zz_4504_ = int_reg_array_35_25_imag;
        _zz_4505_ = int_reg_array_35_25_real;
      end
      6'b011010 : begin
        _zz_4504_ = int_reg_array_35_26_imag;
        _zz_4505_ = int_reg_array_35_26_real;
      end
      6'b011011 : begin
        _zz_4504_ = int_reg_array_35_27_imag;
        _zz_4505_ = int_reg_array_35_27_real;
      end
      6'b011100 : begin
        _zz_4504_ = int_reg_array_35_28_imag;
        _zz_4505_ = int_reg_array_35_28_real;
      end
      6'b011101 : begin
        _zz_4504_ = int_reg_array_35_29_imag;
        _zz_4505_ = int_reg_array_35_29_real;
      end
      6'b011110 : begin
        _zz_4504_ = int_reg_array_35_30_imag;
        _zz_4505_ = int_reg_array_35_30_real;
      end
      6'b011111 : begin
        _zz_4504_ = int_reg_array_35_31_imag;
        _zz_4505_ = int_reg_array_35_31_real;
      end
      6'b100000 : begin
        _zz_4504_ = int_reg_array_35_32_imag;
        _zz_4505_ = int_reg_array_35_32_real;
      end
      6'b100001 : begin
        _zz_4504_ = int_reg_array_35_33_imag;
        _zz_4505_ = int_reg_array_35_33_real;
      end
      6'b100010 : begin
        _zz_4504_ = int_reg_array_35_34_imag;
        _zz_4505_ = int_reg_array_35_34_real;
      end
      6'b100011 : begin
        _zz_4504_ = int_reg_array_35_35_imag;
        _zz_4505_ = int_reg_array_35_35_real;
      end
      6'b100100 : begin
        _zz_4504_ = int_reg_array_35_36_imag;
        _zz_4505_ = int_reg_array_35_36_real;
      end
      6'b100101 : begin
        _zz_4504_ = int_reg_array_35_37_imag;
        _zz_4505_ = int_reg_array_35_37_real;
      end
      6'b100110 : begin
        _zz_4504_ = int_reg_array_35_38_imag;
        _zz_4505_ = int_reg_array_35_38_real;
      end
      6'b100111 : begin
        _zz_4504_ = int_reg_array_35_39_imag;
        _zz_4505_ = int_reg_array_35_39_real;
      end
      6'b101000 : begin
        _zz_4504_ = int_reg_array_35_40_imag;
        _zz_4505_ = int_reg_array_35_40_real;
      end
      6'b101001 : begin
        _zz_4504_ = int_reg_array_35_41_imag;
        _zz_4505_ = int_reg_array_35_41_real;
      end
      6'b101010 : begin
        _zz_4504_ = int_reg_array_35_42_imag;
        _zz_4505_ = int_reg_array_35_42_real;
      end
      6'b101011 : begin
        _zz_4504_ = int_reg_array_35_43_imag;
        _zz_4505_ = int_reg_array_35_43_real;
      end
      6'b101100 : begin
        _zz_4504_ = int_reg_array_35_44_imag;
        _zz_4505_ = int_reg_array_35_44_real;
      end
      6'b101101 : begin
        _zz_4504_ = int_reg_array_35_45_imag;
        _zz_4505_ = int_reg_array_35_45_real;
      end
      6'b101110 : begin
        _zz_4504_ = int_reg_array_35_46_imag;
        _zz_4505_ = int_reg_array_35_46_real;
      end
      6'b101111 : begin
        _zz_4504_ = int_reg_array_35_47_imag;
        _zz_4505_ = int_reg_array_35_47_real;
      end
      6'b110000 : begin
        _zz_4504_ = int_reg_array_35_48_imag;
        _zz_4505_ = int_reg_array_35_48_real;
      end
      6'b110001 : begin
        _zz_4504_ = int_reg_array_35_49_imag;
        _zz_4505_ = int_reg_array_35_49_real;
      end
      6'b110010 : begin
        _zz_4504_ = int_reg_array_35_50_imag;
        _zz_4505_ = int_reg_array_35_50_real;
      end
      6'b110011 : begin
        _zz_4504_ = int_reg_array_35_51_imag;
        _zz_4505_ = int_reg_array_35_51_real;
      end
      6'b110100 : begin
        _zz_4504_ = int_reg_array_35_52_imag;
        _zz_4505_ = int_reg_array_35_52_real;
      end
      6'b110101 : begin
        _zz_4504_ = int_reg_array_35_53_imag;
        _zz_4505_ = int_reg_array_35_53_real;
      end
      6'b110110 : begin
        _zz_4504_ = int_reg_array_35_54_imag;
        _zz_4505_ = int_reg_array_35_54_real;
      end
      6'b110111 : begin
        _zz_4504_ = int_reg_array_35_55_imag;
        _zz_4505_ = int_reg_array_35_55_real;
      end
      6'b111000 : begin
        _zz_4504_ = int_reg_array_35_56_imag;
        _zz_4505_ = int_reg_array_35_56_real;
      end
      6'b111001 : begin
        _zz_4504_ = int_reg_array_35_57_imag;
        _zz_4505_ = int_reg_array_35_57_real;
      end
      6'b111010 : begin
        _zz_4504_ = int_reg_array_35_58_imag;
        _zz_4505_ = int_reg_array_35_58_real;
      end
      6'b111011 : begin
        _zz_4504_ = int_reg_array_35_59_imag;
        _zz_4505_ = int_reg_array_35_59_real;
      end
      6'b111100 : begin
        _zz_4504_ = int_reg_array_35_60_imag;
        _zz_4505_ = int_reg_array_35_60_real;
      end
      6'b111101 : begin
        _zz_4504_ = int_reg_array_35_61_imag;
        _zz_4505_ = int_reg_array_35_61_real;
      end
      6'b111110 : begin
        _zz_4504_ = int_reg_array_35_62_imag;
        _zz_4505_ = int_reg_array_35_62_real;
      end
      default : begin
        _zz_4504_ = int_reg_array_35_63_imag;
        _zz_4505_ = int_reg_array_35_63_real;
      end
    endcase
  end

  always @(*) begin
    case(_zz_2501_)
      6'b000000 : begin
        _zz_4506_ = int_reg_array_36_0_imag;
        _zz_4507_ = int_reg_array_36_0_real;
      end
      6'b000001 : begin
        _zz_4506_ = int_reg_array_36_1_imag;
        _zz_4507_ = int_reg_array_36_1_real;
      end
      6'b000010 : begin
        _zz_4506_ = int_reg_array_36_2_imag;
        _zz_4507_ = int_reg_array_36_2_real;
      end
      6'b000011 : begin
        _zz_4506_ = int_reg_array_36_3_imag;
        _zz_4507_ = int_reg_array_36_3_real;
      end
      6'b000100 : begin
        _zz_4506_ = int_reg_array_36_4_imag;
        _zz_4507_ = int_reg_array_36_4_real;
      end
      6'b000101 : begin
        _zz_4506_ = int_reg_array_36_5_imag;
        _zz_4507_ = int_reg_array_36_5_real;
      end
      6'b000110 : begin
        _zz_4506_ = int_reg_array_36_6_imag;
        _zz_4507_ = int_reg_array_36_6_real;
      end
      6'b000111 : begin
        _zz_4506_ = int_reg_array_36_7_imag;
        _zz_4507_ = int_reg_array_36_7_real;
      end
      6'b001000 : begin
        _zz_4506_ = int_reg_array_36_8_imag;
        _zz_4507_ = int_reg_array_36_8_real;
      end
      6'b001001 : begin
        _zz_4506_ = int_reg_array_36_9_imag;
        _zz_4507_ = int_reg_array_36_9_real;
      end
      6'b001010 : begin
        _zz_4506_ = int_reg_array_36_10_imag;
        _zz_4507_ = int_reg_array_36_10_real;
      end
      6'b001011 : begin
        _zz_4506_ = int_reg_array_36_11_imag;
        _zz_4507_ = int_reg_array_36_11_real;
      end
      6'b001100 : begin
        _zz_4506_ = int_reg_array_36_12_imag;
        _zz_4507_ = int_reg_array_36_12_real;
      end
      6'b001101 : begin
        _zz_4506_ = int_reg_array_36_13_imag;
        _zz_4507_ = int_reg_array_36_13_real;
      end
      6'b001110 : begin
        _zz_4506_ = int_reg_array_36_14_imag;
        _zz_4507_ = int_reg_array_36_14_real;
      end
      6'b001111 : begin
        _zz_4506_ = int_reg_array_36_15_imag;
        _zz_4507_ = int_reg_array_36_15_real;
      end
      6'b010000 : begin
        _zz_4506_ = int_reg_array_36_16_imag;
        _zz_4507_ = int_reg_array_36_16_real;
      end
      6'b010001 : begin
        _zz_4506_ = int_reg_array_36_17_imag;
        _zz_4507_ = int_reg_array_36_17_real;
      end
      6'b010010 : begin
        _zz_4506_ = int_reg_array_36_18_imag;
        _zz_4507_ = int_reg_array_36_18_real;
      end
      6'b010011 : begin
        _zz_4506_ = int_reg_array_36_19_imag;
        _zz_4507_ = int_reg_array_36_19_real;
      end
      6'b010100 : begin
        _zz_4506_ = int_reg_array_36_20_imag;
        _zz_4507_ = int_reg_array_36_20_real;
      end
      6'b010101 : begin
        _zz_4506_ = int_reg_array_36_21_imag;
        _zz_4507_ = int_reg_array_36_21_real;
      end
      6'b010110 : begin
        _zz_4506_ = int_reg_array_36_22_imag;
        _zz_4507_ = int_reg_array_36_22_real;
      end
      6'b010111 : begin
        _zz_4506_ = int_reg_array_36_23_imag;
        _zz_4507_ = int_reg_array_36_23_real;
      end
      6'b011000 : begin
        _zz_4506_ = int_reg_array_36_24_imag;
        _zz_4507_ = int_reg_array_36_24_real;
      end
      6'b011001 : begin
        _zz_4506_ = int_reg_array_36_25_imag;
        _zz_4507_ = int_reg_array_36_25_real;
      end
      6'b011010 : begin
        _zz_4506_ = int_reg_array_36_26_imag;
        _zz_4507_ = int_reg_array_36_26_real;
      end
      6'b011011 : begin
        _zz_4506_ = int_reg_array_36_27_imag;
        _zz_4507_ = int_reg_array_36_27_real;
      end
      6'b011100 : begin
        _zz_4506_ = int_reg_array_36_28_imag;
        _zz_4507_ = int_reg_array_36_28_real;
      end
      6'b011101 : begin
        _zz_4506_ = int_reg_array_36_29_imag;
        _zz_4507_ = int_reg_array_36_29_real;
      end
      6'b011110 : begin
        _zz_4506_ = int_reg_array_36_30_imag;
        _zz_4507_ = int_reg_array_36_30_real;
      end
      6'b011111 : begin
        _zz_4506_ = int_reg_array_36_31_imag;
        _zz_4507_ = int_reg_array_36_31_real;
      end
      6'b100000 : begin
        _zz_4506_ = int_reg_array_36_32_imag;
        _zz_4507_ = int_reg_array_36_32_real;
      end
      6'b100001 : begin
        _zz_4506_ = int_reg_array_36_33_imag;
        _zz_4507_ = int_reg_array_36_33_real;
      end
      6'b100010 : begin
        _zz_4506_ = int_reg_array_36_34_imag;
        _zz_4507_ = int_reg_array_36_34_real;
      end
      6'b100011 : begin
        _zz_4506_ = int_reg_array_36_35_imag;
        _zz_4507_ = int_reg_array_36_35_real;
      end
      6'b100100 : begin
        _zz_4506_ = int_reg_array_36_36_imag;
        _zz_4507_ = int_reg_array_36_36_real;
      end
      6'b100101 : begin
        _zz_4506_ = int_reg_array_36_37_imag;
        _zz_4507_ = int_reg_array_36_37_real;
      end
      6'b100110 : begin
        _zz_4506_ = int_reg_array_36_38_imag;
        _zz_4507_ = int_reg_array_36_38_real;
      end
      6'b100111 : begin
        _zz_4506_ = int_reg_array_36_39_imag;
        _zz_4507_ = int_reg_array_36_39_real;
      end
      6'b101000 : begin
        _zz_4506_ = int_reg_array_36_40_imag;
        _zz_4507_ = int_reg_array_36_40_real;
      end
      6'b101001 : begin
        _zz_4506_ = int_reg_array_36_41_imag;
        _zz_4507_ = int_reg_array_36_41_real;
      end
      6'b101010 : begin
        _zz_4506_ = int_reg_array_36_42_imag;
        _zz_4507_ = int_reg_array_36_42_real;
      end
      6'b101011 : begin
        _zz_4506_ = int_reg_array_36_43_imag;
        _zz_4507_ = int_reg_array_36_43_real;
      end
      6'b101100 : begin
        _zz_4506_ = int_reg_array_36_44_imag;
        _zz_4507_ = int_reg_array_36_44_real;
      end
      6'b101101 : begin
        _zz_4506_ = int_reg_array_36_45_imag;
        _zz_4507_ = int_reg_array_36_45_real;
      end
      6'b101110 : begin
        _zz_4506_ = int_reg_array_36_46_imag;
        _zz_4507_ = int_reg_array_36_46_real;
      end
      6'b101111 : begin
        _zz_4506_ = int_reg_array_36_47_imag;
        _zz_4507_ = int_reg_array_36_47_real;
      end
      6'b110000 : begin
        _zz_4506_ = int_reg_array_36_48_imag;
        _zz_4507_ = int_reg_array_36_48_real;
      end
      6'b110001 : begin
        _zz_4506_ = int_reg_array_36_49_imag;
        _zz_4507_ = int_reg_array_36_49_real;
      end
      6'b110010 : begin
        _zz_4506_ = int_reg_array_36_50_imag;
        _zz_4507_ = int_reg_array_36_50_real;
      end
      6'b110011 : begin
        _zz_4506_ = int_reg_array_36_51_imag;
        _zz_4507_ = int_reg_array_36_51_real;
      end
      6'b110100 : begin
        _zz_4506_ = int_reg_array_36_52_imag;
        _zz_4507_ = int_reg_array_36_52_real;
      end
      6'b110101 : begin
        _zz_4506_ = int_reg_array_36_53_imag;
        _zz_4507_ = int_reg_array_36_53_real;
      end
      6'b110110 : begin
        _zz_4506_ = int_reg_array_36_54_imag;
        _zz_4507_ = int_reg_array_36_54_real;
      end
      6'b110111 : begin
        _zz_4506_ = int_reg_array_36_55_imag;
        _zz_4507_ = int_reg_array_36_55_real;
      end
      6'b111000 : begin
        _zz_4506_ = int_reg_array_36_56_imag;
        _zz_4507_ = int_reg_array_36_56_real;
      end
      6'b111001 : begin
        _zz_4506_ = int_reg_array_36_57_imag;
        _zz_4507_ = int_reg_array_36_57_real;
      end
      6'b111010 : begin
        _zz_4506_ = int_reg_array_36_58_imag;
        _zz_4507_ = int_reg_array_36_58_real;
      end
      6'b111011 : begin
        _zz_4506_ = int_reg_array_36_59_imag;
        _zz_4507_ = int_reg_array_36_59_real;
      end
      6'b111100 : begin
        _zz_4506_ = int_reg_array_36_60_imag;
        _zz_4507_ = int_reg_array_36_60_real;
      end
      6'b111101 : begin
        _zz_4506_ = int_reg_array_36_61_imag;
        _zz_4507_ = int_reg_array_36_61_real;
      end
      6'b111110 : begin
        _zz_4506_ = int_reg_array_36_62_imag;
        _zz_4507_ = int_reg_array_36_62_real;
      end
      default : begin
        _zz_4506_ = int_reg_array_36_63_imag;
        _zz_4507_ = int_reg_array_36_63_real;
      end
    endcase
  end

  always @(*) begin
    case(_zz_2570_)
      6'b000000 : begin
        _zz_4508_ = int_reg_array_37_0_imag;
        _zz_4509_ = int_reg_array_37_0_real;
      end
      6'b000001 : begin
        _zz_4508_ = int_reg_array_37_1_imag;
        _zz_4509_ = int_reg_array_37_1_real;
      end
      6'b000010 : begin
        _zz_4508_ = int_reg_array_37_2_imag;
        _zz_4509_ = int_reg_array_37_2_real;
      end
      6'b000011 : begin
        _zz_4508_ = int_reg_array_37_3_imag;
        _zz_4509_ = int_reg_array_37_3_real;
      end
      6'b000100 : begin
        _zz_4508_ = int_reg_array_37_4_imag;
        _zz_4509_ = int_reg_array_37_4_real;
      end
      6'b000101 : begin
        _zz_4508_ = int_reg_array_37_5_imag;
        _zz_4509_ = int_reg_array_37_5_real;
      end
      6'b000110 : begin
        _zz_4508_ = int_reg_array_37_6_imag;
        _zz_4509_ = int_reg_array_37_6_real;
      end
      6'b000111 : begin
        _zz_4508_ = int_reg_array_37_7_imag;
        _zz_4509_ = int_reg_array_37_7_real;
      end
      6'b001000 : begin
        _zz_4508_ = int_reg_array_37_8_imag;
        _zz_4509_ = int_reg_array_37_8_real;
      end
      6'b001001 : begin
        _zz_4508_ = int_reg_array_37_9_imag;
        _zz_4509_ = int_reg_array_37_9_real;
      end
      6'b001010 : begin
        _zz_4508_ = int_reg_array_37_10_imag;
        _zz_4509_ = int_reg_array_37_10_real;
      end
      6'b001011 : begin
        _zz_4508_ = int_reg_array_37_11_imag;
        _zz_4509_ = int_reg_array_37_11_real;
      end
      6'b001100 : begin
        _zz_4508_ = int_reg_array_37_12_imag;
        _zz_4509_ = int_reg_array_37_12_real;
      end
      6'b001101 : begin
        _zz_4508_ = int_reg_array_37_13_imag;
        _zz_4509_ = int_reg_array_37_13_real;
      end
      6'b001110 : begin
        _zz_4508_ = int_reg_array_37_14_imag;
        _zz_4509_ = int_reg_array_37_14_real;
      end
      6'b001111 : begin
        _zz_4508_ = int_reg_array_37_15_imag;
        _zz_4509_ = int_reg_array_37_15_real;
      end
      6'b010000 : begin
        _zz_4508_ = int_reg_array_37_16_imag;
        _zz_4509_ = int_reg_array_37_16_real;
      end
      6'b010001 : begin
        _zz_4508_ = int_reg_array_37_17_imag;
        _zz_4509_ = int_reg_array_37_17_real;
      end
      6'b010010 : begin
        _zz_4508_ = int_reg_array_37_18_imag;
        _zz_4509_ = int_reg_array_37_18_real;
      end
      6'b010011 : begin
        _zz_4508_ = int_reg_array_37_19_imag;
        _zz_4509_ = int_reg_array_37_19_real;
      end
      6'b010100 : begin
        _zz_4508_ = int_reg_array_37_20_imag;
        _zz_4509_ = int_reg_array_37_20_real;
      end
      6'b010101 : begin
        _zz_4508_ = int_reg_array_37_21_imag;
        _zz_4509_ = int_reg_array_37_21_real;
      end
      6'b010110 : begin
        _zz_4508_ = int_reg_array_37_22_imag;
        _zz_4509_ = int_reg_array_37_22_real;
      end
      6'b010111 : begin
        _zz_4508_ = int_reg_array_37_23_imag;
        _zz_4509_ = int_reg_array_37_23_real;
      end
      6'b011000 : begin
        _zz_4508_ = int_reg_array_37_24_imag;
        _zz_4509_ = int_reg_array_37_24_real;
      end
      6'b011001 : begin
        _zz_4508_ = int_reg_array_37_25_imag;
        _zz_4509_ = int_reg_array_37_25_real;
      end
      6'b011010 : begin
        _zz_4508_ = int_reg_array_37_26_imag;
        _zz_4509_ = int_reg_array_37_26_real;
      end
      6'b011011 : begin
        _zz_4508_ = int_reg_array_37_27_imag;
        _zz_4509_ = int_reg_array_37_27_real;
      end
      6'b011100 : begin
        _zz_4508_ = int_reg_array_37_28_imag;
        _zz_4509_ = int_reg_array_37_28_real;
      end
      6'b011101 : begin
        _zz_4508_ = int_reg_array_37_29_imag;
        _zz_4509_ = int_reg_array_37_29_real;
      end
      6'b011110 : begin
        _zz_4508_ = int_reg_array_37_30_imag;
        _zz_4509_ = int_reg_array_37_30_real;
      end
      6'b011111 : begin
        _zz_4508_ = int_reg_array_37_31_imag;
        _zz_4509_ = int_reg_array_37_31_real;
      end
      6'b100000 : begin
        _zz_4508_ = int_reg_array_37_32_imag;
        _zz_4509_ = int_reg_array_37_32_real;
      end
      6'b100001 : begin
        _zz_4508_ = int_reg_array_37_33_imag;
        _zz_4509_ = int_reg_array_37_33_real;
      end
      6'b100010 : begin
        _zz_4508_ = int_reg_array_37_34_imag;
        _zz_4509_ = int_reg_array_37_34_real;
      end
      6'b100011 : begin
        _zz_4508_ = int_reg_array_37_35_imag;
        _zz_4509_ = int_reg_array_37_35_real;
      end
      6'b100100 : begin
        _zz_4508_ = int_reg_array_37_36_imag;
        _zz_4509_ = int_reg_array_37_36_real;
      end
      6'b100101 : begin
        _zz_4508_ = int_reg_array_37_37_imag;
        _zz_4509_ = int_reg_array_37_37_real;
      end
      6'b100110 : begin
        _zz_4508_ = int_reg_array_37_38_imag;
        _zz_4509_ = int_reg_array_37_38_real;
      end
      6'b100111 : begin
        _zz_4508_ = int_reg_array_37_39_imag;
        _zz_4509_ = int_reg_array_37_39_real;
      end
      6'b101000 : begin
        _zz_4508_ = int_reg_array_37_40_imag;
        _zz_4509_ = int_reg_array_37_40_real;
      end
      6'b101001 : begin
        _zz_4508_ = int_reg_array_37_41_imag;
        _zz_4509_ = int_reg_array_37_41_real;
      end
      6'b101010 : begin
        _zz_4508_ = int_reg_array_37_42_imag;
        _zz_4509_ = int_reg_array_37_42_real;
      end
      6'b101011 : begin
        _zz_4508_ = int_reg_array_37_43_imag;
        _zz_4509_ = int_reg_array_37_43_real;
      end
      6'b101100 : begin
        _zz_4508_ = int_reg_array_37_44_imag;
        _zz_4509_ = int_reg_array_37_44_real;
      end
      6'b101101 : begin
        _zz_4508_ = int_reg_array_37_45_imag;
        _zz_4509_ = int_reg_array_37_45_real;
      end
      6'b101110 : begin
        _zz_4508_ = int_reg_array_37_46_imag;
        _zz_4509_ = int_reg_array_37_46_real;
      end
      6'b101111 : begin
        _zz_4508_ = int_reg_array_37_47_imag;
        _zz_4509_ = int_reg_array_37_47_real;
      end
      6'b110000 : begin
        _zz_4508_ = int_reg_array_37_48_imag;
        _zz_4509_ = int_reg_array_37_48_real;
      end
      6'b110001 : begin
        _zz_4508_ = int_reg_array_37_49_imag;
        _zz_4509_ = int_reg_array_37_49_real;
      end
      6'b110010 : begin
        _zz_4508_ = int_reg_array_37_50_imag;
        _zz_4509_ = int_reg_array_37_50_real;
      end
      6'b110011 : begin
        _zz_4508_ = int_reg_array_37_51_imag;
        _zz_4509_ = int_reg_array_37_51_real;
      end
      6'b110100 : begin
        _zz_4508_ = int_reg_array_37_52_imag;
        _zz_4509_ = int_reg_array_37_52_real;
      end
      6'b110101 : begin
        _zz_4508_ = int_reg_array_37_53_imag;
        _zz_4509_ = int_reg_array_37_53_real;
      end
      6'b110110 : begin
        _zz_4508_ = int_reg_array_37_54_imag;
        _zz_4509_ = int_reg_array_37_54_real;
      end
      6'b110111 : begin
        _zz_4508_ = int_reg_array_37_55_imag;
        _zz_4509_ = int_reg_array_37_55_real;
      end
      6'b111000 : begin
        _zz_4508_ = int_reg_array_37_56_imag;
        _zz_4509_ = int_reg_array_37_56_real;
      end
      6'b111001 : begin
        _zz_4508_ = int_reg_array_37_57_imag;
        _zz_4509_ = int_reg_array_37_57_real;
      end
      6'b111010 : begin
        _zz_4508_ = int_reg_array_37_58_imag;
        _zz_4509_ = int_reg_array_37_58_real;
      end
      6'b111011 : begin
        _zz_4508_ = int_reg_array_37_59_imag;
        _zz_4509_ = int_reg_array_37_59_real;
      end
      6'b111100 : begin
        _zz_4508_ = int_reg_array_37_60_imag;
        _zz_4509_ = int_reg_array_37_60_real;
      end
      6'b111101 : begin
        _zz_4508_ = int_reg_array_37_61_imag;
        _zz_4509_ = int_reg_array_37_61_real;
      end
      6'b111110 : begin
        _zz_4508_ = int_reg_array_37_62_imag;
        _zz_4509_ = int_reg_array_37_62_real;
      end
      default : begin
        _zz_4508_ = int_reg_array_37_63_imag;
        _zz_4509_ = int_reg_array_37_63_real;
      end
    endcase
  end

  always @(*) begin
    case(_zz_2639_)
      6'b000000 : begin
        _zz_4510_ = int_reg_array_38_0_imag;
        _zz_4511_ = int_reg_array_38_0_real;
      end
      6'b000001 : begin
        _zz_4510_ = int_reg_array_38_1_imag;
        _zz_4511_ = int_reg_array_38_1_real;
      end
      6'b000010 : begin
        _zz_4510_ = int_reg_array_38_2_imag;
        _zz_4511_ = int_reg_array_38_2_real;
      end
      6'b000011 : begin
        _zz_4510_ = int_reg_array_38_3_imag;
        _zz_4511_ = int_reg_array_38_3_real;
      end
      6'b000100 : begin
        _zz_4510_ = int_reg_array_38_4_imag;
        _zz_4511_ = int_reg_array_38_4_real;
      end
      6'b000101 : begin
        _zz_4510_ = int_reg_array_38_5_imag;
        _zz_4511_ = int_reg_array_38_5_real;
      end
      6'b000110 : begin
        _zz_4510_ = int_reg_array_38_6_imag;
        _zz_4511_ = int_reg_array_38_6_real;
      end
      6'b000111 : begin
        _zz_4510_ = int_reg_array_38_7_imag;
        _zz_4511_ = int_reg_array_38_7_real;
      end
      6'b001000 : begin
        _zz_4510_ = int_reg_array_38_8_imag;
        _zz_4511_ = int_reg_array_38_8_real;
      end
      6'b001001 : begin
        _zz_4510_ = int_reg_array_38_9_imag;
        _zz_4511_ = int_reg_array_38_9_real;
      end
      6'b001010 : begin
        _zz_4510_ = int_reg_array_38_10_imag;
        _zz_4511_ = int_reg_array_38_10_real;
      end
      6'b001011 : begin
        _zz_4510_ = int_reg_array_38_11_imag;
        _zz_4511_ = int_reg_array_38_11_real;
      end
      6'b001100 : begin
        _zz_4510_ = int_reg_array_38_12_imag;
        _zz_4511_ = int_reg_array_38_12_real;
      end
      6'b001101 : begin
        _zz_4510_ = int_reg_array_38_13_imag;
        _zz_4511_ = int_reg_array_38_13_real;
      end
      6'b001110 : begin
        _zz_4510_ = int_reg_array_38_14_imag;
        _zz_4511_ = int_reg_array_38_14_real;
      end
      6'b001111 : begin
        _zz_4510_ = int_reg_array_38_15_imag;
        _zz_4511_ = int_reg_array_38_15_real;
      end
      6'b010000 : begin
        _zz_4510_ = int_reg_array_38_16_imag;
        _zz_4511_ = int_reg_array_38_16_real;
      end
      6'b010001 : begin
        _zz_4510_ = int_reg_array_38_17_imag;
        _zz_4511_ = int_reg_array_38_17_real;
      end
      6'b010010 : begin
        _zz_4510_ = int_reg_array_38_18_imag;
        _zz_4511_ = int_reg_array_38_18_real;
      end
      6'b010011 : begin
        _zz_4510_ = int_reg_array_38_19_imag;
        _zz_4511_ = int_reg_array_38_19_real;
      end
      6'b010100 : begin
        _zz_4510_ = int_reg_array_38_20_imag;
        _zz_4511_ = int_reg_array_38_20_real;
      end
      6'b010101 : begin
        _zz_4510_ = int_reg_array_38_21_imag;
        _zz_4511_ = int_reg_array_38_21_real;
      end
      6'b010110 : begin
        _zz_4510_ = int_reg_array_38_22_imag;
        _zz_4511_ = int_reg_array_38_22_real;
      end
      6'b010111 : begin
        _zz_4510_ = int_reg_array_38_23_imag;
        _zz_4511_ = int_reg_array_38_23_real;
      end
      6'b011000 : begin
        _zz_4510_ = int_reg_array_38_24_imag;
        _zz_4511_ = int_reg_array_38_24_real;
      end
      6'b011001 : begin
        _zz_4510_ = int_reg_array_38_25_imag;
        _zz_4511_ = int_reg_array_38_25_real;
      end
      6'b011010 : begin
        _zz_4510_ = int_reg_array_38_26_imag;
        _zz_4511_ = int_reg_array_38_26_real;
      end
      6'b011011 : begin
        _zz_4510_ = int_reg_array_38_27_imag;
        _zz_4511_ = int_reg_array_38_27_real;
      end
      6'b011100 : begin
        _zz_4510_ = int_reg_array_38_28_imag;
        _zz_4511_ = int_reg_array_38_28_real;
      end
      6'b011101 : begin
        _zz_4510_ = int_reg_array_38_29_imag;
        _zz_4511_ = int_reg_array_38_29_real;
      end
      6'b011110 : begin
        _zz_4510_ = int_reg_array_38_30_imag;
        _zz_4511_ = int_reg_array_38_30_real;
      end
      6'b011111 : begin
        _zz_4510_ = int_reg_array_38_31_imag;
        _zz_4511_ = int_reg_array_38_31_real;
      end
      6'b100000 : begin
        _zz_4510_ = int_reg_array_38_32_imag;
        _zz_4511_ = int_reg_array_38_32_real;
      end
      6'b100001 : begin
        _zz_4510_ = int_reg_array_38_33_imag;
        _zz_4511_ = int_reg_array_38_33_real;
      end
      6'b100010 : begin
        _zz_4510_ = int_reg_array_38_34_imag;
        _zz_4511_ = int_reg_array_38_34_real;
      end
      6'b100011 : begin
        _zz_4510_ = int_reg_array_38_35_imag;
        _zz_4511_ = int_reg_array_38_35_real;
      end
      6'b100100 : begin
        _zz_4510_ = int_reg_array_38_36_imag;
        _zz_4511_ = int_reg_array_38_36_real;
      end
      6'b100101 : begin
        _zz_4510_ = int_reg_array_38_37_imag;
        _zz_4511_ = int_reg_array_38_37_real;
      end
      6'b100110 : begin
        _zz_4510_ = int_reg_array_38_38_imag;
        _zz_4511_ = int_reg_array_38_38_real;
      end
      6'b100111 : begin
        _zz_4510_ = int_reg_array_38_39_imag;
        _zz_4511_ = int_reg_array_38_39_real;
      end
      6'b101000 : begin
        _zz_4510_ = int_reg_array_38_40_imag;
        _zz_4511_ = int_reg_array_38_40_real;
      end
      6'b101001 : begin
        _zz_4510_ = int_reg_array_38_41_imag;
        _zz_4511_ = int_reg_array_38_41_real;
      end
      6'b101010 : begin
        _zz_4510_ = int_reg_array_38_42_imag;
        _zz_4511_ = int_reg_array_38_42_real;
      end
      6'b101011 : begin
        _zz_4510_ = int_reg_array_38_43_imag;
        _zz_4511_ = int_reg_array_38_43_real;
      end
      6'b101100 : begin
        _zz_4510_ = int_reg_array_38_44_imag;
        _zz_4511_ = int_reg_array_38_44_real;
      end
      6'b101101 : begin
        _zz_4510_ = int_reg_array_38_45_imag;
        _zz_4511_ = int_reg_array_38_45_real;
      end
      6'b101110 : begin
        _zz_4510_ = int_reg_array_38_46_imag;
        _zz_4511_ = int_reg_array_38_46_real;
      end
      6'b101111 : begin
        _zz_4510_ = int_reg_array_38_47_imag;
        _zz_4511_ = int_reg_array_38_47_real;
      end
      6'b110000 : begin
        _zz_4510_ = int_reg_array_38_48_imag;
        _zz_4511_ = int_reg_array_38_48_real;
      end
      6'b110001 : begin
        _zz_4510_ = int_reg_array_38_49_imag;
        _zz_4511_ = int_reg_array_38_49_real;
      end
      6'b110010 : begin
        _zz_4510_ = int_reg_array_38_50_imag;
        _zz_4511_ = int_reg_array_38_50_real;
      end
      6'b110011 : begin
        _zz_4510_ = int_reg_array_38_51_imag;
        _zz_4511_ = int_reg_array_38_51_real;
      end
      6'b110100 : begin
        _zz_4510_ = int_reg_array_38_52_imag;
        _zz_4511_ = int_reg_array_38_52_real;
      end
      6'b110101 : begin
        _zz_4510_ = int_reg_array_38_53_imag;
        _zz_4511_ = int_reg_array_38_53_real;
      end
      6'b110110 : begin
        _zz_4510_ = int_reg_array_38_54_imag;
        _zz_4511_ = int_reg_array_38_54_real;
      end
      6'b110111 : begin
        _zz_4510_ = int_reg_array_38_55_imag;
        _zz_4511_ = int_reg_array_38_55_real;
      end
      6'b111000 : begin
        _zz_4510_ = int_reg_array_38_56_imag;
        _zz_4511_ = int_reg_array_38_56_real;
      end
      6'b111001 : begin
        _zz_4510_ = int_reg_array_38_57_imag;
        _zz_4511_ = int_reg_array_38_57_real;
      end
      6'b111010 : begin
        _zz_4510_ = int_reg_array_38_58_imag;
        _zz_4511_ = int_reg_array_38_58_real;
      end
      6'b111011 : begin
        _zz_4510_ = int_reg_array_38_59_imag;
        _zz_4511_ = int_reg_array_38_59_real;
      end
      6'b111100 : begin
        _zz_4510_ = int_reg_array_38_60_imag;
        _zz_4511_ = int_reg_array_38_60_real;
      end
      6'b111101 : begin
        _zz_4510_ = int_reg_array_38_61_imag;
        _zz_4511_ = int_reg_array_38_61_real;
      end
      6'b111110 : begin
        _zz_4510_ = int_reg_array_38_62_imag;
        _zz_4511_ = int_reg_array_38_62_real;
      end
      default : begin
        _zz_4510_ = int_reg_array_38_63_imag;
        _zz_4511_ = int_reg_array_38_63_real;
      end
    endcase
  end

  always @(*) begin
    case(_zz_2708_)
      6'b000000 : begin
        _zz_4512_ = int_reg_array_39_0_imag;
        _zz_4513_ = int_reg_array_39_0_real;
      end
      6'b000001 : begin
        _zz_4512_ = int_reg_array_39_1_imag;
        _zz_4513_ = int_reg_array_39_1_real;
      end
      6'b000010 : begin
        _zz_4512_ = int_reg_array_39_2_imag;
        _zz_4513_ = int_reg_array_39_2_real;
      end
      6'b000011 : begin
        _zz_4512_ = int_reg_array_39_3_imag;
        _zz_4513_ = int_reg_array_39_3_real;
      end
      6'b000100 : begin
        _zz_4512_ = int_reg_array_39_4_imag;
        _zz_4513_ = int_reg_array_39_4_real;
      end
      6'b000101 : begin
        _zz_4512_ = int_reg_array_39_5_imag;
        _zz_4513_ = int_reg_array_39_5_real;
      end
      6'b000110 : begin
        _zz_4512_ = int_reg_array_39_6_imag;
        _zz_4513_ = int_reg_array_39_6_real;
      end
      6'b000111 : begin
        _zz_4512_ = int_reg_array_39_7_imag;
        _zz_4513_ = int_reg_array_39_7_real;
      end
      6'b001000 : begin
        _zz_4512_ = int_reg_array_39_8_imag;
        _zz_4513_ = int_reg_array_39_8_real;
      end
      6'b001001 : begin
        _zz_4512_ = int_reg_array_39_9_imag;
        _zz_4513_ = int_reg_array_39_9_real;
      end
      6'b001010 : begin
        _zz_4512_ = int_reg_array_39_10_imag;
        _zz_4513_ = int_reg_array_39_10_real;
      end
      6'b001011 : begin
        _zz_4512_ = int_reg_array_39_11_imag;
        _zz_4513_ = int_reg_array_39_11_real;
      end
      6'b001100 : begin
        _zz_4512_ = int_reg_array_39_12_imag;
        _zz_4513_ = int_reg_array_39_12_real;
      end
      6'b001101 : begin
        _zz_4512_ = int_reg_array_39_13_imag;
        _zz_4513_ = int_reg_array_39_13_real;
      end
      6'b001110 : begin
        _zz_4512_ = int_reg_array_39_14_imag;
        _zz_4513_ = int_reg_array_39_14_real;
      end
      6'b001111 : begin
        _zz_4512_ = int_reg_array_39_15_imag;
        _zz_4513_ = int_reg_array_39_15_real;
      end
      6'b010000 : begin
        _zz_4512_ = int_reg_array_39_16_imag;
        _zz_4513_ = int_reg_array_39_16_real;
      end
      6'b010001 : begin
        _zz_4512_ = int_reg_array_39_17_imag;
        _zz_4513_ = int_reg_array_39_17_real;
      end
      6'b010010 : begin
        _zz_4512_ = int_reg_array_39_18_imag;
        _zz_4513_ = int_reg_array_39_18_real;
      end
      6'b010011 : begin
        _zz_4512_ = int_reg_array_39_19_imag;
        _zz_4513_ = int_reg_array_39_19_real;
      end
      6'b010100 : begin
        _zz_4512_ = int_reg_array_39_20_imag;
        _zz_4513_ = int_reg_array_39_20_real;
      end
      6'b010101 : begin
        _zz_4512_ = int_reg_array_39_21_imag;
        _zz_4513_ = int_reg_array_39_21_real;
      end
      6'b010110 : begin
        _zz_4512_ = int_reg_array_39_22_imag;
        _zz_4513_ = int_reg_array_39_22_real;
      end
      6'b010111 : begin
        _zz_4512_ = int_reg_array_39_23_imag;
        _zz_4513_ = int_reg_array_39_23_real;
      end
      6'b011000 : begin
        _zz_4512_ = int_reg_array_39_24_imag;
        _zz_4513_ = int_reg_array_39_24_real;
      end
      6'b011001 : begin
        _zz_4512_ = int_reg_array_39_25_imag;
        _zz_4513_ = int_reg_array_39_25_real;
      end
      6'b011010 : begin
        _zz_4512_ = int_reg_array_39_26_imag;
        _zz_4513_ = int_reg_array_39_26_real;
      end
      6'b011011 : begin
        _zz_4512_ = int_reg_array_39_27_imag;
        _zz_4513_ = int_reg_array_39_27_real;
      end
      6'b011100 : begin
        _zz_4512_ = int_reg_array_39_28_imag;
        _zz_4513_ = int_reg_array_39_28_real;
      end
      6'b011101 : begin
        _zz_4512_ = int_reg_array_39_29_imag;
        _zz_4513_ = int_reg_array_39_29_real;
      end
      6'b011110 : begin
        _zz_4512_ = int_reg_array_39_30_imag;
        _zz_4513_ = int_reg_array_39_30_real;
      end
      6'b011111 : begin
        _zz_4512_ = int_reg_array_39_31_imag;
        _zz_4513_ = int_reg_array_39_31_real;
      end
      6'b100000 : begin
        _zz_4512_ = int_reg_array_39_32_imag;
        _zz_4513_ = int_reg_array_39_32_real;
      end
      6'b100001 : begin
        _zz_4512_ = int_reg_array_39_33_imag;
        _zz_4513_ = int_reg_array_39_33_real;
      end
      6'b100010 : begin
        _zz_4512_ = int_reg_array_39_34_imag;
        _zz_4513_ = int_reg_array_39_34_real;
      end
      6'b100011 : begin
        _zz_4512_ = int_reg_array_39_35_imag;
        _zz_4513_ = int_reg_array_39_35_real;
      end
      6'b100100 : begin
        _zz_4512_ = int_reg_array_39_36_imag;
        _zz_4513_ = int_reg_array_39_36_real;
      end
      6'b100101 : begin
        _zz_4512_ = int_reg_array_39_37_imag;
        _zz_4513_ = int_reg_array_39_37_real;
      end
      6'b100110 : begin
        _zz_4512_ = int_reg_array_39_38_imag;
        _zz_4513_ = int_reg_array_39_38_real;
      end
      6'b100111 : begin
        _zz_4512_ = int_reg_array_39_39_imag;
        _zz_4513_ = int_reg_array_39_39_real;
      end
      6'b101000 : begin
        _zz_4512_ = int_reg_array_39_40_imag;
        _zz_4513_ = int_reg_array_39_40_real;
      end
      6'b101001 : begin
        _zz_4512_ = int_reg_array_39_41_imag;
        _zz_4513_ = int_reg_array_39_41_real;
      end
      6'b101010 : begin
        _zz_4512_ = int_reg_array_39_42_imag;
        _zz_4513_ = int_reg_array_39_42_real;
      end
      6'b101011 : begin
        _zz_4512_ = int_reg_array_39_43_imag;
        _zz_4513_ = int_reg_array_39_43_real;
      end
      6'b101100 : begin
        _zz_4512_ = int_reg_array_39_44_imag;
        _zz_4513_ = int_reg_array_39_44_real;
      end
      6'b101101 : begin
        _zz_4512_ = int_reg_array_39_45_imag;
        _zz_4513_ = int_reg_array_39_45_real;
      end
      6'b101110 : begin
        _zz_4512_ = int_reg_array_39_46_imag;
        _zz_4513_ = int_reg_array_39_46_real;
      end
      6'b101111 : begin
        _zz_4512_ = int_reg_array_39_47_imag;
        _zz_4513_ = int_reg_array_39_47_real;
      end
      6'b110000 : begin
        _zz_4512_ = int_reg_array_39_48_imag;
        _zz_4513_ = int_reg_array_39_48_real;
      end
      6'b110001 : begin
        _zz_4512_ = int_reg_array_39_49_imag;
        _zz_4513_ = int_reg_array_39_49_real;
      end
      6'b110010 : begin
        _zz_4512_ = int_reg_array_39_50_imag;
        _zz_4513_ = int_reg_array_39_50_real;
      end
      6'b110011 : begin
        _zz_4512_ = int_reg_array_39_51_imag;
        _zz_4513_ = int_reg_array_39_51_real;
      end
      6'b110100 : begin
        _zz_4512_ = int_reg_array_39_52_imag;
        _zz_4513_ = int_reg_array_39_52_real;
      end
      6'b110101 : begin
        _zz_4512_ = int_reg_array_39_53_imag;
        _zz_4513_ = int_reg_array_39_53_real;
      end
      6'b110110 : begin
        _zz_4512_ = int_reg_array_39_54_imag;
        _zz_4513_ = int_reg_array_39_54_real;
      end
      6'b110111 : begin
        _zz_4512_ = int_reg_array_39_55_imag;
        _zz_4513_ = int_reg_array_39_55_real;
      end
      6'b111000 : begin
        _zz_4512_ = int_reg_array_39_56_imag;
        _zz_4513_ = int_reg_array_39_56_real;
      end
      6'b111001 : begin
        _zz_4512_ = int_reg_array_39_57_imag;
        _zz_4513_ = int_reg_array_39_57_real;
      end
      6'b111010 : begin
        _zz_4512_ = int_reg_array_39_58_imag;
        _zz_4513_ = int_reg_array_39_58_real;
      end
      6'b111011 : begin
        _zz_4512_ = int_reg_array_39_59_imag;
        _zz_4513_ = int_reg_array_39_59_real;
      end
      6'b111100 : begin
        _zz_4512_ = int_reg_array_39_60_imag;
        _zz_4513_ = int_reg_array_39_60_real;
      end
      6'b111101 : begin
        _zz_4512_ = int_reg_array_39_61_imag;
        _zz_4513_ = int_reg_array_39_61_real;
      end
      6'b111110 : begin
        _zz_4512_ = int_reg_array_39_62_imag;
        _zz_4513_ = int_reg_array_39_62_real;
      end
      default : begin
        _zz_4512_ = int_reg_array_39_63_imag;
        _zz_4513_ = int_reg_array_39_63_real;
      end
    endcase
  end

  always @(*) begin
    case(_zz_2777_)
      6'b000000 : begin
        _zz_4514_ = int_reg_array_40_0_imag;
        _zz_4515_ = int_reg_array_40_0_real;
      end
      6'b000001 : begin
        _zz_4514_ = int_reg_array_40_1_imag;
        _zz_4515_ = int_reg_array_40_1_real;
      end
      6'b000010 : begin
        _zz_4514_ = int_reg_array_40_2_imag;
        _zz_4515_ = int_reg_array_40_2_real;
      end
      6'b000011 : begin
        _zz_4514_ = int_reg_array_40_3_imag;
        _zz_4515_ = int_reg_array_40_3_real;
      end
      6'b000100 : begin
        _zz_4514_ = int_reg_array_40_4_imag;
        _zz_4515_ = int_reg_array_40_4_real;
      end
      6'b000101 : begin
        _zz_4514_ = int_reg_array_40_5_imag;
        _zz_4515_ = int_reg_array_40_5_real;
      end
      6'b000110 : begin
        _zz_4514_ = int_reg_array_40_6_imag;
        _zz_4515_ = int_reg_array_40_6_real;
      end
      6'b000111 : begin
        _zz_4514_ = int_reg_array_40_7_imag;
        _zz_4515_ = int_reg_array_40_7_real;
      end
      6'b001000 : begin
        _zz_4514_ = int_reg_array_40_8_imag;
        _zz_4515_ = int_reg_array_40_8_real;
      end
      6'b001001 : begin
        _zz_4514_ = int_reg_array_40_9_imag;
        _zz_4515_ = int_reg_array_40_9_real;
      end
      6'b001010 : begin
        _zz_4514_ = int_reg_array_40_10_imag;
        _zz_4515_ = int_reg_array_40_10_real;
      end
      6'b001011 : begin
        _zz_4514_ = int_reg_array_40_11_imag;
        _zz_4515_ = int_reg_array_40_11_real;
      end
      6'b001100 : begin
        _zz_4514_ = int_reg_array_40_12_imag;
        _zz_4515_ = int_reg_array_40_12_real;
      end
      6'b001101 : begin
        _zz_4514_ = int_reg_array_40_13_imag;
        _zz_4515_ = int_reg_array_40_13_real;
      end
      6'b001110 : begin
        _zz_4514_ = int_reg_array_40_14_imag;
        _zz_4515_ = int_reg_array_40_14_real;
      end
      6'b001111 : begin
        _zz_4514_ = int_reg_array_40_15_imag;
        _zz_4515_ = int_reg_array_40_15_real;
      end
      6'b010000 : begin
        _zz_4514_ = int_reg_array_40_16_imag;
        _zz_4515_ = int_reg_array_40_16_real;
      end
      6'b010001 : begin
        _zz_4514_ = int_reg_array_40_17_imag;
        _zz_4515_ = int_reg_array_40_17_real;
      end
      6'b010010 : begin
        _zz_4514_ = int_reg_array_40_18_imag;
        _zz_4515_ = int_reg_array_40_18_real;
      end
      6'b010011 : begin
        _zz_4514_ = int_reg_array_40_19_imag;
        _zz_4515_ = int_reg_array_40_19_real;
      end
      6'b010100 : begin
        _zz_4514_ = int_reg_array_40_20_imag;
        _zz_4515_ = int_reg_array_40_20_real;
      end
      6'b010101 : begin
        _zz_4514_ = int_reg_array_40_21_imag;
        _zz_4515_ = int_reg_array_40_21_real;
      end
      6'b010110 : begin
        _zz_4514_ = int_reg_array_40_22_imag;
        _zz_4515_ = int_reg_array_40_22_real;
      end
      6'b010111 : begin
        _zz_4514_ = int_reg_array_40_23_imag;
        _zz_4515_ = int_reg_array_40_23_real;
      end
      6'b011000 : begin
        _zz_4514_ = int_reg_array_40_24_imag;
        _zz_4515_ = int_reg_array_40_24_real;
      end
      6'b011001 : begin
        _zz_4514_ = int_reg_array_40_25_imag;
        _zz_4515_ = int_reg_array_40_25_real;
      end
      6'b011010 : begin
        _zz_4514_ = int_reg_array_40_26_imag;
        _zz_4515_ = int_reg_array_40_26_real;
      end
      6'b011011 : begin
        _zz_4514_ = int_reg_array_40_27_imag;
        _zz_4515_ = int_reg_array_40_27_real;
      end
      6'b011100 : begin
        _zz_4514_ = int_reg_array_40_28_imag;
        _zz_4515_ = int_reg_array_40_28_real;
      end
      6'b011101 : begin
        _zz_4514_ = int_reg_array_40_29_imag;
        _zz_4515_ = int_reg_array_40_29_real;
      end
      6'b011110 : begin
        _zz_4514_ = int_reg_array_40_30_imag;
        _zz_4515_ = int_reg_array_40_30_real;
      end
      6'b011111 : begin
        _zz_4514_ = int_reg_array_40_31_imag;
        _zz_4515_ = int_reg_array_40_31_real;
      end
      6'b100000 : begin
        _zz_4514_ = int_reg_array_40_32_imag;
        _zz_4515_ = int_reg_array_40_32_real;
      end
      6'b100001 : begin
        _zz_4514_ = int_reg_array_40_33_imag;
        _zz_4515_ = int_reg_array_40_33_real;
      end
      6'b100010 : begin
        _zz_4514_ = int_reg_array_40_34_imag;
        _zz_4515_ = int_reg_array_40_34_real;
      end
      6'b100011 : begin
        _zz_4514_ = int_reg_array_40_35_imag;
        _zz_4515_ = int_reg_array_40_35_real;
      end
      6'b100100 : begin
        _zz_4514_ = int_reg_array_40_36_imag;
        _zz_4515_ = int_reg_array_40_36_real;
      end
      6'b100101 : begin
        _zz_4514_ = int_reg_array_40_37_imag;
        _zz_4515_ = int_reg_array_40_37_real;
      end
      6'b100110 : begin
        _zz_4514_ = int_reg_array_40_38_imag;
        _zz_4515_ = int_reg_array_40_38_real;
      end
      6'b100111 : begin
        _zz_4514_ = int_reg_array_40_39_imag;
        _zz_4515_ = int_reg_array_40_39_real;
      end
      6'b101000 : begin
        _zz_4514_ = int_reg_array_40_40_imag;
        _zz_4515_ = int_reg_array_40_40_real;
      end
      6'b101001 : begin
        _zz_4514_ = int_reg_array_40_41_imag;
        _zz_4515_ = int_reg_array_40_41_real;
      end
      6'b101010 : begin
        _zz_4514_ = int_reg_array_40_42_imag;
        _zz_4515_ = int_reg_array_40_42_real;
      end
      6'b101011 : begin
        _zz_4514_ = int_reg_array_40_43_imag;
        _zz_4515_ = int_reg_array_40_43_real;
      end
      6'b101100 : begin
        _zz_4514_ = int_reg_array_40_44_imag;
        _zz_4515_ = int_reg_array_40_44_real;
      end
      6'b101101 : begin
        _zz_4514_ = int_reg_array_40_45_imag;
        _zz_4515_ = int_reg_array_40_45_real;
      end
      6'b101110 : begin
        _zz_4514_ = int_reg_array_40_46_imag;
        _zz_4515_ = int_reg_array_40_46_real;
      end
      6'b101111 : begin
        _zz_4514_ = int_reg_array_40_47_imag;
        _zz_4515_ = int_reg_array_40_47_real;
      end
      6'b110000 : begin
        _zz_4514_ = int_reg_array_40_48_imag;
        _zz_4515_ = int_reg_array_40_48_real;
      end
      6'b110001 : begin
        _zz_4514_ = int_reg_array_40_49_imag;
        _zz_4515_ = int_reg_array_40_49_real;
      end
      6'b110010 : begin
        _zz_4514_ = int_reg_array_40_50_imag;
        _zz_4515_ = int_reg_array_40_50_real;
      end
      6'b110011 : begin
        _zz_4514_ = int_reg_array_40_51_imag;
        _zz_4515_ = int_reg_array_40_51_real;
      end
      6'b110100 : begin
        _zz_4514_ = int_reg_array_40_52_imag;
        _zz_4515_ = int_reg_array_40_52_real;
      end
      6'b110101 : begin
        _zz_4514_ = int_reg_array_40_53_imag;
        _zz_4515_ = int_reg_array_40_53_real;
      end
      6'b110110 : begin
        _zz_4514_ = int_reg_array_40_54_imag;
        _zz_4515_ = int_reg_array_40_54_real;
      end
      6'b110111 : begin
        _zz_4514_ = int_reg_array_40_55_imag;
        _zz_4515_ = int_reg_array_40_55_real;
      end
      6'b111000 : begin
        _zz_4514_ = int_reg_array_40_56_imag;
        _zz_4515_ = int_reg_array_40_56_real;
      end
      6'b111001 : begin
        _zz_4514_ = int_reg_array_40_57_imag;
        _zz_4515_ = int_reg_array_40_57_real;
      end
      6'b111010 : begin
        _zz_4514_ = int_reg_array_40_58_imag;
        _zz_4515_ = int_reg_array_40_58_real;
      end
      6'b111011 : begin
        _zz_4514_ = int_reg_array_40_59_imag;
        _zz_4515_ = int_reg_array_40_59_real;
      end
      6'b111100 : begin
        _zz_4514_ = int_reg_array_40_60_imag;
        _zz_4515_ = int_reg_array_40_60_real;
      end
      6'b111101 : begin
        _zz_4514_ = int_reg_array_40_61_imag;
        _zz_4515_ = int_reg_array_40_61_real;
      end
      6'b111110 : begin
        _zz_4514_ = int_reg_array_40_62_imag;
        _zz_4515_ = int_reg_array_40_62_real;
      end
      default : begin
        _zz_4514_ = int_reg_array_40_63_imag;
        _zz_4515_ = int_reg_array_40_63_real;
      end
    endcase
  end

  always @(*) begin
    case(_zz_2846_)
      6'b000000 : begin
        _zz_4516_ = int_reg_array_41_0_imag;
        _zz_4517_ = int_reg_array_41_0_real;
      end
      6'b000001 : begin
        _zz_4516_ = int_reg_array_41_1_imag;
        _zz_4517_ = int_reg_array_41_1_real;
      end
      6'b000010 : begin
        _zz_4516_ = int_reg_array_41_2_imag;
        _zz_4517_ = int_reg_array_41_2_real;
      end
      6'b000011 : begin
        _zz_4516_ = int_reg_array_41_3_imag;
        _zz_4517_ = int_reg_array_41_3_real;
      end
      6'b000100 : begin
        _zz_4516_ = int_reg_array_41_4_imag;
        _zz_4517_ = int_reg_array_41_4_real;
      end
      6'b000101 : begin
        _zz_4516_ = int_reg_array_41_5_imag;
        _zz_4517_ = int_reg_array_41_5_real;
      end
      6'b000110 : begin
        _zz_4516_ = int_reg_array_41_6_imag;
        _zz_4517_ = int_reg_array_41_6_real;
      end
      6'b000111 : begin
        _zz_4516_ = int_reg_array_41_7_imag;
        _zz_4517_ = int_reg_array_41_7_real;
      end
      6'b001000 : begin
        _zz_4516_ = int_reg_array_41_8_imag;
        _zz_4517_ = int_reg_array_41_8_real;
      end
      6'b001001 : begin
        _zz_4516_ = int_reg_array_41_9_imag;
        _zz_4517_ = int_reg_array_41_9_real;
      end
      6'b001010 : begin
        _zz_4516_ = int_reg_array_41_10_imag;
        _zz_4517_ = int_reg_array_41_10_real;
      end
      6'b001011 : begin
        _zz_4516_ = int_reg_array_41_11_imag;
        _zz_4517_ = int_reg_array_41_11_real;
      end
      6'b001100 : begin
        _zz_4516_ = int_reg_array_41_12_imag;
        _zz_4517_ = int_reg_array_41_12_real;
      end
      6'b001101 : begin
        _zz_4516_ = int_reg_array_41_13_imag;
        _zz_4517_ = int_reg_array_41_13_real;
      end
      6'b001110 : begin
        _zz_4516_ = int_reg_array_41_14_imag;
        _zz_4517_ = int_reg_array_41_14_real;
      end
      6'b001111 : begin
        _zz_4516_ = int_reg_array_41_15_imag;
        _zz_4517_ = int_reg_array_41_15_real;
      end
      6'b010000 : begin
        _zz_4516_ = int_reg_array_41_16_imag;
        _zz_4517_ = int_reg_array_41_16_real;
      end
      6'b010001 : begin
        _zz_4516_ = int_reg_array_41_17_imag;
        _zz_4517_ = int_reg_array_41_17_real;
      end
      6'b010010 : begin
        _zz_4516_ = int_reg_array_41_18_imag;
        _zz_4517_ = int_reg_array_41_18_real;
      end
      6'b010011 : begin
        _zz_4516_ = int_reg_array_41_19_imag;
        _zz_4517_ = int_reg_array_41_19_real;
      end
      6'b010100 : begin
        _zz_4516_ = int_reg_array_41_20_imag;
        _zz_4517_ = int_reg_array_41_20_real;
      end
      6'b010101 : begin
        _zz_4516_ = int_reg_array_41_21_imag;
        _zz_4517_ = int_reg_array_41_21_real;
      end
      6'b010110 : begin
        _zz_4516_ = int_reg_array_41_22_imag;
        _zz_4517_ = int_reg_array_41_22_real;
      end
      6'b010111 : begin
        _zz_4516_ = int_reg_array_41_23_imag;
        _zz_4517_ = int_reg_array_41_23_real;
      end
      6'b011000 : begin
        _zz_4516_ = int_reg_array_41_24_imag;
        _zz_4517_ = int_reg_array_41_24_real;
      end
      6'b011001 : begin
        _zz_4516_ = int_reg_array_41_25_imag;
        _zz_4517_ = int_reg_array_41_25_real;
      end
      6'b011010 : begin
        _zz_4516_ = int_reg_array_41_26_imag;
        _zz_4517_ = int_reg_array_41_26_real;
      end
      6'b011011 : begin
        _zz_4516_ = int_reg_array_41_27_imag;
        _zz_4517_ = int_reg_array_41_27_real;
      end
      6'b011100 : begin
        _zz_4516_ = int_reg_array_41_28_imag;
        _zz_4517_ = int_reg_array_41_28_real;
      end
      6'b011101 : begin
        _zz_4516_ = int_reg_array_41_29_imag;
        _zz_4517_ = int_reg_array_41_29_real;
      end
      6'b011110 : begin
        _zz_4516_ = int_reg_array_41_30_imag;
        _zz_4517_ = int_reg_array_41_30_real;
      end
      6'b011111 : begin
        _zz_4516_ = int_reg_array_41_31_imag;
        _zz_4517_ = int_reg_array_41_31_real;
      end
      6'b100000 : begin
        _zz_4516_ = int_reg_array_41_32_imag;
        _zz_4517_ = int_reg_array_41_32_real;
      end
      6'b100001 : begin
        _zz_4516_ = int_reg_array_41_33_imag;
        _zz_4517_ = int_reg_array_41_33_real;
      end
      6'b100010 : begin
        _zz_4516_ = int_reg_array_41_34_imag;
        _zz_4517_ = int_reg_array_41_34_real;
      end
      6'b100011 : begin
        _zz_4516_ = int_reg_array_41_35_imag;
        _zz_4517_ = int_reg_array_41_35_real;
      end
      6'b100100 : begin
        _zz_4516_ = int_reg_array_41_36_imag;
        _zz_4517_ = int_reg_array_41_36_real;
      end
      6'b100101 : begin
        _zz_4516_ = int_reg_array_41_37_imag;
        _zz_4517_ = int_reg_array_41_37_real;
      end
      6'b100110 : begin
        _zz_4516_ = int_reg_array_41_38_imag;
        _zz_4517_ = int_reg_array_41_38_real;
      end
      6'b100111 : begin
        _zz_4516_ = int_reg_array_41_39_imag;
        _zz_4517_ = int_reg_array_41_39_real;
      end
      6'b101000 : begin
        _zz_4516_ = int_reg_array_41_40_imag;
        _zz_4517_ = int_reg_array_41_40_real;
      end
      6'b101001 : begin
        _zz_4516_ = int_reg_array_41_41_imag;
        _zz_4517_ = int_reg_array_41_41_real;
      end
      6'b101010 : begin
        _zz_4516_ = int_reg_array_41_42_imag;
        _zz_4517_ = int_reg_array_41_42_real;
      end
      6'b101011 : begin
        _zz_4516_ = int_reg_array_41_43_imag;
        _zz_4517_ = int_reg_array_41_43_real;
      end
      6'b101100 : begin
        _zz_4516_ = int_reg_array_41_44_imag;
        _zz_4517_ = int_reg_array_41_44_real;
      end
      6'b101101 : begin
        _zz_4516_ = int_reg_array_41_45_imag;
        _zz_4517_ = int_reg_array_41_45_real;
      end
      6'b101110 : begin
        _zz_4516_ = int_reg_array_41_46_imag;
        _zz_4517_ = int_reg_array_41_46_real;
      end
      6'b101111 : begin
        _zz_4516_ = int_reg_array_41_47_imag;
        _zz_4517_ = int_reg_array_41_47_real;
      end
      6'b110000 : begin
        _zz_4516_ = int_reg_array_41_48_imag;
        _zz_4517_ = int_reg_array_41_48_real;
      end
      6'b110001 : begin
        _zz_4516_ = int_reg_array_41_49_imag;
        _zz_4517_ = int_reg_array_41_49_real;
      end
      6'b110010 : begin
        _zz_4516_ = int_reg_array_41_50_imag;
        _zz_4517_ = int_reg_array_41_50_real;
      end
      6'b110011 : begin
        _zz_4516_ = int_reg_array_41_51_imag;
        _zz_4517_ = int_reg_array_41_51_real;
      end
      6'b110100 : begin
        _zz_4516_ = int_reg_array_41_52_imag;
        _zz_4517_ = int_reg_array_41_52_real;
      end
      6'b110101 : begin
        _zz_4516_ = int_reg_array_41_53_imag;
        _zz_4517_ = int_reg_array_41_53_real;
      end
      6'b110110 : begin
        _zz_4516_ = int_reg_array_41_54_imag;
        _zz_4517_ = int_reg_array_41_54_real;
      end
      6'b110111 : begin
        _zz_4516_ = int_reg_array_41_55_imag;
        _zz_4517_ = int_reg_array_41_55_real;
      end
      6'b111000 : begin
        _zz_4516_ = int_reg_array_41_56_imag;
        _zz_4517_ = int_reg_array_41_56_real;
      end
      6'b111001 : begin
        _zz_4516_ = int_reg_array_41_57_imag;
        _zz_4517_ = int_reg_array_41_57_real;
      end
      6'b111010 : begin
        _zz_4516_ = int_reg_array_41_58_imag;
        _zz_4517_ = int_reg_array_41_58_real;
      end
      6'b111011 : begin
        _zz_4516_ = int_reg_array_41_59_imag;
        _zz_4517_ = int_reg_array_41_59_real;
      end
      6'b111100 : begin
        _zz_4516_ = int_reg_array_41_60_imag;
        _zz_4517_ = int_reg_array_41_60_real;
      end
      6'b111101 : begin
        _zz_4516_ = int_reg_array_41_61_imag;
        _zz_4517_ = int_reg_array_41_61_real;
      end
      6'b111110 : begin
        _zz_4516_ = int_reg_array_41_62_imag;
        _zz_4517_ = int_reg_array_41_62_real;
      end
      default : begin
        _zz_4516_ = int_reg_array_41_63_imag;
        _zz_4517_ = int_reg_array_41_63_real;
      end
    endcase
  end

  always @(*) begin
    case(_zz_2915_)
      6'b000000 : begin
        _zz_4518_ = int_reg_array_42_0_imag;
        _zz_4519_ = int_reg_array_42_0_real;
      end
      6'b000001 : begin
        _zz_4518_ = int_reg_array_42_1_imag;
        _zz_4519_ = int_reg_array_42_1_real;
      end
      6'b000010 : begin
        _zz_4518_ = int_reg_array_42_2_imag;
        _zz_4519_ = int_reg_array_42_2_real;
      end
      6'b000011 : begin
        _zz_4518_ = int_reg_array_42_3_imag;
        _zz_4519_ = int_reg_array_42_3_real;
      end
      6'b000100 : begin
        _zz_4518_ = int_reg_array_42_4_imag;
        _zz_4519_ = int_reg_array_42_4_real;
      end
      6'b000101 : begin
        _zz_4518_ = int_reg_array_42_5_imag;
        _zz_4519_ = int_reg_array_42_5_real;
      end
      6'b000110 : begin
        _zz_4518_ = int_reg_array_42_6_imag;
        _zz_4519_ = int_reg_array_42_6_real;
      end
      6'b000111 : begin
        _zz_4518_ = int_reg_array_42_7_imag;
        _zz_4519_ = int_reg_array_42_7_real;
      end
      6'b001000 : begin
        _zz_4518_ = int_reg_array_42_8_imag;
        _zz_4519_ = int_reg_array_42_8_real;
      end
      6'b001001 : begin
        _zz_4518_ = int_reg_array_42_9_imag;
        _zz_4519_ = int_reg_array_42_9_real;
      end
      6'b001010 : begin
        _zz_4518_ = int_reg_array_42_10_imag;
        _zz_4519_ = int_reg_array_42_10_real;
      end
      6'b001011 : begin
        _zz_4518_ = int_reg_array_42_11_imag;
        _zz_4519_ = int_reg_array_42_11_real;
      end
      6'b001100 : begin
        _zz_4518_ = int_reg_array_42_12_imag;
        _zz_4519_ = int_reg_array_42_12_real;
      end
      6'b001101 : begin
        _zz_4518_ = int_reg_array_42_13_imag;
        _zz_4519_ = int_reg_array_42_13_real;
      end
      6'b001110 : begin
        _zz_4518_ = int_reg_array_42_14_imag;
        _zz_4519_ = int_reg_array_42_14_real;
      end
      6'b001111 : begin
        _zz_4518_ = int_reg_array_42_15_imag;
        _zz_4519_ = int_reg_array_42_15_real;
      end
      6'b010000 : begin
        _zz_4518_ = int_reg_array_42_16_imag;
        _zz_4519_ = int_reg_array_42_16_real;
      end
      6'b010001 : begin
        _zz_4518_ = int_reg_array_42_17_imag;
        _zz_4519_ = int_reg_array_42_17_real;
      end
      6'b010010 : begin
        _zz_4518_ = int_reg_array_42_18_imag;
        _zz_4519_ = int_reg_array_42_18_real;
      end
      6'b010011 : begin
        _zz_4518_ = int_reg_array_42_19_imag;
        _zz_4519_ = int_reg_array_42_19_real;
      end
      6'b010100 : begin
        _zz_4518_ = int_reg_array_42_20_imag;
        _zz_4519_ = int_reg_array_42_20_real;
      end
      6'b010101 : begin
        _zz_4518_ = int_reg_array_42_21_imag;
        _zz_4519_ = int_reg_array_42_21_real;
      end
      6'b010110 : begin
        _zz_4518_ = int_reg_array_42_22_imag;
        _zz_4519_ = int_reg_array_42_22_real;
      end
      6'b010111 : begin
        _zz_4518_ = int_reg_array_42_23_imag;
        _zz_4519_ = int_reg_array_42_23_real;
      end
      6'b011000 : begin
        _zz_4518_ = int_reg_array_42_24_imag;
        _zz_4519_ = int_reg_array_42_24_real;
      end
      6'b011001 : begin
        _zz_4518_ = int_reg_array_42_25_imag;
        _zz_4519_ = int_reg_array_42_25_real;
      end
      6'b011010 : begin
        _zz_4518_ = int_reg_array_42_26_imag;
        _zz_4519_ = int_reg_array_42_26_real;
      end
      6'b011011 : begin
        _zz_4518_ = int_reg_array_42_27_imag;
        _zz_4519_ = int_reg_array_42_27_real;
      end
      6'b011100 : begin
        _zz_4518_ = int_reg_array_42_28_imag;
        _zz_4519_ = int_reg_array_42_28_real;
      end
      6'b011101 : begin
        _zz_4518_ = int_reg_array_42_29_imag;
        _zz_4519_ = int_reg_array_42_29_real;
      end
      6'b011110 : begin
        _zz_4518_ = int_reg_array_42_30_imag;
        _zz_4519_ = int_reg_array_42_30_real;
      end
      6'b011111 : begin
        _zz_4518_ = int_reg_array_42_31_imag;
        _zz_4519_ = int_reg_array_42_31_real;
      end
      6'b100000 : begin
        _zz_4518_ = int_reg_array_42_32_imag;
        _zz_4519_ = int_reg_array_42_32_real;
      end
      6'b100001 : begin
        _zz_4518_ = int_reg_array_42_33_imag;
        _zz_4519_ = int_reg_array_42_33_real;
      end
      6'b100010 : begin
        _zz_4518_ = int_reg_array_42_34_imag;
        _zz_4519_ = int_reg_array_42_34_real;
      end
      6'b100011 : begin
        _zz_4518_ = int_reg_array_42_35_imag;
        _zz_4519_ = int_reg_array_42_35_real;
      end
      6'b100100 : begin
        _zz_4518_ = int_reg_array_42_36_imag;
        _zz_4519_ = int_reg_array_42_36_real;
      end
      6'b100101 : begin
        _zz_4518_ = int_reg_array_42_37_imag;
        _zz_4519_ = int_reg_array_42_37_real;
      end
      6'b100110 : begin
        _zz_4518_ = int_reg_array_42_38_imag;
        _zz_4519_ = int_reg_array_42_38_real;
      end
      6'b100111 : begin
        _zz_4518_ = int_reg_array_42_39_imag;
        _zz_4519_ = int_reg_array_42_39_real;
      end
      6'b101000 : begin
        _zz_4518_ = int_reg_array_42_40_imag;
        _zz_4519_ = int_reg_array_42_40_real;
      end
      6'b101001 : begin
        _zz_4518_ = int_reg_array_42_41_imag;
        _zz_4519_ = int_reg_array_42_41_real;
      end
      6'b101010 : begin
        _zz_4518_ = int_reg_array_42_42_imag;
        _zz_4519_ = int_reg_array_42_42_real;
      end
      6'b101011 : begin
        _zz_4518_ = int_reg_array_42_43_imag;
        _zz_4519_ = int_reg_array_42_43_real;
      end
      6'b101100 : begin
        _zz_4518_ = int_reg_array_42_44_imag;
        _zz_4519_ = int_reg_array_42_44_real;
      end
      6'b101101 : begin
        _zz_4518_ = int_reg_array_42_45_imag;
        _zz_4519_ = int_reg_array_42_45_real;
      end
      6'b101110 : begin
        _zz_4518_ = int_reg_array_42_46_imag;
        _zz_4519_ = int_reg_array_42_46_real;
      end
      6'b101111 : begin
        _zz_4518_ = int_reg_array_42_47_imag;
        _zz_4519_ = int_reg_array_42_47_real;
      end
      6'b110000 : begin
        _zz_4518_ = int_reg_array_42_48_imag;
        _zz_4519_ = int_reg_array_42_48_real;
      end
      6'b110001 : begin
        _zz_4518_ = int_reg_array_42_49_imag;
        _zz_4519_ = int_reg_array_42_49_real;
      end
      6'b110010 : begin
        _zz_4518_ = int_reg_array_42_50_imag;
        _zz_4519_ = int_reg_array_42_50_real;
      end
      6'b110011 : begin
        _zz_4518_ = int_reg_array_42_51_imag;
        _zz_4519_ = int_reg_array_42_51_real;
      end
      6'b110100 : begin
        _zz_4518_ = int_reg_array_42_52_imag;
        _zz_4519_ = int_reg_array_42_52_real;
      end
      6'b110101 : begin
        _zz_4518_ = int_reg_array_42_53_imag;
        _zz_4519_ = int_reg_array_42_53_real;
      end
      6'b110110 : begin
        _zz_4518_ = int_reg_array_42_54_imag;
        _zz_4519_ = int_reg_array_42_54_real;
      end
      6'b110111 : begin
        _zz_4518_ = int_reg_array_42_55_imag;
        _zz_4519_ = int_reg_array_42_55_real;
      end
      6'b111000 : begin
        _zz_4518_ = int_reg_array_42_56_imag;
        _zz_4519_ = int_reg_array_42_56_real;
      end
      6'b111001 : begin
        _zz_4518_ = int_reg_array_42_57_imag;
        _zz_4519_ = int_reg_array_42_57_real;
      end
      6'b111010 : begin
        _zz_4518_ = int_reg_array_42_58_imag;
        _zz_4519_ = int_reg_array_42_58_real;
      end
      6'b111011 : begin
        _zz_4518_ = int_reg_array_42_59_imag;
        _zz_4519_ = int_reg_array_42_59_real;
      end
      6'b111100 : begin
        _zz_4518_ = int_reg_array_42_60_imag;
        _zz_4519_ = int_reg_array_42_60_real;
      end
      6'b111101 : begin
        _zz_4518_ = int_reg_array_42_61_imag;
        _zz_4519_ = int_reg_array_42_61_real;
      end
      6'b111110 : begin
        _zz_4518_ = int_reg_array_42_62_imag;
        _zz_4519_ = int_reg_array_42_62_real;
      end
      default : begin
        _zz_4518_ = int_reg_array_42_63_imag;
        _zz_4519_ = int_reg_array_42_63_real;
      end
    endcase
  end

  always @(*) begin
    case(_zz_2984_)
      6'b000000 : begin
        _zz_4520_ = int_reg_array_43_0_imag;
        _zz_4521_ = int_reg_array_43_0_real;
      end
      6'b000001 : begin
        _zz_4520_ = int_reg_array_43_1_imag;
        _zz_4521_ = int_reg_array_43_1_real;
      end
      6'b000010 : begin
        _zz_4520_ = int_reg_array_43_2_imag;
        _zz_4521_ = int_reg_array_43_2_real;
      end
      6'b000011 : begin
        _zz_4520_ = int_reg_array_43_3_imag;
        _zz_4521_ = int_reg_array_43_3_real;
      end
      6'b000100 : begin
        _zz_4520_ = int_reg_array_43_4_imag;
        _zz_4521_ = int_reg_array_43_4_real;
      end
      6'b000101 : begin
        _zz_4520_ = int_reg_array_43_5_imag;
        _zz_4521_ = int_reg_array_43_5_real;
      end
      6'b000110 : begin
        _zz_4520_ = int_reg_array_43_6_imag;
        _zz_4521_ = int_reg_array_43_6_real;
      end
      6'b000111 : begin
        _zz_4520_ = int_reg_array_43_7_imag;
        _zz_4521_ = int_reg_array_43_7_real;
      end
      6'b001000 : begin
        _zz_4520_ = int_reg_array_43_8_imag;
        _zz_4521_ = int_reg_array_43_8_real;
      end
      6'b001001 : begin
        _zz_4520_ = int_reg_array_43_9_imag;
        _zz_4521_ = int_reg_array_43_9_real;
      end
      6'b001010 : begin
        _zz_4520_ = int_reg_array_43_10_imag;
        _zz_4521_ = int_reg_array_43_10_real;
      end
      6'b001011 : begin
        _zz_4520_ = int_reg_array_43_11_imag;
        _zz_4521_ = int_reg_array_43_11_real;
      end
      6'b001100 : begin
        _zz_4520_ = int_reg_array_43_12_imag;
        _zz_4521_ = int_reg_array_43_12_real;
      end
      6'b001101 : begin
        _zz_4520_ = int_reg_array_43_13_imag;
        _zz_4521_ = int_reg_array_43_13_real;
      end
      6'b001110 : begin
        _zz_4520_ = int_reg_array_43_14_imag;
        _zz_4521_ = int_reg_array_43_14_real;
      end
      6'b001111 : begin
        _zz_4520_ = int_reg_array_43_15_imag;
        _zz_4521_ = int_reg_array_43_15_real;
      end
      6'b010000 : begin
        _zz_4520_ = int_reg_array_43_16_imag;
        _zz_4521_ = int_reg_array_43_16_real;
      end
      6'b010001 : begin
        _zz_4520_ = int_reg_array_43_17_imag;
        _zz_4521_ = int_reg_array_43_17_real;
      end
      6'b010010 : begin
        _zz_4520_ = int_reg_array_43_18_imag;
        _zz_4521_ = int_reg_array_43_18_real;
      end
      6'b010011 : begin
        _zz_4520_ = int_reg_array_43_19_imag;
        _zz_4521_ = int_reg_array_43_19_real;
      end
      6'b010100 : begin
        _zz_4520_ = int_reg_array_43_20_imag;
        _zz_4521_ = int_reg_array_43_20_real;
      end
      6'b010101 : begin
        _zz_4520_ = int_reg_array_43_21_imag;
        _zz_4521_ = int_reg_array_43_21_real;
      end
      6'b010110 : begin
        _zz_4520_ = int_reg_array_43_22_imag;
        _zz_4521_ = int_reg_array_43_22_real;
      end
      6'b010111 : begin
        _zz_4520_ = int_reg_array_43_23_imag;
        _zz_4521_ = int_reg_array_43_23_real;
      end
      6'b011000 : begin
        _zz_4520_ = int_reg_array_43_24_imag;
        _zz_4521_ = int_reg_array_43_24_real;
      end
      6'b011001 : begin
        _zz_4520_ = int_reg_array_43_25_imag;
        _zz_4521_ = int_reg_array_43_25_real;
      end
      6'b011010 : begin
        _zz_4520_ = int_reg_array_43_26_imag;
        _zz_4521_ = int_reg_array_43_26_real;
      end
      6'b011011 : begin
        _zz_4520_ = int_reg_array_43_27_imag;
        _zz_4521_ = int_reg_array_43_27_real;
      end
      6'b011100 : begin
        _zz_4520_ = int_reg_array_43_28_imag;
        _zz_4521_ = int_reg_array_43_28_real;
      end
      6'b011101 : begin
        _zz_4520_ = int_reg_array_43_29_imag;
        _zz_4521_ = int_reg_array_43_29_real;
      end
      6'b011110 : begin
        _zz_4520_ = int_reg_array_43_30_imag;
        _zz_4521_ = int_reg_array_43_30_real;
      end
      6'b011111 : begin
        _zz_4520_ = int_reg_array_43_31_imag;
        _zz_4521_ = int_reg_array_43_31_real;
      end
      6'b100000 : begin
        _zz_4520_ = int_reg_array_43_32_imag;
        _zz_4521_ = int_reg_array_43_32_real;
      end
      6'b100001 : begin
        _zz_4520_ = int_reg_array_43_33_imag;
        _zz_4521_ = int_reg_array_43_33_real;
      end
      6'b100010 : begin
        _zz_4520_ = int_reg_array_43_34_imag;
        _zz_4521_ = int_reg_array_43_34_real;
      end
      6'b100011 : begin
        _zz_4520_ = int_reg_array_43_35_imag;
        _zz_4521_ = int_reg_array_43_35_real;
      end
      6'b100100 : begin
        _zz_4520_ = int_reg_array_43_36_imag;
        _zz_4521_ = int_reg_array_43_36_real;
      end
      6'b100101 : begin
        _zz_4520_ = int_reg_array_43_37_imag;
        _zz_4521_ = int_reg_array_43_37_real;
      end
      6'b100110 : begin
        _zz_4520_ = int_reg_array_43_38_imag;
        _zz_4521_ = int_reg_array_43_38_real;
      end
      6'b100111 : begin
        _zz_4520_ = int_reg_array_43_39_imag;
        _zz_4521_ = int_reg_array_43_39_real;
      end
      6'b101000 : begin
        _zz_4520_ = int_reg_array_43_40_imag;
        _zz_4521_ = int_reg_array_43_40_real;
      end
      6'b101001 : begin
        _zz_4520_ = int_reg_array_43_41_imag;
        _zz_4521_ = int_reg_array_43_41_real;
      end
      6'b101010 : begin
        _zz_4520_ = int_reg_array_43_42_imag;
        _zz_4521_ = int_reg_array_43_42_real;
      end
      6'b101011 : begin
        _zz_4520_ = int_reg_array_43_43_imag;
        _zz_4521_ = int_reg_array_43_43_real;
      end
      6'b101100 : begin
        _zz_4520_ = int_reg_array_43_44_imag;
        _zz_4521_ = int_reg_array_43_44_real;
      end
      6'b101101 : begin
        _zz_4520_ = int_reg_array_43_45_imag;
        _zz_4521_ = int_reg_array_43_45_real;
      end
      6'b101110 : begin
        _zz_4520_ = int_reg_array_43_46_imag;
        _zz_4521_ = int_reg_array_43_46_real;
      end
      6'b101111 : begin
        _zz_4520_ = int_reg_array_43_47_imag;
        _zz_4521_ = int_reg_array_43_47_real;
      end
      6'b110000 : begin
        _zz_4520_ = int_reg_array_43_48_imag;
        _zz_4521_ = int_reg_array_43_48_real;
      end
      6'b110001 : begin
        _zz_4520_ = int_reg_array_43_49_imag;
        _zz_4521_ = int_reg_array_43_49_real;
      end
      6'b110010 : begin
        _zz_4520_ = int_reg_array_43_50_imag;
        _zz_4521_ = int_reg_array_43_50_real;
      end
      6'b110011 : begin
        _zz_4520_ = int_reg_array_43_51_imag;
        _zz_4521_ = int_reg_array_43_51_real;
      end
      6'b110100 : begin
        _zz_4520_ = int_reg_array_43_52_imag;
        _zz_4521_ = int_reg_array_43_52_real;
      end
      6'b110101 : begin
        _zz_4520_ = int_reg_array_43_53_imag;
        _zz_4521_ = int_reg_array_43_53_real;
      end
      6'b110110 : begin
        _zz_4520_ = int_reg_array_43_54_imag;
        _zz_4521_ = int_reg_array_43_54_real;
      end
      6'b110111 : begin
        _zz_4520_ = int_reg_array_43_55_imag;
        _zz_4521_ = int_reg_array_43_55_real;
      end
      6'b111000 : begin
        _zz_4520_ = int_reg_array_43_56_imag;
        _zz_4521_ = int_reg_array_43_56_real;
      end
      6'b111001 : begin
        _zz_4520_ = int_reg_array_43_57_imag;
        _zz_4521_ = int_reg_array_43_57_real;
      end
      6'b111010 : begin
        _zz_4520_ = int_reg_array_43_58_imag;
        _zz_4521_ = int_reg_array_43_58_real;
      end
      6'b111011 : begin
        _zz_4520_ = int_reg_array_43_59_imag;
        _zz_4521_ = int_reg_array_43_59_real;
      end
      6'b111100 : begin
        _zz_4520_ = int_reg_array_43_60_imag;
        _zz_4521_ = int_reg_array_43_60_real;
      end
      6'b111101 : begin
        _zz_4520_ = int_reg_array_43_61_imag;
        _zz_4521_ = int_reg_array_43_61_real;
      end
      6'b111110 : begin
        _zz_4520_ = int_reg_array_43_62_imag;
        _zz_4521_ = int_reg_array_43_62_real;
      end
      default : begin
        _zz_4520_ = int_reg_array_43_63_imag;
        _zz_4521_ = int_reg_array_43_63_real;
      end
    endcase
  end

  always @(*) begin
    case(_zz_3053_)
      6'b000000 : begin
        _zz_4522_ = int_reg_array_44_0_imag;
        _zz_4523_ = int_reg_array_44_0_real;
      end
      6'b000001 : begin
        _zz_4522_ = int_reg_array_44_1_imag;
        _zz_4523_ = int_reg_array_44_1_real;
      end
      6'b000010 : begin
        _zz_4522_ = int_reg_array_44_2_imag;
        _zz_4523_ = int_reg_array_44_2_real;
      end
      6'b000011 : begin
        _zz_4522_ = int_reg_array_44_3_imag;
        _zz_4523_ = int_reg_array_44_3_real;
      end
      6'b000100 : begin
        _zz_4522_ = int_reg_array_44_4_imag;
        _zz_4523_ = int_reg_array_44_4_real;
      end
      6'b000101 : begin
        _zz_4522_ = int_reg_array_44_5_imag;
        _zz_4523_ = int_reg_array_44_5_real;
      end
      6'b000110 : begin
        _zz_4522_ = int_reg_array_44_6_imag;
        _zz_4523_ = int_reg_array_44_6_real;
      end
      6'b000111 : begin
        _zz_4522_ = int_reg_array_44_7_imag;
        _zz_4523_ = int_reg_array_44_7_real;
      end
      6'b001000 : begin
        _zz_4522_ = int_reg_array_44_8_imag;
        _zz_4523_ = int_reg_array_44_8_real;
      end
      6'b001001 : begin
        _zz_4522_ = int_reg_array_44_9_imag;
        _zz_4523_ = int_reg_array_44_9_real;
      end
      6'b001010 : begin
        _zz_4522_ = int_reg_array_44_10_imag;
        _zz_4523_ = int_reg_array_44_10_real;
      end
      6'b001011 : begin
        _zz_4522_ = int_reg_array_44_11_imag;
        _zz_4523_ = int_reg_array_44_11_real;
      end
      6'b001100 : begin
        _zz_4522_ = int_reg_array_44_12_imag;
        _zz_4523_ = int_reg_array_44_12_real;
      end
      6'b001101 : begin
        _zz_4522_ = int_reg_array_44_13_imag;
        _zz_4523_ = int_reg_array_44_13_real;
      end
      6'b001110 : begin
        _zz_4522_ = int_reg_array_44_14_imag;
        _zz_4523_ = int_reg_array_44_14_real;
      end
      6'b001111 : begin
        _zz_4522_ = int_reg_array_44_15_imag;
        _zz_4523_ = int_reg_array_44_15_real;
      end
      6'b010000 : begin
        _zz_4522_ = int_reg_array_44_16_imag;
        _zz_4523_ = int_reg_array_44_16_real;
      end
      6'b010001 : begin
        _zz_4522_ = int_reg_array_44_17_imag;
        _zz_4523_ = int_reg_array_44_17_real;
      end
      6'b010010 : begin
        _zz_4522_ = int_reg_array_44_18_imag;
        _zz_4523_ = int_reg_array_44_18_real;
      end
      6'b010011 : begin
        _zz_4522_ = int_reg_array_44_19_imag;
        _zz_4523_ = int_reg_array_44_19_real;
      end
      6'b010100 : begin
        _zz_4522_ = int_reg_array_44_20_imag;
        _zz_4523_ = int_reg_array_44_20_real;
      end
      6'b010101 : begin
        _zz_4522_ = int_reg_array_44_21_imag;
        _zz_4523_ = int_reg_array_44_21_real;
      end
      6'b010110 : begin
        _zz_4522_ = int_reg_array_44_22_imag;
        _zz_4523_ = int_reg_array_44_22_real;
      end
      6'b010111 : begin
        _zz_4522_ = int_reg_array_44_23_imag;
        _zz_4523_ = int_reg_array_44_23_real;
      end
      6'b011000 : begin
        _zz_4522_ = int_reg_array_44_24_imag;
        _zz_4523_ = int_reg_array_44_24_real;
      end
      6'b011001 : begin
        _zz_4522_ = int_reg_array_44_25_imag;
        _zz_4523_ = int_reg_array_44_25_real;
      end
      6'b011010 : begin
        _zz_4522_ = int_reg_array_44_26_imag;
        _zz_4523_ = int_reg_array_44_26_real;
      end
      6'b011011 : begin
        _zz_4522_ = int_reg_array_44_27_imag;
        _zz_4523_ = int_reg_array_44_27_real;
      end
      6'b011100 : begin
        _zz_4522_ = int_reg_array_44_28_imag;
        _zz_4523_ = int_reg_array_44_28_real;
      end
      6'b011101 : begin
        _zz_4522_ = int_reg_array_44_29_imag;
        _zz_4523_ = int_reg_array_44_29_real;
      end
      6'b011110 : begin
        _zz_4522_ = int_reg_array_44_30_imag;
        _zz_4523_ = int_reg_array_44_30_real;
      end
      6'b011111 : begin
        _zz_4522_ = int_reg_array_44_31_imag;
        _zz_4523_ = int_reg_array_44_31_real;
      end
      6'b100000 : begin
        _zz_4522_ = int_reg_array_44_32_imag;
        _zz_4523_ = int_reg_array_44_32_real;
      end
      6'b100001 : begin
        _zz_4522_ = int_reg_array_44_33_imag;
        _zz_4523_ = int_reg_array_44_33_real;
      end
      6'b100010 : begin
        _zz_4522_ = int_reg_array_44_34_imag;
        _zz_4523_ = int_reg_array_44_34_real;
      end
      6'b100011 : begin
        _zz_4522_ = int_reg_array_44_35_imag;
        _zz_4523_ = int_reg_array_44_35_real;
      end
      6'b100100 : begin
        _zz_4522_ = int_reg_array_44_36_imag;
        _zz_4523_ = int_reg_array_44_36_real;
      end
      6'b100101 : begin
        _zz_4522_ = int_reg_array_44_37_imag;
        _zz_4523_ = int_reg_array_44_37_real;
      end
      6'b100110 : begin
        _zz_4522_ = int_reg_array_44_38_imag;
        _zz_4523_ = int_reg_array_44_38_real;
      end
      6'b100111 : begin
        _zz_4522_ = int_reg_array_44_39_imag;
        _zz_4523_ = int_reg_array_44_39_real;
      end
      6'b101000 : begin
        _zz_4522_ = int_reg_array_44_40_imag;
        _zz_4523_ = int_reg_array_44_40_real;
      end
      6'b101001 : begin
        _zz_4522_ = int_reg_array_44_41_imag;
        _zz_4523_ = int_reg_array_44_41_real;
      end
      6'b101010 : begin
        _zz_4522_ = int_reg_array_44_42_imag;
        _zz_4523_ = int_reg_array_44_42_real;
      end
      6'b101011 : begin
        _zz_4522_ = int_reg_array_44_43_imag;
        _zz_4523_ = int_reg_array_44_43_real;
      end
      6'b101100 : begin
        _zz_4522_ = int_reg_array_44_44_imag;
        _zz_4523_ = int_reg_array_44_44_real;
      end
      6'b101101 : begin
        _zz_4522_ = int_reg_array_44_45_imag;
        _zz_4523_ = int_reg_array_44_45_real;
      end
      6'b101110 : begin
        _zz_4522_ = int_reg_array_44_46_imag;
        _zz_4523_ = int_reg_array_44_46_real;
      end
      6'b101111 : begin
        _zz_4522_ = int_reg_array_44_47_imag;
        _zz_4523_ = int_reg_array_44_47_real;
      end
      6'b110000 : begin
        _zz_4522_ = int_reg_array_44_48_imag;
        _zz_4523_ = int_reg_array_44_48_real;
      end
      6'b110001 : begin
        _zz_4522_ = int_reg_array_44_49_imag;
        _zz_4523_ = int_reg_array_44_49_real;
      end
      6'b110010 : begin
        _zz_4522_ = int_reg_array_44_50_imag;
        _zz_4523_ = int_reg_array_44_50_real;
      end
      6'b110011 : begin
        _zz_4522_ = int_reg_array_44_51_imag;
        _zz_4523_ = int_reg_array_44_51_real;
      end
      6'b110100 : begin
        _zz_4522_ = int_reg_array_44_52_imag;
        _zz_4523_ = int_reg_array_44_52_real;
      end
      6'b110101 : begin
        _zz_4522_ = int_reg_array_44_53_imag;
        _zz_4523_ = int_reg_array_44_53_real;
      end
      6'b110110 : begin
        _zz_4522_ = int_reg_array_44_54_imag;
        _zz_4523_ = int_reg_array_44_54_real;
      end
      6'b110111 : begin
        _zz_4522_ = int_reg_array_44_55_imag;
        _zz_4523_ = int_reg_array_44_55_real;
      end
      6'b111000 : begin
        _zz_4522_ = int_reg_array_44_56_imag;
        _zz_4523_ = int_reg_array_44_56_real;
      end
      6'b111001 : begin
        _zz_4522_ = int_reg_array_44_57_imag;
        _zz_4523_ = int_reg_array_44_57_real;
      end
      6'b111010 : begin
        _zz_4522_ = int_reg_array_44_58_imag;
        _zz_4523_ = int_reg_array_44_58_real;
      end
      6'b111011 : begin
        _zz_4522_ = int_reg_array_44_59_imag;
        _zz_4523_ = int_reg_array_44_59_real;
      end
      6'b111100 : begin
        _zz_4522_ = int_reg_array_44_60_imag;
        _zz_4523_ = int_reg_array_44_60_real;
      end
      6'b111101 : begin
        _zz_4522_ = int_reg_array_44_61_imag;
        _zz_4523_ = int_reg_array_44_61_real;
      end
      6'b111110 : begin
        _zz_4522_ = int_reg_array_44_62_imag;
        _zz_4523_ = int_reg_array_44_62_real;
      end
      default : begin
        _zz_4522_ = int_reg_array_44_63_imag;
        _zz_4523_ = int_reg_array_44_63_real;
      end
    endcase
  end

  always @(*) begin
    case(_zz_3122_)
      6'b000000 : begin
        _zz_4524_ = int_reg_array_45_0_imag;
        _zz_4525_ = int_reg_array_45_0_real;
      end
      6'b000001 : begin
        _zz_4524_ = int_reg_array_45_1_imag;
        _zz_4525_ = int_reg_array_45_1_real;
      end
      6'b000010 : begin
        _zz_4524_ = int_reg_array_45_2_imag;
        _zz_4525_ = int_reg_array_45_2_real;
      end
      6'b000011 : begin
        _zz_4524_ = int_reg_array_45_3_imag;
        _zz_4525_ = int_reg_array_45_3_real;
      end
      6'b000100 : begin
        _zz_4524_ = int_reg_array_45_4_imag;
        _zz_4525_ = int_reg_array_45_4_real;
      end
      6'b000101 : begin
        _zz_4524_ = int_reg_array_45_5_imag;
        _zz_4525_ = int_reg_array_45_5_real;
      end
      6'b000110 : begin
        _zz_4524_ = int_reg_array_45_6_imag;
        _zz_4525_ = int_reg_array_45_6_real;
      end
      6'b000111 : begin
        _zz_4524_ = int_reg_array_45_7_imag;
        _zz_4525_ = int_reg_array_45_7_real;
      end
      6'b001000 : begin
        _zz_4524_ = int_reg_array_45_8_imag;
        _zz_4525_ = int_reg_array_45_8_real;
      end
      6'b001001 : begin
        _zz_4524_ = int_reg_array_45_9_imag;
        _zz_4525_ = int_reg_array_45_9_real;
      end
      6'b001010 : begin
        _zz_4524_ = int_reg_array_45_10_imag;
        _zz_4525_ = int_reg_array_45_10_real;
      end
      6'b001011 : begin
        _zz_4524_ = int_reg_array_45_11_imag;
        _zz_4525_ = int_reg_array_45_11_real;
      end
      6'b001100 : begin
        _zz_4524_ = int_reg_array_45_12_imag;
        _zz_4525_ = int_reg_array_45_12_real;
      end
      6'b001101 : begin
        _zz_4524_ = int_reg_array_45_13_imag;
        _zz_4525_ = int_reg_array_45_13_real;
      end
      6'b001110 : begin
        _zz_4524_ = int_reg_array_45_14_imag;
        _zz_4525_ = int_reg_array_45_14_real;
      end
      6'b001111 : begin
        _zz_4524_ = int_reg_array_45_15_imag;
        _zz_4525_ = int_reg_array_45_15_real;
      end
      6'b010000 : begin
        _zz_4524_ = int_reg_array_45_16_imag;
        _zz_4525_ = int_reg_array_45_16_real;
      end
      6'b010001 : begin
        _zz_4524_ = int_reg_array_45_17_imag;
        _zz_4525_ = int_reg_array_45_17_real;
      end
      6'b010010 : begin
        _zz_4524_ = int_reg_array_45_18_imag;
        _zz_4525_ = int_reg_array_45_18_real;
      end
      6'b010011 : begin
        _zz_4524_ = int_reg_array_45_19_imag;
        _zz_4525_ = int_reg_array_45_19_real;
      end
      6'b010100 : begin
        _zz_4524_ = int_reg_array_45_20_imag;
        _zz_4525_ = int_reg_array_45_20_real;
      end
      6'b010101 : begin
        _zz_4524_ = int_reg_array_45_21_imag;
        _zz_4525_ = int_reg_array_45_21_real;
      end
      6'b010110 : begin
        _zz_4524_ = int_reg_array_45_22_imag;
        _zz_4525_ = int_reg_array_45_22_real;
      end
      6'b010111 : begin
        _zz_4524_ = int_reg_array_45_23_imag;
        _zz_4525_ = int_reg_array_45_23_real;
      end
      6'b011000 : begin
        _zz_4524_ = int_reg_array_45_24_imag;
        _zz_4525_ = int_reg_array_45_24_real;
      end
      6'b011001 : begin
        _zz_4524_ = int_reg_array_45_25_imag;
        _zz_4525_ = int_reg_array_45_25_real;
      end
      6'b011010 : begin
        _zz_4524_ = int_reg_array_45_26_imag;
        _zz_4525_ = int_reg_array_45_26_real;
      end
      6'b011011 : begin
        _zz_4524_ = int_reg_array_45_27_imag;
        _zz_4525_ = int_reg_array_45_27_real;
      end
      6'b011100 : begin
        _zz_4524_ = int_reg_array_45_28_imag;
        _zz_4525_ = int_reg_array_45_28_real;
      end
      6'b011101 : begin
        _zz_4524_ = int_reg_array_45_29_imag;
        _zz_4525_ = int_reg_array_45_29_real;
      end
      6'b011110 : begin
        _zz_4524_ = int_reg_array_45_30_imag;
        _zz_4525_ = int_reg_array_45_30_real;
      end
      6'b011111 : begin
        _zz_4524_ = int_reg_array_45_31_imag;
        _zz_4525_ = int_reg_array_45_31_real;
      end
      6'b100000 : begin
        _zz_4524_ = int_reg_array_45_32_imag;
        _zz_4525_ = int_reg_array_45_32_real;
      end
      6'b100001 : begin
        _zz_4524_ = int_reg_array_45_33_imag;
        _zz_4525_ = int_reg_array_45_33_real;
      end
      6'b100010 : begin
        _zz_4524_ = int_reg_array_45_34_imag;
        _zz_4525_ = int_reg_array_45_34_real;
      end
      6'b100011 : begin
        _zz_4524_ = int_reg_array_45_35_imag;
        _zz_4525_ = int_reg_array_45_35_real;
      end
      6'b100100 : begin
        _zz_4524_ = int_reg_array_45_36_imag;
        _zz_4525_ = int_reg_array_45_36_real;
      end
      6'b100101 : begin
        _zz_4524_ = int_reg_array_45_37_imag;
        _zz_4525_ = int_reg_array_45_37_real;
      end
      6'b100110 : begin
        _zz_4524_ = int_reg_array_45_38_imag;
        _zz_4525_ = int_reg_array_45_38_real;
      end
      6'b100111 : begin
        _zz_4524_ = int_reg_array_45_39_imag;
        _zz_4525_ = int_reg_array_45_39_real;
      end
      6'b101000 : begin
        _zz_4524_ = int_reg_array_45_40_imag;
        _zz_4525_ = int_reg_array_45_40_real;
      end
      6'b101001 : begin
        _zz_4524_ = int_reg_array_45_41_imag;
        _zz_4525_ = int_reg_array_45_41_real;
      end
      6'b101010 : begin
        _zz_4524_ = int_reg_array_45_42_imag;
        _zz_4525_ = int_reg_array_45_42_real;
      end
      6'b101011 : begin
        _zz_4524_ = int_reg_array_45_43_imag;
        _zz_4525_ = int_reg_array_45_43_real;
      end
      6'b101100 : begin
        _zz_4524_ = int_reg_array_45_44_imag;
        _zz_4525_ = int_reg_array_45_44_real;
      end
      6'b101101 : begin
        _zz_4524_ = int_reg_array_45_45_imag;
        _zz_4525_ = int_reg_array_45_45_real;
      end
      6'b101110 : begin
        _zz_4524_ = int_reg_array_45_46_imag;
        _zz_4525_ = int_reg_array_45_46_real;
      end
      6'b101111 : begin
        _zz_4524_ = int_reg_array_45_47_imag;
        _zz_4525_ = int_reg_array_45_47_real;
      end
      6'b110000 : begin
        _zz_4524_ = int_reg_array_45_48_imag;
        _zz_4525_ = int_reg_array_45_48_real;
      end
      6'b110001 : begin
        _zz_4524_ = int_reg_array_45_49_imag;
        _zz_4525_ = int_reg_array_45_49_real;
      end
      6'b110010 : begin
        _zz_4524_ = int_reg_array_45_50_imag;
        _zz_4525_ = int_reg_array_45_50_real;
      end
      6'b110011 : begin
        _zz_4524_ = int_reg_array_45_51_imag;
        _zz_4525_ = int_reg_array_45_51_real;
      end
      6'b110100 : begin
        _zz_4524_ = int_reg_array_45_52_imag;
        _zz_4525_ = int_reg_array_45_52_real;
      end
      6'b110101 : begin
        _zz_4524_ = int_reg_array_45_53_imag;
        _zz_4525_ = int_reg_array_45_53_real;
      end
      6'b110110 : begin
        _zz_4524_ = int_reg_array_45_54_imag;
        _zz_4525_ = int_reg_array_45_54_real;
      end
      6'b110111 : begin
        _zz_4524_ = int_reg_array_45_55_imag;
        _zz_4525_ = int_reg_array_45_55_real;
      end
      6'b111000 : begin
        _zz_4524_ = int_reg_array_45_56_imag;
        _zz_4525_ = int_reg_array_45_56_real;
      end
      6'b111001 : begin
        _zz_4524_ = int_reg_array_45_57_imag;
        _zz_4525_ = int_reg_array_45_57_real;
      end
      6'b111010 : begin
        _zz_4524_ = int_reg_array_45_58_imag;
        _zz_4525_ = int_reg_array_45_58_real;
      end
      6'b111011 : begin
        _zz_4524_ = int_reg_array_45_59_imag;
        _zz_4525_ = int_reg_array_45_59_real;
      end
      6'b111100 : begin
        _zz_4524_ = int_reg_array_45_60_imag;
        _zz_4525_ = int_reg_array_45_60_real;
      end
      6'b111101 : begin
        _zz_4524_ = int_reg_array_45_61_imag;
        _zz_4525_ = int_reg_array_45_61_real;
      end
      6'b111110 : begin
        _zz_4524_ = int_reg_array_45_62_imag;
        _zz_4525_ = int_reg_array_45_62_real;
      end
      default : begin
        _zz_4524_ = int_reg_array_45_63_imag;
        _zz_4525_ = int_reg_array_45_63_real;
      end
    endcase
  end

  always @(*) begin
    case(_zz_3191_)
      6'b000000 : begin
        _zz_4526_ = int_reg_array_46_0_imag;
        _zz_4527_ = int_reg_array_46_0_real;
      end
      6'b000001 : begin
        _zz_4526_ = int_reg_array_46_1_imag;
        _zz_4527_ = int_reg_array_46_1_real;
      end
      6'b000010 : begin
        _zz_4526_ = int_reg_array_46_2_imag;
        _zz_4527_ = int_reg_array_46_2_real;
      end
      6'b000011 : begin
        _zz_4526_ = int_reg_array_46_3_imag;
        _zz_4527_ = int_reg_array_46_3_real;
      end
      6'b000100 : begin
        _zz_4526_ = int_reg_array_46_4_imag;
        _zz_4527_ = int_reg_array_46_4_real;
      end
      6'b000101 : begin
        _zz_4526_ = int_reg_array_46_5_imag;
        _zz_4527_ = int_reg_array_46_5_real;
      end
      6'b000110 : begin
        _zz_4526_ = int_reg_array_46_6_imag;
        _zz_4527_ = int_reg_array_46_6_real;
      end
      6'b000111 : begin
        _zz_4526_ = int_reg_array_46_7_imag;
        _zz_4527_ = int_reg_array_46_7_real;
      end
      6'b001000 : begin
        _zz_4526_ = int_reg_array_46_8_imag;
        _zz_4527_ = int_reg_array_46_8_real;
      end
      6'b001001 : begin
        _zz_4526_ = int_reg_array_46_9_imag;
        _zz_4527_ = int_reg_array_46_9_real;
      end
      6'b001010 : begin
        _zz_4526_ = int_reg_array_46_10_imag;
        _zz_4527_ = int_reg_array_46_10_real;
      end
      6'b001011 : begin
        _zz_4526_ = int_reg_array_46_11_imag;
        _zz_4527_ = int_reg_array_46_11_real;
      end
      6'b001100 : begin
        _zz_4526_ = int_reg_array_46_12_imag;
        _zz_4527_ = int_reg_array_46_12_real;
      end
      6'b001101 : begin
        _zz_4526_ = int_reg_array_46_13_imag;
        _zz_4527_ = int_reg_array_46_13_real;
      end
      6'b001110 : begin
        _zz_4526_ = int_reg_array_46_14_imag;
        _zz_4527_ = int_reg_array_46_14_real;
      end
      6'b001111 : begin
        _zz_4526_ = int_reg_array_46_15_imag;
        _zz_4527_ = int_reg_array_46_15_real;
      end
      6'b010000 : begin
        _zz_4526_ = int_reg_array_46_16_imag;
        _zz_4527_ = int_reg_array_46_16_real;
      end
      6'b010001 : begin
        _zz_4526_ = int_reg_array_46_17_imag;
        _zz_4527_ = int_reg_array_46_17_real;
      end
      6'b010010 : begin
        _zz_4526_ = int_reg_array_46_18_imag;
        _zz_4527_ = int_reg_array_46_18_real;
      end
      6'b010011 : begin
        _zz_4526_ = int_reg_array_46_19_imag;
        _zz_4527_ = int_reg_array_46_19_real;
      end
      6'b010100 : begin
        _zz_4526_ = int_reg_array_46_20_imag;
        _zz_4527_ = int_reg_array_46_20_real;
      end
      6'b010101 : begin
        _zz_4526_ = int_reg_array_46_21_imag;
        _zz_4527_ = int_reg_array_46_21_real;
      end
      6'b010110 : begin
        _zz_4526_ = int_reg_array_46_22_imag;
        _zz_4527_ = int_reg_array_46_22_real;
      end
      6'b010111 : begin
        _zz_4526_ = int_reg_array_46_23_imag;
        _zz_4527_ = int_reg_array_46_23_real;
      end
      6'b011000 : begin
        _zz_4526_ = int_reg_array_46_24_imag;
        _zz_4527_ = int_reg_array_46_24_real;
      end
      6'b011001 : begin
        _zz_4526_ = int_reg_array_46_25_imag;
        _zz_4527_ = int_reg_array_46_25_real;
      end
      6'b011010 : begin
        _zz_4526_ = int_reg_array_46_26_imag;
        _zz_4527_ = int_reg_array_46_26_real;
      end
      6'b011011 : begin
        _zz_4526_ = int_reg_array_46_27_imag;
        _zz_4527_ = int_reg_array_46_27_real;
      end
      6'b011100 : begin
        _zz_4526_ = int_reg_array_46_28_imag;
        _zz_4527_ = int_reg_array_46_28_real;
      end
      6'b011101 : begin
        _zz_4526_ = int_reg_array_46_29_imag;
        _zz_4527_ = int_reg_array_46_29_real;
      end
      6'b011110 : begin
        _zz_4526_ = int_reg_array_46_30_imag;
        _zz_4527_ = int_reg_array_46_30_real;
      end
      6'b011111 : begin
        _zz_4526_ = int_reg_array_46_31_imag;
        _zz_4527_ = int_reg_array_46_31_real;
      end
      6'b100000 : begin
        _zz_4526_ = int_reg_array_46_32_imag;
        _zz_4527_ = int_reg_array_46_32_real;
      end
      6'b100001 : begin
        _zz_4526_ = int_reg_array_46_33_imag;
        _zz_4527_ = int_reg_array_46_33_real;
      end
      6'b100010 : begin
        _zz_4526_ = int_reg_array_46_34_imag;
        _zz_4527_ = int_reg_array_46_34_real;
      end
      6'b100011 : begin
        _zz_4526_ = int_reg_array_46_35_imag;
        _zz_4527_ = int_reg_array_46_35_real;
      end
      6'b100100 : begin
        _zz_4526_ = int_reg_array_46_36_imag;
        _zz_4527_ = int_reg_array_46_36_real;
      end
      6'b100101 : begin
        _zz_4526_ = int_reg_array_46_37_imag;
        _zz_4527_ = int_reg_array_46_37_real;
      end
      6'b100110 : begin
        _zz_4526_ = int_reg_array_46_38_imag;
        _zz_4527_ = int_reg_array_46_38_real;
      end
      6'b100111 : begin
        _zz_4526_ = int_reg_array_46_39_imag;
        _zz_4527_ = int_reg_array_46_39_real;
      end
      6'b101000 : begin
        _zz_4526_ = int_reg_array_46_40_imag;
        _zz_4527_ = int_reg_array_46_40_real;
      end
      6'b101001 : begin
        _zz_4526_ = int_reg_array_46_41_imag;
        _zz_4527_ = int_reg_array_46_41_real;
      end
      6'b101010 : begin
        _zz_4526_ = int_reg_array_46_42_imag;
        _zz_4527_ = int_reg_array_46_42_real;
      end
      6'b101011 : begin
        _zz_4526_ = int_reg_array_46_43_imag;
        _zz_4527_ = int_reg_array_46_43_real;
      end
      6'b101100 : begin
        _zz_4526_ = int_reg_array_46_44_imag;
        _zz_4527_ = int_reg_array_46_44_real;
      end
      6'b101101 : begin
        _zz_4526_ = int_reg_array_46_45_imag;
        _zz_4527_ = int_reg_array_46_45_real;
      end
      6'b101110 : begin
        _zz_4526_ = int_reg_array_46_46_imag;
        _zz_4527_ = int_reg_array_46_46_real;
      end
      6'b101111 : begin
        _zz_4526_ = int_reg_array_46_47_imag;
        _zz_4527_ = int_reg_array_46_47_real;
      end
      6'b110000 : begin
        _zz_4526_ = int_reg_array_46_48_imag;
        _zz_4527_ = int_reg_array_46_48_real;
      end
      6'b110001 : begin
        _zz_4526_ = int_reg_array_46_49_imag;
        _zz_4527_ = int_reg_array_46_49_real;
      end
      6'b110010 : begin
        _zz_4526_ = int_reg_array_46_50_imag;
        _zz_4527_ = int_reg_array_46_50_real;
      end
      6'b110011 : begin
        _zz_4526_ = int_reg_array_46_51_imag;
        _zz_4527_ = int_reg_array_46_51_real;
      end
      6'b110100 : begin
        _zz_4526_ = int_reg_array_46_52_imag;
        _zz_4527_ = int_reg_array_46_52_real;
      end
      6'b110101 : begin
        _zz_4526_ = int_reg_array_46_53_imag;
        _zz_4527_ = int_reg_array_46_53_real;
      end
      6'b110110 : begin
        _zz_4526_ = int_reg_array_46_54_imag;
        _zz_4527_ = int_reg_array_46_54_real;
      end
      6'b110111 : begin
        _zz_4526_ = int_reg_array_46_55_imag;
        _zz_4527_ = int_reg_array_46_55_real;
      end
      6'b111000 : begin
        _zz_4526_ = int_reg_array_46_56_imag;
        _zz_4527_ = int_reg_array_46_56_real;
      end
      6'b111001 : begin
        _zz_4526_ = int_reg_array_46_57_imag;
        _zz_4527_ = int_reg_array_46_57_real;
      end
      6'b111010 : begin
        _zz_4526_ = int_reg_array_46_58_imag;
        _zz_4527_ = int_reg_array_46_58_real;
      end
      6'b111011 : begin
        _zz_4526_ = int_reg_array_46_59_imag;
        _zz_4527_ = int_reg_array_46_59_real;
      end
      6'b111100 : begin
        _zz_4526_ = int_reg_array_46_60_imag;
        _zz_4527_ = int_reg_array_46_60_real;
      end
      6'b111101 : begin
        _zz_4526_ = int_reg_array_46_61_imag;
        _zz_4527_ = int_reg_array_46_61_real;
      end
      6'b111110 : begin
        _zz_4526_ = int_reg_array_46_62_imag;
        _zz_4527_ = int_reg_array_46_62_real;
      end
      default : begin
        _zz_4526_ = int_reg_array_46_63_imag;
        _zz_4527_ = int_reg_array_46_63_real;
      end
    endcase
  end

  always @(*) begin
    case(_zz_3260_)
      6'b000000 : begin
        _zz_4528_ = int_reg_array_47_0_imag;
        _zz_4529_ = int_reg_array_47_0_real;
      end
      6'b000001 : begin
        _zz_4528_ = int_reg_array_47_1_imag;
        _zz_4529_ = int_reg_array_47_1_real;
      end
      6'b000010 : begin
        _zz_4528_ = int_reg_array_47_2_imag;
        _zz_4529_ = int_reg_array_47_2_real;
      end
      6'b000011 : begin
        _zz_4528_ = int_reg_array_47_3_imag;
        _zz_4529_ = int_reg_array_47_3_real;
      end
      6'b000100 : begin
        _zz_4528_ = int_reg_array_47_4_imag;
        _zz_4529_ = int_reg_array_47_4_real;
      end
      6'b000101 : begin
        _zz_4528_ = int_reg_array_47_5_imag;
        _zz_4529_ = int_reg_array_47_5_real;
      end
      6'b000110 : begin
        _zz_4528_ = int_reg_array_47_6_imag;
        _zz_4529_ = int_reg_array_47_6_real;
      end
      6'b000111 : begin
        _zz_4528_ = int_reg_array_47_7_imag;
        _zz_4529_ = int_reg_array_47_7_real;
      end
      6'b001000 : begin
        _zz_4528_ = int_reg_array_47_8_imag;
        _zz_4529_ = int_reg_array_47_8_real;
      end
      6'b001001 : begin
        _zz_4528_ = int_reg_array_47_9_imag;
        _zz_4529_ = int_reg_array_47_9_real;
      end
      6'b001010 : begin
        _zz_4528_ = int_reg_array_47_10_imag;
        _zz_4529_ = int_reg_array_47_10_real;
      end
      6'b001011 : begin
        _zz_4528_ = int_reg_array_47_11_imag;
        _zz_4529_ = int_reg_array_47_11_real;
      end
      6'b001100 : begin
        _zz_4528_ = int_reg_array_47_12_imag;
        _zz_4529_ = int_reg_array_47_12_real;
      end
      6'b001101 : begin
        _zz_4528_ = int_reg_array_47_13_imag;
        _zz_4529_ = int_reg_array_47_13_real;
      end
      6'b001110 : begin
        _zz_4528_ = int_reg_array_47_14_imag;
        _zz_4529_ = int_reg_array_47_14_real;
      end
      6'b001111 : begin
        _zz_4528_ = int_reg_array_47_15_imag;
        _zz_4529_ = int_reg_array_47_15_real;
      end
      6'b010000 : begin
        _zz_4528_ = int_reg_array_47_16_imag;
        _zz_4529_ = int_reg_array_47_16_real;
      end
      6'b010001 : begin
        _zz_4528_ = int_reg_array_47_17_imag;
        _zz_4529_ = int_reg_array_47_17_real;
      end
      6'b010010 : begin
        _zz_4528_ = int_reg_array_47_18_imag;
        _zz_4529_ = int_reg_array_47_18_real;
      end
      6'b010011 : begin
        _zz_4528_ = int_reg_array_47_19_imag;
        _zz_4529_ = int_reg_array_47_19_real;
      end
      6'b010100 : begin
        _zz_4528_ = int_reg_array_47_20_imag;
        _zz_4529_ = int_reg_array_47_20_real;
      end
      6'b010101 : begin
        _zz_4528_ = int_reg_array_47_21_imag;
        _zz_4529_ = int_reg_array_47_21_real;
      end
      6'b010110 : begin
        _zz_4528_ = int_reg_array_47_22_imag;
        _zz_4529_ = int_reg_array_47_22_real;
      end
      6'b010111 : begin
        _zz_4528_ = int_reg_array_47_23_imag;
        _zz_4529_ = int_reg_array_47_23_real;
      end
      6'b011000 : begin
        _zz_4528_ = int_reg_array_47_24_imag;
        _zz_4529_ = int_reg_array_47_24_real;
      end
      6'b011001 : begin
        _zz_4528_ = int_reg_array_47_25_imag;
        _zz_4529_ = int_reg_array_47_25_real;
      end
      6'b011010 : begin
        _zz_4528_ = int_reg_array_47_26_imag;
        _zz_4529_ = int_reg_array_47_26_real;
      end
      6'b011011 : begin
        _zz_4528_ = int_reg_array_47_27_imag;
        _zz_4529_ = int_reg_array_47_27_real;
      end
      6'b011100 : begin
        _zz_4528_ = int_reg_array_47_28_imag;
        _zz_4529_ = int_reg_array_47_28_real;
      end
      6'b011101 : begin
        _zz_4528_ = int_reg_array_47_29_imag;
        _zz_4529_ = int_reg_array_47_29_real;
      end
      6'b011110 : begin
        _zz_4528_ = int_reg_array_47_30_imag;
        _zz_4529_ = int_reg_array_47_30_real;
      end
      6'b011111 : begin
        _zz_4528_ = int_reg_array_47_31_imag;
        _zz_4529_ = int_reg_array_47_31_real;
      end
      6'b100000 : begin
        _zz_4528_ = int_reg_array_47_32_imag;
        _zz_4529_ = int_reg_array_47_32_real;
      end
      6'b100001 : begin
        _zz_4528_ = int_reg_array_47_33_imag;
        _zz_4529_ = int_reg_array_47_33_real;
      end
      6'b100010 : begin
        _zz_4528_ = int_reg_array_47_34_imag;
        _zz_4529_ = int_reg_array_47_34_real;
      end
      6'b100011 : begin
        _zz_4528_ = int_reg_array_47_35_imag;
        _zz_4529_ = int_reg_array_47_35_real;
      end
      6'b100100 : begin
        _zz_4528_ = int_reg_array_47_36_imag;
        _zz_4529_ = int_reg_array_47_36_real;
      end
      6'b100101 : begin
        _zz_4528_ = int_reg_array_47_37_imag;
        _zz_4529_ = int_reg_array_47_37_real;
      end
      6'b100110 : begin
        _zz_4528_ = int_reg_array_47_38_imag;
        _zz_4529_ = int_reg_array_47_38_real;
      end
      6'b100111 : begin
        _zz_4528_ = int_reg_array_47_39_imag;
        _zz_4529_ = int_reg_array_47_39_real;
      end
      6'b101000 : begin
        _zz_4528_ = int_reg_array_47_40_imag;
        _zz_4529_ = int_reg_array_47_40_real;
      end
      6'b101001 : begin
        _zz_4528_ = int_reg_array_47_41_imag;
        _zz_4529_ = int_reg_array_47_41_real;
      end
      6'b101010 : begin
        _zz_4528_ = int_reg_array_47_42_imag;
        _zz_4529_ = int_reg_array_47_42_real;
      end
      6'b101011 : begin
        _zz_4528_ = int_reg_array_47_43_imag;
        _zz_4529_ = int_reg_array_47_43_real;
      end
      6'b101100 : begin
        _zz_4528_ = int_reg_array_47_44_imag;
        _zz_4529_ = int_reg_array_47_44_real;
      end
      6'b101101 : begin
        _zz_4528_ = int_reg_array_47_45_imag;
        _zz_4529_ = int_reg_array_47_45_real;
      end
      6'b101110 : begin
        _zz_4528_ = int_reg_array_47_46_imag;
        _zz_4529_ = int_reg_array_47_46_real;
      end
      6'b101111 : begin
        _zz_4528_ = int_reg_array_47_47_imag;
        _zz_4529_ = int_reg_array_47_47_real;
      end
      6'b110000 : begin
        _zz_4528_ = int_reg_array_47_48_imag;
        _zz_4529_ = int_reg_array_47_48_real;
      end
      6'b110001 : begin
        _zz_4528_ = int_reg_array_47_49_imag;
        _zz_4529_ = int_reg_array_47_49_real;
      end
      6'b110010 : begin
        _zz_4528_ = int_reg_array_47_50_imag;
        _zz_4529_ = int_reg_array_47_50_real;
      end
      6'b110011 : begin
        _zz_4528_ = int_reg_array_47_51_imag;
        _zz_4529_ = int_reg_array_47_51_real;
      end
      6'b110100 : begin
        _zz_4528_ = int_reg_array_47_52_imag;
        _zz_4529_ = int_reg_array_47_52_real;
      end
      6'b110101 : begin
        _zz_4528_ = int_reg_array_47_53_imag;
        _zz_4529_ = int_reg_array_47_53_real;
      end
      6'b110110 : begin
        _zz_4528_ = int_reg_array_47_54_imag;
        _zz_4529_ = int_reg_array_47_54_real;
      end
      6'b110111 : begin
        _zz_4528_ = int_reg_array_47_55_imag;
        _zz_4529_ = int_reg_array_47_55_real;
      end
      6'b111000 : begin
        _zz_4528_ = int_reg_array_47_56_imag;
        _zz_4529_ = int_reg_array_47_56_real;
      end
      6'b111001 : begin
        _zz_4528_ = int_reg_array_47_57_imag;
        _zz_4529_ = int_reg_array_47_57_real;
      end
      6'b111010 : begin
        _zz_4528_ = int_reg_array_47_58_imag;
        _zz_4529_ = int_reg_array_47_58_real;
      end
      6'b111011 : begin
        _zz_4528_ = int_reg_array_47_59_imag;
        _zz_4529_ = int_reg_array_47_59_real;
      end
      6'b111100 : begin
        _zz_4528_ = int_reg_array_47_60_imag;
        _zz_4529_ = int_reg_array_47_60_real;
      end
      6'b111101 : begin
        _zz_4528_ = int_reg_array_47_61_imag;
        _zz_4529_ = int_reg_array_47_61_real;
      end
      6'b111110 : begin
        _zz_4528_ = int_reg_array_47_62_imag;
        _zz_4529_ = int_reg_array_47_62_real;
      end
      default : begin
        _zz_4528_ = int_reg_array_47_63_imag;
        _zz_4529_ = int_reg_array_47_63_real;
      end
    endcase
  end

  always @(*) begin
    case(_zz_3329_)
      6'b000000 : begin
        _zz_4530_ = int_reg_array_48_0_imag;
        _zz_4531_ = int_reg_array_48_0_real;
      end
      6'b000001 : begin
        _zz_4530_ = int_reg_array_48_1_imag;
        _zz_4531_ = int_reg_array_48_1_real;
      end
      6'b000010 : begin
        _zz_4530_ = int_reg_array_48_2_imag;
        _zz_4531_ = int_reg_array_48_2_real;
      end
      6'b000011 : begin
        _zz_4530_ = int_reg_array_48_3_imag;
        _zz_4531_ = int_reg_array_48_3_real;
      end
      6'b000100 : begin
        _zz_4530_ = int_reg_array_48_4_imag;
        _zz_4531_ = int_reg_array_48_4_real;
      end
      6'b000101 : begin
        _zz_4530_ = int_reg_array_48_5_imag;
        _zz_4531_ = int_reg_array_48_5_real;
      end
      6'b000110 : begin
        _zz_4530_ = int_reg_array_48_6_imag;
        _zz_4531_ = int_reg_array_48_6_real;
      end
      6'b000111 : begin
        _zz_4530_ = int_reg_array_48_7_imag;
        _zz_4531_ = int_reg_array_48_7_real;
      end
      6'b001000 : begin
        _zz_4530_ = int_reg_array_48_8_imag;
        _zz_4531_ = int_reg_array_48_8_real;
      end
      6'b001001 : begin
        _zz_4530_ = int_reg_array_48_9_imag;
        _zz_4531_ = int_reg_array_48_9_real;
      end
      6'b001010 : begin
        _zz_4530_ = int_reg_array_48_10_imag;
        _zz_4531_ = int_reg_array_48_10_real;
      end
      6'b001011 : begin
        _zz_4530_ = int_reg_array_48_11_imag;
        _zz_4531_ = int_reg_array_48_11_real;
      end
      6'b001100 : begin
        _zz_4530_ = int_reg_array_48_12_imag;
        _zz_4531_ = int_reg_array_48_12_real;
      end
      6'b001101 : begin
        _zz_4530_ = int_reg_array_48_13_imag;
        _zz_4531_ = int_reg_array_48_13_real;
      end
      6'b001110 : begin
        _zz_4530_ = int_reg_array_48_14_imag;
        _zz_4531_ = int_reg_array_48_14_real;
      end
      6'b001111 : begin
        _zz_4530_ = int_reg_array_48_15_imag;
        _zz_4531_ = int_reg_array_48_15_real;
      end
      6'b010000 : begin
        _zz_4530_ = int_reg_array_48_16_imag;
        _zz_4531_ = int_reg_array_48_16_real;
      end
      6'b010001 : begin
        _zz_4530_ = int_reg_array_48_17_imag;
        _zz_4531_ = int_reg_array_48_17_real;
      end
      6'b010010 : begin
        _zz_4530_ = int_reg_array_48_18_imag;
        _zz_4531_ = int_reg_array_48_18_real;
      end
      6'b010011 : begin
        _zz_4530_ = int_reg_array_48_19_imag;
        _zz_4531_ = int_reg_array_48_19_real;
      end
      6'b010100 : begin
        _zz_4530_ = int_reg_array_48_20_imag;
        _zz_4531_ = int_reg_array_48_20_real;
      end
      6'b010101 : begin
        _zz_4530_ = int_reg_array_48_21_imag;
        _zz_4531_ = int_reg_array_48_21_real;
      end
      6'b010110 : begin
        _zz_4530_ = int_reg_array_48_22_imag;
        _zz_4531_ = int_reg_array_48_22_real;
      end
      6'b010111 : begin
        _zz_4530_ = int_reg_array_48_23_imag;
        _zz_4531_ = int_reg_array_48_23_real;
      end
      6'b011000 : begin
        _zz_4530_ = int_reg_array_48_24_imag;
        _zz_4531_ = int_reg_array_48_24_real;
      end
      6'b011001 : begin
        _zz_4530_ = int_reg_array_48_25_imag;
        _zz_4531_ = int_reg_array_48_25_real;
      end
      6'b011010 : begin
        _zz_4530_ = int_reg_array_48_26_imag;
        _zz_4531_ = int_reg_array_48_26_real;
      end
      6'b011011 : begin
        _zz_4530_ = int_reg_array_48_27_imag;
        _zz_4531_ = int_reg_array_48_27_real;
      end
      6'b011100 : begin
        _zz_4530_ = int_reg_array_48_28_imag;
        _zz_4531_ = int_reg_array_48_28_real;
      end
      6'b011101 : begin
        _zz_4530_ = int_reg_array_48_29_imag;
        _zz_4531_ = int_reg_array_48_29_real;
      end
      6'b011110 : begin
        _zz_4530_ = int_reg_array_48_30_imag;
        _zz_4531_ = int_reg_array_48_30_real;
      end
      6'b011111 : begin
        _zz_4530_ = int_reg_array_48_31_imag;
        _zz_4531_ = int_reg_array_48_31_real;
      end
      6'b100000 : begin
        _zz_4530_ = int_reg_array_48_32_imag;
        _zz_4531_ = int_reg_array_48_32_real;
      end
      6'b100001 : begin
        _zz_4530_ = int_reg_array_48_33_imag;
        _zz_4531_ = int_reg_array_48_33_real;
      end
      6'b100010 : begin
        _zz_4530_ = int_reg_array_48_34_imag;
        _zz_4531_ = int_reg_array_48_34_real;
      end
      6'b100011 : begin
        _zz_4530_ = int_reg_array_48_35_imag;
        _zz_4531_ = int_reg_array_48_35_real;
      end
      6'b100100 : begin
        _zz_4530_ = int_reg_array_48_36_imag;
        _zz_4531_ = int_reg_array_48_36_real;
      end
      6'b100101 : begin
        _zz_4530_ = int_reg_array_48_37_imag;
        _zz_4531_ = int_reg_array_48_37_real;
      end
      6'b100110 : begin
        _zz_4530_ = int_reg_array_48_38_imag;
        _zz_4531_ = int_reg_array_48_38_real;
      end
      6'b100111 : begin
        _zz_4530_ = int_reg_array_48_39_imag;
        _zz_4531_ = int_reg_array_48_39_real;
      end
      6'b101000 : begin
        _zz_4530_ = int_reg_array_48_40_imag;
        _zz_4531_ = int_reg_array_48_40_real;
      end
      6'b101001 : begin
        _zz_4530_ = int_reg_array_48_41_imag;
        _zz_4531_ = int_reg_array_48_41_real;
      end
      6'b101010 : begin
        _zz_4530_ = int_reg_array_48_42_imag;
        _zz_4531_ = int_reg_array_48_42_real;
      end
      6'b101011 : begin
        _zz_4530_ = int_reg_array_48_43_imag;
        _zz_4531_ = int_reg_array_48_43_real;
      end
      6'b101100 : begin
        _zz_4530_ = int_reg_array_48_44_imag;
        _zz_4531_ = int_reg_array_48_44_real;
      end
      6'b101101 : begin
        _zz_4530_ = int_reg_array_48_45_imag;
        _zz_4531_ = int_reg_array_48_45_real;
      end
      6'b101110 : begin
        _zz_4530_ = int_reg_array_48_46_imag;
        _zz_4531_ = int_reg_array_48_46_real;
      end
      6'b101111 : begin
        _zz_4530_ = int_reg_array_48_47_imag;
        _zz_4531_ = int_reg_array_48_47_real;
      end
      6'b110000 : begin
        _zz_4530_ = int_reg_array_48_48_imag;
        _zz_4531_ = int_reg_array_48_48_real;
      end
      6'b110001 : begin
        _zz_4530_ = int_reg_array_48_49_imag;
        _zz_4531_ = int_reg_array_48_49_real;
      end
      6'b110010 : begin
        _zz_4530_ = int_reg_array_48_50_imag;
        _zz_4531_ = int_reg_array_48_50_real;
      end
      6'b110011 : begin
        _zz_4530_ = int_reg_array_48_51_imag;
        _zz_4531_ = int_reg_array_48_51_real;
      end
      6'b110100 : begin
        _zz_4530_ = int_reg_array_48_52_imag;
        _zz_4531_ = int_reg_array_48_52_real;
      end
      6'b110101 : begin
        _zz_4530_ = int_reg_array_48_53_imag;
        _zz_4531_ = int_reg_array_48_53_real;
      end
      6'b110110 : begin
        _zz_4530_ = int_reg_array_48_54_imag;
        _zz_4531_ = int_reg_array_48_54_real;
      end
      6'b110111 : begin
        _zz_4530_ = int_reg_array_48_55_imag;
        _zz_4531_ = int_reg_array_48_55_real;
      end
      6'b111000 : begin
        _zz_4530_ = int_reg_array_48_56_imag;
        _zz_4531_ = int_reg_array_48_56_real;
      end
      6'b111001 : begin
        _zz_4530_ = int_reg_array_48_57_imag;
        _zz_4531_ = int_reg_array_48_57_real;
      end
      6'b111010 : begin
        _zz_4530_ = int_reg_array_48_58_imag;
        _zz_4531_ = int_reg_array_48_58_real;
      end
      6'b111011 : begin
        _zz_4530_ = int_reg_array_48_59_imag;
        _zz_4531_ = int_reg_array_48_59_real;
      end
      6'b111100 : begin
        _zz_4530_ = int_reg_array_48_60_imag;
        _zz_4531_ = int_reg_array_48_60_real;
      end
      6'b111101 : begin
        _zz_4530_ = int_reg_array_48_61_imag;
        _zz_4531_ = int_reg_array_48_61_real;
      end
      6'b111110 : begin
        _zz_4530_ = int_reg_array_48_62_imag;
        _zz_4531_ = int_reg_array_48_62_real;
      end
      default : begin
        _zz_4530_ = int_reg_array_48_63_imag;
        _zz_4531_ = int_reg_array_48_63_real;
      end
    endcase
  end

  always @(*) begin
    case(_zz_3398_)
      6'b000000 : begin
        _zz_4532_ = int_reg_array_49_0_imag;
        _zz_4533_ = int_reg_array_49_0_real;
      end
      6'b000001 : begin
        _zz_4532_ = int_reg_array_49_1_imag;
        _zz_4533_ = int_reg_array_49_1_real;
      end
      6'b000010 : begin
        _zz_4532_ = int_reg_array_49_2_imag;
        _zz_4533_ = int_reg_array_49_2_real;
      end
      6'b000011 : begin
        _zz_4532_ = int_reg_array_49_3_imag;
        _zz_4533_ = int_reg_array_49_3_real;
      end
      6'b000100 : begin
        _zz_4532_ = int_reg_array_49_4_imag;
        _zz_4533_ = int_reg_array_49_4_real;
      end
      6'b000101 : begin
        _zz_4532_ = int_reg_array_49_5_imag;
        _zz_4533_ = int_reg_array_49_5_real;
      end
      6'b000110 : begin
        _zz_4532_ = int_reg_array_49_6_imag;
        _zz_4533_ = int_reg_array_49_6_real;
      end
      6'b000111 : begin
        _zz_4532_ = int_reg_array_49_7_imag;
        _zz_4533_ = int_reg_array_49_7_real;
      end
      6'b001000 : begin
        _zz_4532_ = int_reg_array_49_8_imag;
        _zz_4533_ = int_reg_array_49_8_real;
      end
      6'b001001 : begin
        _zz_4532_ = int_reg_array_49_9_imag;
        _zz_4533_ = int_reg_array_49_9_real;
      end
      6'b001010 : begin
        _zz_4532_ = int_reg_array_49_10_imag;
        _zz_4533_ = int_reg_array_49_10_real;
      end
      6'b001011 : begin
        _zz_4532_ = int_reg_array_49_11_imag;
        _zz_4533_ = int_reg_array_49_11_real;
      end
      6'b001100 : begin
        _zz_4532_ = int_reg_array_49_12_imag;
        _zz_4533_ = int_reg_array_49_12_real;
      end
      6'b001101 : begin
        _zz_4532_ = int_reg_array_49_13_imag;
        _zz_4533_ = int_reg_array_49_13_real;
      end
      6'b001110 : begin
        _zz_4532_ = int_reg_array_49_14_imag;
        _zz_4533_ = int_reg_array_49_14_real;
      end
      6'b001111 : begin
        _zz_4532_ = int_reg_array_49_15_imag;
        _zz_4533_ = int_reg_array_49_15_real;
      end
      6'b010000 : begin
        _zz_4532_ = int_reg_array_49_16_imag;
        _zz_4533_ = int_reg_array_49_16_real;
      end
      6'b010001 : begin
        _zz_4532_ = int_reg_array_49_17_imag;
        _zz_4533_ = int_reg_array_49_17_real;
      end
      6'b010010 : begin
        _zz_4532_ = int_reg_array_49_18_imag;
        _zz_4533_ = int_reg_array_49_18_real;
      end
      6'b010011 : begin
        _zz_4532_ = int_reg_array_49_19_imag;
        _zz_4533_ = int_reg_array_49_19_real;
      end
      6'b010100 : begin
        _zz_4532_ = int_reg_array_49_20_imag;
        _zz_4533_ = int_reg_array_49_20_real;
      end
      6'b010101 : begin
        _zz_4532_ = int_reg_array_49_21_imag;
        _zz_4533_ = int_reg_array_49_21_real;
      end
      6'b010110 : begin
        _zz_4532_ = int_reg_array_49_22_imag;
        _zz_4533_ = int_reg_array_49_22_real;
      end
      6'b010111 : begin
        _zz_4532_ = int_reg_array_49_23_imag;
        _zz_4533_ = int_reg_array_49_23_real;
      end
      6'b011000 : begin
        _zz_4532_ = int_reg_array_49_24_imag;
        _zz_4533_ = int_reg_array_49_24_real;
      end
      6'b011001 : begin
        _zz_4532_ = int_reg_array_49_25_imag;
        _zz_4533_ = int_reg_array_49_25_real;
      end
      6'b011010 : begin
        _zz_4532_ = int_reg_array_49_26_imag;
        _zz_4533_ = int_reg_array_49_26_real;
      end
      6'b011011 : begin
        _zz_4532_ = int_reg_array_49_27_imag;
        _zz_4533_ = int_reg_array_49_27_real;
      end
      6'b011100 : begin
        _zz_4532_ = int_reg_array_49_28_imag;
        _zz_4533_ = int_reg_array_49_28_real;
      end
      6'b011101 : begin
        _zz_4532_ = int_reg_array_49_29_imag;
        _zz_4533_ = int_reg_array_49_29_real;
      end
      6'b011110 : begin
        _zz_4532_ = int_reg_array_49_30_imag;
        _zz_4533_ = int_reg_array_49_30_real;
      end
      6'b011111 : begin
        _zz_4532_ = int_reg_array_49_31_imag;
        _zz_4533_ = int_reg_array_49_31_real;
      end
      6'b100000 : begin
        _zz_4532_ = int_reg_array_49_32_imag;
        _zz_4533_ = int_reg_array_49_32_real;
      end
      6'b100001 : begin
        _zz_4532_ = int_reg_array_49_33_imag;
        _zz_4533_ = int_reg_array_49_33_real;
      end
      6'b100010 : begin
        _zz_4532_ = int_reg_array_49_34_imag;
        _zz_4533_ = int_reg_array_49_34_real;
      end
      6'b100011 : begin
        _zz_4532_ = int_reg_array_49_35_imag;
        _zz_4533_ = int_reg_array_49_35_real;
      end
      6'b100100 : begin
        _zz_4532_ = int_reg_array_49_36_imag;
        _zz_4533_ = int_reg_array_49_36_real;
      end
      6'b100101 : begin
        _zz_4532_ = int_reg_array_49_37_imag;
        _zz_4533_ = int_reg_array_49_37_real;
      end
      6'b100110 : begin
        _zz_4532_ = int_reg_array_49_38_imag;
        _zz_4533_ = int_reg_array_49_38_real;
      end
      6'b100111 : begin
        _zz_4532_ = int_reg_array_49_39_imag;
        _zz_4533_ = int_reg_array_49_39_real;
      end
      6'b101000 : begin
        _zz_4532_ = int_reg_array_49_40_imag;
        _zz_4533_ = int_reg_array_49_40_real;
      end
      6'b101001 : begin
        _zz_4532_ = int_reg_array_49_41_imag;
        _zz_4533_ = int_reg_array_49_41_real;
      end
      6'b101010 : begin
        _zz_4532_ = int_reg_array_49_42_imag;
        _zz_4533_ = int_reg_array_49_42_real;
      end
      6'b101011 : begin
        _zz_4532_ = int_reg_array_49_43_imag;
        _zz_4533_ = int_reg_array_49_43_real;
      end
      6'b101100 : begin
        _zz_4532_ = int_reg_array_49_44_imag;
        _zz_4533_ = int_reg_array_49_44_real;
      end
      6'b101101 : begin
        _zz_4532_ = int_reg_array_49_45_imag;
        _zz_4533_ = int_reg_array_49_45_real;
      end
      6'b101110 : begin
        _zz_4532_ = int_reg_array_49_46_imag;
        _zz_4533_ = int_reg_array_49_46_real;
      end
      6'b101111 : begin
        _zz_4532_ = int_reg_array_49_47_imag;
        _zz_4533_ = int_reg_array_49_47_real;
      end
      6'b110000 : begin
        _zz_4532_ = int_reg_array_49_48_imag;
        _zz_4533_ = int_reg_array_49_48_real;
      end
      6'b110001 : begin
        _zz_4532_ = int_reg_array_49_49_imag;
        _zz_4533_ = int_reg_array_49_49_real;
      end
      6'b110010 : begin
        _zz_4532_ = int_reg_array_49_50_imag;
        _zz_4533_ = int_reg_array_49_50_real;
      end
      6'b110011 : begin
        _zz_4532_ = int_reg_array_49_51_imag;
        _zz_4533_ = int_reg_array_49_51_real;
      end
      6'b110100 : begin
        _zz_4532_ = int_reg_array_49_52_imag;
        _zz_4533_ = int_reg_array_49_52_real;
      end
      6'b110101 : begin
        _zz_4532_ = int_reg_array_49_53_imag;
        _zz_4533_ = int_reg_array_49_53_real;
      end
      6'b110110 : begin
        _zz_4532_ = int_reg_array_49_54_imag;
        _zz_4533_ = int_reg_array_49_54_real;
      end
      6'b110111 : begin
        _zz_4532_ = int_reg_array_49_55_imag;
        _zz_4533_ = int_reg_array_49_55_real;
      end
      6'b111000 : begin
        _zz_4532_ = int_reg_array_49_56_imag;
        _zz_4533_ = int_reg_array_49_56_real;
      end
      6'b111001 : begin
        _zz_4532_ = int_reg_array_49_57_imag;
        _zz_4533_ = int_reg_array_49_57_real;
      end
      6'b111010 : begin
        _zz_4532_ = int_reg_array_49_58_imag;
        _zz_4533_ = int_reg_array_49_58_real;
      end
      6'b111011 : begin
        _zz_4532_ = int_reg_array_49_59_imag;
        _zz_4533_ = int_reg_array_49_59_real;
      end
      6'b111100 : begin
        _zz_4532_ = int_reg_array_49_60_imag;
        _zz_4533_ = int_reg_array_49_60_real;
      end
      6'b111101 : begin
        _zz_4532_ = int_reg_array_49_61_imag;
        _zz_4533_ = int_reg_array_49_61_real;
      end
      6'b111110 : begin
        _zz_4532_ = int_reg_array_49_62_imag;
        _zz_4533_ = int_reg_array_49_62_real;
      end
      default : begin
        _zz_4532_ = int_reg_array_49_63_imag;
        _zz_4533_ = int_reg_array_49_63_real;
      end
    endcase
  end

  always @(*) begin
    case(_zz_3467_)
      6'b000000 : begin
        _zz_4534_ = int_reg_array_50_0_imag;
        _zz_4535_ = int_reg_array_50_0_real;
      end
      6'b000001 : begin
        _zz_4534_ = int_reg_array_50_1_imag;
        _zz_4535_ = int_reg_array_50_1_real;
      end
      6'b000010 : begin
        _zz_4534_ = int_reg_array_50_2_imag;
        _zz_4535_ = int_reg_array_50_2_real;
      end
      6'b000011 : begin
        _zz_4534_ = int_reg_array_50_3_imag;
        _zz_4535_ = int_reg_array_50_3_real;
      end
      6'b000100 : begin
        _zz_4534_ = int_reg_array_50_4_imag;
        _zz_4535_ = int_reg_array_50_4_real;
      end
      6'b000101 : begin
        _zz_4534_ = int_reg_array_50_5_imag;
        _zz_4535_ = int_reg_array_50_5_real;
      end
      6'b000110 : begin
        _zz_4534_ = int_reg_array_50_6_imag;
        _zz_4535_ = int_reg_array_50_6_real;
      end
      6'b000111 : begin
        _zz_4534_ = int_reg_array_50_7_imag;
        _zz_4535_ = int_reg_array_50_7_real;
      end
      6'b001000 : begin
        _zz_4534_ = int_reg_array_50_8_imag;
        _zz_4535_ = int_reg_array_50_8_real;
      end
      6'b001001 : begin
        _zz_4534_ = int_reg_array_50_9_imag;
        _zz_4535_ = int_reg_array_50_9_real;
      end
      6'b001010 : begin
        _zz_4534_ = int_reg_array_50_10_imag;
        _zz_4535_ = int_reg_array_50_10_real;
      end
      6'b001011 : begin
        _zz_4534_ = int_reg_array_50_11_imag;
        _zz_4535_ = int_reg_array_50_11_real;
      end
      6'b001100 : begin
        _zz_4534_ = int_reg_array_50_12_imag;
        _zz_4535_ = int_reg_array_50_12_real;
      end
      6'b001101 : begin
        _zz_4534_ = int_reg_array_50_13_imag;
        _zz_4535_ = int_reg_array_50_13_real;
      end
      6'b001110 : begin
        _zz_4534_ = int_reg_array_50_14_imag;
        _zz_4535_ = int_reg_array_50_14_real;
      end
      6'b001111 : begin
        _zz_4534_ = int_reg_array_50_15_imag;
        _zz_4535_ = int_reg_array_50_15_real;
      end
      6'b010000 : begin
        _zz_4534_ = int_reg_array_50_16_imag;
        _zz_4535_ = int_reg_array_50_16_real;
      end
      6'b010001 : begin
        _zz_4534_ = int_reg_array_50_17_imag;
        _zz_4535_ = int_reg_array_50_17_real;
      end
      6'b010010 : begin
        _zz_4534_ = int_reg_array_50_18_imag;
        _zz_4535_ = int_reg_array_50_18_real;
      end
      6'b010011 : begin
        _zz_4534_ = int_reg_array_50_19_imag;
        _zz_4535_ = int_reg_array_50_19_real;
      end
      6'b010100 : begin
        _zz_4534_ = int_reg_array_50_20_imag;
        _zz_4535_ = int_reg_array_50_20_real;
      end
      6'b010101 : begin
        _zz_4534_ = int_reg_array_50_21_imag;
        _zz_4535_ = int_reg_array_50_21_real;
      end
      6'b010110 : begin
        _zz_4534_ = int_reg_array_50_22_imag;
        _zz_4535_ = int_reg_array_50_22_real;
      end
      6'b010111 : begin
        _zz_4534_ = int_reg_array_50_23_imag;
        _zz_4535_ = int_reg_array_50_23_real;
      end
      6'b011000 : begin
        _zz_4534_ = int_reg_array_50_24_imag;
        _zz_4535_ = int_reg_array_50_24_real;
      end
      6'b011001 : begin
        _zz_4534_ = int_reg_array_50_25_imag;
        _zz_4535_ = int_reg_array_50_25_real;
      end
      6'b011010 : begin
        _zz_4534_ = int_reg_array_50_26_imag;
        _zz_4535_ = int_reg_array_50_26_real;
      end
      6'b011011 : begin
        _zz_4534_ = int_reg_array_50_27_imag;
        _zz_4535_ = int_reg_array_50_27_real;
      end
      6'b011100 : begin
        _zz_4534_ = int_reg_array_50_28_imag;
        _zz_4535_ = int_reg_array_50_28_real;
      end
      6'b011101 : begin
        _zz_4534_ = int_reg_array_50_29_imag;
        _zz_4535_ = int_reg_array_50_29_real;
      end
      6'b011110 : begin
        _zz_4534_ = int_reg_array_50_30_imag;
        _zz_4535_ = int_reg_array_50_30_real;
      end
      6'b011111 : begin
        _zz_4534_ = int_reg_array_50_31_imag;
        _zz_4535_ = int_reg_array_50_31_real;
      end
      6'b100000 : begin
        _zz_4534_ = int_reg_array_50_32_imag;
        _zz_4535_ = int_reg_array_50_32_real;
      end
      6'b100001 : begin
        _zz_4534_ = int_reg_array_50_33_imag;
        _zz_4535_ = int_reg_array_50_33_real;
      end
      6'b100010 : begin
        _zz_4534_ = int_reg_array_50_34_imag;
        _zz_4535_ = int_reg_array_50_34_real;
      end
      6'b100011 : begin
        _zz_4534_ = int_reg_array_50_35_imag;
        _zz_4535_ = int_reg_array_50_35_real;
      end
      6'b100100 : begin
        _zz_4534_ = int_reg_array_50_36_imag;
        _zz_4535_ = int_reg_array_50_36_real;
      end
      6'b100101 : begin
        _zz_4534_ = int_reg_array_50_37_imag;
        _zz_4535_ = int_reg_array_50_37_real;
      end
      6'b100110 : begin
        _zz_4534_ = int_reg_array_50_38_imag;
        _zz_4535_ = int_reg_array_50_38_real;
      end
      6'b100111 : begin
        _zz_4534_ = int_reg_array_50_39_imag;
        _zz_4535_ = int_reg_array_50_39_real;
      end
      6'b101000 : begin
        _zz_4534_ = int_reg_array_50_40_imag;
        _zz_4535_ = int_reg_array_50_40_real;
      end
      6'b101001 : begin
        _zz_4534_ = int_reg_array_50_41_imag;
        _zz_4535_ = int_reg_array_50_41_real;
      end
      6'b101010 : begin
        _zz_4534_ = int_reg_array_50_42_imag;
        _zz_4535_ = int_reg_array_50_42_real;
      end
      6'b101011 : begin
        _zz_4534_ = int_reg_array_50_43_imag;
        _zz_4535_ = int_reg_array_50_43_real;
      end
      6'b101100 : begin
        _zz_4534_ = int_reg_array_50_44_imag;
        _zz_4535_ = int_reg_array_50_44_real;
      end
      6'b101101 : begin
        _zz_4534_ = int_reg_array_50_45_imag;
        _zz_4535_ = int_reg_array_50_45_real;
      end
      6'b101110 : begin
        _zz_4534_ = int_reg_array_50_46_imag;
        _zz_4535_ = int_reg_array_50_46_real;
      end
      6'b101111 : begin
        _zz_4534_ = int_reg_array_50_47_imag;
        _zz_4535_ = int_reg_array_50_47_real;
      end
      6'b110000 : begin
        _zz_4534_ = int_reg_array_50_48_imag;
        _zz_4535_ = int_reg_array_50_48_real;
      end
      6'b110001 : begin
        _zz_4534_ = int_reg_array_50_49_imag;
        _zz_4535_ = int_reg_array_50_49_real;
      end
      6'b110010 : begin
        _zz_4534_ = int_reg_array_50_50_imag;
        _zz_4535_ = int_reg_array_50_50_real;
      end
      6'b110011 : begin
        _zz_4534_ = int_reg_array_50_51_imag;
        _zz_4535_ = int_reg_array_50_51_real;
      end
      6'b110100 : begin
        _zz_4534_ = int_reg_array_50_52_imag;
        _zz_4535_ = int_reg_array_50_52_real;
      end
      6'b110101 : begin
        _zz_4534_ = int_reg_array_50_53_imag;
        _zz_4535_ = int_reg_array_50_53_real;
      end
      6'b110110 : begin
        _zz_4534_ = int_reg_array_50_54_imag;
        _zz_4535_ = int_reg_array_50_54_real;
      end
      6'b110111 : begin
        _zz_4534_ = int_reg_array_50_55_imag;
        _zz_4535_ = int_reg_array_50_55_real;
      end
      6'b111000 : begin
        _zz_4534_ = int_reg_array_50_56_imag;
        _zz_4535_ = int_reg_array_50_56_real;
      end
      6'b111001 : begin
        _zz_4534_ = int_reg_array_50_57_imag;
        _zz_4535_ = int_reg_array_50_57_real;
      end
      6'b111010 : begin
        _zz_4534_ = int_reg_array_50_58_imag;
        _zz_4535_ = int_reg_array_50_58_real;
      end
      6'b111011 : begin
        _zz_4534_ = int_reg_array_50_59_imag;
        _zz_4535_ = int_reg_array_50_59_real;
      end
      6'b111100 : begin
        _zz_4534_ = int_reg_array_50_60_imag;
        _zz_4535_ = int_reg_array_50_60_real;
      end
      6'b111101 : begin
        _zz_4534_ = int_reg_array_50_61_imag;
        _zz_4535_ = int_reg_array_50_61_real;
      end
      6'b111110 : begin
        _zz_4534_ = int_reg_array_50_62_imag;
        _zz_4535_ = int_reg_array_50_62_real;
      end
      default : begin
        _zz_4534_ = int_reg_array_50_63_imag;
        _zz_4535_ = int_reg_array_50_63_real;
      end
    endcase
  end

  always @(*) begin
    case(_zz_3536_)
      6'b000000 : begin
        _zz_4536_ = int_reg_array_51_0_imag;
        _zz_4537_ = int_reg_array_51_0_real;
      end
      6'b000001 : begin
        _zz_4536_ = int_reg_array_51_1_imag;
        _zz_4537_ = int_reg_array_51_1_real;
      end
      6'b000010 : begin
        _zz_4536_ = int_reg_array_51_2_imag;
        _zz_4537_ = int_reg_array_51_2_real;
      end
      6'b000011 : begin
        _zz_4536_ = int_reg_array_51_3_imag;
        _zz_4537_ = int_reg_array_51_3_real;
      end
      6'b000100 : begin
        _zz_4536_ = int_reg_array_51_4_imag;
        _zz_4537_ = int_reg_array_51_4_real;
      end
      6'b000101 : begin
        _zz_4536_ = int_reg_array_51_5_imag;
        _zz_4537_ = int_reg_array_51_5_real;
      end
      6'b000110 : begin
        _zz_4536_ = int_reg_array_51_6_imag;
        _zz_4537_ = int_reg_array_51_6_real;
      end
      6'b000111 : begin
        _zz_4536_ = int_reg_array_51_7_imag;
        _zz_4537_ = int_reg_array_51_7_real;
      end
      6'b001000 : begin
        _zz_4536_ = int_reg_array_51_8_imag;
        _zz_4537_ = int_reg_array_51_8_real;
      end
      6'b001001 : begin
        _zz_4536_ = int_reg_array_51_9_imag;
        _zz_4537_ = int_reg_array_51_9_real;
      end
      6'b001010 : begin
        _zz_4536_ = int_reg_array_51_10_imag;
        _zz_4537_ = int_reg_array_51_10_real;
      end
      6'b001011 : begin
        _zz_4536_ = int_reg_array_51_11_imag;
        _zz_4537_ = int_reg_array_51_11_real;
      end
      6'b001100 : begin
        _zz_4536_ = int_reg_array_51_12_imag;
        _zz_4537_ = int_reg_array_51_12_real;
      end
      6'b001101 : begin
        _zz_4536_ = int_reg_array_51_13_imag;
        _zz_4537_ = int_reg_array_51_13_real;
      end
      6'b001110 : begin
        _zz_4536_ = int_reg_array_51_14_imag;
        _zz_4537_ = int_reg_array_51_14_real;
      end
      6'b001111 : begin
        _zz_4536_ = int_reg_array_51_15_imag;
        _zz_4537_ = int_reg_array_51_15_real;
      end
      6'b010000 : begin
        _zz_4536_ = int_reg_array_51_16_imag;
        _zz_4537_ = int_reg_array_51_16_real;
      end
      6'b010001 : begin
        _zz_4536_ = int_reg_array_51_17_imag;
        _zz_4537_ = int_reg_array_51_17_real;
      end
      6'b010010 : begin
        _zz_4536_ = int_reg_array_51_18_imag;
        _zz_4537_ = int_reg_array_51_18_real;
      end
      6'b010011 : begin
        _zz_4536_ = int_reg_array_51_19_imag;
        _zz_4537_ = int_reg_array_51_19_real;
      end
      6'b010100 : begin
        _zz_4536_ = int_reg_array_51_20_imag;
        _zz_4537_ = int_reg_array_51_20_real;
      end
      6'b010101 : begin
        _zz_4536_ = int_reg_array_51_21_imag;
        _zz_4537_ = int_reg_array_51_21_real;
      end
      6'b010110 : begin
        _zz_4536_ = int_reg_array_51_22_imag;
        _zz_4537_ = int_reg_array_51_22_real;
      end
      6'b010111 : begin
        _zz_4536_ = int_reg_array_51_23_imag;
        _zz_4537_ = int_reg_array_51_23_real;
      end
      6'b011000 : begin
        _zz_4536_ = int_reg_array_51_24_imag;
        _zz_4537_ = int_reg_array_51_24_real;
      end
      6'b011001 : begin
        _zz_4536_ = int_reg_array_51_25_imag;
        _zz_4537_ = int_reg_array_51_25_real;
      end
      6'b011010 : begin
        _zz_4536_ = int_reg_array_51_26_imag;
        _zz_4537_ = int_reg_array_51_26_real;
      end
      6'b011011 : begin
        _zz_4536_ = int_reg_array_51_27_imag;
        _zz_4537_ = int_reg_array_51_27_real;
      end
      6'b011100 : begin
        _zz_4536_ = int_reg_array_51_28_imag;
        _zz_4537_ = int_reg_array_51_28_real;
      end
      6'b011101 : begin
        _zz_4536_ = int_reg_array_51_29_imag;
        _zz_4537_ = int_reg_array_51_29_real;
      end
      6'b011110 : begin
        _zz_4536_ = int_reg_array_51_30_imag;
        _zz_4537_ = int_reg_array_51_30_real;
      end
      6'b011111 : begin
        _zz_4536_ = int_reg_array_51_31_imag;
        _zz_4537_ = int_reg_array_51_31_real;
      end
      6'b100000 : begin
        _zz_4536_ = int_reg_array_51_32_imag;
        _zz_4537_ = int_reg_array_51_32_real;
      end
      6'b100001 : begin
        _zz_4536_ = int_reg_array_51_33_imag;
        _zz_4537_ = int_reg_array_51_33_real;
      end
      6'b100010 : begin
        _zz_4536_ = int_reg_array_51_34_imag;
        _zz_4537_ = int_reg_array_51_34_real;
      end
      6'b100011 : begin
        _zz_4536_ = int_reg_array_51_35_imag;
        _zz_4537_ = int_reg_array_51_35_real;
      end
      6'b100100 : begin
        _zz_4536_ = int_reg_array_51_36_imag;
        _zz_4537_ = int_reg_array_51_36_real;
      end
      6'b100101 : begin
        _zz_4536_ = int_reg_array_51_37_imag;
        _zz_4537_ = int_reg_array_51_37_real;
      end
      6'b100110 : begin
        _zz_4536_ = int_reg_array_51_38_imag;
        _zz_4537_ = int_reg_array_51_38_real;
      end
      6'b100111 : begin
        _zz_4536_ = int_reg_array_51_39_imag;
        _zz_4537_ = int_reg_array_51_39_real;
      end
      6'b101000 : begin
        _zz_4536_ = int_reg_array_51_40_imag;
        _zz_4537_ = int_reg_array_51_40_real;
      end
      6'b101001 : begin
        _zz_4536_ = int_reg_array_51_41_imag;
        _zz_4537_ = int_reg_array_51_41_real;
      end
      6'b101010 : begin
        _zz_4536_ = int_reg_array_51_42_imag;
        _zz_4537_ = int_reg_array_51_42_real;
      end
      6'b101011 : begin
        _zz_4536_ = int_reg_array_51_43_imag;
        _zz_4537_ = int_reg_array_51_43_real;
      end
      6'b101100 : begin
        _zz_4536_ = int_reg_array_51_44_imag;
        _zz_4537_ = int_reg_array_51_44_real;
      end
      6'b101101 : begin
        _zz_4536_ = int_reg_array_51_45_imag;
        _zz_4537_ = int_reg_array_51_45_real;
      end
      6'b101110 : begin
        _zz_4536_ = int_reg_array_51_46_imag;
        _zz_4537_ = int_reg_array_51_46_real;
      end
      6'b101111 : begin
        _zz_4536_ = int_reg_array_51_47_imag;
        _zz_4537_ = int_reg_array_51_47_real;
      end
      6'b110000 : begin
        _zz_4536_ = int_reg_array_51_48_imag;
        _zz_4537_ = int_reg_array_51_48_real;
      end
      6'b110001 : begin
        _zz_4536_ = int_reg_array_51_49_imag;
        _zz_4537_ = int_reg_array_51_49_real;
      end
      6'b110010 : begin
        _zz_4536_ = int_reg_array_51_50_imag;
        _zz_4537_ = int_reg_array_51_50_real;
      end
      6'b110011 : begin
        _zz_4536_ = int_reg_array_51_51_imag;
        _zz_4537_ = int_reg_array_51_51_real;
      end
      6'b110100 : begin
        _zz_4536_ = int_reg_array_51_52_imag;
        _zz_4537_ = int_reg_array_51_52_real;
      end
      6'b110101 : begin
        _zz_4536_ = int_reg_array_51_53_imag;
        _zz_4537_ = int_reg_array_51_53_real;
      end
      6'b110110 : begin
        _zz_4536_ = int_reg_array_51_54_imag;
        _zz_4537_ = int_reg_array_51_54_real;
      end
      6'b110111 : begin
        _zz_4536_ = int_reg_array_51_55_imag;
        _zz_4537_ = int_reg_array_51_55_real;
      end
      6'b111000 : begin
        _zz_4536_ = int_reg_array_51_56_imag;
        _zz_4537_ = int_reg_array_51_56_real;
      end
      6'b111001 : begin
        _zz_4536_ = int_reg_array_51_57_imag;
        _zz_4537_ = int_reg_array_51_57_real;
      end
      6'b111010 : begin
        _zz_4536_ = int_reg_array_51_58_imag;
        _zz_4537_ = int_reg_array_51_58_real;
      end
      6'b111011 : begin
        _zz_4536_ = int_reg_array_51_59_imag;
        _zz_4537_ = int_reg_array_51_59_real;
      end
      6'b111100 : begin
        _zz_4536_ = int_reg_array_51_60_imag;
        _zz_4537_ = int_reg_array_51_60_real;
      end
      6'b111101 : begin
        _zz_4536_ = int_reg_array_51_61_imag;
        _zz_4537_ = int_reg_array_51_61_real;
      end
      6'b111110 : begin
        _zz_4536_ = int_reg_array_51_62_imag;
        _zz_4537_ = int_reg_array_51_62_real;
      end
      default : begin
        _zz_4536_ = int_reg_array_51_63_imag;
        _zz_4537_ = int_reg_array_51_63_real;
      end
    endcase
  end

  always @(*) begin
    case(_zz_3605_)
      6'b000000 : begin
        _zz_4538_ = int_reg_array_52_0_imag;
        _zz_4539_ = int_reg_array_52_0_real;
      end
      6'b000001 : begin
        _zz_4538_ = int_reg_array_52_1_imag;
        _zz_4539_ = int_reg_array_52_1_real;
      end
      6'b000010 : begin
        _zz_4538_ = int_reg_array_52_2_imag;
        _zz_4539_ = int_reg_array_52_2_real;
      end
      6'b000011 : begin
        _zz_4538_ = int_reg_array_52_3_imag;
        _zz_4539_ = int_reg_array_52_3_real;
      end
      6'b000100 : begin
        _zz_4538_ = int_reg_array_52_4_imag;
        _zz_4539_ = int_reg_array_52_4_real;
      end
      6'b000101 : begin
        _zz_4538_ = int_reg_array_52_5_imag;
        _zz_4539_ = int_reg_array_52_5_real;
      end
      6'b000110 : begin
        _zz_4538_ = int_reg_array_52_6_imag;
        _zz_4539_ = int_reg_array_52_6_real;
      end
      6'b000111 : begin
        _zz_4538_ = int_reg_array_52_7_imag;
        _zz_4539_ = int_reg_array_52_7_real;
      end
      6'b001000 : begin
        _zz_4538_ = int_reg_array_52_8_imag;
        _zz_4539_ = int_reg_array_52_8_real;
      end
      6'b001001 : begin
        _zz_4538_ = int_reg_array_52_9_imag;
        _zz_4539_ = int_reg_array_52_9_real;
      end
      6'b001010 : begin
        _zz_4538_ = int_reg_array_52_10_imag;
        _zz_4539_ = int_reg_array_52_10_real;
      end
      6'b001011 : begin
        _zz_4538_ = int_reg_array_52_11_imag;
        _zz_4539_ = int_reg_array_52_11_real;
      end
      6'b001100 : begin
        _zz_4538_ = int_reg_array_52_12_imag;
        _zz_4539_ = int_reg_array_52_12_real;
      end
      6'b001101 : begin
        _zz_4538_ = int_reg_array_52_13_imag;
        _zz_4539_ = int_reg_array_52_13_real;
      end
      6'b001110 : begin
        _zz_4538_ = int_reg_array_52_14_imag;
        _zz_4539_ = int_reg_array_52_14_real;
      end
      6'b001111 : begin
        _zz_4538_ = int_reg_array_52_15_imag;
        _zz_4539_ = int_reg_array_52_15_real;
      end
      6'b010000 : begin
        _zz_4538_ = int_reg_array_52_16_imag;
        _zz_4539_ = int_reg_array_52_16_real;
      end
      6'b010001 : begin
        _zz_4538_ = int_reg_array_52_17_imag;
        _zz_4539_ = int_reg_array_52_17_real;
      end
      6'b010010 : begin
        _zz_4538_ = int_reg_array_52_18_imag;
        _zz_4539_ = int_reg_array_52_18_real;
      end
      6'b010011 : begin
        _zz_4538_ = int_reg_array_52_19_imag;
        _zz_4539_ = int_reg_array_52_19_real;
      end
      6'b010100 : begin
        _zz_4538_ = int_reg_array_52_20_imag;
        _zz_4539_ = int_reg_array_52_20_real;
      end
      6'b010101 : begin
        _zz_4538_ = int_reg_array_52_21_imag;
        _zz_4539_ = int_reg_array_52_21_real;
      end
      6'b010110 : begin
        _zz_4538_ = int_reg_array_52_22_imag;
        _zz_4539_ = int_reg_array_52_22_real;
      end
      6'b010111 : begin
        _zz_4538_ = int_reg_array_52_23_imag;
        _zz_4539_ = int_reg_array_52_23_real;
      end
      6'b011000 : begin
        _zz_4538_ = int_reg_array_52_24_imag;
        _zz_4539_ = int_reg_array_52_24_real;
      end
      6'b011001 : begin
        _zz_4538_ = int_reg_array_52_25_imag;
        _zz_4539_ = int_reg_array_52_25_real;
      end
      6'b011010 : begin
        _zz_4538_ = int_reg_array_52_26_imag;
        _zz_4539_ = int_reg_array_52_26_real;
      end
      6'b011011 : begin
        _zz_4538_ = int_reg_array_52_27_imag;
        _zz_4539_ = int_reg_array_52_27_real;
      end
      6'b011100 : begin
        _zz_4538_ = int_reg_array_52_28_imag;
        _zz_4539_ = int_reg_array_52_28_real;
      end
      6'b011101 : begin
        _zz_4538_ = int_reg_array_52_29_imag;
        _zz_4539_ = int_reg_array_52_29_real;
      end
      6'b011110 : begin
        _zz_4538_ = int_reg_array_52_30_imag;
        _zz_4539_ = int_reg_array_52_30_real;
      end
      6'b011111 : begin
        _zz_4538_ = int_reg_array_52_31_imag;
        _zz_4539_ = int_reg_array_52_31_real;
      end
      6'b100000 : begin
        _zz_4538_ = int_reg_array_52_32_imag;
        _zz_4539_ = int_reg_array_52_32_real;
      end
      6'b100001 : begin
        _zz_4538_ = int_reg_array_52_33_imag;
        _zz_4539_ = int_reg_array_52_33_real;
      end
      6'b100010 : begin
        _zz_4538_ = int_reg_array_52_34_imag;
        _zz_4539_ = int_reg_array_52_34_real;
      end
      6'b100011 : begin
        _zz_4538_ = int_reg_array_52_35_imag;
        _zz_4539_ = int_reg_array_52_35_real;
      end
      6'b100100 : begin
        _zz_4538_ = int_reg_array_52_36_imag;
        _zz_4539_ = int_reg_array_52_36_real;
      end
      6'b100101 : begin
        _zz_4538_ = int_reg_array_52_37_imag;
        _zz_4539_ = int_reg_array_52_37_real;
      end
      6'b100110 : begin
        _zz_4538_ = int_reg_array_52_38_imag;
        _zz_4539_ = int_reg_array_52_38_real;
      end
      6'b100111 : begin
        _zz_4538_ = int_reg_array_52_39_imag;
        _zz_4539_ = int_reg_array_52_39_real;
      end
      6'b101000 : begin
        _zz_4538_ = int_reg_array_52_40_imag;
        _zz_4539_ = int_reg_array_52_40_real;
      end
      6'b101001 : begin
        _zz_4538_ = int_reg_array_52_41_imag;
        _zz_4539_ = int_reg_array_52_41_real;
      end
      6'b101010 : begin
        _zz_4538_ = int_reg_array_52_42_imag;
        _zz_4539_ = int_reg_array_52_42_real;
      end
      6'b101011 : begin
        _zz_4538_ = int_reg_array_52_43_imag;
        _zz_4539_ = int_reg_array_52_43_real;
      end
      6'b101100 : begin
        _zz_4538_ = int_reg_array_52_44_imag;
        _zz_4539_ = int_reg_array_52_44_real;
      end
      6'b101101 : begin
        _zz_4538_ = int_reg_array_52_45_imag;
        _zz_4539_ = int_reg_array_52_45_real;
      end
      6'b101110 : begin
        _zz_4538_ = int_reg_array_52_46_imag;
        _zz_4539_ = int_reg_array_52_46_real;
      end
      6'b101111 : begin
        _zz_4538_ = int_reg_array_52_47_imag;
        _zz_4539_ = int_reg_array_52_47_real;
      end
      6'b110000 : begin
        _zz_4538_ = int_reg_array_52_48_imag;
        _zz_4539_ = int_reg_array_52_48_real;
      end
      6'b110001 : begin
        _zz_4538_ = int_reg_array_52_49_imag;
        _zz_4539_ = int_reg_array_52_49_real;
      end
      6'b110010 : begin
        _zz_4538_ = int_reg_array_52_50_imag;
        _zz_4539_ = int_reg_array_52_50_real;
      end
      6'b110011 : begin
        _zz_4538_ = int_reg_array_52_51_imag;
        _zz_4539_ = int_reg_array_52_51_real;
      end
      6'b110100 : begin
        _zz_4538_ = int_reg_array_52_52_imag;
        _zz_4539_ = int_reg_array_52_52_real;
      end
      6'b110101 : begin
        _zz_4538_ = int_reg_array_52_53_imag;
        _zz_4539_ = int_reg_array_52_53_real;
      end
      6'b110110 : begin
        _zz_4538_ = int_reg_array_52_54_imag;
        _zz_4539_ = int_reg_array_52_54_real;
      end
      6'b110111 : begin
        _zz_4538_ = int_reg_array_52_55_imag;
        _zz_4539_ = int_reg_array_52_55_real;
      end
      6'b111000 : begin
        _zz_4538_ = int_reg_array_52_56_imag;
        _zz_4539_ = int_reg_array_52_56_real;
      end
      6'b111001 : begin
        _zz_4538_ = int_reg_array_52_57_imag;
        _zz_4539_ = int_reg_array_52_57_real;
      end
      6'b111010 : begin
        _zz_4538_ = int_reg_array_52_58_imag;
        _zz_4539_ = int_reg_array_52_58_real;
      end
      6'b111011 : begin
        _zz_4538_ = int_reg_array_52_59_imag;
        _zz_4539_ = int_reg_array_52_59_real;
      end
      6'b111100 : begin
        _zz_4538_ = int_reg_array_52_60_imag;
        _zz_4539_ = int_reg_array_52_60_real;
      end
      6'b111101 : begin
        _zz_4538_ = int_reg_array_52_61_imag;
        _zz_4539_ = int_reg_array_52_61_real;
      end
      6'b111110 : begin
        _zz_4538_ = int_reg_array_52_62_imag;
        _zz_4539_ = int_reg_array_52_62_real;
      end
      default : begin
        _zz_4538_ = int_reg_array_52_63_imag;
        _zz_4539_ = int_reg_array_52_63_real;
      end
    endcase
  end

  always @(*) begin
    case(_zz_3674_)
      6'b000000 : begin
        _zz_4540_ = int_reg_array_53_0_imag;
        _zz_4541_ = int_reg_array_53_0_real;
      end
      6'b000001 : begin
        _zz_4540_ = int_reg_array_53_1_imag;
        _zz_4541_ = int_reg_array_53_1_real;
      end
      6'b000010 : begin
        _zz_4540_ = int_reg_array_53_2_imag;
        _zz_4541_ = int_reg_array_53_2_real;
      end
      6'b000011 : begin
        _zz_4540_ = int_reg_array_53_3_imag;
        _zz_4541_ = int_reg_array_53_3_real;
      end
      6'b000100 : begin
        _zz_4540_ = int_reg_array_53_4_imag;
        _zz_4541_ = int_reg_array_53_4_real;
      end
      6'b000101 : begin
        _zz_4540_ = int_reg_array_53_5_imag;
        _zz_4541_ = int_reg_array_53_5_real;
      end
      6'b000110 : begin
        _zz_4540_ = int_reg_array_53_6_imag;
        _zz_4541_ = int_reg_array_53_6_real;
      end
      6'b000111 : begin
        _zz_4540_ = int_reg_array_53_7_imag;
        _zz_4541_ = int_reg_array_53_7_real;
      end
      6'b001000 : begin
        _zz_4540_ = int_reg_array_53_8_imag;
        _zz_4541_ = int_reg_array_53_8_real;
      end
      6'b001001 : begin
        _zz_4540_ = int_reg_array_53_9_imag;
        _zz_4541_ = int_reg_array_53_9_real;
      end
      6'b001010 : begin
        _zz_4540_ = int_reg_array_53_10_imag;
        _zz_4541_ = int_reg_array_53_10_real;
      end
      6'b001011 : begin
        _zz_4540_ = int_reg_array_53_11_imag;
        _zz_4541_ = int_reg_array_53_11_real;
      end
      6'b001100 : begin
        _zz_4540_ = int_reg_array_53_12_imag;
        _zz_4541_ = int_reg_array_53_12_real;
      end
      6'b001101 : begin
        _zz_4540_ = int_reg_array_53_13_imag;
        _zz_4541_ = int_reg_array_53_13_real;
      end
      6'b001110 : begin
        _zz_4540_ = int_reg_array_53_14_imag;
        _zz_4541_ = int_reg_array_53_14_real;
      end
      6'b001111 : begin
        _zz_4540_ = int_reg_array_53_15_imag;
        _zz_4541_ = int_reg_array_53_15_real;
      end
      6'b010000 : begin
        _zz_4540_ = int_reg_array_53_16_imag;
        _zz_4541_ = int_reg_array_53_16_real;
      end
      6'b010001 : begin
        _zz_4540_ = int_reg_array_53_17_imag;
        _zz_4541_ = int_reg_array_53_17_real;
      end
      6'b010010 : begin
        _zz_4540_ = int_reg_array_53_18_imag;
        _zz_4541_ = int_reg_array_53_18_real;
      end
      6'b010011 : begin
        _zz_4540_ = int_reg_array_53_19_imag;
        _zz_4541_ = int_reg_array_53_19_real;
      end
      6'b010100 : begin
        _zz_4540_ = int_reg_array_53_20_imag;
        _zz_4541_ = int_reg_array_53_20_real;
      end
      6'b010101 : begin
        _zz_4540_ = int_reg_array_53_21_imag;
        _zz_4541_ = int_reg_array_53_21_real;
      end
      6'b010110 : begin
        _zz_4540_ = int_reg_array_53_22_imag;
        _zz_4541_ = int_reg_array_53_22_real;
      end
      6'b010111 : begin
        _zz_4540_ = int_reg_array_53_23_imag;
        _zz_4541_ = int_reg_array_53_23_real;
      end
      6'b011000 : begin
        _zz_4540_ = int_reg_array_53_24_imag;
        _zz_4541_ = int_reg_array_53_24_real;
      end
      6'b011001 : begin
        _zz_4540_ = int_reg_array_53_25_imag;
        _zz_4541_ = int_reg_array_53_25_real;
      end
      6'b011010 : begin
        _zz_4540_ = int_reg_array_53_26_imag;
        _zz_4541_ = int_reg_array_53_26_real;
      end
      6'b011011 : begin
        _zz_4540_ = int_reg_array_53_27_imag;
        _zz_4541_ = int_reg_array_53_27_real;
      end
      6'b011100 : begin
        _zz_4540_ = int_reg_array_53_28_imag;
        _zz_4541_ = int_reg_array_53_28_real;
      end
      6'b011101 : begin
        _zz_4540_ = int_reg_array_53_29_imag;
        _zz_4541_ = int_reg_array_53_29_real;
      end
      6'b011110 : begin
        _zz_4540_ = int_reg_array_53_30_imag;
        _zz_4541_ = int_reg_array_53_30_real;
      end
      6'b011111 : begin
        _zz_4540_ = int_reg_array_53_31_imag;
        _zz_4541_ = int_reg_array_53_31_real;
      end
      6'b100000 : begin
        _zz_4540_ = int_reg_array_53_32_imag;
        _zz_4541_ = int_reg_array_53_32_real;
      end
      6'b100001 : begin
        _zz_4540_ = int_reg_array_53_33_imag;
        _zz_4541_ = int_reg_array_53_33_real;
      end
      6'b100010 : begin
        _zz_4540_ = int_reg_array_53_34_imag;
        _zz_4541_ = int_reg_array_53_34_real;
      end
      6'b100011 : begin
        _zz_4540_ = int_reg_array_53_35_imag;
        _zz_4541_ = int_reg_array_53_35_real;
      end
      6'b100100 : begin
        _zz_4540_ = int_reg_array_53_36_imag;
        _zz_4541_ = int_reg_array_53_36_real;
      end
      6'b100101 : begin
        _zz_4540_ = int_reg_array_53_37_imag;
        _zz_4541_ = int_reg_array_53_37_real;
      end
      6'b100110 : begin
        _zz_4540_ = int_reg_array_53_38_imag;
        _zz_4541_ = int_reg_array_53_38_real;
      end
      6'b100111 : begin
        _zz_4540_ = int_reg_array_53_39_imag;
        _zz_4541_ = int_reg_array_53_39_real;
      end
      6'b101000 : begin
        _zz_4540_ = int_reg_array_53_40_imag;
        _zz_4541_ = int_reg_array_53_40_real;
      end
      6'b101001 : begin
        _zz_4540_ = int_reg_array_53_41_imag;
        _zz_4541_ = int_reg_array_53_41_real;
      end
      6'b101010 : begin
        _zz_4540_ = int_reg_array_53_42_imag;
        _zz_4541_ = int_reg_array_53_42_real;
      end
      6'b101011 : begin
        _zz_4540_ = int_reg_array_53_43_imag;
        _zz_4541_ = int_reg_array_53_43_real;
      end
      6'b101100 : begin
        _zz_4540_ = int_reg_array_53_44_imag;
        _zz_4541_ = int_reg_array_53_44_real;
      end
      6'b101101 : begin
        _zz_4540_ = int_reg_array_53_45_imag;
        _zz_4541_ = int_reg_array_53_45_real;
      end
      6'b101110 : begin
        _zz_4540_ = int_reg_array_53_46_imag;
        _zz_4541_ = int_reg_array_53_46_real;
      end
      6'b101111 : begin
        _zz_4540_ = int_reg_array_53_47_imag;
        _zz_4541_ = int_reg_array_53_47_real;
      end
      6'b110000 : begin
        _zz_4540_ = int_reg_array_53_48_imag;
        _zz_4541_ = int_reg_array_53_48_real;
      end
      6'b110001 : begin
        _zz_4540_ = int_reg_array_53_49_imag;
        _zz_4541_ = int_reg_array_53_49_real;
      end
      6'b110010 : begin
        _zz_4540_ = int_reg_array_53_50_imag;
        _zz_4541_ = int_reg_array_53_50_real;
      end
      6'b110011 : begin
        _zz_4540_ = int_reg_array_53_51_imag;
        _zz_4541_ = int_reg_array_53_51_real;
      end
      6'b110100 : begin
        _zz_4540_ = int_reg_array_53_52_imag;
        _zz_4541_ = int_reg_array_53_52_real;
      end
      6'b110101 : begin
        _zz_4540_ = int_reg_array_53_53_imag;
        _zz_4541_ = int_reg_array_53_53_real;
      end
      6'b110110 : begin
        _zz_4540_ = int_reg_array_53_54_imag;
        _zz_4541_ = int_reg_array_53_54_real;
      end
      6'b110111 : begin
        _zz_4540_ = int_reg_array_53_55_imag;
        _zz_4541_ = int_reg_array_53_55_real;
      end
      6'b111000 : begin
        _zz_4540_ = int_reg_array_53_56_imag;
        _zz_4541_ = int_reg_array_53_56_real;
      end
      6'b111001 : begin
        _zz_4540_ = int_reg_array_53_57_imag;
        _zz_4541_ = int_reg_array_53_57_real;
      end
      6'b111010 : begin
        _zz_4540_ = int_reg_array_53_58_imag;
        _zz_4541_ = int_reg_array_53_58_real;
      end
      6'b111011 : begin
        _zz_4540_ = int_reg_array_53_59_imag;
        _zz_4541_ = int_reg_array_53_59_real;
      end
      6'b111100 : begin
        _zz_4540_ = int_reg_array_53_60_imag;
        _zz_4541_ = int_reg_array_53_60_real;
      end
      6'b111101 : begin
        _zz_4540_ = int_reg_array_53_61_imag;
        _zz_4541_ = int_reg_array_53_61_real;
      end
      6'b111110 : begin
        _zz_4540_ = int_reg_array_53_62_imag;
        _zz_4541_ = int_reg_array_53_62_real;
      end
      default : begin
        _zz_4540_ = int_reg_array_53_63_imag;
        _zz_4541_ = int_reg_array_53_63_real;
      end
    endcase
  end

  always @(*) begin
    case(_zz_3743_)
      6'b000000 : begin
        _zz_4542_ = int_reg_array_54_0_imag;
        _zz_4543_ = int_reg_array_54_0_real;
      end
      6'b000001 : begin
        _zz_4542_ = int_reg_array_54_1_imag;
        _zz_4543_ = int_reg_array_54_1_real;
      end
      6'b000010 : begin
        _zz_4542_ = int_reg_array_54_2_imag;
        _zz_4543_ = int_reg_array_54_2_real;
      end
      6'b000011 : begin
        _zz_4542_ = int_reg_array_54_3_imag;
        _zz_4543_ = int_reg_array_54_3_real;
      end
      6'b000100 : begin
        _zz_4542_ = int_reg_array_54_4_imag;
        _zz_4543_ = int_reg_array_54_4_real;
      end
      6'b000101 : begin
        _zz_4542_ = int_reg_array_54_5_imag;
        _zz_4543_ = int_reg_array_54_5_real;
      end
      6'b000110 : begin
        _zz_4542_ = int_reg_array_54_6_imag;
        _zz_4543_ = int_reg_array_54_6_real;
      end
      6'b000111 : begin
        _zz_4542_ = int_reg_array_54_7_imag;
        _zz_4543_ = int_reg_array_54_7_real;
      end
      6'b001000 : begin
        _zz_4542_ = int_reg_array_54_8_imag;
        _zz_4543_ = int_reg_array_54_8_real;
      end
      6'b001001 : begin
        _zz_4542_ = int_reg_array_54_9_imag;
        _zz_4543_ = int_reg_array_54_9_real;
      end
      6'b001010 : begin
        _zz_4542_ = int_reg_array_54_10_imag;
        _zz_4543_ = int_reg_array_54_10_real;
      end
      6'b001011 : begin
        _zz_4542_ = int_reg_array_54_11_imag;
        _zz_4543_ = int_reg_array_54_11_real;
      end
      6'b001100 : begin
        _zz_4542_ = int_reg_array_54_12_imag;
        _zz_4543_ = int_reg_array_54_12_real;
      end
      6'b001101 : begin
        _zz_4542_ = int_reg_array_54_13_imag;
        _zz_4543_ = int_reg_array_54_13_real;
      end
      6'b001110 : begin
        _zz_4542_ = int_reg_array_54_14_imag;
        _zz_4543_ = int_reg_array_54_14_real;
      end
      6'b001111 : begin
        _zz_4542_ = int_reg_array_54_15_imag;
        _zz_4543_ = int_reg_array_54_15_real;
      end
      6'b010000 : begin
        _zz_4542_ = int_reg_array_54_16_imag;
        _zz_4543_ = int_reg_array_54_16_real;
      end
      6'b010001 : begin
        _zz_4542_ = int_reg_array_54_17_imag;
        _zz_4543_ = int_reg_array_54_17_real;
      end
      6'b010010 : begin
        _zz_4542_ = int_reg_array_54_18_imag;
        _zz_4543_ = int_reg_array_54_18_real;
      end
      6'b010011 : begin
        _zz_4542_ = int_reg_array_54_19_imag;
        _zz_4543_ = int_reg_array_54_19_real;
      end
      6'b010100 : begin
        _zz_4542_ = int_reg_array_54_20_imag;
        _zz_4543_ = int_reg_array_54_20_real;
      end
      6'b010101 : begin
        _zz_4542_ = int_reg_array_54_21_imag;
        _zz_4543_ = int_reg_array_54_21_real;
      end
      6'b010110 : begin
        _zz_4542_ = int_reg_array_54_22_imag;
        _zz_4543_ = int_reg_array_54_22_real;
      end
      6'b010111 : begin
        _zz_4542_ = int_reg_array_54_23_imag;
        _zz_4543_ = int_reg_array_54_23_real;
      end
      6'b011000 : begin
        _zz_4542_ = int_reg_array_54_24_imag;
        _zz_4543_ = int_reg_array_54_24_real;
      end
      6'b011001 : begin
        _zz_4542_ = int_reg_array_54_25_imag;
        _zz_4543_ = int_reg_array_54_25_real;
      end
      6'b011010 : begin
        _zz_4542_ = int_reg_array_54_26_imag;
        _zz_4543_ = int_reg_array_54_26_real;
      end
      6'b011011 : begin
        _zz_4542_ = int_reg_array_54_27_imag;
        _zz_4543_ = int_reg_array_54_27_real;
      end
      6'b011100 : begin
        _zz_4542_ = int_reg_array_54_28_imag;
        _zz_4543_ = int_reg_array_54_28_real;
      end
      6'b011101 : begin
        _zz_4542_ = int_reg_array_54_29_imag;
        _zz_4543_ = int_reg_array_54_29_real;
      end
      6'b011110 : begin
        _zz_4542_ = int_reg_array_54_30_imag;
        _zz_4543_ = int_reg_array_54_30_real;
      end
      6'b011111 : begin
        _zz_4542_ = int_reg_array_54_31_imag;
        _zz_4543_ = int_reg_array_54_31_real;
      end
      6'b100000 : begin
        _zz_4542_ = int_reg_array_54_32_imag;
        _zz_4543_ = int_reg_array_54_32_real;
      end
      6'b100001 : begin
        _zz_4542_ = int_reg_array_54_33_imag;
        _zz_4543_ = int_reg_array_54_33_real;
      end
      6'b100010 : begin
        _zz_4542_ = int_reg_array_54_34_imag;
        _zz_4543_ = int_reg_array_54_34_real;
      end
      6'b100011 : begin
        _zz_4542_ = int_reg_array_54_35_imag;
        _zz_4543_ = int_reg_array_54_35_real;
      end
      6'b100100 : begin
        _zz_4542_ = int_reg_array_54_36_imag;
        _zz_4543_ = int_reg_array_54_36_real;
      end
      6'b100101 : begin
        _zz_4542_ = int_reg_array_54_37_imag;
        _zz_4543_ = int_reg_array_54_37_real;
      end
      6'b100110 : begin
        _zz_4542_ = int_reg_array_54_38_imag;
        _zz_4543_ = int_reg_array_54_38_real;
      end
      6'b100111 : begin
        _zz_4542_ = int_reg_array_54_39_imag;
        _zz_4543_ = int_reg_array_54_39_real;
      end
      6'b101000 : begin
        _zz_4542_ = int_reg_array_54_40_imag;
        _zz_4543_ = int_reg_array_54_40_real;
      end
      6'b101001 : begin
        _zz_4542_ = int_reg_array_54_41_imag;
        _zz_4543_ = int_reg_array_54_41_real;
      end
      6'b101010 : begin
        _zz_4542_ = int_reg_array_54_42_imag;
        _zz_4543_ = int_reg_array_54_42_real;
      end
      6'b101011 : begin
        _zz_4542_ = int_reg_array_54_43_imag;
        _zz_4543_ = int_reg_array_54_43_real;
      end
      6'b101100 : begin
        _zz_4542_ = int_reg_array_54_44_imag;
        _zz_4543_ = int_reg_array_54_44_real;
      end
      6'b101101 : begin
        _zz_4542_ = int_reg_array_54_45_imag;
        _zz_4543_ = int_reg_array_54_45_real;
      end
      6'b101110 : begin
        _zz_4542_ = int_reg_array_54_46_imag;
        _zz_4543_ = int_reg_array_54_46_real;
      end
      6'b101111 : begin
        _zz_4542_ = int_reg_array_54_47_imag;
        _zz_4543_ = int_reg_array_54_47_real;
      end
      6'b110000 : begin
        _zz_4542_ = int_reg_array_54_48_imag;
        _zz_4543_ = int_reg_array_54_48_real;
      end
      6'b110001 : begin
        _zz_4542_ = int_reg_array_54_49_imag;
        _zz_4543_ = int_reg_array_54_49_real;
      end
      6'b110010 : begin
        _zz_4542_ = int_reg_array_54_50_imag;
        _zz_4543_ = int_reg_array_54_50_real;
      end
      6'b110011 : begin
        _zz_4542_ = int_reg_array_54_51_imag;
        _zz_4543_ = int_reg_array_54_51_real;
      end
      6'b110100 : begin
        _zz_4542_ = int_reg_array_54_52_imag;
        _zz_4543_ = int_reg_array_54_52_real;
      end
      6'b110101 : begin
        _zz_4542_ = int_reg_array_54_53_imag;
        _zz_4543_ = int_reg_array_54_53_real;
      end
      6'b110110 : begin
        _zz_4542_ = int_reg_array_54_54_imag;
        _zz_4543_ = int_reg_array_54_54_real;
      end
      6'b110111 : begin
        _zz_4542_ = int_reg_array_54_55_imag;
        _zz_4543_ = int_reg_array_54_55_real;
      end
      6'b111000 : begin
        _zz_4542_ = int_reg_array_54_56_imag;
        _zz_4543_ = int_reg_array_54_56_real;
      end
      6'b111001 : begin
        _zz_4542_ = int_reg_array_54_57_imag;
        _zz_4543_ = int_reg_array_54_57_real;
      end
      6'b111010 : begin
        _zz_4542_ = int_reg_array_54_58_imag;
        _zz_4543_ = int_reg_array_54_58_real;
      end
      6'b111011 : begin
        _zz_4542_ = int_reg_array_54_59_imag;
        _zz_4543_ = int_reg_array_54_59_real;
      end
      6'b111100 : begin
        _zz_4542_ = int_reg_array_54_60_imag;
        _zz_4543_ = int_reg_array_54_60_real;
      end
      6'b111101 : begin
        _zz_4542_ = int_reg_array_54_61_imag;
        _zz_4543_ = int_reg_array_54_61_real;
      end
      6'b111110 : begin
        _zz_4542_ = int_reg_array_54_62_imag;
        _zz_4543_ = int_reg_array_54_62_real;
      end
      default : begin
        _zz_4542_ = int_reg_array_54_63_imag;
        _zz_4543_ = int_reg_array_54_63_real;
      end
    endcase
  end

  always @(*) begin
    case(_zz_3812_)
      6'b000000 : begin
        _zz_4544_ = int_reg_array_55_0_imag;
        _zz_4545_ = int_reg_array_55_0_real;
      end
      6'b000001 : begin
        _zz_4544_ = int_reg_array_55_1_imag;
        _zz_4545_ = int_reg_array_55_1_real;
      end
      6'b000010 : begin
        _zz_4544_ = int_reg_array_55_2_imag;
        _zz_4545_ = int_reg_array_55_2_real;
      end
      6'b000011 : begin
        _zz_4544_ = int_reg_array_55_3_imag;
        _zz_4545_ = int_reg_array_55_3_real;
      end
      6'b000100 : begin
        _zz_4544_ = int_reg_array_55_4_imag;
        _zz_4545_ = int_reg_array_55_4_real;
      end
      6'b000101 : begin
        _zz_4544_ = int_reg_array_55_5_imag;
        _zz_4545_ = int_reg_array_55_5_real;
      end
      6'b000110 : begin
        _zz_4544_ = int_reg_array_55_6_imag;
        _zz_4545_ = int_reg_array_55_6_real;
      end
      6'b000111 : begin
        _zz_4544_ = int_reg_array_55_7_imag;
        _zz_4545_ = int_reg_array_55_7_real;
      end
      6'b001000 : begin
        _zz_4544_ = int_reg_array_55_8_imag;
        _zz_4545_ = int_reg_array_55_8_real;
      end
      6'b001001 : begin
        _zz_4544_ = int_reg_array_55_9_imag;
        _zz_4545_ = int_reg_array_55_9_real;
      end
      6'b001010 : begin
        _zz_4544_ = int_reg_array_55_10_imag;
        _zz_4545_ = int_reg_array_55_10_real;
      end
      6'b001011 : begin
        _zz_4544_ = int_reg_array_55_11_imag;
        _zz_4545_ = int_reg_array_55_11_real;
      end
      6'b001100 : begin
        _zz_4544_ = int_reg_array_55_12_imag;
        _zz_4545_ = int_reg_array_55_12_real;
      end
      6'b001101 : begin
        _zz_4544_ = int_reg_array_55_13_imag;
        _zz_4545_ = int_reg_array_55_13_real;
      end
      6'b001110 : begin
        _zz_4544_ = int_reg_array_55_14_imag;
        _zz_4545_ = int_reg_array_55_14_real;
      end
      6'b001111 : begin
        _zz_4544_ = int_reg_array_55_15_imag;
        _zz_4545_ = int_reg_array_55_15_real;
      end
      6'b010000 : begin
        _zz_4544_ = int_reg_array_55_16_imag;
        _zz_4545_ = int_reg_array_55_16_real;
      end
      6'b010001 : begin
        _zz_4544_ = int_reg_array_55_17_imag;
        _zz_4545_ = int_reg_array_55_17_real;
      end
      6'b010010 : begin
        _zz_4544_ = int_reg_array_55_18_imag;
        _zz_4545_ = int_reg_array_55_18_real;
      end
      6'b010011 : begin
        _zz_4544_ = int_reg_array_55_19_imag;
        _zz_4545_ = int_reg_array_55_19_real;
      end
      6'b010100 : begin
        _zz_4544_ = int_reg_array_55_20_imag;
        _zz_4545_ = int_reg_array_55_20_real;
      end
      6'b010101 : begin
        _zz_4544_ = int_reg_array_55_21_imag;
        _zz_4545_ = int_reg_array_55_21_real;
      end
      6'b010110 : begin
        _zz_4544_ = int_reg_array_55_22_imag;
        _zz_4545_ = int_reg_array_55_22_real;
      end
      6'b010111 : begin
        _zz_4544_ = int_reg_array_55_23_imag;
        _zz_4545_ = int_reg_array_55_23_real;
      end
      6'b011000 : begin
        _zz_4544_ = int_reg_array_55_24_imag;
        _zz_4545_ = int_reg_array_55_24_real;
      end
      6'b011001 : begin
        _zz_4544_ = int_reg_array_55_25_imag;
        _zz_4545_ = int_reg_array_55_25_real;
      end
      6'b011010 : begin
        _zz_4544_ = int_reg_array_55_26_imag;
        _zz_4545_ = int_reg_array_55_26_real;
      end
      6'b011011 : begin
        _zz_4544_ = int_reg_array_55_27_imag;
        _zz_4545_ = int_reg_array_55_27_real;
      end
      6'b011100 : begin
        _zz_4544_ = int_reg_array_55_28_imag;
        _zz_4545_ = int_reg_array_55_28_real;
      end
      6'b011101 : begin
        _zz_4544_ = int_reg_array_55_29_imag;
        _zz_4545_ = int_reg_array_55_29_real;
      end
      6'b011110 : begin
        _zz_4544_ = int_reg_array_55_30_imag;
        _zz_4545_ = int_reg_array_55_30_real;
      end
      6'b011111 : begin
        _zz_4544_ = int_reg_array_55_31_imag;
        _zz_4545_ = int_reg_array_55_31_real;
      end
      6'b100000 : begin
        _zz_4544_ = int_reg_array_55_32_imag;
        _zz_4545_ = int_reg_array_55_32_real;
      end
      6'b100001 : begin
        _zz_4544_ = int_reg_array_55_33_imag;
        _zz_4545_ = int_reg_array_55_33_real;
      end
      6'b100010 : begin
        _zz_4544_ = int_reg_array_55_34_imag;
        _zz_4545_ = int_reg_array_55_34_real;
      end
      6'b100011 : begin
        _zz_4544_ = int_reg_array_55_35_imag;
        _zz_4545_ = int_reg_array_55_35_real;
      end
      6'b100100 : begin
        _zz_4544_ = int_reg_array_55_36_imag;
        _zz_4545_ = int_reg_array_55_36_real;
      end
      6'b100101 : begin
        _zz_4544_ = int_reg_array_55_37_imag;
        _zz_4545_ = int_reg_array_55_37_real;
      end
      6'b100110 : begin
        _zz_4544_ = int_reg_array_55_38_imag;
        _zz_4545_ = int_reg_array_55_38_real;
      end
      6'b100111 : begin
        _zz_4544_ = int_reg_array_55_39_imag;
        _zz_4545_ = int_reg_array_55_39_real;
      end
      6'b101000 : begin
        _zz_4544_ = int_reg_array_55_40_imag;
        _zz_4545_ = int_reg_array_55_40_real;
      end
      6'b101001 : begin
        _zz_4544_ = int_reg_array_55_41_imag;
        _zz_4545_ = int_reg_array_55_41_real;
      end
      6'b101010 : begin
        _zz_4544_ = int_reg_array_55_42_imag;
        _zz_4545_ = int_reg_array_55_42_real;
      end
      6'b101011 : begin
        _zz_4544_ = int_reg_array_55_43_imag;
        _zz_4545_ = int_reg_array_55_43_real;
      end
      6'b101100 : begin
        _zz_4544_ = int_reg_array_55_44_imag;
        _zz_4545_ = int_reg_array_55_44_real;
      end
      6'b101101 : begin
        _zz_4544_ = int_reg_array_55_45_imag;
        _zz_4545_ = int_reg_array_55_45_real;
      end
      6'b101110 : begin
        _zz_4544_ = int_reg_array_55_46_imag;
        _zz_4545_ = int_reg_array_55_46_real;
      end
      6'b101111 : begin
        _zz_4544_ = int_reg_array_55_47_imag;
        _zz_4545_ = int_reg_array_55_47_real;
      end
      6'b110000 : begin
        _zz_4544_ = int_reg_array_55_48_imag;
        _zz_4545_ = int_reg_array_55_48_real;
      end
      6'b110001 : begin
        _zz_4544_ = int_reg_array_55_49_imag;
        _zz_4545_ = int_reg_array_55_49_real;
      end
      6'b110010 : begin
        _zz_4544_ = int_reg_array_55_50_imag;
        _zz_4545_ = int_reg_array_55_50_real;
      end
      6'b110011 : begin
        _zz_4544_ = int_reg_array_55_51_imag;
        _zz_4545_ = int_reg_array_55_51_real;
      end
      6'b110100 : begin
        _zz_4544_ = int_reg_array_55_52_imag;
        _zz_4545_ = int_reg_array_55_52_real;
      end
      6'b110101 : begin
        _zz_4544_ = int_reg_array_55_53_imag;
        _zz_4545_ = int_reg_array_55_53_real;
      end
      6'b110110 : begin
        _zz_4544_ = int_reg_array_55_54_imag;
        _zz_4545_ = int_reg_array_55_54_real;
      end
      6'b110111 : begin
        _zz_4544_ = int_reg_array_55_55_imag;
        _zz_4545_ = int_reg_array_55_55_real;
      end
      6'b111000 : begin
        _zz_4544_ = int_reg_array_55_56_imag;
        _zz_4545_ = int_reg_array_55_56_real;
      end
      6'b111001 : begin
        _zz_4544_ = int_reg_array_55_57_imag;
        _zz_4545_ = int_reg_array_55_57_real;
      end
      6'b111010 : begin
        _zz_4544_ = int_reg_array_55_58_imag;
        _zz_4545_ = int_reg_array_55_58_real;
      end
      6'b111011 : begin
        _zz_4544_ = int_reg_array_55_59_imag;
        _zz_4545_ = int_reg_array_55_59_real;
      end
      6'b111100 : begin
        _zz_4544_ = int_reg_array_55_60_imag;
        _zz_4545_ = int_reg_array_55_60_real;
      end
      6'b111101 : begin
        _zz_4544_ = int_reg_array_55_61_imag;
        _zz_4545_ = int_reg_array_55_61_real;
      end
      6'b111110 : begin
        _zz_4544_ = int_reg_array_55_62_imag;
        _zz_4545_ = int_reg_array_55_62_real;
      end
      default : begin
        _zz_4544_ = int_reg_array_55_63_imag;
        _zz_4545_ = int_reg_array_55_63_real;
      end
    endcase
  end

  always @(*) begin
    case(_zz_3881_)
      6'b000000 : begin
        _zz_4546_ = int_reg_array_56_0_imag;
        _zz_4547_ = int_reg_array_56_0_real;
      end
      6'b000001 : begin
        _zz_4546_ = int_reg_array_56_1_imag;
        _zz_4547_ = int_reg_array_56_1_real;
      end
      6'b000010 : begin
        _zz_4546_ = int_reg_array_56_2_imag;
        _zz_4547_ = int_reg_array_56_2_real;
      end
      6'b000011 : begin
        _zz_4546_ = int_reg_array_56_3_imag;
        _zz_4547_ = int_reg_array_56_3_real;
      end
      6'b000100 : begin
        _zz_4546_ = int_reg_array_56_4_imag;
        _zz_4547_ = int_reg_array_56_4_real;
      end
      6'b000101 : begin
        _zz_4546_ = int_reg_array_56_5_imag;
        _zz_4547_ = int_reg_array_56_5_real;
      end
      6'b000110 : begin
        _zz_4546_ = int_reg_array_56_6_imag;
        _zz_4547_ = int_reg_array_56_6_real;
      end
      6'b000111 : begin
        _zz_4546_ = int_reg_array_56_7_imag;
        _zz_4547_ = int_reg_array_56_7_real;
      end
      6'b001000 : begin
        _zz_4546_ = int_reg_array_56_8_imag;
        _zz_4547_ = int_reg_array_56_8_real;
      end
      6'b001001 : begin
        _zz_4546_ = int_reg_array_56_9_imag;
        _zz_4547_ = int_reg_array_56_9_real;
      end
      6'b001010 : begin
        _zz_4546_ = int_reg_array_56_10_imag;
        _zz_4547_ = int_reg_array_56_10_real;
      end
      6'b001011 : begin
        _zz_4546_ = int_reg_array_56_11_imag;
        _zz_4547_ = int_reg_array_56_11_real;
      end
      6'b001100 : begin
        _zz_4546_ = int_reg_array_56_12_imag;
        _zz_4547_ = int_reg_array_56_12_real;
      end
      6'b001101 : begin
        _zz_4546_ = int_reg_array_56_13_imag;
        _zz_4547_ = int_reg_array_56_13_real;
      end
      6'b001110 : begin
        _zz_4546_ = int_reg_array_56_14_imag;
        _zz_4547_ = int_reg_array_56_14_real;
      end
      6'b001111 : begin
        _zz_4546_ = int_reg_array_56_15_imag;
        _zz_4547_ = int_reg_array_56_15_real;
      end
      6'b010000 : begin
        _zz_4546_ = int_reg_array_56_16_imag;
        _zz_4547_ = int_reg_array_56_16_real;
      end
      6'b010001 : begin
        _zz_4546_ = int_reg_array_56_17_imag;
        _zz_4547_ = int_reg_array_56_17_real;
      end
      6'b010010 : begin
        _zz_4546_ = int_reg_array_56_18_imag;
        _zz_4547_ = int_reg_array_56_18_real;
      end
      6'b010011 : begin
        _zz_4546_ = int_reg_array_56_19_imag;
        _zz_4547_ = int_reg_array_56_19_real;
      end
      6'b010100 : begin
        _zz_4546_ = int_reg_array_56_20_imag;
        _zz_4547_ = int_reg_array_56_20_real;
      end
      6'b010101 : begin
        _zz_4546_ = int_reg_array_56_21_imag;
        _zz_4547_ = int_reg_array_56_21_real;
      end
      6'b010110 : begin
        _zz_4546_ = int_reg_array_56_22_imag;
        _zz_4547_ = int_reg_array_56_22_real;
      end
      6'b010111 : begin
        _zz_4546_ = int_reg_array_56_23_imag;
        _zz_4547_ = int_reg_array_56_23_real;
      end
      6'b011000 : begin
        _zz_4546_ = int_reg_array_56_24_imag;
        _zz_4547_ = int_reg_array_56_24_real;
      end
      6'b011001 : begin
        _zz_4546_ = int_reg_array_56_25_imag;
        _zz_4547_ = int_reg_array_56_25_real;
      end
      6'b011010 : begin
        _zz_4546_ = int_reg_array_56_26_imag;
        _zz_4547_ = int_reg_array_56_26_real;
      end
      6'b011011 : begin
        _zz_4546_ = int_reg_array_56_27_imag;
        _zz_4547_ = int_reg_array_56_27_real;
      end
      6'b011100 : begin
        _zz_4546_ = int_reg_array_56_28_imag;
        _zz_4547_ = int_reg_array_56_28_real;
      end
      6'b011101 : begin
        _zz_4546_ = int_reg_array_56_29_imag;
        _zz_4547_ = int_reg_array_56_29_real;
      end
      6'b011110 : begin
        _zz_4546_ = int_reg_array_56_30_imag;
        _zz_4547_ = int_reg_array_56_30_real;
      end
      6'b011111 : begin
        _zz_4546_ = int_reg_array_56_31_imag;
        _zz_4547_ = int_reg_array_56_31_real;
      end
      6'b100000 : begin
        _zz_4546_ = int_reg_array_56_32_imag;
        _zz_4547_ = int_reg_array_56_32_real;
      end
      6'b100001 : begin
        _zz_4546_ = int_reg_array_56_33_imag;
        _zz_4547_ = int_reg_array_56_33_real;
      end
      6'b100010 : begin
        _zz_4546_ = int_reg_array_56_34_imag;
        _zz_4547_ = int_reg_array_56_34_real;
      end
      6'b100011 : begin
        _zz_4546_ = int_reg_array_56_35_imag;
        _zz_4547_ = int_reg_array_56_35_real;
      end
      6'b100100 : begin
        _zz_4546_ = int_reg_array_56_36_imag;
        _zz_4547_ = int_reg_array_56_36_real;
      end
      6'b100101 : begin
        _zz_4546_ = int_reg_array_56_37_imag;
        _zz_4547_ = int_reg_array_56_37_real;
      end
      6'b100110 : begin
        _zz_4546_ = int_reg_array_56_38_imag;
        _zz_4547_ = int_reg_array_56_38_real;
      end
      6'b100111 : begin
        _zz_4546_ = int_reg_array_56_39_imag;
        _zz_4547_ = int_reg_array_56_39_real;
      end
      6'b101000 : begin
        _zz_4546_ = int_reg_array_56_40_imag;
        _zz_4547_ = int_reg_array_56_40_real;
      end
      6'b101001 : begin
        _zz_4546_ = int_reg_array_56_41_imag;
        _zz_4547_ = int_reg_array_56_41_real;
      end
      6'b101010 : begin
        _zz_4546_ = int_reg_array_56_42_imag;
        _zz_4547_ = int_reg_array_56_42_real;
      end
      6'b101011 : begin
        _zz_4546_ = int_reg_array_56_43_imag;
        _zz_4547_ = int_reg_array_56_43_real;
      end
      6'b101100 : begin
        _zz_4546_ = int_reg_array_56_44_imag;
        _zz_4547_ = int_reg_array_56_44_real;
      end
      6'b101101 : begin
        _zz_4546_ = int_reg_array_56_45_imag;
        _zz_4547_ = int_reg_array_56_45_real;
      end
      6'b101110 : begin
        _zz_4546_ = int_reg_array_56_46_imag;
        _zz_4547_ = int_reg_array_56_46_real;
      end
      6'b101111 : begin
        _zz_4546_ = int_reg_array_56_47_imag;
        _zz_4547_ = int_reg_array_56_47_real;
      end
      6'b110000 : begin
        _zz_4546_ = int_reg_array_56_48_imag;
        _zz_4547_ = int_reg_array_56_48_real;
      end
      6'b110001 : begin
        _zz_4546_ = int_reg_array_56_49_imag;
        _zz_4547_ = int_reg_array_56_49_real;
      end
      6'b110010 : begin
        _zz_4546_ = int_reg_array_56_50_imag;
        _zz_4547_ = int_reg_array_56_50_real;
      end
      6'b110011 : begin
        _zz_4546_ = int_reg_array_56_51_imag;
        _zz_4547_ = int_reg_array_56_51_real;
      end
      6'b110100 : begin
        _zz_4546_ = int_reg_array_56_52_imag;
        _zz_4547_ = int_reg_array_56_52_real;
      end
      6'b110101 : begin
        _zz_4546_ = int_reg_array_56_53_imag;
        _zz_4547_ = int_reg_array_56_53_real;
      end
      6'b110110 : begin
        _zz_4546_ = int_reg_array_56_54_imag;
        _zz_4547_ = int_reg_array_56_54_real;
      end
      6'b110111 : begin
        _zz_4546_ = int_reg_array_56_55_imag;
        _zz_4547_ = int_reg_array_56_55_real;
      end
      6'b111000 : begin
        _zz_4546_ = int_reg_array_56_56_imag;
        _zz_4547_ = int_reg_array_56_56_real;
      end
      6'b111001 : begin
        _zz_4546_ = int_reg_array_56_57_imag;
        _zz_4547_ = int_reg_array_56_57_real;
      end
      6'b111010 : begin
        _zz_4546_ = int_reg_array_56_58_imag;
        _zz_4547_ = int_reg_array_56_58_real;
      end
      6'b111011 : begin
        _zz_4546_ = int_reg_array_56_59_imag;
        _zz_4547_ = int_reg_array_56_59_real;
      end
      6'b111100 : begin
        _zz_4546_ = int_reg_array_56_60_imag;
        _zz_4547_ = int_reg_array_56_60_real;
      end
      6'b111101 : begin
        _zz_4546_ = int_reg_array_56_61_imag;
        _zz_4547_ = int_reg_array_56_61_real;
      end
      6'b111110 : begin
        _zz_4546_ = int_reg_array_56_62_imag;
        _zz_4547_ = int_reg_array_56_62_real;
      end
      default : begin
        _zz_4546_ = int_reg_array_56_63_imag;
        _zz_4547_ = int_reg_array_56_63_real;
      end
    endcase
  end

  always @(*) begin
    case(_zz_3950_)
      6'b000000 : begin
        _zz_4548_ = int_reg_array_57_0_imag;
        _zz_4549_ = int_reg_array_57_0_real;
      end
      6'b000001 : begin
        _zz_4548_ = int_reg_array_57_1_imag;
        _zz_4549_ = int_reg_array_57_1_real;
      end
      6'b000010 : begin
        _zz_4548_ = int_reg_array_57_2_imag;
        _zz_4549_ = int_reg_array_57_2_real;
      end
      6'b000011 : begin
        _zz_4548_ = int_reg_array_57_3_imag;
        _zz_4549_ = int_reg_array_57_3_real;
      end
      6'b000100 : begin
        _zz_4548_ = int_reg_array_57_4_imag;
        _zz_4549_ = int_reg_array_57_4_real;
      end
      6'b000101 : begin
        _zz_4548_ = int_reg_array_57_5_imag;
        _zz_4549_ = int_reg_array_57_5_real;
      end
      6'b000110 : begin
        _zz_4548_ = int_reg_array_57_6_imag;
        _zz_4549_ = int_reg_array_57_6_real;
      end
      6'b000111 : begin
        _zz_4548_ = int_reg_array_57_7_imag;
        _zz_4549_ = int_reg_array_57_7_real;
      end
      6'b001000 : begin
        _zz_4548_ = int_reg_array_57_8_imag;
        _zz_4549_ = int_reg_array_57_8_real;
      end
      6'b001001 : begin
        _zz_4548_ = int_reg_array_57_9_imag;
        _zz_4549_ = int_reg_array_57_9_real;
      end
      6'b001010 : begin
        _zz_4548_ = int_reg_array_57_10_imag;
        _zz_4549_ = int_reg_array_57_10_real;
      end
      6'b001011 : begin
        _zz_4548_ = int_reg_array_57_11_imag;
        _zz_4549_ = int_reg_array_57_11_real;
      end
      6'b001100 : begin
        _zz_4548_ = int_reg_array_57_12_imag;
        _zz_4549_ = int_reg_array_57_12_real;
      end
      6'b001101 : begin
        _zz_4548_ = int_reg_array_57_13_imag;
        _zz_4549_ = int_reg_array_57_13_real;
      end
      6'b001110 : begin
        _zz_4548_ = int_reg_array_57_14_imag;
        _zz_4549_ = int_reg_array_57_14_real;
      end
      6'b001111 : begin
        _zz_4548_ = int_reg_array_57_15_imag;
        _zz_4549_ = int_reg_array_57_15_real;
      end
      6'b010000 : begin
        _zz_4548_ = int_reg_array_57_16_imag;
        _zz_4549_ = int_reg_array_57_16_real;
      end
      6'b010001 : begin
        _zz_4548_ = int_reg_array_57_17_imag;
        _zz_4549_ = int_reg_array_57_17_real;
      end
      6'b010010 : begin
        _zz_4548_ = int_reg_array_57_18_imag;
        _zz_4549_ = int_reg_array_57_18_real;
      end
      6'b010011 : begin
        _zz_4548_ = int_reg_array_57_19_imag;
        _zz_4549_ = int_reg_array_57_19_real;
      end
      6'b010100 : begin
        _zz_4548_ = int_reg_array_57_20_imag;
        _zz_4549_ = int_reg_array_57_20_real;
      end
      6'b010101 : begin
        _zz_4548_ = int_reg_array_57_21_imag;
        _zz_4549_ = int_reg_array_57_21_real;
      end
      6'b010110 : begin
        _zz_4548_ = int_reg_array_57_22_imag;
        _zz_4549_ = int_reg_array_57_22_real;
      end
      6'b010111 : begin
        _zz_4548_ = int_reg_array_57_23_imag;
        _zz_4549_ = int_reg_array_57_23_real;
      end
      6'b011000 : begin
        _zz_4548_ = int_reg_array_57_24_imag;
        _zz_4549_ = int_reg_array_57_24_real;
      end
      6'b011001 : begin
        _zz_4548_ = int_reg_array_57_25_imag;
        _zz_4549_ = int_reg_array_57_25_real;
      end
      6'b011010 : begin
        _zz_4548_ = int_reg_array_57_26_imag;
        _zz_4549_ = int_reg_array_57_26_real;
      end
      6'b011011 : begin
        _zz_4548_ = int_reg_array_57_27_imag;
        _zz_4549_ = int_reg_array_57_27_real;
      end
      6'b011100 : begin
        _zz_4548_ = int_reg_array_57_28_imag;
        _zz_4549_ = int_reg_array_57_28_real;
      end
      6'b011101 : begin
        _zz_4548_ = int_reg_array_57_29_imag;
        _zz_4549_ = int_reg_array_57_29_real;
      end
      6'b011110 : begin
        _zz_4548_ = int_reg_array_57_30_imag;
        _zz_4549_ = int_reg_array_57_30_real;
      end
      6'b011111 : begin
        _zz_4548_ = int_reg_array_57_31_imag;
        _zz_4549_ = int_reg_array_57_31_real;
      end
      6'b100000 : begin
        _zz_4548_ = int_reg_array_57_32_imag;
        _zz_4549_ = int_reg_array_57_32_real;
      end
      6'b100001 : begin
        _zz_4548_ = int_reg_array_57_33_imag;
        _zz_4549_ = int_reg_array_57_33_real;
      end
      6'b100010 : begin
        _zz_4548_ = int_reg_array_57_34_imag;
        _zz_4549_ = int_reg_array_57_34_real;
      end
      6'b100011 : begin
        _zz_4548_ = int_reg_array_57_35_imag;
        _zz_4549_ = int_reg_array_57_35_real;
      end
      6'b100100 : begin
        _zz_4548_ = int_reg_array_57_36_imag;
        _zz_4549_ = int_reg_array_57_36_real;
      end
      6'b100101 : begin
        _zz_4548_ = int_reg_array_57_37_imag;
        _zz_4549_ = int_reg_array_57_37_real;
      end
      6'b100110 : begin
        _zz_4548_ = int_reg_array_57_38_imag;
        _zz_4549_ = int_reg_array_57_38_real;
      end
      6'b100111 : begin
        _zz_4548_ = int_reg_array_57_39_imag;
        _zz_4549_ = int_reg_array_57_39_real;
      end
      6'b101000 : begin
        _zz_4548_ = int_reg_array_57_40_imag;
        _zz_4549_ = int_reg_array_57_40_real;
      end
      6'b101001 : begin
        _zz_4548_ = int_reg_array_57_41_imag;
        _zz_4549_ = int_reg_array_57_41_real;
      end
      6'b101010 : begin
        _zz_4548_ = int_reg_array_57_42_imag;
        _zz_4549_ = int_reg_array_57_42_real;
      end
      6'b101011 : begin
        _zz_4548_ = int_reg_array_57_43_imag;
        _zz_4549_ = int_reg_array_57_43_real;
      end
      6'b101100 : begin
        _zz_4548_ = int_reg_array_57_44_imag;
        _zz_4549_ = int_reg_array_57_44_real;
      end
      6'b101101 : begin
        _zz_4548_ = int_reg_array_57_45_imag;
        _zz_4549_ = int_reg_array_57_45_real;
      end
      6'b101110 : begin
        _zz_4548_ = int_reg_array_57_46_imag;
        _zz_4549_ = int_reg_array_57_46_real;
      end
      6'b101111 : begin
        _zz_4548_ = int_reg_array_57_47_imag;
        _zz_4549_ = int_reg_array_57_47_real;
      end
      6'b110000 : begin
        _zz_4548_ = int_reg_array_57_48_imag;
        _zz_4549_ = int_reg_array_57_48_real;
      end
      6'b110001 : begin
        _zz_4548_ = int_reg_array_57_49_imag;
        _zz_4549_ = int_reg_array_57_49_real;
      end
      6'b110010 : begin
        _zz_4548_ = int_reg_array_57_50_imag;
        _zz_4549_ = int_reg_array_57_50_real;
      end
      6'b110011 : begin
        _zz_4548_ = int_reg_array_57_51_imag;
        _zz_4549_ = int_reg_array_57_51_real;
      end
      6'b110100 : begin
        _zz_4548_ = int_reg_array_57_52_imag;
        _zz_4549_ = int_reg_array_57_52_real;
      end
      6'b110101 : begin
        _zz_4548_ = int_reg_array_57_53_imag;
        _zz_4549_ = int_reg_array_57_53_real;
      end
      6'b110110 : begin
        _zz_4548_ = int_reg_array_57_54_imag;
        _zz_4549_ = int_reg_array_57_54_real;
      end
      6'b110111 : begin
        _zz_4548_ = int_reg_array_57_55_imag;
        _zz_4549_ = int_reg_array_57_55_real;
      end
      6'b111000 : begin
        _zz_4548_ = int_reg_array_57_56_imag;
        _zz_4549_ = int_reg_array_57_56_real;
      end
      6'b111001 : begin
        _zz_4548_ = int_reg_array_57_57_imag;
        _zz_4549_ = int_reg_array_57_57_real;
      end
      6'b111010 : begin
        _zz_4548_ = int_reg_array_57_58_imag;
        _zz_4549_ = int_reg_array_57_58_real;
      end
      6'b111011 : begin
        _zz_4548_ = int_reg_array_57_59_imag;
        _zz_4549_ = int_reg_array_57_59_real;
      end
      6'b111100 : begin
        _zz_4548_ = int_reg_array_57_60_imag;
        _zz_4549_ = int_reg_array_57_60_real;
      end
      6'b111101 : begin
        _zz_4548_ = int_reg_array_57_61_imag;
        _zz_4549_ = int_reg_array_57_61_real;
      end
      6'b111110 : begin
        _zz_4548_ = int_reg_array_57_62_imag;
        _zz_4549_ = int_reg_array_57_62_real;
      end
      default : begin
        _zz_4548_ = int_reg_array_57_63_imag;
        _zz_4549_ = int_reg_array_57_63_real;
      end
    endcase
  end

  always @(*) begin
    case(_zz_4019_)
      6'b000000 : begin
        _zz_4550_ = int_reg_array_58_0_imag;
        _zz_4551_ = int_reg_array_58_0_real;
      end
      6'b000001 : begin
        _zz_4550_ = int_reg_array_58_1_imag;
        _zz_4551_ = int_reg_array_58_1_real;
      end
      6'b000010 : begin
        _zz_4550_ = int_reg_array_58_2_imag;
        _zz_4551_ = int_reg_array_58_2_real;
      end
      6'b000011 : begin
        _zz_4550_ = int_reg_array_58_3_imag;
        _zz_4551_ = int_reg_array_58_3_real;
      end
      6'b000100 : begin
        _zz_4550_ = int_reg_array_58_4_imag;
        _zz_4551_ = int_reg_array_58_4_real;
      end
      6'b000101 : begin
        _zz_4550_ = int_reg_array_58_5_imag;
        _zz_4551_ = int_reg_array_58_5_real;
      end
      6'b000110 : begin
        _zz_4550_ = int_reg_array_58_6_imag;
        _zz_4551_ = int_reg_array_58_6_real;
      end
      6'b000111 : begin
        _zz_4550_ = int_reg_array_58_7_imag;
        _zz_4551_ = int_reg_array_58_7_real;
      end
      6'b001000 : begin
        _zz_4550_ = int_reg_array_58_8_imag;
        _zz_4551_ = int_reg_array_58_8_real;
      end
      6'b001001 : begin
        _zz_4550_ = int_reg_array_58_9_imag;
        _zz_4551_ = int_reg_array_58_9_real;
      end
      6'b001010 : begin
        _zz_4550_ = int_reg_array_58_10_imag;
        _zz_4551_ = int_reg_array_58_10_real;
      end
      6'b001011 : begin
        _zz_4550_ = int_reg_array_58_11_imag;
        _zz_4551_ = int_reg_array_58_11_real;
      end
      6'b001100 : begin
        _zz_4550_ = int_reg_array_58_12_imag;
        _zz_4551_ = int_reg_array_58_12_real;
      end
      6'b001101 : begin
        _zz_4550_ = int_reg_array_58_13_imag;
        _zz_4551_ = int_reg_array_58_13_real;
      end
      6'b001110 : begin
        _zz_4550_ = int_reg_array_58_14_imag;
        _zz_4551_ = int_reg_array_58_14_real;
      end
      6'b001111 : begin
        _zz_4550_ = int_reg_array_58_15_imag;
        _zz_4551_ = int_reg_array_58_15_real;
      end
      6'b010000 : begin
        _zz_4550_ = int_reg_array_58_16_imag;
        _zz_4551_ = int_reg_array_58_16_real;
      end
      6'b010001 : begin
        _zz_4550_ = int_reg_array_58_17_imag;
        _zz_4551_ = int_reg_array_58_17_real;
      end
      6'b010010 : begin
        _zz_4550_ = int_reg_array_58_18_imag;
        _zz_4551_ = int_reg_array_58_18_real;
      end
      6'b010011 : begin
        _zz_4550_ = int_reg_array_58_19_imag;
        _zz_4551_ = int_reg_array_58_19_real;
      end
      6'b010100 : begin
        _zz_4550_ = int_reg_array_58_20_imag;
        _zz_4551_ = int_reg_array_58_20_real;
      end
      6'b010101 : begin
        _zz_4550_ = int_reg_array_58_21_imag;
        _zz_4551_ = int_reg_array_58_21_real;
      end
      6'b010110 : begin
        _zz_4550_ = int_reg_array_58_22_imag;
        _zz_4551_ = int_reg_array_58_22_real;
      end
      6'b010111 : begin
        _zz_4550_ = int_reg_array_58_23_imag;
        _zz_4551_ = int_reg_array_58_23_real;
      end
      6'b011000 : begin
        _zz_4550_ = int_reg_array_58_24_imag;
        _zz_4551_ = int_reg_array_58_24_real;
      end
      6'b011001 : begin
        _zz_4550_ = int_reg_array_58_25_imag;
        _zz_4551_ = int_reg_array_58_25_real;
      end
      6'b011010 : begin
        _zz_4550_ = int_reg_array_58_26_imag;
        _zz_4551_ = int_reg_array_58_26_real;
      end
      6'b011011 : begin
        _zz_4550_ = int_reg_array_58_27_imag;
        _zz_4551_ = int_reg_array_58_27_real;
      end
      6'b011100 : begin
        _zz_4550_ = int_reg_array_58_28_imag;
        _zz_4551_ = int_reg_array_58_28_real;
      end
      6'b011101 : begin
        _zz_4550_ = int_reg_array_58_29_imag;
        _zz_4551_ = int_reg_array_58_29_real;
      end
      6'b011110 : begin
        _zz_4550_ = int_reg_array_58_30_imag;
        _zz_4551_ = int_reg_array_58_30_real;
      end
      6'b011111 : begin
        _zz_4550_ = int_reg_array_58_31_imag;
        _zz_4551_ = int_reg_array_58_31_real;
      end
      6'b100000 : begin
        _zz_4550_ = int_reg_array_58_32_imag;
        _zz_4551_ = int_reg_array_58_32_real;
      end
      6'b100001 : begin
        _zz_4550_ = int_reg_array_58_33_imag;
        _zz_4551_ = int_reg_array_58_33_real;
      end
      6'b100010 : begin
        _zz_4550_ = int_reg_array_58_34_imag;
        _zz_4551_ = int_reg_array_58_34_real;
      end
      6'b100011 : begin
        _zz_4550_ = int_reg_array_58_35_imag;
        _zz_4551_ = int_reg_array_58_35_real;
      end
      6'b100100 : begin
        _zz_4550_ = int_reg_array_58_36_imag;
        _zz_4551_ = int_reg_array_58_36_real;
      end
      6'b100101 : begin
        _zz_4550_ = int_reg_array_58_37_imag;
        _zz_4551_ = int_reg_array_58_37_real;
      end
      6'b100110 : begin
        _zz_4550_ = int_reg_array_58_38_imag;
        _zz_4551_ = int_reg_array_58_38_real;
      end
      6'b100111 : begin
        _zz_4550_ = int_reg_array_58_39_imag;
        _zz_4551_ = int_reg_array_58_39_real;
      end
      6'b101000 : begin
        _zz_4550_ = int_reg_array_58_40_imag;
        _zz_4551_ = int_reg_array_58_40_real;
      end
      6'b101001 : begin
        _zz_4550_ = int_reg_array_58_41_imag;
        _zz_4551_ = int_reg_array_58_41_real;
      end
      6'b101010 : begin
        _zz_4550_ = int_reg_array_58_42_imag;
        _zz_4551_ = int_reg_array_58_42_real;
      end
      6'b101011 : begin
        _zz_4550_ = int_reg_array_58_43_imag;
        _zz_4551_ = int_reg_array_58_43_real;
      end
      6'b101100 : begin
        _zz_4550_ = int_reg_array_58_44_imag;
        _zz_4551_ = int_reg_array_58_44_real;
      end
      6'b101101 : begin
        _zz_4550_ = int_reg_array_58_45_imag;
        _zz_4551_ = int_reg_array_58_45_real;
      end
      6'b101110 : begin
        _zz_4550_ = int_reg_array_58_46_imag;
        _zz_4551_ = int_reg_array_58_46_real;
      end
      6'b101111 : begin
        _zz_4550_ = int_reg_array_58_47_imag;
        _zz_4551_ = int_reg_array_58_47_real;
      end
      6'b110000 : begin
        _zz_4550_ = int_reg_array_58_48_imag;
        _zz_4551_ = int_reg_array_58_48_real;
      end
      6'b110001 : begin
        _zz_4550_ = int_reg_array_58_49_imag;
        _zz_4551_ = int_reg_array_58_49_real;
      end
      6'b110010 : begin
        _zz_4550_ = int_reg_array_58_50_imag;
        _zz_4551_ = int_reg_array_58_50_real;
      end
      6'b110011 : begin
        _zz_4550_ = int_reg_array_58_51_imag;
        _zz_4551_ = int_reg_array_58_51_real;
      end
      6'b110100 : begin
        _zz_4550_ = int_reg_array_58_52_imag;
        _zz_4551_ = int_reg_array_58_52_real;
      end
      6'b110101 : begin
        _zz_4550_ = int_reg_array_58_53_imag;
        _zz_4551_ = int_reg_array_58_53_real;
      end
      6'b110110 : begin
        _zz_4550_ = int_reg_array_58_54_imag;
        _zz_4551_ = int_reg_array_58_54_real;
      end
      6'b110111 : begin
        _zz_4550_ = int_reg_array_58_55_imag;
        _zz_4551_ = int_reg_array_58_55_real;
      end
      6'b111000 : begin
        _zz_4550_ = int_reg_array_58_56_imag;
        _zz_4551_ = int_reg_array_58_56_real;
      end
      6'b111001 : begin
        _zz_4550_ = int_reg_array_58_57_imag;
        _zz_4551_ = int_reg_array_58_57_real;
      end
      6'b111010 : begin
        _zz_4550_ = int_reg_array_58_58_imag;
        _zz_4551_ = int_reg_array_58_58_real;
      end
      6'b111011 : begin
        _zz_4550_ = int_reg_array_58_59_imag;
        _zz_4551_ = int_reg_array_58_59_real;
      end
      6'b111100 : begin
        _zz_4550_ = int_reg_array_58_60_imag;
        _zz_4551_ = int_reg_array_58_60_real;
      end
      6'b111101 : begin
        _zz_4550_ = int_reg_array_58_61_imag;
        _zz_4551_ = int_reg_array_58_61_real;
      end
      6'b111110 : begin
        _zz_4550_ = int_reg_array_58_62_imag;
        _zz_4551_ = int_reg_array_58_62_real;
      end
      default : begin
        _zz_4550_ = int_reg_array_58_63_imag;
        _zz_4551_ = int_reg_array_58_63_real;
      end
    endcase
  end

  always @(*) begin
    case(_zz_4088_)
      6'b000000 : begin
        _zz_4552_ = int_reg_array_59_0_imag;
        _zz_4553_ = int_reg_array_59_0_real;
      end
      6'b000001 : begin
        _zz_4552_ = int_reg_array_59_1_imag;
        _zz_4553_ = int_reg_array_59_1_real;
      end
      6'b000010 : begin
        _zz_4552_ = int_reg_array_59_2_imag;
        _zz_4553_ = int_reg_array_59_2_real;
      end
      6'b000011 : begin
        _zz_4552_ = int_reg_array_59_3_imag;
        _zz_4553_ = int_reg_array_59_3_real;
      end
      6'b000100 : begin
        _zz_4552_ = int_reg_array_59_4_imag;
        _zz_4553_ = int_reg_array_59_4_real;
      end
      6'b000101 : begin
        _zz_4552_ = int_reg_array_59_5_imag;
        _zz_4553_ = int_reg_array_59_5_real;
      end
      6'b000110 : begin
        _zz_4552_ = int_reg_array_59_6_imag;
        _zz_4553_ = int_reg_array_59_6_real;
      end
      6'b000111 : begin
        _zz_4552_ = int_reg_array_59_7_imag;
        _zz_4553_ = int_reg_array_59_7_real;
      end
      6'b001000 : begin
        _zz_4552_ = int_reg_array_59_8_imag;
        _zz_4553_ = int_reg_array_59_8_real;
      end
      6'b001001 : begin
        _zz_4552_ = int_reg_array_59_9_imag;
        _zz_4553_ = int_reg_array_59_9_real;
      end
      6'b001010 : begin
        _zz_4552_ = int_reg_array_59_10_imag;
        _zz_4553_ = int_reg_array_59_10_real;
      end
      6'b001011 : begin
        _zz_4552_ = int_reg_array_59_11_imag;
        _zz_4553_ = int_reg_array_59_11_real;
      end
      6'b001100 : begin
        _zz_4552_ = int_reg_array_59_12_imag;
        _zz_4553_ = int_reg_array_59_12_real;
      end
      6'b001101 : begin
        _zz_4552_ = int_reg_array_59_13_imag;
        _zz_4553_ = int_reg_array_59_13_real;
      end
      6'b001110 : begin
        _zz_4552_ = int_reg_array_59_14_imag;
        _zz_4553_ = int_reg_array_59_14_real;
      end
      6'b001111 : begin
        _zz_4552_ = int_reg_array_59_15_imag;
        _zz_4553_ = int_reg_array_59_15_real;
      end
      6'b010000 : begin
        _zz_4552_ = int_reg_array_59_16_imag;
        _zz_4553_ = int_reg_array_59_16_real;
      end
      6'b010001 : begin
        _zz_4552_ = int_reg_array_59_17_imag;
        _zz_4553_ = int_reg_array_59_17_real;
      end
      6'b010010 : begin
        _zz_4552_ = int_reg_array_59_18_imag;
        _zz_4553_ = int_reg_array_59_18_real;
      end
      6'b010011 : begin
        _zz_4552_ = int_reg_array_59_19_imag;
        _zz_4553_ = int_reg_array_59_19_real;
      end
      6'b010100 : begin
        _zz_4552_ = int_reg_array_59_20_imag;
        _zz_4553_ = int_reg_array_59_20_real;
      end
      6'b010101 : begin
        _zz_4552_ = int_reg_array_59_21_imag;
        _zz_4553_ = int_reg_array_59_21_real;
      end
      6'b010110 : begin
        _zz_4552_ = int_reg_array_59_22_imag;
        _zz_4553_ = int_reg_array_59_22_real;
      end
      6'b010111 : begin
        _zz_4552_ = int_reg_array_59_23_imag;
        _zz_4553_ = int_reg_array_59_23_real;
      end
      6'b011000 : begin
        _zz_4552_ = int_reg_array_59_24_imag;
        _zz_4553_ = int_reg_array_59_24_real;
      end
      6'b011001 : begin
        _zz_4552_ = int_reg_array_59_25_imag;
        _zz_4553_ = int_reg_array_59_25_real;
      end
      6'b011010 : begin
        _zz_4552_ = int_reg_array_59_26_imag;
        _zz_4553_ = int_reg_array_59_26_real;
      end
      6'b011011 : begin
        _zz_4552_ = int_reg_array_59_27_imag;
        _zz_4553_ = int_reg_array_59_27_real;
      end
      6'b011100 : begin
        _zz_4552_ = int_reg_array_59_28_imag;
        _zz_4553_ = int_reg_array_59_28_real;
      end
      6'b011101 : begin
        _zz_4552_ = int_reg_array_59_29_imag;
        _zz_4553_ = int_reg_array_59_29_real;
      end
      6'b011110 : begin
        _zz_4552_ = int_reg_array_59_30_imag;
        _zz_4553_ = int_reg_array_59_30_real;
      end
      6'b011111 : begin
        _zz_4552_ = int_reg_array_59_31_imag;
        _zz_4553_ = int_reg_array_59_31_real;
      end
      6'b100000 : begin
        _zz_4552_ = int_reg_array_59_32_imag;
        _zz_4553_ = int_reg_array_59_32_real;
      end
      6'b100001 : begin
        _zz_4552_ = int_reg_array_59_33_imag;
        _zz_4553_ = int_reg_array_59_33_real;
      end
      6'b100010 : begin
        _zz_4552_ = int_reg_array_59_34_imag;
        _zz_4553_ = int_reg_array_59_34_real;
      end
      6'b100011 : begin
        _zz_4552_ = int_reg_array_59_35_imag;
        _zz_4553_ = int_reg_array_59_35_real;
      end
      6'b100100 : begin
        _zz_4552_ = int_reg_array_59_36_imag;
        _zz_4553_ = int_reg_array_59_36_real;
      end
      6'b100101 : begin
        _zz_4552_ = int_reg_array_59_37_imag;
        _zz_4553_ = int_reg_array_59_37_real;
      end
      6'b100110 : begin
        _zz_4552_ = int_reg_array_59_38_imag;
        _zz_4553_ = int_reg_array_59_38_real;
      end
      6'b100111 : begin
        _zz_4552_ = int_reg_array_59_39_imag;
        _zz_4553_ = int_reg_array_59_39_real;
      end
      6'b101000 : begin
        _zz_4552_ = int_reg_array_59_40_imag;
        _zz_4553_ = int_reg_array_59_40_real;
      end
      6'b101001 : begin
        _zz_4552_ = int_reg_array_59_41_imag;
        _zz_4553_ = int_reg_array_59_41_real;
      end
      6'b101010 : begin
        _zz_4552_ = int_reg_array_59_42_imag;
        _zz_4553_ = int_reg_array_59_42_real;
      end
      6'b101011 : begin
        _zz_4552_ = int_reg_array_59_43_imag;
        _zz_4553_ = int_reg_array_59_43_real;
      end
      6'b101100 : begin
        _zz_4552_ = int_reg_array_59_44_imag;
        _zz_4553_ = int_reg_array_59_44_real;
      end
      6'b101101 : begin
        _zz_4552_ = int_reg_array_59_45_imag;
        _zz_4553_ = int_reg_array_59_45_real;
      end
      6'b101110 : begin
        _zz_4552_ = int_reg_array_59_46_imag;
        _zz_4553_ = int_reg_array_59_46_real;
      end
      6'b101111 : begin
        _zz_4552_ = int_reg_array_59_47_imag;
        _zz_4553_ = int_reg_array_59_47_real;
      end
      6'b110000 : begin
        _zz_4552_ = int_reg_array_59_48_imag;
        _zz_4553_ = int_reg_array_59_48_real;
      end
      6'b110001 : begin
        _zz_4552_ = int_reg_array_59_49_imag;
        _zz_4553_ = int_reg_array_59_49_real;
      end
      6'b110010 : begin
        _zz_4552_ = int_reg_array_59_50_imag;
        _zz_4553_ = int_reg_array_59_50_real;
      end
      6'b110011 : begin
        _zz_4552_ = int_reg_array_59_51_imag;
        _zz_4553_ = int_reg_array_59_51_real;
      end
      6'b110100 : begin
        _zz_4552_ = int_reg_array_59_52_imag;
        _zz_4553_ = int_reg_array_59_52_real;
      end
      6'b110101 : begin
        _zz_4552_ = int_reg_array_59_53_imag;
        _zz_4553_ = int_reg_array_59_53_real;
      end
      6'b110110 : begin
        _zz_4552_ = int_reg_array_59_54_imag;
        _zz_4553_ = int_reg_array_59_54_real;
      end
      6'b110111 : begin
        _zz_4552_ = int_reg_array_59_55_imag;
        _zz_4553_ = int_reg_array_59_55_real;
      end
      6'b111000 : begin
        _zz_4552_ = int_reg_array_59_56_imag;
        _zz_4553_ = int_reg_array_59_56_real;
      end
      6'b111001 : begin
        _zz_4552_ = int_reg_array_59_57_imag;
        _zz_4553_ = int_reg_array_59_57_real;
      end
      6'b111010 : begin
        _zz_4552_ = int_reg_array_59_58_imag;
        _zz_4553_ = int_reg_array_59_58_real;
      end
      6'b111011 : begin
        _zz_4552_ = int_reg_array_59_59_imag;
        _zz_4553_ = int_reg_array_59_59_real;
      end
      6'b111100 : begin
        _zz_4552_ = int_reg_array_59_60_imag;
        _zz_4553_ = int_reg_array_59_60_real;
      end
      6'b111101 : begin
        _zz_4552_ = int_reg_array_59_61_imag;
        _zz_4553_ = int_reg_array_59_61_real;
      end
      6'b111110 : begin
        _zz_4552_ = int_reg_array_59_62_imag;
        _zz_4553_ = int_reg_array_59_62_real;
      end
      default : begin
        _zz_4552_ = int_reg_array_59_63_imag;
        _zz_4553_ = int_reg_array_59_63_real;
      end
    endcase
  end

  always @(*) begin
    case(_zz_4157_)
      6'b000000 : begin
        _zz_4554_ = int_reg_array_60_0_imag;
        _zz_4555_ = int_reg_array_60_0_real;
      end
      6'b000001 : begin
        _zz_4554_ = int_reg_array_60_1_imag;
        _zz_4555_ = int_reg_array_60_1_real;
      end
      6'b000010 : begin
        _zz_4554_ = int_reg_array_60_2_imag;
        _zz_4555_ = int_reg_array_60_2_real;
      end
      6'b000011 : begin
        _zz_4554_ = int_reg_array_60_3_imag;
        _zz_4555_ = int_reg_array_60_3_real;
      end
      6'b000100 : begin
        _zz_4554_ = int_reg_array_60_4_imag;
        _zz_4555_ = int_reg_array_60_4_real;
      end
      6'b000101 : begin
        _zz_4554_ = int_reg_array_60_5_imag;
        _zz_4555_ = int_reg_array_60_5_real;
      end
      6'b000110 : begin
        _zz_4554_ = int_reg_array_60_6_imag;
        _zz_4555_ = int_reg_array_60_6_real;
      end
      6'b000111 : begin
        _zz_4554_ = int_reg_array_60_7_imag;
        _zz_4555_ = int_reg_array_60_7_real;
      end
      6'b001000 : begin
        _zz_4554_ = int_reg_array_60_8_imag;
        _zz_4555_ = int_reg_array_60_8_real;
      end
      6'b001001 : begin
        _zz_4554_ = int_reg_array_60_9_imag;
        _zz_4555_ = int_reg_array_60_9_real;
      end
      6'b001010 : begin
        _zz_4554_ = int_reg_array_60_10_imag;
        _zz_4555_ = int_reg_array_60_10_real;
      end
      6'b001011 : begin
        _zz_4554_ = int_reg_array_60_11_imag;
        _zz_4555_ = int_reg_array_60_11_real;
      end
      6'b001100 : begin
        _zz_4554_ = int_reg_array_60_12_imag;
        _zz_4555_ = int_reg_array_60_12_real;
      end
      6'b001101 : begin
        _zz_4554_ = int_reg_array_60_13_imag;
        _zz_4555_ = int_reg_array_60_13_real;
      end
      6'b001110 : begin
        _zz_4554_ = int_reg_array_60_14_imag;
        _zz_4555_ = int_reg_array_60_14_real;
      end
      6'b001111 : begin
        _zz_4554_ = int_reg_array_60_15_imag;
        _zz_4555_ = int_reg_array_60_15_real;
      end
      6'b010000 : begin
        _zz_4554_ = int_reg_array_60_16_imag;
        _zz_4555_ = int_reg_array_60_16_real;
      end
      6'b010001 : begin
        _zz_4554_ = int_reg_array_60_17_imag;
        _zz_4555_ = int_reg_array_60_17_real;
      end
      6'b010010 : begin
        _zz_4554_ = int_reg_array_60_18_imag;
        _zz_4555_ = int_reg_array_60_18_real;
      end
      6'b010011 : begin
        _zz_4554_ = int_reg_array_60_19_imag;
        _zz_4555_ = int_reg_array_60_19_real;
      end
      6'b010100 : begin
        _zz_4554_ = int_reg_array_60_20_imag;
        _zz_4555_ = int_reg_array_60_20_real;
      end
      6'b010101 : begin
        _zz_4554_ = int_reg_array_60_21_imag;
        _zz_4555_ = int_reg_array_60_21_real;
      end
      6'b010110 : begin
        _zz_4554_ = int_reg_array_60_22_imag;
        _zz_4555_ = int_reg_array_60_22_real;
      end
      6'b010111 : begin
        _zz_4554_ = int_reg_array_60_23_imag;
        _zz_4555_ = int_reg_array_60_23_real;
      end
      6'b011000 : begin
        _zz_4554_ = int_reg_array_60_24_imag;
        _zz_4555_ = int_reg_array_60_24_real;
      end
      6'b011001 : begin
        _zz_4554_ = int_reg_array_60_25_imag;
        _zz_4555_ = int_reg_array_60_25_real;
      end
      6'b011010 : begin
        _zz_4554_ = int_reg_array_60_26_imag;
        _zz_4555_ = int_reg_array_60_26_real;
      end
      6'b011011 : begin
        _zz_4554_ = int_reg_array_60_27_imag;
        _zz_4555_ = int_reg_array_60_27_real;
      end
      6'b011100 : begin
        _zz_4554_ = int_reg_array_60_28_imag;
        _zz_4555_ = int_reg_array_60_28_real;
      end
      6'b011101 : begin
        _zz_4554_ = int_reg_array_60_29_imag;
        _zz_4555_ = int_reg_array_60_29_real;
      end
      6'b011110 : begin
        _zz_4554_ = int_reg_array_60_30_imag;
        _zz_4555_ = int_reg_array_60_30_real;
      end
      6'b011111 : begin
        _zz_4554_ = int_reg_array_60_31_imag;
        _zz_4555_ = int_reg_array_60_31_real;
      end
      6'b100000 : begin
        _zz_4554_ = int_reg_array_60_32_imag;
        _zz_4555_ = int_reg_array_60_32_real;
      end
      6'b100001 : begin
        _zz_4554_ = int_reg_array_60_33_imag;
        _zz_4555_ = int_reg_array_60_33_real;
      end
      6'b100010 : begin
        _zz_4554_ = int_reg_array_60_34_imag;
        _zz_4555_ = int_reg_array_60_34_real;
      end
      6'b100011 : begin
        _zz_4554_ = int_reg_array_60_35_imag;
        _zz_4555_ = int_reg_array_60_35_real;
      end
      6'b100100 : begin
        _zz_4554_ = int_reg_array_60_36_imag;
        _zz_4555_ = int_reg_array_60_36_real;
      end
      6'b100101 : begin
        _zz_4554_ = int_reg_array_60_37_imag;
        _zz_4555_ = int_reg_array_60_37_real;
      end
      6'b100110 : begin
        _zz_4554_ = int_reg_array_60_38_imag;
        _zz_4555_ = int_reg_array_60_38_real;
      end
      6'b100111 : begin
        _zz_4554_ = int_reg_array_60_39_imag;
        _zz_4555_ = int_reg_array_60_39_real;
      end
      6'b101000 : begin
        _zz_4554_ = int_reg_array_60_40_imag;
        _zz_4555_ = int_reg_array_60_40_real;
      end
      6'b101001 : begin
        _zz_4554_ = int_reg_array_60_41_imag;
        _zz_4555_ = int_reg_array_60_41_real;
      end
      6'b101010 : begin
        _zz_4554_ = int_reg_array_60_42_imag;
        _zz_4555_ = int_reg_array_60_42_real;
      end
      6'b101011 : begin
        _zz_4554_ = int_reg_array_60_43_imag;
        _zz_4555_ = int_reg_array_60_43_real;
      end
      6'b101100 : begin
        _zz_4554_ = int_reg_array_60_44_imag;
        _zz_4555_ = int_reg_array_60_44_real;
      end
      6'b101101 : begin
        _zz_4554_ = int_reg_array_60_45_imag;
        _zz_4555_ = int_reg_array_60_45_real;
      end
      6'b101110 : begin
        _zz_4554_ = int_reg_array_60_46_imag;
        _zz_4555_ = int_reg_array_60_46_real;
      end
      6'b101111 : begin
        _zz_4554_ = int_reg_array_60_47_imag;
        _zz_4555_ = int_reg_array_60_47_real;
      end
      6'b110000 : begin
        _zz_4554_ = int_reg_array_60_48_imag;
        _zz_4555_ = int_reg_array_60_48_real;
      end
      6'b110001 : begin
        _zz_4554_ = int_reg_array_60_49_imag;
        _zz_4555_ = int_reg_array_60_49_real;
      end
      6'b110010 : begin
        _zz_4554_ = int_reg_array_60_50_imag;
        _zz_4555_ = int_reg_array_60_50_real;
      end
      6'b110011 : begin
        _zz_4554_ = int_reg_array_60_51_imag;
        _zz_4555_ = int_reg_array_60_51_real;
      end
      6'b110100 : begin
        _zz_4554_ = int_reg_array_60_52_imag;
        _zz_4555_ = int_reg_array_60_52_real;
      end
      6'b110101 : begin
        _zz_4554_ = int_reg_array_60_53_imag;
        _zz_4555_ = int_reg_array_60_53_real;
      end
      6'b110110 : begin
        _zz_4554_ = int_reg_array_60_54_imag;
        _zz_4555_ = int_reg_array_60_54_real;
      end
      6'b110111 : begin
        _zz_4554_ = int_reg_array_60_55_imag;
        _zz_4555_ = int_reg_array_60_55_real;
      end
      6'b111000 : begin
        _zz_4554_ = int_reg_array_60_56_imag;
        _zz_4555_ = int_reg_array_60_56_real;
      end
      6'b111001 : begin
        _zz_4554_ = int_reg_array_60_57_imag;
        _zz_4555_ = int_reg_array_60_57_real;
      end
      6'b111010 : begin
        _zz_4554_ = int_reg_array_60_58_imag;
        _zz_4555_ = int_reg_array_60_58_real;
      end
      6'b111011 : begin
        _zz_4554_ = int_reg_array_60_59_imag;
        _zz_4555_ = int_reg_array_60_59_real;
      end
      6'b111100 : begin
        _zz_4554_ = int_reg_array_60_60_imag;
        _zz_4555_ = int_reg_array_60_60_real;
      end
      6'b111101 : begin
        _zz_4554_ = int_reg_array_60_61_imag;
        _zz_4555_ = int_reg_array_60_61_real;
      end
      6'b111110 : begin
        _zz_4554_ = int_reg_array_60_62_imag;
        _zz_4555_ = int_reg_array_60_62_real;
      end
      default : begin
        _zz_4554_ = int_reg_array_60_63_imag;
        _zz_4555_ = int_reg_array_60_63_real;
      end
    endcase
  end

  always @(*) begin
    case(_zz_4226_)
      6'b000000 : begin
        _zz_4556_ = int_reg_array_61_0_imag;
        _zz_4557_ = int_reg_array_61_0_real;
      end
      6'b000001 : begin
        _zz_4556_ = int_reg_array_61_1_imag;
        _zz_4557_ = int_reg_array_61_1_real;
      end
      6'b000010 : begin
        _zz_4556_ = int_reg_array_61_2_imag;
        _zz_4557_ = int_reg_array_61_2_real;
      end
      6'b000011 : begin
        _zz_4556_ = int_reg_array_61_3_imag;
        _zz_4557_ = int_reg_array_61_3_real;
      end
      6'b000100 : begin
        _zz_4556_ = int_reg_array_61_4_imag;
        _zz_4557_ = int_reg_array_61_4_real;
      end
      6'b000101 : begin
        _zz_4556_ = int_reg_array_61_5_imag;
        _zz_4557_ = int_reg_array_61_5_real;
      end
      6'b000110 : begin
        _zz_4556_ = int_reg_array_61_6_imag;
        _zz_4557_ = int_reg_array_61_6_real;
      end
      6'b000111 : begin
        _zz_4556_ = int_reg_array_61_7_imag;
        _zz_4557_ = int_reg_array_61_7_real;
      end
      6'b001000 : begin
        _zz_4556_ = int_reg_array_61_8_imag;
        _zz_4557_ = int_reg_array_61_8_real;
      end
      6'b001001 : begin
        _zz_4556_ = int_reg_array_61_9_imag;
        _zz_4557_ = int_reg_array_61_9_real;
      end
      6'b001010 : begin
        _zz_4556_ = int_reg_array_61_10_imag;
        _zz_4557_ = int_reg_array_61_10_real;
      end
      6'b001011 : begin
        _zz_4556_ = int_reg_array_61_11_imag;
        _zz_4557_ = int_reg_array_61_11_real;
      end
      6'b001100 : begin
        _zz_4556_ = int_reg_array_61_12_imag;
        _zz_4557_ = int_reg_array_61_12_real;
      end
      6'b001101 : begin
        _zz_4556_ = int_reg_array_61_13_imag;
        _zz_4557_ = int_reg_array_61_13_real;
      end
      6'b001110 : begin
        _zz_4556_ = int_reg_array_61_14_imag;
        _zz_4557_ = int_reg_array_61_14_real;
      end
      6'b001111 : begin
        _zz_4556_ = int_reg_array_61_15_imag;
        _zz_4557_ = int_reg_array_61_15_real;
      end
      6'b010000 : begin
        _zz_4556_ = int_reg_array_61_16_imag;
        _zz_4557_ = int_reg_array_61_16_real;
      end
      6'b010001 : begin
        _zz_4556_ = int_reg_array_61_17_imag;
        _zz_4557_ = int_reg_array_61_17_real;
      end
      6'b010010 : begin
        _zz_4556_ = int_reg_array_61_18_imag;
        _zz_4557_ = int_reg_array_61_18_real;
      end
      6'b010011 : begin
        _zz_4556_ = int_reg_array_61_19_imag;
        _zz_4557_ = int_reg_array_61_19_real;
      end
      6'b010100 : begin
        _zz_4556_ = int_reg_array_61_20_imag;
        _zz_4557_ = int_reg_array_61_20_real;
      end
      6'b010101 : begin
        _zz_4556_ = int_reg_array_61_21_imag;
        _zz_4557_ = int_reg_array_61_21_real;
      end
      6'b010110 : begin
        _zz_4556_ = int_reg_array_61_22_imag;
        _zz_4557_ = int_reg_array_61_22_real;
      end
      6'b010111 : begin
        _zz_4556_ = int_reg_array_61_23_imag;
        _zz_4557_ = int_reg_array_61_23_real;
      end
      6'b011000 : begin
        _zz_4556_ = int_reg_array_61_24_imag;
        _zz_4557_ = int_reg_array_61_24_real;
      end
      6'b011001 : begin
        _zz_4556_ = int_reg_array_61_25_imag;
        _zz_4557_ = int_reg_array_61_25_real;
      end
      6'b011010 : begin
        _zz_4556_ = int_reg_array_61_26_imag;
        _zz_4557_ = int_reg_array_61_26_real;
      end
      6'b011011 : begin
        _zz_4556_ = int_reg_array_61_27_imag;
        _zz_4557_ = int_reg_array_61_27_real;
      end
      6'b011100 : begin
        _zz_4556_ = int_reg_array_61_28_imag;
        _zz_4557_ = int_reg_array_61_28_real;
      end
      6'b011101 : begin
        _zz_4556_ = int_reg_array_61_29_imag;
        _zz_4557_ = int_reg_array_61_29_real;
      end
      6'b011110 : begin
        _zz_4556_ = int_reg_array_61_30_imag;
        _zz_4557_ = int_reg_array_61_30_real;
      end
      6'b011111 : begin
        _zz_4556_ = int_reg_array_61_31_imag;
        _zz_4557_ = int_reg_array_61_31_real;
      end
      6'b100000 : begin
        _zz_4556_ = int_reg_array_61_32_imag;
        _zz_4557_ = int_reg_array_61_32_real;
      end
      6'b100001 : begin
        _zz_4556_ = int_reg_array_61_33_imag;
        _zz_4557_ = int_reg_array_61_33_real;
      end
      6'b100010 : begin
        _zz_4556_ = int_reg_array_61_34_imag;
        _zz_4557_ = int_reg_array_61_34_real;
      end
      6'b100011 : begin
        _zz_4556_ = int_reg_array_61_35_imag;
        _zz_4557_ = int_reg_array_61_35_real;
      end
      6'b100100 : begin
        _zz_4556_ = int_reg_array_61_36_imag;
        _zz_4557_ = int_reg_array_61_36_real;
      end
      6'b100101 : begin
        _zz_4556_ = int_reg_array_61_37_imag;
        _zz_4557_ = int_reg_array_61_37_real;
      end
      6'b100110 : begin
        _zz_4556_ = int_reg_array_61_38_imag;
        _zz_4557_ = int_reg_array_61_38_real;
      end
      6'b100111 : begin
        _zz_4556_ = int_reg_array_61_39_imag;
        _zz_4557_ = int_reg_array_61_39_real;
      end
      6'b101000 : begin
        _zz_4556_ = int_reg_array_61_40_imag;
        _zz_4557_ = int_reg_array_61_40_real;
      end
      6'b101001 : begin
        _zz_4556_ = int_reg_array_61_41_imag;
        _zz_4557_ = int_reg_array_61_41_real;
      end
      6'b101010 : begin
        _zz_4556_ = int_reg_array_61_42_imag;
        _zz_4557_ = int_reg_array_61_42_real;
      end
      6'b101011 : begin
        _zz_4556_ = int_reg_array_61_43_imag;
        _zz_4557_ = int_reg_array_61_43_real;
      end
      6'b101100 : begin
        _zz_4556_ = int_reg_array_61_44_imag;
        _zz_4557_ = int_reg_array_61_44_real;
      end
      6'b101101 : begin
        _zz_4556_ = int_reg_array_61_45_imag;
        _zz_4557_ = int_reg_array_61_45_real;
      end
      6'b101110 : begin
        _zz_4556_ = int_reg_array_61_46_imag;
        _zz_4557_ = int_reg_array_61_46_real;
      end
      6'b101111 : begin
        _zz_4556_ = int_reg_array_61_47_imag;
        _zz_4557_ = int_reg_array_61_47_real;
      end
      6'b110000 : begin
        _zz_4556_ = int_reg_array_61_48_imag;
        _zz_4557_ = int_reg_array_61_48_real;
      end
      6'b110001 : begin
        _zz_4556_ = int_reg_array_61_49_imag;
        _zz_4557_ = int_reg_array_61_49_real;
      end
      6'b110010 : begin
        _zz_4556_ = int_reg_array_61_50_imag;
        _zz_4557_ = int_reg_array_61_50_real;
      end
      6'b110011 : begin
        _zz_4556_ = int_reg_array_61_51_imag;
        _zz_4557_ = int_reg_array_61_51_real;
      end
      6'b110100 : begin
        _zz_4556_ = int_reg_array_61_52_imag;
        _zz_4557_ = int_reg_array_61_52_real;
      end
      6'b110101 : begin
        _zz_4556_ = int_reg_array_61_53_imag;
        _zz_4557_ = int_reg_array_61_53_real;
      end
      6'b110110 : begin
        _zz_4556_ = int_reg_array_61_54_imag;
        _zz_4557_ = int_reg_array_61_54_real;
      end
      6'b110111 : begin
        _zz_4556_ = int_reg_array_61_55_imag;
        _zz_4557_ = int_reg_array_61_55_real;
      end
      6'b111000 : begin
        _zz_4556_ = int_reg_array_61_56_imag;
        _zz_4557_ = int_reg_array_61_56_real;
      end
      6'b111001 : begin
        _zz_4556_ = int_reg_array_61_57_imag;
        _zz_4557_ = int_reg_array_61_57_real;
      end
      6'b111010 : begin
        _zz_4556_ = int_reg_array_61_58_imag;
        _zz_4557_ = int_reg_array_61_58_real;
      end
      6'b111011 : begin
        _zz_4556_ = int_reg_array_61_59_imag;
        _zz_4557_ = int_reg_array_61_59_real;
      end
      6'b111100 : begin
        _zz_4556_ = int_reg_array_61_60_imag;
        _zz_4557_ = int_reg_array_61_60_real;
      end
      6'b111101 : begin
        _zz_4556_ = int_reg_array_61_61_imag;
        _zz_4557_ = int_reg_array_61_61_real;
      end
      6'b111110 : begin
        _zz_4556_ = int_reg_array_61_62_imag;
        _zz_4557_ = int_reg_array_61_62_real;
      end
      default : begin
        _zz_4556_ = int_reg_array_61_63_imag;
        _zz_4557_ = int_reg_array_61_63_real;
      end
    endcase
  end

  always @(*) begin
    case(_zz_4295_)
      6'b000000 : begin
        _zz_4558_ = int_reg_array_62_0_imag;
        _zz_4559_ = int_reg_array_62_0_real;
      end
      6'b000001 : begin
        _zz_4558_ = int_reg_array_62_1_imag;
        _zz_4559_ = int_reg_array_62_1_real;
      end
      6'b000010 : begin
        _zz_4558_ = int_reg_array_62_2_imag;
        _zz_4559_ = int_reg_array_62_2_real;
      end
      6'b000011 : begin
        _zz_4558_ = int_reg_array_62_3_imag;
        _zz_4559_ = int_reg_array_62_3_real;
      end
      6'b000100 : begin
        _zz_4558_ = int_reg_array_62_4_imag;
        _zz_4559_ = int_reg_array_62_4_real;
      end
      6'b000101 : begin
        _zz_4558_ = int_reg_array_62_5_imag;
        _zz_4559_ = int_reg_array_62_5_real;
      end
      6'b000110 : begin
        _zz_4558_ = int_reg_array_62_6_imag;
        _zz_4559_ = int_reg_array_62_6_real;
      end
      6'b000111 : begin
        _zz_4558_ = int_reg_array_62_7_imag;
        _zz_4559_ = int_reg_array_62_7_real;
      end
      6'b001000 : begin
        _zz_4558_ = int_reg_array_62_8_imag;
        _zz_4559_ = int_reg_array_62_8_real;
      end
      6'b001001 : begin
        _zz_4558_ = int_reg_array_62_9_imag;
        _zz_4559_ = int_reg_array_62_9_real;
      end
      6'b001010 : begin
        _zz_4558_ = int_reg_array_62_10_imag;
        _zz_4559_ = int_reg_array_62_10_real;
      end
      6'b001011 : begin
        _zz_4558_ = int_reg_array_62_11_imag;
        _zz_4559_ = int_reg_array_62_11_real;
      end
      6'b001100 : begin
        _zz_4558_ = int_reg_array_62_12_imag;
        _zz_4559_ = int_reg_array_62_12_real;
      end
      6'b001101 : begin
        _zz_4558_ = int_reg_array_62_13_imag;
        _zz_4559_ = int_reg_array_62_13_real;
      end
      6'b001110 : begin
        _zz_4558_ = int_reg_array_62_14_imag;
        _zz_4559_ = int_reg_array_62_14_real;
      end
      6'b001111 : begin
        _zz_4558_ = int_reg_array_62_15_imag;
        _zz_4559_ = int_reg_array_62_15_real;
      end
      6'b010000 : begin
        _zz_4558_ = int_reg_array_62_16_imag;
        _zz_4559_ = int_reg_array_62_16_real;
      end
      6'b010001 : begin
        _zz_4558_ = int_reg_array_62_17_imag;
        _zz_4559_ = int_reg_array_62_17_real;
      end
      6'b010010 : begin
        _zz_4558_ = int_reg_array_62_18_imag;
        _zz_4559_ = int_reg_array_62_18_real;
      end
      6'b010011 : begin
        _zz_4558_ = int_reg_array_62_19_imag;
        _zz_4559_ = int_reg_array_62_19_real;
      end
      6'b010100 : begin
        _zz_4558_ = int_reg_array_62_20_imag;
        _zz_4559_ = int_reg_array_62_20_real;
      end
      6'b010101 : begin
        _zz_4558_ = int_reg_array_62_21_imag;
        _zz_4559_ = int_reg_array_62_21_real;
      end
      6'b010110 : begin
        _zz_4558_ = int_reg_array_62_22_imag;
        _zz_4559_ = int_reg_array_62_22_real;
      end
      6'b010111 : begin
        _zz_4558_ = int_reg_array_62_23_imag;
        _zz_4559_ = int_reg_array_62_23_real;
      end
      6'b011000 : begin
        _zz_4558_ = int_reg_array_62_24_imag;
        _zz_4559_ = int_reg_array_62_24_real;
      end
      6'b011001 : begin
        _zz_4558_ = int_reg_array_62_25_imag;
        _zz_4559_ = int_reg_array_62_25_real;
      end
      6'b011010 : begin
        _zz_4558_ = int_reg_array_62_26_imag;
        _zz_4559_ = int_reg_array_62_26_real;
      end
      6'b011011 : begin
        _zz_4558_ = int_reg_array_62_27_imag;
        _zz_4559_ = int_reg_array_62_27_real;
      end
      6'b011100 : begin
        _zz_4558_ = int_reg_array_62_28_imag;
        _zz_4559_ = int_reg_array_62_28_real;
      end
      6'b011101 : begin
        _zz_4558_ = int_reg_array_62_29_imag;
        _zz_4559_ = int_reg_array_62_29_real;
      end
      6'b011110 : begin
        _zz_4558_ = int_reg_array_62_30_imag;
        _zz_4559_ = int_reg_array_62_30_real;
      end
      6'b011111 : begin
        _zz_4558_ = int_reg_array_62_31_imag;
        _zz_4559_ = int_reg_array_62_31_real;
      end
      6'b100000 : begin
        _zz_4558_ = int_reg_array_62_32_imag;
        _zz_4559_ = int_reg_array_62_32_real;
      end
      6'b100001 : begin
        _zz_4558_ = int_reg_array_62_33_imag;
        _zz_4559_ = int_reg_array_62_33_real;
      end
      6'b100010 : begin
        _zz_4558_ = int_reg_array_62_34_imag;
        _zz_4559_ = int_reg_array_62_34_real;
      end
      6'b100011 : begin
        _zz_4558_ = int_reg_array_62_35_imag;
        _zz_4559_ = int_reg_array_62_35_real;
      end
      6'b100100 : begin
        _zz_4558_ = int_reg_array_62_36_imag;
        _zz_4559_ = int_reg_array_62_36_real;
      end
      6'b100101 : begin
        _zz_4558_ = int_reg_array_62_37_imag;
        _zz_4559_ = int_reg_array_62_37_real;
      end
      6'b100110 : begin
        _zz_4558_ = int_reg_array_62_38_imag;
        _zz_4559_ = int_reg_array_62_38_real;
      end
      6'b100111 : begin
        _zz_4558_ = int_reg_array_62_39_imag;
        _zz_4559_ = int_reg_array_62_39_real;
      end
      6'b101000 : begin
        _zz_4558_ = int_reg_array_62_40_imag;
        _zz_4559_ = int_reg_array_62_40_real;
      end
      6'b101001 : begin
        _zz_4558_ = int_reg_array_62_41_imag;
        _zz_4559_ = int_reg_array_62_41_real;
      end
      6'b101010 : begin
        _zz_4558_ = int_reg_array_62_42_imag;
        _zz_4559_ = int_reg_array_62_42_real;
      end
      6'b101011 : begin
        _zz_4558_ = int_reg_array_62_43_imag;
        _zz_4559_ = int_reg_array_62_43_real;
      end
      6'b101100 : begin
        _zz_4558_ = int_reg_array_62_44_imag;
        _zz_4559_ = int_reg_array_62_44_real;
      end
      6'b101101 : begin
        _zz_4558_ = int_reg_array_62_45_imag;
        _zz_4559_ = int_reg_array_62_45_real;
      end
      6'b101110 : begin
        _zz_4558_ = int_reg_array_62_46_imag;
        _zz_4559_ = int_reg_array_62_46_real;
      end
      6'b101111 : begin
        _zz_4558_ = int_reg_array_62_47_imag;
        _zz_4559_ = int_reg_array_62_47_real;
      end
      6'b110000 : begin
        _zz_4558_ = int_reg_array_62_48_imag;
        _zz_4559_ = int_reg_array_62_48_real;
      end
      6'b110001 : begin
        _zz_4558_ = int_reg_array_62_49_imag;
        _zz_4559_ = int_reg_array_62_49_real;
      end
      6'b110010 : begin
        _zz_4558_ = int_reg_array_62_50_imag;
        _zz_4559_ = int_reg_array_62_50_real;
      end
      6'b110011 : begin
        _zz_4558_ = int_reg_array_62_51_imag;
        _zz_4559_ = int_reg_array_62_51_real;
      end
      6'b110100 : begin
        _zz_4558_ = int_reg_array_62_52_imag;
        _zz_4559_ = int_reg_array_62_52_real;
      end
      6'b110101 : begin
        _zz_4558_ = int_reg_array_62_53_imag;
        _zz_4559_ = int_reg_array_62_53_real;
      end
      6'b110110 : begin
        _zz_4558_ = int_reg_array_62_54_imag;
        _zz_4559_ = int_reg_array_62_54_real;
      end
      6'b110111 : begin
        _zz_4558_ = int_reg_array_62_55_imag;
        _zz_4559_ = int_reg_array_62_55_real;
      end
      6'b111000 : begin
        _zz_4558_ = int_reg_array_62_56_imag;
        _zz_4559_ = int_reg_array_62_56_real;
      end
      6'b111001 : begin
        _zz_4558_ = int_reg_array_62_57_imag;
        _zz_4559_ = int_reg_array_62_57_real;
      end
      6'b111010 : begin
        _zz_4558_ = int_reg_array_62_58_imag;
        _zz_4559_ = int_reg_array_62_58_real;
      end
      6'b111011 : begin
        _zz_4558_ = int_reg_array_62_59_imag;
        _zz_4559_ = int_reg_array_62_59_real;
      end
      6'b111100 : begin
        _zz_4558_ = int_reg_array_62_60_imag;
        _zz_4559_ = int_reg_array_62_60_real;
      end
      6'b111101 : begin
        _zz_4558_ = int_reg_array_62_61_imag;
        _zz_4559_ = int_reg_array_62_61_real;
      end
      6'b111110 : begin
        _zz_4558_ = int_reg_array_62_62_imag;
        _zz_4559_ = int_reg_array_62_62_real;
      end
      default : begin
        _zz_4558_ = int_reg_array_62_63_imag;
        _zz_4559_ = int_reg_array_62_63_real;
      end
    endcase
  end

  always @(*) begin
    case(_zz_4364_)
      6'b000000 : begin
        _zz_4560_ = int_reg_array_63_0_imag;
        _zz_4561_ = int_reg_array_63_0_real;
      end
      6'b000001 : begin
        _zz_4560_ = int_reg_array_63_1_imag;
        _zz_4561_ = int_reg_array_63_1_real;
      end
      6'b000010 : begin
        _zz_4560_ = int_reg_array_63_2_imag;
        _zz_4561_ = int_reg_array_63_2_real;
      end
      6'b000011 : begin
        _zz_4560_ = int_reg_array_63_3_imag;
        _zz_4561_ = int_reg_array_63_3_real;
      end
      6'b000100 : begin
        _zz_4560_ = int_reg_array_63_4_imag;
        _zz_4561_ = int_reg_array_63_4_real;
      end
      6'b000101 : begin
        _zz_4560_ = int_reg_array_63_5_imag;
        _zz_4561_ = int_reg_array_63_5_real;
      end
      6'b000110 : begin
        _zz_4560_ = int_reg_array_63_6_imag;
        _zz_4561_ = int_reg_array_63_6_real;
      end
      6'b000111 : begin
        _zz_4560_ = int_reg_array_63_7_imag;
        _zz_4561_ = int_reg_array_63_7_real;
      end
      6'b001000 : begin
        _zz_4560_ = int_reg_array_63_8_imag;
        _zz_4561_ = int_reg_array_63_8_real;
      end
      6'b001001 : begin
        _zz_4560_ = int_reg_array_63_9_imag;
        _zz_4561_ = int_reg_array_63_9_real;
      end
      6'b001010 : begin
        _zz_4560_ = int_reg_array_63_10_imag;
        _zz_4561_ = int_reg_array_63_10_real;
      end
      6'b001011 : begin
        _zz_4560_ = int_reg_array_63_11_imag;
        _zz_4561_ = int_reg_array_63_11_real;
      end
      6'b001100 : begin
        _zz_4560_ = int_reg_array_63_12_imag;
        _zz_4561_ = int_reg_array_63_12_real;
      end
      6'b001101 : begin
        _zz_4560_ = int_reg_array_63_13_imag;
        _zz_4561_ = int_reg_array_63_13_real;
      end
      6'b001110 : begin
        _zz_4560_ = int_reg_array_63_14_imag;
        _zz_4561_ = int_reg_array_63_14_real;
      end
      6'b001111 : begin
        _zz_4560_ = int_reg_array_63_15_imag;
        _zz_4561_ = int_reg_array_63_15_real;
      end
      6'b010000 : begin
        _zz_4560_ = int_reg_array_63_16_imag;
        _zz_4561_ = int_reg_array_63_16_real;
      end
      6'b010001 : begin
        _zz_4560_ = int_reg_array_63_17_imag;
        _zz_4561_ = int_reg_array_63_17_real;
      end
      6'b010010 : begin
        _zz_4560_ = int_reg_array_63_18_imag;
        _zz_4561_ = int_reg_array_63_18_real;
      end
      6'b010011 : begin
        _zz_4560_ = int_reg_array_63_19_imag;
        _zz_4561_ = int_reg_array_63_19_real;
      end
      6'b010100 : begin
        _zz_4560_ = int_reg_array_63_20_imag;
        _zz_4561_ = int_reg_array_63_20_real;
      end
      6'b010101 : begin
        _zz_4560_ = int_reg_array_63_21_imag;
        _zz_4561_ = int_reg_array_63_21_real;
      end
      6'b010110 : begin
        _zz_4560_ = int_reg_array_63_22_imag;
        _zz_4561_ = int_reg_array_63_22_real;
      end
      6'b010111 : begin
        _zz_4560_ = int_reg_array_63_23_imag;
        _zz_4561_ = int_reg_array_63_23_real;
      end
      6'b011000 : begin
        _zz_4560_ = int_reg_array_63_24_imag;
        _zz_4561_ = int_reg_array_63_24_real;
      end
      6'b011001 : begin
        _zz_4560_ = int_reg_array_63_25_imag;
        _zz_4561_ = int_reg_array_63_25_real;
      end
      6'b011010 : begin
        _zz_4560_ = int_reg_array_63_26_imag;
        _zz_4561_ = int_reg_array_63_26_real;
      end
      6'b011011 : begin
        _zz_4560_ = int_reg_array_63_27_imag;
        _zz_4561_ = int_reg_array_63_27_real;
      end
      6'b011100 : begin
        _zz_4560_ = int_reg_array_63_28_imag;
        _zz_4561_ = int_reg_array_63_28_real;
      end
      6'b011101 : begin
        _zz_4560_ = int_reg_array_63_29_imag;
        _zz_4561_ = int_reg_array_63_29_real;
      end
      6'b011110 : begin
        _zz_4560_ = int_reg_array_63_30_imag;
        _zz_4561_ = int_reg_array_63_30_real;
      end
      6'b011111 : begin
        _zz_4560_ = int_reg_array_63_31_imag;
        _zz_4561_ = int_reg_array_63_31_real;
      end
      6'b100000 : begin
        _zz_4560_ = int_reg_array_63_32_imag;
        _zz_4561_ = int_reg_array_63_32_real;
      end
      6'b100001 : begin
        _zz_4560_ = int_reg_array_63_33_imag;
        _zz_4561_ = int_reg_array_63_33_real;
      end
      6'b100010 : begin
        _zz_4560_ = int_reg_array_63_34_imag;
        _zz_4561_ = int_reg_array_63_34_real;
      end
      6'b100011 : begin
        _zz_4560_ = int_reg_array_63_35_imag;
        _zz_4561_ = int_reg_array_63_35_real;
      end
      6'b100100 : begin
        _zz_4560_ = int_reg_array_63_36_imag;
        _zz_4561_ = int_reg_array_63_36_real;
      end
      6'b100101 : begin
        _zz_4560_ = int_reg_array_63_37_imag;
        _zz_4561_ = int_reg_array_63_37_real;
      end
      6'b100110 : begin
        _zz_4560_ = int_reg_array_63_38_imag;
        _zz_4561_ = int_reg_array_63_38_real;
      end
      6'b100111 : begin
        _zz_4560_ = int_reg_array_63_39_imag;
        _zz_4561_ = int_reg_array_63_39_real;
      end
      6'b101000 : begin
        _zz_4560_ = int_reg_array_63_40_imag;
        _zz_4561_ = int_reg_array_63_40_real;
      end
      6'b101001 : begin
        _zz_4560_ = int_reg_array_63_41_imag;
        _zz_4561_ = int_reg_array_63_41_real;
      end
      6'b101010 : begin
        _zz_4560_ = int_reg_array_63_42_imag;
        _zz_4561_ = int_reg_array_63_42_real;
      end
      6'b101011 : begin
        _zz_4560_ = int_reg_array_63_43_imag;
        _zz_4561_ = int_reg_array_63_43_real;
      end
      6'b101100 : begin
        _zz_4560_ = int_reg_array_63_44_imag;
        _zz_4561_ = int_reg_array_63_44_real;
      end
      6'b101101 : begin
        _zz_4560_ = int_reg_array_63_45_imag;
        _zz_4561_ = int_reg_array_63_45_real;
      end
      6'b101110 : begin
        _zz_4560_ = int_reg_array_63_46_imag;
        _zz_4561_ = int_reg_array_63_46_real;
      end
      6'b101111 : begin
        _zz_4560_ = int_reg_array_63_47_imag;
        _zz_4561_ = int_reg_array_63_47_real;
      end
      6'b110000 : begin
        _zz_4560_ = int_reg_array_63_48_imag;
        _zz_4561_ = int_reg_array_63_48_real;
      end
      6'b110001 : begin
        _zz_4560_ = int_reg_array_63_49_imag;
        _zz_4561_ = int_reg_array_63_49_real;
      end
      6'b110010 : begin
        _zz_4560_ = int_reg_array_63_50_imag;
        _zz_4561_ = int_reg_array_63_50_real;
      end
      6'b110011 : begin
        _zz_4560_ = int_reg_array_63_51_imag;
        _zz_4561_ = int_reg_array_63_51_real;
      end
      6'b110100 : begin
        _zz_4560_ = int_reg_array_63_52_imag;
        _zz_4561_ = int_reg_array_63_52_real;
      end
      6'b110101 : begin
        _zz_4560_ = int_reg_array_63_53_imag;
        _zz_4561_ = int_reg_array_63_53_real;
      end
      6'b110110 : begin
        _zz_4560_ = int_reg_array_63_54_imag;
        _zz_4561_ = int_reg_array_63_54_real;
      end
      6'b110111 : begin
        _zz_4560_ = int_reg_array_63_55_imag;
        _zz_4561_ = int_reg_array_63_55_real;
      end
      6'b111000 : begin
        _zz_4560_ = int_reg_array_63_56_imag;
        _zz_4561_ = int_reg_array_63_56_real;
      end
      6'b111001 : begin
        _zz_4560_ = int_reg_array_63_57_imag;
        _zz_4561_ = int_reg_array_63_57_real;
      end
      6'b111010 : begin
        _zz_4560_ = int_reg_array_63_58_imag;
        _zz_4561_ = int_reg_array_63_58_real;
      end
      6'b111011 : begin
        _zz_4560_ = int_reg_array_63_59_imag;
        _zz_4561_ = int_reg_array_63_59_real;
      end
      6'b111100 : begin
        _zz_4560_ = int_reg_array_63_60_imag;
        _zz_4561_ = int_reg_array_63_60_real;
      end
      6'b111101 : begin
        _zz_4560_ = int_reg_array_63_61_imag;
        _zz_4561_ = int_reg_array_63_61_real;
      end
      6'b111110 : begin
        _zz_4560_ = int_reg_array_63_62_imag;
        _zz_4561_ = int_reg_array_63_62_real;
      end
      default : begin
        _zz_4560_ = int_reg_array_63_63_imag;
        _zz_4561_ = int_reg_array_63_63_real;
      end
    endcase
  end

  assign _zz_10_ = _zz_7_;
  assign _zz_11_ = _zz_15_;
  assign _zz_12_ = (2'b00);
  assign _zz_2_ = 1'b1;
  assign _zz_8_ = 1'b1;
  assign Axi4Incr_highCat = _zz_13_[31 : 12];
  assign Axi4Incr_sizeValue = 1'b1;
  assign Axi4Incr_alignMask = 12'h0;
  assign Axi4Incr_base = (_zz_4563_ & (~ Axi4Incr_alignMask));
  assign Axi4Incr_baseIncr = (Axi4Incr_base + _zz_4564_);
  always @ (*) begin
    if((((_zz_14_ & 8'h08) == 8'h08))) begin
        _zz_16_ = (2'b11);
    end else if((((_zz_14_ & 8'h04) == 8'h04))) begin
        _zz_16_ = (2'b10);
    end else if((((_zz_14_ & 8'h02) == 8'h02))) begin
        _zz_16_ = (2'b01);
    end else begin
        _zz_16_ = (2'b00);
    end
  end

  assign Axi4Incr_wrapCase = ((2'b00) + _zz_16_);
  always @ (*) begin
    case(_zz_6_)
      2'b00 : begin
        Axi4Incr_result = _zz_13_;
      end
      2'b10 : begin
        Axi4Incr_result = {Axi4Incr_highCat,_zz_4433_};
      end
      default : begin
        Axi4Incr_result = {Axi4Incr_highCat,Axi4Incr_baseIncr};
      end
    endcase
  end

  assign _zz_17_ = _zz_4566_[5:0];
  assign _zz_18_ = ({63'd0,(1'b1)} <<< _zz_17_);
  assign _zz_19_ = _zz_18_[0];
  assign _zz_20_ = _zz_18_[1];
  assign _zz_21_ = _zz_18_[2];
  assign _zz_22_ = _zz_18_[3];
  assign _zz_23_ = _zz_18_[4];
  assign _zz_24_ = _zz_18_[5];
  assign _zz_25_ = _zz_18_[6];
  assign _zz_26_ = _zz_18_[7];
  assign _zz_27_ = _zz_18_[8];
  assign _zz_28_ = _zz_18_[9];
  assign _zz_29_ = _zz_18_[10];
  assign _zz_30_ = _zz_18_[11];
  assign _zz_31_ = _zz_18_[12];
  assign _zz_32_ = _zz_18_[13];
  assign _zz_33_ = _zz_18_[14];
  assign _zz_34_ = _zz_18_[15];
  assign _zz_35_ = _zz_18_[16];
  assign _zz_36_ = _zz_18_[17];
  assign _zz_37_ = _zz_18_[18];
  assign _zz_38_ = _zz_18_[19];
  assign _zz_39_ = _zz_18_[20];
  assign _zz_40_ = _zz_18_[21];
  assign _zz_41_ = _zz_18_[22];
  assign _zz_42_ = _zz_18_[23];
  assign _zz_43_ = _zz_18_[24];
  assign _zz_44_ = _zz_18_[25];
  assign _zz_45_ = _zz_18_[26];
  assign _zz_46_ = _zz_18_[27];
  assign _zz_47_ = _zz_18_[28];
  assign _zz_48_ = _zz_18_[29];
  assign _zz_49_ = _zz_18_[30];
  assign _zz_50_ = _zz_18_[31];
  assign _zz_51_ = _zz_18_[32];
  assign _zz_52_ = _zz_18_[33];
  assign _zz_53_ = _zz_18_[34];
  assign _zz_54_ = _zz_18_[35];
  assign _zz_55_ = _zz_18_[36];
  assign _zz_56_ = _zz_18_[37];
  assign _zz_57_ = _zz_18_[38];
  assign _zz_58_ = _zz_18_[39];
  assign _zz_59_ = _zz_18_[40];
  assign _zz_60_ = _zz_18_[41];
  assign _zz_61_ = _zz_18_[42];
  assign _zz_62_ = _zz_18_[43];
  assign _zz_63_ = _zz_18_[44];
  assign _zz_64_ = _zz_18_[45];
  assign _zz_65_ = _zz_18_[46];
  assign _zz_66_ = _zz_18_[47];
  assign _zz_67_ = _zz_18_[48];
  assign _zz_68_ = _zz_18_[49];
  assign _zz_69_ = _zz_18_[50];
  assign _zz_70_ = _zz_18_[51];
  assign _zz_71_ = _zz_18_[52];
  assign _zz_72_ = _zz_18_[53];
  assign _zz_73_ = _zz_18_[54];
  assign _zz_74_ = _zz_18_[55];
  assign _zz_75_ = _zz_18_[56];
  assign _zz_76_ = _zz_18_[57];
  assign _zz_77_ = _zz_18_[58];
  assign _zz_78_ = _zz_18_[59];
  assign _zz_79_ = _zz_18_[60];
  assign _zz_80_ = _zz_18_[61];
  assign _zz_81_ = _zz_18_[62];
  assign _zz_82_ = _zz_18_[63];
  assign _zz_83_ = (((32'h0 <= load_data_area_current_addr) && (load_data_area_current_addr < 32'h00000040)) ? _zz_9__regNext : {_zz_4434_,_zz_4435_});
  assign _zz_84_ = _zz_83_[15 : 0];
  assign _zz_85_ = _zz_83_[31 : 16];
  assign _zz_86_ = _zz_4567_[5:0];
  assign _zz_87_ = ({63'd0,(1'b1)} <<< _zz_86_);
  assign _zz_88_ = _zz_87_[0];
  assign _zz_89_ = _zz_87_[1];
  assign _zz_90_ = _zz_87_[2];
  assign _zz_91_ = _zz_87_[3];
  assign _zz_92_ = _zz_87_[4];
  assign _zz_93_ = _zz_87_[5];
  assign _zz_94_ = _zz_87_[6];
  assign _zz_95_ = _zz_87_[7];
  assign _zz_96_ = _zz_87_[8];
  assign _zz_97_ = _zz_87_[9];
  assign _zz_98_ = _zz_87_[10];
  assign _zz_99_ = _zz_87_[11];
  assign _zz_100_ = _zz_87_[12];
  assign _zz_101_ = _zz_87_[13];
  assign _zz_102_ = _zz_87_[14];
  assign _zz_103_ = _zz_87_[15];
  assign _zz_104_ = _zz_87_[16];
  assign _zz_105_ = _zz_87_[17];
  assign _zz_106_ = _zz_87_[18];
  assign _zz_107_ = _zz_87_[19];
  assign _zz_108_ = _zz_87_[20];
  assign _zz_109_ = _zz_87_[21];
  assign _zz_110_ = _zz_87_[22];
  assign _zz_111_ = _zz_87_[23];
  assign _zz_112_ = _zz_87_[24];
  assign _zz_113_ = _zz_87_[25];
  assign _zz_114_ = _zz_87_[26];
  assign _zz_115_ = _zz_87_[27];
  assign _zz_116_ = _zz_87_[28];
  assign _zz_117_ = _zz_87_[29];
  assign _zz_118_ = _zz_87_[30];
  assign _zz_119_ = _zz_87_[31];
  assign _zz_120_ = _zz_87_[32];
  assign _zz_121_ = _zz_87_[33];
  assign _zz_122_ = _zz_87_[34];
  assign _zz_123_ = _zz_87_[35];
  assign _zz_124_ = _zz_87_[36];
  assign _zz_125_ = _zz_87_[37];
  assign _zz_126_ = _zz_87_[38];
  assign _zz_127_ = _zz_87_[39];
  assign _zz_128_ = _zz_87_[40];
  assign _zz_129_ = _zz_87_[41];
  assign _zz_130_ = _zz_87_[42];
  assign _zz_131_ = _zz_87_[43];
  assign _zz_132_ = _zz_87_[44];
  assign _zz_133_ = _zz_87_[45];
  assign _zz_134_ = _zz_87_[46];
  assign _zz_135_ = _zz_87_[47];
  assign _zz_136_ = _zz_87_[48];
  assign _zz_137_ = _zz_87_[49];
  assign _zz_138_ = _zz_87_[50];
  assign _zz_139_ = _zz_87_[51];
  assign _zz_140_ = _zz_87_[52];
  assign _zz_141_ = _zz_87_[53];
  assign _zz_142_ = _zz_87_[54];
  assign _zz_143_ = _zz_87_[55];
  assign _zz_144_ = _zz_87_[56];
  assign _zz_145_ = _zz_87_[57];
  assign _zz_146_ = _zz_87_[58];
  assign _zz_147_ = _zz_87_[59];
  assign _zz_148_ = _zz_87_[60];
  assign _zz_149_ = _zz_87_[61];
  assign _zz_150_ = _zz_87_[62];
  assign _zz_151_ = _zz_87_[63];
  assign _zz_152_ = (((32'h00000f00 <= load_data_area_current_addr) && (load_data_area_current_addr < 32'h00000f40)) ? _zz_9__regNext : {_zz_4436_,_zz_4437_});
  assign _zz_153_ = _zz_152_[15 : 0];
  assign _zz_154_ = _zz_152_[31 : 16];
  assign _zz_155_ = _zz_4568_[5:0];
  assign _zz_156_ = ({63'd0,(1'b1)} <<< _zz_155_);
  assign _zz_157_ = _zz_156_[0];
  assign _zz_158_ = _zz_156_[1];
  assign _zz_159_ = _zz_156_[2];
  assign _zz_160_ = _zz_156_[3];
  assign _zz_161_ = _zz_156_[4];
  assign _zz_162_ = _zz_156_[5];
  assign _zz_163_ = _zz_156_[6];
  assign _zz_164_ = _zz_156_[7];
  assign _zz_165_ = _zz_156_[8];
  assign _zz_166_ = _zz_156_[9];
  assign _zz_167_ = _zz_156_[10];
  assign _zz_168_ = _zz_156_[11];
  assign _zz_169_ = _zz_156_[12];
  assign _zz_170_ = _zz_156_[13];
  assign _zz_171_ = _zz_156_[14];
  assign _zz_172_ = _zz_156_[15];
  assign _zz_173_ = _zz_156_[16];
  assign _zz_174_ = _zz_156_[17];
  assign _zz_175_ = _zz_156_[18];
  assign _zz_176_ = _zz_156_[19];
  assign _zz_177_ = _zz_156_[20];
  assign _zz_178_ = _zz_156_[21];
  assign _zz_179_ = _zz_156_[22];
  assign _zz_180_ = _zz_156_[23];
  assign _zz_181_ = _zz_156_[24];
  assign _zz_182_ = _zz_156_[25];
  assign _zz_183_ = _zz_156_[26];
  assign _zz_184_ = _zz_156_[27];
  assign _zz_185_ = _zz_156_[28];
  assign _zz_186_ = _zz_156_[29];
  assign _zz_187_ = _zz_156_[30];
  assign _zz_188_ = _zz_156_[31];
  assign _zz_189_ = _zz_156_[32];
  assign _zz_190_ = _zz_156_[33];
  assign _zz_191_ = _zz_156_[34];
  assign _zz_192_ = _zz_156_[35];
  assign _zz_193_ = _zz_156_[36];
  assign _zz_194_ = _zz_156_[37];
  assign _zz_195_ = _zz_156_[38];
  assign _zz_196_ = _zz_156_[39];
  assign _zz_197_ = _zz_156_[40];
  assign _zz_198_ = _zz_156_[41];
  assign _zz_199_ = _zz_156_[42];
  assign _zz_200_ = _zz_156_[43];
  assign _zz_201_ = _zz_156_[44];
  assign _zz_202_ = _zz_156_[45];
  assign _zz_203_ = _zz_156_[46];
  assign _zz_204_ = _zz_156_[47];
  assign _zz_205_ = _zz_156_[48];
  assign _zz_206_ = _zz_156_[49];
  assign _zz_207_ = _zz_156_[50];
  assign _zz_208_ = _zz_156_[51];
  assign _zz_209_ = _zz_156_[52];
  assign _zz_210_ = _zz_156_[53];
  assign _zz_211_ = _zz_156_[54];
  assign _zz_212_ = _zz_156_[55];
  assign _zz_213_ = _zz_156_[56];
  assign _zz_214_ = _zz_156_[57];
  assign _zz_215_ = _zz_156_[58];
  assign _zz_216_ = _zz_156_[59];
  assign _zz_217_ = _zz_156_[60];
  assign _zz_218_ = _zz_156_[61];
  assign _zz_219_ = _zz_156_[62];
  assign _zz_220_ = _zz_156_[63];
  assign _zz_221_ = (((32'h00000b80 <= load_data_area_current_addr) && (load_data_area_current_addr < 32'h00000bc0)) ? _zz_9__regNext : {_zz_4438_,_zz_4439_});
  assign _zz_222_ = _zz_221_[15 : 0];
  assign _zz_223_ = _zz_221_[31 : 16];
  assign _zz_224_ = _zz_4569_[5:0];
  assign _zz_225_ = ({63'd0,(1'b1)} <<< _zz_224_);
  assign _zz_226_ = _zz_225_[0];
  assign _zz_227_ = _zz_225_[1];
  assign _zz_228_ = _zz_225_[2];
  assign _zz_229_ = _zz_225_[3];
  assign _zz_230_ = _zz_225_[4];
  assign _zz_231_ = _zz_225_[5];
  assign _zz_232_ = _zz_225_[6];
  assign _zz_233_ = _zz_225_[7];
  assign _zz_234_ = _zz_225_[8];
  assign _zz_235_ = _zz_225_[9];
  assign _zz_236_ = _zz_225_[10];
  assign _zz_237_ = _zz_225_[11];
  assign _zz_238_ = _zz_225_[12];
  assign _zz_239_ = _zz_225_[13];
  assign _zz_240_ = _zz_225_[14];
  assign _zz_241_ = _zz_225_[15];
  assign _zz_242_ = _zz_225_[16];
  assign _zz_243_ = _zz_225_[17];
  assign _zz_244_ = _zz_225_[18];
  assign _zz_245_ = _zz_225_[19];
  assign _zz_246_ = _zz_225_[20];
  assign _zz_247_ = _zz_225_[21];
  assign _zz_248_ = _zz_225_[22];
  assign _zz_249_ = _zz_225_[23];
  assign _zz_250_ = _zz_225_[24];
  assign _zz_251_ = _zz_225_[25];
  assign _zz_252_ = _zz_225_[26];
  assign _zz_253_ = _zz_225_[27];
  assign _zz_254_ = _zz_225_[28];
  assign _zz_255_ = _zz_225_[29];
  assign _zz_256_ = _zz_225_[30];
  assign _zz_257_ = _zz_225_[31];
  assign _zz_258_ = _zz_225_[32];
  assign _zz_259_ = _zz_225_[33];
  assign _zz_260_ = _zz_225_[34];
  assign _zz_261_ = _zz_225_[35];
  assign _zz_262_ = _zz_225_[36];
  assign _zz_263_ = _zz_225_[37];
  assign _zz_264_ = _zz_225_[38];
  assign _zz_265_ = _zz_225_[39];
  assign _zz_266_ = _zz_225_[40];
  assign _zz_267_ = _zz_225_[41];
  assign _zz_268_ = _zz_225_[42];
  assign _zz_269_ = _zz_225_[43];
  assign _zz_270_ = _zz_225_[44];
  assign _zz_271_ = _zz_225_[45];
  assign _zz_272_ = _zz_225_[46];
  assign _zz_273_ = _zz_225_[47];
  assign _zz_274_ = _zz_225_[48];
  assign _zz_275_ = _zz_225_[49];
  assign _zz_276_ = _zz_225_[50];
  assign _zz_277_ = _zz_225_[51];
  assign _zz_278_ = _zz_225_[52];
  assign _zz_279_ = _zz_225_[53];
  assign _zz_280_ = _zz_225_[54];
  assign _zz_281_ = _zz_225_[55];
  assign _zz_282_ = _zz_225_[56];
  assign _zz_283_ = _zz_225_[57];
  assign _zz_284_ = _zz_225_[58];
  assign _zz_285_ = _zz_225_[59];
  assign _zz_286_ = _zz_225_[60];
  assign _zz_287_ = _zz_225_[61];
  assign _zz_288_ = _zz_225_[62];
  assign _zz_289_ = _zz_225_[63];
  assign _zz_290_ = (((32'h000009c0 <= load_data_area_current_addr) && (load_data_area_current_addr < 32'h00000a00)) ? _zz_9__regNext : {_zz_4440_,_zz_4441_});
  assign _zz_291_ = _zz_290_[15 : 0];
  assign _zz_292_ = _zz_290_[31 : 16];
  assign _zz_293_ = _zz_4570_[5:0];
  assign _zz_294_ = ({63'd0,(1'b1)} <<< _zz_293_);
  assign _zz_295_ = _zz_294_[0];
  assign _zz_296_ = _zz_294_[1];
  assign _zz_297_ = _zz_294_[2];
  assign _zz_298_ = _zz_294_[3];
  assign _zz_299_ = _zz_294_[4];
  assign _zz_300_ = _zz_294_[5];
  assign _zz_301_ = _zz_294_[6];
  assign _zz_302_ = _zz_294_[7];
  assign _zz_303_ = _zz_294_[8];
  assign _zz_304_ = _zz_294_[9];
  assign _zz_305_ = _zz_294_[10];
  assign _zz_306_ = _zz_294_[11];
  assign _zz_307_ = _zz_294_[12];
  assign _zz_308_ = _zz_294_[13];
  assign _zz_309_ = _zz_294_[14];
  assign _zz_310_ = _zz_294_[15];
  assign _zz_311_ = _zz_294_[16];
  assign _zz_312_ = _zz_294_[17];
  assign _zz_313_ = _zz_294_[18];
  assign _zz_314_ = _zz_294_[19];
  assign _zz_315_ = _zz_294_[20];
  assign _zz_316_ = _zz_294_[21];
  assign _zz_317_ = _zz_294_[22];
  assign _zz_318_ = _zz_294_[23];
  assign _zz_319_ = _zz_294_[24];
  assign _zz_320_ = _zz_294_[25];
  assign _zz_321_ = _zz_294_[26];
  assign _zz_322_ = _zz_294_[27];
  assign _zz_323_ = _zz_294_[28];
  assign _zz_324_ = _zz_294_[29];
  assign _zz_325_ = _zz_294_[30];
  assign _zz_326_ = _zz_294_[31];
  assign _zz_327_ = _zz_294_[32];
  assign _zz_328_ = _zz_294_[33];
  assign _zz_329_ = _zz_294_[34];
  assign _zz_330_ = _zz_294_[35];
  assign _zz_331_ = _zz_294_[36];
  assign _zz_332_ = _zz_294_[37];
  assign _zz_333_ = _zz_294_[38];
  assign _zz_334_ = _zz_294_[39];
  assign _zz_335_ = _zz_294_[40];
  assign _zz_336_ = _zz_294_[41];
  assign _zz_337_ = _zz_294_[42];
  assign _zz_338_ = _zz_294_[43];
  assign _zz_339_ = _zz_294_[44];
  assign _zz_340_ = _zz_294_[45];
  assign _zz_341_ = _zz_294_[46];
  assign _zz_342_ = _zz_294_[47];
  assign _zz_343_ = _zz_294_[48];
  assign _zz_344_ = _zz_294_[49];
  assign _zz_345_ = _zz_294_[50];
  assign _zz_346_ = _zz_294_[51];
  assign _zz_347_ = _zz_294_[52];
  assign _zz_348_ = _zz_294_[53];
  assign _zz_349_ = _zz_294_[54];
  assign _zz_350_ = _zz_294_[55];
  assign _zz_351_ = _zz_294_[56];
  assign _zz_352_ = _zz_294_[57];
  assign _zz_353_ = _zz_294_[58];
  assign _zz_354_ = _zz_294_[59];
  assign _zz_355_ = _zz_294_[60];
  assign _zz_356_ = _zz_294_[61];
  assign _zz_357_ = _zz_294_[62];
  assign _zz_358_ = _zz_294_[63];
  assign _zz_359_ = (((32'h00000b00 <= load_data_area_current_addr) && (load_data_area_current_addr < 32'h00000b40)) ? _zz_9__regNext : {_zz_4442_,_zz_4443_});
  assign _zz_360_ = _zz_359_[15 : 0];
  assign _zz_361_ = _zz_359_[31 : 16];
  assign _zz_362_ = _zz_4571_[5:0];
  assign _zz_363_ = ({63'd0,(1'b1)} <<< _zz_362_);
  assign _zz_364_ = _zz_363_[0];
  assign _zz_365_ = _zz_363_[1];
  assign _zz_366_ = _zz_363_[2];
  assign _zz_367_ = _zz_363_[3];
  assign _zz_368_ = _zz_363_[4];
  assign _zz_369_ = _zz_363_[5];
  assign _zz_370_ = _zz_363_[6];
  assign _zz_371_ = _zz_363_[7];
  assign _zz_372_ = _zz_363_[8];
  assign _zz_373_ = _zz_363_[9];
  assign _zz_374_ = _zz_363_[10];
  assign _zz_375_ = _zz_363_[11];
  assign _zz_376_ = _zz_363_[12];
  assign _zz_377_ = _zz_363_[13];
  assign _zz_378_ = _zz_363_[14];
  assign _zz_379_ = _zz_363_[15];
  assign _zz_380_ = _zz_363_[16];
  assign _zz_381_ = _zz_363_[17];
  assign _zz_382_ = _zz_363_[18];
  assign _zz_383_ = _zz_363_[19];
  assign _zz_384_ = _zz_363_[20];
  assign _zz_385_ = _zz_363_[21];
  assign _zz_386_ = _zz_363_[22];
  assign _zz_387_ = _zz_363_[23];
  assign _zz_388_ = _zz_363_[24];
  assign _zz_389_ = _zz_363_[25];
  assign _zz_390_ = _zz_363_[26];
  assign _zz_391_ = _zz_363_[27];
  assign _zz_392_ = _zz_363_[28];
  assign _zz_393_ = _zz_363_[29];
  assign _zz_394_ = _zz_363_[30];
  assign _zz_395_ = _zz_363_[31];
  assign _zz_396_ = _zz_363_[32];
  assign _zz_397_ = _zz_363_[33];
  assign _zz_398_ = _zz_363_[34];
  assign _zz_399_ = _zz_363_[35];
  assign _zz_400_ = _zz_363_[36];
  assign _zz_401_ = _zz_363_[37];
  assign _zz_402_ = _zz_363_[38];
  assign _zz_403_ = _zz_363_[39];
  assign _zz_404_ = _zz_363_[40];
  assign _zz_405_ = _zz_363_[41];
  assign _zz_406_ = _zz_363_[42];
  assign _zz_407_ = _zz_363_[43];
  assign _zz_408_ = _zz_363_[44];
  assign _zz_409_ = _zz_363_[45];
  assign _zz_410_ = _zz_363_[46];
  assign _zz_411_ = _zz_363_[47];
  assign _zz_412_ = _zz_363_[48];
  assign _zz_413_ = _zz_363_[49];
  assign _zz_414_ = _zz_363_[50];
  assign _zz_415_ = _zz_363_[51];
  assign _zz_416_ = _zz_363_[52];
  assign _zz_417_ = _zz_363_[53];
  assign _zz_418_ = _zz_363_[54];
  assign _zz_419_ = _zz_363_[55];
  assign _zz_420_ = _zz_363_[56];
  assign _zz_421_ = _zz_363_[57];
  assign _zz_422_ = _zz_363_[58];
  assign _zz_423_ = _zz_363_[59];
  assign _zz_424_ = _zz_363_[60];
  assign _zz_425_ = _zz_363_[61];
  assign _zz_426_ = _zz_363_[62];
  assign _zz_427_ = _zz_363_[63];
  assign _zz_428_ = (((32'h000005c0 <= load_data_area_current_addr) && (load_data_area_current_addr < 32'h00000600)) ? _zz_9__regNext : {_zz_4444_,_zz_4445_});
  assign _zz_429_ = _zz_428_[15 : 0];
  assign _zz_430_ = _zz_428_[31 : 16];
  assign _zz_431_ = _zz_4572_[5:0];
  assign _zz_432_ = ({63'd0,(1'b1)} <<< _zz_431_);
  assign _zz_433_ = _zz_432_[0];
  assign _zz_434_ = _zz_432_[1];
  assign _zz_435_ = _zz_432_[2];
  assign _zz_436_ = _zz_432_[3];
  assign _zz_437_ = _zz_432_[4];
  assign _zz_438_ = _zz_432_[5];
  assign _zz_439_ = _zz_432_[6];
  assign _zz_440_ = _zz_432_[7];
  assign _zz_441_ = _zz_432_[8];
  assign _zz_442_ = _zz_432_[9];
  assign _zz_443_ = _zz_432_[10];
  assign _zz_444_ = _zz_432_[11];
  assign _zz_445_ = _zz_432_[12];
  assign _zz_446_ = _zz_432_[13];
  assign _zz_447_ = _zz_432_[14];
  assign _zz_448_ = _zz_432_[15];
  assign _zz_449_ = _zz_432_[16];
  assign _zz_450_ = _zz_432_[17];
  assign _zz_451_ = _zz_432_[18];
  assign _zz_452_ = _zz_432_[19];
  assign _zz_453_ = _zz_432_[20];
  assign _zz_454_ = _zz_432_[21];
  assign _zz_455_ = _zz_432_[22];
  assign _zz_456_ = _zz_432_[23];
  assign _zz_457_ = _zz_432_[24];
  assign _zz_458_ = _zz_432_[25];
  assign _zz_459_ = _zz_432_[26];
  assign _zz_460_ = _zz_432_[27];
  assign _zz_461_ = _zz_432_[28];
  assign _zz_462_ = _zz_432_[29];
  assign _zz_463_ = _zz_432_[30];
  assign _zz_464_ = _zz_432_[31];
  assign _zz_465_ = _zz_432_[32];
  assign _zz_466_ = _zz_432_[33];
  assign _zz_467_ = _zz_432_[34];
  assign _zz_468_ = _zz_432_[35];
  assign _zz_469_ = _zz_432_[36];
  assign _zz_470_ = _zz_432_[37];
  assign _zz_471_ = _zz_432_[38];
  assign _zz_472_ = _zz_432_[39];
  assign _zz_473_ = _zz_432_[40];
  assign _zz_474_ = _zz_432_[41];
  assign _zz_475_ = _zz_432_[42];
  assign _zz_476_ = _zz_432_[43];
  assign _zz_477_ = _zz_432_[44];
  assign _zz_478_ = _zz_432_[45];
  assign _zz_479_ = _zz_432_[46];
  assign _zz_480_ = _zz_432_[47];
  assign _zz_481_ = _zz_432_[48];
  assign _zz_482_ = _zz_432_[49];
  assign _zz_483_ = _zz_432_[50];
  assign _zz_484_ = _zz_432_[51];
  assign _zz_485_ = _zz_432_[52];
  assign _zz_486_ = _zz_432_[53];
  assign _zz_487_ = _zz_432_[54];
  assign _zz_488_ = _zz_432_[55];
  assign _zz_489_ = _zz_432_[56];
  assign _zz_490_ = _zz_432_[57];
  assign _zz_491_ = _zz_432_[58];
  assign _zz_492_ = _zz_432_[59];
  assign _zz_493_ = _zz_432_[60];
  assign _zz_494_ = _zz_432_[61];
  assign _zz_495_ = _zz_432_[62];
  assign _zz_496_ = _zz_432_[63];
  assign _zz_497_ = (((32'h00000c80 <= load_data_area_current_addr) && (load_data_area_current_addr < 32'h00000cc0)) ? _zz_9__regNext : {_zz_4446_,_zz_4447_});
  assign _zz_498_ = _zz_497_[15 : 0];
  assign _zz_499_ = _zz_497_[31 : 16];
  assign _zz_500_ = _zz_4573_[5:0];
  assign _zz_501_ = ({63'd0,(1'b1)} <<< _zz_500_);
  assign _zz_502_ = _zz_501_[0];
  assign _zz_503_ = _zz_501_[1];
  assign _zz_504_ = _zz_501_[2];
  assign _zz_505_ = _zz_501_[3];
  assign _zz_506_ = _zz_501_[4];
  assign _zz_507_ = _zz_501_[5];
  assign _zz_508_ = _zz_501_[6];
  assign _zz_509_ = _zz_501_[7];
  assign _zz_510_ = _zz_501_[8];
  assign _zz_511_ = _zz_501_[9];
  assign _zz_512_ = _zz_501_[10];
  assign _zz_513_ = _zz_501_[11];
  assign _zz_514_ = _zz_501_[12];
  assign _zz_515_ = _zz_501_[13];
  assign _zz_516_ = _zz_501_[14];
  assign _zz_517_ = _zz_501_[15];
  assign _zz_518_ = _zz_501_[16];
  assign _zz_519_ = _zz_501_[17];
  assign _zz_520_ = _zz_501_[18];
  assign _zz_521_ = _zz_501_[19];
  assign _zz_522_ = _zz_501_[20];
  assign _zz_523_ = _zz_501_[21];
  assign _zz_524_ = _zz_501_[22];
  assign _zz_525_ = _zz_501_[23];
  assign _zz_526_ = _zz_501_[24];
  assign _zz_527_ = _zz_501_[25];
  assign _zz_528_ = _zz_501_[26];
  assign _zz_529_ = _zz_501_[27];
  assign _zz_530_ = _zz_501_[28];
  assign _zz_531_ = _zz_501_[29];
  assign _zz_532_ = _zz_501_[30];
  assign _zz_533_ = _zz_501_[31];
  assign _zz_534_ = _zz_501_[32];
  assign _zz_535_ = _zz_501_[33];
  assign _zz_536_ = _zz_501_[34];
  assign _zz_537_ = _zz_501_[35];
  assign _zz_538_ = _zz_501_[36];
  assign _zz_539_ = _zz_501_[37];
  assign _zz_540_ = _zz_501_[38];
  assign _zz_541_ = _zz_501_[39];
  assign _zz_542_ = _zz_501_[40];
  assign _zz_543_ = _zz_501_[41];
  assign _zz_544_ = _zz_501_[42];
  assign _zz_545_ = _zz_501_[43];
  assign _zz_546_ = _zz_501_[44];
  assign _zz_547_ = _zz_501_[45];
  assign _zz_548_ = _zz_501_[46];
  assign _zz_549_ = _zz_501_[47];
  assign _zz_550_ = _zz_501_[48];
  assign _zz_551_ = _zz_501_[49];
  assign _zz_552_ = _zz_501_[50];
  assign _zz_553_ = _zz_501_[51];
  assign _zz_554_ = _zz_501_[52];
  assign _zz_555_ = _zz_501_[53];
  assign _zz_556_ = _zz_501_[54];
  assign _zz_557_ = _zz_501_[55];
  assign _zz_558_ = _zz_501_[56];
  assign _zz_559_ = _zz_501_[57];
  assign _zz_560_ = _zz_501_[58];
  assign _zz_561_ = _zz_501_[59];
  assign _zz_562_ = _zz_501_[60];
  assign _zz_563_ = _zz_501_[61];
  assign _zz_564_ = _zz_501_[62];
  assign _zz_565_ = _zz_501_[63];
  assign _zz_566_ = (((32'h00000a40 <= load_data_area_current_addr) && (load_data_area_current_addr < 32'h00000a80)) ? _zz_9__regNext : {_zz_4448_,_zz_4449_});
  assign _zz_567_ = _zz_566_[15 : 0];
  assign _zz_568_ = _zz_566_[31 : 16];
  assign _zz_569_ = _zz_4574_[5:0];
  assign _zz_570_ = ({63'd0,(1'b1)} <<< _zz_569_);
  assign _zz_571_ = _zz_570_[0];
  assign _zz_572_ = _zz_570_[1];
  assign _zz_573_ = _zz_570_[2];
  assign _zz_574_ = _zz_570_[3];
  assign _zz_575_ = _zz_570_[4];
  assign _zz_576_ = _zz_570_[5];
  assign _zz_577_ = _zz_570_[6];
  assign _zz_578_ = _zz_570_[7];
  assign _zz_579_ = _zz_570_[8];
  assign _zz_580_ = _zz_570_[9];
  assign _zz_581_ = _zz_570_[10];
  assign _zz_582_ = _zz_570_[11];
  assign _zz_583_ = _zz_570_[12];
  assign _zz_584_ = _zz_570_[13];
  assign _zz_585_ = _zz_570_[14];
  assign _zz_586_ = _zz_570_[15];
  assign _zz_587_ = _zz_570_[16];
  assign _zz_588_ = _zz_570_[17];
  assign _zz_589_ = _zz_570_[18];
  assign _zz_590_ = _zz_570_[19];
  assign _zz_591_ = _zz_570_[20];
  assign _zz_592_ = _zz_570_[21];
  assign _zz_593_ = _zz_570_[22];
  assign _zz_594_ = _zz_570_[23];
  assign _zz_595_ = _zz_570_[24];
  assign _zz_596_ = _zz_570_[25];
  assign _zz_597_ = _zz_570_[26];
  assign _zz_598_ = _zz_570_[27];
  assign _zz_599_ = _zz_570_[28];
  assign _zz_600_ = _zz_570_[29];
  assign _zz_601_ = _zz_570_[30];
  assign _zz_602_ = _zz_570_[31];
  assign _zz_603_ = _zz_570_[32];
  assign _zz_604_ = _zz_570_[33];
  assign _zz_605_ = _zz_570_[34];
  assign _zz_606_ = _zz_570_[35];
  assign _zz_607_ = _zz_570_[36];
  assign _zz_608_ = _zz_570_[37];
  assign _zz_609_ = _zz_570_[38];
  assign _zz_610_ = _zz_570_[39];
  assign _zz_611_ = _zz_570_[40];
  assign _zz_612_ = _zz_570_[41];
  assign _zz_613_ = _zz_570_[42];
  assign _zz_614_ = _zz_570_[43];
  assign _zz_615_ = _zz_570_[44];
  assign _zz_616_ = _zz_570_[45];
  assign _zz_617_ = _zz_570_[46];
  assign _zz_618_ = _zz_570_[47];
  assign _zz_619_ = _zz_570_[48];
  assign _zz_620_ = _zz_570_[49];
  assign _zz_621_ = _zz_570_[50];
  assign _zz_622_ = _zz_570_[51];
  assign _zz_623_ = _zz_570_[52];
  assign _zz_624_ = _zz_570_[53];
  assign _zz_625_ = _zz_570_[54];
  assign _zz_626_ = _zz_570_[55];
  assign _zz_627_ = _zz_570_[56];
  assign _zz_628_ = _zz_570_[57];
  assign _zz_629_ = _zz_570_[58];
  assign _zz_630_ = _zz_570_[59];
  assign _zz_631_ = _zz_570_[60];
  assign _zz_632_ = _zz_570_[61];
  assign _zz_633_ = _zz_570_[62];
  assign _zz_634_ = _zz_570_[63];
  assign _zz_635_ = (((32'h000002c0 <= load_data_area_current_addr) && (load_data_area_current_addr < 32'h00000300)) ? _zz_9__regNext : {_zz_4450_,_zz_4451_});
  assign _zz_636_ = _zz_635_[15 : 0];
  assign _zz_637_ = _zz_635_[31 : 16];
  assign _zz_638_ = _zz_4575_[5:0];
  assign _zz_639_ = ({63'd0,(1'b1)} <<< _zz_638_);
  assign _zz_640_ = _zz_639_[0];
  assign _zz_641_ = _zz_639_[1];
  assign _zz_642_ = _zz_639_[2];
  assign _zz_643_ = _zz_639_[3];
  assign _zz_644_ = _zz_639_[4];
  assign _zz_645_ = _zz_639_[5];
  assign _zz_646_ = _zz_639_[6];
  assign _zz_647_ = _zz_639_[7];
  assign _zz_648_ = _zz_639_[8];
  assign _zz_649_ = _zz_639_[9];
  assign _zz_650_ = _zz_639_[10];
  assign _zz_651_ = _zz_639_[11];
  assign _zz_652_ = _zz_639_[12];
  assign _zz_653_ = _zz_639_[13];
  assign _zz_654_ = _zz_639_[14];
  assign _zz_655_ = _zz_639_[15];
  assign _zz_656_ = _zz_639_[16];
  assign _zz_657_ = _zz_639_[17];
  assign _zz_658_ = _zz_639_[18];
  assign _zz_659_ = _zz_639_[19];
  assign _zz_660_ = _zz_639_[20];
  assign _zz_661_ = _zz_639_[21];
  assign _zz_662_ = _zz_639_[22];
  assign _zz_663_ = _zz_639_[23];
  assign _zz_664_ = _zz_639_[24];
  assign _zz_665_ = _zz_639_[25];
  assign _zz_666_ = _zz_639_[26];
  assign _zz_667_ = _zz_639_[27];
  assign _zz_668_ = _zz_639_[28];
  assign _zz_669_ = _zz_639_[29];
  assign _zz_670_ = _zz_639_[30];
  assign _zz_671_ = _zz_639_[31];
  assign _zz_672_ = _zz_639_[32];
  assign _zz_673_ = _zz_639_[33];
  assign _zz_674_ = _zz_639_[34];
  assign _zz_675_ = _zz_639_[35];
  assign _zz_676_ = _zz_639_[36];
  assign _zz_677_ = _zz_639_[37];
  assign _zz_678_ = _zz_639_[38];
  assign _zz_679_ = _zz_639_[39];
  assign _zz_680_ = _zz_639_[40];
  assign _zz_681_ = _zz_639_[41];
  assign _zz_682_ = _zz_639_[42];
  assign _zz_683_ = _zz_639_[43];
  assign _zz_684_ = _zz_639_[44];
  assign _zz_685_ = _zz_639_[45];
  assign _zz_686_ = _zz_639_[46];
  assign _zz_687_ = _zz_639_[47];
  assign _zz_688_ = _zz_639_[48];
  assign _zz_689_ = _zz_639_[49];
  assign _zz_690_ = _zz_639_[50];
  assign _zz_691_ = _zz_639_[51];
  assign _zz_692_ = _zz_639_[52];
  assign _zz_693_ = _zz_639_[53];
  assign _zz_694_ = _zz_639_[54];
  assign _zz_695_ = _zz_639_[55];
  assign _zz_696_ = _zz_639_[56];
  assign _zz_697_ = _zz_639_[57];
  assign _zz_698_ = _zz_639_[58];
  assign _zz_699_ = _zz_639_[59];
  assign _zz_700_ = _zz_639_[60];
  assign _zz_701_ = _zz_639_[61];
  assign _zz_702_ = _zz_639_[62];
  assign _zz_703_ = _zz_639_[63];
  assign _zz_704_ = (((32'h00000f80 <= load_data_area_current_addr) && (load_data_area_current_addr < 32'h00000fc0)) ? _zz_9__regNext : {_zz_4452_,_zz_4453_});
  assign _zz_705_ = _zz_704_[15 : 0];
  assign _zz_706_ = _zz_704_[31 : 16];
  assign _zz_707_ = _zz_4576_[5:0];
  assign _zz_708_ = ({63'd0,(1'b1)} <<< _zz_707_);
  assign _zz_709_ = _zz_708_[0];
  assign _zz_710_ = _zz_708_[1];
  assign _zz_711_ = _zz_708_[2];
  assign _zz_712_ = _zz_708_[3];
  assign _zz_713_ = _zz_708_[4];
  assign _zz_714_ = _zz_708_[5];
  assign _zz_715_ = _zz_708_[6];
  assign _zz_716_ = _zz_708_[7];
  assign _zz_717_ = _zz_708_[8];
  assign _zz_718_ = _zz_708_[9];
  assign _zz_719_ = _zz_708_[10];
  assign _zz_720_ = _zz_708_[11];
  assign _zz_721_ = _zz_708_[12];
  assign _zz_722_ = _zz_708_[13];
  assign _zz_723_ = _zz_708_[14];
  assign _zz_724_ = _zz_708_[15];
  assign _zz_725_ = _zz_708_[16];
  assign _zz_726_ = _zz_708_[17];
  assign _zz_727_ = _zz_708_[18];
  assign _zz_728_ = _zz_708_[19];
  assign _zz_729_ = _zz_708_[20];
  assign _zz_730_ = _zz_708_[21];
  assign _zz_731_ = _zz_708_[22];
  assign _zz_732_ = _zz_708_[23];
  assign _zz_733_ = _zz_708_[24];
  assign _zz_734_ = _zz_708_[25];
  assign _zz_735_ = _zz_708_[26];
  assign _zz_736_ = _zz_708_[27];
  assign _zz_737_ = _zz_708_[28];
  assign _zz_738_ = _zz_708_[29];
  assign _zz_739_ = _zz_708_[30];
  assign _zz_740_ = _zz_708_[31];
  assign _zz_741_ = _zz_708_[32];
  assign _zz_742_ = _zz_708_[33];
  assign _zz_743_ = _zz_708_[34];
  assign _zz_744_ = _zz_708_[35];
  assign _zz_745_ = _zz_708_[36];
  assign _zz_746_ = _zz_708_[37];
  assign _zz_747_ = _zz_708_[38];
  assign _zz_748_ = _zz_708_[39];
  assign _zz_749_ = _zz_708_[40];
  assign _zz_750_ = _zz_708_[41];
  assign _zz_751_ = _zz_708_[42];
  assign _zz_752_ = _zz_708_[43];
  assign _zz_753_ = _zz_708_[44];
  assign _zz_754_ = _zz_708_[45];
  assign _zz_755_ = _zz_708_[46];
  assign _zz_756_ = _zz_708_[47];
  assign _zz_757_ = _zz_708_[48];
  assign _zz_758_ = _zz_708_[49];
  assign _zz_759_ = _zz_708_[50];
  assign _zz_760_ = _zz_708_[51];
  assign _zz_761_ = _zz_708_[52];
  assign _zz_762_ = _zz_708_[53];
  assign _zz_763_ = _zz_708_[54];
  assign _zz_764_ = _zz_708_[55];
  assign _zz_765_ = _zz_708_[56];
  assign _zz_766_ = _zz_708_[57];
  assign _zz_767_ = _zz_708_[58];
  assign _zz_768_ = _zz_708_[59];
  assign _zz_769_ = _zz_708_[60];
  assign _zz_770_ = _zz_708_[61];
  assign _zz_771_ = _zz_708_[62];
  assign _zz_772_ = _zz_708_[63];
  assign _zz_773_ = (((32'h00000780 <= load_data_area_current_addr) && (load_data_area_current_addr < 32'h000007c0)) ? _zz_9__regNext : {_zz_4454_,_zz_4455_});
  assign _zz_774_ = _zz_773_[15 : 0];
  assign _zz_775_ = _zz_773_[31 : 16];
  assign _zz_776_ = _zz_4577_[5:0];
  assign _zz_777_ = ({63'd0,(1'b1)} <<< _zz_776_);
  assign _zz_778_ = _zz_777_[0];
  assign _zz_779_ = _zz_777_[1];
  assign _zz_780_ = _zz_777_[2];
  assign _zz_781_ = _zz_777_[3];
  assign _zz_782_ = _zz_777_[4];
  assign _zz_783_ = _zz_777_[5];
  assign _zz_784_ = _zz_777_[6];
  assign _zz_785_ = _zz_777_[7];
  assign _zz_786_ = _zz_777_[8];
  assign _zz_787_ = _zz_777_[9];
  assign _zz_788_ = _zz_777_[10];
  assign _zz_789_ = _zz_777_[11];
  assign _zz_790_ = _zz_777_[12];
  assign _zz_791_ = _zz_777_[13];
  assign _zz_792_ = _zz_777_[14];
  assign _zz_793_ = _zz_777_[15];
  assign _zz_794_ = _zz_777_[16];
  assign _zz_795_ = _zz_777_[17];
  assign _zz_796_ = _zz_777_[18];
  assign _zz_797_ = _zz_777_[19];
  assign _zz_798_ = _zz_777_[20];
  assign _zz_799_ = _zz_777_[21];
  assign _zz_800_ = _zz_777_[22];
  assign _zz_801_ = _zz_777_[23];
  assign _zz_802_ = _zz_777_[24];
  assign _zz_803_ = _zz_777_[25];
  assign _zz_804_ = _zz_777_[26];
  assign _zz_805_ = _zz_777_[27];
  assign _zz_806_ = _zz_777_[28];
  assign _zz_807_ = _zz_777_[29];
  assign _zz_808_ = _zz_777_[30];
  assign _zz_809_ = _zz_777_[31];
  assign _zz_810_ = _zz_777_[32];
  assign _zz_811_ = _zz_777_[33];
  assign _zz_812_ = _zz_777_[34];
  assign _zz_813_ = _zz_777_[35];
  assign _zz_814_ = _zz_777_[36];
  assign _zz_815_ = _zz_777_[37];
  assign _zz_816_ = _zz_777_[38];
  assign _zz_817_ = _zz_777_[39];
  assign _zz_818_ = _zz_777_[40];
  assign _zz_819_ = _zz_777_[41];
  assign _zz_820_ = _zz_777_[42];
  assign _zz_821_ = _zz_777_[43];
  assign _zz_822_ = _zz_777_[44];
  assign _zz_823_ = _zz_777_[45];
  assign _zz_824_ = _zz_777_[46];
  assign _zz_825_ = _zz_777_[47];
  assign _zz_826_ = _zz_777_[48];
  assign _zz_827_ = _zz_777_[49];
  assign _zz_828_ = _zz_777_[50];
  assign _zz_829_ = _zz_777_[51];
  assign _zz_830_ = _zz_777_[52];
  assign _zz_831_ = _zz_777_[53];
  assign _zz_832_ = _zz_777_[54];
  assign _zz_833_ = _zz_777_[55];
  assign _zz_834_ = _zz_777_[56];
  assign _zz_835_ = _zz_777_[57];
  assign _zz_836_ = _zz_777_[58];
  assign _zz_837_ = _zz_777_[59];
  assign _zz_838_ = _zz_777_[60];
  assign _zz_839_ = _zz_777_[61];
  assign _zz_840_ = _zz_777_[62];
  assign _zz_841_ = _zz_777_[63];
  assign _zz_842_ = (((32'h00000580 <= load_data_area_current_addr) && (load_data_area_current_addr < 32'h000005c0)) ? _zz_9__regNext : {_zz_4456_,_zz_4457_});
  assign _zz_843_ = _zz_842_[15 : 0];
  assign _zz_844_ = _zz_842_[31 : 16];
  assign _zz_845_ = _zz_4578_[5:0];
  assign _zz_846_ = ({63'd0,(1'b1)} <<< _zz_845_);
  assign _zz_847_ = _zz_846_[0];
  assign _zz_848_ = _zz_846_[1];
  assign _zz_849_ = _zz_846_[2];
  assign _zz_850_ = _zz_846_[3];
  assign _zz_851_ = _zz_846_[4];
  assign _zz_852_ = _zz_846_[5];
  assign _zz_853_ = _zz_846_[6];
  assign _zz_854_ = _zz_846_[7];
  assign _zz_855_ = _zz_846_[8];
  assign _zz_856_ = _zz_846_[9];
  assign _zz_857_ = _zz_846_[10];
  assign _zz_858_ = _zz_846_[11];
  assign _zz_859_ = _zz_846_[12];
  assign _zz_860_ = _zz_846_[13];
  assign _zz_861_ = _zz_846_[14];
  assign _zz_862_ = _zz_846_[15];
  assign _zz_863_ = _zz_846_[16];
  assign _zz_864_ = _zz_846_[17];
  assign _zz_865_ = _zz_846_[18];
  assign _zz_866_ = _zz_846_[19];
  assign _zz_867_ = _zz_846_[20];
  assign _zz_868_ = _zz_846_[21];
  assign _zz_869_ = _zz_846_[22];
  assign _zz_870_ = _zz_846_[23];
  assign _zz_871_ = _zz_846_[24];
  assign _zz_872_ = _zz_846_[25];
  assign _zz_873_ = _zz_846_[26];
  assign _zz_874_ = _zz_846_[27];
  assign _zz_875_ = _zz_846_[28];
  assign _zz_876_ = _zz_846_[29];
  assign _zz_877_ = _zz_846_[30];
  assign _zz_878_ = _zz_846_[31];
  assign _zz_879_ = _zz_846_[32];
  assign _zz_880_ = _zz_846_[33];
  assign _zz_881_ = _zz_846_[34];
  assign _zz_882_ = _zz_846_[35];
  assign _zz_883_ = _zz_846_[36];
  assign _zz_884_ = _zz_846_[37];
  assign _zz_885_ = _zz_846_[38];
  assign _zz_886_ = _zz_846_[39];
  assign _zz_887_ = _zz_846_[40];
  assign _zz_888_ = _zz_846_[41];
  assign _zz_889_ = _zz_846_[42];
  assign _zz_890_ = _zz_846_[43];
  assign _zz_891_ = _zz_846_[44];
  assign _zz_892_ = _zz_846_[45];
  assign _zz_893_ = _zz_846_[46];
  assign _zz_894_ = _zz_846_[47];
  assign _zz_895_ = _zz_846_[48];
  assign _zz_896_ = _zz_846_[49];
  assign _zz_897_ = _zz_846_[50];
  assign _zz_898_ = _zz_846_[51];
  assign _zz_899_ = _zz_846_[52];
  assign _zz_900_ = _zz_846_[53];
  assign _zz_901_ = _zz_846_[54];
  assign _zz_902_ = _zz_846_[55];
  assign _zz_903_ = _zz_846_[56];
  assign _zz_904_ = _zz_846_[57];
  assign _zz_905_ = _zz_846_[58];
  assign _zz_906_ = _zz_846_[59];
  assign _zz_907_ = _zz_846_[60];
  assign _zz_908_ = _zz_846_[61];
  assign _zz_909_ = _zz_846_[62];
  assign _zz_910_ = _zz_846_[63];
  assign _zz_911_ = (((32'h00000500 <= load_data_area_current_addr) && (load_data_area_current_addr < 32'h00000540)) ? _zz_9__regNext : {_zz_4458_,_zz_4459_});
  assign _zz_912_ = _zz_911_[15 : 0];
  assign _zz_913_ = _zz_911_[31 : 16];
  assign _zz_914_ = _zz_4579_[5:0];
  assign _zz_915_ = ({63'd0,(1'b1)} <<< _zz_914_);
  assign _zz_916_ = _zz_915_[0];
  assign _zz_917_ = _zz_915_[1];
  assign _zz_918_ = _zz_915_[2];
  assign _zz_919_ = _zz_915_[3];
  assign _zz_920_ = _zz_915_[4];
  assign _zz_921_ = _zz_915_[5];
  assign _zz_922_ = _zz_915_[6];
  assign _zz_923_ = _zz_915_[7];
  assign _zz_924_ = _zz_915_[8];
  assign _zz_925_ = _zz_915_[9];
  assign _zz_926_ = _zz_915_[10];
  assign _zz_927_ = _zz_915_[11];
  assign _zz_928_ = _zz_915_[12];
  assign _zz_929_ = _zz_915_[13];
  assign _zz_930_ = _zz_915_[14];
  assign _zz_931_ = _zz_915_[15];
  assign _zz_932_ = _zz_915_[16];
  assign _zz_933_ = _zz_915_[17];
  assign _zz_934_ = _zz_915_[18];
  assign _zz_935_ = _zz_915_[19];
  assign _zz_936_ = _zz_915_[20];
  assign _zz_937_ = _zz_915_[21];
  assign _zz_938_ = _zz_915_[22];
  assign _zz_939_ = _zz_915_[23];
  assign _zz_940_ = _zz_915_[24];
  assign _zz_941_ = _zz_915_[25];
  assign _zz_942_ = _zz_915_[26];
  assign _zz_943_ = _zz_915_[27];
  assign _zz_944_ = _zz_915_[28];
  assign _zz_945_ = _zz_915_[29];
  assign _zz_946_ = _zz_915_[30];
  assign _zz_947_ = _zz_915_[31];
  assign _zz_948_ = _zz_915_[32];
  assign _zz_949_ = _zz_915_[33];
  assign _zz_950_ = _zz_915_[34];
  assign _zz_951_ = _zz_915_[35];
  assign _zz_952_ = _zz_915_[36];
  assign _zz_953_ = _zz_915_[37];
  assign _zz_954_ = _zz_915_[38];
  assign _zz_955_ = _zz_915_[39];
  assign _zz_956_ = _zz_915_[40];
  assign _zz_957_ = _zz_915_[41];
  assign _zz_958_ = _zz_915_[42];
  assign _zz_959_ = _zz_915_[43];
  assign _zz_960_ = _zz_915_[44];
  assign _zz_961_ = _zz_915_[45];
  assign _zz_962_ = _zz_915_[46];
  assign _zz_963_ = _zz_915_[47];
  assign _zz_964_ = _zz_915_[48];
  assign _zz_965_ = _zz_915_[49];
  assign _zz_966_ = _zz_915_[50];
  assign _zz_967_ = _zz_915_[51];
  assign _zz_968_ = _zz_915_[52];
  assign _zz_969_ = _zz_915_[53];
  assign _zz_970_ = _zz_915_[54];
  assign _zz_971_ = _zz_915_[55];
  assign _zz_972_ = _zz_915_[56];
  assign _zz_973_ = _zz_915_[57];
  assign _zz_974_ = _zz_915_[58];
  assign _zz_975_ = _zz_915_[59];
  assign _zz_976_ = _zz_915_[60];
  assign _zz_977_ = _zz_915_[61];
  assign _zz_978_ = _zz_915_[62];
  assign _zz_979_ = _zz_915_[63];
  assign _zz_980_ = (((32'h00000880 <= load_data_area_current_addr) && (load_data_area_current_addr < 32'h000008c0)) ? _zz_9__regNext : {_zz_4460_,_zz_4461_});
  assign _zz_981_ = _zz_980_[15 : 0];
  assign _zz_982_ = _zz_980_[31 : 16];
  assign _zz_983_ = _zz_4580_[5:0];
  assign _zz_984_ = ({63'd0,(1'b1)} <<< _zz_983_);
  assign _zz_985_ = _zz_984_[0];
  assign _zz_986_ = _zz_984_[1];
  assign _zz_987_ = _zz_984_[2];
  assign _zz_988_ = _zz_984_[3];
  assign _zz_989_ = _zz_984_[4];
  assign _zz_990_ = _zz_984_[5];
  assign _zz_991_ = _zz_984_[6];
  assign _zz_992_ = _zz_984_[7];
  assign _zz_993_ = _zz_984_[8];
  assign _zz_994_ = _zz_984_[9];
  assign _zz_995_ = _zz_984_[10];
  assign _zz_996_ = _zz_984_[11];
  assign _zz_997_ = _zz_984_[12];
  assign _zz_998_ = _zz_984_[13];
  assign _zz_999_ = _zz_984_[14];
  assign _zz_1000_ = _zz_984_[15];
  assign _zz_1001_ = _zz_984_[16];
  assign _zz_1002_ = _zz_984_[17];
  assign _zz_1003_ = _zz_984_[18];
  assign _zz_1004_ = _zz_984_[19];
  assign _zz_1005_ = _zz_984_[20];
  assign _zz_1006_ = _zz_984_[21];
  assign _zz_1007_ = _zz_984_[22];
  assign _zz_1008_ = _zz_984_[23];
  assign _zz_1009_ = _zz_984_[24];
  assign _zz_1010_ = _zz_984_[25];
  assign _zz_1011_ = _zz_984_[26];
  assign _zz_1012_ = _zz_984_[27];
  assign _zz_1013_ = _zz_984_[28];
  assign _zz_1014_ = _zz_984_[29];
  assign _zz_1015_ = _zz_984_[30];
  assign _zz_1016_ = _zz_984_[31];
  assign _zz_1017_ = _zz_984_[32];
  assign _zz_1018_ = _zz_984_[33];
  assign _zz_1019_ = _zz_984_[34];
  assign _zz_1020_ = _zz_984_[35];
  assign _zz_1021_ = _zz_984_[36];
  assign _zz_1022_ = _zz_984_[37];
  assign _zz_1023_ = _zz_984_[38];
  assign _zz_1024_ = _zz_984_[39];
  assign _zz_1025_ = _zz_984_[40];
  assign _zz_1026_ = _zz_984_[41];
  assign _zz_1027_ = _zz_984_[42];
  assign _zz_1028_ = _zz_984_[43];
  assign _zz_1029_ = _zz_984_[44];
  assign _zz_1030_ = _zz_984_[45];
  assign _zz_1031_ = _zz_984_[46];
  assign _zz_1032_ = _zz_984_[47];
  assign _zz_1033_ = _zz_984_[48];
  assign _zz_1034_ = _zz_984_[49];
  assign _zz_1035_ = _zz_984_[50];
  assign _zz_1036_ = _zz_984_[51];
  assign _zz_1037_ = _zz_984_[52];
  assign _zz_1038_ = _zz_984_[53];
  assign _zz_1039_ = _zz_984_[54];
  assign _zz_1040_ = _zz_984_[55];
  assign _zz_1041_ = _zz_984_[56];
  assign _zz_1042_ = _zz_984_[57];
  assign _zz_1043_ = _zz_984_[58];
  assign _zz_1044_ = _zz_984_[59];
  assign _zz_1045_ = _zz_984_[60];
  assign _zz_1046_ = _zz_984_[61];
  assign _zz_1047_ = _zz_984_[62];
  assign _zz_1048_ = _zz_984_[63];
  assign _zz_1049_ = (((32'h00000180 <= load_data_area_current_addr) && (load_data_area_current_addr < 32'h000001c0)) ? _zz_9__regNext : {_zz_4462_,_zz_4463_});
  assign _zz_1050_ = _zz_1049_[15 : 0];
  assign _zz_1051_ = _zz_1049_[31 : 16];
  assign _zz_1052_ = _zz_4581_[5:0];
  assign _zz_1053_ = ({63'd0,(1'b1)} <<< _zz_1052_);
  assign _zz_1054_ = _zz_1053_[0];
  assign _zz_1055_ = _zz_1053_[1];
  assign _zz_1056_ = _zz_1053_[2];
  assign _zz_1057_ = _zz_1053_[3];
  assign _zz_1058_ = _zz_1053_[4];
  assign _zz_1059_ = _zz_1053_[5];
  assign _zz_1060_ = _zz_1053_[6];
  assign _zz_1061_ = _zz_1053_[7];
  assign _zz_1062_ = _zz_1053_[8];
  assign _zz_1063_ = _zz_1053_[9];
  assign _zz_1064_ = _zz_1053_[10];
  assign _zz_1065_ = _zz_1053_[11];
  assign _zz_1066_ = _zz_1053_[12];
  assign _zz_1067_ = _zz_1053_[13];
  assign _zz_1068_ = _zz_1053_[14];
  assign _zz_1069_ = _zz_1053_[15];
  assign _zz_1070_ = _zz_1053_[16];
  assign _zz_1071_ = _zz_1053_[17];
  assign _zz_1072_ = _zz_1053_[18];
  assign _zz_1073_ = _zz_1053_[19];
  assign _zz_1074_ = _zz_1053_[20];
  assign _zz_1075_ = _zz_1053_[21];
  assign _zz_1076_ = _zz_1053_[22];
  assign _zz_1077_ = _zz_1053_[23];
  assign _zz_1078_ = _zz_1053_[24];
  assign _zz_1079_ = _zz_1053_[25];
  assign _zz_1080_ = _zz_1053_[26];
  assign _zz_1081_ = _zz_1053_[27];
  assign _zz_1082_ = _zz_1053_[28];
  assign _zz_1083_ = _zz_1053_[29];
  assign _zz_1084_ = _zz_1053_[30];
  assign _zz_1085_ = _zz_1053_[31];
  assign _zz_1086_ = _zz_1053_[32];
  assign _zz_1087_ = _zz_1053_[33];
  assign _zz_1088_ = _zz_1053_[34];
  assign _zz_1089_ = _zz_1053_[35];
  assign _zz_1090_ = _zz_1053_[36];
  assign _zz_1091_ = _zz_1053_[37];
  assign _zz_1092_ = _zz_1053_[38];
  assign _zz_1093_ = _zz_1053_[39];
  assign _zz_1094_ = _zz_1053_[40];
  assign _zz_1095_ = _zz_1053_[41];
  assign _zz_1096_ = _zz_1053_[42];
  assign _zz_1097_ = _zz_1053_[43];
  assign _zz_1098_ = _zz_1053_[44];
  assign _zz_1099_ = _zz_1053_[45];
  assign _zz_1100_ = _zz_1053_[46];
  assign _zz_1101_ = _zz_1053_[47];
  assign _zz_1102_ = _zz_1053_[48];
  assign _zz_1103_ = _zz_1053_[49];
  assign _zz_1104_ = _zz_1053_[50];
  assign _zz_1105_ = _zz_1053_[51];
  assign _zz_1106_ = _zz_1053_[52];
  assign _zz_1107_ = _zz_1053_[53];
  assign _zz_1108_ = _zz_1053_[54];
  assign _zz_1109_ = _zz_1053_[55];
  assign _zz_1110_ = _zz_1053_[56];
  assign _zz_1111_ = _zz_1053_[57];
  assign _zz_1112_ = _zz_1053_[58];
  assign _zz_1113_ = _zz_1053_[59];
  assign _zz_1114_ = _zz_1053_[60];
  assign _zz_1115_ = _zz_1053_[61];
  assign _zz_1116_ = _zz_1053_[62];
  assign _zz_1117_ = _zz_1053_[63];
  assign _zz_1118_ = (((32'h00000200 <= load_data_area_current_addr) && (load_data_area_current_addr < 32'h00000240)) ? _zz_9__regNext : {_zz_4464_,_zz_4465_});
  assign _zz_1119_ = _zz_1118_[15 : 0];
  assign _zz_1120_ = _zz_1118_[31 : 16];
  assign _zz_1121_ = _zz_4582_[5:0];
  assign _zz_1122_ = ({63'd0,(1'b1)} <<< _zz_1121_);
  assign _zz_1123_ = _zz_1122_[0];
  assign _zz_1124_ = _zz_1122_[1];
  assign _zz_1125_ = _zz_1122_[2];
  assign _zz_1126_ = _zz_1122_[3];
  assign _zz_1127_ = _zz_1122_[4];
  assign _zz_1128_ = _zz_1122_[5];
  assign _zz_1129_ = _zz_1122_[6];
  assign _zz_1130_ = _zz_1122_[7];
  assign _zz_1131_ = _zz_1122_[8];
  assign _zz_1132_ = _zz_1122_[9];
  assign _zz_1133_ = _zz_1122_[10];
  assign _zz_1134_ = _zz_1122_[11];
  assign _zz_1135_ = _zz_1122_[12];
  assign _zz_1136_ = _zz_1122_[13];
  assign _zz_1137_ = _zz_1122_[14];
  assign _zz_1138_ = _zz_1122_[15];
  assign _zz_1139_ = _zz_1122_[16];
  assign _zz_1140_ = _zz_1122_[17];
  assign _zz_1141_ = _zz_1122_[18];
  assign _zz_1142_ = _zz_1122_[19];
  assign _zz_1143_ = _zz_1122_[20];
  assign _zz_1144_ = _zz_1122_[21];
  assign _zz_1145_ = _zz_1122_[22];
  assign _zz_1146_ = _zz_1122_[23];
  assign _zz_1147_ = _zz_1122_[24];
  assign _zz_1148_ = _zz_1122_[25];
  assign _zz_1149_ = _zz_1122_[26];
  assign _zz_1150_ = _zz_1122_[27];
  assign _zz_1151_ = _zz_1122_[28];
  assign _zz_1152_ = _zz_1122_[29];
  assign _zz_1153_ = _zz_1122_[30];
  assign _zz_1154_ = _zz_1122_[31];
  assign _zz_1155_ = _zz_1122_[32];
  assign _zz_1156_ = _zz_1122_[33];
  assign _zz_1157_ = _zz_1122_[34];
  assign _zz_1158_ = _zz_1122_[35];
  assign _zz_1159_ = _zz_1122_[36];
  assign _zz_1160_ = _zz_1122_[37];
  assign _zz_1161_ = _zz_1122_[38];
  assign _zz_1162_ = _zz_1122_[39];
  assign _zz_1163_ = _zz_1122_[40];
  assign _zz_1164_ = _zz_1122_[41];
  assign _zz_1165_ = _zz_1122_[42];
  assign _zz_1166_ = _zz_1122_[43];
  assign _zz_1167_ = _zz_1122_[44];
  assign _zz_1168_ = _zz_1122_[45];
  assign _zz_1169_ = _zz_1122_[46];
  assign _zz_1170_ = _zz_1122_[47];
  assign _zz_1171_ = _zz_1122_[48];
  assign _zz_1172_ = _zz_1122_[49];
  assign _zz_1173_ = _zz_1122_[50];
  assign _zz_1174_ = _zz_1122_[51];
  assign _zz_1175_ = _zz_1122_[52];
  assign _zz_1176_ = _zz_1122_[53];
  assign _zz_1177_ = _zz_1122_[54];
  assign _zz_1178_ = _zz_1122_[55];
  assign _zz_1179_ = _zz_1122_[56];
  assign _zz_1180_ = _zz_1122_[57];
  assign _zz_1181_ = _zz_1122_[58];
  assign _zz_1182_ = _zz_1122_[59];
  assign _zz_1183_ = _zz_1122_[60];
  assign _zz_1184_ = _zz_1122_[61];
  assign _zz_1185_ = _zz_1122_[62];
  assign _zz_1186_ = _zz_1122_[63];
  assign _zz_1187_ = (((32'h000006c0 <= load_data_area_current_addr) && (load_data_area_current_addr < 32'h00000700)) ? _zz_9__regNext : {_zz_4466_,_zz_4467_});
  assign _zz_1188_ = _zz_1187_[15 : 0];
  assign _zz_1189_ = _zz_1187_[31 : 16];
  assign _zz_1190_ = _zz_4583_[5:0];
  assign _zz_1191_ = ({63'd0,(1'b1)} <<< _zz_1190_);
  assign _zz_1192_ = _zz_1191_[0];
  assign _zz_1193_ = _zz_1191_[1];
  assign _zz_1194_ = _zz_1191_[2];
  assign _zz_1195_ = _zz_1191_[3];
  assign _zz_1196_ = _zz_1191_[4];
  assign _zz_1197_ = _zz_1191_[5];
  assign _zz_1198_ = _zz_1191_[6];
  assign _zz_1199_ = _zz_1191_[7];
  assign _zz_1200_ = _zz_1191_[8];
  assign _zz_1201_ = _zz_1191_[9];
  assign _zz_1202_ = _zz_1191_[10];
  assign _zz_1203_ = _zz_1191_[11];
  assign _zz_1204_ = _zz_1191_[12];
  assign _zz_1205_ = _zz_1191_[13];
  assign _zz_1206_ = _zz_1191_[14];
  assign _zz_1207_ = _zz_1191_[15];
  assign _zz_1208_ = _zz_1191_[16];
  assign _zz_1209_ = _zz_1191_[17];
  assign _zz_1210_ = _zz_1191_[18];
  assign _zz_1211_ = _zz_1191_[19];
  assign _zz_1212_ = _zz_1191_[20];
  assign _zz_1213_ = _zz_1191_[21];
  assign _zz_1214_ = _zz_1191_[22];
  assign _zz_1215_ = _zz_1191_[23];
  assign _zz_1216_ = _zz_1191_[24];
  assign _zz_1217_ = _zz_1191_[25];
  assign _zz_1218_ = _zz_1191_[26];
  assign _zz_1219_ = _zz_1191_[27];
  assign _zz_1220_ = _zz_1191_[28];
  assign _zz_1221_ = _zz_1191_[29];
  assign _zz_1222_ = _zz_1191_[30];
  assign _zz_1223_ = _zz_1191_[31];
  assign _zz_1224_ = _zz_1191_[32];
  assign _zz_1225_ = _zz_1191_[33];
  assign _zz_1226_ = _zz_1191_[34];
  assign _zz_1227_ = _zz_1191_[35];
  assign _zz_1228_ = _zz_1191_[36];
  assign _zz_1229_ = _zz_1191_[37];
  assign _zz_1230_ = _zz_1191_[38];
  assign _zz_1231_ = _zz_1191_[39];
  assign _zz_1232_ = _zz_1191_[40];
  assign _zz_1233_ = _zz_1191_[41];
  assign _zz_1234_ = _zz_1191_[42];
  assign _zz_1235_ = _zz_1191_[43];
  assign _zz_1236_ = _zz_1191_[44];
  assign _zz_1237_ = _zz_1191_[45];
  assign _zz_1238_ = _zz_1191_[46];
  assign _zz_1239_ = _zz_1191_[47];
  assign _zz_1240_ = _zz_1191_[48];
  assign _zz_1241_ = _zz_1191_[49];
  assign _zz_1242_ = _zz_1191_[50];
  assign _zz_1243_ = _zz_1191_[51];
  assign _zz_1244_ = _zz_1191_[52];
  assign _zz_1245_ = _zz_1191_[53];
  assign _zz_1246_ = _zz_1191_[54];
  assign _zz_1247_ = _zz_1191_[55];
  assign _zz_1248_ = _zz_1191_[56];
  assign _zz_1249_ = _zz_1191_[57];
  assign _zz_1250_ = _zz_1191_[58];
  assign _zz_1251_ = _zz_1191_[59];
  assign _zz_1252_ = _zz_1191_[60];
  assign _zz_1253_ = _zz_1191_[61];
  assign _zz_1254_ = _zz_1191_[62];
  assign _zz_1255_ = _zz_1191_[63];
  assign _zz_1256_ = (((32'h000004c0 <= load_data_area_current_addr) && (load_data_area_current_addr < 32'h00000500)) ? _zz_9__regNext : {_zz_4468_,_zz_4469_});
  assign _zz_1257_ = _zz_1256_[15 : 0];
  assign _zz_1258_ = _zz_1256_[31 : 16];
  assign _zz_1259_ = _zz_4584_[5:0];
  assign _zz_1260_ = ({63'd0,(1'b1)} <<< _zz_1259_);
  assign _zz_1261_ = _zz_1260_[0];
  assign _zz_1262_ = _zz_1260_[1];
  assign _zz_1263_ = _zz_1260_[2];
  assign _zz_1264_ = _zz_1260_[3];
  assign _zz_1265_ = _zz_1260_[4];
  assign _zz_1266_ = _zz_1260_[5];
  assign _zz_1267_ = _zz_1260_[6];
  assign _zz_1268_ = _zz_1260_[7];
  assign _zz_1269_ = _zz_1260_[8];
  assign _zz_1270_ = _zz_1260_[9];
  assign _zz_1271_ = _zz_1260_[10];
  assign _zz_1272_ = _zz_1260_[11];
  assign _zz_1273_ = _zz_1260_[12];
  assign _zz_1274_ = _zz_1260_[13];
  assign _zz_1275_ = _zz_1260_[14];
  assign _zz_1276_ = _zz_1260_[15];
  assign _zz_1277_ = _zz_1260_[16];
  assign _zz_1278_ = _zz_1260_[17];
  assign _zz_1279_ = _zz_1260_[18];
  assign _zz_1280_ = _zz_1260_[19];
  assign _zz_1281_ = _zz_1260_[20];
  assign _zz_1282_ = _zz_1260_[21];
  assign _zz_1283_ = _zz_1260_[22];
  assign _zz_1284_ = _zz_1260_[23];
  assign _zz_1285_ = _zz_1260_[24];
  assign _zz_1286_ = _zz_1260_[25];
  assign _zz_1287_ = _zz_1260_[26];
  assign _zz_1288_ = _zz_1260_[27];
  assign _zz_1289_ = _zz_1260_[28];
  assign _zz_1290_ = _zz_1260_[29];
  assign _zz_1291_ = _zz_1260_[30];
  assign _zz_1292_ = _zz_1260_[31];
  assign _zz_1293_ = _zz_1260_[32];
  assign _zz_1294_ = _zz_1260_[33];
  assign _zz_1295_ = _zz_1260_[34];
  assign _zz_1296_ = _zz_1260_[35];
  assign _zz_1297_ = _zz_1260_[36];
  assign _zz_1298_ = _zz_1260_[37];
  assign _zz_1299_ = _zz_1260_[38];
  assign _zz_1300_ = _zz_1260_[39];
  assign _zz_1301_ = _zz_1260_[40];
  assign _zz_1302_ = _zz_1260_[41];
  assign _zz_1303_ = _zz_1260_[42];
  assign _zz_1304_ = _zz_1260_[43];
  assign _zz_1305_ = _zz_1260_[44];
  assign _zz_1306_ = _zz_1260_[45];
  assign _zz_1307_ = _zz_1260_[46];
  assign _zz_1308_ = _zz_1260_[47];
  assign _zz_1309_ = _zz_1260_[48];
  assign _zz_1310_ = _zz_1260_[49];
  assign _zz_1311_ = _zz_1260_[50];
  assign _zz_1312_ = _zz_1260_[51];
  assign _zz_1313_ = _zz_1260_[52];
  assign _zz_1314_ = _zz_1260_[53];
  assign _zz_1315_ = _zz_1260_[54];
  assign _zz_1316_ = _zz_1260_[55];
  assign _zz_1317_ = _zz_1260_[56];
  assign _zz_1318_ = _zz_1260_[57];
  assign _zz_1319_ = _zz_1260_[58];
  assign _zz_1320_ = _zz_1260_[59];
  assign _zz_1321_ = _zz_1260_[60];
  assign _zz_1322_ = _zz_1260_[61];
  assign _zz_1323_ = _zz_1260_[62];
  assign _zz_1324_ = _zz_1260_[63];
  assign _zz_1325_ = (((32'h00000c40 <= load_data_area_current_addr) && (load_data_area_current_addr < 32'h00000c80)) ? _zz_9__regNext : {_zz_4470_,_zz_4471_});
  assign _zz_1326_ = _zz_1325_[15 : 0];
  assign _zz_1327_ = _zz_1325_[31 : 16];
  assign _zz_1328_ = _zz_4585_[5:0];
  assign _zz_1329_ = ({63'd0,(1'b1)} <<< _zz_1328_);
  assign _zz_1330_ = _zz_1329_[0];
  assign _zz_1331_ = _zz_1329_[1];
  assign _zz_1332_ = _zz_1329_[2];
  assign _zz_1333_ = _zz_1329_[3];
  assign _zz_1334_ = _zz_1329_[4];
  assign _zz_1335_ = _zz_1329_[5];
  assign _zz_1336_ = _zz_1329_[6];
  assign _zz_1337_ = _zz_1329_[7];
  assign _zz_1338_ = _zz_1329_[8];
  assign _zz_1339_ = _zz_1329_[9];
  assign _zz_1340_ = _zz_1329_[10];
  assign _zz_1341_ = _zz_1329_[11];
  assign _zz_1342_ = _zz_1329_[12];
  assign _zz_1343_ = _zz_1329_[13];
  assign _zz_1344_ = _zz_1329_[14];
  assign _zz_1345_ = _zz_1329_[15];
  assign _zz_1346_ = _zz_1329_[16];
  assign _zz_1347_ = _zz_1329_[17];
  assign _zz_1348_ = _zz_1329_[18];
  assign _zz_1349_ = _zz_1329_[19];
  assign _zz_1350_ = _zz_1329_[20];
  assign _zz_1351_ = _zz_1329_[21];
  assign _zz_1352_ = _zz_1329_[22];
  assign _zz_1353_ = _zz_1329_[23];
  assign _zz_1354_ = _zz_1329_[24];
  assign _zz_1355_ = _zz_1329_[25];
  assign _zz_1356_ = _zz_1329_[26];
  assign _zz_1357_ = _zz_1329_[27];
  assign _zz_1358_ = _zz_1329_[28];
  assign _zz_1359_ = _zz_1329_[29];
  assign _zz_1360_ = _zz_1329_[30];
  assign _zz_1361_ = _zz_1329_[31];
  assign _zz_1362_ = _zz_1329_[32];
  assign _zz_1363_ = _zz_1329_[33];
  assign _zz_1364_ = _zz_1329_[34];
  assign _zz_1365_ = _zz_1329_[35];
  assign _zz_1366_ = _zz_1329_[36];
  assign _zz_1367_ = _zz_1329_[37];
  assign _zz_1368_ = _zz_1329_[38];
  assign _zz_1369_ = _zz_1329_[39];
  assign _zz_1370_ = _zz_1329_[40];
  assign _zz_1371_ = _zz_1329_[41];
  assign _zz_1372_ = _zz_1329_[42];
  assign _zz_1373_ = _zz_1329_[43];
  assign _zz_1374_ = _zz_1329_[44];
  assign _zz_1375_ = _zz_1329_[45];
  assign _zz_1376_ = _zz_1329_[46];
  assign _zz_1377_ = _zz_1329_[47];
  assign _zz_1378_ = _zz_1329_[48];
  assign _zz_1379_ = _zz_1329_[49];
  assign _zz_1380_ = _zz_1329_[50];
  assign _zz_1381_ = _zz_1329_[51];
  assign _zz_1382_ = _zz_1329_[52];
  assign _zz_1383_ = _zz_1329_[53];
  assign _zz_1384_ = _zz_1329_[54];
  assign _zz_1385_ = _zz_1329_[55];
  assign _zz_1386_ = _zz_1329_[56];
  assign _zz_1387_ = _zz_1329_[57];
  assign _zz_1388_ = _zz_1329_[58];
  assign _zz_1389_ = _zz_1329_[59];
  assign _zz_1390_ = _zz_1329_[60];
  assign _zz_1391_ = _zz_1329_[61];
  assign _zz_1392_ = _zz_1329_[62];
  assign _zz_1393_ = _zz_1329_[63];
  assign _zz_1394_ = (((32'h000001c0 <= load_data_area_current_addr) && (load_data_area_current_addr < 32'h00000200)) ? _zz_9__regNext : {_zz_4472_,_zz_4473_});
  assign _zz_1395_ = _zz_1394_[15 : 0];
  assign _zz_1396_ = _zz_1394_[31 : 16];
  assign _zz_1397_ = _zz_4586_[5:0];
  assign _zz_1398_ = ({63'd0,(1'b1)} <<< _zz_1397_);
  assign _zz_1399_ = _zz_1398_[0];
  assign _zz_1400_ = _zz_1398_[1];
  assign _zz_1401_ = _zz_1398_[2];
  assign _zz_1402_ = _zz_1398_[3];
  assign _zz_1403_ = _zz_1398_[4];
  assign _zz_1404_ = _zz_1398_[5];
  assign _zz_1405_ = _zz_1398_[6];
  assign _zz_1406_ = _zz_1398_[7];
  assign _zz_1407_ = _zz_1398_[8];
  assign _zz_1408_ = _zz_1398_[9];
  assign _zz_1409_ = _zz_1398_[10];
  assign _zz_1410_ = _zz_1398_[11];
  assign _zz_1411_ = _zz_1398_[12];
  assign _zz_1412_ = _zz_1398_[13];
  assign _zz_1413_ = _zz_1398_[14];
  assign _zz_1414_ = _zz_1398_[15];
  assign _zz_1415_ = _zz_1398_[16];
  assign _zz_1416_ = _zz_1398_[17];
  assign _zz_1417_ = _zz_1398_[18];
  assign _zz_1418_ = _zz_1398_[19];
  assign _zz_1419_ = _zz_1398_[20];
  assign _zz_1420_ = _zz_1398_[21];
  assign _zz_1421_ = _zz_1398_[22];
  assign _zz_1422_ = _zz_1398_[23];
  assign _zz_1423_ = _zz_1398_[24];
  assign _zz_1424_ = _zz_1398_[25];
  assign _zz_1425_ = _zz_1398_[26];
  assign _zz_1426_ = _zz_1398_[27];
  assign _zz_1427_ = _zz_1398_[28];
  assign _zz_1428_ = _zz_1398_[29];
  assign _zz_1429_ = _zz_1398_[30];
  assign _zz_1430_ = _zz_1398_[31];
  assign _zz_1431_ = _zz_1398_[32];
  assign _zz_1432_ = _zz_1398_[33];
  assign _zz_1433_ = _zz_1398_[34];
  assign _zz_1434_ = _zz_1398_[35];
  assign _zz_1435_ = _zz_1398_[36];
  assign _zz_1436_ = _zz_1398_[37];
  assign _zz_1437_ = _zz_1398_[38];
  assign _zz_1438_ = _zz_1398_[39];
  assign _zz_1439_ = _zz_1398_[40];
  assign _zz_1440_ = _zz_1398_[41];
  assign _zz_1441_ = _zz_1398_[42];
  assign _zz_1442_ = _zz_1398_[43];
  assign _zz_1443_ = _zz_1398_[44];
  assign _zz_1444_ = _zz_1398_[45];
  assign _zz_1445_ = _zz_1398_[46];
  assign _zz_1446_ = _zz_1398_[47];
  assign _zz_1447_ = _zz_1398_[48];
  assign _zz_1448_ = _zz_1398_[49];
  assign _zz_1449_ = _zz_1398_[50];
  assign _zz_1450_ = _zz_1398_[51];
  assign _zz_1451_ = _zz_1398_[52];
  assign _zz_1452_ = _zz_1398_[53];
  assign _zz_1453_ = _zz_1398_[54];
  assign _zz_1454_ = _zz_1398_[55];
  assign _zz_1455_ = _zz_1398_[56];
  assign _zz_1456_ = _zz_1398_[57];
  assign _zz_1457_ = _zz_1398_[58];
  assign _zz_1458_ = _zz_1398_[59];
  assign _zz_1459_ = _zz_1398_[60];
  assign _zz_1460_ = _zz_1398_[61];
  assign _zz_1461_ = _zz_1398_[62];
  assign _zz_1462_ = _zz_1398_[63];
  assign _zz_1463_ = (((32'h00000e80 <= load_data_area_current_addr) && (load_data_area_current_addr < 32'h00000ec0)) ? _zz_9__regNext : {_zz_4474_,_zz_4475_});
  assign _zz_1464_ = _zz_1463_[15 : 0];
  assign _zz_1465_ = _zz_1463_[31 : 16];
  assign _zz_1466_ = _zz_4587_[5:0];
  assign _zz_1467_ = ({63'd0,(1'b1)} <<< _zz_1466_);
  assign _zz_1468_ = _zz_1467_[0];
  assign _zz_1469_ = _zz_1467_[1];
  assign _zz_1470_ = _zz_1467_[2];
  assign _zz_1471_ = _zz_1467_[3];
  assign _zz_1472_ = _zz_1467_[4];
  assign _zz_1473_ = _zz_1467_[5];
  assign _zz_1474_ = _zz_1467_[6];
  assign _zz_1475_ = _zz_1467_[7];
  assign _zz_1476_ = _zz_1467_[8];
  assign _zz_1477_ = _zz_1467_[9];
  assign _zz_1478_ = _zz_1467_[10];
  assign _zz_1479_ = _zz_1467_[11];
  assign _zz_1480_ = _zz_1467_[12];
  assign _zz_1481_ = _zz_1467_[13];
  assign _zz_1482_ = _zz_1467_[14];
  assign _zz_1483_ = _zz_1467_[15];
  assign _zz_1484_ = _zz_1467_[16];
  assign _zz_1485_ = _zz_1467_[17];
  assign _zz_1486_ = _zz_1467_[18];
  assign _zz_1487_ = _zz_1467_[19];
  assign _zz_1488_ = _zz_1467_[20];
  assign _zz_1489_ = _zz_1467_[21];
  assign _zz_1490_ = _zz_1467_[22];
  assign _zz_1491_ = _zz_1467_[23];
  assign _zz_1492_ = _zz_1467_[24];
  assign _zz_1493_ = _zz_1467_[25];
  assign _zz_1494_ = _zz_1467_[26];
  assign _zz_1495_ = _zz_1467_[27];
  assign _zz_1496_ = _zz_1467_[28];
  assign _zz_1497_ = _zz_1467_[29];
  assign _zz_1498_ = _zz_1467_[30];
  assign _zz_1499_ = _zz_1467_[31];
  assign _zz_1500_ = _zz_1467_[32];
  assign _zz_1501_ = _zz_1467_[33];
  assign _zz_1502_ = _zz_1467_[34];
  assign _zz_1503_ = _zz_1467_[35];
  assign _zz_1504_ = _zz_1467_[36];
  assign _zz_1505_ = _zz_1467_[37];
  assign _zz_1506_ = _zz_1467_[38];
  assign _zz_1507_ = _zz_1467_[39];
  assign _zz_1508_ = _zz_1467_[40];
  assign _zz_1509_ = _zz_1467_[41];
  assign _zz_1510_ = _zz_1467_[42];
  assign _zz_1511_ = _zz_1467_[43];
  assign _zz_1512_ = _zz_1467_[44];
  assign _zz_1513_ = _zz_1467_[45];
  assign _zz_1514_ = _zz_1467_[46];
  assign _zz_1515_ = _zz_1467_[47];
  assign _zz_1516_ = _zz_1467_[48];
  assign _zz_1517_ = _zz_1467_[49];
  assign _zz_1518_ = _zz_1467_[50];
  assign _zz_1519_ = _zz_1467_[51];
  assign _zz_1520_ = _zz_1467_[52];
  assign _zz_1521_ = _zz_1467_[53];
  assign _zz_1522_ = _zz_1467_[54];
  assign _zz_1523_ = _zz_1467_[55];
  assign _zz_1524_ = _zz_1467_[56];
  assign _zz_1525_ = _zz_1467_[57];
  assign _zz_1526_ = _zz_1467_[58];
  assign _zz_1527_ = _zz_1467_[59];
  assign _zz_1528_ = _zz_1467_[60];
  assign _zz_1529_ = _zz_1467_[61];
  assign _zz_1530_ = _zz_1467_[62];
  assign _zz_1531_ = _zz_1467_[63];
  assign _zz_1532_ = (((32'h00000700 <= load_data_area_current_addr) && (load_data_area_current_addr < 32'h00000740)) ? _zz_9__regNext : {_zz_4476_,_zz_4477_});
  assign _zz_1533_ = _zz_1532_[15 : 0];
  assign _zz_1534_ = _zz_1532_[31 : 16];
  assign _zz_1535_ = _zz_4588_[5:0];
  assign _zz_1536_ = ({63'd0,(1'b1)} <<< _zz_1535_);
  assign _zz_1537_ = _zz_1536_[0];
  assign _zz_1538_ = _zz_1536_[1];
  assign _zz_1539_ = _zz_1536_[2];
  assign _zz_1540_ = _zz_1536_[3];
  assign _zz_1541_ = _zz_1536_[4];
  assign _zz_1542_ = _zz_1536_[5];
  assign _zz_1543_ = _zz_1536_[6];
  assign _zz_1544_ = _zz_1536_[7];
  assign _zz_1545_ = _zz_1536_[8];
  assign _zz_1546_ = _zz_1536_[9];
  assign _zz_1547_ = _zz_1536_[10];
  assign _zz_1548_ = _zz_1536_[11];
  assign _zz_1549_ = _zz_1536_[12];
  assign _zz_1550_ = _zz_1536_[13];
  assign _zz_1551_ = _zz_1536_[14];
  assign _zz_1552_ = _zz_1536_[15];
  assign _zz_1553_ = _zz_1536_[16];
  assign _zz_1554_ = _zz_1536_[17];
  assign _zz_1555_ = _zz_1536_[18];
  assign _zz_1556_ = _zz_1536_[19];
  assign _zz_1557_ = _zz_1536_[20];
  assign _zz_1558_ = _zz_1536_[21];
  assign _zz_1559_ = _zz_1536_[22];
  assign _zz_1560_ = _zz_1536_[23];
  assign _zz_1561_ = _zz_1536_[24];
  assign _zz_1562_ = _zz_1536_[25];
  assign _zz_1563_ = _zz_1536_[26];
  assign _zz_1564_ = _zz_1536_[27];
  assign _zz_1565_ = _zz_1536_[28];
  assign _zz_1566_ = _zz_1536_[29];
  assign _zz_1567_ = _zz_1536_[30];
  assign _zz_1568_ = _zz_1536_[31];
  assign _zz_1569_ = _zz_1536_[32];
  assign _zz_1570_ = _zz_1536_[33];
  assign _zz_1571_ = _zz_1536_[34];
  assign _zz_1572_ = _zz_1536_[35];
  assign _zz_1573_ = _zz_1536_[36];
  assign _zz_1574_ = _zz_1536_[37];
  assign _zz_1575_ = _zz_1536_[38];
  assign _zz_1576_ = _zz_1536_[39];
  assign _zz_1577_ = _zz_1536_[40];
  assign _zz_1578_ = _zz_1536_[41];
  assign _zz_1579_ = _zz_1536_[42];
  assign _zz_1580_ = _zz_1536_[43];
  assign _zz_1581_ = _zz_1536_[44];
  assign _zz_1582_ = _zz_1536_[45];
  assign _zz_1583_ = _zz_1536_[46];
  assign _zz_1584_ = _zz_1536_[47];
  assign _zz_1585_ = _zz_1536_[48];
  assign _zz_1586_ = _zz_1536_[49];
  assign _zz_1587_ = _zz_1536_[50];
  assign _zz_1588_ = _zz_1536_[51];
  assign _zz_1589_ = _zz_1536_[52];
  assign _zz_1590_ = _zz_1536_[53];
  assign _zz_1591_ = _zz_1536_[54];
  assign _zz_1592_ = _zz_1536_[55];
  assign _zz_1593_ = _zz_1536_[56];
  assign _zz_1594_ = _zz_1536_[57];
  assign _zz_1595_ = _zz_1536_[58];
  assign _zz_1596_ = _zz_1536_[59];
  assign _zz_1597_ = _zz_1536_[60];
  assign _zz_1598_ = _zz_1536_[61];
  assign _zz_1599_ = _zz_1536_[62];
  assign _zz_1600_ = _zz_1536_[63];
  assign _zz_1601_ = (((32'h00000d80 <= load_data_area_current_addr) && (load_data_area_current_addr < 32'h00000dc0)) ? _zz_9__regNext : {_zz_4478_,_zz_4479_});
  assign _zz_1602_ = _zz_1601_[15 : 0];
  assign _zz_1603_ = _zz_1601_[31 : 16];
  assign _zz_1604_ = _zz_4589_[5:0];
  assign _zz_1605_ = ({63'd0,(1'b1)} <<< _zz_1604_);
  assign _zz_1606_ = _zz_1605_[0];
  assign _zz_1607_ = _zz_1605_[1];
  assign _zz_1608_ = _zz_1605_[2];
  assign _zz_1609_ = _zz_1605_[3];
  assign _zz_1610_ = _zz_1605_[4];
  assign _zz_1611_ = _zz_1605_[5];
  assign _zz_1612_ = _zz_1605_[6];
  assign _zz_1613_ = _zz_1605_[7];
  assign _zz_1614_ = _zz_1605_[8];
  assign _zz_1615_ = _zz_1605_[9];
  assign _zz_1616_ = _zz_1605_[10];
  assign _zz_1617_ = _zz_1605_[11];
  assign _zz_1618_ = _zz_1605_[12];
  assign _zz_1619_ = _zz_1605_[13];
  assign _zz_1620_ = _zz_1605_[14];
  assign _zz_1621_ = _zz_1605_[15];
  assign _zz_1622_ = _zz_1605_[16];
  assign _zz_1623_ = _zz_1605_[17];
  assign _zz_1624_ = _zz_1605_[18];
  assign _zz_1625_ = _zz_1605_[19];
  assign _zz_1626_ = _zz_1605_[20];
  assign _zz_1627_ = _zz_1605_[21];
  assign _zz_1628_ = _zz_1605_[22];
  assign _zz_1629_ = _zz_1605_[23];
  assign _zz_1630_ = _zz_1605_[24];
  assign _zz_1631_ = _zz_1605_[25];
  assign _zz_1632_ = _zz_1605_[26];
  assign _zz_1633_ = _zz_1605_[27];
  assign _zz_1634_ = _zz_1605_[28];
  assign _zz_1635_ = _zz_1605_[29];
  assign _zz_1636_ = _zz_1605_[30];
  assign _zz_1637_ = _zz_1605_[31];
  assign _zz_1638_ = _zz_1605_[32];
  assign _zz_1639_ = _zz_1605_[33];
  assign _zz_1640_ = _zz_1605_[34];
  assign _zz_1641_ = _zz_1605_[35];
  assign _zz_1642_ = _zz_1605_[36];
  assign _zz_1643_ = _zz_1605_[37];
  assign _zz_1644_ = _zz_1605_[38];
  assign _zz_1645_ = _zz_1605_[39];
  assign _zz_1646_ = _zz_1605_[40];
  assign _zz_1647_ = _zz_1605_[41];
  assign _zz_1648_ = _zz_1605_[42];
  assign _zz_1649_ = _zz_1605_[43];
  assign _zz_1650_ = _zz_1605_[44];
  assign _zz_1651_ = _zz_1605_[45];
  assign _zz_1652_ = _zz_1605_[46];
  assign _zz_1653_ = _zz_1605_[47];
  assign _zz_1654_ = _zz_1605_[48];
  assign _zz_1655_ = _zz_1605_[49];
  assign _zz_1656_ = _zz_1605_[50];
  assign _zz_1657_ = _zz_1605_[51];
  assign _zz_1658_ = _zz_1605_[52];
  assign _zz_1659_ = _zz_1605_[53];
  assign _zz_1660_ = _zz_1605_[54];
  assign _zz_1661_ = _zz_1605_[55];
  assign _zz_1662_ = _zz_1605_[56];
  assign _zz_1663_ = _zz_1605_[57];
  assign _zz_1664_ = _zz_1605_[58];
  assign _zz_1665_ = _zz_1605_[59];
  assign _zz_1666_ = _zz_1605_[60];
  assign _zz_1667_ = _zz_1605_[61];
  assign _zz_1668_ = _zz_1605_[62];
  assign _zz_1669_ = _zz_1605_[63];
  assign _zz_1670_ = (((32'h00000ac0 <= load_data_area_current_addr) && (load_data_area_current_addr < 32'h00000b00)) ? _zz_9__regNext : {_zz_4480_,_zz_4481_});
  assign _zz_1671_ = _zz_1670_[15 : 0];
  assign _zz_1672_ = _zz_1670_[31 : 16];
  assign _zz_1673_ = _zz_4590_[5:0];
  assign _zz_1674_ = ({63'd0,(1'b1)} <<< _zz_1673_);
  assign _zz_1675_ = _zz_1674_[0];
  assign _zz_1676_ = _zz_1674_[1];
  assign _zz_1677_ = _zz_1674_[2];
  assign _zz_1678_ = _zz_1674_[3];
  assign _zz_1679_ = _zz_1674_[4];
  assign _zz_1680_ = _zz_1674_[5];
  assign _zz_1681_ = _zz_1674_[6];
  assign _zz_1682_ = _zz_1674_[7];
  assign _zz_1683_ = _zz_1674_[8];
  assign _zz_1684_ = _zz_1674_[9];
  assign _zz_1685_ = _zz_1674_[10];
  assign _zz_1686_ = _zz_1674_[11];
  assign _zz_1687_ = _zz_1674_[12];
  assign _zz_1688_ = _zz_1674_[13];
  assign _zz_1689_ = _zz_1674_[14];
  assign _zz_1690_ = _zz_1674_[15];
  assign _zz_1691_ = _zz_1674_[16];
  assign _zz_1692_ = _zz_1674_[17];
  assign _zz_1693_ = _zz_1674_[18];
  assign _zz_1694_ = _zz_1674_[19];
  assign _zz_1695_ = _zz_1674_[20];
  assign _zz_1696_ = _zz_1674_[21];
  assign _zz_1697_ = _zz_1674_[22];
  assign _zz_1698_ = _zz_1674_[23];
  assign _zz_1699_ = _zz_1674_[24];
  assign _zz_1700_ = _zz_1674_[25];
  assign _zz_1701_ = _zz_1674_[26];
  assign _zz_1702_ = _zz_1674_[27];
  assign _zz_1703_ = _zz_1674_[28];
  assign _zz_1704_ = _zz_1674_[29];
  assign _zz_1705_ = _zz_1674_[30];
  assign _zz_1706_ = _zz_1674_[31];
  assign _zz_1707_ = _zz_1674_[32];
  assign _zz_1708_ = _zz_1674_[33];
  assign _zz_1709_ = _zz_1674_[34];
  assign _zz_1710_ = _zz_1674_[35];
  assign _zz_1711_ = _zz_1674_[36];
  assign _zz_1712_ = _zz_1674_[37];
  assign _zz_1713_ = _zz_1674_[38];
  assign _zz_1714_ = _zz_1674_[39];
  assign _zz_1715_ = _zz_1674_[40];
  assign _zz_1716_ = _zz_1674_[41];
  assign _zz_1717_ = _zz_1674_[42];
  assign _zz_1718_ = _zz_1674_[43];
  assign _zz_1719_ = _zz_1674_[44];
  assign _zz_1720_ = _zz_1674_[45];
  assign _zz_1721_ = _zz_1674_[46];
  assign _zz_1722_ = _zz_1674_[47];
  assign _zz_1723_ = _zz_1674_[48];
  assign _zz_1724_ = _zz_1674_[49];
  assign _zz_1725_ = _zz_1674_[50];
  assign _zz_1726_ = _zz_1674_[51];
  assign _zz_1727_ = _zz_1674_[52];
  assign _zz_1728_ = _zz_1674_[53];
  assign _zz_1729_ = _zz_1674_[54];
  assign _zz_1730_ = _zz_1674_[55];
  assign _zz_1731_ = _zz_1674_[56];
  assign _zz_1732_ = _zz_1674_[57];
  assign _zz_1733_ = _zz_1674_[58];
  assign _zz_1734_ = _zz_1674_[59];
  assign _zz_1735_ = _zz_1674_[60];
  assign _zz_1736_ = _zz_1674_[61];
  assign _zz_1737_ = _zz_1674_[62];
  assign _zz_1738_ = _zz_1674_[63];
  assign _zz_1739_ = (((32'h00000380 <= load_data_area_current_addr) && (load_data_area_current_addr < 32'h000003c0)) ? _zz_9__regNext : {_zz_4482_,_zz_4483_});
  assign _zz_1740_ = _zz_1739_[15 : 0];
  assign _zz_1741_ = _zz_1739_[31 : 16];
  assign _zz_1742_ = _zz_4591_[5:0];
  assign _zz_1743_ = ({63'd0,(1'b1)} <<< _zz_1742_);
  assign _zz_1744_ = _zz_1743_[0];
  assign _zz_1745_ = _zz_1743_[1];
  assign _zz_1746_ = _zz_1743_[2];
  assign _zz_1747_ = _zz_1743_[3];
  assign _zz_1748_ = _zz_1743_[4];
  assign _zz_1749_ = _zz_1743_[5];
  assign _zz_1750_ = _zz_1743_[6];
  assign _zz_1751_ = _zz_1743_[7];
  assign _zz_1752_ = _zz_1743_[8];
  assign _zz_1753_ = _zz_1743_[9];
  assign _zz_1754_ = _zz_1743_[10];
  assign _zz_1755_ = _zz_1743_[11];
  assign _zz_1756_ = _zz_1743_[12];
  assign _zz_1757_ = _zz_1743_[13];
  assign _zz_1758_ = _zz_1743_[14];
  assign _zz_1759_ = _zz_1743_[15];
  assign _zz_1760_ = _zz_1743_[16];
  assign _zz_1761_ = _zz_1743_[17];
  assign _zz_1762_ = _zz_1743_[18];
  assign _zz_1763_ = _zz_1743_[19];
  assign _zz_1764_ = _zz_1743_[20];
  assign _zz_1765_ = _zz_1743_[21];
  assign _zz_1766_ = _zz_1743_[22];
  assign _zz_1767_ = _zz_1743_[23];
  assign _zz_1768_ = _zz_1743_[24];
  assign _zz_1769_ = _zz_1743_[25];
  assign _zz_1770_ = _zz_1743_[26];
  assign _zz_1771_ = _zz_1743_[27];
  assign _zz_1772_ = _zz_1743_[28];
  assign _zz_1773_ = _zz_1743_[29];
  assign _zz_1774_ = _zz_1743_[30];
  assign _zz_1775_ = _zz_1743_[31];
  assign _zz_1776_ = _zz_1743_[32];
  assign _zz_1777_ = _zz_1743_[33];
  assign _zz_1778_ = _zz_1743_[34];
  assign _zz_1779_ = _zz_1743_[35];
  assign _zz_1780_ = _zz_1743_[36];
  assign _zz_1781_ = _zz_1743_[37];
  assign _zz_1782_ = _zz_1743_[38];
  assign _zz_1783_ = _zz_1743_[39];
  assign _zz_1784_ = _zz_1743_[40];
  assign _zz_1785_ = _zz_1743_[41];
  assign _zz_1786_ = _zz_1743_[42];
  assign _zz_1787_ = _zz_1743_[43];
  assign _zz_1788_ = _zz_1743_[44];
  assign _zz_1789_ = _zz_1743_[45];
  assign _zz_1790_ = _zz_1743_[46];
  assign _zz_1791_ = _zz_1743_[47];
  assign _zz_1792_ = _zz_1743_[48];
  assign _zz_1793_ = _zz_1743_[49];
  assign _zz_1794_ = _zz_1743_[50];
  assign _zz_1795_ = _zz_1743_[51];
  assign _zz_1796_ = _zz_1743_[52];
  assign _zz_1797_ = _zz_1743_[53];
  assign _zz_1798_ = _zz_1743_[54];
  assign _zz_1799_ = _zz_1743_[55];
  assign _zz_1800_ = _zz_1743_[56];
  assign _zz_1801_ = _zz_1743_[57];
  assign _zz_1802_ = _zz_1743_[58];
  assign _zz_1803_ = _zz_1743_[59];
  assign _zz_1804_ = _zz_1743_[60];
  assign _zz_1805_ = _zz_1743_[61];
  assign _zz_1806_ = _zz_1743_[62];
  assign _zz_1807_ = _zz_1743_[63];
  assign _zz_1808_ = (((32'h00000800 <= load_data_area_current_addr) && (load_data_area_current_addr < 32'h00000840)) ? _zz_9__regNext : {_zz_4484_,_zz_4485_});
  assign _zz_1809_ = _zz_1808_[15 : 0];
  assign _zz_1810_ = _zz_1808_[31 : 16];
  assign _zz_1811_ = _zz_4592_[5:0];
  assign _zz_1812_ = ({63'd0,(1'b1)} <<< _zz_1811_);
  assign _zz_1813_ = _zz_1812_[0];
  assign _zz_1814_ = _zz_1812_[1];
  assign _zz_1815_ = _zz_1812_[2];
  assign _zz_1816_ = _zz_1812_[3];
  assign _zz_1817_ = _zz_1812_[4];
  assign _zz_1818_ = _zz_1812_[5];
  assign _zz_1819_ = _zz_1812_[6];
  assign _zz_1820_ = _zz_1812_[7];
  assign _zz_1821_ = _zz_1812_[8];
  assign _zz_1822_ = _zz_1812_[9];
  assign _zz_1823_ = _zz_1812_[10];
  assign _zz_1824_ = _zz_1812_[11];
  assign _zz_1825_ = _zz_1812_[12];
  assign _zz_1826_ = _zz_1812_[13];
  assign _zz_1827_ = _zz_1812_[14];
  assign _zz_1828_ = _zz_1812_[15];
  assign _zz_1829_ = _zz_1812_[16];
  assign _zz_1830_ = _zz_1812_[17];
  assign _zz_1831_ = _zz_1812_[18];
  assign _zz_1832_ = _zz_1812_[19];
  assign _zz_1833_ = _zz_1812_[20];
  assign _zz_1834_ = _zz_1812_[21];
  assign _zz_1835_ = _zz_1812_[22];
  assign _zz_1836_ = _zz_1812_[23];
  assign _zz_1837_ = _zz_1812_[24];
  assign _zz_1838_ = _zz_1812_[25];
  assign _zz_1839_ = _zz_1812_[26];
  assign _zz_1840_ = _zz_1812_[27];
  assign _zz_1841_ = _zz_1812_[28];
  assign _zz_1842_ = _zz_1812_[29];
  assign _zz_1843_ = _zz_1812_[30];
  assign _zz_1844_ = _zz_1812_[31];
  assign _zz_1845_ = _zz_1812_[32];
  assign _zz_1846_ = _zz_1812_[33];
  assign _zz_1847_ = _zz_1812_[34];
  assign _zz_1848_ = _zz_1812_[35];
  assign _zz_1849_ = _zz_1812_[36];
  assign _zz_1850_ = _zz_1812_[37];
  assign _zz_1851_ = _zz_1812_[38];
  assign _zz_1852_ = _zz_1812_[39];
  assign _zz_1853_ = _zz_1812_[40];
  assign _zz_1854_ = _zz_1812_[41];
  assign _zz_1855_ = _zz_1812_[42];
  assign _zz_1856_ = _zz_1812_[43];
  assign _zz_1857_ = _zz_1812_[44];
  assign _zz_1858_ = _zz_1812_[45];
  assign _zz_1859_ = _zz_1812_[46];
  assign _zz_1860_ = _zz_1812_[47];
  assign _zz_1861_ = _zz_1812_[48];
  assign _zz_1862_ = _zz_1812_[49];
  assign _zz_1863_ = _zz_1812_[50];
  assign _zz_1864_ = _zz_1812_[51];
  assign _zz_1865_ = _zz_1812_[52];
  assign _zz_1866_ = _zz_1812_[53];
  assign _zz_1867_ = _zz_1812_[54];
  assign _zz_1868_ = _zz_1812_[55];
  assign _zz_1869_ = _zz_1812_[56];
  assign _zz_1870_ = _zz_1812_[57];
  assign _zz_1871_ = _zz_1812_[58];
  assign _zz_1872_ = _zz_1812_[59];
  assign _zz_1873_ = _zz_1812_[60];
  assign _zz_1874_ = _zz_1812_[61];
  assign _zz_1875_ = _zz_1812_[62];
  assign _zz_1876_ = _zz_1812_[63];
  assign _zz_1877_ = (((32'h00000f40 <= load_data_area_current_addr) && (load_data_area_current_addr < 32'h00000f80)) ? _zz_9__regNext : {_zz_4486_,_zz_4487_});
  assign _zz_1878_ = _zz_1877_[15 : 0];
  assign _zz_1879_ = _zz_1877_[31 : 16];
  assign _zz_1880_ = _zz_4593_[5:0];
  assign _zz_1881_ = ({63'd0,(1'b1)} <<< _zz_1880_);
  assign _zz_1882_ = _zz_1881_[0];
  assign _zz_1883_ = _zz_1881_[1];
  assign _zz_1884_ = _zz_1881_[2];
  assign _zz_1885_ = _zz_1881_[3];
  assign _zz_1886_ = _zz_1881_[4];
  assign _zz_1887_ = _zz_1881_[5];
  assign _zz_1888_ = _zz_1881_[6];
  assign _zz_1889_ = _zz_1881_[7];
  assign _zz_1890_ = _zz_1881_[8];
  assign _zz_1891_ = _zz_1881_[9];
  assign _zz_1892_ = _zz_1881_[10];
  assign _zz_1893_ = _zz_1881_[11];
  assign _zz_1894_ = _zz_1881_[12];
  assign _zz_1895_ = _zz_1881_[13];
  assign _zz_1896_ = _zz_1881_[14];
  assign _zz_1897_ = _zz_1881_[15];
  assign _zz_1898_ = _zz_1881_[16];
  assign _zz_1899_ = _zz_1881_[17];
  assign _zz_1900_ = _zz_1881_[18];
  assign _zz_1901_ = _zz_1881_[19];
  assign _zz_1902_ = _zz_1881_[20];
  assign _zz_1903_ = _zz_1881_[21];
  assign _zz_1904_ = _zz_1881_[22];
  assign _zz_1905_ = _zz_1881_[23];
  assign _zz_1906_ = _zz_1881_[24];
  assign _zz_1907_ = _zz_1881_[25];
  assign _zz_1908_ = _zz_1881_[26];
  assign _zz_1909_ = _zz_1881_[27];
  assign _zz_1910_ = _zz_1881_[28];
  assign _zz_1911_ = _zz_1881_[29];
  assign _zz_1912_ = _zz_1881_[30];
  assign _zz_1913_ = _zz_1881_[31];
  assign _zz_1914_ = _zz_1881_[32];
  assign _zz_1915_ = _zz_1881_[33];
  assign _zz_1916_ = _zz_1881_[34];
  assign _zz_1917_ = _zz_1881_[35];
  assign _zz_1918_ = _zz_1881_[36];
  assign _zz_1919_ = _zz_1881_[37];
  assign _zz_1920_ = _zz_1881_[38];
  assign _zz_1921_ = _zz_1881_[39];
  assign _zz_1922_ = _zz_1881_[40];
  assign _zz_1923_ = _zz_1881_[41];
  assign _zz_1924_ = _zz_1881_[42];
  assign _zz_1925_ = _zz_1881_[43];
  assign _zz_1926_ = _zz_1881_[44];
  assign _zz_1927_ = _zz_1881_[45];
  assign _zz_1928_ = _zz_1881_[46];
  assign _zz_1929_ = _zz_1881_[47];
  assign _zz_1930_ = _zz_1881_[48];
  assign _zz_1931_ = _zz_1881_[49];
  assign _zz_1932_ = _zz_1881_[50];
  assign _zz_1933_ = _zz_1881_[51];
  assign _zz_1934_ = _zz_1881_[52];
  assign _zz_1935_ = _zz_1881_[53];
  assign _zz_1936_ = _zz_1881_[54];
  assign _zz_1937_ = _zz_1881_[55];
  assign _zz_1938_ = _zz_1881_[56];
  assign _zz_1939_ = _zz_1881_[57];
  assign _zz_1940_ = _zz_1881_[58];
  assign _zz_1941_ = _zz_1881_[59];
  assign _zz_1942_ = _zz_1881_[60];
  assign _zz_1943_ = _zz_1881_[61];
  assign _zz_1944_ = _zz_1881_[62];
  assign _zz_1945_ = _zz_1881_[63];
  assign _zz_1946_ = (((32'h00000680 <= load_data_area_current_addr) && (load_data_area_current_addr < 32'h000006c0)) ? _zz_9__regNext : {_zz_4488_,_zz_4489_});
  assign _zz_1947_ = _zz_1946_[15 : 0];
  assign _zz_1948_ = _zz_1946_[31 : 16];
  assign _zz_1949_ = _zz_4594_[5:0];
  assign _zz_1950_ = ({63'd0,(1'b1)} <<< _zz_1949_);
  assign _zz_1951_ = _zz_1950_[0];
  assign _zz_1952_ = _zz_1950_[1];
  assign _zz_1953_ = _zz_1950_[2];
  assign _zz_1954_ = _zz_1950_[3];
  assign _zz_1955_ = _zz_1950_[4];
  assign _zz_1956_ = _zz_1950_[5];
  assign _zz_1957_ = _zz_1950_[6];
  assign _zz_1958_ = _zz_1950_[7];
  assign _zz_1959_ = _zz_1950_[8];
  assign _zz_1960_ = _zz_1950_[9];
  assign _zz_1961_ = _zz_1950_[10];
  assign _zz_1962_ = _zz_1950_[11];
  assign _zz_1963_ = _zz_1950_[12];
  assign _zz_1964_ = _zz_1950_[13];
  assign _zz_1965_ = _zz_1950_[14];
  assign _zz_1966_ = _zz_1950_[15];
  assign _zz_1967_ = _zz_1950_[16];
  assign _zz_1968_ = _zz_1950_[17];
  assign _zz_1969_ = _zz_1950_[18];
  assign _zz_1970_ = _zz_1950_[19];
  assign _zz_1971_ = _zz_1950_[20];
  assign _zz_1972_ = _zz_1950_[21];
  assign _zz_1973_ = _zz_1950_[22];
  assign _zz_1974_ = _zz_1950_[23];
  assign _zz_1975_ = _zz_1950_[24];
  assign _zz_1976_ = _zz_1950_[25];
  assign _zz_1977_ = _zz_1950_[26];
  assign _zz_1978_ = _zz_1950_[27];
  assign _zz_1979_ = _zz_1950_[28];
  assign _zz_1980_ = _zz_1950_[29];
  assign _zz_1981_ = _zz_1950_[30];
  assign _zz_1982_ = _zz_1950_[31];
  assign _zz_1983_ = _zz_1950_[32];
  assign _zz_1984_ = _zz_1950_[33];
  assign _zz_1985_ = _zz_1950_[34];
  assign _zz_1986_ = _zz_1950_[35];
  assign _zz_1987_ = _zz_1950_[36];
  assign _zz_1988_ = _zz_1950_[37];
  assign _zz_1989_ = _zz_1950_[38];
  assign _zz_1990_ = _zz_1950_[39];
  assign _zz_1991_ = _zz_1950_[40];
  assign _zz_1992_ = _zz_1950_[41];
  assign _zz_1993_ = _zz_1950_[42];
  assign _zz_1994_ = _zz_1950_[43];
  assign _zz_1995_ = _zz_1950_[44];
  assign _zz_1996_ = _zz_1950_[45];
  assign _zz_1997_ = _zz_1950_[46];
  assign _zz_1998_ = _zz_1950_[47];
  assign _zz_1999_ = _zz_1950_[48];
  assign _zz_2000_ = _zz_1950_[49];
  assign _zz_2001_ = _zz_1950_[50];
  assign _zz_2002_ = _zz_1950_[51];
  assign _zz_2003_ = _zz_1950_[52];
  assign _zz_2004_ = _zz_1950_[53];
  assign _zz_2005_ = _zz_1950_[54];
  assign _zz_2006_ = _zz_1950_[55];
  assign _zz_2007_ = _zz_1950_[56];
  assign _zz_2008_ = _zz_1950_[57];
  assign _zz_2009_ = _zz_1950_[58];
  assign _zz_2010_ = _zz_1950_[59];
  assign _zz_2011_ = _zz_1950_[60];
  assign _zz_2012_ = _zz_1950_[61];
  assign _zz_2013_ = _zz_1950_[62];
  assign _zz_2014_ = _zz_1950_[63];
  assign _zz_2015_ = (((32'h00000400 <= load_data_area_current_addr) && (load_data_area_current_addr < 32'h00000440)) ? _zz_9__regNext : {_zz_4490_,_zz_4491_});
  assign _zz_2016_ = _zz_2015_[15 : 0];
  assign _zz_2017_ = _zz_2015_[31 : 16];
  assign _zz_2018_ = _zz_4595_[5:0];
  assign _zz_2019_ = ({63'd0,(1'b1)} <<< _zz_2018_);
  assign _zz_2020_ = _zz_2019_[0];
  assign _zz_2021_ = _zz_2019_[1];
  assign _zz_2022_ = _zz_2019_[2];
  assign _zz_2023_ = _zz_2019_[3];
  assign _zz_2024_ = _zz_2019_[4];
  assign _zz_2025_ = _zz_2019_[5];
  assign _zz_2026_ = _zz_2019_[6];
  assign _zz_2027_ = _zz_2019_[7];
  assign _zz_2028_ = _zz_2019_[8];
  assign _zz_2029_ = _zz_2019_[9];
  assign _zz_2030_ = _zz_2019_[10];
  assign _zz_2031_ = _zz_2019_[11];
  assign _zz_2032_ = _zz_2019_[12];
  assign _zz_2033_ = _zz_2019_[13];
  assign _zz_2034_ = _zz_2019_[14];
  assign _zz_2035_ = _zz_2019_[15];
  assign _zz_2036_ = _zz_2019_[16];
  assign _zz_2037_ = _zz_2019_[17];
  assign _zz_2038_ = _zz_2019_[18];
  assign _zz_2039_ = _zz_2019_[19];
  assign _zz_2040_ = _zz_2019_[20];
  assign _zz_2041_ = _zz_2019_[21];
  assign _zz_2042_ = _zz_2019_[22];
  assign _zz_2043_ = _zz_2019_[23];
  assign _zz_2044_ = _zz_2019_[24];
  assign _zz_2045_ = _zz_2019_[25];
  assign _zz_2046_ = _zz_2019_[26];
  assign _zz_2047_ = _zz_2019_[27];
  assign _zz_2048_ = _zz_2019_[28];
  assign _zz_2049_ = _zz_2019_[29];
  assign _zz_2050_ = _zz_2019_[30];
  assign _zz_2051_ = _zz_2019_[31];
  assign _zz_2052_ = _zz_2019_[32];
  assign _zz_2053_ = _zz_2019_[33];
  assign _zz_2054_ = _zz_2019_[34];
  assign _zz_2055_ = _zz_2019_[35];
  assign _zz_2056_ = _zz_2019_[36];
  assign _zz_2057_ = _zz_2019_[37];
  assign _zz_2058_ = _zz_2019_[38];
  assign _zz_2059_ = _zz_2019_[39];
  assign _zz_2060_ = _zz_2019_[40];
  assign _zz_2061_ = _zz_2019_[41];
  assign _zz_2062_ = _zz_2019_[42];
  assign _zz_2063_ = _zz_2019_[43];
  assign _zz_2064_ = _zz_2019_[44];
  assign _zz_2065_ = _zz_2019_[45];
  assign _zz_2066_ = _zz_2019_[46];
  assign _zz_2067_ = _zz_2019_[47];
  assign _zz_2068_ = _zz_2019_[48];
  assign _zz_2069_ = _zz_2019_[49];
  assign _zz_2070_ = _zz_2019_[50];
  assign _zz_2071_ = _zz_2019_[51];
  assign _zz_2072_ = _zz_2019_[52];
  assign _zz_2073_ = _zz_2019_[53];
  assign _zz_2074_ = _zz_2019_[54];
  assign _zz_2075_ = _zz_2019_[55];
  assign _zz_2076_ = _zz_2019_[56];
  assign _zz_2077_ = _zz_2019_[57];
  assign _zz_2078_ = _zz_2019_[58];
  assign _zz_2079_ = _zz_2019_[59];
  assign _zz_2080_ = _zz_2019_[60];
  assign _zz_2081_ = _zz_2019_[61];
  assign _zz_2082_ = _zz_2019_[62];
  assign _zz_2083_ = _zz_2019_[63];
  assign _zz_2084_ = (((32'h00000980 <= load_data_area_current_addr) && (load_data_area_current_addr < 32'h000009c0)) ? _zz_9__regNext : {_zz_4492_,_zz_4493_});
  assign _zz_2085_ = _zz_2084_[15 : 0];
  assign _zz_2086_ = _zz_2084_[31 : 16];
  assign _zz_2087_ = _zz_4596_[5:0];
  assign _zz_2088_ = ({63'd0,(1'b1)} <<< _zz_2087_);
  assign _zz_2089_ = _zz_2088_[0];
  assign _zz_2090_ = _zz_2088_[1];
  assign _zz_2091_ = _zz_2088_[2];
  assign _zz_2092_ = _zz_2088_[3];
  assign _zz_2093_ = _zz_2088_[4];
  assign _zz_2094_ = _zz_2088_[5];
  assign _zz_2095_ = _zz_2088_[6];
  assign _zz_2096_ = _zz_2088_[7];
  assign _zz_2097_ = _zz_2088_[8];
  assign _zz_2098_ = _zz_2088_[9];
  assign _zz_2099_ = _zz_2088_[10];
  assign _zz_2100_ = _zz_2088_[11];
  assign _zz_2101_ = _zz_2088_[12];
  assign _zz_2102_ = _zz_2088_[13];
  assign _zz_2103_ = _zz_2088_[14];
  assign _zz_2104_ = _zz_2088_[15];
  assign _zz_2105_ = _zz_2088_[16];
  assign _zz_2106_ = _zz_2088_[17];
  assign _zz_2107_ = _zz_2088_[18];
  assign _zz_2108_ = _zz_2088_[19];
  assign _zz_2109_ = _zz_2088_[20];
  assign _zz_2110_ = _zz_2088_[21];
  assign _zz_2111_ = _zz_2088_[22];
  assign _zz_2112_ = _zz_2088_[23];
  assign _zz_2113_ = _zz_2088_[24];
  assign _zz_2114_ = _zz_2088_[25];
  assign _zz_2115_ = _zz_2088_[26];
  assign _zz_2116_ = _zz_2088_[27];
  assign _zz_2117_ = _zz_2088_[28];
  assign _zz_2118_ = _zz_2088_[29];
  assign _zz_2119_ = _zz_2088_[30];
  assign _zz_2120_ = _zz_2088_[31];
  assign _zz_2121_ = _zz_2088_[32];
  assign _zz_2122_ = _zz_2088_[33];
  assign _zz_2123_ = _zz_2088_[34];
  assign _zz_2124_ = _zz_2088_[35];
  assign _zz_2125_ = _zz_2088_[36];
  assign _zz_2126_ = _zz_2088_[37];
  assign _zz_2127_ = _zz_2088_[38];
  assign _zz_2128_ = _zz_2088_[39];
  assign _zz_2129_ = _zz_2088_[40];
  assign _zz_2130_ = _zz_2088_[41];
  assign _zz_2131_ = _zz_2088_[42];
  assign _zz_2132_ = _zz_2088_[43];
  assign _zz_2133_ = _zz_2088_[44];
  assign _zz_2134_ = _zz_2088_[45];
  assign _zz_2135_ = _zz_2088_[46];
  assign _zz_2136_ = _zz_2088_[47];
  assign _zz_2137_ = _zz_2088_[48];
  assign _zz_2138_ = _zz_2088_[49];
  assign _zz_2139_ = _zz_2088_[50];
  assign _zz_2140_ = _zz_2088_[51];
  assign _zz_2141_ = _zz_2088_[52];
  assign _zz_2142_ = _zz_2088_[53];
  assign _zz_2143_ = _zz_2088_[54];
  assign _zz_2144_ = _zz_2088_[55];
  assign _zz_2145_ = _zz_2088_[56];
  assign _zz_2146_ = _zz_2088_[57];
  assign _zz_2147_ = _zz_2088_[58];
  assign _zz_2148_ = _zz_2088_[59];
  assign _zz_2149_ = _zz_2088_[60];
  assign _zz_2150_ = _zz_2088_[61];
  assign _zz_2151_ = _zz_2088_[62];
  assign _zz_2152_ = _zz_2088_[63];
  assign _zz_2153_ = (((32'h00000e00 <= load_data_area_current_addr) && (load_data_area_current_addr < 32'h00000e40)) ? _zz_9__regNext : {_zz_4494_,_zz_4495_});
  assign _zz_2154_ = _zz_2153_[15 : 0];
  assign _zz_2155_ = _zz_2153_[31 : 16];
  assign _zz_2156_ = _zz_4597_[5:0];
  assign _zz_2157_ = ({63'd0,(1'b1)} <<< _zz_2156_);
  assign _zz_2158_ = _zz_2157_[0];
  assign _zz_2159_ = _zz_2157_[1];
  assign _zz_2160_ = _zz_2157_[2];
  assign _zz_2161_ = _zz_2157_[3];
  assign _zz_2162_ = _zz_2157_[4];
  assign _zz_2163_ = _zz_2157_[5];
  assign _zz_2164_ = _zz_2157_[6];
  assign _zz_2165_ = _zz_2157_[7];
  assign _zz_2166_ = _zz_2157_[8];
  assign _zz_2167_ = _zz_2157_[9];
  assign _zz_2168_ = _zz_2157_[10];
  assign _zz_2169_ = _zz_2157_[11];
  assign _zz_2170_ = _zz_2157_[12];
  assign _zz_2171_ = _zz_2157_[13];
  assign _zz_2172_ = _zz_2157_[14];
  assign _zz_2173_ = _zz_2157_[15];
  assign _zz_2174_ = _zz_2157_[16];
  assign _zz_2175_ = _zz_2157_[17];
  assign _zz_2176_ = _zz_2157_[18];
  assign _zz_2177_ = _zz_2157_[19];
  assign _zz_2178_ = _zz_2157_[20];
  assign _zz_2179_ = _zz_2157_[21];
  assign _zz_2180_ = _zz_2157_[22];
  assign _zz_2181_ = _zz_2157_[23];
  assign _zz_2182_ = _zz_2157_[24];
  assign _zz_2183_ = _zz_2157_[25];
  assign _zz_2184_ = _zz_2157_[26];
  assign _zz_2185_ = _zz_2157_[27];
  assign _zz_2186_ = _zz_2157_[28];
  assign _zz_2187_ = _zz_2157_[29];
  assign _zz_2188_ = _zz_2157_[30];
  assign _zz_2189_ = _zz_2157_[31];
  assign _zz_2190_ = _zz_2157_[32];
  assign _zz_2191_ = _zz_2157_[33];
  assign _zz_2192_ = _zz_2157_[34];
  assign _zz_2193_ = _zz_2157_[35];
  assign _zz_2194_ = _zz_2157_[36];
  assign _zz_2195_ = _zz_2157_[37];
  assign _zz_2196_ = _zz_2157_[38];
  assign _zz_2197_ = _zz_2157_[39];
  assign _zz_2198_ = _zz_2157_[40];
  assign _zz_2199_ = _zz_2157_[41];
  assign _zz_2200_ = _zz_2157_[42];
  assign _zz_2201_ = _zz_2157_[43];
  assign _zz_2202_ = _zz_2157_[44];
  assign _zz_2203_ = _zz_2157_[45];
  assign _zz_2204_ = _zz_2157_[46];
  assign _zz_2205_ = _zz_2157_[47];
  assign _zz_2206_ = _zz_2157_[48];
  assign _zz_2207_ = _zz_2157_[49];
  assign _zz_2208_ = _zz_2157_[50];
  assign _zz_2209_ = _zz_2157_[51];
  assign _zz_2210_ = _zz_2157_[52];
  assign _zz_2211_ = _zz_2157_[53];
  assign _zz_2212_ = _zz_2157_[54];
  assign _zz_2213_ = _zz_2157_[55];
  assign _zz_2214_ = _zz_2157_[56];
  assign _zz_2215_ = _zz_2157_[57];
  assign _zz_2216_ = _zz_2157_[58];
  assign _zz_2217_ = _zz_2157_[59];
  assign _zz_2218_ = _zz_2157_[60];
  assign _zz_2219_ = _zz_2157_[61];
  assign _zz_2220_ = _zz_2157_[62];
  assign _zz_2221_ = _zz_2157_[63];
  assign _zz_2222_ = (((32'h00000e40 <= load_data_area_current_addr) && (load_data_area_current_addr < 32'h00000e80)) ? _zz_9__regNext : {_zz_4496_,_zz_4497_});
  assign _zz_2223_ = _zz_2222_[15 : 0];
  assign _zz_2224_ = _zz_2222_[31 : 16];
  assign _zz_2225_ = _zz_4598_[5:0];
  assign _zz_2226_ = ({63'd0,(1'b1)} <<< _zz_2225_);
  assign _zz_2227_ = _zz_2226_[0];
  assign _zz_2228_ = _zz_2226_[1];
  assign _zz_2229_ = _zz_2226_[2];
  assign _zz_2230_ = _zz_2226_[3];
  assign _zz_2231_ = _zz_2226_[4];
  assign _zz_2232_ = _zz_2226_[5];
  assign _zz_2233_ = _zz_2226_[6];
  assign _zz_2234_ = _zz_2226_[7];
  assign _zz_2235_ = _zz_2226_[8];
  assign _zz_2236_ = _zz_2226_[9];
  assign _zz_2237_ = _zz_2226_[10];
  assign _zz_2238_ = _zz_2226_[11];
  assign _zz_2239_ = _zz_2226_[12];
  assign _zz_2240_ = _zz_2226_[13];
  assign _zz_2241_ = _zz_2226_[14];
  assign _zz_2242_ = _zz_2226_[15];
  assign _zz_2243_ = _zz_2226_[16];
  assign _zz_2244_ = _zz_2226_[17];
  assign _zz_2245_ = _zz_2226_[18];
  assign _zz_2246_ = _zz_2226_[19];
  assign _zz_2247_ = _zz_2226_[20];
  assign _zz_2248_ = _zz_2226_[21];
  assign _zz_2249_ = _zz_2226_[22];
  assign _zz_2250_ = _zz_2226_[23];
  assign _zz_2251_ = _zz_2226_[24];
  assign _zz_2252_ = _zz_2226_[25];
  assign _zz_2253_ = _zz_2226_[26];
  assign _zz_2254_ = _zz_2226_[27];
  assign _zz_2255_ = _zz_2226_[28];
  assign _zz_2256_ = _zz_2226_[29];
  assign _zz_2257_ = _zz_2226_[30];
  assign _zz_2258_ = _zz_2226_[31];
  assign _zz_2259_ = _zz_2226_[32];
  assign _zz_2260_ = _zz_2226_[33];
  assign _zz_2261_ = _zz_2226_[34];
  assign _zz_2262_ = _zz_2226_[35];
  assign _zz_2263_ = _zz_2226_[36];
  assign _zz_2264_ = _zz_2226_[37];
  assign _zz_2265_ = _zz_2226_[38];
  assign _zz_2266_ = _zz_2226_[39];
  assign _zz_2267_ = _zz_2226_[40];
  assign _zz_2268_ = _zz_2226_[41];
  assign _zz_2269_ = _zz_2226_[42];
  assign _zz_2270_ = _zz_2226_[43];
  assign _zz_2271_ = _zz_2226_[44];
  assign _zz_2272_ = _zz_2226_[45];
  assign _zz_2273_ = _zz_2226_[46];
  assign _zz_2274_ = _zz_2226_[47];
  assign _zz_2275_ = _zz_2226_[48];
  assign _zz_2276_ = _zz_2226_[49];
  assign _zz_2277_ = _zz_2226_[50];
  assign _zz_2278_ = _zz_2226_[51];
  assign _zz_2279_ = _zz_2226_[52];
  assign _zz_2280_ = _zz_2226_[53];
  assign _zz_2281_ = _zz_2226_[54];
  assign _zz_2282_ = _zz_2226_[55];
  assign _zz_2283_ = _zz_2226_[56];
  assign _zz_2284_ = _zz_2226_[57];
  assign _zz_2285_ = _zz_2226_[58];
  assign _zz_2286_ = _zz_2226_[59];
  assign _zz_2287_ = _zz_2226_[60];
  assign _zz_2288_ = _zz_2226_[61];
  assign _zz_2289_ = _zz_2226_[62];
  assign _zz_2290_ = _zz_2226_[63];
  assign _zz_2291_ = (((32'h00000600 <= load_data_area_current_addr) && (load_data_area_current_addr < 32'h00000640)) ? _zz_9__regNext : {_zz_4498_,_zz_4499_});
  assign _zz_2292_ = _zz_2291_[15 : 0];
  assign _zz_2293_ = _zz_2291_[31 : 16];
  assign _zz_2294_ = _zz_4599_[5:0];
  assign _zz_2295_ = ({63'd0,(1'b1)} <<< _zz_2294_);
  assign _zz_2296_ = _zz_2295_[0];
  assign _zz_2297_ = _zz_2295_[1];
  assign _zz_2298_ = _zz_2295_[2];
  assign _zz_2299_ = _zz_2295_[3];
  assign _zz_2300_ = _zz_2295_[4];
  assign _zz_2301_ = _zz_2295_[5];
  assign _zz_2302_ = _zz_2295_[6];
  assign _zz_2303_ = _zz_2295_[7];
  assign _zz_2304_ = _zz_2295_[8];
  assign _zz_2305_ = _zz_2295_[9];
  assign _zz_2306_ = _zz_2295_[10];
  assign _zz_2307_ = _zz_2295_[11];
  assign _zz_2308_ = _zz_2295_[12];
  assign _zz_2309_ = _zz_2295_[13];
  assign _zz_2310_ = _zz_2295_[14];
  assign _zz_2311_ = _zz_2295_[15];
  assign _zz_2312_ = _zz_2295_[16];
  assign _zz_2313_ = _zz_2295_[17];
  assign _zz_2314_ = _zz_2295_[18];
  assign _zz_2315_ = _zz_2295_[19];
  assign _zz_2316_ = _zz_2295_[20];
  assign _zz_2317_ = _zz_2295_[21];
  assign _zz_2318_ = _zz_2295_[22];
  assign _zz_2319_ = _zz_2295_[23];
  assign _zz_2320_ = _zz_2295_[24];
  assign _zz_2321_ = _zz_2295_[25];
  assign _zz_2322_ = _zz_2295_[26];
  assign _zz_2323_ = _zz_2295_[27];
  assign _zz_2324_ = _zz_2295_[28];
  assign _zz_2325_ = _zz_2295_[29];
  assign _zz_2326_ = _zz_2295_[30];
  assign _zz_2327_ = _zz_2295_[31];
  assign _zz_2328_ = _zz_2295_[32];
  assign _zz_2329_ = _zz_2295_[33];
  assign _zz_2330_ = _zz_2295_[34];
  assign _zz_2331_ = _zz_2295_[35];
  assign _zz_2332_ = _zz_2295_[36];
  assign _zz_2333_ = _zz_2295_[37];
  assign _zz_2334_ = _zz_2295_[38];
  assign _zz_2335_ = _zz_2295_[39];
  assign _zz_2336_ = _zz_2295_[40];
  assign _zz_2337_ = _zz_2295_[41];
  assign _zz_2338_ = _zz_2295_[42];
  assign _zz_2339_ = _zz_2295_[43];
  assign _zz_2340_ = _zz_2295_[44];
  assign _zz_2341_ = _zz_2295_[45];
  assign _zz_2342_ = _zz_2295_[46];
  assign _zz_2343_ = _zz_2295_[47];
  assign _zz_2344_ = _zz_2295_[48];
  assign _zz_2345_ = _zz_2295_[49];
  assign _zz_2346_ = _zz_2295_[50];
  assign _zz_2347_ = _zz_2295_[51];
  assign _zz_2348_ = _zz_2295_[52];
  assign _zz_2349_ = _zz_2295_[53];
  assign _zz_2350_ = _zz_2295_[54];
  assign _zz_2351_ = _zz_2295_[55];
  assign _zz_2352_ = _zz_2295_[56];
  assign _zz_2353_ = _zz_2295_[57];
  assign _zz_2354_ = _zz_2295_[58];
  assign _zz_2355_ = _zz_2295_[59];
  assign _zz_2356_ = _zz_2295_[60];
  assign _zz_2357_ = _zz_2295_[61];
  assign _zz_2358_ = _zz_2295_[62];
  assign _zz_2359_ = _zz_2295_[63];
  assign _zz_2360_ = (((32'h00000040 <= load_data_area_current_addr) && (load_data_area_current_addr < 32'h00000080)) ? _zz_9__regNext : {_zz_4500_,_zz_4501_});
  assign _zz_2361_ = _zz_2360_[15 : 0];
  assign _zz_2362_ = _zz_2360_[31 : 16];
  assign _zz_2363_ = _zz_4600_[5:0];
  assign _zz_2364_ = ({63'd0,(1'b1)} <<< _zz_2363_);
  assign _zz_2365_ = _zz_2364_[0];
  assign _zz_2366_ = _zz_2364_[1];
  assign _zz_2367_ = _zz_2364_[2];
  assign _zz_2368_ = _zz_2364_[3];
  assign _zz_2369_ = _zz_2364_[4];
  assign _zz_2370_ = _zz_2364_[5];
  assign _zz_2371_ = _zz_2364_[6];
  assign _zz_2372_ = _zz_2364_[7];
  assign _zz_2373_ = _zz_2364_[8];
  assign _zz_2374_ = _zz_2364_[9];
  assign _zz_2375_ = _zz_2364_[10];
  assign _zz_2376_ = _zz_2364_[11];
  assign _zz_2377_ = _zz_2364_[12];
  assign _zz_2378_ = _zz_2364_[13];
  assign _zz_2379_ = _zz_2364_[14];
  assign _zz_2380_ = _zz_2364_[15];
  assign _zz_2381_ = _zz_2364_[16];
  assign _zz_2382_ = _zz_2364_[17];
  assign _zz_2383_ = _zz_2364_[18];
  assign _zz_2384_ = _zz_2364_[19];
  assign _zz_2385_ = _zz_2364_[20];
  assign _zz_2386_ = _zz_2364_[21];
  assign _zz_2387_ = _zz_2364_[22];
  assign _zz_2388_ = _zz_2364_[23];
  assign _zz_2389_ = _zz_2364_[24];
  assign _zz_2390_ = _zz_2364_[25];
  assign _zz_2391_ = _zz_2364_[26];
  assign _zz_2392_ = _zz_2364_[27];
  assign _zz_2393_ = _zz_2364_[28];
  assign _zz_2394_ = _zz_2364_[29];
  assign _zz_2395_ = _zz_2364_[30];
  assign _zz_2396_ = _zz_2364_[31];
  assign _zz_2397_ = _zz_2364_[32];
  assign _zz_2398_ = _zz_2364_[33];
  assign _zz_2399_ = _zz_2364_[34];
  assign _zz_2400_ = _zz_2364_[35];
  assign _zz_2401_ = _zz_2364_[36];
  assign _zz_2402_ = _zz_2364_[37];
  assign _zz_2403_ = _zz_2364_[38];
  assign _zz_2404_ = _zz_2364_[39];
  assign _zz_2405_ = _zz_2364_[40];
  assign _zz_2406_ = _zz_2364_[41];
  assign _zz_2407_ = _zz_2364_[42];
  assign _zz_2408_ = _zz_2364_[43];
  assign _zz_2409_ = _zz_2364_[44];
  assign _zz_2410_ = _zz_2364_[45];
  assign _zz_2411_ = _zz_2364_[46];
  assign _zz_2412_ = _zz_2364_[47];
  assign _zz_2413_ = _zz_2364_[48];
  assign _zz_2414_ = _zz_2364_[49];
  assign _zz_2415_ = _zz_2364_[50];
  assign _zz_2416_ = _zz_2364_[51];
  assign _zz_2417_ = _zz_2364_[52];
  assign _zz_2418_ = _zz_2364_[53];
  assign _zz_2419_ = _zz_2364_[54];
  assign _zz_2420_ = _zz_2364_[55];
  assign _zz_2421_ = _zz_2364_[56];
  assign _zz_2422_ = _zz_2364_[57];
  assign _zz_2423_ = _zz_2364_[58];
  assign _zz_2424_ = _zz_2364_[59];
  assign _zz_2425_ = _zz_2364_[60];
  assign _zz_2426_ = _zz_2364_[61];
  assign _zz_2427_ = _zz_2364_[62];
  assign _zz_2428_ = _zz_2364_[63];
  assign _zz_2429_ = (((32'h00000d00 <= load_data_area_current_addr) && (load_data_area_current_addr < 32'h00000d40)) ? _zz_9__regNext : {_zz_4502_,_zz_4503_});
  assign _zz_2430_ = _zz_2429_[15 : 0];
  assign _zz_2431_ = _zz_2429_[31 : 16];
  assign _zz_2432_ = _zz_4601_[5:0];
  assign _zz_2433_ = ({63'd0,(1'b1)} <<< _zz_2432_);
  assign _zz_2434_ = _zz_2433_[0];
  assign _zz_2435_ = _zz_2433_[1];
  assign _zz_2436_ = _zz_2433_[2];
  assign _zz_2437_ = _zz_2433_[3];
  assign _zz_2438_ = _zz_2433_[4];
  assign _zz_2439_ = _zz_2433_[5];
  assign _zz_2440_ = _zz_2433_[6];
  assign _zz_2441_ = _zz_2433_[7];
  assign _zz_2442_ = _zz_2433_[8];
  assign _zz_2443_ = _zz_2433_[9];
  assign _zz_2444_ = _zz_2433_[10];
  assign _zz_2445_ = _zz_2433_[11];
  assign _zz_2446_ = _zz_2433_[12];
  assign _zz_2447_ = _zz_2433_[13];
  assign _zz_2448_ = _zz_2433_[14];
  assign _zz_2449_ = _zz_2433_[15];
  assign _zz_2450_ = _zz_2433_[16];
  assign _zz_2451_ = _zz_2433_[17];
  assign _zz_2452_ = _zz_2433_[18];
  assign _zz_2453_ = _zz_2433_[19];
  assign _zz_2454_ = _zz_2433_[20];
  assign _zz_2455_ = _zz_2433_[21];
  assign _zz_2456_ = _zz_2433_[22];
  assign _zz_2457_ = _zz_2433_[23];
  assign _zz_2458_ = _zz_2433_[24];
  assign _zz_2459_ = _zz_2433_[25];
  assign _zz_2460_ = _zz_2433_[26];
  assign _zz_2461_ = _zz_2433_[27];
  assign _zz_2462_ = _zz_2433_[28];
  assign _zz_2463_ = _zz_2433_[29];
  assign _zz_2464_ = _zz_2433_[30];
  assign _zz_2465_ = _zz_2433_[31];
  assign _zz_2466_ = _zz_2433_[32];
  assign _zz_2467_ = _zz_2433_[33];
  assign _zz_2468_ = _zz_2433_[34];
  assign _zz_2469_ = _zz_2433_[35];
  assign _zz_2470_ = _zz_2433_[36];
  assign _zz_2471_ = _zz_2433_[37];
  assign _zz_2472_ = _zz_2433_[38];
  assign _zz_2473_ = _zz_2433_[39];
  assign _zz_2474_ = _zz_2433_[40];
  assign _zz_2475_ = _zz_2433_[41];
  assign _zz_2476_ = _zz_2433_[42];
  assign _zz_2477_ = _zz_2433_[43];
  assign _zz_2478_ = _zz_2433_[44];
  assign _zz_2479_ = _zz_2433_[45];
  assign _zz_2480_ = _zz_2433_[46];
  assign _zz_2481_ = _zz_2433_[47];
  assign _zz_2482_ = _zz_2433_[48];
  assign _zz_2483_ = _zz_2433_[49];
  assign _zz_2484_ = _zz_2433_[50];
  assign _zz_2485_ = _zz_2433_[51];
  assign _zz_2486_ = _zz_2433_[52];
  assign _zz_2487_ = _zz_2433_[53];
  assign _zz_2488_ = _zz_2433_[54];
  assign _zz_2489_ = _zz_2433_[55];
  assign _zz_2490_ = _zz_2433_[56];
  assign _zz_2491_ = _zz_2433_[57];
  assign _zz_2492_ = _zz_2433_[58];
  assign _zz_2493_ = _zz_2433_[59];
  assign _zz_2494_ = _zz_2433_[60];
  assign _zz_2495_ = _zz_2433_[61];
  assign _zz_2496_ = _zz_2433_[62];
  assign _zz_2497_ = _zz_2433_[63];
  assign _zz_2498_ = (((32'h00000240 <= load_data_area_current_addr) && (load_data_area_current_addr < 32'h00000280)) ? _zz_9__regNext : {_zz_4504_,_zz_4505_});
  assign _zz_2499_ = _zz_2498_[15 : 0];
  assign _zz_2500_ = _zz_2498_[31 : 16];
  assign _zz_2501_ = _zz_4602_[5:0];
  assign _zz_2502_ = ({63'd0,(1'b1)} <<< _zz_2501_);
  assign _zz_2503_ = _zz_2502_[0];
  assign _zz_2504_ = _zz_2502_[1];
  assign _zz_2505_ = _zz_2502_[2];
  assign _zz_2506_ = _zz_2502_[3];
  assign _zz_2507_ = _zz_2502_[4];
  assign _zz_2508_ = _zz_2502_[5];
  assign _zz_2509_ = _zz_2502_[6];
  assign _zz_2510_ = _zz_2502_[7];
  assign _zz_2511_ = _zz_2502_[8];
  assign _zz_2512_ = _zz_2502_[9];
  assign _zz_2513_ = _zz_2502_[10];
  assign _zz_2514_ = _zz_2502_[11];
  assign _zz_2515_ = _zz_2502_[12];
  assign _zz_2516_ = _zz_2502_[13];
  assign _zz_2517_ = _zz_2502_[14];
  assign _zz_2518_ = _zz_2502_[15];
  assign _zz_2519_ = _zz_2502_[16];
  assign _zz_2520_ = _zz_2502_[17];
  assign _zz_2521_ = _zz_2502_[18];
  assign _zz_2522_ = _zz_2502_[19];
  assign _zz_2523_ = _zz_2502_[20];
  assign _zz_2524_ = _zz_2502_[21];
  assign _zz_2525_ = _zz_2502_[22];
  assign _zz_2526_ = _zz_2502_[23];
  assign _zz_2527_ = _zz_2502_[24];
  assign _zz_2528_ = _zz_2502_[25];
  assign _zz_2529_ = _zz_2502_[26];
  assign _zz_2530_ = _zz_2502_[27];
  assign _zz_2531_ = _zz_2502_[28];
  assign _zz_2532_ = _zz_2502_[29];
  assign _zz_2533_ = _zz_2502_[30];
  assign _zz_2534_ = _zz_2502_[31];
  assign _zz_2535_ = _zz_2502_[32];
  assign _zz_2536_ = _zz_2502_[33];
  assign _zz_2537_ = _zz_2502_[34];
  assign _zz_2538_ = _zz_2502_[35];
  assign _zz_2539_ = _zz_2502_[36];
  assign _zz_2540_ = _zz_2502_[37];
  assign _zz_2541_ = _zz_2502_[38];
  assign _zz_2542_ = _zz_2502_[39];
  assign _zz_2543_ = _zz_2502_[40];
  assign _zz_2544_ = _zz_2502_[41];
  assign _zz_2545_ = _zz_2502_[42];
  assign _zz_2546_ = _zz_2502_[43];
  assign _zz_2547_ = _zz_2502_[44];
  assign _zz_2548_ = _zz_2502_[45];
  assign _zz_2549_ = _zz_2502_[46];
  assign _zz_2550_ = _zz_2502_[47];
  assign _zz_2551_ = _zz_2502_[48];
  assign _zz_2552_ = _zz_2502_[49];
  assign _zz_2553_ = _zz_2502_[50];
  assign _zz_2554_ = _zz_2502_[51];
  assign _zz_2555_ = _zz_2502_[52];
  assign _zz_2556_ = _zz_2502_[53];
  assign _zz_2557_ = _zz_2502_[54];
  assign _zz_2558_ = _zz_2502_[55];
  assign _zz_2559_ = _zz_2502_[56];
  assign _zz_2560_ = _zz_2502_[57];
  assign _zz_2561_ = _zz_2502_[58];
  assign _zz_2562_ = _zz_2502_[59];
  assign _zz_2563_ = _zz_2502_[60];
  assign _zz_2564_ = _zz_2502_[61];
  assign _zz_2565_ = _zz_2502_[62];
  assign _zz_2566_ = _zz_2502_[63];
  assign _zz_2567_ = (((32'h00000a00 <= load_data_area_current_addr) && (load_data_area_current_addr < 32'h00000a40)) ? _zz_9__regNext : {_zz_4506_,_zz_4507_});
  assign _zz_2568_ = _zz_2567_[15 : 0];
  assign _zz_2569_ = _zz_2567_[31 : 16];
  assign _zz_2570_ = _zz_4603_[5:0];
  assign _zz_2571_ = ({63'd0,(1'b1)} <<< _zz_2570_);
  assign _zz_2572_ = _zz_2571_[0];
  assign _zz_2573_ = _zz_2571_[1];
  assign _zz_2574_ = _zz_2571_[2];
  assign _zz_2575_ = _zz_2571_[3];
  assign _zz_2576_ = _zz_2571_[4];
  assign _zz_2577_ = _zz_2571_[5];
  assign _zz_2578_ = _zz_2571_[6];
  assign _zz_2579_ = _zz_2571_[7];
  assign _zz_2580_ = _zz_2571_[8];
  assign _zz_2581_ = _zz_2571_[9];
  assign _zz_2582_ = _zz_2571_[10];
  assign _zz_2583_ = _zz_2571_[11];
  assign _zz_2584_ = _zz_2571_[12];
  assign _zz_2585_ = _zz_2571_[13];
  assign _zz_2586_ = _zz_2571_[14];
  assign _zz_2587_ = _zz_2571_[15];
  assign _zz_2588_ = _zz_2571_[16];
  assign _zz_2589_ = _zz_2571_[17];
  assign _zz_2590_ = _zz_2571_[18];
  assign _zz_2591_ = _zz_2571_[19];
  assign _zz_2592_ = _zz_2571_[20];
  assign _zz_2593_ = _zz_2571_[21];
  assign _zz_2594_ = _zz_2571_[22];
  assign _zz_2595_ = _zz_2571_[23];
  assign _zz_2596_ = _zz_2571_[24];
  assign _zz_2597_ = _zz_2571_[25];
  assign _zz_2598_ = _zz_2571_[26];
  assign _zz_2599_ = _zz_2571_[27];
  assign _zz_2600_ = _zz_2571_[28];
  assign _zz_2601_ = _zz_2571_[29];
  assign _zz_2602_ = _zz_2571_[30];
  assign _zz_2603_ = _zz_2571_[31];
  assign _zz_2604_ = _zz_2571_[32];
  assign _zz_2605_ = _zz_2571_[33];
  assign _zz_2606_ = _zz_2571_[34];
  assign _zz_2607_ = _zz_2571_[35];
  assign _zz_2608_ = _zz_2571_[36];
  assign _zz_2609_ = _zz_2571_[37];
  assign _zz_2610_ = _zz_2571_[38];
  assign _zz_2611_ = _zz_2571_[39];
  assign _zz_2612_ = _zz_2571_[40];
  assign _zz_2613_ = _zz_2571_[41];
  assign _zz_2614_ = _zz_2571_[42];
  assign _zz_2615_ = _zz_2571_[43];
  assign _zz_2616_ = _zz_2571_[44];
  assign _zz_2617_ = _zz_2571_[45];
  assign _zz_2618_ = _zz_2571_[46];
  assign _zz_2619_ = _zz_2571_[47];
  assign _zz_2620_ = _zz_2571_[48];
  assign _zz_2621_ = _zz_2571_[49];
  assign _zz_2622_ = _zz_2571_[50];
  assign _zz_2623_ = _zz_2571_[51];
  assign _zz_2624_ = _zz_2571_[52];
  assign _zz_2625_ = _zz_2571_[53];
  assign _zz_2626_ = _zz_2571_[54];
  assign _zz_2627_ = _zz_2571_[55];
  assign _zz_2628_ = _zz_2571_[56];
  assign _zz_2629_ = _zz_2571_[57];
  assign _zz_2630_ = _zz_2571_[58];
  assign _zz_2631_ = _zz_2571_[59];
  assign _zz_2632_ = _zz_2571_[60];
  assign _zz_2633_ = _zz_2571_[61];
  assign _zz_2634_ = _zz_2571_[62];
  assign _zz_2635_ = _zz_2571_[63];
  assign _zz_2636_ = (((32'h00000640 <= load_data_area_current_addr) && (load_data_area_current_addr < 32'h00000680)) ? _zz_9__regNext : {_zz_4508_,_zz_4509_});
  assign _zz_2637_ = _zz_2636_[15 : 0];
  assign _zz_2638_ = _zz_2636_[31 : 16];
  assign _zz_2639_ = _zz_4604_[5:0];
  assign _zz_2640_ = ({63'd0,(1'b1)} <<< _zz_2639_);
  assign _zz_2641_ = _zz_2640_[0];
  assign _zz_2642_ = _zz_2640_[1];
  assign _zz_2643_ = _zz_2640_[2];
  assign _zz_2644_ = _zz_2640_[3];
  assign _zz_2645_ = _zz_2640_[4];
  assign _zz_2646_ = _zz_2640_[5];
  assign _zz_2647_ = _zz_2640_[6];
  assign _zz_2648_ = _zz_2640_[7];
  assign _zz_2649_ = _zz_2640_[8];
  assign _zz_2650_ = _zz_2640_[9];
  assign _zz_2651_ = _zz_2640_[10];
  assign _zz_2652_ = _zz_2640_[11];
  assign _zz_2653_ = _zz_2640_[12];
  assign _zz_2654_ = _zz_2640_[13];
  assign _zz_2655_ = _zz_2640_[14];
  assign _zz_2656_ = _zz_2640_[15];
  assign _zz_2657_ = _zz_2640_[16];
  assign _zz_2658_ = _zz_2640_[17];
  assign _zz_2659_ = _zz_2640_[18];
  assign _zz_2660_ = _zz_2640_[19];
  assign _zz_2661_ = _zz_2640_[20];
  assign _zz_2662_ = _zz_2640_[21];
  assign _zz_2663_ = _zz_2640_[22];
  assign _zz_2664_ = _zz_2640_[23];
  assign _zz_2665_ = _zz_2640_[24];
  assign _zz_2666_ = _zz_2640_[25];
  assign _zz_2667_ = _zz_2640_[26];
  assign _zz_2668_ = _zz_2640_[27];
  assign _zz_2669_ = _zz_2640_[28];
  assign _zz_2670_ = _zz_2640_[29];
  assign _zz_2671_ = _zz_2640_[30];
  assign _zz_2672_ = _zz_2640_[31];
  assign _zz_2673_ = _zz_2640_[32];
  assign _zz_2674_ = _zz_2640_[33];
  assign _zz_2675_ = _zz_2640_[34];
  assign _zz_2676_ = _zz_2640_[35];
  assign _zz_2677_ = _zz_2640_[36];
  assign _zz_2678_ = _zz_2640_[37];
  assign _zz_2679_ = _zz_2640_[38];
  assign _zz_2680_ = _zz_2640_[39];
  assign _zz_2681_ = _zz_2640_[40];
  assign _zz_2682_ = _zz_2640_[41];
  assign _zz_2683_ = _zz_2640_[42];
  assign _zz_2684_ = _zz_2640_[43];
  assign _zz_2685_ = _zz_2640_[44];
  assign _zz_2686_ = _zz_2640_[45];
  assign _zz_2687_ = _zz_2640_[46];
  assign _zz_2688_ = _zz_2640_[47];
  assign _zz_2689_ = _zz_2640_[48];
  assign _zz_2690_ = _zz_2640_[49];
  assign _zz_2691_ = _zz_2640_[50];
  assign _zz_2692_ = _zz_2640_[51];
  assign _zz_2693_ = _zz_2640_[52];
  assign _zz_2694_ = _zz_2640_[53];
  assign _zz_2695_ = _zz_2640_[54];
  assign _zz_2696_ = _zz_2640_[55];
  assign _zz_2697_ = _zz_2640_[56];
  assign _zz_2698_ = _zz_2640_[57];
  assign _zz_2699_ = _zz_2640_[58];
  assign _zz_2700_ = _zz_2640_[59];
  assign _zz_2701_ = _zz_2640_[60];
  assign _zz_2702_ = _zz_2640_[61];
  assign _zz_2703_ = _zz_2640_[62];
  assign _zz_2704_ = _zz_2640_[63];
  assign _zz_2705_ = (((32'h00000080 <= load_data_area_current_addr) && (load_data_area_current_addr < 32'h000000c0)) ? _zz_9__regNext : {_zz_4510_,_zz_4511_});
  assign _zz_2706_ = _zz_2705_[15 : 0];
  assign _zz_2707_ = _zz_2705_[31 : 16];
  assign _zz_2708_ = _zz_4605_[5:0];
  assign _zz_2709_ = ({63'd0,(1'b1)} <<< _zz_2708_);
  assign _zz_2710_ = _zz_2709_[0];
  assign _zz_2711_ = _zz_2709_[1];
  assign _zz_2712_ = _zz_2709_[2];
  assign _zz_2713_ = _zz_2709_[3];
  assign _zz_2714_ = _zz_2709_[4];
  assign _zz_2715_ = _zz_2709_[5];
  assign _zz_2716_ = _zz_2709_[6];
  assign _zz_2717_ = _zz_2709_[7];
  assign _zz_2718_ = _zz_2709_[8];
  assign _zz_2719_ = _zz_2709_[9];
  assign _zz_2720_ = _zz_2709_[10];
  assign _zz_2721_ = _zz_2709_[11];
  assign _zz_2722_ = _zz_2709_[12];
  assign _zz_2723_ = _zz_2709_[13];
  assign _zz_2724_ = _zz_2709_[14];
  assign _zz_2725_ = _zz_2709_[15];
  assign _zz_2726_ = _zz_2709_[16];
  assign _zz_2727_ = _zz_2709_[17];
  assign _zz_2728_ = _zz_2709_[18];
  assign _zz_2729_ = _zz_2709_[19];
  assign _zz_2730_ = _zz_2709_[20];
  assign _zz_2731_ = _zz_2709_[21];
  assign _zz_2732_ = _zz_2709_[22];
  assign _zz_2733_ = _zz_2709_[23];
  assign _zz_2734_ = _zz_2709_[24];
  assign _zz_2735_ = _zz_2709_[25];
  assign _zz_2736_ = _zz_2709_[26];
  assign _zz_2737_ = _zz_2709_[27];
  assign _zz_2738_ = _zz_2709_[28];
  assign _zz_2739_ = _zz_2709_[29];
  assign _zz_2740_ = _zz_2709_[30];
  assign _zz_2741_ = _zz_2709_[31];
  assign _zz_2742_ = _zz_2709_[32];
  assign _zz_2743_ = _zz_2709_[33];
  assign _zz_2744_ = _zz_2709_[34];
  assign _zz_2745_ = _zz_2709_[35];
  assign _zz_2746_ = _zz_2709_[36];
  assign _zz_2747_ = _zz_2709_[37];
  assign _zz_2748_ = _zz_2709_[38];
  assign _zz_2749_ = _zz_2709_[39];
  assign _zz_2750_ = _zz_2709_[40];
  assign _zz_2751_ = _zz_2709_[41];
  assign _zz_2752_ = _zz_2709_[42];
  assign _zz_2753_ = _zz_2709_[43];
  assign _zz_2754_ = _zz_2709_[44];
  assign _zz_2755_ = _zz_2709_[45];
  assign _zz_2756_ = _zz_2709_[46];
  assign _zz_2757_ = _zz_2709_[47];
  assign _zz_2758_ = _zz_2709_[48];
  assign _zz_2759_ = _zz_2709_[49];
  assign _zz_2760_ = _zz_2709_[50];
  assign _zz_2761_ = _zz_2709_[51];
  assign _zz_2762_ = _zz_2709_[52];
  assign _zz_2763_ = _zz_2709_[53];
  assign _zz_2764_ = _zz_2709_[54];
  assign _zz_2765_ = _zz_2709_[55];
  assign _zz_2766_ = _zz_2709_[56];
  assign _zz_2767_ = _zz_2709_[57];
  assign _zz_2768_ = _zz_2709_[58];
  assign _zz_2769_ = _zz_2709_[59];
  assign _zz_2770_ = _zz_2709_[60];
  assign _zz_2771_ = _zz_2709_[61];
  assign _zz_2772_ = _zz_2709_[62];
  assign _zz_2773_ = _zz_2709_[63];
  assign _zz_2774_ = (((32'h00000840 <= load_data_area_current_addr) && (load_data_area_current_addr < 32'h00000880)) ? _zz_9__regNext : {_zz_4512_,_zz_4513_});
  assign _zz_2775_ = _zz_2774_[15 : 0];
  assign _zz_2776_ = _zz_2774_[31 : 16];
  assign _zz_2777_ = _zz_4606_[5:0];
  assign _zz_2778_ = ({63'd0,(1'b1)} <<< _zz_2777_);
  assign _zz_2779_ = _zz_2778_[0];
  assign _zz_2780_ = _zz_2778_[1];
  assign _zz_2781_ = _zz_2778_[2];
  assign _zz_2782_ = _zz_2778_[3];
  assign _zz_2783_ = _zz_2778_[4];
  assign _zz_2784_ = _zz_2778_[5];
  assign _zz_2785_ = _zz_2778_[6];
  assign _zz_2786_ = _zz_2778_[7];
  assign _zz_2787_ = _zz_2778_[8];
  assign _zz_2788_ = _zz_2778_[9];
  assign _zz_2789_ = _zz_2778_[10];
  assign _zz_2790_ = _zz_2778_[11];
  assign _zz_2791_ = _zz_2778_[12];
  assign _zz_2792_ = _zz_2778_[13];
  assign _zz_2793_ = _zz_2778_[14];
  assign _zz_2794_ = _zz_2778_[15];
  assign _zz_2795_ = _zz_2778_[16];
  assign _zz_2796_ = _zz_2778_[17];
  assign _zz_2797_ = _zz_2778_[18];
  assign _zz_2798_ = _zz_2778_[19];
  assign _zz_2799_ = _zz_2778_[20];
  assign _zz_2800_ = _zz_2778_[21];
  assign _zz_2801_ = _zz_2778_[22];
  assign _zz_2802_ = _zz_2778_[23];
  assign _zz_2803_ = _zz_2778_[24];
  assign _zz_2804_ = _zz_2778_[25];
  assign _zz_2805_ = _zz_2778_[26];
  assign _zz_2806_ = _zz_2778_[27];
  assign _zz_2807_ = _zz_2778_[28];
  assign _zz_2808_ = _zz_2778_[29];
  assign _zz_2809_ = _zz_2778_[30];
  assign _zz_2810_ = _zz_2778_[31];
  assign _zz_2811_ = _zz_2778_[32];
  assign _zz_2812_ = _zz_2778_[33];
  assign _zz_2813_ = _zz_2778_[34];
  assign _zz_2814_ = _zz_2778_[35];
  assign _zz_2815_ = _zz_2778_[36];
  assign _zz_2816_ = _zz_2778_[37];
  assign _zz_2817_ = _zz_2778_[38];
  assign _zz_2818_ = _zz_2778_[39];
  assign _zz_2819_ = _zz_2778_[40];
  assign _zz_2820_ = _zz_2778_[41];
  assign _zz_2821_ = _zz_2778_[42];
  assign _zz_2822_ = _zz_2778_[43];
  assign _zz_2823_ = _zz_2778_[44];
  assign _zz_2824_ = _zz_2778_[45];
  assign _zz_2825_ = _zz_2778_[46];
  assign _zz_2826_ = _zz_2778_[47];
  assign _zz_2827_ = _zz_2778_[48];
  assign _zz_2828_ = _zz_2778_[49];
  assign _zz_2829_ = _zz_2778_[50];
  assign _zz_2830_ = _zz_2778_[51];
  assign _zz_2831_ = _zz_2778_[52];
  assign _zz_2832_ = _zz_2778_[53];
  assign _zz_2833_ = _zz_2778_[54];
  assign _zz_2834_ = _zz_2778_[55];
  assign _zz_2835_ = _zz_2778_[56];
  assign _zz_2836_ = _zz_2778_[57];
  assign _zz_2837_ = _zz_2778_[58];
  assign _zz_2838_ = _zz_2778_[59];
  assign _zz_2839_ = _zz_2778_[60];
  assign _zz_2840_ = _zz_2778_[61];
  assign _zz_2841_ = _zz_2778_[62];
  assign _zz_2842_ = _zz_2778_[63];
  assign _zz_2843_ = (((32'h00000140 <= load_data_area_current_addr) && (load_data_area_current_addr < 32'h00000180)) ? _zz_9__regNext : {_zz_4514_,_zz_4515_});
  assign _zz_2844_ = _zz_2843_[15 : 0];
  assign _zz_2845_ = _zz_2843_[31 : 16];
  assign _zz_2846_ = _zz_4607_[5:0];
  assign _zz_2847_ = ({63'd0,(1'b1)} <<< _zz_2846_);
  assign _zz_2848_ = _zz_2847_[0];
  assign _zz_2849_ = _zz_2847_[1];
  assign _zz_2850_ = _zz_2847_[2];
  assign _zz_2851_ = _zz_2847_[3];
  assign _zz_2852_ = _zz_2847_[4];
  assign _zz_2853_ = _zz_2847_[5];
  assign _zz_2854_ = _zz_2847_[6];
  assign _zz_2855_ = _zz_2847_[7];
  assign _zz_2856_ = _zz_2847_[8];
  assign _zz_2857_ = _zz_2847_[9];
  assign _zz_2858_ = _zz_2847_[10];
  assign _zz_2859_ = _zz_2847_[11];
  assign _zz_2860_ = _zz_2847_[12];
  assign _zz_2861_ = _zz_2847_[13];
  assign _zz_2862_ = _zz_2847_[14];
  assign _zz_2863_ = _zz_2847_[15];
  assign _zz_2864_ = _zz_2847_[16];
  assign _zz_2865_ = _zz_2847_[17];
  assign _zz_2866_ = _zz_2847_[18];
  assign _zz_2867_ = _zz_2847_[19];
  assign _zz_2868_ = _zz_2847_[20];
  assign _zz_2869_ = _zz_2847_[21];
  assign _zz_2870_ = _zz_2847_[22];
  assign _zz_2871_ = _zz_2847_[23];
  assign _zz_2872_ = _zz_2847_[24];
  assign _zz_2873_ = _zz_2847_[25];
  assign _zz_2874_ = _zz_2847_[26];
  assign _zz_2875_ = _zz_2847_[27];
  assign _zz_2876_ = _zz_2847_[28];
  assign _zz_2877_ = _zz_2847_[29];
  assign _zz_2878_ = _zz_2847_[30];
  assign _zz_2879_ = _zz_2847_[31];
  assign _zz_2880_ = _zz_2847_[32];
  assign _zz_2881_ = _zz_2847_[33];
  assign _zz_2882_ = _zz_2847_[34];
  assign _zz_2883_ = _zz_2847_[35];
  assign _zz_2884_ = _zz_2847_[36];
  assign _zz_2885_ = _zz_2847_[37];
  assign _zz_2886_ = _zz_2847_[38];
  assign _zz_2887_ = _zz_2847_[39];
  assign _zz_2888_ = _zz_2847_[40];
  assign _zz_2889_ = _zz_2847_[41];
  assign _zz_2890_ = _zz_2847_[42];
  assign _zz_2891_ = _zz_2847_[43];
  assign _zz_2892_ = _zz_2847_[44];
  assign _zz_2893_ = _zz_2847_[45];
  assign _zz_2894_ = _zz_2847_[46];
  assign _zz_2895_ = _zz_2847_[47];
  assign _zz_2896_ = _zz_2847_[48];
  assign _zz_2897_ = _zz_2847_[49];
  assign _zz_2898_ = _zz_2847_[50];
  assign _zz_2899_ = _zz_2847_[51];
  assign _zz_2900_ = _zz_2847_[52];
  assign _zz_2901_ = _zz_2847_[53];
  assign _zz_2902_ = _zz_2847_[54];
  assign _zz_2903_ = _zz_2847_[55];
  assign _zz_2904_ = _zz_2847_[56];
  assign _zz_2905_ = _zz_2847_[57];
  assign _zz_2906_ = _zz_2847_[58];
  assign _zz_2907_ = _zz_2847_[59];
  assign _zz_2908_ = _zz_2847_[60];
  assign _zz_2909_ = _zz_2847_[61];
  assign _zz_2910_ = _zz_2847_[62];
  assign _zz_2911_ = _zz_2847_[63];
  assign _zz_2912_ = (((32'h000000c0 <= load_data_area_current_addr) && (load_data_area_current_addr < 32'h00000100)) ? _zz_9__regNext : {_zz_4516_,_zz_4517_});
  assign _zz_2913_ = _zz_2912_[15 : 0];
  assign _zz_2914_ = _zz_2912_[31 : 16];
  assign _zz_2915_ = _zz_4608_[5:0];
  assign _zz_2916_ = ({63'd0,(1'b1)} <<< _zz_2915_);
  assign _zz_2917_ = _zz_2916_[0];
  assign _zz_2918_ = _zz_2916_[1];
  assign _zz_2919_ = _zz_2916_[2];
  assign _zz_2920_ = _zz_2916_[3];
  assign _zz_2921_ = _zz_2916_[4];
  assign _zz_2922_ = _zz_2916_[5];
  assign _zz_2923_ = _zz_2916_[6];
  assign _zz_2924_ = _zz_2916_[7];
  assign _zz_2925_ = _zz_2916_[8];
  assign _zz_2926_ = _zz_2916_[9];
  assign _zz_2927_ = _zz_2916_[10];
  assign _zz_2928_ = _zz_2916_[11];
  assign _zz_2929_ = _zz_2916_[12];
  assign _zz_2930_ = _zz_2916_[13];
  assign _zz_2931_ = _zz_2916_[14];
  assign _zz_2932_ = _zz_2916_[15];
  assign _zz_2933_ = _zz_2916_[16];
  assign _zz_2934_ = _zz_2916_[17];
  assign _zz_2935_ = _zz_2916_[18];
  assign _zz_2936_ = _zz_2916_[19];
  assign _zz_2937_ = _zz_2916_[20];
  assign _zz_2938_ = _zz_2916_[21];
  assign _zz_2939_ = _zz_2916_[22];
  assign _zz_2940_ = _zz_2916_[23];
  assign _zz_2941_ = _zz_2916_[24];
  assign _zz_2942_ = _zz_2916_[25];
  assign _zz_2943_ = _zz_2916_[26];
  assign _zz_2944_ = _zz_2916_[27];
  assign _zz_2945_ = _zz_2916_[28];
  assign _zz_2946_ = _zz_2916_[29];
  assign _zz_2947_ = _zz_2916_[30];
  assign _zz_2948_ = _zz_2916_[31];
  assign _zz_2949_ = _zz_2916_[32];
  assign _zz_2950_ = _zz_2916_[33];
  assign _zz_2951_ = _zz_2916_[34];
  assign _zz_2952_ = _zz_2916_[35];
  assign _zz_2953_ = _zz_2916_[36];
  assign _zz_2954_ = _zz_2916_[37];
  assign _zz_2955_ = _zz_2916_[38];
  assign _zz_2956_ = _zz_2916_[39];
  assign _zz_2957_ = _zz_2916_[40];
  assign _zz_2958_ = _zz_2916_[41];
  assign _zz_2959_ = _zz_2916_[42];
  assign _zz_2960_ = _zz_2916_[43];
  assign _zz_2961_ = _zz_2916_[44];
  assign _zz_2962_ = _zz_2916_[45];
  assign _zz_2963_ = _zz_2916_[46];
  assign _zz_2964_ = _zz_2916_[47];
  assign _zz_2965_ = _zz_2916_[48];
  assign _zz_2966_ = _zz_2916_[49];
  assign _zz_2967_ = _zz_2916_[50];
  assign _zz_2968_ = _zz_2916_[51];
  assign _zz_2969_ = _zz_2916_[52];
  assign _zz_2970_ = _zz_2916_[53];
  assign _zz_2971_ = _zz_2916_[54];
  assign _zz_2972_ = _zz_2916_[55];
  assign _zz_2973_ = _zz_2916_[56];
  assign _zz_2974_ = _zz_2916_[57];
  assign _zz_2975_ = _zz_2916_[58];
  assign _zz_2976_ = _zz_2916_[59];
  assign _zz_2977_ = _zz_2916_[60];
  assign _zz_2978_ = _zz_2916_[61];
  assign _zz_2979_ = _zz_2916_[62];
  assign _zz_2980_ = _zz_2916_[63];
  assign _zz_2981_ = (((32'h00000340 <= load_data_area_current_addr) && (load_data_area_current_addr < 32'h00000380)) ? _zz_9__regNext : {_zz_4518_,_zz_4519_});
  assign _zz_2982_ = _zz_2981_[15 : 0];
  assign _zz_2983_ = _zz_2981_[31 : 16];
  assign _zz_2984_ = _zz_4609_[5:0];
  assign _zz_2985_ = ({63'd0,(1'b1)} <<< _zz_2984_);
  assign _zz_2986_ = _zz_2985_[0];
  assign _zz_2987_ = _zz_2985_[1];
  assign _zz_2988_ = _zz_2985_[2];
  assign _zz_2989_ = _zz_2985_[3];
  assign _zz_2990_ = _zz_2985_[4];
  assign _zz_2991_ = _zz_2985_[5];
  assign _zz_2992_ = _zz_2985_[6];
  assign _zz_2993_ = _zz_2985_[7];
  assign _zz_2994_ = _zz_2985_[8];
  assign _zz_2995_ = _zz_2985_[9];
  assign _zz_2996_ = _zz_2985_[10];
  assign _zz_2997_ = _zz_2985_[11];
  assign _zz_2998_ = _zz_2985_[12];
  assign _zz_2999_ = _zz_2985_[13];
  assign _zz_3000_ = _zz_2985_[14];
  assign _zz_3001_ = _zz_2985_[15];
  assign _zz_3002_ = _zz_2985_[16];
  assign _zz_3003_ = _zz_2985_[17];
  assign _zz_3004_ = _zz_2985_[18];
  assign _zz_3005_ = _zz_2985_[19];
  assign _zz_3006_ = _zz_2985_[20];
  assign _zz_3007_ = _zz_2985_[21];
  assign _zz_3008_ = _zz_2985_[22];
  assign _zz_3009_ = _zz_2985_[23];
  assign _zz_3010_ = _zz_2985_[24];
  assign _zz_3011_ = _zz_2985_[25];
  assign _zz_3012_ = _zz_2985_[26];
  assign _zz_3013_ = _zz_2985_[27];
  assign _zz_3014_ = _zz_2985_[28];
  assign _zz_3015_ = _zz_2985_[29];
  assign _zz_3016_ = _zz_2985_[30];
  assign _zz_3017_ = _zz_2985_[31];
  assign _zz_3018_ = _zz_2985_[32];
  assign _zz_3019_ = _zz_2985_[33];
  assign _zz_3020_ = _zz_2985_[34];
  assign _zz_3021_ = _zz_2985_[35];
  assign _zz_3022_ = _zz_2985_[36];
  assign _zz_3023_ = _zz_2985_[37];
  assign _zz_3024_ = _zz_2985_[38];
  assign _zz_3025_ = _zz_2985_[39];
  assign _zz_3026_ = _zz_2985_[40];
  assign _zz_3027_ = _zz_2985_[41];
  assign _zz_3028_ = _zz_2985_[42];
  assign _zz_3029_ = _zz_2985_[43];
  assign _zz_3030_ = _zz_2985_[44];
  assign _zz_3031_ = _zz_2985_[45];
  assign _zz_3032_ = _zz_2985_[46];
  assign _zz_3033_ = _zz_2985_[47];
  assign _zz_3034_ = _zz_2985_[48];
  assign _zz_3035_ = _zz_2985_[49];
  assign _zz_3036_ = _zz_2985_[50];
  assign _zz_3037_ = _zz_2985_[51];
  assign _zz_3038_ = _zz_2985_[52];
  assign _zz_3039_ = _zz_2985_[53];
  assign _zz_3040_ = _zz_2985_[54];
  assign _zz_3041_ = _zz_2985_[55];
  assign _zz_3042_ = _zz_2985_[56];
  assign _zz_3043_ = _zz_2985_[57];
  assign _zz_3044_ = _zz_2985_[58];
  assign _zz_3045_ = _zz_2985_[59];
  assign _zz_3046_ = _zz_2985_[60];
  assign _zz_3047_ = _zz_2985_[61];
  assign _zz_3048_ = _zz_2985_[62];
  assign _zz_3049_ = _zz_2985_[63];
  assign _zz_3050_ = (((32'h00000dc0 <= load_data_area_current_addr) && (load_data_area_current_addr < 32'h00000e00)) ? _zz_9__regNext : {_zz_4520_,_zz_4521_});
  assign _zz_3051_ = _zz_3050_[15 : 0];
  assign _zz_3052_ = _zz_3050_[31 : 16];
  assign _zz_3053_ = _zz_4610_[5:0];
  assign _zz_3054_ = ({63'd0,(1'b1)} <<< _zz_3053_);
  assign _zz_3055_ = _zz_3054_[0];
  assign _zz_3056_ = _zz_3054_[1];
  assign _zz_3057_ = _zz_3054_[2];
  assign _zz_3058_ = _zz_3054_[3];
  assign _zz_3059_ = _zz_3054_[4];
  assign _zz_3060_ = _zz_3054_[5];
  assign _zz_3061_ = _zz_3054_[6];
  assign _zz_3062_ = _zz_3054_[7];
  assign _zz_3063_ = _zz_3054_[8];
  assign _zz_3064_ = _zz_3054_[9];
  assign _zz_3065_ = _zz_3054_[10];
  assign _zz_3066_ = _zz_3054_[11];
  assign _zz_3067_ = _zz_3054_[12];
  assign _zz_3068_ = _zz_3054_[13];
  assign _zz_3069_ = _zz_3054_[14];
  assign _zz_3070_ = _zz_3054_[15];
  assign _zz_3071_ = _zz_3054_[16];
  assign _zz_3072_ = _zz_3054_[17];
  assign _zz_3073_ = _zz_3054_[18];
  assign _zz_3074_ = _zz_3054_[19];
  assign _zz_3075_ = _zz_3054_[20];
  assign _zz_3076_ = _zz_3054_[21];
  assign _zz_3077_ = _zz_3054_[22];
  assign _zz_3078_ = _zz_3054_[23];
  assign _zz_3079_ = _zz_3054_[24];
  assign _zz_3080_ = _zz_3054_[25];
  assign _zz_3081_ = _zz_3054_[26];
  assign _zz_3082_ = _zz_3054_[27];
  assign _zz_3083_ = _zz_3054_[28];
  assign _zz_3084_ = _zz_3054_[29];
  assign _zz_3085_ = _zz_3054_[30];
  assign _zz_3086_ = _zz_3054_[31];
  assign _zz_3087_ = _zz_3054_[32];
  assign _zz_3088_ = _zz_3054_[33];
  assign _zz_3089_ = _zz_3054_[34];
  assign _zz_3090_ = _zz_3054_[35];
  assign _zz_3091_ = _zz_3054_[36];
  assign _zz_3092_ = _zz_3054_[37];
  assign _zz_3093_ = _zz_3054_[38];
  assign _zz_3094_ = _zz_3054_[39];
  assign _zz_3095_ = _zz_3054_[40];
  assign _zz_3096_ = _zz_3054_[41];
  assign _zz_3097_ = _zz_3054_[42];
  assign _zz_3098_ = _zz_3054_[43];
  assign _zz_3099_ = _zz_3054_[44];
  assign _zz_3100_ = _zz_3054_[45];
  assign _zz_3101_ = _zz_3054_[46];
  assign _zz_3102_ = _zz_3054_[47];
  assign _zz_3103_ = _zz_3054_[48];
  assign _zz_3104_ = _zz_3054_[49];
  assign _zz_3105_ = _zz_3054_[50];
  assign _zz_3106_ = _zz_3054_[51];
  assign _zz_3107_ = _zz_3054_[52];
  assign _zz_3108_ = _zz_3054_[53];
  assign _zz_3109_ = _zz_3054_[54];
  assign _zz_3110_ = _zz_3054_[55];
  assign _zz_3111_ = _zz_3054_[56];
  assign _zz_3112_ = _zz_3054_[57];
  assign _zz_3113_ = _zz_3054_[58];
  assign _zz_3114_ = _zz_3054_[59];
  assign _zz_3115_ = _zz_3054_[60];
  assign _zz_3116_ = _zz_3054_[61];
  assign _zz_3117_ = _zz_3054_[62];
  assign _zz_3118_ = _zz_3054_[63];
  assign _zz_3119_ = (((32'h00000d40 <= load_data_area_current_addr) && (load_data_area_current_addr < 32'h00000d80)) ? _zz_9__regNext : {_zz_4522_,_zz_4523_});
  assign _zz_3120_ = _zz_3119_[15 : 0];
  assign _zz_3121_ = _zz_3119_[31 : 16];
  assign _zz_3122_ = _zz_4611_[5:0];
  assign _zz_3123_ = ({63'd0,(1'b1)} <<< _zz_3122_);
  assign _zz_3124_ = _zz_3123_[0];
  assign _zz_3125_ = _zz_3123_[1];
  assign _zz_3126_ = _zz_3123_[2];
  assign _zz_3127_ = _zz_3123_[3];
  assign _zz_3128_ = _zz_3123_[4];
  assign _zz_3129_ = _zz_3123_[5];
  assign _zz_3130_ = _zz_3123_[6];
  assign _zz_3131_ = _zz_3123_[7];
  assign _zz_3132_ = _zz_3123_[8];
  assign _zz_3133_ = _zz_3123_[9];
  assign _zz_3134_ = _zz_3123_[10];
  assign _zz_3135_ = _zz_3123_[11];
  assign _zz_3136_ = _zz_3123_[12];
  assign _zz_3137_ = _zz_3123_[13];
  assign _zz_3138_ = _zz_3123_[14];
  assign _zz_3139_ = _zz_3123_[15];
  assign _zz_3140_ = _zz_3123_[16];
  assign _zz_3141_ = _zz_3123_[17];
  assign _zz_3142_ = _zz_3123_[18];
  assign _zz_3143_ = _zz_3123_[19];
  assign _zz_3144_ = _zz_3123_[20];
  assign _zz_3145_ = _zz_3123_[21];
  assign _zz_3146_ = _zz_3123_[22];
  assign _zz_3147_ = _zz_3123_[23];
  assign _zz_3148_ = _zz_3123_[24];
  assign _zz_3149_ = _zz_3123_[25];
  assign _zz_3150_ = _zz_3123_[26];
  assign _zz_3151_ = _zz_3123_[27];
  assign _zz_3152_ = _zz_3123_[28];
  assign _zz_3153_ = _zz_3123_[29];
  assign _zz_3154_ = _zz_3123_[30];
  assign _zz_3155_ = _zz_3123_[31];
  assign _zz_3156_ = _zz_3123_[32];
  assign _zz_3157_ = _zz_3123_[33];
  assign _zz_3158_ = _zz_3123_[34];
  assign _zz_3159_ = _zz_3123_[35];
  assign _zz_3160_ = _zz_3123_[36];
  assign _zz_3161_ = _zz_3123_[37];
  assign _zz_3162_ = _zz_3123_[38];
  assign _zz_3163_ = _zz_3123_[39];
  assign _zz_3164_ = _zz_3123_[40];
  assign _zz_3165_ = _zz_3123_[41];
  assign _zz_3166_ = _zz_3123_[42];
  assign _zz_3167_ = _zz_3123_[43];
  assign _zz_3168_ = _zz_3123_[44];
  assign _zz_3169_ = _zz_3123_[45];
  assign _zz_3170_ = _zz_3123_[46];
  assign _zz_3171_ = _zz_3123_[47];
  assign _zz_3172_ = _zz_3123_[48];
  assign _zz_3173_ = _zz_3123_[49];
  assign _zz_3174_ = _zz_3123_[50];
  assign _zz_3175_ = _zz_3123_[51];
  assign _zz_3176_ = _zz_3123_[52];
  assign _zz_3177_ = _zz_3123_[53];
  assign _zz_3178_ = _zz_3123_[54];
  assign _zz_3179_ = _zz_3123_[55];
  assign _zz_3180_ = _zz_3123_[56];
  assign _zz_3181_ = _zz_3123_[57];
  assign _zz_3182_ = _zz_3123_[58];
  assign _zz_3183_ = _zz_3123_[59];
  assign _zz_3184_ = _zz_3123_[60];
  assign _zz_3185_ = _zz_3123_[61];
  assign _zz_3186_ = _zz_3123_[62];
  assign _zz_3187_ = _zz_3123_[63];
  assign _zz_3188_ = (((32'h00000280 <= load_data_area_current_addr) && (load_data_area_current_addr < 32'h000002c0)) ? _zz_9__regNext : {_zz_4524_,_zz_4525_});
  assign _zz_3189_ = _zz_3188_[15 : 0];
  assign _zz_3190_ = _zz_3188_[31 : 16];
  assign _zz_3191_ = _zz_4612_[5:0];
  assign _zz_3192_ = ({63'd0,(1'b1)} <<< _zz_3191_);
  assign _zz_3193_ = _zz_3192_[0];
  assign _zz_3194_ = _zz_3192_[1];
  assign _zz_3195_ = _zz_3192_[2];
  assign _zz_3196_ = _zz_3192_[3];
  assign _zz_3197_ = _zz_3192_[4];
  assign _zz_3198_ = _zz_3192_[5];
  assign _zz_3199_ = _zz_3192_[6];
  assign _zz_3200_ = _zz_3192_[7];
  assign _zz_3201_ = _zz_3192_[8];
  assign _zz_3202_ = _zz_3192_[9];
  assign _zz_3203_ = _zz_3192_[10];
  assign _zz_3204_ = _zz_3192_[11];
  assign _zz_3205_ = _zz_3192_[12];
  assign _zz_3206_ = _zz_3192_[13];
  assign _zz_3207_ = _zz_3192_[14];
  assign _zz_3208_ = _zz_3192_[15];
  assign _zz_3209_ = _zz_3192_[16];
  assign _zz_3210_ = _zz_3192_[17];
  assign _zz_3211_ = _zz_3192_[18];
  assign _zz_3212_ = _zz_3192_[19];
  assign _zz_3213_ = _zz_3192_[20];
  assign _zz_3214_ = _zz_3192_[21];
  assign _zz_3215_ = _zz_3192_[22];
  assign _zz_3216_ = _zz_3192_[23];
  assign _zz_3217_ = _zz_3192_[24];
  assign _zz_3218_ = _zz_3192_[25];
  assign _zz_3219_ = _zz_3192_[26];
  assign _zz_3220_ = _zz_3192_[27];
  assign _zz_3221_ = _zz_3192_[28];
  assign _zz_3222_ = _zz_3192_[29];
  assign _zz_3223_ = _zz_3192_[30];
  assign _zz_3224_ = _zz_3192_[31];
  assign _zz_3225_ = _zz_3192_[32];
  assign _zz_3226_ = _zz_3192_[33];
  assign _zz_3227_ = _zz_3192_[34];
  assign _zz_3228_ = _zz_3192_[35];
  assign _zz_3229_ = _zz_3192_[36];
  assign _zz_3230_ = _zz_3192_[37];
  assign _zz_3231_ = _zz_3192_[38];
  assign _zz_3232_ = _zz_3192_[39];
  assign _zz_3233_ = _zz_3192_[40];
  assign _zz_3234_ = _zz_3192_[41];
  assign _zz_3235_ = _zz_3192_[42];
  assign _zz_3236_ = _zz_3192_[43];
  assign _zz_3237_ = _zz_3192_[44];
  assign _zz_3238_ = _zz_3192_[45];
  assign _zz_3239_ = _zz_3192_[46];
  assign _zz_3240_ = _zz_3192_[47];
  assign _zz_3241_ = _zz_3192_[48];
  assign _zz_3242_ = _zz_3192_[49];
  assign _zz_3243_ = _zz_3192_[50];
  assign _zz_3244_ = _zz_3192_[51];
  assign _zz_3245_ = _zz_3192_[52];
  assign _zz_3246_ = _zz_3192_[53];
  assign _zz_3247_ = _zz_3192_[54];
  assign _zz_3248_ = _zz_3192_[55];
  assign _zz_3249_ = _zz_3192_[56];
  assign _zz_3250_ = _zz_3192_[57];
  assign _zz_3251_ = _zz_3192_[58];
  assign _zz_3252_ = _zz_3192_[59];
  assign _zz_3253_ = _zz_3192_[60];
  assign _zz_3254_ = _zz_3192_[61];
  assign _zz_3255_ = _zz_3192_[62];
  assign _zz_3256_ = _zz_3192_[63];
  assign _zz_3257_ = (((32'h00000740 <= load_data_area_current_addr) && (load_data_area_current_addr < 32'h00000780)) ? _zz_9__regNext : {_zz_4526_,_zz_4527_});
  assign _zz_3258_ = _zz_3257_[15 : 0];
  assign _zz_3259_ = _zz_3257_[31 : 16];
  assign _zz_3260_ = _zz_4613_[5:0];
  assign _zz_3261_ = ({63'd0,(1'b1)} <<< _zz_3260_);
  assign _zz_3262_ = _zz_3261_[0];
  assign _zz_3263_ = _zz_3261_[1];
  assign _zz_3264_ = _zz_3261_[2];
  assign _zz_3265_ = _zz_3261_[3];
  assign _zz_3266_ = _zz_3261_[4];
  assign _zz_3267_ = _zz_3261_[5];
  assign _zz_3268_ = _zz_3261_[6];
  assign _zz_3269_ = _zz_3261_[7];
  assign _zz_3270_ = _zz_3261_[8];
  assign _zz_3271_ = _zz_3261_[9];
  assign _zz_3272_ = _zz_3261_[10];
  assign _zz_3273_ = _zz_3261_[11];
  assign _zz_3274_ = _zz_3261_[12];
  assign _zz_3275_ = _zz_3261_[13];
  assign _zz_3276_ = _zz_3261_[14];
  assign _zz_3277_ = _zz_3261_[15];
  assign _zz_3278_ = _zz_3261_[16];
  assign _zz_3279_ = _zz_3261_[17];
  assign _zz_3280_ = _zz_3261_[18];
  assign _zz_3281_ = _zz_3261_[19];
  assign _zz_3282_ = _zz_3261_[20];
  assign _zz_3283_ = _zz_3261_[21];
  assign _zz_3284_ = _zz_3261_[22];
  assign _zz_3285_ = _zz_3261_[23];
  assign _zz_3286_ = _zz_3261_[24];
  assign _zz_3287_ = _zz_3261_[25];
  assign _zz_3288_ = _zz_3261_[26];
  assign _zz_3289_ = _zz_3261_[27];
  assign _zz_3290_ = _zz_3261_[28];
  assign _zz_3291_ = _zz_3261_[29];
  assign _zz_3292_ = _zz_3261_[30];
  assign _zz_3293_ = _zz_3261_[31];
  assign _zz_3294_ = _zz_3261_[32];
  assign _zz_3295_ = _zz_3261_[33];
  assign _zz_3296_ = _zz_3261_[34];
  assign _zz_3297_ = _zz_3261_[35];
  assign _zz_3298_ = _zz_3261_[36];
  assign _zz_3299_ = _zz_3261_[37];
  assign _zz_3300_ = _zz_3261_[38];
  assign _zz_3301_ = _zz_3261_[39];
  assign _zz_3302_ = _zz_3261_[40];
  assign _zz_3303_ = _zz_3261_[41];
  assign _zz_3304_ = _zz_3261_[42];
  assign _zz_3305_ = _zz_3261_[43];
  assign _zz_3306_ = _zz_3261_[44];
  assign _zz_3307_ = _zz_3261_[45];
  assign _zz_3308_ = _zz_3261_[46];
  assign _zz_3309_ = _zz_3261_[47];
  assign _zz_3310_ = _zz_3261_[48];
  assign _zz_3311_ = _zz_3261_[49];
  assign _zz_3312_ = _zz_3261_[50];
  assign _zz_3313_ = _zz_3261_[51];
  assign _zz_3314_ = _zz_3261_[52];
  assign _zz_3315_ = _zz_3261_[53];
  assign _zz_3316_ = _zz_3261_[54];
  assign _zz_3317_ = _zz_3261_[55];
  assign _zz_3318_ = _zz_3261_[56];
  assign _zz_3319_ = _zz_3261_[57];
  assign _zz_3320_ = _zz_3261_[58];
  assign _zz_3321_ = _zz_3261_[59];
  assign _zz_3322_ = _zz_3261_[60];
  assign _zz_3323_ = _zz_3261_[61];
  assign _zz_3324_ = _zz_3261_[62];
  assign _zz_3325_ = _zz_3261_[63];
  assign _zz_3326_ = (((32'h00000ec0 <= load_data_area_current_addr) && (load_data_area_current_addr < 32'h00000f00)) ? _zz_9__regNext : {_zz_4528_,_zz_4529_});
  assign _zz_3327_ = _zz_3326_[15 : 0];
  assign _zz_3328_ = _zz_3326_[31 : 16];
  assign _zz_3329_ = _zz_4614_[5:0];
  assign _zz_3330_ = ({63'd0,(1'b1)} <<< _zz_3329_);
  assign _zz_3331_ = _zz_3330_[0];
  assign _zz_3332_ = _zz_3330_[1];
  assign _zz_3333_ = _zz_3330_[2];
  assign _zz_3334_ = _zz_3330_[3];
  assign _zz_3335_ = _zz_3330_[4];
  assign _zz_3336_ = _zz_3330_[5];
  assign _zz_3337_ = _zz_3330_[6];
  assign _zz_3338_ = _zz_3330_[7];
  assign _zz_3339_ = _zz_3330_[8];
  assign _zz_3340_ = _zz_3330_[9];
  assign _zz_3341_ = _zz_3330_[10];
  assign _zz_3342_ = _zz_3330_[11];
  assign _zz_3343_ = _zz_3330_[12];
  assign _zz_3344_ = _zz_3330_[13];
  assign _zz_3345_ = _zz_3330_[14];
  assign _zz_3346_ = _zz_3330_[15];
  assign _zz_3347_ = _zz_3330_[16];
  assign _zz_3348_ = _zz_3330_[17];
  assign _zz_3349_ = _zz_3330_[18];
  assign _zz_3350_ = _zz_3330_[19];
  assign _zz_3351_ = _zz_3330_[20];
  assign _zz_3352_ = _zz_3330_[21];
  assign _zz_3353_ = _zz_3330_[22];
  assign _zz_3354_ = _zz_3330_[23];
  assign _zz_3355_ = _zz_3330_[24];
  assign _zz_3356_ = _zz_3330_[25];
  assign _zz_3357_ = _zz_3330_[26];
  assign _zz_3358_ = _zz_3330_[27];
  assign _zz_3359_ = _zz_3330_[28];
  assign _zz_3360_ = _zz_3330_[29];
  assign _zz_3361_ = _zz_3330_[30];
  assign _zz_3362_ = _zz_3330_[31];
  assign _zz_3363_ = _zz_3330_[32];
  assign _zz_3364_ = _zz_3330_[33];
  assign _zz_3365_ = _zz_3330_[34];
  assign _zz_3366_ = _zz_3330_[35];
  assign _zz_3367_ = _zz_3330_[36];
  assign _zz_3368_ = _zz_3330_[37];
  assign _zz_3369_ = _zz_3330_[38];
  assign _zz_3370_ = _zz_3330_[39];
  assign _zz_3371_ = _zz_3330_[40];
  assign _zz_3372_ = _zz_3330_[41];
  assign _zz_3373_ = _zz_3330_[42];
  assign _zz_3374_ = _zz_3330_[43];
  assign _zz_3375_ = _zz_3330_[44];
  assign _zz_3376_ = _zz_3330_[45];
  assign _zz_3377_ = _zz_3330_[46];
  assign _zz_3378_ = _zz_3330_[47];
  assign _zz_3379_ = _zz_3330_[48];
  assign _zz_3380_ = _zz_3330_[49];
  assign _zz_3381_ = _zz_3330_[50];
  assign _zz_3382_ = _zz_3330_[51];
  assign _zz_3383_ = _zz_3330_[52];
  assign _zz_3384_ = _zz_3330_[53];
  assign _zz_3385_ = _zz_3330_[54];
  assign _zz_3386_ = _zz_3330_[55];
  assign _zz_3387_ = _zz_3330_[56];
  assign _zz_3388_ = _zz_3330_[57];
  assign _zz_3389_ = _zz_3330_[58];
  assign _zz_3390_ = _zz_3330_[59];
  assign _zz_3391_ = _zz_3330_[60];
  assign _zz_3392_ = _zz_3330_[61];
  assign _zz_3393_ = _zz_3330_[62];
  assign _zz_3394_ = _zz_3330_[63];
  assign _zz_3395_ = (((32'h00000b40 <= load_data_area_current_addr) && (load_data_area_current_addr < 32'h00000b80)) ? _zz_9__regNext : {_zz_4530_,_zz_4531_});
  assign _zz_3396_ = _zz_3395_[15 : 0];
  assign _zz_3397_ = _zz_3395_[31 : 16];
  assign _zz_3398_ = _zz_4615_[5:0];
  assign _zz_3399_ = ({63'd0,(1'b1)} <<< _zz_3398_);
  assign _zz_3400_ = _zz_3399_[0];
  assign _zz_3401_ = _zz_3399_[1];
  assign _zz_3402_ = _zz_3399_[2];
  assign _zz_3403_ = _zz_3399_[3];
  assign _zz_3404_ = _zz_3399_[4];
  assign _zz_3405_ = _zz_3399_[5];
  assign _zz_3406_ = _zz_3399_[6];
  assign _zz_3407_ = _zz_3399_[7];
  assign _zz_3408_ = _zz_3399_[8];
  assign _zz_3409_ = _zz_3399_[9];
  assign _zz_3410_ = _zz_3399_[10];
  assign _zz_3411_ = _zz_3399_[11];
  assign _zz_3412_ = _zz_3399_[12];
  assign _zz_3413_ = _zz_3399_[13];
  assign _zz_3414_ = _zz_3399_[14];
  assign _zz_3415_ = _zz_3399_[15];
  assign _zz_3416_ = _zz_3399_[16];
  assign _zz_3417_ = _zz_3399_[17];
  assign _zz_3418_ = _zz_3399_[18];
  assign _zz_3419_ = _zz_3399_[19];
  assign _zz_3420_ = _zz_3399_[20];
  assign _zz_3421_ = _zz_3399_[21];
  assign _zz_3422_ = _zz_3399_[22];
  assign _zz_3423_ = _zz_3399_[23];
  assign _zz_3424_ = _zz_3399_[24];
  assign _zz_3425_ = _zz_3399_[25];
  assign _zz_3426_ = _zz_3399_[26];
  assign _zz_3427_ = _zz_3399_[27];
  assign _zz_3428_ = _zz_3399_[28];
  assign _zz_3429_ = _zz_3399_[29];
  assign _zz_3430_ = _zz_3399_[30];
  assign _zz_3431_ = _zz_3399_[31];
  assign _zz_3432_ = _zz_3399_[32];
  assign _zz_3433_ = _zz_3399_[33];
  assign _zz_3434_ = _zz_3399_[34];
  assign _zz_3435_ = _zz_3399_[35];
  assign _zz_3436_ = _zz_3399_[36];
  assign _zz_3437_ = _zz_3399_[37];
  assign _zz_3438_ = _zz_3399_[38];
  assign _zz_3439_ = _zz_3399_[39];
  assign _zz_3440_ = _zz_3399_[40];
  assign _zz_3441_ = _zz_3399_[41];
  assign _zz_3442_ = _zz_3399_[42];
  assign _zz_3443_ = _zz_3399_[43];
  assign _zz_3444_ = _zz_3399_[44];
  assign _zz_3445_ = _zz_3399_[45];
  assign _zz_3446_ = _zz_3399_[46];
  assign _zz_3447_ = _zz_3399_[47];
  assign _zz_3448_ = _zz_3399_[48];
  assign _zz_3449_ = _zz_3399_[49];
  assign _zz_3450_ = _zz_3399_[50];
  assign _zz_3451_ = _zz_3399_[51];
  assign _zz_3452_ = _zz_3399_[52];
  assign _zz_3453_ = _zz_3399_[53];
  assign _zz_3454_ = _zz_3399_[54];
  assign _zz_3455_ = _zz_3399_[55];
  assign _zz_3456_ = _zz_3399_[56];
  assign _zz_3457_ = _zz_3399_[57];
  assign _zz_3458_ = _zz_3399_[58];
  assign _zz_3459_ = _zz_3399_[59];
  assign _zz_3460_ = _zz_3399_[60];
  assign _zz_3461_ = _zz_3399_[61];
  assign _zz_3462_ = _zz_3399_[62];
  assign _zz_3463_ = _zz_3399_[63];
  assign _zz_3464_ = (((32'h00000100 <= load_data_area_current_addr) && (load_data_area_current_addr < 32'h00000140)) ? _zz_9__regNext : {_zz_4532_,_zz_4533_});
  assign _zz_3465_ = _zz_3464_[15 : 0];
  assign _zz_3466_ = _zz_3464_[31 : 16];
  assign _zz_3467_ = _zz_4616_[5:0];
  assign _zz_3468_ = ({63'd0,(1'b1)} <<< _zz_3467_);
  assign _zz_3469_ = _zz_3468_[0];
  assign _zz_3470_ = _zz_3468_[1];
  assign _zz_3471_ = _zz_3468_[2];
  assign _zz_3472_ = _zz_3468_[3];
  assign _zz_3473_ = _zz_3468_[4];
  assign _zz_3474_ = _zz_3468_[5];
  assign _zz_3475_ = _zz_3468_[6];
  assign _zz_3476_ = _zz_3468_[7];
  assign _zz_3477_ = _zz_3468_[8];
  assign _zz_3478_ = _zz_3468_[9];
  assign _zz_3479_ = _zz_3468_[10];
  assign _zz_3480_ = _zz_3468_[11];
  assign _zz_3481_ = _zz_3468_[12];
  assign _zz_3482_ = _zz_3468_[13];
  assign _zz_3483_ = _zz_3468_[14];
  assign _zz_3484_ = _zz_3468_[15];
  assign _zz_3485_ = _zz_3468_[16];
  assign _zz_3486_ = _zz_3468_[17];
  assign _zz_3487_ = _zz_3468_[18];
  assign _zz_3488_ = _zz_3468_[19];
  assign _zz_3489_ = _zz_3468_[20];
  assign _zz_3490_ = _zz_3468_[21];
  assign _zz_3491_ = _zz_3468_[22];
  assign _zz_3492_ = _zz_3468_[23];
  assign _zz_3493_ = _zz_3468_[24];
  assign _zz_3494_ = _zz_3468_[25];
  assign _zz_3495_ = _zz_3468_[26];
  assign _zz_3496_ = _zz_3468_[27];
  assign _zz_3497_ = _zz_3468_[28];
  assign _zz_3498_ = _zz_3468_[29];
  assign _zz_3499_ = _zz_3468_[30];
  assign _zz_3500_ = _zz_3468_[31];
  assign _zz_3501_ = _zz_3468_[32];
  assign _zz_3502_ = _zz_3468_[33];
  assign _zz_3503_ = _zz_3468_[34];
  assign _zz_3504_ = _zz_3468_[35];
  assign _zz_3505_ = _zz_3468_[36];
  assign _zz_3506_ = _zz_3468_[37];
  assign _zz_3507_ = _zz_3468_[38];
  assign _zz_3508_ = _zz_3468_[39];
  assign _zz_3509_ = _zz_3468_[40];
  assign _zz_3510_ = _zz_3468_[41];
  assign _zz_3511_ = _zz_3468_[42];
  assign _zz_3512_ = _zz_3468_[43];
  assign _zz_3513_ = _zz_3468_[44];
  assign _zz_3514_ = _zz_3468_[45];
  assign _zz_3515_ = _zz_3468_[46];
  assign _zz_3516_ = _zz_3468_[47];
  assign _zz_3517_ = _zz_3468_[48];
  assign _zz_3518_ = _zz_3468_[49];
  assign _zz_3519_ = _zz_3468_[50];
  assign _zz_3520_ = _zz_3468_[51];
  assign _zz_3521_ = _zz_3468_[52];
  assign _zz_3522_ = _zz_3468_[53];
  assign _zz_3523_ = _zz_3468_[54];
  assign _zz_3524_ = _zz_3468_[55];
  assign _zz_3525_ = _zz_3468_[56];
  assign _zz_3526_ = _zz_3468_[57];
  assign _zz_3527_ = _zz_3468_[58];
  assign _zz_3528_ = _zz_3468_[59];
  assign _zz_3529_ = _zz_3468_[60];
  assign _zz_3530_ = _zz_3468_[61];
  assign _zz_3531_ = _zz_3468_[62];
  assign _zz_3532_ = _zz_3468_[63];
  assign _zz_3533_ = (((32'h00000cc0 <= load_data_area_current_addr) && (load_data_area_current_addr < 32'h00000d00)) ? _zz_9__regNext : {_zz_4534_,_zz_4535_});
  assign _zz_3534_ = _zz_3533_[15 : 0];
  assign _zz_3535_ = _zz_3533_[31 : 16];
  assign _zz_3536_ = _zz_4617_[5:0];
  assign _zz_3537_ = ({63'd0,(1'b1)} <<< _zz_3536_);
  assign _zz_3538_ = _zz_3537_[0];
  assign _zz_3539_ = _zz_3537_[1];
  assign _zz_3540_ = _zz_3537_[2];
  assign _zz_3541_ = _zz_3537_[3];
  assign _zz_3542_ = _zz_3537_[4];
  assign _zz_3543_ = _zz_3537_[5];
  assign _zz_3544_ = _zz_3537_[6];
  assign _zz_3545_ = _zz_3537_[7];
  assign _zz_3546_ = _zz_3537_[8];
  assign _zz_3547_ = _zz_3537_[9];
  assign _zz_3548_ = _zz_3537_[10];
  assign _zz_3549_ = _zz_3537_[11];
  assign _zz_3550_ = _zz_3537_[12];
  assign _zz_3551_ = _zz_3537_[13];
  assign _zz_3552_ = _zz_3537_[14];
  assign _zz_3553_ = _zz_3537_[15];
  assign _zz_3554_ = _zz_3537_[16];
  assign _zz_3555_ = _zz_3537_[17];
  assign _zz_3556_ = _zz_3537_[18];
  assign _zz_3557_ = _zz_3537_[19];
  assign _zz_3558_ = _zz_3537_[20];
  assign _zz_3559_ = _zz_3537_[21];
  assign _zz_3560_ = _zz_3537_[22];
  assign _zz_3561_ = _zz_3537_[23];
  assign _zz_3562_ = _zz_3537_[24];
  assign _zz_3563_ = _zz_3537_[25];
  assign _zz_3564_ = _zz_3537_[26];
  assign _zz_3565_ = _zz_3537_[27];
  assign _zz_3566_ = _zz_3537_[28];
  assign _zz_3567_ = _zz_3537_[29];
  assign _zz_3568_ = _zz_3537_[30];
  assign _zz_3569_ = _zz_3537_[31];
  assign _zz_3570_ = _zz_3537_[32];
  assign _zz_3571_ = _zz_3537_[33];
  assign _zz_3572_ = _zz_3537_[34];
  assign _zz_3573_ = _zz_3537_[35];
  assign _zz_3574_ = _zz_3537_[36];
  assign _zz_3575_ = _zz_3537_[37];
  assign _zz_3576_ = _zz_3537_[38];
  assign _zz_3577_ = _zz_3537_[39];
  assign _zz_3578_ = _zz_3537_[40];
  assign _zz_3579_ = _zz_3537_[41];
  assign _zz_3580_ = _zz_3537_[42];
  assign _zz_3581_ = _zz_3537_[43];
  assign _zz_3582_ = _zz_3537_[44];
  assign _zz_3583_ = _zz_3537_[45];
  assign _zz_3584_ = _zz_3537_[46];
  assign _zz_3585_ = _zz_3537_[47];
  assign _zz_3586_ = _zz_3537_[48];
  assign _zz_3587_ = _zz_3537_[49];
  assign _zz_3588_ = _zz_3537_[50];
  assign _zz_3589_ = _zz_3537_[51];
  assign _zz_3590_ = _zz_3537_[52];
  assign _zz_3591_ = _zz_3537_[53];
  assign _zz_3592_ = _zz_3537_[54];
  assign _zz_3593_ = _zz_3537_[55];
  assign _zz_3594_ = _zz_3537_[56];
  assign _zz_3595_ = _zz_3537_[57];
  assign _zz_3596_ = _zz_3537_[58];
  assign _zz_3597_ = _zz_3537_[59];
  assign _zz_3598_ = _zz_3537_[60];
  assign _zz_3599_ = _zz_3537_[61];
  assign _zz_3600_ = _zz_3537_[62];
  assign _zz_3601_ = _zz_3537_[63];
  assign _zz_3602_ = (((32'h00000440 <= load_data_area_current_addr) && (load_data_area_current_addr < 32'h00000480)) ? _zz_9__regNext : {_zz_4536_,_zz_4537_});
  assign _zz_3603_ = _zz_3602_[15 : 0];
  assign _zz_3604_ = _zz_3602_[31 : 16];
  assign _zz_3605_ = _zz_4618_[5:0];
  assign _zz_3606_ = ({63'd0,(1'b1)} <<< _zz_3605_);
  assign _zz_3607_ = _zz_3606_[0];
  assign _zz_3608_ = _zz_3606_[1];
  assign _zz_3609_ = _zz_3606_[2];
  assign _zz_3610_ = _zz_3606_[3];
  assign _zz_3611_ = _zz_3606_[4];
  assign _zz_3612_ = _zz_3606_[5];
  assign _zz_3613_ = _zz_3606_[6];
  assign _zz_3614_ = _zz_3606_[7];
  assign _zz_3615_ = _zz_3606_[8];
  assign _zz_3616_ = _zz_3606_[9];
  assign _zz_3617_ = _zz_3606_[10];
  assign _zz_3618_ = _zz_3606_[11];
  assign _zz_3619_ = _zz_3606_[12];
  assign _zz_3620_ = _zz_3606_[13];
  assign _zz_3621_ = _zz_3606_[14];
  assign _zz_3622_ = _zz_3606_[15];
  assign _zz_3623_ = _zz_3606_[16];
  assign _zz_3624_ = _zz_3606_[17];
  assign _zz_3625_ = _zz_3606_[18];
  assign _zz_3626_ = _zz_3606_[19];
  assign _zz_3627_ = _zz_3606_[20];
  assign _zz_3628_ = _zz_3606_[21];
  assign _zz_3629_ = _zz_3606_[22];
  assign _zz_3630_ = _zz_3606_[23];
  assign _zz_3631_ = _zz_3606_[24];
  assign _zz_3632_ = _zz_3606_[25];
  assign _zz_3633_ = _zz_3606_[26];
  assign _zz_3634_ = _zz_3606_[27];
  assign _zz_3635_ = _zz_3606_[28];
  assign _zz_3636_ = _zz_3606_[29];
  assign _zz_3637_ = _zz_3606_[30];
  assign _zz_3638_ = _zz_3606_[31];
  assign _zz_3639_ = _zz_3606_[32];
  assign _zz_3640_ = _zz_3606_[33];
  assign _zz_3641_ = _zz_3606_[34];
  assign _zz_3642_ = _zz_3606_[35];
  assign _zz_3643_ = _zz_3606_[36];
  assign _zz_3644_ = _zz_3606_[37];
  assign _zz_3645_ = _zz_3606_[38];
  assign _zz_3646_ = _zz_3606_[39];
  assign _zz_3647_ = _zz_3606_[40];
  assign _zz_3648_ = _zz_3606_[41];
  assign _zz_3649_ = _zz_3606_[42];
  assign _zz_3650_ = _zz_3606_[43];
  assign _zz_3651_ = _zz_3606_[44];
  assign _zz_3652_ = _zz_3606_[45];
  assign _zz_3653_ = _zz_3606_[46];
  assign _zz_3654_ = _zz_3606_[47];
  assign _zz_3655_ = _zz_3606_[48];
  assign _zz_3656_ = _zz_3606_[49];
  assign _zz_3657_ = _zz_3606_[50];
  assign _zz_3658_ = _zz_3606_[51];
  assign _zz_3659_ = _zz_3606_[52];
  assign _zz_3660_ = _zz_3606_[53];
  assign _zz_3661_ = _zz_3606_[54];
  assign _zz_3662_ = _zz_3606_[55];
  assign _zz_3663_ = _zz_3606_[56];
  assign _zz_3664_ = _zz_3606_[57];
  assign _zz_3665_ = _zz_3606_[58];
  assign _zz_3666_ = _zz_3606_[59];
  assign _zz_3667_ = _zz_3606_[60];
  assign _zz_3668_ = _zz_3606_[61];
  assign _zz_3669_ = _zz_3606_[62];
  assign _zz_3670_ = _zz_3606_[63];
  assign _zz_3671_ = (((32'h00000540 <= load_data_area_current_addr) && (load_data_area_current_addr < 32'h00000580)) ? _zz_9__regNext : {_zz_4538_,_zz_4539_});
  assign _zz_3672_ = _zz_3671_[15 : 0];
  assign _zz_3673_ = _zz_3671_[31 : 16];
  assign _zz_3674_ = _zz_4619_[5:0];
  assign _zz_3675_ = ({63'd0,(1'b1)} <<< _zz_3674_);
  assign _zz_3676_ = _zz_3675_[0];
  assign _zz_3677_ = _zz_3675_[1];
  assign _zz_3678_ = _zz_3675_[2];
  assign _zz_3679_ = _zz_3675_[3];
  assign _zz_3680_ = _zz_3675_[4];
  assign _zz_3681_ = _zz_3675_[5];
  assign _zz_3682_ = _zz_3675_[6];
  assign _zz_3683_ = _zz_3675_[7];
  assign _zz_3684_ = _zz_3675_[8];
  assign _zz_3685_ = _zz_3675_[9];
  assign _zz_3686_ = _zz_3675_[10];
  assign _zz_3687_ = _zz_3675_[11];
  assign _zz_3688_ = _zz_3675_[12];
  assign _zz_3689_ = _zz_3675_[13];
  assign _zz_3690_ = _zz_3675_[14];
  assign _zz_3691_ = _zz_3675_[15];
  assign _zz_3692_ = _zz_3675_[16];
  assign _zz_3693_ = _zz_3675_[17];
  assign _zz_3694_ = _zz_3675_[18];
  assign _zz_3695_ = _zz_3675_[19];
  assign _zz_3696_ = _zz_3675_[20];
  assign _zz_3697_ = _zz_3675_[21];
  assign _zz_3698_ = _zz_3675_[22];
  assign _zz_3699_ = _zz_3675_[23];
  assign _zz_3700_ = _zz_3675_[24];
  assign _zz_3701_ = _zz_3675_[25];
  assign _zz_3702_ = _zz_3675_[26];
  assign _zz_3703_ = _zz_3675_[27];
  assign _zz_3704_ = _zz_3675_[28];
  assign _zz_3705_ = _zz_3675_[29];
  assign _zz_3706_ = _zz_3675_[30];
  assign _zz_3707_ = _zz_3675_[31];
  assign _zz_3708_ = _zz_3675_[32];
  assign _zz_3709_ = _zz_3675_[33];
  assign _zz_3710_ = _zz_3675_[34];
  assign _zz_3711_ = _zz_3675_[35];
  assign _zz_3712_ = _zz_3675_[36];
  assign _zz_3713_ = _zz_3675_[37];
  assign _zz_3714_ = _zz_3675_[38];
  assign _zz_3715_ = _zz_3675_[39];
  assign _zz_3716_ = _zz_3675_[40];
  assign _zz_3717_ = _zz_3675_[41];
  assign _zz_3718_ = _zz_3675_[42];
  assign _zz_3719_ = _zz_3675_[43];
  assign _zz_3720_ = _zz_3675_[44];
  assign _zz_3721_ = _zz_3675_[45];
  assign _zz_3722_ = _zz_3675_[46];
  assign _zz_3723_ = _zz_3675_[47];
  assign _zz_3724_ = _zz_3675_[48];
  assign _zz_3725_ = _zz_3675_[49];
  assign _zz_3726_ = _zz_3675_[50];
  assign _zz_3727_ = _zz_3675_[51];
  assign _zz_3728_ = _zz_3675_[52];
  assign _zz_3729_ = _zz_3675_[53];
  assign _zz_3730_ = _zz_3675_[54];
  assign _zz_3731_ = _zz_3675_[55];
  assign _zz_3732_ = _zz_3675_[56];
  assign _zz_3733_ = _zz_3675_[57];
  assign _zz_3734_ = _zz_3675_[58];
  assign _zz_3735_ = _zz_3675_[59];
  assign _zz_3736_ = _zz_3675_[60];
  assign _zz_3737_ = _zz_3675_[61];
  assign _zz_3738_ = _zz_3675_[62];
  assign _zz_3739_ = _zz_3675_[63];
  assign _zz_3740_ = (((32'h000008c0 <= load_data_area_current_addr) && (load_data_area_current_addr < 32'h00000900)) ? _zz_9__regNext : {_zz_4540_,_zz_4541_});
  assign _zz_3741_ = _zz_3740_[15 : 0];
  assign _zz_3742_ = _zz_3740_[31 : 16];
  assign _zz_3743_ = _zz_4620_[5:0];
  assign _zz_3744_ = ({63'd0,(1'b1)} <<< _zz_3743_);
  assign _zz_3745_ = _zz_3744_[0];
  assign _zz_3746_ = _zz_3744_[1];
  assign _zz_3747_ = _zz_3744_[2];
  assign _zz_3748_ = _zz_3744_[3];
  assign _zz_3749_ = _zz_3744_[4];
  assign _zz_3750_ = _zz_3744_[5];
  assign _zz_3751_ = _zz_3744_[6];
  assign _zz_3752_ = _zz_3744_[7];
  assign _zz_3753_ = _zz_3744_[8];
  assign _zz_3754_ = _zz_3744_[9];
  assign _zz_3755_ = _zz_3744_[10];
  assign _zz_3756_ = _zz_3744_[11];
  assign _zz_3757_ = _zz_3744_[12];
  assign _zz_3758_ = _zz_3744_[13];
  assign _zz_3759_ = _zz_3744_[14];
  assign _zz_3760_ = _zz_3744_[15];
  assign _zz_3761_ = _zz_3744_[16];
  assign _zz_3762_ = _zz_3744_[17];
  assign _zz_3763_ = _zz_3744_[18];
  assign _zz_3764_ = _zz_3744_[19];
  assign _zz_3765_ = _zz_3744_[20];
  assign _zz_3766_ = _zz_3744_[21];
  assign _zz_3767_ = _zz_3744_[22];
  assign _zz_3768_ = _zz_3744_[23];
  assign _zz_3769_ = _zz_3744_[24];
  assign _zz_3770_ = _zz_3744_[25];
  assign _zz_3771_ = _zz_3744_[26];
  assign _zz_3772_ = _zz_3744_[27];
  assign _zz_3773_ = _zz_3744_[28];
  assign _zz_3774_ = _zz_3744_[29];
  assign _zz_3775_ = _zz_3744_[30];
  assign _zz_3776_ = _zz_3744_[31];
  assign _zz_3777_ = _zz_3744_[32];
  assign _zz_3778_ = _zz_3744_[33];
  assign _zz_3779_ = _zz_3744_[34];
  assign _zz_3780_ = _zz_3744_[35];
  assign _zz_3781_ = _zz_3744_[36];
  assign _zz_3782_ = _zz_3744_[37];
  assign _zz_3783_ = _zz_3744_[38];
  assign _zz_3784_ = _zz_3744_[39];
  assign _zz_3785_ = _zz_3744_[40];
  assign _zz_3786_ = _zz_3744_[41];
  assign _zz_3787_ = _zz_3744_[42];
  assign _zz_3788_ = _zz_3744_[43];
  assign _zz_3789_ = _zz_3744_[44];
  assign _zz_3790_ = _zz_3744_[45];
  assign _zz_3791_ = _zz_3744_[46];
  assign _zz_3792_ = _zz_3744_[47];
  assign _zz_3793_ = _zz_3744_[48];
  assign _zz_3794_ = _zz_3744_[49];
  assign _zz_3795_ = _zz_3744_[50];
  assign _zz_3796_ = _zz_3744_[51];
  assign _zz_3797_ = _zz_3744_[52];
  assign _zz_3798_ = _zz_3744_[53];
  assign _zz_3799_ = _zz_3744_[54];
  assign _zz_3800_ = _zz_3744_[55];
  assign _zz_3801_ = _zz_3744_[56];
  assign _zz_3802_ = _zz_3744_[57];
  assign _zz_3803_ = _zz_3744_[58];
  assign _zz_3804_ = _zz_3744_[59];
  assign _zz_3805_ = _zz_3744_[60];
  assign _zz_3806_ = _zz_3744_[61];
  assign _zz_3807_ = _zz_3744_[62];
  assign _zz_3808_ = _zz_3744_[63];
  assign _zz_3809_ = (((32'h00000a80 <= load_data_area_current_addr) && (load_data_area_current_addr < 32'h00000ac0)) ? _zz_9__regNext : {_zz_4542_,_zz_4543_});
  assign _zz_3810_ = _zz_3809_[15 : 0];
  assign _zz_3811_ = _zz_3809_[31 : 16];
  assign _zz_3812_ = _zz_4621_[5:0];
  assign _zz_3813_ = ({63'd0,(1'b1)} <<< _zz_3812_);
  assign _zz_3814_ = _zz_3813_[0];
  assign _zz_3815_ = _zz_3813_[1];
  assign _zz_3816_ = _zz_3813_[2];
  assign _zz_3817_ = _zz_3813_[3];
  assign _zz_3818_ = _zz_3813_[4];
  assign _zz_3819_ = _zz_3813_[5];
  assign _zz_3820_ = _zz_3813_[6];
  assign _zz_3821_ = _zz_3813_[7];
  assign _zz_3822_ = _zz_3813_[8];
  assign _zz_3823_ = _zz_3813_[9];
  assign _zz_3824_ = _zz_3813_[10];
  assign _zz_3825_ = _zz_3813_[11];
  assign _zz_3826_ = _zz_3813_[12];
  assign _zz_3827_ = _zz_3813_[13];
  assign _zz_3828_ = _zz_3813_[14];
  assign _zz_3829_ = _zz_3813_[15];
  assign _zz_3830_ = _zz_3813_[16];
  assign _zz_3831_ = _zz_3813_[17];
  assign _zz_3832_ = _zz_3813_[18];
  assign _zz_3833_ = _zz_3813_[19];
  assign _zz_3834_ = _zz_3813_[20];
  assign _zz_3835_ = _zz_3813_[21];
  assign _zz_3836_ = _zz_3813_[22];
  assign _zz_3837_ = _zz_3813_[23];
  assign _zz_3838_ = _zz_3813_[24];
  assign _zz_3839_ = _zz_3813_[25];
  assign _zz_3840_ = _zz_3813_[26];
  assign _zz_3841_ = _zz_3813_[27];
  assign _zz_3842_ = _zz_3813_[28];
  assign _zz_3843_ = _zz_3813_[29];
  assign _zz_3844_ = _zz_3813_[30];
  assign _zz_3845_ = _zz_3813_[31];
  assign _zz_3846_ = _zz_3813_[32];
  assign _zz_3847_ = _zz_3813_[33];
  assign _zz_3848_ = _zz_3813_[34];
  assign _zz_3849_ = _zz_3813_[35];
  assign _zz_3850_ = _zz_3813_[36];
  assign _zz_3851_ = _zz_3813_[37];
  assign _zz_3852_ = _zz_3813_[38];
  assign _zz_3853_ = _zz_3813_[39];
  assign _zz_3854_ = _zz_3813_[40];
  assign _zz_3855_ = _zz_3813_[41];
  assign _zz_3856_ = _zz_3813_[42];
  assign _zz_3857_ = _zz_3813_[43];
  assign _zz_3858_ = _zz_3813_[44];
  assign _zz_3859_ = _zz_3813_[45];
  assign _zz_3860_ = _zz_3813_[46];
  assign _zz_3861_ = _zz_3813_[47];
  assign _zz_3862_ = _zz_3813_[48];
  assign _zz_3863_ = _zz_3813_[49];
  assign _zz_3864_ = _zz_3813_[50];
  assign _zz_3865_ = _zz_3813_[51];
  assign _zz_3866_ = _zz_3813_[52];
  assign _zz_3867_ = _zz_3813_[53];
  assign _zz_3868_ = _zz_3813_[54];
  assign _zz_3869_ = _zz_3813_[55];
  assign _zz_3870_ = _zz_3813_[56];
  assign _zz_3871_ = _zz_3813_[57];
  assign _zz_3872_ = _zz_3813_[58];
  assign _zz_3873_ = _zz_3813_[59];
  assign _zz_3874_ = _zz_3813_[60];
  assign _zz_3875_ = _zz_3813_[61];
  assign _zz_3876_ = _zz_3813_[62];
  assign _zz_3877_ = _zz_3813_[63];
  assign _zz_3878_ = (((32'h000007c0 <= load_data_area_current_addr) && (load_data_area_current_addr < 32'h00000800)) ? _zz_9__regNext : {_zz_4544_,_zz_4545_});
  assign _zz_3879_ = _zz_3878_[15 : 0];
  assign _zz_3880_ = _zz_3878_[31 : 16];
  assign _zz_3881_ = _zz_4622_[5:0];
  assign _zz_3882_ = ({63'd0,(1'b1)} <<< _zz_3881_);
  assign _zz_3883_ = _zz_3882_[0];
  assign _zz_3884_ = _zz_3882_[1];
  assign _zz_3885_ = _zz_3882_[2];
  assign _zz_3886_ = _zz_3882_[3];
  assign _zz_3887_ = _zz_3882_[4];
  assign _zz_3888_ = _zz_3882_[5];
  assign _zz_3889_ = _zz_3882_[6];
  assign _zz_3890_ = _zz_3882_[7];
  assign _zz_3891_ = _zz_3882_[8];
  assign _zz_3892_ = _zz_3882_[9];
  assign _zz_3893_ = _zz_3882_[10];
  assign _zz_3894_ = _zz_3882_[11];
  assign _zz_3895_ = _zz_3882_[12];
  assign _zz_3896_ = _zz_3882_[13];
  assign _zz_3897_ = _zz_3882_[14];
  assign _zz_3898_ = _zz_3882_[15];
  assign _zz_3899_ = _zz_3882_[16];
  assign _zz_3900_ = _zz_3882_[17];
  assign _zz_3901_ = _zz_3882_[18];
  assign _zz_3902_ = _zz_3882_[19];
  assign _zz_3903_ = _zz_3882_[20];
  assign _zz_3904_ = _zz_3882_[21];
  assign _zz_3905_ = _zz_3882_[22];
  assign _zz_3906_ = _zz_3882_[23];
  assign _zz_3907_ = _zz_3882_[24];
  assign _zz_3908_ = _zz_3882_[25];
  assign _zz_3909_ = _zz_3882_[26];
  assign _zz_3910_ = _zz_3882_[27];
  assign _zz_3911_ = _zz_3882_[28];
  assign _zz_3912_ = _zz_3882_[29];
  assign _zz_3913_ = _zz_3882_[30];
  assign _zz_3914_ = _zz_3882_[31];
  assign _zz_3915_ = _zz_3882_[32];
  assign _zz_3916_ = _zz_3882_[33];
  assign _zz_3917_ = _zz_3882_[34];
  assign _zz_3918_ = _zz_3882_[35];
  assign _zz_3919_ = _zz_3882_[36];
  assign _zz_3920_ = _zz_3882_[37];
  assign _zz_3921_ = _zz_3882_[38];
  assign _zz_3922_ = _zz_3882_[39];
  assign _zz_3923_ = _zz_3882_[40];
  assign _zz_3924_ = _zz_3882_[41];
  assign _zz_3925_ = _zz_3882_[42];
  assign _zz_3926_ = _zz_3882_[43];
  assign _zz_3927_ = _zz_3882_[44];
  assign _zz_3928_ = _zz_3882_[45];
  assign _zz_3929_ = _zz_3882_[46];
  assign _zz_3930_ = _zz_3882_[47];
  assign _zz_3931_ = _zz_3882_[48];
  assign _zz_3932_ = _zz_3882_[49];
  assign _zz_3933_ = _zz_3882_[50];
  assign _zz_3934_ = _zz_3882_[51];
  assign _zz_3935_ = _zz_3882_[52];
  assign _zz_3936_ = _zz_3882_[53];
  assign _zz_3937_ = _zz_3882_[54];
  assign _zz_3938_ = _zz_3882_[55];
  assign _zz_3939_ = _zz_3882_[56];
  assign _zz_3940_ = _zz_3882_[57];
  assign _zz_3941_ = _zz_3882_[58];
  assign _zz_3942_ = _zz_3882_[59];
  assign _zz_3943_ = _zz_3882_[60];
  assign _zz_3944_ = _zz_3882_[61];
  assign _zz_3945_ = _zz_3882_[62];
  assign _zz_3946_ = _zz_3882_[63];
  assign _zz_3947_ = (((32'h00000c00 <= load_data_area_current_addr) && (load_data_area_current_addr < 32'h00000c40)) ? _zz_9__regNext : {_zz_4546_,_zz_4547_});
  assign _zz_3948_ = _zz_3947_[15 : 0];
  assign _zz_3949_ = _zz_3947_[31 : 16];
  assign _zz_3950_ = _zz_4623_[5:0];
  assign _zz_3951_ = ({63'd0,(1'b1)} <<< _zz_3950_);
  assign _zz_3952_ = _zz_3951_[0];
  assign _zz_3953_ = _zz_3951_[1];
  assign _zz_3954_ = _zz_3951_[2];
  assign _zz_3955_ = _zz_3951_[3];
  assign _zz_3956_ = _zz_3951_[4];
  assign _zz_3957_ = _zz_3951_[5];
  assign _zz_3958_ = _zz_3951_[6];
  assign _zz_3959_ = _zz_3951_[7];
  assign _zz_3960_ = _zz_3951_[8];
  assign _zz_3961_ = _zz_3951_[9];
  assign _zz_3962_ = _zz_3951_[10];
  assign _zz_3963_ = _zz_3951_[11];
  assign _zz_3964_ = _zz_3951_[12];
  assign _zz_3965_ = _zz_3951_[13];
  assign _zz_3966_ = _zz_3951_[14];
  assign _zz_3967_ = _zz_3951_[15];
  assign _zz_3968_ = _zz_3951_[16];
  assign _zz_3969_ = _zz_3951_[17];
  assign _zz_3970_ = _zz_3951_[18];
  assign _zz_3971_ = _zz_3951_[19];
  assign _zz_3972_ = _zz_3951_[20];
  assign _zz_3973_ = _zz_3951_[21];
  assign _zz_3974_ = _zz_3951_[22];
  assign _zz_3975_ = _zz_3951_[23];
  assign _zz_3976_ = _zz_3951_[24];
  assign _zz_3977_ = _zz_3951_[25];
  assign _zz_3978_ = _zz_3951_[26];
  assign _zz_3979_ = _zz_3951_[27];
  assign _zz_3980_ = _zz_3951_[28];
  assign _zz_3981_ = _zz_3951_[29];
  assign _zz_3982_ = _zz_3951_[30];
  assign _zz_3983_ = _zz_3951_[31];
  assign _zz_3984_ = _zz_3951_[32];
  assign _zz_3985_ = _zz_3951_[33];
  assign _zz_3986_ = _zz_3951_[34];
  assign _zz_3987_ = _zz_3951_[35];
  assign _zz_3988_ = _zz_3951_[36];
  assign _zz_3989_ = _zz_3951_[37];
  assign _zz_3990_ = _zz_3951_[38];
  assign _zz_3991_ = _zz_3951_[39];
  assign _zz_3992_ = _zz_3951_[40];
  assign _zz_3993_ = _zz_3951_[41];
  assign _zz_3994_ = _zz_3951_[42];
  assign _zz_3995_ = _zz_3951_[43];
  assign _zz_3996_ = _zz_3951_[44];
  assign _zz_3997_ = _zz_3951_[45];
  assign _zz_3998_ = _zz_3951_[46];
  assign _zz_3999_ = _zz_3951_[47];
  assign _zz_4000_ = _zz_3951_[48];
  assign _zz_4001_ = _zz_3951_[49];
  assign _zz_4002_ = _zz_3951_[50];
  assign _zz_4003_ = _zz_3951_[51];
  assign _zz_4004_ = _zz_3951_[52];
  assign _zz_4005_ = _zz_3951_[53];
  assign _zz_4006_ = _zz_3951_[54];
  assign _zz_4007_ = _zz_3951_[55];
  assign _zz_4008_ = _zz_3951_[56];
  assign _zz_4009_ = _zz_3951_[57];
  assign _zz_4010_ = _zz_3951_[58];
  assign _zz_4011_ = _zz_3951_[59];
  assign _zz_4012_ = _zz_3951_[60];
  assign _zz_4013_ = _zz_3951_[61];
  assign _zz_4014_ = _zz_3951_[62];
  assign _zz_4015_ = _zz_3951_[63];
  assign _zz_4016_ = (((32'h00000940 <= load_data_area_current_addr) && (load_data_area_current_addr < 32'h00000980)) ? _zz_9__regNext : {_zz_4548_,_zz_4549_});
  assign _zz_4017_ = _zz_4016_[15 : 0];
  assign _zz_4018_ = _zz_4016_[31 : 16];
  assign _zz_4019_ = _zz_4624_[5:0];
  assign _zz_4020_ = ({63'd0,(1'b1)} <<< _zz_4019_);
  assign _zz_4021_ = _zz_4020_[0];
  assign _zz_4022_ = _zz_4020_[1];
  assign _zz_4023_ = _zz_4020_[2];
  assign _zz_4024_ = _zz_4020_[3];
  assign _zz_4025_ = _zz_4020_[4];
  assign _zz_4026_ = _zz_4020_[5];
  assign _zz_4027_ = _zz_4020_[6];
  assign _zz_4028_ = _zz_4020_[7];
  assign _zz_4029_ = _zz_4020_[8];
  assign _zz_4030_ = _zz_4020_[9];
  assign _zz_4031_ = _zz_4020_[10];
  assign _zz_4032_ = _zz_4020_[11];
  assign _zz_4033_ = _zz_4020_[12];
  assign _zz_4034_ = _zz_4020_[13];
  assign _zz_4035_ = _zz_4020_[14];
  assign _zz_4036_ = _zz_4020_[15];
  assign _zz_4037_ = _zz_4020_[16];
  assign _zz_4038_ = _zz_4020_[17];
  assign _zz_4039_ = _zz_4020_[18];
  assign _zz_4040_ = _zz_4020_[19];
  assign _zz_4041_ = _zz_4020_[20];
  assign _zz_4042_ = _zz_4020_[21];
  assign _zz_4043_ = _zz_4020_[22];
  assign _zz_4044_ = _zz_4020_[23];
  assign _zz_4045_ = _zz_4020_[24];
  assign _zz_4046_ = _zz_4020_[25];
  assign _zz_4047_ = _zz_4020_[26];
  assign _zz_4048_ = _zz_4020_[27];
  assign _zz_4049_ = _zz_4020_[28];
  assign _zz_4050_ = _zz_4020_[29];
  assign _zz_4051_ = _zz_4020_[30];
  assign _zz_4052_ = _zz_4020_[31];
  assign _zz_4053_ = _zz_4020_[32];
  assign _zz_4054_ = _zz_4020_[33];
  assign _zz_4055_ = _zz_4020_[34];
  assign _zz_4056_ = _zz_4020_[35];
  assign _zz_4057_ = _zz_4020_[36];
  assign _zz_4058_ = _zz_4020_[37];
  assign _zz_4059_ = _zz_4020_[38];
  assign _zz_4060_ = _zz_4020_[39];
  assign _zz_4061_ = _zz_4020_[40];
  assign _zz_4062_ = _zz_4020_[41];
  assign _zz_4063_ = _zz_4020_[42];
  assign _zz_4064_ = _zz_4020_[43];
  assign _zz_4065_ = _zz_4020_[44];
  assign _zz_4066_ = _zz_4020_[45];
  assign _zz_4067_ = _zz_4020_[46];
  assign _zz_4068_ = _zz_4020_[47];
  assign _zz_4069_ = _zz_4020_[48];
  assign _zz_4070_ = _zz_4020_[49];
  assign _zz_4071_ = _zz_4020_[50];
  assign _zz_4072_ = _zz_4020_[51];
  assign _zz_4073_ = _zz_4020_[52];
  assign _zz_4074_ = _zz_4020_[53];
  assign _zz_4075_ = _zz_4020_[54];
  assign _zz_4076_ = _zz_4020_[55];
  assign _zz_4077_ = _zz_4020_[56];
  assign _zz_4078_ = _zz_4020_[57];
  assign _zz_4079_ = _zz_4020_[58];
  assign _zz_4080_ = _zz_4020_[59];
  assign _zz_4081_ = _zz_4020_[60];
  assign _zz_4082_ = _zz_4020_[61];
  assign _zz_4083_ = _zz_4020_[62];
  assign _zz_4084_ = _zz_4020_[63];
  assign _zz_4085_ = (((32'h00000300 <= load_data_area_current_addr) && (load_data_area_current_addr < 32'h00000340)) ? _zz_9__regNext : {_zz_4550_,_zz_4551_});
  assign _zz_4086_ = _zz_4085_[15 : 0];
  assign _zz_4087_ = _zz_4085_[31 : 16];
  assign _zz_4088_ = _zz_4625_[5:0];
  assign _zz_4089_ = ({63'd0,(1'b1)} <<< _zz_4088_);
  assign _zz_4090_ = _zz_4089_[0];
  assign _zz_4091_ = _zz_4089_[1];
  assign _zz_4092_ = _zz_4089_[2];
  assign _zz_4093_ = _zz_4089_[3];
  assign _zz_4094_ = _zz_4089_[4];
  assign _zz_4095_ = _zz_4089_[5];
  assign _zz_4096_ = _zz_4089_[6];
  assign _zz_4097_ = _zz_4089_[7];
  assign _zz_4098_ = _zz_4089_[8];
  assign _zz_4099_ = _zz_4089_[9];
  assign _zz_4100_ = _zz_4089_[10];
  assign _zz_4101_ = _zz_4089_[11];
  assign _zz_4102_ = _zz_4089_[12];
  assign _zz_4103_ = _zz_4089_[13];
  assign _zz_4104_ = _zz_4089_[14];
  assign _zz_4105_ = _zz_4089_[15];
  assign _zz_4106_ = _zz_4089_[16];
  assign _zz_4107_ = _zz_4089_[17];
  assign _zz_4108_ = _zz_4089_[18];
  assign _zz_4109_ = _zz_4089_[19];
  assign _zz_4110_ = _zz_4089_[20];
  assign _zz_4111_ = _zz_4089_[21];
  assign _zz_4112_ = _zz_4089_[22];
  assign _zz_4113_ = _zz_4089_[23];
  assign _zz_4114_ = _zz_4089_[24];
  assign _zz_4115_ = _zz_4089_[25];
  assign _zz_4116_ = _zz_4089_[26];
  assign _zz_4117_ = _zz_4089_[27];
  assign _zz_4118_ = _zz_4089_[28];
  assign _zz_4119_ = _zz_4089_[29];
  assign _zz_4120_ = _zz_4089_[30];
  assign _zz_4121_ = _zz_4089_[31];
  assign _zz_4122_ = _zz_4089_[32];
  assign _zz_4123_ = _zz_4089_[33];
  assign _zz_4124_ = _zz_4089_[34];
  assign _zz_4125_ = _zz_4089_[35];
  assign _zz_4126_ = _zz_4089_[36];
  assign _zz_4127_ = _zz_4089_[37];
  assign _zz_4128_ = _zz_4089_[38];
  assign _zz_4129_ = _zz_4089_[39];
  assign _zz_4130_ = _zz_4089_[40];
  assign _zz_4131_ = _zz_4089_[41];
  assign _zz_4132_ = _zz_4089_[42];
  assign _zz_4133_ = _zz_4089_[43];
  assign _zz_4134_ = _zz_4089_[44];
  assign _zz_4135_ = _zz_4089_[45];
  assign _zz_4136_ = _zz_4089_[46];
  assign _zz_4137_ = _zz_4089_[47];
  assign _zz_4138_ = _zz_4089_[48];
  assign _zz_4139_ = _zz_4089_[49];
  assign _zz_4140_ = _zz_4089_[50];
  assign _zz_4141_ = _zz_4089_[51];
  assign _zz_4142_ = _zz_4089_[52];
  assign _zz_4143_ = _zz_4089_[53];
  assign _zz_4144_ = _zz_4089_[54];
  assign _zz_4145_ = _zz_4089_[55];
  assign _zz_4146_ = _zz_4089_[56];
  assign _zz_4147_ = _zz_4089_[57];
  assign _zz_4148_ = _zz_4089_[58];
  assign _zz_4149_ = _zz_4089_[59];
  assign _zz_4150_ = _zz_4089_[60];
  assign _zz_4151_ = _zz_4089_[61];
  assign _zz_4152_ = _zz_4089_[62];
  assign _zz_4153_ = _zz_4089_[63];
  assign _zz_4154_ = (((32'h00000900 <= load_data_area_current_addr) && (load_data_area_current_addr < 32'h00000940)) ? _zz_9__regNext : {_zz_4552_,_zz_4553_});
  assign _zz_4155_ = _zz_4154_[15 : 0];
  assign _zz_4156_ = _zz_4154_[31 : 16];
  assign _zz_4157_ = _zz_4626_[5:0];
  assign _zz_4158_ = ({63'd0,(1'b1)} <<< _zz_4157_);
  assign _zz_4159_ = _zz_4158_[0];
  assign _zz_4160_ = _zz_4158_[1];
  assign _zz_4161_ = _zz_4158_[2];
  assign _zz_4162_ = _zz_4158_[3];
  assign _zz_4163_ = _zz_4158_[4];
  assign _zz_4164_ = _zz_4158_[5];
  assign _zz_4165_ = _zz_4158_[6];
  assign _zz_4166_ = _zz_4158_[7];
  assign _zz_4167_ = _zz_4158_[8];
  assign _zz_4168_ = _zz_4158_[9];
  assign _zz_4169_ = _zz_4158_[10];
  assign _zz_4170_ = _zz_4158_[11];
  assign _zz_4171_ = _zz_4158_[12];
  assign _zz_4172_ = _zz_4158_[13];
  assign _zz_4173_ = _zz_4158_[14];
  assign _zz_4174_ = _zz_4158_[15];
  assign _zz_4175_ = _zz_4158_[16];
  assign _zz_4176_ = _zz_4158_[17];
  assign _zz_4177_ = _zz_4158_[18];
  assign _zz_4178_ = _zz_4158_[19];
  assign _zz_4179_ = _zz_4158_[20];
  assign _zz_4180_ = _zz_4158_[21];
  assign _zz_4181_ = _zz_4158_[22];
  assign _zz_4182_ = _zz_4158_[23];
  assign _zz_4183_ = _zz_4158_[24];
  assign _zz_4184_ = _zz_4158_[25];
  assign _zz_4185_ = _zz_4158_[26];
  assign _zz_4186_ = _zz_4158_[27];
  assign _zz_4187_ = _zz_4158_[28];
  assign _zz_4188_ = _zz_4158_[29];
  assign _zz_4189_ = _zz_4158_[30];
  assign _zz_4190_ = _zz_4158_[31];
  assign _zz_4191_ = _zz_4158_[32];
  assign _zz_4192_ = _zz_4158_[33];
  assign _zz_4193_ = _zz_4158_[34];
  assign _zz_4194_ = _zz_4158_[35];
  assign _zz_4195_ = _zz_4158_[36];
  assign _zz_4196_ = _zz_4158_[37];
  assign _zz_4197_ = _zz_4158_[38];
  assign _zz_4198_ = _zz_4158_[39];
  assign _zz_4199_ = _zz_4158_[40];
  assign _zz_4200_ = _zz_4158_[41];
  assign _zz_4201_ = _zz_4158_[42];
  assign _zz_4202_ = _zz_4158_[43];
  assign _zz_4203_ = _zz_4158_[44];
  assign _zz_4204_ = _zz_4158_[45];
  assign _zz_4205_ = _zz_4158_[46];
  assign _zz_4206_ = _zz_4158_[47];
  assign _zz_4207_ = _zz_4158_[48];
  assign _zz_4208_ = _zz_4158_[49];
  assign _zz_4209_ = _zz_4158_[50];
  assign _zz_4210_ = _zz_4158_[51];
  assign _zz_4211_ = _zz_4158_[52];
  assign _zz_4212_ = _zz_4158_[53];
  assign _zz_4213_ = _zz_4158_[54];
  assign _zz_4214_ = _zz_4158_[55];
  assign _zz_4215_ = _zz_4158_[56];
  assign _zz_4216_ = _zz_4158_[57];
  assign _zz_4217_ = _zz_4158_[58];
  assign _zz_4218_ = _zz_4158_[59];
  assign _zz_4219_ = _zz_4158_[60];
  assign _zz_4220_ = _zz_4158_[61];
  assign _zz_4221_ = _zz_4158_[62];
  assign _zz_4222_ = _zz_4158_[63];
  assign _zz_4223_ = (((32'h00000fc0 <= load_data_area_current_addr) && (load_data_area_current_addr < 32'h00001000)) ? _zz_9__regNext : {_zz_4554_,_zz_4555_});
  assign _zz_4224_ = _zz_4223_[15 : 0];
  assign _zz_4225_ = _zz_4223_[31 : 16];
  assign _zz_4226_ = _zz_4627_[5:0];
  assign _zz_4227_ = ({63'd0,(1'b1)} <<< _zz_4226_);
  assign _zz_4228_ = _zz_4227_[0];
  assign _zz_4229_ = _zz_4227_[1];
  assign _zz_4230_ = _zz_4227_[2];
  assign _zz_4231_ = _zz_4227_[3];
  assign _zz_4232_ = _zz_4227_[4];
  assign _zz_4233_ = _zz_4227_[5];
  assign _zz_4234_ = _zz_4227_[6];
  assign _zz_4235_ = _zz_4227_[7];
  assign _zz_4236_ = _zz_4227_[8];
  assign _zz_4237_ = _zz_4227_[9];
  assign _zz_4238_ = _zz_4227_[10];
  assign _zz_4239_ = _zz_4227_[11];
  assign _zz_4240_ = _zz_4227_[12];
  assign _zz_4241_ = _zz_4227_[13];
  assign _zz_4242_ = _zz_4227_[14];
  assign _zz_4243_ = _zz_4227_[15];
  assign _zz_4244_ = _zz_4227_[16];
  assign _zz_4245_ = _zz_4227_[17];
  assign _zz_4246_ = _zz_4227_[18];
  assign _zz_4247_ = _zz_4227_[19];
  assign _zz_4248_ = _zz_4227_[20];
  assign _zz_4249_ = _zz_4227_[21];
  assign _zz_4250_ = _zz_4227_[22];
  assign _zz_4251_ = _zz_4227_[23];
  assign _zz_4252_ = _zz_4227_[24];
  assign _zz_4253_ = _zz_4227_[25];
  assign _zz_4254_ = _zz_4227_[26];
  assign _zz_4255_ = _zz_4227_[27];
  assign _zz_4256_ = _zz_4227_[28];
  assign _zz_4257_ = _zz_4227_[29];
  assign _zz_4258_ = _zz_4227_[30];
  assign _zz_4259_ = _zz_4227_[31];
  assign _zz_4260_ = _zz_4227_[32];
  assign _zz_4261_ = _zz_4227_[33];
  assign _zz_4262_ = _zz_4227_[34];
  assign _zz_4263_ = _zz_4227_[35];
  assign _zz_4264_ = _zz_4227_[36];
  assign _zz_4265_ = _zz_4227_[37];
  assign _zz_4266_ = _zz_4227_[38];
  assign _zz_4267_ = _zz_4227_[39];
  assign _zz_4268_ = _zz_4227_[40];
  assign _zz_4269_ = _zz_4227_[41];
  assign _zz_4270_ = _zz_4227_[42];
  assign _zz_4271_ = _zz_4227_[43];
  assign _zz_4272_ = _zz_4227_[44];
  assign _zz_4273_ = _zz_4227_[45];
  assign _zz_4274_ = _zz_4227_[46];
  assign _zz_4275_ = _zz_4227_[47];
  assign _zz_4276_ = _zz_4227_[48];
  assign _zz_4277_ = _zz_4227_[49];
  assign _zz_4278_ = _zz_4227_[50];
  assign _zz_4279_ = _zz_4227_[51];
  assign _zz_4280_ = _zz_4227_[52];
  assign _zz_4281_ = _zz_4227_[53];
  assign _zz_4282_ = _zz_4227_[54];
  assign _zz_4283_ = _zz_4227_[55];
  assign _zz_4284_ = _zz_4227_[56];
  assign _zz_4285_ = _zz_4227_[57];
  assign _zz_4286_ = _zz_4227_[58];
  assign _zz_4287_ = _zz_4227_[59];
  assign _zz_4288_ = _zz_4227_[60];
  assign _zz_4289_ = _zz_4227_[61];
  assign _zz_4290_ = _zz_4227_[62];
  assign _zz_4291_ = _zz_4227_[63];
  assign _zz_4292_ = (((32'h000003c0 <= load_data_area_current_addr) && (load_data_area_current_addr < 32'h00000400)) ? _zz_9__regNext : {_zz_4556_,_zz_4557_});
  assign _zz_4293_ = _zz_4292_[15 : 0];
  assign _zz_4294_ = _zz_4292_[31 : 16];
  assign _zz_4295_ = _zz_4628_[5:0];
  assign _zz_4296_ = ({63'd0,(1'b1)} <<< _zz_4295_);
  assign _zz_4297_ = _zz_4296_[0];
  assign _zz_4298_ = _zz_4296_[1];
  assign _zz_4299_ = _zz_4296_[2];
  assign _zz_4300_ = _zz_4296_[3];
  assign _zz_4301_ = _zz_4296_[4];
  assign _zz_4302_ = _zz_4296_[5];
  assign _zz_4303_ = _zz_4296_[6];
  assign _zz_4304_ = _zz_4296_[7];
  assign _zz_4305_ = _zz_4296_[8];
  assign _zz_4306_ = _zz_4296_[9];
  assign _zz_4307_ = _zz_4296_[10];
  assign _zz_4308_ = _zz_4296_[11];
  assign _zz_4309_ = _zz_4296_[12];
  assign _zz_4310_ = _zz_4296_[13];
  assign _zz_4311_ = _zz_4296_[14];
  assign _zz_4312_ = _zz_4296_[15];
  assign _zz_4313_ = _zz_4296_[16];
  assign _zz_4314_ = _zz_4296_[17];
  assign _zz_4315_ = _zz_4296_[18];
  assign _zz_4316_ = _zz_4296_[19];
  assign _zz_4317_ = _zz_4296_[20];
  assign _zz_4318_ = _zz_4296_[21];
  assign _zz_4319_ = _zz_4296_[22];
  assign _zz_4320_ = _zz_4296_[23];
  assign _zz_4321_ = _zz_4296_[24];
  assign _zz_4322_ = _zz_4296_[25];
  assign _zz_4323_ = _zz_4296_[26];
  assign _zz_4324_ = _zz_4296_[27];
  assign _zz_4325_ = _zz_4296_[28];
  assign _zz_4326_ = _zz_4296_[29];
  assign _zz_4327_ = _zz_4296_[30];
  assign _zz_4328_ = _zz_4296_[31];
  assign _zz_4329_ = _zz_4296_[32];
  assign _zz_4330_ = _zz_4296_[33];
  assign _zz_4331_ = _zz_4296_[34];
  assign _zz_4332_ = _zz_4296_[35];
  assign _zz_4333_ = _zz_4296_[36];
  assign _zz_4334_ = _zz_4296_[37];
  assign _zz_4335_ = _zz_4296_[38];
  assign _zz_4336_ = _zz_4296_[39];
  assign _zz_4337_ = _zz_4296_[40];
  assign _zz_4338_ = _zz_4296_[41];
  assign _zz_4339_ = _zz_4296_[42];
  assign _zz_4340_ = _zz_4296_[43];
  assign _zz_4341_ = _zz_4296_[44];
  assign _zz_4342_ = _zz_4296_[45];
  assign _zz_4343_ = _zz_4296_[46];
  assign _zz_4344_ = _zz_4296_[47];
  assign _zz_4345_ = _zz_4296_[48];
  assign _zz_4346_ = _zz_4296_[49];
  assign _zz_4347_ = _zz_4296_[50];
  assign _zz_4348_ = _zz_4296_[51];
  assign _zz_4349_ = _zz_4296_[52];
  assign _zz_4350_ = _zz_4296_[53];
  assign _zz_4351_ = _zz_4296_[54];
  assign _zz_4352_ = _zz_4296_[55];
  assign _zz_4353_ = _zz_4296_[56];
  assign _zz_4354_ = _zz_4296_[57];
  assign _zz_4355_ = _zz_4296_[58];
  assign _zz_4356_ = _zz_4296_[59];
  assign _zz_4357_ = _zz_4296_[60];
  assign _zz_4358_ = _zz_4296_[61];
  assign _zz_4359_ = _zz_4296_[62];
  assign _zz_4360_ = _zz_4296_[63];
  assign _zz_4361_ = (((32'h00000bc0 <= load_data_area_current_addr) && (load_data_area_current_addr < 32'h00000c00)) ? _zz_9__regNext : {_zz_4558_,_zz_4559_});
  assign _zz_4362_ = _zz_4361_[15 : 0];
  assign _zz_4363_ = _zz_4361_[31 : 16];
  assign _zz_4364_ = _zz_4629_[5:0];
  assign _zz_4365_ = ({63'd0,(1'b1)} <<< _zz_4364_);
  assign _zz_4366_ = _zz_4365_[0];
  assign _zz_4367_ = _zz_4365_[1];
  assign _zz_4368_ = _zz_4365_[2];
  assign _zz_4369_ = _zz_4365_[3];
  assign _zz_4370_ = _zz_4365_[4];
  assign _zz_4371_ = _zz_4365_[5];
  assign _zz_4372_ = _zz_4365_[6];
  assign _zz_4373_ = _zz_4365_[7];
  assign _zz_4374_ = _zz_4365_[8];
  assign _zz_4375_ = _zz_4365_[9];
  assign _zz_4376_ = _zz_4365_[10];
  assign _zz_4377_ = _zz_4365_[11];
  assign _zz_4378_ = _zz_4365_[12];
  assign _zz_4379_ = _zz_4365_[13];
  assign _zz_4380_ = _zz_4365_[14];
  assign _zz_4381_ = _zz_4365_[15];
  assign _zz_4382_ = _zz_4365_[16];
  assign _zz_4383_ = _zz_4365_[17];
  assign _zz_4384_ = _zz_4365_[18];
  assign _zz_4385_ = _zz_4365_[19];
  assign _zz_4386_ = _zz_4365_[20];
  assign _zz_4387_ = _zz_4365_[21];
  assign _zz_4388_ = _zz_4365_[22];
  assign _zz_4389_ = _zz_4365_[23];
  assign _zz_4390_ = _zz_4365_[24];
  assign _zz_4391_ = _zz_4365_[25];
  assign _zz_4392_ = _zz_4365_[26];
  assign _zz_4393_ = _zz_4365_[27];
  assign _zz_4394_ = _zz_4365_[28];
  assign _zz_4395_ = _zz_4365_[29];
  assign _zz_4396_ = _zz_4365_[30];
  assign _zz_4397_ = _zz_4365_[31];
  assign _zz_4398_ = _zz_4365_[32];
  assign _zz_4399_ = _zz_4365_[33];
  assign _zz_4400_ = _zz_4365_[34];
  assign _zz_4401_ = _zz_4365_[35];
  assign _zz_4402_ = _zz_4365_[36];
  assign _zz_4403_ = _zz_4365_[37];
  assign _zz_4404_ = _zz_4365_[38];
  assign _zz_4405_ = _zz_4365_[39];
  assign _zz_4406_ = _zz_4365_[40];
  assign _zz_4407_ = _zz_4365_[41];
  assign _zz_4408_ = _zz_4365_[42];
  assign _zz_4409_ = _zz_4365_[43];
  assign _zz_4410_ = _zz_4365_[44];
  assign _zz_4411_ = _zz_4365_[45];
  assign _zz_4412_ = _zz_4365_[46];
  assign _zz_4413_ = _zz_4365_[47];
  assign _zz_4414_ = _zz_4365_[48];
  assign _zz_4415_ = _zz_4365_[49];
  assign _zz_4416_ = _zz_4365_[50];
  assign _zz_4417_ = _zz_4365_[51];
  assign _zz_4418_ = _zz_4365_[52];
  assign _zz_4419_ = _zz_4365_[53];
  assign _zz_4420_ = _zz_4365_[54];
  assign _zz_4421_ = _zz_4365_[55];
  assign _zz_4422_ = _zz_4365_[56];
  assign _zz_4423_ = _zz_4365_[57];
  assign _zz_4424_ = _zz_4365_[58];
  assign _zz_4425_ = _zz_4365_[59];
  assign _zz_4426_ = _zz_4365_[60];
  assign _zz_4427_ = _zz_4365_[61];
  assign _zz_4428_ = _zz_4365_[62];
  assign _zz_4429_ = _zz_4365_[63];
  assign _zz_4430_ = (((32'h00000480 <= load_data_area_current_addr) && (load_data_area_current_addr < 32'h000004c0)) ? _zz_9__regNext : {_zz_4560_,_zz_4561_});
  assign _zz_4431_ = _zz_4430_[15 : 0];
  assign _zz_4432_ = _zz_4430_[31 : 16];
  assign io_coef_out_valid = transfer_done;
  assign io_coef_out_payload_0_0_0_real = int_reg_array_0_0_real;
  assign io_coef_out_payload_0_0_0_imag = int_reg_array_0_0_imag;
  assign io_coef_out_payload_0_0_1_real = int_reg_array_0_1_real;
  assign io_coef_out_payload_0_0_1_imag = int_reg_array_0_1_imag;
  assign io_coef_out_payload_0_0_2_real = int_reg_array_0_2_real;
  assign io_coef_out_payload_0_0_2_imag = int_reg_array_0_2_imag;
  assign io_coef_out_payload_0_0_3_real = int_reg_array_0_3_real;
  assign io_coef_out_payload_0_0_3_imag = int_reg_array_0_3_imag;
  assign io_coef_out_payload_0_0_4_real = int_reg_array_0_4_real;
  assign io_coef_out_payload_0_0_4_imag = int_reg_array_0_4_imag;
  assign io_coef_out_payload_0_0_5_real = int_reg_array_0_5_real;
  assign io_coef_out_payload_0_0_5_imag = int_reg_array_0_5_imag;
  assign io_coef_out_payload_0_0_6_real = int_reg_array_0_6_real;
  assign io_coef_out_payload_0_0_6_imag = int_reg_array_0_6_imag;
  assign io_coef_out_payload_0_0_7_real = int_reg_array_0_7_real;
  assign io_coef_out_payload_0_0_7_imag = int_reg_array_0_7_imag;
  assign io_coef_out_payload_0_0_8_real = int_reg_array_0_8_real;
  assign io_coef_out_payload_0_0_8_imag = int_reg_array_0_8_imag;
  assign io_coef_out_payload_0_0_9_real = int_reg_array_0_9_real;
  assign io_coef_out_payload_0_0_9_imag = int_reg_array_0_9_imag;
  assign io_coef_out_payload_0_0_10_real = int_reg_array_0_10_real;
  assign io_coef_out_payload_0_0_10_imag = int_reg_array_0_10_imag;
  assign io_coef_out_payload_0_0_11_real = int_reg_array_0_11_real;
  assign io_coef_out_payload_0_0_11_imag = int_reg_array_0_11_imag;
  assign io_coef_out_payload_0_0_12_real = int_reg_array_0_12_real;
  assign io_coef_out_payload_0_0_12_imag = int_reg_array_0_12_imag;
  assign io_coef_out_payload_0_0_13_real = int_reg_array_0_13_real;
  assign io_coef_out_payload_0_0_13_imag = int_reg_array_0_13_imag;
  assign io_coef_out_payload_0_0_14_real = int_reg_array_0_14_real;
  assign io_coef_out_payload_0_0_14_imag = int_reg_array_0_14_imag;
  assign io_coef_out_payload_0_0_15_real = int_reg_array_0_15_real;
  assign io_coef_out_payload_0_0_15_imag = int_reg_array_0_15_imag;
  assign io_coef_out_payload_0_0_16_real = int_reg_array_0_16_real;
  assign io_coef_out_payload_0_0_16_imag = int_reg_array_0_16_imag;
  assign io_coef_out_payload_0_0_17_real = int_reg_array_0_17_real;
  assign io_coef_out_payload_0_0_17_imag = int_reg_array_0_17_imag;
  assign io_coef_out_payload_0_0_18_real = int_reg_array_0_18_real;
  assign io_coef_out_payload_0_0_18_imag = int_reg_array_0_18_imag;
  assign io_coef_out_payload_0_0_19_real = int_reg_array_0_19_real;
  assign io_coef_out_payload_0_0_19_imag = int_reg_array_0_19_imag;
  assign io_coef_out_payload_0_0_20_real = int_reg_array_0_20_real;
  assign io_coef_out_payload_0_0_20_imag = int_reg_array_0_20_imag;
  assign io_coef_out_payload_0_0_21_real = int_reg_array_0_21_real;
  assign io_coef_out_payload_0_0_21_imag = int_reg_array_0_21_imag;
  assign io_coef_out_payload_0_0_22_real = int_reg_array_0_22_real;
  assign io_coef_out_payload_0_0_22_imag = int_reg_array_0_22_imag;
  assign io_coef_out_payload_0_0_23_real = int_reg_array_0_23_real;
  assign io_coef_out_payload_0_0_23_imag = int_reg_array_0_23_imag;
  assign io_coef_out_payload_0_0_24_real = int_reg_array_0_24_real;
  assign io_coef_out_payload_0_0_24_imag = int_reg_array_0_24_imag;
  assign io_coef_out_payload_0_0_25_real = int_reg_array_0_25_real;
  assign io_coef_out_payload_0_0_25_imag = int_reg_array_0_25_imag;
  assign io_coef_out_payload_0_0_26_real = int_reg_array_0_26_real;
  assign io_coef_out_payload_0_0_26_imag = int_reg_array_0_26_imag;
  assign io_coef_out_payload_0_0_27_real = int_reg_array_0_27_real;
  assign io_coef_out_payload_0_0_27_imag = int_reg_array_0_27_imag;
  assign io_coef_out_payload_0_0_28_real = int_reg_array_0_28_real;
  assign io_coef_out_payload_0_0_28_imag = int_reg_array_0_28_imag;
  assign io_coef_out_payload_0_0_29_real = int_reg_array_0_29_real;
  assign io_coef_out_payload_0_0_29_imag = int_reg_array_0_29_imag;
  assign io_coef_out_payload_0_0_30_real = int_reg_array_0_30_real;
  assign io_coef_out_payload_0_0_30_imag = int_reg_array_0_30_imag;
  assign io_coef_out_payload_0_0_31_real = int_reg_array_0_31_real;
  assign io_coef_out_payload_0_0_31_imag = int_reg_array_0_31_imag;
  assign io_coef_out_payload_0_0_32_real = int_reg_array_0_32_real;
  assign io_coef_out_payload_0_0_32_imag = int_reg_array_0_32_imag;
  assign io_coef_out_payload_0_0_33_real = int_reg_array_0_33_real;
  assign io_coef_out_payload_0_0_33_imag = int_reg_array_0_33_imag;
  assign io_coef_out_payload_0_0_34_real = int_reg_array_0_34_real;
  assign io_coef_out_payload_0_0_34_imag = int_reg_array_0_34_imag;
  assign io_coef_out_payload_0_0_35_real = int_reg_array_0_35_real;
  assign io_coef_out_payload_0_0_35_imag = int_reg_array_0_35_imag;
  assign io_coef_out_payload_0_0_36_real = int_reg_array_0_36_real;
  assign io_coef_out_payload_0_0_36_imag = int_reg_array_0_36_imag;
  assign io_coef_out_payload_0_0_37_real = int_reg_array_0_37_real;
  assign io_coef_out_payload_0_0_37_imag = int_reg_array_0_37_imag;
  assign io_coef_out_payload_0_0_38_real = int_reg_array_0_38_real;
  assign io_coef_out_payload_0_0_38_imag = int_reg_array_0_38_imag;
  assign io_coef_out_payload_0_0_39_real = int_reg_array_0_39_real;
  assign io_coef_out_payload_0_0_39_imag = int_reg_array_0_39_imag;
  assign io_coef_out_payload_0_0_40_real = int_reg_array_0_40_real;
  assign io_coef_out_payload_0_0_40_imag = int_reg_array_0_40_imag;
  assign io_coef_out_payload_0_0_41_real = int_reg_array_0_41_real;
  assign io_coef_out_payload_0_0_41_imag = int_reg_array_0_41_imag;
  assign io_coef_out_payload_0_0_42_real = int_reg_array_0_42_real;
  assign io_coef_out_payload_0_0_42_imag = int_reg_array_0_42_imag;
  assign io_coef_out_payload_0_0_43_real = int_reg_array_0_43_real;
  assign io_coef_out_payload_0_0_43_imag = int_reg_array_0_43_imag;
  assign io_coef_out_payload_0_0_44_real = int_reg_array_0_44_real;
  assign io_coef_out_payload_0_0_44_imag = int_reg_array_0_44_imag;
  assign io_coef_out_payload_0_0_45_real = int_reg_array_0_45_real;
  assign io_coef_out_payload_0_0_45_imag = int_reg_array_0_45_imag;
  assign io_coef_out_payload_0_0_46_real = int_reg_array_0_46_real;
  assign io_coef_out_payload_0_0_46_imag = int_reg_array_0_46_imag;
  assign io_coef_out_payload_0_0_47_real = int_reg_array_0_47_real;
  assign io_coef_out_payload_0_0_47_imag = int_reg_array_0_47_imag;
  assign io_coef_out_payload_0_0_48_real = int_reg_array_0_48_real;
  assign io_coef_out_payload_0_0_48_imag = int_reg_array_0_48_imag;
  assign io_coef_out_payload_0_0_49_real = int_reg_array_0_49_real;
  assign io_coef_out_payload_0_0_49_imag = int_reg_array_0_49_imag;
  assign io_coef_out_payload_0_1_0_real = int_reg_array_1_0_real;
  assign io_coef_out_payload_0_1_0_imag = int_reg_array_1_0_imag;
  assign io_coef_out_payload_0_1_1_real = int_reg_array_1_1_real;
  assign io_coef_out_payload_0_1_1_imag = int_reg_array_1_1_imag;
  assign io_coef_out_payload_0_1_2_real = int_reg_array_1_2_real;
  assign io_coef_out_payload_0_1_2_imag = int_reg_array_1_2_imag;
  assign io_coef_out_payload_0_1_3_real = int_reg_array_1_3_real;
  assign io_coef_out_payload_0_1_3_imag = int_reg_array_1_3_imag;
  assign io_coef_out_payload_0_1_4_real = int_reg_array_1_4_real;
  assign io_coef_out_payload_0_1_4_imag = int_reg_array_1_4_imag;
  assign io_coef_out_payload_0_1_5_real = int_reg_array_1_5_real;
  assign io_coef_out_payload_0_1_5_imag = int_reg_array_1_5_imag;
  assign io_coef_out_payload_0_1_6_real = int_reg_array_1_6_real;
  assign io_coef_out_payload_0_1_6_imag = int_reg_array_1_6_imag;
  assign io_coef_out_payload_0_1_7_real = int_reg_array_1_7_real;
  assign io_coef_out_payload_0_1_7_imag = int_reg_array_1_7_imag;
  assign io_coef_out_payload_0_1_8_real = int_reg_array_1_8_real;
  assign io_coef_out_payload_0_1_8_imag = int_reg_array_1_8_imag;
  assign io_coef_out_payload_0_1_9_real = int_reg_array_1_9_real;
  assign io_coef_out_payload_0_1_9_imag = int_reg_array_1_9_imag;
  assign io_coef_out_payload_0_1_10_real = int_reg_array_1_10_real;
  assign io_coef_out_payload_0_1_10_imag = int_reg_array_1_10_imag;
  assign io_coef_out_payload_0_1_11_real = int_reg_array_1_11_real;
  assign io_coef_out_payload_0_1_11_imag = int_reg_array_1_11_imag;
  assign io_coef_out_payload_0_1_12_real = int_reg_array_1_12_real;
  assign io_coef_out_payload_0_1_12_imag = int_reg_array_1_12_imag;
  assign io_coef_out_payload_0_1_13_real = int_reg_array_1_13_real;
  assign io_coef_out_payload_0_1_13_imag = int_reg_array_1_13_imag;
  assign io_coef_out_payload_0_1_14_real = int_reg_array_1_14_real;
  assign io_coef_out_payload_0_1_14_imag = int_reg_array_1_14_imag;
  assign io_coef_out_payload_0_1_15_real = int_reg_array_1_15_real;
  assign io_coef_out_payload_0_1_15_imag = int_reg_array_1_15_imag;
  assign io_coef_out_payload_0_1_16_real = int_reg_array_1_16_real;
  assign io_coef_out_payload_0_1_16_imag = int_reg_array_1_16_imag;
  assign io_coef_out_payload_0_1_17_real = int_reg_array_1_17_real;
  assign io_coef_out_payload_0_1_17_imag = int_reg_array_1_17_imag;
  assign io_coef_out_payload_0_1_18_real = int_reg_array_1_18_real;
  assign io_coef_out_payload_0_1_18_imag = int_reg_array_1_18_imag;
  assign io_coef_out_payload_0_1_19_real = int_reg_array_1_19_real;
  assign io_coef_out_payload_0_1_19_imag = int_reg_array_1_19_imag;
  assign io_coef_out_payload_0_1_20_real = int_reg_array_1_20_real;
  assign io_coef_out_payload_0_1_20_imag = int_reg_array_1_20_imag;
  assign io_coef_out_payload_0_1_21_real = int_reg_array_1_21_real;
  assign io_coef_out_payload_0_1_21_imag = int_reg_array_1_21_imag;
  assign io_coef_out_payload_0_1_22_real = int_reg_array_1_22_real;
  assign io_coef_out_payload_0_1_22_imag = int_reg_array_1_22_imag;
  assign io_coef_out_payload_0_1_23_real = int_reg_array_1_23_real;
  assign io_coef_out_payload_0_1_23_imag = int_reg_array_1_23_imag;
  assign io_coef_out_payload_0_1_24_real = int_reg_array_1_24_real;
  assign io_coef_out_payload_0_1_24_imag = int_reg_array_1_24_imag;
  assign io_coef_out_payload_0_1_25_real = int_reg_array_1_25_real;
  assign io_coef_out_payload_0_1_25_imag = int_reg_array_1_25_imag;
  assign io_coef_out_payload_0_1_26_real = int_reg_array_1_26_real;
  assign io_coef_out_payload_0_1_26_imag = int_reg_array_1_26_imag;
  assign io_coef_out_payload_0_1_27_real = int_reg_array_1_27_real;
  assign io_coef_out_payload_0_1_27_imag = int_reg_array_1_27_imag;
  assign io_coef_out_payload_0_1_28_real = int_reg_array_1_28_real;
  assign io_coef_out_payload_0_1_28_imag = int_reg_array_1_28_imag;
  assign io_coef_out_payload_0_1_29_real = int_reg_array_1_29_real;
  assign io_coef_out_payload_0_1_29_imag = int_reg_array_1_29_imag;
  assign io_coef_out_payload_0_1_30_real = int_reg_array_1_30_real;
  assign io_coef_out_payload_0_1_30_imag = int_reg_array_1_30_imag;
  assign io_coef_out_payload_0_1_31_real = int_reg_array_1_31_real;
  assign io_coef_out_payload_0_1_31_imag = int_reg_array_1_31_imag;
  assign io_coef_out_payload_0_1_32_real = int_reg_array_1_32_real;
  assign io_coef_out_payload_0_1_32_imag = int_reg_array_1_32_imag;
  assign io_coef_out_payload_0_1_33_real = int_reg_array_1_33_real;
  assign io_coef_out_payload_0_1_33_imag = int_reg_array_1_33_imag;
  assign io_coef_out_payload_0_1_34_real = int_reg_array_1_34_real;
  assign io_coef_out_payload_0_1_34_imag = int_reg_array_1_34_imag;
  assign io_coef_out_payload_0_1_35_real = int_reg_array_1_35_real;
  assign io_coef_out_payload_0_1_35_imag = int_reg_array_1_35_imag;
  assign io_coef_out_payload_0_1_36_real = int_reg_array_1_36_real;
  assign io_coef_out_payload_0_1_36_imag = int_reg_array_1_36_imag;
  assign io_coef_out_payload_0_1_37_real = int_reg_array_1_37_real;
  assign io_coef_out_payload_0_1_37_imag = int_reg_array_1_37_imag;
  assign io_coef_out_payload_0_1_38_real = int_reg_array_1_38_real;
  assign io_coef_out_payload_0_1_38_imag = int_reg_array_1_38_imag;
  assign io_coef_out_payload_0_1_39_real = int_reg_array_1_39_real;
  assign io_coef_out_payload_0_1_39_imag = int_reg_array_1_39_imag;
  assign io_coef_out_payload_0_1_40_real = int_reg_array_1_40_real;
  assign io_coef_out_payload_0_1_40_imag = int_reg_array_1_40_imag;
  assign io_coef_out_payload_0_1_41_real = int_reg_array_1_41_real;
  assign io_coef_out_payload_0_1_41_imag = int_reg_array_1_41_imag;
  assign io_coef_out_payload_0_1_42_real = int_reg_array_1_42_real;
  assign io_coef_out_payload_0_1_42_imag = int_reg_array_1_42_imag;
  assign io_coef_out_payload_0_1_43_real = int_reg_array_1_43_real;
  assign io_coef_out_payload_0_1_43_imag = int_reg_array_1_43_imag;
  assign io_coef_out_payload_0_1_44_real = int_reg_array_1_44_real;
  assign io_coef_out_payload_0_1_44_imag = int_reg_array_1_44_imag;
  assign io_coef_out_payload_0_1_45_real = int_reg_array_1_45_real;
  assign io_coef_out_payload_0_1_45_imag = int_reg_array_1_45_imag;
  assign io_coef_out_payload_0_1_46_real = int_reg_array_1_46_real;
  assign io_coef_out_payload_0_1_46_imag = int_reg_array_1_46_imag;
  assign io_coef_out_payload_0_1_47_real = int_reg_array_1_47_real;
  assign io_coef_out_payload_0_1_47_imag = int_reg_array_1_47_imag;
  assign io_coef_out_payload_0_1_48_real = int_reg_array_1_48_real;
  assign io_coef_out_payload_0_1_48_imag = int_reg_array_1_48_imag;
  assign io_coef_out_payload_0_1_49_real = int_reg_array_1_49_real;
  assign io_coef_out_payload_0_1_49_imag = int_reg_array_1_49_imag;
  assign io_coef_out_payload_0_2_0_real = int_reg_array_2_0_real;
  assign io_coef_out_payload_0_2_0_imag = int_reg_array_2_0_imag;
  assign io_coef_out_payload_0_2_1_real = int_reg_array_2_1_real;
  assign io_coef_out_payload_0_2_1_imag = int_reg_array_2_1_imag;
  assign io_coef_out_payload_0_2_2_real = int_reg_array_2_2_real;
  assign io_coef_out_payload_0_2_2_imag = int_reg_array_2_2_imag;
  assign io_coef_out_payload_0_2_3_real = int_reg_array_2_3_real;
  assign io_coef_out_payload_0_2_3_imag = int_reg_array_2_3_imag;
  assign io_coef_out_payload_0_2_4_real = int_reg_array_2_4_real;
  assign io_coef_out_payload_0_2_4_imag = int_reg_array_2_4_imag;
  assign io_coef_out_payload_0_2_5_real = int_reg_array_2_5_real;
  assign io_coef_out_payload_0_2_5_imag = int_reg_array_2_5_imag;
  assign io_coef_out_payload_0_2_6_real = int_reg_array_2_6_real;
  assign io_coef_out_payload_0_2_6_imag = int_reg_array_2_6_imag;
  assign io_coef_out_payload_0_2_7_real = int_reg_array_2_7_real;
  assign io_coef_out_payload_0_2_7_imag = int_reg_array_2_7_imag;
  assign io_coef_out_payload_0_2_8_real = int_reg_array_2_8_real;
  assign io_coef_out_payload_0_2_8_imag = int_reg_array_2_8_imag;
  assign io_coef_out_payload_0_2_9_real = int_reg_array_2_9_real;
  assign io_coef_out_payload_0_2_9_imag = int_reg_array_2_9_imag;
  assign io_coef_out_payload_0_2_10_real = int_reg_array_2_10_real;
  assign io_coef_out_payload_0_2_10_imag = int_reg_array_2_10_imag;
  assign io_coef_out_payload_0_2_11_real = int_reg_array_2_11_real;
  assign io_coef_out_payload_0_2_11_imag = int_reg_array_2_11_imag;
  assign io_coef_out_payload_0_2_12_real = int_reg_array_2_12_real;
  assign io_coef_out_payload_0_2_12_imag = int_reg_array_2_12_imag;
  assign io_coef_out_payload_0_2_13_real = int_reg_array_2_13_real;
  assign io_coef_out_payload_0_2_13_imag = int_reg_array_2_13_imag;
  assign io_coef_out_payload_0_2_14_real = int_reg_array_2_14_real;
  assign io_coef_out_payload_0_2_14_imag = int_reg_array_2_14_imag;
  assign io_coef_out_payload_0_2_15_real = int_reg_array_2_15_real;
  assign io_coef_out_payload_0_2_15_imag = int_reg_array_2_15_imag;
  assign io_coef_out_payload_0_2_16_real = int_reg_array_2_16_real;
  assign io_coef_out_payload_0_2_16_imag = int_reg_array_2_16_imag;
  assign io_coef_out_payload_0_2_17_real = int_reg_array_2_17_real;
  assign io_coef_out_payload_0_2_17_imag = int_reg_array_2_17_imag;
  assign io_coef_out_payload_0_2_18_real = int_reg_array_2_18_real;
  assign io_coef_out_payload_0_2_18_imag = int_reg_array_2_18_imag;
  assign io_coef_out_payload_0_2_19_real = int_reg_array_2_19_real;
  assign io_coef_out_payload_0_2_19_imag = int_reg_array_2_19_imag;
  assign io_coef_out_payload_0_2_20_real = int_reg_array_2_20_real;
  assign io_coef_out_payload_0_2_20_imag = int_reg_array_2_20_imag;
  assign io_coef_out_payload_0_2_21_real = int_reg_array_2_21_real;
  assign io_coef_out_payload_0_2_21_imag = int_reg_array_2_21_imag;
  assign io_coef_out_payload_0_2_22_real = int_reg_array_2_22_real;
  assign io_coef_out_payload_0_2_22_imag = int_reg_array_2_22_imag;
  assign io_coef_out_payload_0_2_23_real = int_reg_array_2_23_real;
  assign io_coef_out_payload_0_2_23_imag = int_reg_array_2_23_imag;
  assign io_coef_out_payload_0_2_24_real = int_reg_array_2_24_real;
  assign io_coef_out_payload_0_2_24_imag = int_reg_array_2_24_imag;
  assign io_coef_out_payload_0_2_25_real = int_reg_array_2_25_real;
  assign io_coef_out_payload_0_2_25_imag = int_reg_array_2_25_imag;
  assign io_coef_out_payload_0_2_26_real = int_reg_array_2_26_real;
  assign io_coef_out_payload_0_2_26_imag = int_reg_array_2_26_imag;
  assign io_coef_out_payload_0_2_27_real = int_reg_array_2_27_real;
  assign io_coef_out_payload_0_2_27_imag = int_reg_array_2_27_imag;
  assign io_coef_out_payload_0_2_28_real = int_reg_array_2_28_real;
  assign io_coef_out_payload_0_2_28_imag = int_reg_array_2_28_imag;
  assign io_coef_out_payload_0_2_29_real = int_reg_array_2_29_real;
  assign io_coef_out_payload_0_2_29_imag = int_reg_array_2_29_imag;
  assign io_coef_out_payload_0_2_30_real = int_reg_array_2_30_real;
  assign io_coef_out_payload_0_2_30_imag = int_reg_array_2_30_imag;
  assign io_coef_out_payload_0_2_31_real = int_reg_array_2_31_real;
  assign io_coef_out_payload_0_2_31_imag = int_reg_array_2_31_imag;
  assign io_coef_out_payload_0_2_32_real = int_reg_array_2_32_real;
  assign io_coef_out_payload_0_2_32_imag = int_reg_array_2_32_imag;
  assign io_coef_out_payload_0_2_33_real = int_reg_array_2_33_real;
  assign io_coef_out_payload_0_2_33_imag = int_reg_array_2_33_imag;
  assign io_coef_out_payload_0_2_34_real = int_reg_array_2_34_real;
  assign io_coef_out_payload_0_2_34_imag = int_reg_array_2_34_imag;
  assign io_coef_out_payload_0_2_35_real = int_reg_array_2_35_real;
  assign io_coef_out_payload_0_2_35_imag = int_reg_array_2_35_imag;
  assign io_coef_out_payload_0_2_36_real = int_reg_array_2_36_real;
  assign io_coef_out_payload_0_2_36_imag = int_reg_array_2_36_imag;
  assign io_coef_out_payload_0_2_37_real = int_reg_array_2_37_real;
  assign io_coef_out_payload_0_2_37_imag = int_reg_array_2_37_imag;
  assign io_coef_out_payload_0_2_38_real = int_reg_array_2_38_real;
  assign io_coef_out_payload_0_2_38_imag = int_reg_array_2_38_imag;
  assign io_coef_out_payload_0_2_39_real = int_reg_array_2_39_real;
  assign io_coef_out_payload_0_2_39_imag = int_reg_array_2_39_imag;
  assign io_coef_out_payload_0_2_40_real = int_reg_array_2_40_real;
  assign io_coef_out_payload_0_2_40_imag = int_reg_array_2_40_imag;
  assign io_coef_out_payload_0_2_41_real = int_reg_array_2_41_real;
  assign io_coef_out_payload_0_2_41_imag = int_reg_array_2_41_imag;
  assign io_coef_out_payload_0_2_42_real = int_reg_array_2_42_real;
  assign io_coef_out_payload_0_2_42_imag = int_reg_array_2_42_imag;
  assign io_coef_out_payload_0_2_43_real = int_reg_array_2_43_real;
  assign io_coef_out_payload_0_2_43_imag = int_reg_array_2_43_imag;
  assign io_coef_out_payload_0_2_44_real = int_reg_array_2_44_real;
  assign io_coef_out_payload_0_2_44_imag = int_reg_array_2_44_imag;
  assign io_coef_out_payload_0_2_45_real = int_reg_array_2_45_real;
  assign io_coef_out_payload_0_2_45_imag = int_reg_array_2_45_imag;
  assign io_coef_out_payload_0_2_46_real = int_reg_array_2_46_real;
  assign io_coef_out_payload_0_2_46_imag = int_reg_array_2_46_imag;
  assign io_coef_out_payload_0_2_47_real = int_reg_array_2_47_real;
  assign io_coef_out_payload_0_2_47_imag = int_reg_array_2_47_imag;
  assign io_coef_out_payload_0_2_48_real = int_reg_array_2_48_real;
  assign io_coef_out_payload_0_2_48_imag = int_reg_array_2_48_imag;
  assign io_coef_out_payload_0_2_49_real = int_reg_array_2_49_real;
  assign io_coef_out_payload_0_2_49_imag = int_reg_array_2_49_imag;
  assign io_coef_out_payload_0_3_0_real = int_reg_array_3_0_real;
  assign io_coef_out_payload_0_3_0_imag = int_reg_array_3_0_imag;
  assign io_coef_out_payload_0_3_1_real = int_reg_array_3_1_real;
  assign io_coef_out_payload_0_3_1_imag = int_reg_array_3_1_imag;
  assign io_coef_out_payload_0_3_2_real = int_reg_array_3_2_real;
  assign io_coef_out_payload_0_3_2_imag = int_reg_array_3_2_imag;
  assign io_coef_out_payload_0_3_3_real = int_reg_array_3_3_real;
  assign io_coef_out_payload_0_3_3_imag = int_reg_array_3_3_imag;
  assign io_coef_out_payload_0_3_4_real = int_reg_array_3_4_real;
  assign io_coef_out_payload_0_3_4_imag = int_reg_array_3_4_imag;
  assign io_coef_out_payload_0_3_5_real = int_reg_array_3_5_real;
  assign io_coef_out_payload_0_3_5_imag = int_reg_array_3_5_imag;
  assign io_coef_out_payload_0_3_6_real = int_reg_array_3_6_real;
  assign io_coef_out_payload_0_3_6_imag = int_reg_array_3_6_imag;
  assign io_coef_out_payload_0_3_7_real = int_reg_array_3_7_real;
  assign io_coef_out_payload_0_3_7_imag = int_reg_array_3_7_imag;
  assign io_coef_out_payload_0_3_8_real = int_reg_array_3_8_real;
  assign io_coef_out_payload_0_3_8_imag = int_reg_array_3_8_imag;
  assign io_coef_out_payload_0_3_9_real = int_reg_array_3_9_real;
  assign io_coef_out_payload_0_3_9_imag = int_reg_array_3_9_imag;
  assign io_coef_out_payload_0_3_10_real = int_reg_array_3_10_real;
  assign io_coef_out_payload_0_3_10_imag = int_reg_array_3_10_imag;
  assign io_coef_out_payload_0_3_11_real = int_reg_array_3_11_real;
  assign io_coef_out_payload_0_3_11_imag = int_reg_array_3_11_imag;
  assign io_coef_out_payload_0_3_12_real = int_reg_array_3_12_real;
  assign io_coef_out_payload_0_3_12_imag = int_reg_array_3_12_imag;
  assign io_coef_out_payload_0_3_13_real = int_reg_array_3_13_real;
  assign io_coef_out_payload_0_3_13_imag = int_reg_array_3_13_imag;
  assign io_coef_out_payload_0_3_14_real = int_reg_array_3_14_real;
  assign io_coef_out_payload_0_3_14_imag = int_reg_array_3_14_imag;
  assign io_coef_out_payload_0_3_15_real = int_reg_array_3_15_real;
  assign io_coef_out_payload_0_3_15_imag = int_reg_array_3_15_imag;
  assign io_coef_out_payload_0_3_16_real = int_reg_array_3_16_real;
  assign io_coef_out_payload_0_3_16_imag = int_reg_array_3_16_imag;
  assign io_coef_out_payload_0_3_17_real = int_reg_array_3_17_real;
  assign io_coef_out_payload_0_3_17_imag = int_reg_array_3_17_imag;
  assign io_coef_out_payload_0_3_18_real = int_reg_array_3_18_real;
  assign io_coef_out_payload_0_3_18_imag = int_reg_array_3_18_imag;
  assign io_coef_out_payload_0_3_19_real = int_reg_array_3_19_real;
  assign io_coef_out_payload_0_3_19_imag = int_reg_array_3_19_imag;
  assign io_coef_out_payload_0_3_20_real = int_reg_array_3_20_real;
  assign io_coef_out_payload_0_3_20_imag = int_reg_array_3_20_imag;
  assign io_coef_out_payload_0_3_21_real = int_reg_array_3_21_real;
  assign io_coef_out_payload_0_3_21_imag = int_reg_array_3_21_imag;
  assign io_coef_out_payload_0_3_22_real = int_reg_array_3_22_real;
  assign io_coef_out_payload_0_3_22_imag = int_reg_array_3_22_imag;
  assign io_coef_out_payload_0_3_23_real = int_reg_array_3_23_real;
  assign io_coef_out_payload_0_3_23_imag = int_reg_array_3_23_imag;
  assign io_coef_out_payload_0_3_24_real = int_reg_array_3_24_real;
  assign io_coef_out_payload_0_3_24_imag = int_reg_array_3_24_imag;
  assign io_coef_out_payload_0_3_25_real = int_reg_array_3_25_real;
  assign io_coef_out_payload_0_3_25_imag = int_reg_array_3_25_imag;
  assign io_coef_out_payload_0_3_26_real = int_reg_array_3_26_real;
  assign io_coef_out_payload_0_3_26_imag = int_reg_array_3_26_imag;
  assign io_coef_out_payload_0_3_27_real = int_reg_array_3_27_real;
  assign io_coef_out_payload_0_3_27_imag = int_reg_array_3_27_imag;
  assign io_coef_out_payload_0_3_28_real = int_reg_array_3_28_real;
  assign io_coef_out_payload_0_3_28_imag = int_reg_array_3_28_imag;
  assign io_coef_out_payload_0_3_29_real = int_reg_array_3_29_real;
  assign io_coef_out_payload_0_3_29_imag = int_reg_array_3_29_imag;
  assign io_coef_out_payload_0_3_30_real = int_reg_array_3_30_real;
  assign io_coef_out_payload_0_3_30_imag = int_reg_array_3_30_imag;
  assign io_coef_out_payload_0_3_31_real = int_reg_array_3_31_real;
  assign io_coef_out_payload_0_3_31_imag = int_reg_array_3_31_imag;
  assign io_coef_out_payload_0_3_32_real = int_reg_array_3_32_real;
  assign io_coef_out_payload_0_3_32_imag = int_reg_array_3_32_imag;
  assign io_coef_out_payload_0_3_33_real = int_reg_array_3_33_real;
  assign io_coef_out_payload_0_3_33_imag = int_reg_array_3_33_imag;
  assign io_coef_out_payload_0_3_34_real = int_reg_array_3_34_real;
  assign io_coef_out_payload_0_3_34_imag = int_reg_array_3_34_imag;
  assign io_coef_out_payload_0_3_35_real = int_reg_array_3_35_real;
  assign io_coef_out_payload_0_3_35_imag = int_reg_array_3_35_imag;
  assign io_coef_out_payload_0_3_36_real = int_reg_array_3_36_real;
  assign io_coef_out_payload_0_3_36_imag = int_reg_array_3_36_imag;
  assign io_coef_out_payload_0_3_37_real = int_reg_array_3_37_real;
  assign io_coef_out_payload_0_3_37_imag = int_reg_array_3_37_imag;
  assign io_coef_out_payload_0_3_38_real = int_reg_array_3_38_real;
  assign io_coef_out_payload_0_3_38_imag = int_reg_array_3_38_imag;
  assign io_coef_out_payload_0_3_39_real = int_reg_array_3_39_real;
  assign io_coef_out_payload_0_3_39_imag = int_reg_array_3_39_imag;
  assign io_coef_out_payload_0_3_40_real = int_reg_array_3_40_real;
  assign io_coef_out_payload_0_3_40_imag = int_reg_array_3_40_imag;
  assign io_coef_out_payload_0_3_41_real = int_reg_array_3_41_real;
  assign io_coef_out_payload_0_3_41_imag = int_reg_array_3_41_imag;
  assign io_coef_out_payload_0_3_42_real = int_reg_array_3_42_real;
  assign io_coef_out_payload_0_3_42_imag = int_reg_array_3_42_imag;
  assign io_coef_out_payload_0_3_43_real = int_reg_array_3_43_real;
  assign io_coef_out_payload_0_3_43_imag = int_reg_array_3_43_imag;
  assign io_coef_out_payload_0_3_44_real = int_reg_array_3_44_real;
  assign io_coef_out_payload_0_3_44_imag = int_reg_array_3_44_imag;
  assign io_coef_out_payload_0_3_45_real = int_reg_array_3_45_real;
  assign io_coef_out_payload_0_3_45_imag = int_reg_array_3_45_imag;
  assign io_coef_out_payload_0_3_46_real = int_reg_array_3_46_real;
  assign io_coef_out_payload_0_3_46_imag = int_reg_array_3_46_imag;
  assign io_coef_out_payload_0_3_47_real = int_reg_array_3_47_real;
  assign io_coef_out_payload_0_3_47_imag = int_reg_array_3_47_imag;
  assign io_coef_out_payload_0_3_48_real = int_reg_array_3_48_real;
  assign io_coef_out_payload_0_3_48_imag = int_reg_array_3_48_imag;
  assign io_coef_out_payload_0_3_49_real = int_reg_array_3_49_real;
  assign io_coef_out_payload_0_3_49_imag = int_reg_array_3_49_imag;
  assign io_coef_out_payload_0_4_0_real = int_reg_array_4_0_real;
  assign io_coef_out_payload_0_4_0_imag = int_reg_array_4_0_imag;
  assign io_coef_out_payload_0_4_1_real = int_reg_array_4_1_real;
  assign io_coef_out_payload_0_4_1_imag = int_reg_array_4_1_imag;
  assign io_coef_out_payload_0_4_2_real = int_reg_array_4_2_real;
  assign io_coef_out_payload_0_4_2_imag = int_reg_array_4_2_imag;
  assign io_coef_out_payload_0_4_3_real = int_reg_array_4_3_real;
  assign io_coef_out_payload_0_4_3_imag = int_reg_array_4_3_imag;
  assign io_coef_out_payload_0_4_4_real = int_reg_array_4_4_real;
  assign io_coef_out_payload_0_4_4_imag = int_reg_array_4_4_imag;
  assign io_coef_out_payload_0_4_5_real = int_reg_array_4_5_real;
  assign io_coef_out_payload_0_4_5_imag = int_reg_array_4_5_imag;
  assign io_coef_out_payload_0_4_6_real = int_reg_array_4_6_real;
  assign io_coef_out_payload_0_4_6_imag = int_reg_array_4_6_imag;
  assign io_coef_out_payload_0_4_7_real = int_reg_array_4_7_real;
  assign io_coef_out_payload_0_4_7_imag = int_reg_array_4_7_imag;
  assign io_coef_out_payload_0_4_8_real = int_reg_array_4_8_real;
  assign io_coef_out_payload_0_4_8_imag = int_reg_array_4_8_imag;
  assign io_coef_out_payload_0_4_9_real = int_reg_array_4_9_real;
  assign io_coef_out_payload_0_4_9_imag = int_reg_array_4_9_imag;
  assign io_coef_out_payload_0_4_10_real = int_reg_array_4_10_real;
  assign io_coef_out_payload_0_4_10_imag = int_reg_array_4_10_imag;
  assign io_coef_out_payload_0_4_11_real = int_reg_array_4_11_real;
  assign io_coef_out_payload_0_4_11_imag = int_reg_array_4_11_imag;
  assign io_coef_out_payload_0_4_12_real = int_reg_array_4_12_real;
  assign io_coef_out_payload_0_4_12_imag = int_reg_array_4_12_imag;
  assign io_coef_out_payload_0_4_13_real = int_reg_array_4_13_real;
  assign io_coef_out_payload_0_4_13_imag = int_reg_array_4_13_imag;
  assign io_coef_out_payload_0_4_14_real = int_reg_array_4_14_real;
  assign io_coef_out_payload_0_4_14_imag = int_reg_array_4_14_imag;
  assign io_coef_out_payload_0_4_15_real = int_reg_array_4_15_real;
  assign io_coef_out_payload_0_4_15_imag = int_reg_array_4_15_imag;
  assign io_coef_out_payload_0_4_16_real = int_reg_array_4_16_real;
  assign io_coef_out_payload_0_4_16_imag = int_reg_array_4_16_imag;
  assign io_coef_out_payload_0_4_17_real = int_reg_array_4_17_real;
  assign io_coef_out_payload_0_4_17_imag = int_reg_array_4_17_imag;
  assign io_coef_out_payload_0_4_18_real = int_reg_array_4_18_real;
  assign io_coef_out_payload_0_4_18_imag = int_reg_array_4_18_imag;
  assign io_coef_out_payload_0_4_19_real = int_reg_array_4_19_real;
  assign io_coef_out_payload_0_4_19_imag = int_reg_array_4_19_imag;
  assign io_coef_out_payload_0_4_20_real = int_reg_array_4_20_real;
  assign io_coef_out_payload_0_4_20_imag = int_reg_array_4_20_imag;
  assign io_coef_out_payload_0_4_21_real = int_reg_array_4_21_real;
  assign io_coef_out_payload_0_4_21_imag = int_reg_array_4_21_imag;
  assign io_coef_out_payload_0_4_22_real = int_reg_array_4_22_real;
  assign io_coef_out_payload_0_4_22_imag = int_reg_array_4_22_imag;
  assign io_coef_out_payload_0_4_23_real = int_reg_array_4_23_real;
  assign io_coef_out_payload_0_4_23_imag = int_reg_array_4_23_imag;
  assign io_coef_out_payload_0_4_24_real = int_reg_array_4_24_real;
  assign io_coef_out_payload_0_4_24_imag = int_reg_array_4_24_imag;
  assign io_coef_out_payload_0_4_25_real = int_reg_array_4_25_real;
  assign io_coef_out_payload_0_4_25_imag = int_reg_array_4_25_imag;
  assign io_coef_out_payload_0_4_26_real = int_reg_array_4_26_real;
  assign io_coef_out_payload_0_4_26_imag = int_reg_array_4_26_imag;
  assign io_coef_out_payload_0_4_27_real = int_reg_array_4_27_real;
  assign io_coef_out_payload_0_4_27_imag = int_reg_array_4_27_imag;
  assign io_coef_out_payload_0_4_28_real = int_reg_array_4_28_real;
  assign io_coef_out_payload_0_4_28_imag = int_reg_array_4_28_imag;
  assign io_coef_out_payload_0_4_29_real = int_reg_array_4_29_real;
  assign io_coef_out_payload_0_4_29_imag = int_reg_array_4_29_imag;
  assign io_coef_out_payload_0_4_30_real = int_reg_array_4_30_real;
  assign io_coef_out_payload_0_4_30_imag = int_reg_array_4_30_imag;
  assign io_coef_out_payload_0_4_31_real = int_reg_array_4_31_real;
  assign io_coef_out_payload_0_4_31_imag = int_reg_array_4_31_imag;
  assign io_coef_out_payload_0_4_32_real = int_reg_array_4_32_real;
  assign io_coef_out_payload_0_4_32_imag = int_reg_array_4_32_imag;
  assign io_coef_out_payload_0_4_33_real = int_reg_array_4_33_real;
  assign io_coef_out_payload_0_4_33_imag = int_reg_array_4_33_imag;
  assign io_coef_out_payload_0_4_34_real = int_reg_array_4_34_real;
  assign io_coef_out_payload_0_4_34_imag = int_reg_array_4_34_imag;
  assign io_coef_out_payload_0_4_35_real = int_reg_array_4_35_real;
  assign io_coef_out_payload_0_4_35_imag = int_reg_array_4_35_imag;
  assign io_coef_out_payload_0_4_36_real = int_reg_array_4_36_real;
  assign io_coef_out_payload_0_4_36_imag = int_reg_array_4_36_imag;
  assign io_coef_out_payload_0_4_37_real = int_reg_array_4_37_real;
  assign io_coef_out_payload_0_4_37_imag = int_reg_array_4_37_imag;
  assign io_coef_out_payload_0_4_38_real = int_reg_array_4_38_real;
  assign io_coef_out_payload_0_4_38_imag = int_reg_array_4_38_imag;
  assign io_coef_out_payload_0_4_39_real = int_reg_array_4_39_real;
  assign io_coef_out_payload_0_4_39_imag = int_reg_array_4_39_imag;
  assign io_coef_out_payload_0_4_40_real = int_reg_array_4_40_real;
  assign io_coef_out_payload_0_4_40_imag = int_reg_array_4_40_imag;
  assign io_coef_out_payload_0_4_41_real = int_reg_array_4_41_real;
  assign io_coef_out_payload_0_4_41_imag = int_reg_array_4_41_imag;
  assign io_coef_out_payload_0_4_42_real = int_reg_array_4_42_real;
  assign io_coef_out_payload_0_4_42_imag = int_reg_array_4_42_imag;
  assign io_coef_out_payload_0_4_43_real = int_reg_array_4_43_real;
  assign io_coef_out_payload_0_4_43_imag = int_reg_array_4_43_imag;
  assign io_coef_out_payload_0_4_44_real = int_reg_array_4_44_real;
  assign io_coef_out_payload_0_4_44_imag = int_reg_array_4_44_imag;
  assign io_coef_out_payload_0_4_45_real = int_reg_array_4_45_real;
  assign io_coef_out_payload_0_4_45_imag = int_reg_array_4_45_imag;
  assign io_coef_out_payload_0_4_46_real = int_reg_array_4_46_real;
  assign io_coef_out_payload_0_4_46_imag = int_reg_array_4_46_imag;
  assign io_coef_out_payload_0_4_47_real = int_reg_array_4_47_real;
  assign io_coef_out_payload_0_4_47_imag = int_reg_array_4_47_imag;
  assign io_coef_out_payload_0_4_48_real = int_reg_array_4_48_real;
  assign io_coef_out_payload_0_4_48_imag = int_reg_array_4_48_imag;
  assign io_coef_out_payload_0_4_49_real = int_reg_array_4_49_real;
  assign io_coef_out_payload_0_4_49_imag = int_reg_array_4_49_imag;
  assign io_coef_out_payload_0_5_0_real = int_reg_array_5_0_real;
  assign io_coef_out_payload_0_5_0_imag = int_reg_array_5_0_imag;
  assign io_coef_out_payload_0_5_1_real = int_reg_array_5_1_real;
  assign io_coef_out_payload_0_5_1_imag = int_reg_array_5_1_imag;
  assign io_coef_out_payload_0_5_2_real = int_reg_array_5_2_real;
  assign io_coef_out_payload_0_5_2_imag = int_reg_array_5_2_imag;
  assign io_coef_out_payload_0_5_3_real = int_reg_array_5_3_real;
  assign io_coef_out_payload_0_5_3_imag = int_reg_array_5_3_imag;
  assign io_coef_out_payload_0_5_4_real = int_reg_array_5_4_real;
  assign io_coef_out_payload_0_5_4_imag = int_reg_array_5_4_imag;
  assign io_coef_out_payload_0_5_5_real = int_reg_array_5_5_real;
  assign io_coef_out_payload_0_5_5_imag = int_reg_array_5_5_imag;
  assign io_coef_out_payload_0_5_6_real = int_reg_array_5_6_real;
  assign io_coef_out_payload_0_5_6_imag = int_reg_array_5_6_imag;
  assign io_coef_out_payload_0_5_7_real = int_reg_array_5_7_real;
  assign io_coef_out_payload_0_5_7_imag = int_reg_array_5_7_imag;
  assign io_coef_out_payload_0_5_8_real = int_reg_array_5_8_real;
  assign io_coef_out_payload_0_5_8_imag = int_reg_array_5_8_imag;
  assign io_coef_out_payload_0_5_9_real = int_reg_array_5_9_real;
  assign io_coef_out_payload_0_5_9_imag = int_reg_array_5_9_imag;
  assign io_coef_out_payload_0_5_10_real = int_reg_array_5_10_real;
  assign io_coef_out_payload_0_5_10_imag = int_reg_array_5_10_imag;
  assign io_coef_out_payload_0_5_11_real = int_reg_array_5_11_real;
  assign io_coef_out_payload_0_5_11_imag = int_reg_array_5_11_imag;
  assign io_coef_out_payload_0_5_12_real = int_reg_array_5_12_real;
  assign io_coef_out_payload_0_5_12_imag = int_reg_array_5_12_imag;
  assign io_coef_out_payload_0_5_13_real = int_reg_array_5_13_real;
  assign io_coef_out_payload_0_5_13_imag = int_reg_array_5_13_imag;
  assign io_coef_out_payload_0_5_14_real = int_reg_array_5_14_real;
  assign io_coef_out_payload_0_5_14_imag = int_reg_array_5_14_imag;
  assign io_coef_out_payload_0_5_15_real = int_reg_array_5_15_real;
  assign io_coef_out_payload_0_5_15_imag = int_reg_array_5_15_imag;
  assign io_coef_out_payload_0_5_16_real = int_reg_array_5_16_real;
  assign io_coef_out_payload_0_5_16_imag = int_reg_array_5_16_imag;
  assign io_coef_out_payload_0_5_17_real = int_reg_array_5_17_real;
  assign io_coef_out_payload_0_5_17_imag = int_reg_array_5_17_imag;
  assign io_coef_out_payload_0_5_18_real = int_reg_array_5_18_real;
  assign io_coef_out_payload_0_5_18_imag = int_reg_array_5_18_imag;
  assign io_coef_out_payload_0_5_19_real = int_reg_array_5_19_real;
  assign io_coef_out_payload_0_5_19_imag = int_reg_array_5_19_imag;
  assign io_coef_out_payload_0_5_20_real = int_reg_array_5_20_real;
  assign io_coef_out_payload_0_5_20_imag = int_reg_array_5_20_imag;
  assign io_coef_out_payload_0_5_21_real = int_reg_array_5_21_real;
  assign io_coef_out_payload_0_5_21_imag = int_reg_array_5_21_imag;
  assign io_coef_out_payload_0_5_22_real = int_reg_array_5_22_real;
  assign io_coef_out_payload_0_5_22_imag = int_reg_array_5_22_imag;
  assign io_coef_out_payload_0_5_23_real = int_reg_array_5_23_real;
  assign io_coef_out_payload_0_5_23_imag = int_reg_array_5_23_imag;
  assign io_coef_out_payload_0_5_24_real = int_reg_array_5_24_real;
  assign io_coef_out_payload_0_5_24_imag = int_reg_array_5_24_imag;
  assign io_coef_out_payload_0_5_25_real = int_reg_array_5_25_real;
  assign io_coef_out_payload_0_5_25_imag = int_reg_array_5_25_imag;
  assign io_coef_out_payload_0_5_26_real = int_reg_array_5_26_real;
  assign io_coef_out_payload_0_5_26_imag = int_reg_array_5_26_imag;
  assign io_coef_out_payload_0_5_27_real = int_reg_array_5_27_real;
  assign io_coef_out_payload_0_5_27_imag = int_reg_array_5_27_imag;
  assign io_coef_out_payload_0_5_28_real = int_reg_array_5_28_real;
  assign io_coef_out_payload_0_5_28_imag = int_reg_array_5_28_imag;
  assign io_coef_out_payload_0_5_29_real = int_reg_array_5_29_real;
  assign io_coef_out_payload_0_5_29_imag = int_reg_array_5_29_imag;
  assign io_coef_out_payload_0_5_30_real = int_reg_array_5_30_real;
  assign io_coef_out_payload_0_5_30_imag = int_reg_array_5_30_imag;
  assign io_coef_out_payload_0_5_31_real = int_reg_array_5_31_real;
  assign io_coef_out_payload_0_5_31_imag = int_reg_array_5_31_imag;
  assign io_coef_out_payload_0_5_32_real = int_reg_array_5_32_real;
  assign io_coef_out_payload_0_5_32_imag = int_reg_array_5_32_imag;
  assign io_coef_out_payload_0_5_33_real = int_reg_array_5_33_real;
  assign io_coef_out_payload_0_5_33_imag = int_reg_array_5_33_imag;
  assign io_coef_out_payload_0_5_34_real = int_reg_array_5_34_real;
  assign io_coef_out_payload_0_5_34_imag = int_reg_array_5_34_imag;
  assign io_coef_out_payload_0_5_35_real = int_reg_array_5_35_real;
  assign io_coef_out_payload_0_5_35_imag = int_reg_array_5_35_imag;
  assign io_coef_out_payload_0_5_36_real = int_reg_array_5_36_real;
  assign io_coef_out_payload_0_5_36_imag = int_reg_array_5_36_imag;
  assign io_coef_out_payload_0_5_37_real = int_reg_array_5_37_real;
  assign io_coef_out_payload_0_5_37_imag = int_reg_array_5_37_imag;
  assign io_coef_out_payload_0_5_38_real = int_reg_array_5_38_real;
  assign io_coef_out_payload_0_5_38_imag = int_reg_array_5_38_imag;
  assign io_coef_out_payload_0_5_39_real = int_reg_array_5_39_real;
  assign io_coef_out_payload_0_5_39_imag = int_reg_array_5_39_imag;
  assign io_coef_out_payload_0_5_40_real = int_reg_array_5_40_real;
  assign io_coef_out_payload_0_5_40_imag = int_reg_array_5_40_imag;
  assign io_coef_out_payload_0_5_41_real = int_reg_array_5_41_real;
  assign io_coef_out_payload_0_5_41_imag = int_reg_array_5_41_imag;
  assign io_coef_out_payload_0_5_42_real = int_reg_array_5_42_real;
  assign io_coef_out_payload_0_5_42_imag = int_reg_array_5_42_imag;
  assign io_coef_out_payload_0_5_43_real = int_reg_array_5_43_real;
  assign io_coef_out_payload_0_5_43_imag = int_reg_array_5_43_imag;
  assign io_coef_out_payload_0_5_44_real = int_reg_array_5_44_real;
  assign io_coef_out_payload_0_5_44_imag = int_reg_array_5_44_imag;
  assign io_coef_out_payload_0_5_45_real = int_reg_array_5_45_real;
  assign io_coef_out_payload_0_5_45_imag = int_reg_array_5_45_imag;
  assign io_coef_out_payload_0_5_46_real = int_reg_array_5_46_real;
  assign io_coef_out_payload_0_5_46_imag = int_reg_array_5_46_imag;
  assign io_coef_out_payload_0_5_47_real = int_reg_array_5_47_real;
  assign io_coef_out_payload_0_5_47_imag = int_reg_array_5_47_imag;
  assign io_coef_out_payload_0_5_48_real = int_reg_array_5_48_real;
  assign io_coef_out_payload_0_5_48_imag = int_reg_array_5_48_imag;
  assign io_coef_out_payload_0_5_49_real = int_reg_array_5_49_real;
  assign io_coef_out_payload_0_5_49_imag = int_reg_array_5_49_imag;
  assign io_coef_out_payload_0_6_0_real = int_reg_array_6_0_real;
  assign io_coef_out_payload_0_6_0_imag = int_reg_array_6_0_imag;
  assign io_coef_out_payload_0_6_1_real = int_reg_array_6_1_real;
  assign io_coef_out_payload_0_6_1_imag = int_reg_array_6_1_imag;
  assign io_coef_out_payload_0_6_2_real = int_reg_array_6_2_real;
  assign io_coef_out_payload_0_6_2_imag = int_reg_array_6_2_imag;
  assign io_coef_out_payload_0_6_3_real = int_reg_array_6_3_real;
  assign io_coef_out_payload_0_6_3_imag = int_reg_array_6_3_imag;
  assign io_coef_out_payload_0_6_4_real = int_reg_array_6_4_real;
  assign io_coef_out_payload_0_6_4_imag = int_reg_array_6_4_imag;
  assign io_coef_out_payload_0_6_5_real = int_reg_array_6_5_real;
  assign io_coef_out_payload_0_6_5_imag = int_reg_array_6_5_imag;
  assign io_coef_out_payload_0_6_6_real = int_reg_array_6_6_real;
  assign io_coef_out_payload_0_6_6_imag = int_reg_array_6_6_imag;
  assign io_coef_out_payload_0_6_7_real = int_reg_array_6_7_real;
  assign io_coef_out_payload_0_6_7_imag = int_reg_array_6_7_imag;
  assign io_coef_out_payload_0_6_8_real = int_reg_array_6_8_real;
  assign io_coef_out_payload_0_6_8_imag = int_reg_array_6_8_imag;
  assign io_coef_out_payload_0_6_9_real = int_reg_array_6_9_real;
  assign io_coef_out_payload_0_6_9_imag = int_reg_array_6_9_imag;
  assign io_coef_out_payload_0_6_10_real = int_reg_array_6_10_real;
  assign io_coef_out_payload_0_6_10_imag = int_reg_array_6_10_imag;
  assign io_coef_out_payload_0_6_11_real = int_reg_array_6_11_real;
  assign io_coef_out_payload_0_6_11_imag = int_reg_array_6_11_imag;
  assign io_coef_out_payload_0_6_12_real = int_reg_array_6_12_real;
  assign io_coef_out_payload_0_6_12_imag = int_reg_array_6_12_imag;
  assign io_coef_out_payload_0_6_13_real = int_reg_array_6_13_real;
  assign io_coef_out_payload_0_6_13_imag = int_reg_array_6_13_imag;
  assign io_coef_out_payload_0_6_14_real = int_reg_array_6_14_real;
  assign io_coef_out_payload_0_6_14_imag = int_reg_array_6_14_imag;
  assign io_coef_out_payload_0_6_15_real = int_reg_array_6_15_real;
  assign io_coef_out_payload_0_6_15_imag = int_reg_array_6_15_imag;
  assign io_coef_out_payload_0_6_16_real = int_reg_array_6_16_real;
  assign io_coef_out_payload_0_6_16_imag = int_reg_array_6_16_imag;
  assign io_coef_out_payload_0_6_17_real = int_reg_array_6_17_real;
  assign io_coef_out_payload_0_6_17_imag = int_reg_array_6_17_imag;
  assign io_coef_out_payload_0_6_18_real = int_reg_array_6_18_real;
  assign io_coef_out_payload_0_6_18_imag = int_reg_array_6_18_imag;
  assign io_coef_out_payload_0_6_19_real = int_reg_array_6_19_real;
  assign io_coef_out_payload_0_6_19_imag = int_reg_array_6_19_imag;
  assign io_coef_out_payload_0_6_20_real = int_reg_array_6_20_real;
  assign io_coef_out_payload_0_6_20_imag = int_reg_array_6_20_imag;
  assign io_coef_out_payload_0_6_21_real = int_reg_array_6_21_real;
  assign io_coef_out_payload_0_6_21_imag = int_reg_array_6_21_imag;
  assign io_coef_out_payload_0_6_22_real = int_reg_array_6_22_real;
  assign io_coef_out_payload_0_6_22_imag = int_reg_array_6_22_imag;
  assign io_coef_out_payload_0_6_23_real = int_reg_array_6_23_real;
  assign io_coef_out_payload_0_6_23_imag = int_reg_array_6_23_imag;
  assign io_coef_out_payload_0_6_24_real = int_reg_array_6_24_real;
  assign io_coef_out_payload_0_6_24_imag = int_reg_array_6_24_imag;
  assign io_coef_out_payload_0_6_25_real = int_reg_array_6_25_real;
  assign io_coef_out_payload_0_6_25_imag = int_reg_array_6_25_imag;
  assign io_coef_out_payload_0_6_26_real = int_reg_array_6_26_real;
  assign io_coef_out_payload_0_6_26_imag = int_reg_array_6_26_imag;
  assign io_coef_out_payload_0_6_27_real = int_reg_array_6_27_real;
  assign io_coef_out_payload_0_6_27_imag = int_reg_array_6_27_imag;
  assign io_coef_out_payload_0_6_28_real = int_reg_array_6_28_real;
  assign io_coef_out_payload_0_6_28_imag = int_reg_array_6_28_imag;
  assign io_coef_out_payload_0_6_29_real = int_reg_array_6_29_real;
  assign io_coef_out_payload_0_6_29_imag = int_reg_array_6_29_imag;
  assign io_coef_out_payload_0_6_30_real = int_reg_array_6_30_real;
  assign io_coef_out_payload_0_6_30_imag = int_reg_array_6_30_imag;
  assign io_coef_out_payload_0_6_31_real = int_reg_array_6_31_real;
  assign io_coef_out_payload_0_6_31_imag = int_reg_array_6_31_imag;
  assign io_coef_out_payload_0_6_32_real = int_reg_array_6_32_real;
  assign io_coef_out_payload_0_6_32_imag = int_reg_array_6_32_imag;
  assign io_coef_out_payload_0_6_33_real = int_reg_array_6_33_real;
  assign io_coef_out_payload_0_6_33_imag = int_reg_array_6_33_imag;
  assign io_coef_out_payload_0_6_34_real = int_reg_array_6_34_real;
  assign io_coef_out_payload_0_6_34_imag = int_reg_array_6_34_imag;
  assign io_coef_out_payload_0_6_35_real = int_reg_array_6_35_real;
  assign io_coef_out_payload_0_6_35_imag = int_reg_array_6_35_imag;
  assign io_coef_out_payload_0_6_36_real = int_reg_array_6_36_real;
  assign io_coef_out_payload_0_6_36_imag = int_reg_array_6_36_imag;
  assign io_coef_out_payload_0_6_37_real = int_reg_array_6_37_real;
  assign io_coef_out_payload_0_6_37_imag = int_reg_array_6_37_imag;
  assign io_coef_out_payload_0_6_38_real = int_reg_array_6_38_real;
  assign io_coef_out_payload_0_6_38_imag = int_reg_array_6_38_imag;
  assign io_coef_out_payload_0_6_39_real = int_reg_array_6_39_real;
  assign io_coef_out_payload_0_6_39_imag = int_reg_array_6_39_imag;
  assign io_coef_out_payload_0_6_40_real = int_reg_array_6_40_real;
  assign io_coef_out_payload_0_6_40_imag = int_reg_array_6_40_imag;
  assign io_coef_out_payload_0_6_41_real = int_reg_array_6_41_real;
  assign io_coef_out_payload_0_6_41_imag = int_reg_array_6_41_imag;
  assign io_coef_out_payload_0_6_42_real = int_reg_array_6_42_real;
  assign io_coef_out_payload_0_6_42_imag = int_reg_array_6_42_imag;
  assign io_coef_out_payload_0_6_43_real = int_reg_array_6_43_real;
  assign io_coef_out_payload_0_6_43_imag = int_reg_array_6_43_imag;
  assign io_coef_out_payload_0_6_44_real = int_reg_array_6_44_real;
  assign io_coef_out_payload_0_6_44_imag = int_reg_array_6_44_imag;
  assign io_coef_out_payload_0_6_45_real = int_reg_array_6_45_real;
  assign io_coef_out_payload_0_6_45_imag = int_reg_array_6_45_imag;
  assign io_coef_out_payload_0_6_46_real = int_reg_array_6_46_real;
  assign io_coef_out_payload_0_6_46_imag = int_reg_array_6_46_imag;
  assign io_coef_out_payload_0_6_47_real = int_reg_array_6_47_real;
  assign io_coef_out_payload_0_6_47_imag = int_reg_array_6_47_imag;
  assign io_coef_out_payload_0_6_48_real = int_reg_array_6_48_real;
  assign io_coef_out_payload_0_6_48_imag = int_reg_array_6_48_imag;
  assign io_coef_out_payload_0_6_49_real = int_reg_array_6_49_real;
  assign io_coef_out_payload_0_6_49_imag = int_reg_array_6_49_imag;
  assign io_coef_out_payload_0_7_0_real = int_reg_array_7_0_real;
  assign io_coef_out_payload_0_7_0_imag = int_reg_array_7_0_imag;
  assign io_coef_out_payload_0_7_1_real = int_reg_array_7_1_real;
  assign io_coef_out_payload_0_7_1_imag = int_reg_array_7_1_imag;
  assign io_coef_out_payload_0_7_2_real = int_reg_array_7_2_real;
  assign io_coef_out_payload_0_7_2_imag = int_reg_array_7_2_imag;
  assign io_coef_out_payload_0_7_3_real = int_reg_array_7_3_real;
  assign io_coef_out_payload_0_7_3_imag = int_reg_array_7_3_imag;
  assign io_coef_out_payload_0_7_4_real = int_reg_array_7_4_real;
  assign io_coef_out_payload_0_7_4_imag = int_reg_array_7_4_imag;
  assign io_coef_out_payload_0_7_5_real = int_reg_array_7_5_real;
  assign io_coef_out_payload_0_7_5_imag = int_reg_array_7_5_imag;
  assign io_coef_out_payload_0_7_6_real = int_reg_array_7_6_real;
  assign io_coef_out_payload_0_7_6_imag = int_reg_array_7_6_imag;
  assign io_coef_out_payload_0_7_7_real = int_reg_array_7_7_real;
  assign io_coef_out_payload_0_7_7_imag = int_reg_array_7_7_imag;
  assign io_coef_out_payload_0_7_8_real = int_reg_array_7_8_real;
  assign io_coef_out_payload_0_7_8_imag = int_reg_array_7_8_imag;
  assign io_coef_out_payload_0_7_9_real = int_reg_array_7_9_real;
  assign io_coef_out_payload_0_7_9_imag = int_reg_array_7_9_imag;
  assign io_coef_out_payload_0_7_10_real = int_reg_array_7_10_real;
  assign io_coef_out_payload_0_7_10_imag = int_reg_array_7_10_imag;
  assign io_coef_out_payload_0_7_11_real = int_reg_array_7_11_real;
  assign io_coef_out_payload_0_7_11_imag = int_reg_array_7_11_imag;
  assign io_coef_out_payload_0_7_12_real = int_reg_array_7_12_real;
  assign io_coef_out_payload_0_7_12_imag = int_reg_array_7_12_imag;
  assign io_coef_out_payload_0_7_13_real = int_reg_array_7_13_real;
  assign io_coef_out_payload_0_7_13_imag = int_reg_array_7_13_imag;
  assign io_coef_out_payload_0_7_14_real = int_reg_array_7_14_real;
  assign io_coef_out_payload_0_7_14_imag = int_reg_array_7_14_imag;
  assign io_coef_out_payload_0_7_15_real = int_reg_array_7_15_real;
  assign io_coef_out_payload_0_7_15_imag = int_reg_array_7_15_imag;
  assign io_coef_out_payload_0_7_16_real = int_reg_array_7_16_real;
  assign io_coef_out_payload_0_7_16_imag = int_reg_array_7_16_imag;
  assign io_coef_out_payload_0_7_17_real = int_reg_array_7_17_real;
  assign io_coef_out_payload_0_7_17_imag = int_reg_array_7_17_imag;
  assign io_coef_out_payload_0_7_18_real = int_reg_array_7_18_real;
  assign io_coef_out_payload_0_7_18_imag = int_reg_array_7_18_imag;
  assign io_coef_out_payload_0_7_19_real = int_reg_array_7_19_real;
  assign io_coef_out_payload_0_7_19_imag = int_reg_array_7_19_imag;
  assign io_coef_out_payload_0_7_20_real = int_reg_array_7_20_real;
  assign io_coef_out_payload_0_7_20_imag = int_reg_array_7_20_imag;
  assign io_coef_out_payload_0_7_21_real = int_reg_array_7_21_real;
  assign io_coef_out_payload_0_7_21_imag = int_reg_array_7_21_imag;
  assign io_coef_out_payload_0_7_22_real = int_reg_array_7_22_real;
  assign io_coef_out_payload_0_7_22_imag = int_reg_array_7_22_imag;
  assign io_coef_out_payload_0_7_23_real = int_reg_array_7_23_real;
  assign io_coef_out_payload_0_7_23_imag = int_reg_array_7_23_imag;
  assign io_coef_out_payload_0_7_24_real = int_reg_array_7_24_real;
  assign io_coef_out_payload_0_7_24_imag = int_reg_array_7_24_imag;
  assign io_coef_out_payload_0_7_25_real = int_reg_array_7_25_real;
  assign io_coef_out_payload_0_7_25_imag = int_reg_array_7_25_imag;
  assign io_coef_out_payload_0_7_26_real = int_reg_array_7_26_real;
  assign io_coef_out_payload_0_7_26_imag = int_reg_array_7_26_imag;
  assign io_coef_out_payload_0_7_27_real = int_reg_array_7_27_real;
  assign io_coef_out_payload_0_7_27_imag = int_reg_array_7_27_imag;
  assign io_coef_out_payload_0_7_28_real = int_reg_array_7_28_real;
  assign io_coef_out_payload_0_7_28_imag = int_reg_array_7_28_imag;
  assign io_coef_out_payload_0_7_29_real = int_reg_array_7_29_real;
  assign io_coef_out_payload_0_7_29_imag = int_reg_array_7_29_imag;
  assign io_coef_out_payload_0_7_30_real = int_reg_array_7_30_real;
  assign io_coef_out_payload_0_7_30_imag = int_reg_array_7_30_imag;
  assign io_coef_out_payload_0_7_31_real = int_reg_array_7_31_real;
  assign io_coef_out_payload_0_7_31_imag = int_reg_array_7_31_imag;
  assign io_coef_out_payload_0_7_32_real = int_reg_array_7_32_real;
  assign io_coef_out_payload_0_7_32_imag = int_reg_array_7_32_imag;
  assign io_coef_out_payload_0_7_33_real = int_reg_array_7_33_real;
  assign io_coef_out_payload_0_7_33_imag = int_reg_array_7_33_imag;
  assign io_coef_out_payload_0_7_34_real = int_reg_array_7_34_real;
  assign io_coef_out_payload_0_7_34_imag = int_reg_array_7_34_imag;
  assign io_coef_out_payload_0_7_35_real = int_reg_array_7_35_real;
  assign io_coef_out_payload_0_7_35_imag = int_reg_array_7_35_imag;
  assign io_coef_out_payload_0_7_36_real = int_reg_array_7_36_real;
  assign io_coef_out_payload_0_7_36_imag = int_reg_array_7_36_imag;
  assign io_coef_out_payload_0_7_37_real = int_reg_array_7_37_real;
  assign io_coef_out_payload_0_7_37_imag = int_reg_array_7_37_imag;
  assign io_coef_out_payload_0_7_38_real = int_reg_array_7_38_real;
  assign io_coef_out_payload_0_7_38_imag = int_reg_array_7_38_imag;
  assign io_coef_out_payload_0_7_39_real = int_reg_array_7_39_real;
  assign io_coef_out_payload_0_7_39_imag = int_reg_array_7_39_imag;
  assign io_coef_out_payload_0_7_40_real = int_reg_array_7_40_real;
  assign io_coef_out_payload_0_7_40_imag = int_reg_array_7_40_imag;
  assign io_coef_out_payload_0_7_41_real = int_reg_array_7_41_real;
  assign io_coef_out_payload_0_7_41_imag = int_reg_array_7_41_imag;
  assign io_coef_out_payload_0_7_42_real = int_reg_array_7_42_real;
  assign io_coef_out_payload_0_7_42_imag = int_reg_array_7_42_imag;
  assign io_coef_out_payload_0_7_43_real = int_reg_array_7_43_real;
  assign io_coef_out_payload_0_7_43_imag = int_reg_array_7_43_imag;
  assign io_coef_out_payload_0_7_44_real = int_reg_array_7_44_real;
  assign io_coef_out_payload_0_7_44_imag = int_reg_array_7_44_imag;
  assign io_coef_out_payload_0_7_45_real = int_reg_array_7_45_real;
  assign io_coef_out_payload_0_7_45_imag = int_reg_array_7_45_imag;
  assign io_coef_out_payload_0_7_46_real = int_reg_array_7_46_real;
  assign io_coef_out_payload_0_7_46_imag = int_reg_array_7_46_imag;
  assign io_coef_out_payload_0_7_47_real = int_reg_array_7_47_real;
  assign io_coef_out_payload_0_7_47_imag = int_reg_array_7_47_imag;
  assign io_coef_out_payload_0_7_48_real = int_reg_array_7_48_real;
  assign io_coef_out_payload_0_7_48_imag = int_reg_array_7_48_imag;
  assign io_coef_out_payload_0_7_49_real = int_reg_array_7_49_real;
  assign io_coef_out_payload_0_7_49_imag = int_reg_array_7_49_imag;
  assign io_coef_out_payload_0_8_0_real = int_reg_array_8_0_real;
  assign io_coef_out_payload_0_8_0_imag = int_reg_array_8_0_imag;
  assign io_coef_out_payload_0_8_1_real = int_reg_array_8_1_real;
  assign io_coef_out_payload_0_8_1_imag = int_reg_array_8_1_imag;
  assign io_coef_out_payload_0_8_2_real = int_reg_array_8_2_real;
  assign io_coef_out_payload_0_8_2_imag = int_reg_array_8_2_imag;
  assign io_coef_out_payload_0_8_3_real = int_reg_array_8_3_real;
  assign io_coef_out_payload_0_8_3_imag = int_reg_array_8_3_imag;
  assign io_coef_out_payload_0_8_4_real = int_reg_array_8_4_real;
  assign io_coef_out_payload_0_8_4_imag = int_reg_array_8_4_imag;
  assign io_coef_out_payload_0_8_5_real = int_reg_array_8_5_real;
  assign io_coef_out_payload_0_8_5_imag = int_reg_array_8_5_imag;
  assign io_coef_out_payload_0_8_6_real = int_reg_array_8_6_real;
  assign io_coef_out_payload_0_8_6_imag = int_reg_array_8_6_imag;
  assign io_coef_out_payload_0_8_7_real = int_reg_array_8_7_real;
  assign io_coef_out_payload_0_8_7_imag = int_reg_array_8_7_imag;
  assign io_coef_out_payload_0_8_8_real = int_reg_array_8_8_real;
  assign io_coef_out_payload_0_8_8_imag = int_reg_array_8_8_imag;
  assign io_coef_out_payload_0_8_9_real = int_reg_array_8_9_real;
  assign io_coef_out_payload_0_8_9_imag = int_reg_array_8_9_imag;
  assign io_coef_out_payload_0_8_10_real = int_reg_array_8_10_real;
  assign io_coef_out_payload_0_8_10_imag = int_reg_array_8_10_imag;
  assign io_coef_out_payload_0_8_11_real = int_reg_array_8_11_real;
  assign io_coef_out_payload_0_8_11_imag = int_reg_array_8_11_imag;
  assign io_coef_out_payload_0_8_12_real = int_reg_array_8_12_real;
  assign io_coef_out_payload_0_8_12_imag = int_reg_array_8_12_imag;
  assign io_coef_out_payload_0_8_13_real = int_reg_array_8_13_real;
  assign io_coef_out_payload_0_8_13_imag = int_reg_array_8_13_imag;
  assign io_coef_out_payload_0_8_14_real = int_reg_array_8_14_real;
  assign io_coef_out_payload_0_8_14_imag = int_reg_array_8_14_imag;
  assign io_coef_out_payload_0_8_15_real = int_reg_array_8_15_real;
  assign io_coef_out_payload_0_8_15_imag = int_reg_array_8_15_imag;
  assign io_coef_out_payload_0_8_16_real = int_reg_array_8_16_real;
  assign io_coef_out_payload_0_8_16_imag = int_reg_array_8_16_imag;
  assign io_coef_out_payload_0_8_17_real = int_reg_array_8_17_real;
  assign io_coef_out_payload_0_8_17_imag = int_reg_array_8_17_imag;
  assign io_coef_out_payload_0_8_18_real = int_reg_array_8_18_real;
  assign io_coef_out_payload_0_8_18_imag = int_reg_array_8_18_imag;
  assign io_coef_out_payload_0_8_19_real = int_reg_array_8_19_real;
  assign io_coef_out_payload_0_8_19_imag = int_reg_array_8_19_imag;
  assign io_coef_out_payload_0_8_20_real = int_reg_array_8_20_real;
  assign io_coef_out_payload_0_8_20_imag = int_reg_array_8_20_imag;
  assign io_coef_out_payload_0_8_21_real = int_reg_array_8_21_real;
  assign io_coef_out_payload_0_8_21_imag = int_reg_array_8_21_imag;
  assign io_coef_out_payload_0_8_22_real = int_reg_array_8_22_real;
  assign io_coef_out_payload_0_8_22_imag = int_reg_array_8_22_imag;
  assign io_coef_out_payload_0_8_23_real = int_reg_array_8_23_real;
  assign io_coef_out_payload_0_8_23_imag = int_reg_array_8_23_imag;
  assign io_coef_out_payload_0_8_24_real = int_reg_array_8_24_real;
  assign io_coef_out_payload_0_8_24_imag = int_reg_array_8_24_imag;
  assign io_coef_out_payload_0_8_25_real = int_reg_array_8_25_real;
  assign io_coef_out_payload_0_8_25_imag = int_reg_array_8_25_imag;
  assign io_coef_out_payload_0_8_26_real = int_reg_array_8_26_real;
  assign io_coef_out_payload_0_8_26_imag = int_reg_array_8_26_imag;
  assign io_coef_out_payload_0_8_27_real = int_reg_array_8_27_real;
  assign io_coef_out_payload_0_8_27_imag = int_reg_array_8_27_imag;
  assign io_coef_out_payload_0_8_28_real = int_reg_array_8_28_real;
  assign io_coef_out_payload_0_8_28_imag = int_reg_array_8_28_imag;
  assign io_coef_out_payload_0_8_29_real = int_reg_array_8_29_real;
  assign io_coef_out_payload_0_8_29_imag = int_reg_array_8_29_imag;
  assign io_coef_out_payload_0_8_30_real = int_reg_array_8_30_real;
  assign io_coef_out_payload_0_8_30_imag = int_reg_array_8_30_imag;
  assign io_coef_out_payload_0_8_31_real = int_reg_array_8_31_real;
  assign io_coef_out_payload_0_8_31_imag = int_reg_array_8_31_imag;
  assign io_coef_out_payload_0_8_32_real = int_reg_array_8_32_real;
  assign io_coef_out_payload_0_8_32_imag = int_reg_array_8_32_imag;
  assign io_coef_out_payload_0_8_33_real = int_reg_array_8_33_real;
  assign io_coef_out_payload_0_8_33_imag = int_reg_array_8_33_imag;
  assign io_coef_out_payload_0_8_34_real = int_reg_array_8_34_real;
  assign io_coef_out_payload_0_8_34_imag = int_reg_array_8_34_imag;
  assign io_coef_out_payload_0_8_35_real = int_reg_array_8_35_real;
  assign io_coef_out_payload_0_8_35_imag = int_reg_array_8_35_imag;
  assign io_coef_out_payload_0_8_36_real = int_reg_array_8_36_real;
  assign io_coef_out_payload_0_8_36_imag = int_reg_array_8_36_imag;
  assign io_coef_out_payload_0_8_37_real = int_reg_array_8_37_real;
  assign io_coef_out_payload_0_8_37_imag = int_reg_array_8_37_imag;
  assign io_coef_out_payload_0_8_38_real = int_reg_array_8_38_real;
  assign io_coef_out_payload_0_8_38_imag = int_reg_array_8_38_imag;
  assign io_coef_out_payload_0_8_39_real = int_reg_array_8_39_real;
  assign io_coef_out_payload_0_8_39_imag = int_reg_array_8_39_imag;
  assign io_coef_out_payload_0_8_40_real = int_reg_array_8_40_real;
  assign io_coef_out_payload_0_8_40_imag = int_reg_array_8_40_imag;
  assign io_coef_out_payload_0_8_41_real = int_reg_array_8_41_real;
  assign io_coef_out_payload_0_8_41_imag = int_reg_array_8_41_imag;
  assign io_coef_out_payload_0_8_42_real = int_reg_array_8_42_real;
  assign io_coef_out_payload_0_8_42_imag = int_reg_array_8_42_imag;
  assign io_coef_out_payload_0_8_43_real = int_reg_array_8_43_real;
  assign io_coef_out_payload_0_8_43_imag = int_reg_array_8_43_imag;
  assign io_coef_out_payload_0_8_44_real = int_reg_array_8_44_real;
  assign io_coef_out_payload_0_8_44_imag = int_reg_array_8_44_imag;
  assign io_coef_out_payload_0_8_45_real = int_reg_array_8_45_real;
  assign io_coef_out_payload_0_8_45_imag = int_reg_array_8_45_imag;
  assign io_coef_out_payload_0_8_46_real = int_reg_array_8_46_real;
  assign io_coef_out_payload_0_8_46_imag = int_reg_array_8_46_imag;
  assign io_coef_out_payload_0_8_47_real = int_reg_array_8_47_real;
  assign io_coef_out_payload_0_8_47_imag = int_reg_array_8_47_imag;
  assign io_coef_out_payload_0_8_48_real = int_reg_array_8_48_real;
  assign io_coef_out_payload_0_8_48_imag = int_reg_array_8_48_imag;
  assign io_coef_out_payload_0_8_49_real = int_reg_array_8_49_real;
  assign io_coef_out_payload_0_8_49_imag = int_reg_array_8_49_imag;
  assign io_coef_out_payload_0_9_0_real = int_reg_array_9_0_real;
  assign io_coef_out_payload_0_9_0_imag = int_reg_array_9_0_imag;
  assign io_coef_out_payload_0_9_1_real = int_reg_array_9_1_real;
  assign io_coef_out_payload_0_9_1_imag = int_reg_array_9_1_imag;
  assign io_coef_out_payload_0_9_2_real = int_reg_array_9_2_real;
  assign io_coef_out_payload_0_9_2_imag = int_reg_array_9_2_imag;
  assign io_coef_out_payload_0_9_3_real = int_reg_array_9_3_real;
  assign io_coef_out_payload_0_9_3_imag = int_reg_array_9_3_imag;
  assign io_coef_out_payload_0_9_4_real = int_reg_array_9_4_real;
  assign io_coef_out_payload_0_9_4_imag = int_reg_array_9_4_imag;
  assign io_coef_out_payload_0_9_5_real = int_reg_array_9_5_real;
  assign io_coef_out_payload_0_9_5_imag = int_reg_array_9_5_imag;
  assign io_coef_out_payload_0_9_6_real = int_reg_array_9_6_real;
  assign io_coef_out_payload_0_9_6_imag = int_reg_array_9_6_imag;
  assign io_coef_out_payload_0_9_7_real = int_reg_array_9_7_real;
  assign io_coef_out_payload_0_9_7_imag = int_reg_array_9_7_imag;
  assign io_coef_out_payload_0_9_8_real = int_reg_array_9_8_real;
  assign io_coef_out_payload_0_9_8_imag = int_reg_array_9_8_imag;
  assign io_coef_out_payload_0_9_9_real = int_reg_array_9_9_real;
  assign io_coef_out_payload_0_9_9_imag = int_reg_array_9_9_imag;
  assign io_coef_out_payload_0_9_10_real = int_reg_array_9_10_real;
  assign io_coef_out_payload_0_9_10_imag = int_reg_array_9_10_imag;
  assign io_coef_out_payload_0_9_11_real = int_reg_array_9_11_real;
  assign io_coef_out_payload_0_9_11_imag = int_reg_array_9_11_imag;
  assign io_coef_out_payload_0_9_12_real = int_reg_array_9_12_real;
  assign io_coef_out_payload_0_9_12_imag = int_reg_array_9_12_imag;
  assign io_coef_out_payload_0_9_13_real = int_reg_array_9_13_real;
  assign io_coef_out_payload_0_9_13_imag = int_reg_array_9_13_imag;
  assign io_coef_out_payload_0_9_14_real = int_reg_array_9_14_real;
  assign io_coef_out_payload_0_9_14_imag = int_reg_array_9_14_imag;
  assign io_coef_out_payload_0_9_15_real = int_reg_array_9_15_real;
  assign io_coef_out_payload_0_9_15_imag = int_reg_array_9_15_imag;
  assign io_coef_out_payload_0_9_16_real = int_reg_array_9_16_real;
  assign io_coef_out_payload_0_9_16_imag = int_reg_array_9_16_imag;
  assign io_coef_out_payload_0_9_17_real = int_reg_array_9_17_real;
  assign io_coef_out_payload_0_9_17_imag = int_reg_array_9_17_imag;
  assign io_coef_out_payload_0_9_18_real = int_reg_array_9_18_real;
  assign io_coef_out_payload_0_9_18_imag = int_reg_array_9_18_imag;
  assign io_coef_out_payload_0_9_19_real = int_reg_array_9_19_real;
  assign io_coef_out_payload_0_9_19_imag = int_reg_array_9_19_imag;
  assign io_coef_out_payload_0_9_20_real = int_reg_array_9_20_real;
  assign io_coef_out_payload_0_9_20_imag = int_reg_array_9_20_imag;
  assign io_coef_out_payload_0_9_21_real = int_reg_array_9_21_real;
  assign io_coef_out_payload_0_9_21_imag = int_reg_array_9_21_imag;
  assign io_coef_out_payload_0_9_22_real = int_reg_array_9_22_real;
  assign io_coef_out_payload_0_9_22_imag = int_reg_array_9_22_imag;
  assign io_coef_out_payload_0_9_23_real = int_reg_array_9_23_real;
  assign io_coef_out_payload_0_9_23_imag = int_reg_array_9_23_imag;
  assign io_coef_out_payload_0_9_24_real = int_reg_array_9_24_real;
  assign io_coef_out_payload_0_9_24_imag = int_reg_array_9_24_imag;
  assign io_coef_out_payload_0_9_25_real = int_reg_array_9_25_real;
  assign io_coef_out_payload_0_9_25_imag = int_reg_array_9_25_imag;
  assign io_coef_out_payload_0_9_26_real = int_reg_array_9_26_real;
  assign io_coef_out_payload_0_9_26_imag = int_reg_array_9_26_imag;
  assign io_coef_out_payload_0_9_27_real = int_reg_array_9_27_real;
  assign io_coef_out_payload_0_9_27_imag = int_reg_array_9_27_imag;
  assign io_coef_out_payload_0_9_28_real = int_reg_array_9_28_real;
  assign io_coef_out_payload_0_9_28_imag = int_reg_array_9_28_imag;
  assign io_coef_out_payload_0_9_29_real = int_reg_array_9_29_real;
  assign io_coef_out_payload_0_9_29_imag = int_reg_array_9_29_imag;
  assign io_coef_out_payload_0_9_30_real = int_reg_array_9_30_real;
  assign io_coef_out_payload_0_9_30_imag = int_reg_array_9_30_imag;
  assign io_coef_out_payload_0_9_31_real = int_reg_array_9_31_real;
  assign io_coef_out_payload_0_9_31_imag = int_reg_array_9_31_imag;
  assign io_coef_out_payload_0_9_32_real = int_reg_array_9_32_real;
  assign io_coef_out_payload_0_9_32_imag = int_reg_array_9_32_imag;
  assign io_coef_out_payload_0_9_33_real = int_reg_array_9_33_real;
  assign io_coef_out_payload_0_9_33_imag = int_reg_array_9_33_imag;
  assign io_coef_out_payload_0_9_34_real = int_reg_array_9_34_real;
  assign io_coef_out_payload_0_9_34_imag = int_reg_array_9_34_imag;
  assign io_coef_out_payload_0_9_35_real = int_reg_array_9_35_real;
  assign io_coef_out_payload_0_9_35_imag = int_reg_array_9_35_imag;
  assign io_coef_out_payload_0_9_36_real = int_reg_array_9_36_real;
  assign io_coef_out_payload_0_9_36_imag = int_reg_array_9_36_imag;
  assign io_coef_out_payload_0_9_37_real = int_reg_array_9_37_real;
  assign io_coef_out_payload_0_9_37_imag = int_reg_array_9_37_imag;
  assign io_coef_out_payload_0_9_38_real = int_reg_array_9_38_real;
  assign io_coef_out_payload_0_9_38_imag = int_reg_array_9_38_imag;
  assign io_coef_out_payload_0_9_39_real = int_reg_array_9_39_real;
  assign io_coef_out_payload_0_9_39_imag = int_reg_array_9_39_imag;
  assign io_coef_out_payload_0_9_40_real = int_reg_array_9_40_real;
  assign io_coef_out_payload_0_9_40_imag = int_reg_array_9_40_imag;
  assign io_coef_out_payload_0_9_41_real = int_reg_array_9_41_real;
  assign io_coef_out_payload_0_9_41_imag = int_reg_array_9_41_imag;
  assign io_coef_out_payload_0_9_42_real = int_reg_array_9_42_real;
  assign io_coef_out_payload_0_9_42_imag = int_reg_array_9_42_imag;
  assign io_coef_out_payload_0_9_43_real = int_reg_array_9_43_real;
  assign io_coef_out_payload_0_9_43_imag = int_reg_array_9_43_imag;
  assign io_coef_out_payload_0_9_44_real = int_reg_array_9_44_real;
  assign io_coef_out_payload_0_9_44_imag = int_reg_array_9_44_imag;
  assign io_coef_out_payload_0_9_45_real = int_reg_array_9_45_real;
  assign io_coef_out_payload_0_9_45_imag = int_reg_array_9_45_imag;
  assign io_coef_out_payload_0_9_46_real = int_reg_array_9_46_real;
  assign io_coef_out_payload_0_9_46_imag = int_reg_array_9_46_imag;
  assign io_coef_out_payload_0_9_47_real = int_reg_array_9_47_real;
  assign io_coef_out_payload_0_9_47_imag = int_reg_array_9_47_imag;
  assign io_coef_out_payload_0_9_48_real = int_reg_array_9_48_real;
  assign io_coef_out_payload_0_9_48_imag = int_reg_array_9_48_imag;
  assign io_coef_out_payload_0_9_49_real = int_reg_array_9_49_real;
  assign io_coef_out_payload_0_9_49_imag = int_reg_array_9_49_imag;
  assign io_coef_out_payload_0_10_0_real = int_reg_array_10_0_real;
  assign io_coef_out_payload_0_10_0_imag = int_reg_array_10_0_imag;
  assign io_coef_out_payload_0_10_1_real = int_reg_array_10_1_real;
  assign io_coef_out_payload_0_10_1_imag = int_reg_array_10_1_imag;
  assign io_coef_out_payload_0_10_2_real = int_reg_array_10_2_real;
  assign io_coef_out_payload_0_10_2_imag = int_reg_array_10_2_imag;
  assign io_coef_out_payload_0_10_3_real = int_reg_array_10_3_real;
  assign io_coef_out_payload_0_10_3_imag = int_reg_array_10_3_imag;
  assign io_coef_out_payload_0_10_4_real = int_reg_array_10_4_real;
  assign io_coef_out_payload_0_10_4_imag = int_reg_array_10_4_imag;
  assign io_coef_out_payload_0_10_5_real = int_reg_array_10_5_real;
  assign io_coef_out_payload_0_10_5_imag = int_reg_array_10_5_imag;
  assign io_coef_out_payload_0_10_6_real = int_reg_array_10_6_real;
  assign io_coef_out_payload_0_10_6_imag = int_reg_array_10_6_imag;
  assign io_coef_out_payload_0_10_7_real = int_reg_array_10_7_real;
  assign io_coef_out_payload_0_10_7_imag = int_reg_array_10_7_imag;
  assign io_coef_out_payload_0_10_8_real = int_reg_array_10_8_real;
  assign io_coef_out_payload_0_10_8_imag = int_reg_array_10_8_imag;
  assign io_coef_out_payload_0_10_9_real = int_reg_array_10_9_real;
  assign io_coef_out_payload_0_10_9_imag = int_reg_array_10_9_imag;
  assign io_coef_out_payload_0_10_10_real = int_reg_array_10_10_real;
  assign io_coef_out_payload_0_10_10_imag = int_reg_array_10_10_imag;
  assign io_coef_out_payload_0_10_11_real = int_reg_array_10_11_real;
  assign io_coef_out_payload_0_10_11_imag = int_reg_array_10_11_imag;
  assign io_coef_out_payload_0_10_12_real = int_reg_array_10_12_real;
  assign io_coef_out_payload_0_10_12_imag = int_reg_array_10_12_imag;
  assign io_coef_out_payload_0_10_13_real = int_reg_array_10_13_real;
  assign io_coef_out_payload_0_10_13_imag = int_reg_array_10_13_imag;
  assign io_coef_out_payload_0_10_14_real = int_reg_array_10_14_real;
  assign io_coef_out_payload_0_10_14_imag = int_reg_array_10_14_imag;
  assign io_coef_out_payload_0_10_15_real = int_reg_array_10_15_real;
  assign io_coef_out_payload_0_10_15_imag = int_reg_array_10_15_imag;
  assign io_coef_out_payload_0_10_16_real = int_reg_array_10_16_real;
  assign io_coef_out_payload_0_10_16_imag = int_reg_array_10_16_imag;
  assign io_coef_out_payload_0_10_17_real = int_reg_array_10_17_real;
  assign io_coef_out_payload_0_10_17_imag = int_reg_array_10_17_imag;
  assign io_coef_out_payload_0_10_18_real = int_reg_array_10_18_real;
  assign io_coef_out_payload_0_10_18_imag = int_reg_array_10_18_imag;
  assign io_coef_out_payload_0_10_19_real = int_reg_array_10_19_real;
  assign io_coef_out_payload_0_10_19_imag = int_reg_array_10_19_imag;
  assign io_coef_out_payload_0_10_20_real = int_reg_array_10_20_real;
  assign io_coef_out_payload_0_10_20_imag = int_reg_array_10_20_imag;
  assign io_coef_out_payload_0_10_21_real = int_reg_array_10_21_real;
  assign io_coef_out_payload_0_10_21_imag = int_reg_array_10_21_imag;
  assign io_coef_out_payload_0_10_22_real = int_reg_array_10_22_real;
  assign io_coef_out_payload_0_10_22_imag = int_reg_array_10_22_imag;
  assign io_coef_out_payload_0_10_23_real = int_reg_array_10_23_real;
  assign io_coef_out_payload_0_10_23_imag = int_reg_array_10_23_imag;
  assign io_coef_out_payload_0_10_24_real = int_reg_array_10_24_real;
  assign io_coef_out_payload_0_10_24_imag = int_reg_array_10_24_imag;
  assign io_coef_out_payload_0_10_25_real = int_reg_array_10_25_real;
  assign io_coef_out_payload_0_10_25_imag = int_reg_array_10_25_imag;
  assign io_coef_out_payload_0_10_26_real = int_reg_array_10_26_real;
  assign io_coef_out_payload_0_10_26_imag = int_reg_array_10_26_imag;
  assign io_coef_out_payload_0_10_27_real = int_reg_array_10_27_real;
  assign io_coef_out_payload_0_10_27_imag = int_reg_array_10_27_imag;
  assign io_coef_out_payload_0_10_28_real = int_reg_array_10_28_real;
  assign io_coef_out_payload_0_10_28_imag = int_reg_array_10_28_imag;
  assign io_coef_out_payload_0_10_29_real = int_reg_array_10_29_real;
  assign io_coef_out_payload_0_10_29_imag = int_reg_array_10_29_imag;
  assign io_coef_out_payload_0_10_30_real = int_reg_array_10_30_real;
  assign io_coef_out_payload_0_10_30_imag = int_reg_array_10_30_imag;
  assign io_coef_out_payload_0_10_31_real = int_reg_array_10_31_real;
  assign io_coef_out_payload_0_10_31_imag = int_reg_array_10_31_imag;
  assign io_coef_out_payload_0_10_32_real = int_reg_array_10_32_real;
  assign io_coef_out_payload_0_10_32_imag = int_reg_array_10_32_imag;
  assign io_coef_out_payload_0_10_33_real = int_reg_array_10_33_real;
  assign io_coef_out_payload_0_10_33_imag = int_reg_array_10_33_imag;
  assign io_coef_out_payload_0_10_34_real = int_reg_array_10_34_real;
  assign io_coef_out_payload_0_10_34_imag = int_reg_array_10_34_imag;
  assign io_coef_out_payload_0_10_35_real = int_reg_array_10_35_real;
  assign io_coef_out_payload_0_10_35_imag = int_reg_array_10_35_imag;
  assign io_coef_out_payload_0_10_36_real = int_reg_array_10_36_real;
  assign io_coef_out_payload_0_10_36_imag = int_reg_array_10_36_imag;
  assign io_coef_out_payload_0_10_37_real = int_reg_array_10_37_real;
  assign io_coef_out_payload_0_10_37_imag = int_reg_array_10_37_imag;
  assign io_coef_out_payload_0_10_38_real = int_reg_array_10_38_real;
  assign io_coef_out_payload_0_10_38_imag = int_reg_array_10_38_imag;
  assign io_coef_out_payload_0_10_39_real = int_reg_array_10_39_real;
  assign io_coef_out_payload_0_10_39_imag = int_reg_array_10_39_imag;
  assign io_coef_out_payload_0_10_40_real = int_reg_array_10_40_real;
  assign io_coef_out_payload_0_10_40_imag = int_reg_array_10_40_imag;
  assign io_coef_out_payload_0_10_41_real = int_reg_array_10_41_real;
  assign io_coef_out_payload_0_10_41_imag = int_reg_array_10_41_imag;
  assign io_coef_out_payload_0_10_42_real = int_reg_array_10_42_real;
  assign io_coef_out_payload_0_10_42_imag = int_reg_array_10_42_imag;
  assign io_coef_out_payload_0_10_43_real = int_reg_array_10_43_real;
  assign io_coef_out_payload_0_10_43_imag = int_reg_array_10_43_imag;
  assign io_coef_out_payload_0_10_44_real = int_reg_array_10_44_real;
  assign io_coef_out_payload_0_10_44_imag = int_reg_array_10_44_imag;
  assign io_coef_out_payload_0_10_45_real = int_reg_array_10_45_real;
  assign io_coef_out_payload_0_10_45_imag = int_reg_array_10_45_imag;
  assign io_coef_out_payload_0_10_46_real = int_reg_array_10_46_real;
  assign io_coef_out_payload_0_10_46_imag = int_reg_array_10_46_imag;
  assign io_coef_out_payload_0_10_47_real = int_reg_array_10_47_real;
  assign io_coef_out_payload_0_10_47_imag = int_reg_array_10_47_imag;
  assign io_coef_out_payload_0_10_48_real = int_reg_array_10_48_real;
  assign io_coef_out_payload_0_10_48_imag = int_reg_array_10_48_imag;
  assign io_coef_out_payload_0_10_49_real = int_reg_array_10_49_real;
  assign io_coef_out_payload_0_10_49_imag = int_reg_array_10_49_imag;
  assign io_coef_out_payload_0_11_0_real = int_reg_array_11_0_real;
  assign io_coef_out_payload_0_11_0_imag = int_reg_array_11_0_imag;
  assign io_coef_out_payload_0_11_1_real = int_reg_array_11_1_real;
  assign io_coef_out_payload_0_11_1_imag = int_reg_array_11_1_imag;
  assign io_coef_out_payload_0_11_2_real = int_reg_array_11_2_real;
  assign io_coef_out_payload_0_11_2_imag = int_reg_array_11_2_imag;
  assign io_coef_out_payload_0_11_3_real = int_reg_array_11_3_real;
  assign io_coef_out_payload_0_11_3_imag = int_reg_array_11_3_imag;
  assign io_coef_out_payload_0_11_4_real = int_reg_array_11_4_real;
  assign io_coef_out_payload_0_11_4_imag = int_reg_array_11_4_imag;
  assign io_coef_out_payload_0_11_5_real = int_reg_array_11_5_real;
  assign io_coef_out_payload_0_11_5_imag = int_reg_array_11_5_imag;
  assign io_coef_out_payload_0_11_6_real = int_reg_array_11_6_real;
  assign io_coef_out_payload_0_11_6_imag = int_reg_array_11_6_imag;
  assign io_coef_out_payload_0_11_7_real = int_reg_array_11_7_real;
  assign io_coef_out_payload_0_11_7_imag = int_reg_array_11_7_imag;
  assign io_coef_out_payload_0_11_8_real = int_reg_array_11_8_real;
  assign io_coef_out_payload_0_11_8_imag = int_reg_array_11_8_imag;
  assign io_coef_out_payload_0_11_9_real = int_reg_array_11_9_real;
  assign io_coef_out_payload_0_11_9_imag = int_reg_array_11_9_imag;
  assign io_coef_out_payload_0_11_10_real = int_reg_array_11_10_real;
  assign io_coef_out_payload_0_11_10_imag = int_reg_array_11_10_imag;
  assign io_coef_out_payload_0_11_11_real = int_reg_array_11_11_real;
  assign io_coef_out_payload_0_11_11_imag = int_reg_array_11_11_imag;
  assign io_coef_out_payload_0_11_12_real = int_reg_array_11_12_real;
  assign io_coef_out_payload_0_11_12_imag = int_reg_array_11_12_imag;
  assign io_coef_out_payload_0_11_13_real = int_reg_array_11_13_real;
  assign io_coef_out_payload_0_11_13_imag = int_reg_array_11_13_imag;
  assign io_coef_out_payload_0_11_14_real = int_reg_array_11_14_real;
  assign io_coef_out_payload_0_11_14_imag = int_reg_array_11_14_imag;
  assign io_coef_out_payload_0_11_15_real = int_reg_array_11_15_real;
  assign io_coef_out_payload_0_11_15_imag = int_reg_array_11_15_imag;
  assign io_coef_out_payload_0_11_16_real = int_reg_array_11_16_real;
  assign io_coef_out_payload_0_11_16_imag = int_reg_array_11_16_imag;
  assign io_coef_out_payload_0_11_17_real = int_reg_array_11_17_real;
  assign io_coef_out_payload_0_11_17_imag = int_reg_array_11_17_imag;
  assign io_coef_out_payload_0_11_18_real = int_reg_array_11_18_real;
  assign io_coef_out_payload_0_11_18_imag = int_reg_array_11_18_imag;
  assign io_coef_out_payload_0_11_19_real = int_reg_array_11_19_real;
  assign io_coef_out_payload_0_11_19_imag = int_reg_array_11_19_imag;
  assign io_coef_out_payload_0_11_20_real = int_reg_array_11_20_real;
  assign io_coef_out_payload_0_11_20_imag = int_reg_array_11_20_imag;
  assign io_coef_out_payload_0_11_21_real = int_reg_array_11_21_real;
  assign io_coef_out_payload_0_11_21_imag = int_reg_array_11_21_imag;
  assign io_coef_out_payload_0_11_22_real = int_reg_array_11_22_real;
  assign io_coef_out_payload_0_11_22_imag = int_reg_array_11_22_imag;
  assign io_coef_out_payload_0_11_23_real = int_reg_array_11_23_real;
  assign io_coef_out_payload_0_11_23_imag = int_reg_array_11_23_imag;
  assign io_coef_out_payload_0_11_24_real = int_reg_array_11_24_real;
  assign io_coef_out_payload_0_11_24_imag = int_reg_array_11_24_imag;
  assign io_coef_out_payload_0_11_25_real = int_reg_array_11_25_real;
  assign io_coef_out_payload_0_11_25_imag = int_reg_array_11_25_imag;
  assign io_coef_out_payload_0_11_26_real = int_reg_array_11_26_real;
  assign io_coef_out_payload_0_11_26_imag = int_reg_array_11_26_imag;
  assign io_coef_out_payload_0_11_27_real = int_reg_array_11_27_real;
  assign io_coef_out_payload_0_11_27_imag = int_reg_array_11_27_imag;
  assign io_coef_out_payload_0_11_28_real = int_reg_array_11_28_real;
  assign io_coef_out_payload_0_11_28_imag = int_reg_array_11_28_imag;
  assign io_coef_out_payload_0_11_29_real = int_reg_array_11_29_real;
  assign io_coef_out_payload_0_11_29_imag = int_reg_array_11_29_imag;
  assign io_coef_out_payload_0_11_30_real = int_reg_array_11_30_real;
  assign io_coef_out_payload_0_11_30_imag = int_reg_array_11_30_imag;
  assign io_coef_out_payload_0_11_31_real = int_reg_array_11_31_real;
  assign io_coef_out_payload_0_11_31_imag = int_reg_array_11_31_imag;
  assign io_coef_out_payload_0_11_32_real = int_reg_array_11_32_real;
  assign io_coef_out_payload_0_11_32_imag = int_reg_array_11_32_imag;
  assign io_coef_out_payload_0_11_33_real = int_reg_array_11_33_real;
  assign io_coef_out_payload_0_11_33_imag = int_reg_array_11_33_imag;
  assign io_coef_out_payload_0_11_34_real = int_reg_array_11_34_real;
  assign io_coef_out_payload_0_11_34_imag = int_reg_array_11_34_imag;
  assign io_coef_out_payload_0_11_35_real = int_reg_array_11_35_real;
  assign io_coef_out_payload_0_11_35_imag = int_reg_array_11_35_imag;
  assign io_coef_out_payload_0_11_36_real = int_reg_array_11_36_real;
  assign io_coef_out_payload_0_11_36_imag = int_reg_array_11_36_imag;
  assign io_coef_out_payload_0_11_37_real = int_reg_array_11_37_real;
  assign io_coef_out_payload_0_11_37_imag = int_reg_array_11_37_imag;
  assign io_coef_out_payload_0_11_38_real = int_reg_array_11_38_real;
  assign io_coef_out_payload_0_11_38_imag = int_reg_array_11_38_imag;
  assign io_coef_out_payload_0_11_39_real = int_reg_array_11_39_real;
  assign io_coef_out_payload_0_11_39_imag = int_reg_array_11_39_imag;
  assign io_coef_out_payload_0_11_40_real = int_reg_array_11_40_real;
  assign io_coef_out_payload_0_11_40_imag = int_reg_array_11_40_imag;
  assign io_coef_out_payload_0_11_41_real = int_reg_array_11_41_real;
  assign io_coef_out_payload_0_11_41_imag = int_reg_array_11_41_imag;
  assign io_coef_out_payload_0_11_42_real = int_reg_array_11_42_real;
  assign io_coef_out_payload_0_11_42_imag = int_reg_array_11_42_imag;
  assign io_coef_out_payload_0_11_43_real = int_reg_array_11_43_real;
  assign io_coef_out_payload_0_11_43_imag = int_reg_array_11_43_imag;
  assign io_coef_out_payload_0_11_44_real = int_reg_array_11_44_real;
  assign io_coef_out_payload_0_11_44_imag = int_reg_array_11_44_imag;
  assign io_coef_out_payload_0_11_45_real = int_reg_array_11_45_real;
  assign io_coef_out_payload_0_11_45_imag = int_reg_array_11_45_imag;
  assign io_coef_out_payload_0_11_46_real = int_reg_array_11_46_real;
  assign io_coef_out_payload_0_11_46_imag = int_reg_array_11_46_imag;
  assign io_coef_out_payload_0_11_47_real = int_reg_array_11_47_real;
  assign io_coef_out_payload_0_11_47_imag = int_reg_array_11_47_imag;
  assign io_coef_out_payload_0_11_48_real = int_reg_array_11_48_real;
  assign io_coef_out_payload_0_11_48_imag = int_reg_array_11_48_imag;
  assign io_coef_out_payload_0_11_49_real = int_reg_array_11_49_real;
  assign io_coef_out_payload_0_11_49_imag = int_reg_array_11_49_imag;
  assign io_coef_out_payload_0_12_0_real = int_reg_array_12_0_real;
  assign io_coef_out_payload_0_12_0_imag = int_reg_array_12_0_imag;
  assign io_coef_out_payload_0_12_1_real = int_reg_array_12_1_real;
  assign io_coef_out_payload_0_12_1_imag = int_reg_array_12_1_imag;
  assign io_coef_out_payload_0_12_2_real = int_reg_array_12_2_real;
  assign io_coef_out_payload_0_12_2_imag = int_reg_array_12_2_imag;
  assign io_coef_out_payload_0_12_3_real = int_reg_array_12_3_real;
  assign io_coef_out_payload_0_12_3_imag = int_reg_array_12_3_imag;
  assign io_coef_out_payload_0_12_4_real = int_reg_array_12_4_real;
  assign io_coef_out_payload_0_12_4_imag = int_reg_array_12_4_imag;
  assign io_coef_out_payload_0_12_5_real = int_reg_array_12_5_real;
  assign io_coef_out_payload_0_12_5_imag = int_reg_array_12_5_imag;
  assign io_coef_out_payload_0_12_6_real = int_reg_array_12_6_real;
  assign io_coef_out_payload_0_12_6_imag = int_reg_array_12_6_imag;
  assign io_coef_out_payload_0_12_7_real = int_reg_array_12_7_real;
  assign io_coef_out_payload_0_12_7_imag = int_reg_array_12_7_imag;
  assign io_coef_out_payload_0_12_8_real = int_reg_array_12_8_real;
  assign io_coef_out_payload_0_12_8_imag = int_reg_array_12_8_imag;
  assign io_coef_out_payload_0_12_9_real = int_reg_array_12_9_real;
  assign io_coef_out_payload_0_12_9_imag = int_reg_array_12_9_imag;
  assign io_coef_out_payload_0_12_10_real = int_reg_array_12_10_real;
  assign io_coef_out_payload_0_12_10_imag = int_reg_array_12_10_imag;
  assign io_coef_out_payload_0_12_11_real = int_reg_array_12_11_real;
  assign io_coef_out_payload_0_12_11_imag = int_reg_array_12_11_imag;
  assign io_coef_out_payload_0_12_12_real = int_reg_array_12_12_real;
  assign io_coef_out_payload_0_12_12_imag = int_reg_array_12_12_imag;
  assign io_coef_out_payload_0_12_13_real = int_reg_array_12_13_real;
  assign io_coef_out_payload_0_12_13_imag = int_reg_array_12_13_imag;
  assign io_coef_out_payload_0_12_14_real = int_reg_array_12_14_real;
  assign io_coef_out_payload_0_12_14_imag = int_reg_array_12_14_imag;
  assign io_coef_out_payload_0_12_15_real = int_reg_array_12_15_real;
  assign io_coef_out_payload_0_12_15_imag = int_reg_array_12_15_imag;
  assign io_coef_out_payload_0_12_16_real = int_reg_array_12_16_real;
  assign io_coef_out_payload_0_12_16_imag = int_reg_array_12_16_imag;
  assign io_coef_out_payload_0_12_17_real = int_reg_array_12_17_real;
  assign io_coef_out_payload_0_12_17_imag = int_reg_array_12_17_imag;
  assign io_coef_out_payload_0_12_18_real = int_reg_array_12_18_real;
  assign io_coef_out_payload_0_12_18_imag = int_reg_array_12_18_imag;
  assign io_coef_out_payload_0_12_19_real = int_reg_array_12_19_real;
  assign io_coef_out_payload_0_12_19_imag = int_reg_array_12_19_imag;
  assign io_coef_out_payload_0_12_20_real = int_reg_array_12_20_real;
  assign io_coef_out_payload_0_12_20_imag = int_reg_array_12_20_imag;
  assign io_coef_out_payload_0_12_21_real = int_reg_array_12_21_real;
  assign io_coef_out_payload_0_12_21_imag = int_reg_array_12_21_imag;
  assign io_coef_out_payload_0_12_22_real = int_reg_array_12_22_real;
  assign io_coef_out_payload_0_12_22_imag = int_reg_array_12_22_imag;
  assign io_coef_out_payload_0_12_23_real = int_reg_array_12_23_real;
  assign io_coef_out_payload_0_12_23_imag = int_reg_array_12_23_imag;
  assign io_coef_out_payload_0_12_24_real = int_reg_array_12_24_real;
  assign io_coef_out_payload_0_12_24_imag = int_reg_array_12_24_imag;
  assign io_coef_out_payload_0_12_25_real = int_reg_array_12_25_real;
  assign io_coef_out_payload_0_12_25_imag = int_reg_array_12_25_imag;
  assign io_coef_out_payload_0_12_26_real = int_reg_array_12_26_real;
  assign io_coef_out_payload_0_12_26_imag = int_reg_array_12_26_imag;
  assign io_coef_out_payload_0_12_27_real = int_reg_array_12_27_real;
  assign io_coef_out_payload_0_12_27_imag = int_reg_array_12_27_imag;
  assign io_coef_out_payload_0_12_28_real = int_reg_array_12_28_real;
  assign io_coef_out_payload_0_12_28_imag = int_reg_array_12_28_imag;
  assign io_coef_out_payload_0_12_29_real = int_reg_array_12_29_real;
  assign io_coef_out_payload_0_12_29_imag = int_reg_array_12_29_imag;
  assign io_coef_out_payload_0_12_30_real = int_reg_array_12_30_real;
  assign io_coef_out_payload_0_12_30_imag = int_reg_array_12_30_imag;
  assign io_coef_out_payload_0_12_31_real = int_reg_array_12_31_real;
  assign io_coef_out_payload_0_12_31_imag = int_reg_array_12_31_imag;
  assign io_coef_out_payload_0_12_32_real = int_reg_array_12_32_real;
  assign io_coef_out_payload_0_12_32_imag = int_reg_array_12_32_imag;
  assign io_coef_out_payload_0_12_33_real = int_reg_array_12_33_real;
  assign io_coef_out_payload_0_12_33_imag = int_reg_array_12_33_imag;
  assign io_coef_out_payload_0_12_34_real = int_reg_array_12_34_real;
  assign io_coef_out_payload_0_12_34_imag = int_reg_array_12_34_imag;
  assign io_coef_out_payload_0_12_35_real = int_reg_array_12_35_real;
  assign io_coef_out_payload_0_12_35_imag = int_reg_array_12_35_imag;
  assign io_coef_out_payload_0_12_36_real = int_reg_array_12_36_real;
  assign io_coef_out_payload_0_12_36_imag = int_reg_array_12_36_imag;
  assign io_coef_out_payload_0_12_37_real = int_reg_array_12_37_real;
  assign io_coef_out_payload_0_12_37_imag = int_reg_array_12_37_imag;
  assign io_coef_out_payload_0_12_38_real = int_reg_array_12_38_real;
  assign io_coef_out_payload_0_12_38_imag = int_reg_array_12_38_imag;
  assign io_coef_out_payload_0_12_39_real = int_reg_array_12_39_real;
  assign io_coef_out_payload_0_12_39_imag = int_reg_array_12_39_imag;
  assign io_coef_out_payload_0_12_40_real = int_reg_array_12_40_real;
  assign io_coef_out_payload_0_12_40_imag = int_reg_array_12_40_imag;
  assign io_coef_out_payload_0_12_41_real = int_reg_array_12_41_real;
  assign io_coef_out_payload_0_12_41_imag = int_reg_array_12_41_imag;
  assign io_coef_out_payload_0_12_42_real = int_reg_array_12_42_real;
  assign io_coef_out_payload_0_12_42_imag = int_reg_array_12_42_imag;
  assign io_coef_out_payload_0_12_43_real = int_reg_array_12_43_real;
  assign io_coef_out_payload_0_12_43_imag = int_reg_array_12_43_imag;
  assign io_coef_out_payload_0_12_44_real = int_reg_array_12_44_real;
  assign io_coef_out_payload_0_12_44_imag = int_reg_array_12_44_imag;
  assign io_coef_out_payload_0_12_45_real = int_reg_array_12_45_real;
  assign io_coef_out_payload_0_12_45_imag = int_reg_array_12_45_imag;
  assign io_coef_out_payload_0_12_46_real = int_reg_array_12_46_real;
  assign io_coef_out_payload_0_12_46_imag = int_reg_array_12_46_imag;
  assign io_coef_out_payload_0_12_47_real = int_reg_array_12_47_real;
  assign io_coef_out_payload_0_12_47_imag = int_reg_array_12_47_imag;
  assign io_coef_out_payload_0_12_48_real = int_reg_array_12_48_real;
  assign io_coef_out_payload_0_12_48_imag = int_reg_array_12_48_imag;
  assign io_coef_out_payload_0_12_49_real = int_reg_array_12_49_real;
  assign io_coef_out_payload_0_12_49_imag = int_reg_array_12_49_imag;
  assign io_coef_out_payload_0_13_0_real = int_reg_array_13_0_real;
  assign io_coef_out_payload_0_13_0_imag = int_reg_array_13_0_imag;
  assign io_coef_out_payload_0_13_1_real = int_reg_array_13_1_real;
  assign io_coef_out_payload_0_13_1_imag = int_reg_array_13_1_imag;
  assign io_coef_out_payload_0_13_2_real = int_reg_array_13_2_real;
  assign io_coef_out_payload_0_13_2_imag = int_reg_array_13_2_imag;
  assign io_coef_out_payload_0_13_3_real = int_reg_array_13_3_real;
  assign io_coef_out_payload_0_13_3_imag = int_reg_array_13_3_imag;
  assign io_coef_out_payload_0_13_4_real = int_reg_array_13_4_real;
  assign io_coef_out_payload_0_13_4_imag = int_reg_array_13_4_imag;
  assign io_coef_out_payload_0_13_5_real = int_reg_array_13_5_real;
  assign io_coef_out_payload_0_13_5_imag = int_reg_array_13_5_imag;
  assign io_coef_out_payload_0_13_6_real = int_reg_array_13_6_real;
  assign io_coef_out_payload_0_13_6_imag = int_reg_array_13_6_imag;
  assign io_coef_out_payload_0_13_7_real = int_reg_array_13_7_real;
  assign io_coef_out_payload_0_13_7_imag = int_reg_array_13_7_imag;
  assign io_coef_out_payload_0_13_8_real = int_reg_array_13_8_real;
  assign io_coef_out_payload_0_13_8_imag = int_reg_array_13_8_imag;
  assign io_coef_out_payload_0_13_9_real = int_reg_array_13_9_real;
  assign io_coef_out_payload_0_13_9_imag = int_reg_array_13_9_imag;
  assign io_coef_out_payload_0_13_10_real = int_reg_array_13_10_real;
  assign io_coef_out_payload_0_13_10_imag = int_reg_array_13_10_imag;
  assign io_coef_out_payload_0_13_11_real = int_reg_array_13_11_real;
  assign io_coef_out_payload_0_13_11_imag = int_reg_array_13_11_imag;
  assign io_coef_out_payload_0_13_12_real = int_reg_array_13_12_real;
  assign io_coef_out_payload_0_13_12_imag = int_reg_array_13_12_imag;
  assign io_coef_out_payload_0_13_13_real = int_reg_array_13_13_real;
  assign io_coef_out_payload_0_13_13_imag = int_reg_array_13_13_imag;
  assign io_coef_out_payload_0_13_14_real = int_reg_array_13_14_real;
  assign io_coef_out_payload_0_13_14_imag = int_reg_array_13_14_imag;
  assign io_coef_out_payload_0_13_15_real = int_reg_array_13_15_real;
  assign io_coef_out_payload_0_13_15_imag = int_reg_array_13_15_imag;
  assign io_coef_out_payload_0_13_16_real = int_reg_array_13_16_real;
  assign io_coef_out_payload_0_13_16_imag = int_reg_array_13_16_imag;
  assign io_coef_out_payload_0_13_17_real = int_reg_array_13_17_real;
  assign io_coef_out_payload_0_13_17_imag = int_reg_array_13_17_imag;
  assign io_coef_out_payload_0_13_18_real = int_reg_array_13_18_real;
  assign io_coef_out_payload_0_13_18_imag = int_reg_array_13_18_imag;
  assign io_coef_out_payload_0_13_19_real = int_reg_array_13_19_real;
  assign io_coef_out_payload_0_13_19_imag = int_reg_array_13_19_imag;
  assign io_coef_out_payload_0_13_20_real = int_reg_array_13_20_real;
  assign io_coef_out_payload_0_13_20_imag = int_reg_array_13_20_imag;
  assign io_coef_out_payload_0_13_21_real = int_reg_array_13_21_real;
  assign io_coef_out_payload_0_13_21_imag = int_reg_array_13_21_imag;
  assign io_coef_out_payload_0_13_22_real = int_reg_array_13_22_real;
  assign io_coef_out_payload_0_13_22_imag = int_reg_array_13_22_imag;
  assign io_coef_out_payload_0_13_23_real = int_reg_array_13_23_real;
  assign io_coef_out_payload_0_13_23_imag = int_reg_array_13_23_imag;
  assign io_coef_out_payload_0_13_24_real = int_reg_array_13_24_real;
  assign io_coef_out_payload_0_13_24_imag = int_reg_array_13_24_imag;
  assign io_coef_out_payload_0_13_25_real = int_reg_array_13_25_real;
  assign io_coef_out_payload_0_13_25_imag = int_reg_array_13_25_imag;
  assign io_coef_out_payload_0_13_26_real = int_reg_array_13_26_real;
  assign io_coef_out_payload_0_13_26_imag = int_reg_array_13_26_imag;
  assign io_coef_out_payload_0_13_27_real = int_reg_array_13_27_real;
  assign io_coef_out_payload_0_13_27_imag = int_reg_array_13_27_imag;
  assign io_coef_out_payload_0_13_28_real = int_reg_array_13_28_real;
  assign io_coef_out_payload_0_13_28_imag = int_reg_array_13_28_imag;
  assign io_coef_out_payload_0_13_29_real = int_reg_array_13_29_real;
  assign io_coef_out_payload_0_13_29_imag = int_reg_array_13_29_imag;
  assign io_coef_out_payload_0_13_30_real = int_reg_array_13_30_real;
  assign io_coef_out_payload_0_13_30_imag = int_reg_array_13_30_imag;
  assign io_coef_out_payload_0_13_31_real = int_reg_array_13_31_real;
  assign io_coef_out_payload_0_13_31_imag = int_reg_array_13_31_imag;
  assign io_coef_out_payload_0_13_32_real = int_reg_array_13_32_real;
  assign io_coef_out_payload_0_13_32_imag = int_reg_array_13_32_imag;
  assign io_coef_out_payload_0_13_33_real = int_reg_array_13_33_real;
  assign io_coef_out_payload_0_13_33_imag = int_reg_array_13_33_imag;
  assign io_coef_out_payload_0_13_34_real = int_reg_array_13_34_real;
  assign io_coef_out_payload_0_13_34_imag = int_reg_array_13_34_imag;
  assign io_coef_out_payload_0_13_35_real = int_reg_array_13_35_real;
  assign io_coef_out_payload_0_13_35_imag = int_reg_array_13_35_imag;
  assign io_coef_out_payload_0_13_36_real = int_reg_array_13_36_real;
  assign io_coef_out_payload_0_13_36_imag = int_reg_array_13_36_imag;
  assign io_coef_out_payload_0_13_37_real = int_reg_array_13_37_real;
  assign io_coef_out_payload_0_13_37_imag = int_reg_array_13_37_imag;
  assign io_coef_out_payload_0_13_38_real = int_reg_array_13_38_real;
  assign io_coef_out_payload_0_13_38_imag = int_reg_array_13_38_imag;
  assign io_coef_out_payload_0_13_39_real = int_reg_array_13_39_real;
  assign io_coef_out_payload_0_13_39_imag = int_reg_array_13_39_imag;
  assign io_coef_out_payload_0_13_40_real = int_reg_array_13_40_real;
  assign io_coef_out_payload_0_13_40_imag = int_reg_array_13_40_imag;
  assign io_coef_out_payload_0_13_41_real = int_reg_array_13_41_real;
  assign io_coef_out_payload_0_13_41_imag = int_reg_array_13_41_imag;
  assign io_coef_out_payload_0_13_42_real = int_reg_array_13_42_real;
  assign io_coef_out_payload_0_13_42_imag = int_reg_array_13_42_imag;
  assign io_coef_out_payload_0_13_43_real = int_reg_array_13_43_real;
  assign io_coef_out_payload_0_13_43_imag = int_reg_array_13_43_imag;
  assign io_coef_out_payload_0_13_44_real = int_reg_array_13_44_real;
  assign io_coef_out_payload_0_13_44_imag = int_reg_array_13_44_imag;
  assign io_coef_out_payload_0_13_45_real = int_reg_array_13_45_real;
  assign io_coef_out_payload_0_13_45_imag = int_reg_array_13_45_imag;
  assign io_coef_out_payload_0_13_46_real = int_reg_array_13_46_real;
  assign io_coef_out_payload_0_13_46_imag = int_reg_array_13_46_imag;
  assign io_coef_out_payload_0_13_47_real = int_reg_array_13_47_real;
  assign io_coef_out_payload_0_13_47_imag = int_reg_array_13_47_imag;
  assign io_coef_out_payload_0_13_48_real = int_reg_array_13_48_real;
  assign io_coef_out_payload_0_13_48_imag = int_reg_array_13_48_imag;
  assign io_coef_out_payload_0_13_49_real = int_reg_array_13_49_real;
  assign io_coef_out_payload_0_13_49_imag = int_reg_array_13_49_imag;
  assign io_coef_out_payload_0_14_0_real = int_reg_array_14_0_real;
  assign io_coef_out_payload_0_14_0_imag = int_reg_array_14_0_imag;
  assign io_coef_out_payload_0_14_1_real = int_reg_array_14_1_real;
  assign io_coef_out_payload_0_14_1_imag = int_reg_array_14_1_imag;
  assign io_coef_out_payload_0_14_2_real = int_reg_array_14_2_real;
  assign io_coef_out_payload_0_14_2_imag = int_reg_array_14_2_imag;
  assign io_coef_out_payload_0_14_3_real = int_reg_array_14_3_real;
  assign io_coef_out_payload_0_14_3_imag = int_reg_array_14_3_imag;
  assign io_coef_out_payload_0_14_4_real = int_reg_array_14_4_real;
  assign io_coef_out_payload_0_14_4_imag = int_reg_array_14_4_imag;
  assign io_coef_out_payload_0_14_5_real = int_reg_array_14_5_real;
  assign io_coef_out_payload_0_14_5_imag = int_reg_array_14_5_imag;
  assign io_coef_out_payload_0_14_6_real = int_reg_array_14_6_real;
  assign io_coef_out_payload_0_14_6_imag = int_reg_array_14_6_imag;
  assign io_coef_out_payload_0_14_7_real = int_reg_array_14_7_real;
  assign io_coef_out_payload_0_14_7_imag = int_reg_array_14_7_imag;
  assign io_coef_out_payload_0_14_8_real = int_reg_array_14_8_real;
  assign io_coef_out_payload_0_14_8_imag = int_reg_array_14_8_imag;
  assign io_coef_out_payload_0_14_9_real = int_reg_array_14_9_real;
  assign io_coef_out_payload_0_14_9_imag = int_reg_array_14_9_imag;
  assign io_coef_out_payload_0_14_10_real = int_reg_array_14_10_real;
  assign io_coef_out_payload_0_14_10_imag = int_reg_array_14_10_imag;
  assign io_coef_out_payload_0_14_11_real = int_reg_array_14_11_real;
  assign io_coef_out_payload_0_14_11_imag = int_reg_array_14_11_imag;
  assign io_coef_out_payload_0_14_12_real = int_reg_array_14_12_real;
  assign io_coef_out_payload_0_14_12_imag = int_reg_array_14_12_imag;
  assign io_coef_out_payload_0_14_13_real = int_reg_array_14_13_real;
  assign io_coef_out_payload_0_14_13_imag = int_reg_array_14_13_imag;
  assign io_coef_out_payload_0_14_14_real = int_reg_array_14_14_real;
  assign io_coef_out_payload_0_14_14_imag = int_reg_array_14_14_imag;
  assign io_coef_out_payload_0_14_15_real = int_reg_array_14_15_real;
  assign io_coef_out_payload_0_14_15_imag = int_reg_array_14_15_imag;
  assign io_coef_out_payload_0_14_16_real = int_reg_array_14_16_real;
  assign io_coef_out_payload_0_14_16_imag = int_reg_array_14_16_imag;
  assign io_coef_out_payload_0_14_17_real = int_reg_array_14_17_real;
  assign io_coef_out_payload_0_14_17_imag = int_reg_array_14_17_imag;
  assign io_coef_out_payload_0_14_18_real = int_reg_array_14_18_real;
  assign io_coef_out_payload_0_14_18_imag = int_reg_array_14_18_imag;
  assign io_coef_out_payload_0_14_19_real = int_reg_array_14_19_real;
  assign io_coef_out_payload_0_14_19_imag = int_reg_array_14_19_imag;
  assign io_coef_out_payload_0_14_20_real = int_reg_array_14_20_real;
  assign io_coef_out_payload_0_14_20_imag = int_reg_array_14_20_imag;
  assign io_coef_out_payload_0_14_21_real = int_reg_array_14_21_real;
  assign io_coef_out_payload_0_14_21_imag = int_reg_array_14_21_imag;
  assign io_coef_out_payload_0_14_22_real = int_reg_array_14_22_real;
  assign io_coef_out_payload_0_14_22_imag = int_reg_array_14_22_imag;
  assign io_coef_out_payload_0_14_23_real = int_reg_array_14_23_real;
  assign io_coef_out_payload_0_14_23_imag = int_reg_array_14_23_imag;
  assign io_coef_out_payload_0_14_24_real = int_reg_array_14_24_real;
  assign io_coef_out_payload_0_14_24_imag = int_reg_array_14_24_imag;
  assign io_coef_out_payload_0_14_25_real = int_reg_array_14_25_real;
  assign io_coef_out_payload_0_14_25_imag = int_reg_array_14_25_imag;
  assign io_coef_out_payload_0_14_26_real = int_reg_array_14_26_real;
  assign io_coef_out_payload_0_14_26_imag = int_reg_array_14_26_imag;
  assign io_coef_out_payload_0_14_27_real = int_reg_array_14_27_real;
  assign io_coef_out_payload_0_14_27_imag = int_reg_array_14_27_imag;
  assign io_coef_out_payload_0_14_28_real = int_reg_array_14_28_real;
  assign io_coef_out_payload_0_14_28_imag = int_reg_array_14_28_imag;
  assign io_coef_out_payload_0_14_29_real = int_reg_array_14_29_real;
  assign io_coef_out_payload_0_14_29_imag = int_reg_array_14_29_imag;
  assign io_coef_out_payload_0_14_30_real = int_reg_array_14_30_real;
  assign io_coef_out_payload_0_14_30_imag = int_reg_array_14_30_imag;
  assign io_coef_out_payload_0_14_31_real = int_reg_array_14_31_real;
  assign io_coef_out_payload_0_14_31_imag = int_reg_array_14_31_imag;
  assign io_coef_out_payload_0_14_32_real = int_reg_array_14_32_real;
  assign io_coef_out_payload_0_14_32_imag = int_reg_array_14_32_imag;
  assign io_coef_out_payload_0_14_33_real = int_reg_array_14_33_real;
  assign io_coef_out_payload_0_14_33_imag = int_reg_array_14_33_imag;
  assign io_coef_out_payload_0_14_34_real = int_reg_array_14_34_real;
  assign io_coef_out_payload_0_14_34_imag = int_reg_array_14_34_imag;
  assign io_coef_out_payload_0_14_35_real = int_reg_array_14_35_real;
  assign io_coef_out_payload_0_14_35_imag = int_reg_array_14_35_imag;
  assign io_coef_out_payload_0_14_36_real = int_reg_array_14_36_real;
  assign io_coef_out_payload_0_14_36_imag = int_reg_array_14_36_imag;
  assign io_coef_out_payload_0_14_37_real = int_reg_array_14_37_real;
  assign io_coef_out_payload_0_14_37_imag = int_reg_array_14_37_imag;
  assign io_coef_out_payload_0_14_38_real = int_reg_array_14_38_real;
  assign io_coef_out_payload_0_14_38_imag = int_reg_array_14_38_imag;
  assign io_coef_out_payload_0_14_39_real = int_reg_array_14_39_real;
  assign io_coef_out_payload_0_14_39_imag = int_reg_array_14_39_imag;
  assign io_coef_out_payload_0_14_40_real = int_reg_array_14_40_real;
  assign io_coef_out_payload_0_14_40_imag = int_reg_array_14_40_imag;
  assign io_coef_out_payload_0_14_41_real = int_reg_array_14_41_real;
  assign io_coef_out_payload_0_14_41_imag = int_reg_array_14_41_imag;
  assign io_coef_out_payload_0_14_42_real = int_reg_array_14_42_real;
  assign io_coef_out_payload_0_14_42_imag = int_reg_array_14_42_imag;
  assign io_coef_out_payload_0_14_43_real = int_reg_array_14_43_real;
  assign io_coef_out_payload_0_14_43_imag = int_reg_array_14_43_imag;
  assign io_coef_out_payload_0_14_44_real = int_reg_array_14_44_real;
  assign io_coef_out_payload_0_14_44_imag = int_reg_array_14_44_imag;
  assign io_coef_out_payload_0_14_45_real = int_reg_array_14_45_real;
  assign io_coef_out_payload_0_14_45_imag = int_reg_array_14_45_imag;
  assign io_coef_out_payload_0_14_46_real = int_reg_array_14_46_real;
  assign io_coef_out_payload_0_14_46_imag = int_reg_array_14_46_imag;
  assign io_coef_out_payload_0_14_47_real = int_reg_array_14_47_real;
  assign io_coef_out_payload_0_14_47_imag = int_reg_array_14_47_imag;
  assign io_coef_out_payload_0_14_48_real = int_reg_array_14_48_real;
  assign io_coef_out_payload_0_14_48_imag = int_reg_array_14_48_imag;
  assign io_coef_out_payload_0_14_49_real = int_reg_array_14_49_real;
  assign io_coef_out_payload_0_14_49_imag = int_reg_array_14_49_imag;
  assign io_coef_out_payload_0_15_0_real = int_reg_array_15_0_real;
  assign io_coef_out_payload_0_15_0_imag = int_reg_array_15_0_imag;
  assign io_coef_out_payload_0_15_1_real = int_reg_array_15_1_real;
  assign io_coef_out_payload_0_15_1_imag = int_reg_array_15_1_imag;
  assign io_coef_out_payload_0_15_2_real = int_reg_array_15_2_real;
  assign io_coef_out_payload_0_15_2_imag = int_reg_array_15_2_imag;
  assign io_coef_out_payload_0_15_3_real = int_reg_array_15_3_real;
  assign io_coef_out_payload_0_15_3_imag = int_reg_array_15_3_imag;
  assign io_coef_out_payload_0_15_4_real = int_reg_array_15_4_real;
  assign io_coef_out_payload_0_15_4_imag = int_reg_array_15_4_imag;
  assign io_coef_out_payload_0_15_5_real = int_reg_array_15_5_real;
  assign io_coef_out_payload_0_15_5_imag = int_reg_array_15_5_imag;
  assign io_coef_out_payload_0_15_6_real = int_reg_array_15_6_real;
  assign io_coef_out_payload_0_15_6_imag = int_reg_array_15_6_imag;
  assign io_coef_out_payload_0_15_7_real = int_reg_array_15_7_real;
  assign io_coef_out_payload_0_15_7_imag = int_reg_array_15_7_imag;
  assign io_coef_out_payload_0_15_8_real = int_reg_array_15_8_real;
  assign io_coef_out_payload_0_15_8_imag = int_reg_array_15_8_imag;
  assign io_coef_out_payload_0_15_9_real = int_reg_array_15_9_real;
  assign io_coef_out_payload_0_15_9_imag = int_reg_array_15_9_imag;
  assign io_coef_out_payload_0_15_10_real = int_reg_array_15_10_real;
  assign io_coef_out_payload_0_15_10_imag = int_reg_array_15_10_imag;
  assign io_coef_out_payload_0_15_11_real = int_reg_array_15_11_real;
  assign io_coef_out_payload_0_15_11_imag = int_reg_array_15_11_imag;
  assign io_coef_out_payload_0_15_12_real = int_reg_array_15_12_real;
  assign io_coef_out_payload_0_15_12_imag = int_reg_array_15_12_imag;
  assign io_coef_out_payload_0_15_13_real = int_reg_array_15_13_real;
  assign io_coef_out_payload_0_15_13_imag = int_reg_array_15_13_imag;
  assign io_coef_out_payload_0_15_14_real = int_reg_array_15_14_real;
  assign io_coef_out_payload_0_15_14_imag = int_reg_array_15_14_imag;
  assign io_coef_out_payload_0_15_15_real = int_reg_array_15_15_real;
  assign io_coef_out_payload_0_15_15_imag = int_reg_array_15_15_imag;
  assign io_coef_out_payload_0_15_16_real = int_reg_array_15_16_real;
  assign io_coef_out_payload_0_15_16_imag = int_reg_array_15_16_imag;
  assign io_coef_out_payload_0_15_17_real = int_reg_array_15_17_real;
  assign io_coef_out_payload_0_15_17_imag = int_reg_array_15_17_imag;
  assign io_coef_out_payload_0_15_18_real = int_reg_array_15_18_real;
  assign io_coef_out_payload_0_15_18_imag = int_reg_array_15_18_imag;
  assign io_coef_out_payload_0_15_19_real = int_reg_array_15_19_real;
  assign io_coef_out_payload_0_15_19_imag = int_reg_array_15_19_imag;
  assign io_coef_out_payload_0_15_20_real = int_reg_array_15_20_real;
  assign io_coef_out_payload_0_15_20_imag = int_reg_array_15_20_imag;
  assign io_coef_out_payload_0_15_21_real = int_reg_array_15_21_real;
  assign io_coef_out_payload_0_15_21_imag = int_reg_array_15_21_imag;
  assign io_coef_out_payload_0_15_22_real = int_reg_array_15_22_real;
  assign io_coef_out_payload_0_15_22_imag = int_reg_array_15_22_imag;
  assign io_coef_out_payload_0_15_23_real = int_reg_array_15_23_real;
  assign io_coef_out_payload_0_15_23_imag = int_reg_array_15_23_imag;
  assign io_coef_out_payload_0_15_24_real = int_reg_array_15_24_real;
  assign io_coef_out_payload_0_15_24_imag = int_reg_array_15_24_imag;
  assign io_coef_out_payload_0_15_25_real = int_reg_array_15_25_real;
  assign io_coef_out_payload_0_15_25_imag = int_reg_array_15_25_imag;
  assign io_coef_out_payload_0_15_26_real = int_reg_array_15_26_real;
  assign io_coef_out_payload_0_15_26_imag = int_reg_array_15_26_imag;
  assign io_coef_out_payload_0_15_27_real = int_reg_array_15_27_real;
  assign io_coef_out_payload_0_15_27_imag = int_reg_array_15_27_imag;
  assign io_coef_out_payload_0_15_28_real = int_reg_array_15_28_real;
  assign io_coef_out_payload_0_15_28_imag = int_reg_array_15_28_imag;
  assign io_coef_out_payload_0_15_29_real = int_reg_array_15_29_real;
  assign io_coef_out_payload_0_15_29_imag = int_reg_array_15_29_imag;
  assign io_coef_out_payload_0_15_30_real = int_reg_array_15_30_real;
  assign io_coef_out_payload_0_15_30_imag = int_reg_array_15_30_imag;
  assign io_coef_out_payload_0_15_31_real = int_reg_array_15_31_real;
  assign io_coef_out_payload_0_15_31_imag = int_reg_array_15_31_imag;
  assign io_coef_out_payload_0_15_32_real = int_reg_array_15_32_real;
  assign io_coef_out_payload_0_15_32_imag = int_reg_array_15_32_imag;
  assign io_coef_out_payload_0_15_33_real = int_reg_array_15_33_real;
  assign io_coef_out_payload_0_15_33_imag = int_reg_array_15_33_imag;
  assign io_coef_out_payload_0_15_34_real = int_reg_array_15_34_real;
  assign io_coef_out_payload_0_15_34_imag = int_reg_array_15_34_imag;
  assign io_coef_out_payload_0_15_35_real = int_reg_array_15_35_real;
  assign io_coef_out_payload_0_15_35_imag = int_reg_array_15_35_imag;
  assign io_coef_out_payload_0_15_36_real = int_reg_array_15_36_real;
  assign io_coef_out_payload_0_15_36_imag = int_reg_array_15_36_imag;
  assign io_coef_out_payload_0_15_37_real = int_reg_array_15_37_real;
  assign io_coef_out_payload_0_15_37_imag = int_reg_array_15_37_imag;
  assign io_coef_out_payload_0_15_38_real = int_reg_array_15_38_real;
  assign io_coef_out_payload_0_15_38_imag = int_reg_array_15_38_imag;
  assign io_coef_out_payload_0_15_39_real = int_reg_array_15_39_real;
  assign io_coef_out_payload_0_15_39_imag = int_reg_array_15_39_imag;
  assign io_coef_out_payload_0_15_40_real = int_reg_array_15_40_real;
  assign io_coef_out_payload_0_15_40_imag = int_reg_array_15_40_imag;
  assign io_coef_out_payload_0_15_41_real = int_reg_array_15_41_real;
  assign io_coef_out_payload_0_15_41_imag = int_reg_array_15_41_imag;
  assign io_coef_out_payload_0_15_42_real = int_reg_array_15_42_real;
  assign io_coef_out_payload_0_15_42_imag = int_reg_array_15_42_imag;
  assign io_coef_out_payload_0_15_43_real = int_reg_array_15_43_real;
  assign io_coef_out_payload_0_15_43_imag = int_reg_array_15_43_imag;
  assign io_coef_out_payload_0_15_44_real = int_reg_array_15_44_real;
  assign io_coef_out_payload_0_15_44_imag = int_reg_array_15_44_imag;
  assign io_coef_out_payload_0_15_45_real = int_reg_array_15_45_real;
  assign io_coef_out_payload_0_15_45_imag = int_reg_array_15_45_imag;
  assign io_coef_out_payload_0_15_46_real = int_reg_array_15_46_real;
  assign io_coef_out_payload_0_15_46_imag = int_reg_array_15_46_imag;
  assign io_coef_out_payload_0_15_47_real = int_reg_array_15_47_real;
  assign io_coef_out_payload_0_15_47_imag = int_reg_array_15_47_imag;
  assign io_coef_out_payload_0_15_48_real = int_reg_array_15_48_real;
  assign io_coef_out_payload_0_15_48_imag = int_reg_array_15_48_imag;
  assign io_coef_out_payload_0_15_49_real = int_reg_array_15_49_real;
  assign io_coef_out_payload_0_15_49_imag = int_reg_array_15_49_imag;
  assign io_coef_out_payload_0_16_0_real = int_reg_array_16_0_real;
  assign io_coef_out_payload_0_16_0_imag = int_reg_array_16_0_imag;
  assign io_coef_out_payload_0_16_1_real = int_reg_array_16_1_real;
  assign io_coef_out_payload_0_16_1_imag = int_reg_array_16_1_imag;
  assign io_coef_out_payload_0_16_2_real = int_reg_array_16_2_real;
  assign io_coef_out_payload_0_16_2_imag = int_reg_array_16_2_imag;
  assign io_coef_out_payload_0_16_3_real = int_reg_array_16_3_real;
  assign io_coef_out_payload_0_16_3_imag = int_reg_array_16_3_imag;
  assign io_coef_out_payload_0_16_4_real = int_reg_array_16_4_real;
  assign io_coef_out_payload_0_16_4_imag = int_reg_array_16_4_imag;
  assign io_coef_out_payload_0_16_5_real = int_reg_array_16_5_real;
  assign io_coef_out_payload_0_16_5_imag = int_reg_array_16_5_imag;
  assign io_coef_out_payload_0_16_6_real = int_reg_array_16_6_real;
  assign io_coef_out_payload_0_16_6_imag = int_reg_array_16_6_imag;
  assign io_coef_out_payload_0_16_7_real = int_reg_array_16_7_real;
  assign io_coef_out_payload_0_16_7_imag = int_reg_array_16_7_imag;
  assign io_coef_out_payload_0_16_8_real = int_reg_array_16_8_real;
  assign io_coef_out_payload_0_16_8_imag = int_reg_array_16_8_imag;
  assign io_coef_out_payload_0_16_9_real = int_reg_array_16_9_real;
  assign io_coef_out_payload_0_16_9_imag = int_reg_array_16_9_imag;
  assign io_coef_out_payload_0_16_10_real = int_reg_array_16_10_real;
  assign io_coef_out_payload_0_16_10_imag = int_reg_array_16_10_imag;
  assign io_coef_out_payload_0_16_11_real = int_reg_array_16_11_real;
  assign io_coef_out_payload_0_16_11_imag = int_reg_array_16_11_imag;
  assign io_coef_out_payload_0_16_12_real = int_reg_array_16_12_real;
  assign io_coef_out_payload_0_16_12_imag = int_reg_array_16_12_imag;
  assign io_coef_out_payload_0_16_13_real = int_reg_array_16_13_real;
  assign io_coef_out_payload_0_16_13_imag = int_reg_array_16_13_imag;
  assign io_coef_out_payload_0_16_14_real = int_reg_array_16_14_real;
  assign io_coef_out_payload_0_16_14_imag = int_reg_array_16_14_imag;
  assign io_coef_out_payload_0_16_15_real = int_reg_array_16_15_real;
  assign io_coef_out_payload_0_16_15_imag = int_reg_array_16_15_imag;
  assign io_coef_out_payload_0_16_16_real = int_reg_array_16_16_real;
  assign io_coef_out_payload_0_16_16_imag = int_reg_array_16_16_imag;
  assign io_coef_out_payload_0_16_17_real = int_reg_array_16_17_real;
  assign io_coef_out_payload_0_16_17_imag = int_reg_array_16_17_imag;
  assign io_coef_out_payload_0_16_18_real = int_reg_array_16_18_real;
  assign io_coef_out_payload_0_16_18_imag = int_reg_array_16_18_imag;
  assign io_coef_out_payload_0_16_19_real = int_reg_array_16_19_real;
  assign io_coef_out_payload_0_16_19_imag = int_reg_array_16_19_imag;
  assign io_coef_out_payload_0_16_20_real = int_reg_array_16_20_real;
  assign io_coef_out_payload_0_16_20_imag = int_reg_array_16_20_imag;
  assign io_coef_out_payload_0_16_21_real = int_reg_array_16_21_real;
  assign io_coef_out_payload_0_16_21_imag = int_reg_array_16_21_imag;
  assign io_coef_out_payload_0_16_22_real = int_reg_array_16_22_real;
  assign io_coef_out_payload_0_16_22_imag = int_reg_array_16_22_imag;
  assign io_coef_out_payload_0_16_23_real = int_reg_array_16_23_real;
  assign io_coef_out_payload_0_16_23_imag = int_reg_array_16_23_imag;
  assign io_coef_out_payload_0_16_24_real = int_reg_array_16_24_real;
  assign io_coef_out_payload_0_16_24_imag = int_reg_array_16_24_imag;
  assign io_coef_out_payload_0_16_25_real = int_reg_array_16_25_real;
  assign io_coef_out_payload_0_16_25_imag = int_reg_array_16_25_imag;
  assign io_coef_out_payload_0_16_26_real = int_reg_array_16_26_real;
  assign io_coef_out_payload_0_16_26_imag = int_reg_array_16_26_imag;
  assign io_coef_out_payload_0_16_27_real = int_reg_array_16_27_real;
  assign io_coef_out_payload_0_16_27_imag = int_reg_array_16_27_imag;
  assign io_coef_out_payload_0_16_28_real = int_reg_array_16_28_real;
  assign io_coef_out_payload_0_16_28_imag = int_reg_array_16_28_imag;
  assign io_coef_out_payload_0_16_29_real = int_reg_array_16_29_real;
  assign io_coef_out_payload_0_16_29_imag = int_reg_array_16_29_imag;
  assign io_coef_out_payload_0_16_30_real = int_reg_array_16_30_real;
  assign io_coef_out_payload_0_16_30_imag = int_reg_array_16_30_imag;
  assign io_coef_out_payload_0_16_31_real = int_reg_array_16_31_real;
  assign io_coef_out_payload_0_16_31_imag = int_reg_array_16_31_imag;
  assign io_coef_out_payload_0_16_32_real = int_reg_array_16_32_real;
  assign io_coef_out_payload_0_16_32_imag = int_reg_array_16_32_imag;
  assign io_coef_out_payload_0_16_33_real = int_reg_array_16_33_real;
  assign io_coef_out_payload_0_16_33_imag = int_reg_array_16_33_imag;
  assign io_coef_out_payload_0_16_34_real = int_reg_array_16_34_real;
  assign io_coef_out_payload_0_16_34_imag = int_reg_array_16_34_imag;
  assign io_coef_out_payload_0_16_35_real = int_reg_array_16_35_real;
  assign io_coef_out_payload_0_16_35_imag = int_reg_array_16_35_imag;
  assign io_coef_out_payload_0_16_36_real = int_reg_array_16_36_real;
  assign io_coef_out_payload_0_16_36_imag = int_reg_array_16_36_imag;
  assign io_coef_out_payload_0_16_37_real = int_reg_array_16_37_real;
  assign io_coef_out_payload_0_16_37_imag = int_reg_array_16_37_imag;
  assign io_coef_out_payload_0_16_38_real = int_reg_array_16_38_real;
  assign io_coef_out_payload_0_16_38_imag = int_reg_array_16_38_imag;
  assign io_coef_out_payload_0_16_39_real = int_reg_array_16_39_real;
  assign io_coef_out_payload_0_16_39_imag = int_reg_array_16_39_imag;
  assign io_coef_out_payload_0_16_40_real = int_reg_array_16_40_real;
  assign io_coef_out_payload_0_16_40_imag = int_reg_array_16_40_imag;
  assign io_coef_out_payload_0_16_41_real = int_reg_array_16_41_real;
  assign io_coef_out_payload_0_16_41_imag = int_reg_array_16_41_imag;
  assign io_coef_out_payload_0_16_42_real = int_reg_array_16_42_real;
  assign io_coef_out_payload_0_16_42_imag = int_reg_array_16_42_imag;
  assign io_coef_out_payload_0_16_43_real = int_reg_array_16_43_real;
  assign io_coef_out_payload_0_16_43_imag = int_reg_array_16_43_imag;
  assign io_coef_out_payload_0_16_44_real = int_reg_array_16_44_real;
  assign io_coef_out_payload_0_16_44_imag = int_reg_array_16_44_imag;
  assign io_coef_out_payload_0_16_45_real = int_reg_array_16_45_real;
  assign io_coef_out_payload_0_16_45_imag = int_reg_array_16_45_imag;
  assign io_coef_out_payload_0_16_46_real = int_reg_array_16_46_real;
  assign io_coef_out_payload_0_16_46_imag = int_reg_array_16_46_imag;
  assign io_coef_out_payload_0_16_47_real = int_reg_array_16_47_real;
  assign io_coef_out_payload_0_16_47_imag = int_reg_array_16_47_imag;
  assign io_coef_out_payload_0_16_48_real = int_reg_array_16_48_real;
  assign io_coef_out_payload_0_16_48_imag = int_reg_array_16_48_imag;
  assign io_coef_out_payload_0_16_49_real = int_reg_array_16_49_real;
  assign io_coef_out_payload_0_16_49_imag = int_reg_array_16_49_imag;
  assign io_coef_out_payload_0_17_0_real = int_reg_array_17_0_real;
  assign io_coef_out_payload_0_17_0_imag = int_reg_array_17_0_imag;
  assign io_coef_out_payload_0_17_1_real = int_reg_array_17_1_real;
  assign io_coef_out_payload_0_17_1_imag = int_reg_array_17_1_imag;
  assign io_coef_out_payload_0_17_2_real = int_reg_array_17_2_real;
  assign io_coef_out_payload_0_17_2_imag = int_reg_array_17_2_imag;
  assign io_coef_out_payload_0_17_3_real = int_reg_array_17_3_real;
  assign io_coef_out_payload_0_17_3_imag = int_reg_array_17_3_imag;
  assign io_coef_out_payload_0_17_4_real = int_reg_array_17_4_real;
  assign io_coef_out_payload_0_17_4_imag = int_reg_array_17_4_imag;
  assign io_coef_out_payload_0_17_5_real = int_reg_array_17_5_real;
  assign io_coef_out_payload_0_17_5_imag = int_reg_array_17_5_imag;
  assign io_coef_out_payload_0_17_6_real = int_reg_array_17_6_real;
  assign io_coef_out_payload_0_17_6_imag = int_reg_array_17_6_imag;
  assign io_coef_out_payload_0_17_7_real = int_reg_array_17_7_real;
  assign io_coef_out_payload_0_17_7_imag = int_reg_array_17_7_imag;
  assign io_coef_out_payload_0_17_8_real = int_reg_array_17_8_real;
  assign io_coef_out_payload_0_17_8_imag = int_reg_array_17_8_imag;
  assign io_coef_out_payload_0_17_9_real = int_reg_array_17_9_real;
  assign io_coef_out_payload_0_17_9_imag = int_reg_array_17_9_imag;
  assign io_coef_out_payload_0_17_10_real = int_reg_array_17_10_real;
  assign io_coef_out_payload_0_17_10_imag = int_reg_array_17_10_imag;
  assign io_coef_out_payload_0_17_11_real = int_reg_array_17_11_real;
  assign io_coef_out_payload_0_17_11_imag = int_reg_array_17_11_imag;
  assign io_coef_out_payload_0_17_12_real = int_reg_array_17_12_real;
  assign io_coef_out_payload_0_17_12_imag = int_reg_array_17_12_imag;
  assign io_coef_out_payload_0_17_13_real = int_reg_array_17_13_real;
  assign io_coef_out_payload_0_17_13_imag = int_reg_array_17_13_imag;
  assign io_coef_out_payload_0_17_14_real = int_reg_array_17_14_real;
  assign io_coef_out_payload_0_17_14_imag = int_reg_array_17_14_imag;
  assign io_coef_out_payload_0_17_15_real = int_reg_array_17_15_real;
  assign io_coef_out_payload_0_17_15_imag = int_reg_array_17_15_imag;
  assign io_coef_out_payload_0_17_16_real = int_reg_array_17_16_real;
  assign io_coef_out_payload_0_17_16_imag = int_reg_array_17_16_imag;
  assign io_coef_out_payload_0_17_17_real = int_reg_array_17_17_real;
  assign io_coef_out_payload_0_17_17_imag = int_reg_array_17_17_imag;
  assign io_coef_out_payload_0_17_18_real = int_reg_array_17_18_real;
  assign io_coef_out_payload_0_17_18_imag = int_reg_array_17_18_imag;
  assign io_coef_out_payload_0_17_19_real = int_reg_array_17_19_real;
  assign io_coef_out_payload_0_17_19_imag = int_reg_array_17_19_imag;
  assign io_coef_out_payload_0_17_20_real = int_reg_array_17_20_real;
  assign io_coef_out_payload_0_17_20_imag = int_reg_array_17_20_imag;
  assign io_coef_out_payload_0_17_21_real = int_reg_array_17_21_real;
  assign io_coef_out_payload_0_17_21_imag = int_reg_array_17_21_imag;
  assign io_coef_out_payload_0_17_22_real = int_reg_array_17_22_real;
  assign io_coef_out_payload_0_17_22_imag = int_reg_array_17_22_imag;
  assign io_coef_out_payload_0_17_23_real = int_reg_array_17_23_real;
  assign io_coef_out_payload_0_17_23_imag = int_reg_array_17_23_imag;
  assign io_coef_out_payload_0_17_24_real = int_reg_array_17_24_real;
  assign io_coef_out_payload_0_17_24_imag = int_reg_array_17_24_imag;
  assign io_coef_out_payload_0_17_25_real = int_reg_array_17_25_real;
  assign io_coef_out_payload_0_17_25_imag = int_reg_array_17_25_imag;
  assign io_coef_out_payload_0_17_26_real = int_reg_array_17_26_real;
  assign io_coef_out_payload_0_17_26_imag = int_reg_array_17_26_imag;
  assign io_coef_out_payload_0_17_27_real = int_reg_array_17_27_real;
  assign io_coef_out_payload_0_17_27_imag = int_reg_array_17_27_imag;
  assign io_coef_out_payload_0_17_28_real = int_reg_array_17_28_real;
  assign io_coef_out_payload_0_17_28_imag = int_reg_array_17_28_imag;
  assign io_coef_out_payload_0_17_29_real = int_reg_array_17_29_real;
  assign io_coef_out_payload_0_17_29_imag = int_reg_array_17_29_imag;
  assign io_coef_out_payload_0_17_30_real = int_reg_array_17_30_real;
  assign io_coef_out_payload_0_17_30_imag = int_reg_array_17_30_imag;
  assign io_coef_out_payload_0_17_31_real = int_reg_array_17_31_real;
  assign io_coef_out_payload_0_17_31_imag = int_reg_array_17_31_imag;
  assign io_coef_out_payload_0_17_32_real = int_reg_array_17_32_real;
  assign io_coef_out_payload_0_17_32_imag = int_reg_array_17_32_imag;
  assign io_coef_out_payload_0_17_33_real = int_reg_array_17_33_real;
  assign io_coef_out_payload_0_17_33_imag = int_reg_array_17_33_imag;
  assign io_coef_out_payload_0_17_34_real = int_reg_array_17_34_real;
  assign io_coef_out_payload_0_17_34_imag = int_reg_array_17_34_imag;
  assign io_coef_out_payload_0_17_35_real = int_reg_array_17_35_real;
  assign io_coef_out_payload_0_17_35_imag = int_reg_array_17_35_imag;
  assign io_coef_out_payload_0_17_36_real = int_reg_array_17_36_real;
  assign io_coef_out_payload_0_17_36_imag = int_reg_array_17_36_imag;
  assign io_coef_out_payload_0_17_37_real = int_reg_array_17_37_real;
  assign io_coef_out_payload_0_17_37_imag = int_reg_array_17_37_imag;
  assign io_coef_out_payload_0_17_38_real = int_reg_array_17_38_real;
  assign io_coef_out_payload_0_17_38_imag = int_reg_array_17_38_imag;
  assign io_coef_out_payload_0_17_39_real = int_reg_array_17_39_real;
  assign io_coef_out_payload_0_17_39_imag = int_reg_array_17_39_imag;
  assign io_coef_out_payload_0_17_40_real = int_reg_array_17_40_real;
  assign io_coef_out_payload_0_17_40_imag = int_reg_array_17_40_imag;
  assign io_coef_out_payload_0_17_41_real = int_reg_array_17_41_real;
  assign io_coef_out_payload_0_17_41_imag = int_reg_array_17_41_imag;
  assign io_coef_out_payload_0_17_42_real = int_reg_array_17_42_real;
  assign io_coef_out_payload_0_17_42_imag = int_reg_array_17_42_imag;
  assign io_coef_out_payload_0_17_43_real = int_reg_array_17_43_real;
  assign io_coef_out_payload_0_17_43_imag = int_reg_array_17_43_imag;
  assign io_coef_out_payload_0_17_44_real = int_reg_array_17_44_real;
  assign io_coef_out_payload_0_17_44_imag = int_reg_array_17_44_imag;
  assign io_coef_out_payload_0_17_45_real = int_reg_array_17_45_real;
  assign io_coef_out_payload_0_17_45_imag = int_reg_array_17_45_imag;
  assign io_coef_out_payload_0_17_46_real = int_reg_array_17_46_real;
  assign io_coef_out_payload_0_17_46_imag = int_reg_array_17_46_imag;
  assign io_coef_out_payload_0_17_47_real = int_reg_array_17_47_real;
  assign io_coef_out_payload_0_17_47_imag = int_reg_array_17_47_imag;
  assign io_coef_out_payload_0_17_48_real = int_reg_array_17_48_real;
  assign io_coef_out_payload_0_17_48_imag = int_reg_array_17_48_imag;
  assign io_coef_out_payload_0_17_49_real = int_reg_array_17_49_real;
  assign io_coef_out_payload_0_17_49_imag = int_reg_array_17_49_imag;
  assign io_coef_out_payload_0_18_0_real = int_reg_array_18_0_real;
  assign io_coef_out_payload_0_18_0_imag = int_reg_array_18_0_imag;
  assign io_coef_out_payload_0_18_1_real = int_reg_array_18_1_real;
  assign io_coef_out_payload_0_18_1_imag = int_reg_array_18_1_imag;
  assign io_coef_out_payload_0_18_2_real = int_reg_array_18_2_real;
  assign io_coef_out_payload_0_18_2_imag = int_reg_array_18_2_imag;
  assign io_coef_out_payload_0_18_3_real = int_reg_array_18_3_real;
  assign io_coef_out_payload_0_18_3_imag = int_reg_array_18_3_imag;
  assign io_coef_out_payload_0_18_4_real = int_reg_array_18_4_real;
  assign io_coef_out_payload_0_18_4_imag = int_reg_array_18_4_imag;
  assign io_coef_out_payload_0_18_5_real = int_reg_array_18_5_real;
  assign io_coef_out_payload_0_18_5_imag = int_reg_array_18_5_imag;
  assign io_coef_out_payload_0_18_6_real = int_reg_array_18_6_real;
  assign io_coef_out_payload_0_18_6_imag = int_reg_array_18_6_imag;
  assign io_coef_out_payload_0_18_7_real = int_reg_array_18_7_real;
  assign io_coef_out_payload_0_18_7_imag = int_reg_array_18_7_imag;
  assign io_coef_out_payload_0_18_8_real = int_reg_array_18_8_real;
  assign io_coef_out_payload_0_18_8_imag = int_reg_array_18_8_imag;
  assign io_coef_out_payload_0_18_9_real = int_reg_array_18_9_real;
  assign io_coef_out_payload_0_18_9_imag = int_reg_array_18_9_imag;
  assign io_coef_out_payload_0_18_10_real = int_reg_array_18_10_real;
  assign io_coef_out_payload_0_18_10_imag = int_reg_array_18_10_imag;
  assign io_coef_out_payload_0_18_11_real = int_reg_array_18_11_real;
  assign io_coef_out_payload_0_18_11_imag = int_reg_array_18_11_imag;
  assign io_coef_out_payload_0_18_12_real = int_reg_array_18_12_real;
  assign io_coef_out_payload_0_18_12_imag = int_reg_array_18_12_imag;
  assign io_coef_out_payload_0_18_13_real = int_reg_array_18_13_real;
  assign io_coef_out_payload_0_18_13_imag = int_reg_array_18_13_imag;
  assign io_coef_out_payload_0_18_14_real = int_reg_array_18_14_real;
  assign io_coef_out_payload_0_18_14_imag = int_reg_array_18_14_imag;
  assign io_coef_out_payload_0_18_15_real = int_reg_array_18_15_real;
  assign io_coef_out_payload_0_18_15_imag = int_reg_array_18_15_imag;
  assign io_coef_out_payload_0_18_16_real = int_reg_array_18_16_real;
  assign io_coef_out_payload_0_18_16_imag = int_reg_array_18_16_imag;
  assign io_coef_out_payload_0_18_17_real = int_reg_array_18_17_real;
  assign io_coef_out_payload_0_18_17_imag = int_reg_array_18_17_imag;
  assign io_coef_out_payload_0_18_18_real = int_reg_array_18_18_real;
  assign io_coef_out_payload_0_18_18_imag = int_reg_array_18_18_imag;
  assign io_coef_out_payload_0_18_19_real = int_reg_array_18_19_real;
  assign io_coef_out_payload_0_18_19_imag = int_reg_array_18_19_imag;
  assign io_coef_out_payload_0_18_20_real = int_reg_array_18_20_real;
  assign io_coef_out_payload_0_18_20_imag = int_reg_array_18_20_imag;
  assign io_coef_out_payload_0_18_21_real = int_reg_array_18_21_real;
  assign io_coef_out_payload_0_18_21_imag = int_reg_array_18_21_imag;
  assign io_coef_out_payload_0_18_22_real = int_reg_array_18_22_real;
  assign io_coef_out_payload_0_18_22_imag = int_reg_array_18_22_imag;
  assign io_coef_out_payload_0_18_23_real = int_reg_array_18_23_real;
  assign io_coef_out_payload_0_18_23_imag = int_reg_array_18_23_imag;
  assign io_coef_out_payload_0_18_24_real = int_reg_array_18_24_real;
  assign io_coef_out_payload_0_18_24_imag = int_reg_array_18_24_imag;
  assign io_coef_out_payload_0_18_25_real = int_reg_array_18_25_real;
  assign io_coef_out_payload_0_18_25_imag = int_reg_array_18_25_imag;
  assign io_coef_out_payload_0_18_26_real = int_reg_array_18_26_real;
  assign io_coef_out_payload_0_18_26_imag = int_reg_array_18_26_imag;
  assign io_coef_out_payload_0_18_27_real = int_reg_array_18_27_real;
  assign io_coef_out_payload_0_18_27_imag = int_reg_array_18_27_imag;
  assign io_coef_out_payload_0_18_28_real = int_reg_array_18_28_real;
  assign io_coef_out_payload_0_18_28_imag = int_reg_array_18_28_imag;
  assign io_coef_out_payload_0_18_29_real = int_reg_array_18_29_real;
  assign io_coef_out_payload_0_18_29_imag = int_reg_array_18_29_imag;
  assign io_coef_out_payload_0_18_30_real = int_reg_array_18_30_real;
  assign io_coef_out_payload_0_18_30_imag = int_reg_array_18_30_imag;
  assign io_coef_out_payload_0_18_31_real = int_reg_array_18_31_real;
  assign io_coef_out_payload_0_18_31_imag = int_reg_array_18_31_imag;
  assign io_coef_out_payload_0_18_32_real = int_reg_array_18_32_real;
  assign io_coef_out_payload_0_18_32_imag = int_reg_array_18_32_imag;
  assign io_coef_out_payload_0_18_33_real = int_reg_array_18_33_real;
  assign io_coef_out_payload_0_18_33_imag = int_reg_array_18_33_imag;
  assign io_coef_out_payload_0_18_34_real = int_reg_array_18_34_real;
  assign io_coef_out_payload_0_18_34_imag = int_reg_array_18_34_imag;
  assign io_coef_out_payload_0_18_35_real = int_reg_array_18_35_real;
  assign io_coef_out_payload_0_18_35_imag = int_reg_array_18_35_imag;
  assign io_coef_out_payload_0_18_36_real = int_reg_array_18_36_real;
  assign io_coef_out_payload_0_18_36_imag = int_reg_array_18_36_imag;
  assign io_coef_out_payload_0_18_37_real = int_reg_array_18_37_real;
  assign io_coef_out_payload_0_18_37_imag = int_reg_array_18_37_imag;
  assign io_coef_out_payload_0_18_38_real = int_reg_array_18_38_real;
  assign io_coef_out_payload_0_18_38_imag = int_reg_array_18_38_imag;
  assign io_coef_out_payload_0_18_39_real = int_reg_array_18_39_real;
  assign io_coef_out_payload_0_18_39_imag = int_reg_array_18_39_imag;
  assign io_coef_out_payload_0_18_40_real = int_reg_array_18_40_real;
  assign io_coef_out_payload_0_18_40_imag = int_reg_array_18_40_imag;
  assign io_coef_out_payload_0_18_41_real = int_reg_array_18_41_real;
  assign io_coef_out_payload_0_18_41_imag = int_reg_array_18_41_imag;
  assign io_coef_out_payload_0_18_42_real = int_reg_array_18_42_real;
  assign io_coef_out_payload_0_18_42_imag = int_reg_array_18_42_imag;
  assign io_coef_out_payload_0_18_43_real = int_reg_array_18_43_real;
  assign io_coef_out_payload_0_18_43_imag = int_reg_array_18_43_imag;
  assign io_coef_out_payload_0_18_44_real = int_reg_array_18_44_real;
  assign io_coef_out_payload_0_18_44_imag = int_reg_array_18_44_imag;
  assign io_coef_out_payload_0_18_45_real = int_reg_array_18_45_real;
  assign io_coef_out_payload_0_18_45_imag = int_reg_array_18_45_imag;
  assign io_coef_out_payload_0_18_46_real = int_reg_array_18_46_real;
  assign io_coef_out_payload_0_18_46_imag = int_reg_array_18_46_imag;
  assign io_coef_out_payload_0_18_47_real = int_reg_array_18_47_real;
  assign io_coef_out_payload_0_18_47_imag = int_reg_array_18_47_imag;
  assign io_coef_out_payload_0_18_48_real = int_reg_array_18_48_real;
  assign io_coef_out_payload_0_18_48_imag = int_reg_array_18_48_imag;
  assign io_coef_out_payload_0_18_49_real = int_reg_array_18_49_real;
  assign io_coef_out_payload_0_18_49_imag = int_reg_array_18_49_imag;
  assign io_coef_out_payload_0_19_0_real = int_reg_array_19_0_real;
  assign io_coef_out_payload_0_19_0_imag = int_reg_array_19_0_imag;
  assign io_coef_out_payload_0_19_1_real = int_reg_array_19_1_real;
  assign io_coef_out_payload_0_19_1_imag = int_reg_array_19_1_imag;
  assign io_coef_out_payload_0_19_2_real = int_reg_array_19_2_real;
  assign io_coef_out_payload_0_19_2_imag = int_reg_array_19_2_imag;
  assign io_coef_out_payload_0_19_3_real = int_reg_array_19_3_real;
  assign io_coef_out_payload_0_19_3_imag = int_reg_array_19_3_imag;
  assign io_coef_out_payload_0_19_4_real = int_reg_array_19_4_real;
  assign io_coef_out_payload_0_19_4_imag = int_reg_array_19_4_imag;
  assign io_coef_out_payload_0_19_5_real = int_reg_array_19_5_real;
  assign io_coef_out_payload_0_19_5_imag = int_reg_array_19_5_imag;
  assign io_coef_out_payload_0_19_6_real = int_reg_array_19_6_real;
  assign io_coef_out_payload_0_19_6_imag = int_reg_array_19_6_imag;
  assign io_coef_out_payload_0_19_7_real = int_reg_array_19_7_real;
  assign io_coef_out_payload_0_19_7_imag = int_reg_array_19_7_imag;
  assign io_coef_out_payload_0_19_8_real = int_reg_array_19_8_real;
  assign io_coef_out_payload_0_19_8_imag = int_reg_array_19_8_imag;
  assign io_coef_out_payload_0_19_9_real = int_reg_array_19_9_real;
  assign io_coef_out_payload_0_19_9_imag = int_reg_array_19_9_imag;
  assign io_coef_out_payload_0_19_10_real = int_reg_array_19_10_real;
  assign io_coef_out_payload_0_19_10_imag = int_reg_array_19_10_imag;
  assign io_coef_out_payload_0_19_11_real = int_reg_array_19_11_real;
  assign io_coef_out_payload_0_19_11_imag = int_reg_array_19_11_imag;
  assign io_coef_out_payload_0_19_12_real = int_reg_array_19_12_real;
  assign io_coef_out_payload_0_19_12_imag = int_reg_array_19_12_imag;
  assign io_coef_out_payload_0_19_13_real = int_reg_array_19_13_real;
  assign io_coef_out_payload_0_19_13_imag = int_reg_array_19_13_imag;
  assign io_coef_out_payload_0_19_14_real = int_reg_array_19_14_real;
  assign io_coef_out_payload_0_19_14_imag = int_reg_array_19_14_imag;
  assign io_coef_out_payload_0_19_15_real = int_reg_array_19_15_real;
  assign io_coef_out_payload_0_19_15_imag = int_reg_array_19_15_imag;
  assign io_coef_out_payload_0_19_16_real = int_reg_array_19_16_real;
  assign io_coef_out_payload_0_19_16_imag = int_reg_array_19_16_imag;
  assign io_coef_out_payload_0_19_17_real = int_reg_array_19_17_real;
  assign io_coef_out_payload_0_19_17_imag = int_reg_array_19_17_imag;
  assign io_coef_out_payload_0_19_18_real = int_reg_array_19_18_real;
  assign io_coef_out_payload_0_19_18_imag = int_reg_array_19_18_imag;
  assign io_coef_out_payload_0_19_19_real = int_reg_array_19_19_real;
  assign io_coef_out_payload_0_19_19_imag = int_reg_array_19_19_imag;
  assign io_coef_out_payload_0_19_20_real = int_reg_array_19_20_real;
  assign io_coef_out_payload_0_19_20_imag = int_reg_array_19_20_imag;
  assign io_coef_out_payload_0_19_21_real = int_reg_array_19_21_real;
  assign io_coef_out_payload_0_19_21_imag = int_reg_array_19_21_imag;
  assign io_coef_out_payload_0_19_22_real = int_reg_array_19_22_real;
  assign io_coef_out_payload_0_19_22_imag = int_reg_array_19_22_imag;
  assign io_coef_out_payload_0_19_23_real = int_reg_array_19_23_real;
  assign io_coef_out_payload_0_19_23_imag = int_reg_array_19_23_imag;
  assign io_coef_out_payload_0_19_24_real = int_reg_array_19_24_real;
  assign io_coef_out_payload_0_19_24_imag = int_reg_array_19_24_imag;
  assign io_coef_out_payload_0_19_25_real = int_reg_array_19_25_real;
  assign io_coef_out_payload_0_19_25_imag = int_reg_array_19_25_imag;
  assign io_coef_out_payload_0_19_26_real = int_reg_array_19_26_real;
  assign io_coef_out_payload_0_19_26_imag = int_reg_array_19_26_imag;
  assign io_coef_out_payload_0_19_27_real = int_reg_array_19_27_real;
  assign io_coef_out_payload_0_19_27_imag = int_reg_array_19_27_imag;
  assign io_coef_out_payload_0_19_28_real = int_reg_array_19_28_real;
  assign io_coef_out_payload_0_19_28_imag = int_reg_array_19_28_imag;
  assign io_coef_out_payload_0_19_29_real = int_reg_array_19_29_real;
  assign io_coef_out_payload_0_19_29_imag = int_reg_array_19_29_imag;
  assign io_coef_out_payload_0_19_30_real = int_reg_array_19_30_real;
  assign io_coef_out_payload_0_19_30_imag = int_reg_array_19_30_imag;
  assign io_coef_out_payload_0_19_31_real = int_reg_array_19_31_real;
  assign io_coef_out_payload_0_19_31_imag = int_reg_array_19_31_imag;
  assign io_coef_out_payload_0_19_32_real = int_reg_array_19_32_real;
  assign io_coef_out_payload_0_19_32_imag = int_reg_array_19_32_imag;
  assign io_coef_out_payload_0_19_33_real = int_reg_array_19_33_real;
  assign io_coef_out_payload_0_19_33_imag = int_reg_array_19_33_imag;
  assign io_coef_out_payload_0_19_34_real = int_reg_array_19_34_real;
  assign io_coef_out_payload_0_19_34_imag = int_reg_array_19_34_imag;
  assign io_coef_out_payload_0_19_35_real = int_reg_array_19_35_real;
  assign io_coef_out_payload_0_19_35_imag = int_reg_array_19_35_imag;
  assign io_coef_out_payload_0_19_36_real = int_reg_array_19_36_real;
  assign io_coef_out_payload_0_19_36_imag = int_reg_array_19_36_imag;
  assign io_coef_out_payload_0_19_37_real = int_reg_array_19_37_real;
  assign io_coef_out_payload_0_19_37_imag = int_reg_array_19_37_imag;
  assign io_coef_out_payload_0_19_38_real = int_reg_array_19_38_real;
  assign io_coef_out_payload_0_19_38_imag = int_reg_array_19_38_imag;
  assign io_coef_out_payload_0_19_39_real = int_reg_array_19_39_real;
  assign io_coef_out_payload_0_19_39_imag = int_reg_array_19_39_imag;
  assign io_coef_out_payload_0_19_40_real = int_reg_array_19_40_real;
  assign io_coef_out_payload_0_19_40_imag = int_reg_array_19_40_imag;
  assign io_coef_out_payload_0_19_41_real = int_reg_array_19_41_real;
  assign io_coef_out_payload_0_19_41_imag = int_reg_array_19_41_imag;
  assign io_coef_out_payload_0_19_42_real = int_reg_array_19_42_real;
  assign io_coef_out_payload_0_19_42_imag = int_reg_array_19_42_imag;
  assign io_coef_out_payload_0_19_43_real = int_reg_array_19_43_real;
  assign io_coef_out_payload_0_19_43_imag = int_reg_array_19_43_imag;
  assign io_coef_out_payload_0_19_44_real = int_reg_array_19_44_real;
  assign io_coef_out_payload_0_19_44_imag = int_reg_array_19_44_imag;
  assign io_coef_out_payload_0_19_45_real = int_reg_array_19_45_real;
  assign io_coef_out_payload_0_19_45_imag = int_reg_array_19_45_imag;
  assign io_coef_out_payload_0_19_46_real = int_reg_array_19_46_real;
  assign io_coef_out_payload_0_19_46_imag = int_reg_array_19_46_imag;
  assign io_coef_out_payload_0_19_47_real = int_reg_array_19_47_real;
  assign io_coef_out_payload_0_19_47_imag = int_reg_array_19_47_imag;
  assign io_coef_out_payload_0_19_48_real = int_reg_array_19_48_real;
  assign io_coef_out_payload_0_19_48_imag = int_reg_array_19_48_imag;
  assign io_coef_out_payload_0_19_49_real = int_reg_array_19_49_real;
  assign io_coef_out_payload_0_19_49_imag = int_reg_array_19_49_imag;
  assign io_coef_out_payload_0_20_0_real = int_reg_array_20_0_real;
  assign io_coef_out_payload_0_20_0_imag = int_reg_array_20_0_imag;
  assign io_coef_out_payload_0_20_1_real = int_reg_array_20_1_real;
  assign io_coef_out_payload_0_20_1_imag = int_reg_array_20_1_imag;
  assign io_coef_out_payload_0_20_2_real = int_reg_array_20_2_real;
  assign io_coef_out_payload_0_20_2_imag = int_reg_array_20_2_imag;
  assign io_coef_out_payload_0_20_3_real = int_reg_array_20_3_real;
  assign io_coef_out_payload_0_20_3_imag = int_reg_array_20_3_imag;
  assign io_coef_out_payload_0_20_4_real = int_reg_array_20_4_real;
  assign io_coef_out_payload_0_20_4_imag = int_reg_array_20_4_imag;
  assign io_coef_out_payload_0_20_5_real = int_reg_array_20_5_real;
  assign io_coef_out_payload_0_20_5_imag = int_reg_array_20_5_imag;
  assign io_coef_out_payload_0_20_6_real = int_reg_array_20_6_real;
  assign io_coef_out_payload_0_20_6_imag = int_reg_array_20_6_imag;
  assign io_coef_out_payload_0_20_7_real = int_reg_array_20_7_real;
  assign io_coef_out_payload_0_20_7_imag = int_reg_array_20_7_imag;
  assign io_coef_out_payload_0_20_8_real = int_reg_array_20_8_real;
  assign io_coef_out_payload_0_20_8_imag = int_reg_array_20_8_imag;
  assign io_coef_out_payload_0_20_9_real = int_reg_array_20_9_real;
  assign io_coef_out_payload_0_20_9_imag = int_reg_array_20_9_imag;
  assign io_coef_out_payload_0_20_10_real = int_reg_array_20_10_real;
  assign io_coef_out_payload_0_20_10_imag = int_reg_array_20_10_imag;
  assign io_coef_out_payload_0_20_11_real = int_reg_array_20_11_real;
  assign io_coef_out_payload_0_20_11_imag = int_reg_array_20_11_imag;
  assign io_coef_out_payload_0_20_12_real = int_reg_array_20_12_real;
  assign io_coef_out_payload_0_20_12_imag = int_reg_array_20_12_imag;
  assign io_coef_out_payload_0_20_13_real = int_reg_array_20_13_real;
  assign io_coef_out_payload_0_20_13_imag = int_reg_array_20_13_imag;
  assign io_coef_out_payload_0_20_14_real = int_reg_array_20_14_real;
  assign io_coef_out_payload_0_20_14_imag = int_reg_array_20_14_imag;
  assign io_coef_out_payload_0_20_15_real = int_reg_array_20_15_real;
  assign io_coef_out_payload_0_20_15_imag = int_reg_array_20_15_imag;
  assign io_coef_out_payload_0_20_16_real = int_reg_array_20_16_real;
  assign io_coef_out_payload_0_20_16_imag = int_reg_array_20_16_imag;
  assign io_coef_out_payload_0_20_17_real = int_reg_array_20_17_real;
  assign io_coef_out_payload_0_20_17_imag = int_reg_array_20_17_imag;
  assign io_coef_out_payload_0_20_18_real = int_reg_array_20_18_real;
  assign io_coef_out_payload_0_20_18_imag = int_reg_array_20_18_imag;
  assign io_coef_out_payload_0_20_19_real = int_reg_array_20_19_real;
  assign io_coef_out_payload_0_20_19_imag = int_reg_array_20_19_imag;
  assign io_coef_out_payload_0_20_20_real = int_reg_array_20_20_real;
  assign io_coef_out_payload_0_20_20_imag = int_reg_array_20_20_imag;
  assign io_coef_out_payload_0_20_21_real = int_reg_array_20_21_real;
  assign io_coef_out_payload_0_20_21_imag = int_reg_array_20_21_imag;
  assign io_coef_out_payload_0_20_22_real = int_reg_array_20_22_real;
  assign io_coef_out_payload_0_20_22_imag = int_reg_array_20_22_imag;
  assign io_coef_out_payload_0_20_23_real = int_reg_array_20_23_real;
  assign io_coef_out_payload_0_20_23_imag = int_reg_array_20_23_imag;
  assign io_coef_out_payload_0_20_24_real = int_reg_array_20_24_real;
  assign io_coef_out_payload_0_20_24_imag = int_reg_array_20_24_imag;
  assign io_coef_out_payload_0_20_25_real = int_reg_array_20_25_real;
  assign io_coef_out_payload_0_20_25_imag = int_reg_array_20_25_imag;
  assign io_coef_out_payload_0_20_26_real = int_reg_array_20_26_real;
  assign io_coef_out_payload_0_20_26_imag = int_reg_array_20_26_imag;
  assign io_coef_out_payload_0_20_27_real = int_reg_array_20_27_real;
  assign io_coef_out_payload_0_20_27_imag = int_reg_array_20_27_imag;
  assign io_coef_out_payload_0_20_28_real = int_reg_array_20_28_real;
  assign io_coef_out_payload_0_20_28_imag = int_reg_array_20_28_imag;
  assign io_coef_out_payload_0_20_29_real = int_reg_array_20_29_real;
  assign io_coef_out_payload_0_20_29_imag = int_reg_array_20_29_imag;
  assign io_coef_out_payload_0_20_30_real = int_reg_array_20_30_real;
  assign io_coef_out_payload_0_20_30_imag = int_reg_array_20_30_imag;
  assign io_coef_out_payload_0_20_31_real = int_reg_array_20_31_real;
  assign io_coef_out_payload_0_20_31_imag = int_reg_array_20_31_imag;
  assign io_coef_out_payload_0_20_32_real = int_reg_array_20_32_real;
  assign io_coef_out_payload_0_20_32_imag = int_reg_array_20_32_imag;
  assign io_coef_out_payload_0_20_33_real = int_reg_array_20_33_real;
  assign io_coef_out_payload_0_20_33_imag = int_reg_array_20_33_imag;
  assign io_coef_out_payload_0_20_34_real = int_reg_array_20_34_real;
  assign io_coef_out_payload_0_20_34_imag = int_reg_array_20_34_imag;
  assign io_coef_out_payload_0_20_35_real = int_reg_array_20_35_real;
  assign io_coef_out_payload_0_20_35_imag = int_reg_array_20_35_imag;
  assign io_coef_out_payload_0_20_36_real = int_reg_array_20_36_real;
  assign io_coef_out_payload_0_20_36_imag = int_reg_array_20_36_imag;
  assign io_coef_out_payload_0_20_37_real = int_reg_array_20_37_real;
  assign io_coef_out_payload_0_20_37_imag = int_reg_array_20_37_imag;
  assign io_coef_out_payload_0_20_38_real = int_reg_array_20_38_real;
  assign io_coef_out_payload_0_20_38_imag = int_reg_array_20_38_imag;
  assign io_coef_out_payload_0_20_39_real = int_reg_array_20_39_real;
  assign io_coef_out_payload_0_20_39_imag = int_reg_array_20_39_imag;
  assign io_coef_out_payload_0_20_40_real = int_reg_array_20_40_real;
  assign io_coef_out_payload_0_20_40_imag = int_reg_array_20_40_imag;
  assign io_coef_out_payload_0_20_41_real = int_reg_array_20_41_real;
  assign io_coef_out_payload_0_20_41_imag = int_reg_array_20_41_imag;
  assign io_coef_out_payload_0_20_42_real = int_reg_array_20_42_real;
  assign io_coef_out_payload_0_20_42_imag = int_reg_array_20_42_imag;
  assign io_coef_out_payload_0_20_43_real = int_reg_array_20_43_real;
  assign io_coef_out_payload_0_20_43_imag = int_reg_array_20_43_imag;
  assign io_coef_out_payload_0_20_44_real = int_reg_array_20_44_real;
  assign io_coef_out_payload_0_20_44_imag = int_reg_array_20_44_imag;
  assign io_coef_out_payload_0_20_45_real = int_reg_array_20_45_real;
  assign io_coef_out_payload_0_20_45_imag = int_reg_array_20_45_imag;
  assign io_coef_out_payload_0_20_46_real = int_reg_array_20_46_real;
  assign io_coef_out_payload_0_20_46_imag = int_reg_array_20_46_imag;
  assign io_coef_out_payload_0_20_47_real = int_reg_array_20_47_real;
  assign io_coef_out_payload_0_20_47_imag = int_reg_array_20_47_imag;
  assign io_coef_out_payload_0_20_48_real = int_reg_array_20_48_real;
  assign io_coef_out_payload_0_20_48_imag = int_reg_array_20_48_imag;
  assign io_coef_out_payload_0_20_49_real = int_reg_array_20_49_real;
  assign io_coef_out_payload_0_20_49_imag = int_reg_array_20_49_imag;
  assign io_coef_out_payload_0_21_0_real = int_reg_array_21_0_real;
  assign io_coef_out_payload_0_21_0_imag = int_reg_array_21_0_imag;
  assign io_coef_out_payload_0_21_1_real = int_reg_array_21_1_real;
  assign io_coef_out_payload_0_21_1_imag = int_reg_array_21_1_imag;
  assign io_coef_out_payload_0_21_2_real = int_reg_array_21_2_real;
  assign io_coef_out_payload_0_21_2_imag = int_reg_array_21_2_imag;
  assign io_coef_out_payload_0_21_3_real = int_reg_array_21_3_real;
  assign io_coef_out_payload_0_21_3_imag = int_reg_array_21_3_imag;
  assign io_coef_out_payload_0_21_4_real = int_reg_array_21_4_real;
  assign io_coef_out_payload_0_21_4_imag = int_reg_array_21_4_imag;
  assign io_coef_out_payload_0_21_5_real = int_reg_array_21_5_real;
  assign io_coef_out_payload_0_21_5_imag = int_reg_array_21_5_imag;
  assign io_coef_out_payload_0_21_6_real = int_reg_array_21_6_real;
  assign io_coef_out_payload_0_21_6_imag = int_reg_array_21_6_imag;
  assign io_coef_out_payload_0_21_7_real = int_reg_array_21_7_real;
  assign io_coef_out_payload_0_21_7_imag = int_reg_array_21_7_imag;
  assign io_coef_out_payload_0_21_8_real = int_reg_array_21_8_real;
  assign io_coef_out_payload_0_21_8_imag = int_reg_array_21_8_imag;
  assign io_coef_out_payload_0_21_9_real = int_reg_array_21_9_real;
  assign io_coef_out_payload_0_21_9_imag = int_reg_array_21_9_imag;
  assign io_coef_out_payload_0_21_10_real = int_reg_array_21_10_real;
  assign io_coef_out_payload_0_21_10_imag = int_reg_array_21_10_imag;
  assign io_coef_out_payload_0_21_11_real = int_reg_array_21_11_real;
  assign io_coef_out_payload_0_21_11_imag = int_reg_array_21_11_imag;
  assign io_coef_out_payload_0_21_12_real = int_reg_array_21_12_real;
  assign io_coef_out_payload_0_21_12_imag = int_reg_array_21_12_imag;
  assign io_coef_out_payload_0_21_13_real = int_reg_array_21_13_real;
  assign io_coef_out_payload_0_21_13_imag = int_reg_array_21_13_imag;
  assign io_coef_out_payload_0_21_14_real = int_reg_array_21_14_real;
  assign io_coef_out_payload_0_21_14_imag = int_reg_array_21_14_imag;
  assign io_coef_out_payload_0_21_15_real = int_reg_array_21_15_real;
  assign io_coef_out_payload_0_21_15_imag = int_reg_array_21_15_imag;
  assign io_coef_out_payload_0_21_16_real = int_reg_array_21_16_real;
  assign io_coef_out_payload_0_21_16_imag = int_reg_array_21_16_imag;
  assign io_coef_out_payload_0_21_17_real = int_reg_array_21_17_real;
  assign io_coef_out_payload_0_21_17_imag = int_reg_array_21_17_imag;
  assign io_coef_out_payload_0_21_18_real = int_reg_array_21_18_real;
  assign io_coef_out_payload_0_21_18_imag = int_reg_array_21_18_imag;
  assign io_coef_out_payload_0_21_19_real = int_reg_array_21_19_real;
  assign io_coef_out_payload_0_21_19_imag = int_reg_array_21_19_imag;
  assign io_coef_out_payload_0_21_20_real = int_reg_array_21_20_real;
  assign io_coef_out_payload_0_21_20_imag = int_reg_array_21_20_imag;
  assign io_coef_out_payload_0_21_21_real = int_reg_array_21_21_real;
  assign io_coef_out_payload_0_21_21_imag = int_reg_array_21_21_imag;
  assign io_coef_out_payload_0_21_22_real = int_reg_array_21_22_real;
  assign io_coef_out_payload_0_21_22_imag = int_reg_array_21_22_imag;
  assign io_coef_out_payload_0_21_23_real = int_reg_array_21_23_real;
  assign io_coef_out_payload_0_21_23_imag = int_reg_array_21_23_imag;
  assign io_coef_out_payload_0_21_24_real = int_reg_array_21_24_real;
  assign io_coef_out_payload_0_21_24_imag = int_reg_array_21_24_imag;
  assign io_coef_out_payload_0_21_25_real = int_reg_array_21_25_real;
  assign io_coef_out_payload_0_21_25_imag = int_reg_array_21_25_imag;
  assign io_coef_out_payload_0_21_26_real = int_reg_array_21_26_real;
  assign io_coef_out_payload_0_21_26_imag = int_reg_array_21_26_imag;
  assign io_coef_out_payload_0_21_27_real = int_reg_array_21_27_real;
  assign io_coef_out_payload_0_21_27_imag = int_reg_array_21_27_imag;
  assign io_coef_out_payload_0_21_28_real = int_reg_array_21_28_real;
  assign io_coef_out_payload_0_21_28_imag = int_reg_array_21_28_imag;
  assign io_coef_out_payload_0_21_29_real = int_reg_array_21_29_real;
  assign io_coef_out_payload_0_21_29_imag = int_reg_array_21_29_imag;
  assign io_coef_out_payload_0_21_30_real = int_reg_array_21_30_real;
  assign io_coef_out_payload_0_21_30_imag = int_reg_array_21_30_imag;
  assign io_coef_out_payload_0_21_31_real = int_reg_array_21_31_real;
  assign io_coef_out_payload_0_21_31_imag = int_reg_array_21_31_imag;
  assign io_coef_out_payload_0_21_32_real = int_reg_array_21_32_real;
  assign io_coef_out_payload_0_21_32_imag = int_reg_array_21_32_imag;
  assign io_coef_out_payload_0_21_33_real = int_reg_array_21_33_real;
  assign io_coef_out_payload_0_21_33_imag = int_reg_array_21_33_imag;
  assign io_coef_out_payload_0_21_34_real = int_reg_array_21_34_real;
  assign io_coef_out_payload_0_21_34_imag = int_reg_array_21_34_imag;
  assign io_coef_out_payload_0_21_35_real = int_reg_array_21_35_real;
  assign io_coef_out_payload_0_21_35_imag = int_reg_array_21_35_imag;
  assign io_coef_out_payload_0_21_36_real = int_reg_array_21_36_real;
  assign io_coef_out_payload_0_21_36_imag = int_reg_array_21_36_imag;
  assign io_coef_out_payload_0_21_37_real = int_reg_array_21_37_real;
  assign io_coef_out_payload_0_21_37_imag = int_reg_array_21_37_imag;
  assign io_coef_out_payload_0_21_38_real = int_reg_array_21_38_real;
  assign io_coef_out_payload_0_21_38_imag = int_reg_array_21_38_imag;
  assign io_coef_out_payload_0_21_39_real = int_reg_array_21_39_real;
  assign io_coef_out_payload_0_21_39_imag = int_reg_array_21_39_imag;
  assign io_coef_out_payload_0_21_40_real = int_reg_array_21_40_real;
  assign io_coef_out_payload_0_21_40_imag = int_reg_array_21_40_imag;
  assign io_coef_out_payload_0_21_41_real = int_reg_array_21_41_real;
  assign io_coef_out_payload_0_21_41_imag = int_reg_array_21_41_imag;
  assign io_coef_out_payload_0_21_42_real = int_reg_array_21_42_real;
  assign io_coef_out_payload_0_21_42_imag = int_reg_array_21_42_imag;
  assign io_coef_out_payload_0_21_43_real = int_reg_array_21_43_real;
  assign io_coef_out_payload_0_21_43_imag = int_reg_array_21_43_imag;
  assign io_coef_out_payload_0_21_44_real = int_reg_array_21_44_real;
  assign io_coef_out_payload_0_21_44_imag = int_reg_array_21_44_imag;
  assign io_coef_out_payload_0_21_45_real = int_reg_array_21_45_real;
  assign io_coef_out_payload_0_21_45_imag = int_reg_array_21_45_imag;
  assign io_coef_out_payload_0_21_46_real = int_reg_array_21_46_real;
  assign io_coef_out_payload_0_21_46_imag = int_reg_array_21_46_imag;
  assign io_coef_out_payload_0_21_47_real = int_reg_array_21_47_real;
  assign io_coef_out_payload_0_21_47_imag = int_reg_array_21_47_imag;
  assign io_coef_out_payload_0_21_48_real = int_reg_array_21_48_real;
  assign io_coef_out_payload_0_21_48_imag = int_reg_array_21_48_imag;
  assign io_coef_out_payload_0_21_49_real = int_reg_array_21_49_real;
  assign io_coef_out_payload_0_21_49_imag = int_reg_array_21_49_imag;
  assign io_coef_out_payload_0_22_0_real = int_reg_array_22_0_real;
  assign io_coef_out_payload_0_22_0_imag = int_reg_array_22_0_imag;
  assign io_coef_out_payload_0_22_1_real = int_reg_array_22_1_real;
  assign io_coef_out_payload_0_22_1_imag = int_reg_array_22_1_imag;
  assign io_coef_out_payload_0_22_2_real = int_reg_array_22_2_real;
  assign io_coef_out_payload_0_22_2_imag = int_reg_array_22_2_imag;
  assign io_coef_out_payload_0_22_3_real = int_reg_array_22_3_real;
  assign io_coef_out_payload_0_22_3_imag = int_reg_array_22_3_imag;
  assign io_coef_out_payload_0_22_4_real = int_reg_array_22_4_real;
  assign io_coef_out_payload_0_22_4_imag = int_reg_array_22_4_imag;
  assign io_coef_out_payload_0_22_5_real = int_reg_array_22_5_real;
  assign io_coef_out_payload_0_22_5_imag = int_reg_array_22_5_imag;
  assign io_coef_out_payload_0_22_6_real = int_reg_array_22_6_real;
  assign io_coef_out_payload_0_22_6_imag = int_reg_array_22_6_imag;
  assign io_coef_out_payload_0_22_7_real = int_reg_array_22_7_real;
  assign io_coef_out_payload_0_22_7_imag = int_reg_array_22_7_imag;
  assign io_coef_out_payload_0_22_8_real = int_reg_array_22_8_real;
  assign io_coef_out_payload_0_22_8_imag = int_reg_array_22_8_imag;
  assign io_coef_out_payload_0_22_9_real = int_reg_array_22_9_real;
  assign io_coef_out_payload_0_22_9_imag = int_reg_array_22_9_imag;
  assign io_coef_out_payload_0_22_10_real = int_reg_array_22_10_real;
  assign io_coef_out_payload_0_22_10_imag = int_reg_array_22_10_imag;
  assign io_coef_out_payload_0_22_11_real = int_reg_array_22_11_real;
  assign io_coef_out_payload_0_22_11_imag = int_reg_array_22_11_imag;
  assign io_coef_out_payload_0_22_12_real = int_reg_array_22_12_real;
  assign io_coef_out_payload_0_22_12_imag = int_reg_array_22_12_imag;
  assign io_coef_out_payload_0_22_13_real = int_reg_array_22_13_real;
  assign io_coef_out_payload_0_22_13_imag = int_reg_array_22_13_imag;
  assign io_coef_out_payload_0_22_14_real = int_reg_array_22_14_real;
  assign io_coef_out_payload_0_22_14_imag = int_reg_array_22_14_imag;
  assign io_coef_out_payload_0_22_15_real = int_reg_array_22_15_real;
  assign io_coef_out_payload_0_22_15_imag = int_reg_array_22_15_imag;
  assign io_coef_out_payload_0_22_16_real = int_reg_array_22_16_real;
  assign io_coef_out_payload_0_22_16_imag = int_reg_array_22_16_imag;
  assign io_coef_out_payload_0_22_17_real = int_reg_array_22_17_real;
  assign io_coef_out_payload_0_22_17_imag = int_reg_array_22_17_imag;
  assign io_coef_out_payload_0_22_18_real = int_reg_array_22_18_real;
  assign io_coef_out_payload_0_22_18_imag = int_reg_array_22_18_imag;
  assign io_coef_out_payload_0_22_19_real = int_reg_array_22_19_real;
  assign io_coef_out_payload_0_22_19_imag = int_reg_array_22_19_imag;
  assign io_coef_out_payload_0_22_20_real = int_reg_array_22_20_real;
  assign io_coef_out_payload_0_22_20_imag = int_reg_array_22_20_imag;
  assign io_coef_out_payload_0_22_21_real = int_reg_array_22_21_real;
  assign io_coef_out_payload_0_22_21_imag = int_reg_array_22_21_imag;
  assign io_coef_out_payload_0_22_22_real = int_reg_array_22_22_real;
  assign io_coef_out_payload_0_22_22_imag = int_reg_array_22_22_imag;
  assign io_coef_out_payload_0_22_23_real = int_reg_array_22_23_real;
  assign io_coef_out_payload_0_22_23_imag = int_reg_array_22_23_imag;
  assign io_coef_out_payload_0_22_24_real = int_reg_array_22_24_real;
  assign io_coef_out_payload_0_22_24_imag = int_reg_array_22_24_imag;
  assign io_coef_out_payload_0_22_25_real = int_reg_array_22_25_real;
  assign io_coef_out_payload_0_22_25_imag = int_reg_array_22_25_imag;
  assign io_coef_out_payload_0_22_26_real = int_reg_array_22_26_real;
  assign io_coef_out_payload_0_22_26_imag = int_reg_array_22_26_imag;
  assign io_coef_out_payload_0_22_27_real = int_reg_array_22_27_real;
  assign io_coef_out_payload_0_22_27_imag = int_reg_array_22_27_imag;
  assign io_coef_out_payload_0_22_28_real = int_reg_array_22_28_real;
  assign io_coef_out_payload_0_22_28_imag = int_reg_array_22_28_imag;
  assign io_coef_out_payload_0_22_29_real = int_reg_array_22_29_real;
  assign io_coef_out_payload_0_22_29_imag = int_reg_array_22_29_imag;
  assign io_coef_out_payload_0_22_30_real = int_reg_array_22_30_real;
  assign io_coef_out_payload_0_22_30_imag = int_reg_array_22_30_imag;
  assign io_coef_out_payload_0_22_31_real = int_reg_array_22_31_real;
  assign io_coef_out_payload_0_22_31_imag = int_reg_array_22_31_imag;
  assign io_coef_out_payload_0_22_32_real = int_reg_array_22_32_real;
  assign io_coef_out_payload_0_22_32_imag = int_reg_array_22_32_imag;
  assign io_coef_out_payload_0_22_33_real = int_reg_array_22_33_real;
  assign io_coef_out_payload_0_22_33_imag = int_reg_array_22_33_imag;
  assign io_coef_out_payload_0_22_34_real = int_reg_array_22_34_real;
  assign io_coef_out_payload_0_22_34_imag = int_reg_array_22_34_imag;
  assign io_coef_out_payload_0_22_35_real = int_reg_array_22_35_real;
  assign io_coef_out_payload_0_22_35_imag = int_reg_array_22_35_imag;
  assign io_coef_out_payload_0_22_36_real = int_reg_array_22_36_real;
  assign io_coef_out_payload_0_22_36_imag = int_reg_array_22_36_imag;
  assign io_coef_out_payload_0_22_37_real = int_reg_array_22_37_real;
  assign io_coef_out_payload_0_22_37_imag = int_reg_array_22_37_imag;
  assign io_coef_out_payload_0_22_38_real = int_reg_array_22_38_real;
  assign io_coef_out_payload_0_22_38_imag = int_reg_array_22_38_imag;
  assign io_coef_out_payload_0_22_39_real = int_reg_array_22_39_real;
  assign io_coef_out_payload_0_22_39_imag = int_reg_array_22_39_imag;
  assign io_coef_out_payload_0_22_40_real = int_reg_array_22_40_real;
  assign io_coef_out_payload_0_22_40_imag = int_reg_array_22_40_imag;
  assign io_coef_out_payload_0_22_41_real = int_reg_array_22_41_real;
  assign io_coef_out_payload_0_22_41_imag = int_reg_array_22_41_imag;
  assign io_coef_out_payload_0_22_42_real = int_reg_array_22_42_real;
  assign io_coef_out_payload_0_22_42_imag = int_reg_array_22_42_imag;
  assign io_coef_out_payload_0_22_43_real = int_reg_array_22_43_real;
  assign io_coef_out_payload_0_22_43_imag = int_reg_array_22_43_imag;
  assign io_coef_out_payload_0_22_44_real = int_reg_array_22_44_real;
  assign io_coef_out_payload_0_22_44_imag = int_reg_array_22_44_imag;
  assign io_coef_out_payload_0_22_45_real = int_reg_array_22_45_real;
  assign io_coef_out_payload_0_22_45_imag = int_reg_array_22_45_imag;
  assign io_coef_out_payload_0_22_46_real = int_reg_array_22_46_real;
  assign io_coef_out_payload_0_22_46_imag = int_reg_array_22_46_imag;
  assign io_coef_out_payload_0_22_47_real = int_reg_array_22_47_real;
  assign io_coef_out_payload_0_22_47_imag = int_reg_array_22_47_imag;
  assign io_coef_out_payload_0_22_48_real = int_reg_array_22_48_real;
  assign io_coef_out_payload_0_22_48_imag = int_reg_array_22_48_imag;
  assign io_coef_out_payload_0_22_49_real = int_reg_array_22_49_real;
  assign io_coef_out_payload_0_22_49_imag = int_reg_array_22_49_imag;
  assign io_coef_out_payload_0_23_0_real = int_reg_array_23_0_real;
  assign io_coef_out_payload_0_23_0_imag = int_reg_array_23_0_imag;
  assign io_coef_out_payload_0_23_1_real = int_reg_array_23_1_real;
  assign io_coef_out_payload_0_23_1_imag = int_reg_array_23_1_imag;
  assign io_coef_out_payload_0_23_2_real = int_reg_array_23_2_real;
  assign io_coef_out_payload_0_23_2_imag = int_reg_array_23_2_imag;
  assign io_coef_out_payload_0_23_3_real = int_reg_array_23_3_real;
  assign io_coef_out_payload_0_23_3_imag = int_reg_array_23_3_imag;
  assign io_coef_out_payload_0_23_4_real = int_reg_array_23_4_real;
  assign io_coef_out_payload_0_23_4_imag = int_reg_array_23_4_imag;
  assign io_coef_out_payload_0_23_5_real = int_reg_array_23_5_real;
  assign io_coef_out_payload_0_23_5_imag = int_reg_array_23_5_imag;
  assign io_coef_out_payload_0_23_6_real = int_reg_array_23_6_real;
  assign io_coef_out_payload_0_23_6_imag = int_reg_array_23_6_imag;
  assign io_coef_out_payload_0_23_7_real = int_reg_array_23_7_real;
  assign io_coef_out_payload_0_23_7_imag = int_reg_array_23_7_imag;
  assign io_coef_out_payload_0_23_8_real = int_reg_array_23_8_real;
  assign io_coef_out_payload_0_23_8_imag = int_reg_array_23_8_imag;
  assign io_coef_out_payload_0_23_9_real = int_reg_array_23_9_real;
  assign io_coef_out_payload_0_23_9_imag = int_reg_array_23_9_imag;
  assign io_coef_out_payload_0_23_10_real = int_reg_array_23_10_real;
  assign io_coef_out_payload_0_23_10_imag = int_reg_array_23_10_imag;
  assign io_coef_out_payload_0_23_11_real = int_reg_array_23_11_real;
  assign io_coef_out_payload_0_23_11_imag = int_reg_array_23_11_imag;
  assign io_coef_out_payload_0_23_12_real = int_reg_array_23_12_real;
  assign io_coef_out_payload_0_23_12_imag = int_reg_array_23_12_imag;
  assign io_coef_out_payload_0_23_13_real = int_reg_array_23_13_real;
  assign io_coef_out_payload_0_23_13_imag = int_reg_array_23_13_imag;
  assign io_coef_out_payload_0_23_14_real = int_reg_array_23_14_real;
  assign io_coef_out_payload_0_23_14_imag = int_reg_array_23_14_imag;
  assign io_coef_out_payload_0_23_15_real = int_reg_array_23_15_real;
  assign io_coef_out_payload_0_23_15_imag = int_reg_array_23_15_imag;
  assign io_coef_out_payload_0_23_16_real = int_reg_array_23_16_real;
  assign io_coef_out_payload_0_23_16_imag = int_reg_array_23_16_imag;
  assign io_coef_out_payload_0_23_17_real = int_reg_array_23_17_real;
  assign io_coef_out_payload_0_23_17_imag = int_reg_array_23_17_imag;
  assign io_coef_out_payload_0_23_18_real = int_reg_array_23_18_real;
  assign io_coef_out_payload_0_23_18_imag = int_reg_array_23_18_imag;
  assign io_coef_out_payload_0_23_19_real = int_reg_array_23_19_real;
  assign io_coef_out_payload_0_23_19_imag = int_reg_array_23_19_imag;
  assign io_coef_out_payload_0_23_20_real = int_reg_array_23_20_real;
  assign io_coef_out_payload_0_23_20_imag = int_reg_array_23_20_imag;
  assign io_coef_out_payload_0_23_21_real = int_reg_array_23_21_real;
  assign io_coef_out_payload_0_23_21_imag = int_reg_array_23_21_imag;
  assign io_coef_out_payload_0_23_22_real = int_reg_array_23_22_real;
  assign io_coef_out_payload_0_23_22_imag = int_reg_array_23_22_imag;
  assign io_coef_out_payload_0_23_23_real = int_reg_array_23_23_real;
  assign io_coef_out_payload_0_23_23_imag = int_reg_array_23_23_imag;
  assign io_coef_out_payload_0_23_24_real = int_reg_array_23_24_real;
  assign io_coef_out_payload_0_23_24_imag = int_reg_array_23_24_imag;
  assign io_coef_out_payload_0_23_25_real = int_reg_array_23_25_real;
  assign io_coef_out_payload_0_23_25_imag = int_reg_array_23_25_imag;
  assign io_coef_out_payload_0_23_26_real = int_reg_array_23_26_real;
  assign io_coef_out_payload_0_23_26_imag = int_reg_array_23_26_imag;
  assign io_coef_out_payload_0_23_27_real = int_reg_array_23_27_real;
  assign io_coef_out_payload_0_23_27_imag = int_reg_array_23_27_imag;
  assign io_coef_out_payload_0_23_28_real = int_reg_array_23_28_real;
  assign io_coef_out_payload_0_23_28_imag = int_reg_array_23_28_imag;
  assign io_coef_out_payload_0_23_29_real = int_reg_array_23_29_real;
  assign io_coef_out_payload_0_23_29_imag = int_reg_array_23_29_imag;
  assign io_coef_out_payload_0_23_30_real = int_reg_array_23_30_real;
  assign io_coef_out_payload_0_23_30_imag = int_reg_array_23_30_imag;
  assign io_coef_out_payload_0_23_31_real = int_reg_array_23_31_real;
  assign io_coef_out_payload_0_23_31_imag = int_reg_array_23_31_imag;
  assign io_coef_out_payload_0_23_32_real = int_reg_array_23_32_real;
  assign io_coef_out_payload_0_23_32_imag = int_reg_array_23_32_imag;
  assign io_coef_out_payload_0_23_33_real = int_reg_array_23_33_real;
  assign io_coef_out_payload_0_23_33_imag = int_reg_array_23_33_imag;
  assign io_coef_out_payload_0_23_34_real = int_reg_array_23_34_real;
  assign io_coef_out_payload_0_23_34_imag = int_reg_array_23_34_imag;
  assign io_coef_out_payload_0_23_35_real = int_reg_array_23_35_real;
  assign io_coef_out_payload_0_23_35_imag = int_reg_array_23_35_imag;
  assign io_coef_out_payload_0_23_36_real = int_reg_array_23_36_real;
  assign io_coef_out_payload_0_23_36_imag = int_reg_array_23_36_imag;
  assign io_coef_out_payload_0_23_37_real = int_reg_array_23_37_real;
  assign io_coef_out_payload_0_23_37_imag = int_reg_array_23_37_imag;
  assign io_coef_out_payload_0_23_38_real = int_reg_array_23_38_real;
  assign io_coef_out_payload_0_23_38_imag = int_reg_array_23_38_imag;
  assign io_coef_out_payload_0_23_39_real = int_reg_array_23_39_real;
  assign io_coef_out_payload_0_23_39_imag = int_reg_array_23_39_imag;
  assign io_coef_out_payload_0_23_40_real = int_reg_array_23_40_real;
  assign io_coef_out_payload_0_23_40_imag = int_reg_array_23_40_imag;
  assign io_coef_out_payload_0_23_41_real = int_reg_array_23_41_real;
  assign io_coef_out_payload_0_23_41_imag = int_reg_array_23_41_imag;
  assign io_coef_out_payload_0_23_42_real = int_reg_array_23_42_real;
  assign io_coef_out_payload_0_23_42_imag = int_reg_array_23_42_imag;
  assign io_coef_out_payload_0_23_43_real = int_reg_array_23_43_real;
  assign io_coef_out_payload_0_23_43_imag = int_reg_array_23_43_imag;
  assign io_coef_out_payload_0_23_44_real = int_reg_array_23_44_real;
  assign io_coef_out_payload_0_23_44_imag = int_reg_array_23_44_imag;
  assign io_coef_out_payload_0_23_45_real = int_reg_array_23_45_real;
  assign io_coef_out_payload_0_23_45_imag = int_reg_array_23_45_imag;
  assign io_coef_out_payload_0_23_46_real = int_reg_array_23_46_real;
  assign io_coef_out_payload_0_23_46_imag = int_reg_array_23_46_imag;
  assign io_coef_out_payload_0_23_47_real = int_reg_array_23_47_real;
  assign io_coef_out_payload_0_23_47_imag = int_reg_array_23_47_imag;
  assign io_coef_out_payload_0_23_48_real = int_reg_array_23_48_real;
  assign io_coef_out_payload_0_23_48_imag = int_reg_array_23_48_imag;
  assign io_coef_out_payload_0_23_49_real = int_reg_array_23_49_real;
  assign io_coef_out_payload_0_23_49_imag = int_reg_array_23_49_imag;
  assign io_coef_out_payload_0_24_0_real = int_reg_array_24_0_real;
  assign io_coef_out_payload_0_24_0_imag = int_reg_array_24_0_imag;
  assign io_coef_out_payload_0_24_1_real = int_reg_array_24_1_real;
  assign io_coef_out_payload_0_24_1_imag = int_reg_array_24_1_imag;
  assign io_coef_out_payload_0_24_2_real = int_reg_array_24_2_real;
  assign io_coef_out_payload_0_24_2_imag = int_reg_array_24_2_imag;
  assign io_coef_out_payload_0_24_3_real = int_reg_array_24_3_real;
  assign io_coef_out_payload_0_24_3_imag = int_reg_array_24_3_imag;
  assign io_coef_out_payload_0_24_4_real = int_reg_array_24_4_real;
  assign io_coef_out_payload_0_24_4_imag = int_reg_array_24_4_imag;
  assign io_coef_out_payload_0_24_5_real = int_reg_array_24_5_real;
  assign io_coef_out_payload_0_24_5_imag = int_reg_array_24_5_imag;
  assign io_coef_out_payload_0_24_6_real = int_reg_array_24_6_real;
  assign io_coef_out_payload_0_24_6_imag = int_reg_array_24_6_imag;
  assign io_coef_out_payload_0_24_7_real = int_reg_array_24_7_real;
  assign io_coef_out_payload_0_24_7_imag = int_reg_array_24_7_imag;
  assign io_coef_out_payload_0_24_8_real = int_reg_array_24_8_real;
  assign io_coef_out_payload_0_24_8_imag = int_reg_array_24_8_imag;
  assign io_coef_out_payload_0_24_9_real = int_reg_array_24_9_real;
  assign io_coef_out_payload_0_24_9_imag = int_reg_array_24_9_imag;
  assign io_coef_out_payload_0_24_10_real = int_reg_array_24_10_real;
  assign io_coef_out_payload_0_24_10_imag = int_reg_array_24_10_imag;
  assign io_coef_out_payload_0_24_11_real = int_reg_array_24_11_real;
  assign io_coef_out_payload_0_24_11_imag = int_reg_array_24_11_imag;
  assign io_coef_out_payload_0_24_12_real = int_reg_array_24_12_real;
  assign io_coef_out_payload_0_24_12_imag = int_reg_array_24_12_imag;
  assign io_coef_out_payload_0_24_13_real = int_reg_array_24_13_real;
  assign io_coef_out_payload_0_24_13_imag = int_reg_array_24_13_imag;
  assign io_coef_out_payload_0_24_14_real = int_reg_array_24_14_real;
  assign io_coef_out_payload_0_24_14_imag = int_reg_array_24_14_imag;
  assign io_coef_out_payload_0_24_15_real = int_reg_array_24_15_real;
  assign io_coef_out_payload_0_24_15_imag = int_reg_array_24_15_imag;
  assign io_coef_out_payload_0_24_16_real = int_reg_array_24_16_real;
  assign io_coef_out_payload_0_24_16_imag = int_reg_array_24_16_imag;
  assign io_coef_out_payload_0_24_17_real = int_reg_array_24_17_real;
  assign io_coef_out_payload_0_24_17_imag = int_reg_array_24_17_imag;
  assign io_coef_out_payload_0_24_18_real = int_reg_array_24_18_real;
  assign io_coef_out_payload_0_24_18_imag = int_reg_array_24_18_imag;
  assign io_coef_out_payload_0_24_19_real = int_reg_array_24_19_real;
  assign io_coef_out_payload_0_24_19_imag = int_reg_array_24_19_imag;
  assign io_coef_out_payload_0_24_20_real = int_reg_array_24_20_real;
  assign io_coef_out_payload_0_24_20_imag = int_reg_array_24_20_imag;
  assign io_coef_out_payload_0_24_21_real = int_reg_array_24_21_real;
  assign io_coef_out_payload_0_24_21_imag = int_reg_array_24_21_imag;
  assign io_coef_out_payload_0_24_22_real = int_reg_array_24_22_real;
  assign io_coef_out_payload_0_24_22_imag = int_reg_array_24_22_imag;
  assign io_coef_out_payload_0_24_23_real = int_reg_array_24_23_real;
  assign io_coef_out_payload_0_24_23_imag = int_reg_array_24_23_imag;
  assign io_coef_out_payload_0_24_24_real = int_reg_array_24_24_real;
  assign io_coef_out_payload_0_24_24_imag = int_reg_array_24_24_imag;
  assign io_coef_out_payload_0_24_25_real = int_reg_array_24_25_real;
  assign io_coef_out_payload_0_24_25_imag = int_reg_array_24_25_imag;
  assign io_coef_out_payload_0_24_26_real = int_reg_array_24_26_real;
  assign io_coef_out_payload_0_24_26_imag = int_reg_array_24_26_imag;
  assign io_coef_out_payload_0_24_27_real = int_reg_array_24_27_real;
  assign io_coef_out_payload_0_24_27_imag = int_reg_array_24_27_imag;
  assign io_coef_out_payload_0_24_28_real = int_reg_array_24_28_real;
  assign io_coef_out_payload_0_24_28_imag = int_reg_array_24_28_imag;
  assign io_coef_out_payload_0_24_29_real = int_reg_array_24_29_real;
  assign io_coef_out_payload_0_24_29_imag = int_reg_array_24_29_imag;
  assign io_coef_out_payload_0_24_30_real = int_reg_array_24_30_real;
  assign io_coef_out_payload_0_24_30_imag = int_reg_array_24_30_imag;
  assign io_coef_out_payload_0_24_31_real = int_reg_array_24_31_real;
  assign io_coef_out_payload_0_24_31_imag = int_reg_array_24_31_imag;
  assign io_coef_out_payload_0_24_32_real = int_reg_array_24_32_real;
  assign io_coef_out_payload_0_24_32_imag = int_reg_array_24_32_imag;
  assign io_coef_out_payload_0_24_33_real = int_reg_array_24_33_real;
  assign io_coef_out_payload_0_24_33_imag = int_reg_array_24_33_imag;
  assign io_coef_out_payload_0_24_34_real = int_reg_array_24_34_real;
  assign io_coef_out_payload_0_24_34_imag = int_reg_array_24_34_imag;
  assign io_coef_out_payload_0_24_35_real = int_reg_array_24_35_real;
  assign io_coef_out_payload_0_24_35_imag = int_reg_array_24_35_imag;
  assign io_coef_out_payload_0_24_36_real = int_reg_array_24_36_real;
  assign io_coef_out_payload_0_24_36_imag = int_reg_array_24_36_imag;
  assign io_coef_out_payload_0_24_37_real = int_reg_array_24_37_real;
  assign io_coef_out_payload_0_24_37_imag = int_reg_array_24_37_imag;
  assign io_coef_out_payload_0_24_38_real = int_reg_array_24_38_real;
  assign io_coef_out_payload_0_24_38_imag = int_reg_array_24_38_imag;
  assign io_coef_out_payload_0_24_39_real = int_reg_array_24_39_real;
  assign io_coef_out_payload_0_24_39_imag = int_reg_array_24_39_imag;
  assign io_coef_out_payload_0_24_40_real = int_reg_array_24_40_real;
  assign io_coef_out_payload_0_24_40_imag = int_reg_array_24_40_imag;
  assign io_coef_out_payload_0_24_41_real = int_reg_array_24_41_real;
  assign io_coef_out_payload_0_24_41_imag = int_reg_array_24_41_imag;
  assign io_coef_out_payload_0_24_42_real = int_reg_array_24_42_real;
  assign io_coef_out_payload_0_24_42_imag = int_reg_array_24_42_imag;
  assign io_coef_out_payload_0_24_43_real = int_reg_array_24_43_real;
  assign io_coef_out_payload_0_24_43_imag = int_reg_array_24_43_imag;
  assign io_coef_out_payload_0_24_44_real = int_reg_array_24_44_real;
  assign io_coef_out_payload_0_24_44_imag = int_reg_array_24_44_imag;
  assign io_coef_out_payload_0_24_45_real = int_reg_array_24_45_real;
  assign io_coef_out_payload_0_24_45_imag = int_reg_array_24_45_imag;
  assign io_coef_out_payload_0_24_46_real = int_reg_array_24_46_real;
  assign io_coef_out_payload_0_24_46_imag = int_reg_array_24_46_imag;
  assign io_coef_out_payload_0_24_47_real = int_reg_array_24_47_real;
  assign io_coef_out_payload_0_24_47_imag = int_reg_array_24_47_imag;
  assign io_coef_out_payload_0_24_48_real = int_reg_array_24_48_real;
  assign io_coef_out_payload_0_24_48_imag = int_reg_array_24_48_imag;
  assign io_coef_out_payload_0_24_49_real = int_reg_array_24_49_real;
  assign io_coef_out_payload_0_24_49_imag = int_reg_array_24_49_imag;
  assign io_coef_out_payload_0_25_0_real = int_reg_array_25_0_real;
  assign io_coef_out_payload_0_25_0_imag = int_reg_array_25_0_imag;
  assign io_coef_out_payload_0_25_1_real = int_reg_array_25_1_real;
  assign io_coef_out_payload_0_25_1_imag = int_reg_array_25_1_imag;
  assign io_coef_out_payload_0_25_2_real = int_reg_array_25_2_real;
  assign io_coef_out_payload_0_25_2_imag = int_reg_array_25_2_imag;
  assign io_coef_out_payload_0_25_3_real = int_reg_array_25_3_real;
  assign io_coef_out_payload_0_25_3_imag = int_reg_array_25_3_imag;
  assign io_coef_out_payload_0_25_4_real = int_reg_array_25_4_real;
  assign io_coef_out_payload_0_25_4_imag = int_reg_array_25_4_imag;
  assign io_coef_out_payload_0_25_5_real = int_reg_array_25_5_real;
  assign io_coef_out_payload_0_25_5_imag = int_reg_array_25_5_imag;
  assign io_coef_out_payload_0_25_6_real = int_reg_array_25_6_real;
  assign io_coef_out_payload_0_25_6_imag = int_reg_array_25_6_imag;
  assign io_coef_out_payload_0_25_7_real = int_reg_array_25_7_real;
  assign io_coef_out_payload_0_25_7_imag = int_reg_array_25_7_imag;
  assign io_coef_out_payload_0_25_8_real = int_reg_array_25_8_real;
  assign io_coef_out_payload_0_25_8_imag = int_reg_array_25_8_imag;
  assign io_coef_out_payload_0_25_9_real = int_reg_array_25_9_real;
  assign io_coef_out_payload_0_25_9_imag = int_reg_array_25_9_imag;
  assign io_coef_out_payload_0_25_10_real = int_reg_array_25_10_real;
  assign io_coef_out_payload_0_25_10_imag = int_reg_array_25_10_imag;
  assign io_coef_out_payload_0_25_11_real = int_reg_array_25_11_real;
  assign io_coef_out_payload_0_25_11_imag = int_reg_array_25_11_imag;
  assign io_coef_out_payload_0_25_12_real = int_reg_array_25_12_real;
  assign io_coef_out_payload_0_25_12_imag = int_reg_array_25_12_imag;
  assign io_coef_out_payload_0_25_13_real = int_reg_array_25_13_real;
  assign io_coef_out_payload_0_25_13_imag = int_reg_array_25_13_imag;
  assign io_coef_out_payload_0_25_14_real = int_reg_array_25_14_real;
  assign io_coef_out_payload_0_25_14_imag = int_reg_array_25_14_imag;
  assign io_coef_out_payload_0_25_15_real = int_reg_array_25_15_real;
  assign io_coef_out_payload_0_25_15_imag = int_reg_array_25_15_imag;
  assign io_coef_out_payload_0_25_16_real = int_reg_array_25_16_real;
  assign io_coef_out_payload_0_25_16_imag = int_reg_array_25_16_imag;
  assign io_coef_out_payload_0_25_17_real = int_reg_array_25_17_real;
  assign io_coef_out_payload_0_25_17_imag = int_reg_array_25_17_imag;
  assign io_coef_out_payload_0_25_18_real = int_reg_array_25_18_real;
  assign io_coef_out_payload_0_25_18_imag = int_reg_array_25_18_imag;
  assign io_coef_out_payload_0_25_19_real = int_reg_array_25_19_real;
  assign io_coef_out_payload_0_25_19_imag = int_reg_array_25_19_imag;
  assign io_coef_out_payload_0_25_20_real = int_reg_array_25_20_real;
  assign io_coef_out_payload_0_25_20_imag = int_reg_array_25_20_imag;
  assign io_coef_out_payload_0_25_21_real = int_reg_array_25_21_real;
  assign io_coef_out_payload_0_25_21_imag = int_reg_array_25_21_imag;
  assign io_coef_out_payload_0_25_22_real = int_reg_array_25_22_real;
  assign io_coef_out_payload_0_25_22_imag = int_reg_array_25_22_imag;
  assign io_coef_out_payload_0_25_23_real = int_reg_array_25_23_real;
  assign io_coef_out_payload_0_25_23_imag = int_reg_array_25_23_imag;
  assign io_coef_out_payload_0_25_24_real = int_reg_array_25_24_real;
  assign io_coef_out_payload_0_25_24_imag = int_reg_array_25_24_imag;
  assign io_coef_out_payload_0_25_25_real = int_reg_array_25_25_real;
  assign io_coef_out_payload_0_25_25_imag = int_reg_array_25_25_imag;
  assign io_coef_out_payload_0_25_26_real = int_reg_array_25_26_real;
  assign io_coef_out_payload_0_25_26_imag = int_reg_array_25_26_imag;
  assign io_coef_out_payload_0_25_27_real = int_reg_array_25_27_real;
  assign io_coef_out_payload_0_25_27_imag = int_reg_array_25_27_imag;
  assign io_coef_out_payload_0_25_28_real = int_reg_array_25_28_real;
  assign io_coef_out_payload_0_25_28_imag = int_reg_array_25_28_imag;
  assign io_coef_out_payload_0_25_29_real = int_reg_array_25_29_real;
  assign io_coef_out_payload_0_25_29_imag = int_reg_array_25_29_imag;
  assign io_coef_out_payload_0_25_30_real = int_reg_array_25_30_real;
  assign io_coef_out_payload_0_25_30_imag = int_reg_array_25_30_imag;
  assign io_coef_out_payload_0_25_31_real = int_reg_array_25_31_real;
  assign io_coef_out_payload_0_25_31_imag = int_reg_array_25_31_imag;
  assign io_coef_out_payload_0_25_32_real = int_reg_array_25_32_real;
  assign io_coef_out_payload_0_25_32_imag = int_reg_array_25_32_imag;
  assign io_coef_out_payload_0_25_33_real = int_reg_array_25_33_real;
  assign io_coef_out_payload_0_25_33_imag = int_reg_array_25_33_imag;
  assign io_coef_out_payload_0_25_34_real = int_reg_array_25_34_real;
  assign io_coef_out_payload_0_25_34_imag = int_reg_array_25_34_imag;
  assign io_coef_out_payload_0_25_35_real = int_reg_array_25_35_real;
  assign io_coef_out_payload_0_25_35_imag = int_reg_array_25_35_imag;
  assign io_coef_out_payload_0_25_36_real = int_reg_array_25_36_real;
  assign io_coef_out_payload_0_25_36_imag = int_reg_array_25_36_imag;
  assign io_coef_out_payload_0_25_37_real = int_reg_array_25_37_real;
  assign io_coef_out_payload_0_25_37_imag = int_reg_array_25_37_imag;
  assign io_coef_out_payload_0_25_38_real = int_reg_array_25_38_real;
  assign io_coef_out_payload_0_25_38_imag = int_reg_array_25_38_imag;
  assign io_coef_out_payload_0_25_39_real = int_reg_array_25_39_real;
  assign io_coef_out_payload_0_25_39_imag = int_reg_array_25_39_imag;
  assign io_coef_out_payload_0_25_40_real = int_reg_array_25_40_real;
  assign io_coef_out_payload_0_25_40_imag = int_reg_array_25_40_imag;
  assign io_coef_out_payload_0_25_41_real = int_reg_array_25_41_real;
  assign io_coef_out_payload_0_25_41_imag = int_reg_array_25_41_imag;
  assign io_coef_out_payload_0_25_42_real = int_reg_array_25_42_real;
  assign io_coef_out_payload_0_25_42_imag = int_reg_array_25_42_imag;
  assign io_coef_out_payload_0_25_43_real = int_reg_array_25_43_real;
  assign io_coef_out_payload_0_25_43_imag = int_reg_array_25_43_imag;
  assign io_coef_out_payload_0_25_44_real = int_reg_array_25_44_real;
  assign io_coef_out_payload_0_25_44_imag = int_reg_array_25_44_imag;
  assign io_coef_out_payload_0_25_45_real = int_reg_array_25_45_real;
  assign io_coef_out_payload_0_25_45_imag = int_reg_array_25_45_imag;
  assign io_coef_out_payload_0_25_46_real = int_reg_array_25_46_real;
  assign io_coef_out_payload_0_25_46_imag = int_reg_array_25_46_imag;
  assign io_coef_out_payload_0_25_47_real = int_reg_array_25_47_real;
  assign io_coef_out_payload_0_25_47_imag = int_reg_array_25_47_imag;
  assign io_coef_out_payload_0_25_48_real = int_reg_array_25_48_real;
  assign io_coef_out_payload_0_25_48_imag = int_reg_array_25_48_imag;
  assign io_coef_out_payload_0_25_49_real = int_reg_array_25_49_real;
  assign io_coef_out_payload_0_25_49_imag = int_reg_array_25_49_imag;
  assign io_coef_out_payload_0_26_0_real = int_reg_array_26_0_real;
  assign io_coef_out_payload_0_26_0_imag = int_reg_array_26_0_imag;
  assign io_coef_out_payload_0_26_1_real = int_reg_array_26_1_real;
  assign io_coef_out_payload_0_26_1_imag = int_reg_array_26_1_imag;
  assign io_coef_out_payload_0_26_2_real = int_reg_array_26_2_real;
  assign io_coef_out_payload_0_26_2_imag = int_reg_array_26_2_imag;
  assign io_coef_out_payload_0_26_3_real = int_reg_array_26_3_real;
  assign io_coef_out_payload_0_26_3_imag = int_reg_array_26_3_imag;
  assign io_coef_out_payload_0_26_4_real = int_reg_array_26_4_real;
  assign io_coef_out_payload_0_26_4_imag = int_reg_array_26_4_imag;
  assign io_coef_out_payload_0_26_5_real = int_reg_array_26_5_real;
  assign io_coef_out_payload_0_26_5_imag = int_reg_array_26_5_imag;
  assign io_coef_out_payload_0_26_6_real = int_reg_array_26_6_real;
  assign io_coef_out_payload_0_26_6_imag = int_reg_array_26_6_imag;
  assign io_coef_out_payload_0_26_7_real = int_reg_array_26_7_real;
  assign io_coef_out_payload_0_26_7_imag = int_reg_array_26_7_imag;
  assign io_coef_out_payload_0_26_8_real = int_reg_array_26_8_real;
  assign io_coef_out_payload_0_26_8_imag = int_reg_array_26_8_imag;
  assign io_coef_out_payload_0_26_9_real = int_reg_array_26_9_real;
  assign io_coef_out_payload_0_26_9_imag = int_reg_array_26_9_imag;
  assign io_coef_out_payload_0_26_10_real = int_reg_array_26_10_real;
  assign io_coef_out_payload_0_26_10_imag = int_reg_array_26_10_imag;
  assign io_coef_out_payload_0_26_11_real = int_reg_array_26_11_real;
  assign io_coef_out_payload_0_26_11_imag = int_reg_array_26_11_imag;
  assign io_coef_out_payload_0_26_12_real = int_reg_array_26_12_real;
  assign io_coef_out_payload_0_26_12_imag = int_reg_array_26_12_imag;
  assign io_coef_out_payload_0_26_13_real = int_reg_array_26_13_real;
  assign io_coef_out_payload_0_26_13_imag = int_reg_array_26_13_imag;
  assign io_coef_out_payload_0_26_14_real = int_reg_array_26_14_real;
  assign io_coef_out_payload_0_26_14_imag = int_reg_array_26_14_imag;
  assign io_coef_out_payload_0_26_15_real = int_reg_array_26_15_real;
  assign io_coef_out_payload_0_26_15_imag = int_reg_array_26_15_imag;
  assign io_coef_out_payload_0_26_16_real = int_reg_array_26_16_real;
  assign io_coef_out_payload_0_26_16_imag = int_reg_array_26_16_imag;
  assign io_coef_out_payload_0_26_17_real = int_reg_array_26_17_real;
  assign io_coef_out_payload_0_26_17_imag = int_reg_array_26_17_imag;
  assign io_coef_out_payload_0_26_18_real = int_reg_array_26_18_real;
  assign io_coef_out_payload_0_26_18_imag = int_reg_array_26_18_imag;
  assign io_coef_out_payload_0_26_19_real = int_reg_array_26_19_real;
  assign io_coef_out_payload_0_26_19_imag = int_reg_array_26_19_imag;
  assign io_coef_out_payload_0_26_20_real = int_reg_array_26_20_real;
  assign io_coef_out_payload_0_26_20_imag = int_reg_array_26_20_imag;
  assign io_coef_out_payload_0_26_21_real = int_reg_array_26_21_real;
  assign io_coef_out_payload_0_26_21_imag = int_reg_array_26_21_imag;
  assign io_coef_out_payload_0_26_22_real = int_reg_array_26_22_real;
  assign io_coef_out_payload_0_26_22_imag = int_reg_array_26_22_imag;
  assign io_coef_out_payload_0_26_23_real = int_reg_array_26_23_real;
  assign io_coef_out_payload_0_26_23_imag = int_reg_array_26_23_imag;
  assign io_coef_out_payload_0_26_24_real = int_reg_array_26_24_real;
  assign io_coef_out_payload_0_26_24_imag = int_reg_array_26_24_imag;
  assign io_coef_out_payload_0_26_25_real = int_reg_array_26_25_real;
  assign io_coef_out_payload_0_26_25_imag = int_reg_array_26_25_imag;
  assign io_coef_out_payload_0_26_26_real = int_reg_array_26_26_real;
  assign io_coef_out_payload_0_26_26_imag = int_reg_array_26_26_imag;
  assign io_coef_out_payload_0_26_27_real = int_reg_array_26_27_real;
  assign io_coef_out_payload_0_26_27_imag = int_reg_array_26_27_imag;
  assign io_coef_out_payload_0_26_28_real = int_reg_array_26_28_real;
  assign io_coef_out_payload_0_26_28_imag = int_reg_array_26_28_imag;
  assign io_coef_out_payload_0_26_29_real = int_reg_array_26_29_real;
  assign io_coef_out_payload_0_26_29_imag = int_reg_array_26_29_imag;
  assign io_coef_out_payload_0_26_30_real = int_reg_array_26_30_real;
  assign io_coef_out_payload_0_26_30_imag = int_reg_array_26_30_imag;
  assign io_coef_out_payload_0_26_31_real = int_reg_array_26_31_real;
  assign io_coef_out_payload_0_26_31_imag = int_reg_array_26_31_imag;
  assign io_coef_out_payload_0_26_32_real = int_reg_array_26_32_real;
  assign io_coef_out_payload_0_26_32_imag = int_reg_array_26_32_imag;
  assign io_coef_out_payload_0_26_33_real = int_reg_array_26_33_real;
  assign io_coef_out_payload_0_26_33_imag = int_reg_array_26_33_imag;
  assign io_coef_out_payload_0_26_34_real = int_reg_array_26_34_real;
  assign io_coef_out_payload_0_26_34_imag = int_reg_array_26_34_imag;
  assign io_coef_out_payload_0_26_35_real = int_reg_array_26_35_real;
  assign io_coef_out_payload_0_26_35_imag = int_reg_array_26_35_imag;
  assign io_coef_out_payload_0_26_36_real = int_reg_array_26_36_real;
  assign io_coef_out_payload_0_26_36_imag = int_reg_array_26_36_imag;
  assign io_coef_out_payload_0_26_37_real = int_reg_array_26_37_real;
  assign io_coef_out_payload_0_26_37_imag = int_reg_array_26_37_imag;
  assign io_coef_out_payload_0_26_38_real = int_reg_array_26_38_real;
  assign io_coef_out_payload_0_26_38_imag = int_reg_array_26_38_imag;
  assign io_coef_out_payload_0_26_39_real = int_reg_array_26_39_real;
  assign io_coef_out_payload_0_26_39_imag = int_reg_array_26_39_imag;
  assign io_coef_out_payload_0_26_40_real = int_reg_array_26_40_real;
  assign io_coef_out_payload_0_26_40_imag = int_reg_array_26_40_imag;
  assign io_coef_out_payload_0_26_41_real = int_reg_array_26_41_real;
  assign io_coef_out_payload_0_26_41_imag = int_reg_array_26_41_imag;
  assign io_coef_out_payload_0_26_42_real = int_reg_array_26_42_real;
  assign io_coef_out_payload_0_26_42_imag = int_reg_array_26_42_imag;
  assign io_coef_out_payload_0_26_43_real = int_reg_array_26_43_real;
  assign io_coef_out_payload_0_26_43_imag = int_reg_array_26_43_imag;
  assign io_coef_out_payload_0_26_44_real = int_reg_array_26_44_real;
  assign io_coef_out_payload_0_26_44_imag = int_reg_array_26_44_imag;
  assign io_coef_out_payload_0_26_45_real = int_reg_array_26_45_real;
  assign io_coef_out_payload_0_26_45_imag = int_reg_array_26_45_imag;
  assign io_coef_out_payload_0_26_46_real = int_reg_array_26_46_real;
  assign io_coef_out_payload_0_26_46_imag = int_reg_array_26_46_imag;
  assign io_coef_out_payload_0_26_47_real = int_reg_array_26_47_real;
  assign io_coef_out_payload_0_26_47_imag = int_reg_array_26_47_imag;
  assign io_coef_out_payload_0_26_48_real = int_reg_array_26_48_real;
  assign io_coef_out_payload_0_26_48_imag = int_reg_array_26_48_imag;
  assign io_coef_out_payload_0_26_49_real = int_reg_array_26_49_real;
  assign io_coef_out_payload_0_26_49_imag = int_reg_array_26_49_imag;
  assign io_coef_out_payload_0_27_0_real = int_reg_array_27_0_real;
  assign io_coef_out_payload_0_27_0_imag = int_reg_array_27_0_imag;
  assign io_coef_out_payload_0_27_1_real = int_reg_array_27_1_real;
  assign io_coef_out_payload_0_27_1_imag = int_reg_array_27_1_imag;
  assign io_coef_out_payload_0_27_2_real = int_reg_array_27_2_real;
  assign io_coef_out_payload_0_27_2_imag = int_reg_array_27_2_imag;
  assign io_coef_out_payload_0_27_3_real = int_reg_array_27_3_real;
  assign io_coef_out_payload_0_27_3_imag = int_reg_array_27_3_imag;
  assign io_coef_out_payload_0_27_4_real = int_reg_array_27_4_real;
  assign io_coef_out_payload_0_27_4_imag = int_reg_array_27_4_imag;
  assign io_coef_out_payload_0_27_5_real = int_reg_array_27_5_real;
  assign io_coef_out_payload_0_27_5_imag = int_reg_array_27_5_imag;
  assign io_coef_out_payload_0_27_6_real = int_reg_array_27_6_real;
  assign io_coef_out_payload_0_27_6_imag = int_reg_array_27_6_imag;
  assign io_coef_out_payload_0_27_7_real = int_reg_array_27_7_real;
  assign io_coef_out_payload_0_27_7_imag = int_reg_array_27_7_imag;
  assign io_coef_out_payload_0_27_8_real = int_reg_array_27_8_real;
  assign io_coef_out_payload_0_27_8_imag = int_reg_array_27_8_imag;
  assign io_coef_out_payload_0_27_9_real = int_reg_array_27_9_real;
  assign io_coef_out_payload_0_27_9_imag = int_reg_array_27_9_imag;
  assign io_coef_out_payload_0_27_10_real = int_reg_array_27_10_real;
  assign io_coef_out_payload_0_27_10_imag = int_reg_array_27_10_imag;
  assign io_coef_out_payload_0_27_11_real = int_reg_array_27_11_real;
  assign io_coef_out_payload_0_27_11_imag = int_reg_array_27_11_imag;
  assign io_coef_out_payload_0_27_12_real = int_reg_array_27_12_real;
  assign io_coef_out_payload_0_27_12_imag = int_reg_array_27_12_imag;
  assign io_coef_out_payload_0_27_13_real = int_reg_array_27_13_real;
  assign io_coef_out_payload_0_27_13_imag = int_reg_array_27_13_imag;
  assign io_coef_out_payload_0_27_14_real = int_reg_array_27_14_real;
  assign io_coef_out_payload_0_27_14_imag = int_reg_array_27_14_imag;
  assign io_coef_out_payload_0_27_15_real = int_reg_array_27_15_real;
  assign io_coef_out_payload_0_27_15_imag = int_reg_array_27_15_imag;
  assign io_coef_out_payload_0_27_16_real = int_reg_array_27_16_real;
  assign io_coef_out_payload_0_27_16_imag = int_reg_array_27_16_imag;
  assign io_coef_out_payload_0_27_17_real = int_reg_array_27_17_real;
  assign io_coef_out_payload_0_27_17_imag = int_reg_array_27_17_imag;
  assign io_coef_out_payload_0_27_18_real = int_reg_array_27_18_real;
  assign io_coef_out_payload_0_27_18_imag = int_reg_array_27_18_imag;
  assign io_coef_out_payload_0_27_19_real = int_reg_array_27_19_real;
  assign io_coef_out_payload_0_27_19_imag = int_reg_array_27_19_imag;
  assign io_coef_out_payload_0_27_20_real = int_reg_array_27_20_real;
  assign io_coef_out_payload_0_27_20_imag = int_reg_array_27_20_imag;
  assign io_coef_out_payload_0_27_21_real = int_reg_array_27_21_real;
  assign io_coef_out_payload_0_27_21_imag = int_reg_array_27_21_imag;
  assign io_coef_out_payload_0_27_22_real = int_reg_array_27_22_real;
  assign io_coef_out_payload_0_27_22_imag = int_reg_array_27_22_imag;
  assign io_coef_out_payload_0_27_23_real = int_reg_array_27_23_real;
  assign io_coef_out_payload_0_27_23_imag = int_reg_array_27_23_imag;
  assign io_coef_out_payload_0_27_24_real = int_reg_array_27_24_real;
  assign io_coef_out_payload_0_27_24_imag = int_reg_array_27_24_imag;
  assign io_coef_out_payload_0_27_25_real = int_reg_array_27_25_real;
  assign io_coef_out_payload_0_27_25_imag = int_reg_array_27_25_imag;
  assign io_coef_out_payload_0_27_26_real = int_reg_array_27_26_real;
  assign io_coef_out_payload_0_27_26_imag = int_reg_array_27_26_imag;
  assign io_coef_out_payload_0_27_27_real = int_reg_array_27_27_real;
  assign io_coef_out_payload_0_27_27_imag = int_reg_array_27_27_imag;
  assign io_coef_out_payload_0_27_28_real = int_reg_array_27_28_real;
  assign io_coef_out_payload_0_27_28_imag = int_reg_array_27_28_imag;
  assign io_coef_out_payload_0_27_29_real = int_reg_array_27_29_real;
  assign io_coef_out_payload_0_27_29_imag = int_reg_array_27_29_imag;
  assign io_coef_out_payload_0_27_30_real = int_reg_array_27_30_real;
  assign io_coef_out_payload_0_27_30_imag = int_reg_array_27_30_imag;
  assign io_coef_out_payload_0_27_31_real = int_reg_array_27_31_real;
  assign io_coef_out_payload_0_27_31_imag = int_reg_array_27_31_imag;
  assign io_coef_out_payload_0_27_32_real = int_reg_array_27_32_real;
  assign io_coef_out_payload_0_27_32_imag = int_reg_array_27_32_imag;
  assign io_coef_out_payload_0_27_33_real = int_reg_array_27_33_real;
  assign io_coef_out_payload_0_27_33_imag = int_reg_array_27_33_imag;
  assign io_coef_out_payload_0_27_34_real = int_reg_array_27_34_real;
  assign io_coef_out_payload_0_27_34_imag = int_reg_array_27_34_imag;
  assign io_coef_out_payload_0_27_35_real = int_reg_array_27_35_real;
  assign io_coef_out_payload_0_27_35_imag = int_reg_array_27_35_imag;
  assign io_coef_out_payload_0_27_36_real = int_reg_array_27_36_real;
  assign io_coef_out_payload_0_27_36_imag = int_reg_array_27_36_imag;
  assign io_coef_out_payload_0_27_37_real = int_reg_array_27_37_real;
  assign io_coef_out_payload_0_27_37_imag = int_reg_array_27_37_imag;
  assign io_coef_out_payload_0_27_38_real = int_reg_array_27_38_real;
  assign io_coef_out_payload_0_27_38_imag = int_reg_array_27_38_imag;
  assign io_coef_out_payload_0_27_39_real = int_reg_array_27_39_real;
  assign io_coef_out_payload_0_27_39_imag = int_reg_array_27_39_imag;
  assign io_coef_out_payload_0_27_40_real = int_reg_array_27_40_real;
  assign io_coef_out_payload_0_27_40_imag = int_reg_array_27_40_imag;
  assign io_coef_out_payload_0_27_41_real = int_reg_array_27_41_real;
  assign io_coef_out_payload_0_27_41_imag = int_reg_array_27_41_imag;
  assign io_coef_out_payload_0_27_42_real = int_reg_array_27_42_real;
  assign io_coef_out_payload_0_27_42_imag = int_reg_array_27_42_imag;
  assign io_coef_out_payload_0_27_43_real = int_reg_array_27_43_real;
  assign io_coef_out_payload_0_27_43_imag = int_reg_array_27_43_imag;
  assign io_coef_out_payload_0_27_44_real = int_reg_array_27_44_real;
  assign io_coef_out_payload_0_27_44_imag = int_reg_array_27_44_imag;
  assign io_coef_out_payload_0_27_45_real = int_reg_array_27_45_real;
  assign io_coef_out_payload_0_27_45_imag = int_reg_array_27_45_imag;
  assign io_coef_out_payload_0_27_46_real = int_reg_array_27_46_real;
  assign io_coef_out_payload_0_27_46_imag = int_reg_array_27_46_imag;
  assign io_coef_out_payload_0_27_47_real = int_reg_array_27_47_real;
  assign io_coef_out_payload_0_27_47_imag = int_reg_array_27_47_imag;
  assign io_coef_out_payload_0_27_48_real = int_reg_array_27_48_real;
  assign io_coef_out_payload_0_27_48_imag = int_reg_array_27_48_imag;
  assign io_coef_out_payload_0_27_49_real = int_reg_array_27_49_real;
  assign io_coef_out_payload_0_27_49_imag = int_reg_array_27_49_imag;
  assign io_coef_out_payload_0_28_0_real = int_reg_array_28_0_real;
  assign io_coef_out_payload_0_28_0_imag = int_reg_array_28_0_imag;
  assign io_coef_out_payload_0_28_1_real = int_reg_array_28_1_real;
  assign io_coef_out_payload_0_28_1_imag = int_reg_array_28_1_imag;
  assign io_coef_out_payload_0_28_2_real = int_reg_array_28_2_real;
  assign io_coef_out_payload_0_28_2_imag = int_reg_array_28_2_imag;
  assign io_coef_out_payload_0_28_3_real = int_reg_array_28_3_real;
  assign io_coef_out_payload_0_28_3_imag = int_reg_array_28_3_imag;
  assign io_coef_out_payload_0_28_4_real = int_reg_array_28_4_real;
  assign io_coef_out_payload_0_28_4_imag = int_reg_array_28_4_imag;
  assign io_coef_out_payload_0_28_5_real = int_reg_array_28_5_real;
  assign io_coef_out_payload_0_28_5_imag = int_reg_array_28_5_imag;
  assign io_coef_out_payload_0_28_6_real = int_reg_array_28_6_real;
  assign io_coef_out_payload_0_28_6_imag = int_reg_array_28_6_imag;
  assign io_coef_out_payload_0_28_7_real = int_reg_array_28_7_real;
  assign io_coef_out_payload_0_28_7_imag = int_reg_array_28_7_imag;
  assign io_coef_out_payload_0_28_8_real = int_reg_array_28_8_real;
  assign io_coef_out_payload_0_28_8_imag = int_reg_array_28_8_imag;
  assign io_coef_out_payload_0_28_9_real = int_reg_array_28_9_real;
  assign io_coef_out_payload_0_28_9_imag = int_reg_array_28_9_imag;
  assign io_coef_out_payload_0_28_10_real = int_reg_array_28_10_real;
  assign io_coef_out_payload_0_28_10_imag = int_reg_array_28_10_imag;
  assign io_coef_out_payload_0_28_11_real = int_reg_array_28_11_real;
  assign io_coef_out_payload_0_28_11_imag = int_reg_array_28_11_imag;
  assign io_coef_out_payload_0_28_12_real = int_reg_array_28_12_real;
  assign io_coef_out_payload_0_28_12_imag = int_reg_array_28_12_imag;
  assign io_coef_out_payload_0_28_13_real = int_reg_array_28_13_real;
  assign io_coef_out_payload_0_28_13_imag = int_reg_array_28_13_imag;
  assign io_coef_out_payload_0_28_14_real = int_reg_array_28_14_real;
  assign io_coef_out_payload_0_28_14_imag = int_reg_array_28_14_imag;
  assign io_coef_out_payload_0_28_15_real = int_reg_array_28_15_real;
  assign io_coef_out_payload_0_28_15_imag = int_reg_array_28_15_imag;
  assign io_coef_out_payload_0_28_16_real = int_reg_array_28_16_real;
  assign io_coef_out_payload_0_28_16_imag = int_reg_array_28_16_imag;
  assign io_coef_out_payload_0_28_17_real = int_reg_array_28_17_real;
  assign io_coef_out_payload_0_28_17_imag = int_reg_array_28_17_imag;
  assign io_coef_out_payload_0_28_18_real = int_reg_array_28_18_real;
  assign io_coef_out_payload_0_28_18_imag = int_reg_array_28_18_imag;
  assign io_coef_out_payload_0_28_19_real = int_reg_array_28_19_real;
  assign io_coef_out_payload_0_28_19_imag = int_reg_array_28_19_imag;
  assign io_coef_out_payload_0_28_20_real = int_reg_array_28_20_real;
  assign io_coef_out_payload_0_28_20_imag = int_reg_array_28_20_imag;
  assign io_coef_out_payload_0_28_21_real = int_reg_array_28_21_real;
  assign io_coef_out_payload_0_28_21_imag = int_reg_array_28_21_imag;
  assign io_coef_out_payload_0_28_22_real = int_reg_array_28_22_real;
  assign io_coef_out_payload_0_28_22_imag = int_reg_array_28_22_imag;
  assign io_coef_out_payload_0_28_23_real = int_reg_array_28_23_real;
  assign io_coef_out_payload_0_28_23_imag = int_reg_array_28_23_imag;
  assign io_coef_out_payload_0_28_24_real = int_reg_array_28_24_real;
  assign io_coef_out_payload_0_28_24_imag = int_reg_array_28_24_imag;
  assign io_coef_out_payload_0_28_25_real = int_reg_array_28_25_real;
  assign io_coef_out_payload_0_28_25_imag = int_reg_array_28_25_imag;
  assign io_coef_out_payload_0_28_26_real = int_reg_array_28_26_real;
  assign io_coef_out_payload_0_28_26_imag = int_reg_array_28_26_imag;
  assign io_coef_out_payload_0_28_27_real = int_reg_array_28_27_real;
  assign io_coef_out_payload_0_28_27_imag = int_reg_array_28_27_imag;
  assign io_coef_out_payload_0_28_28_real = int_reg_array_28_28_real;
  assign io_coef_out_payload_0_28_28_imag = int_reg_array_28_28_imag;
  assign io_coef_out_payload_0_28_29_real = int_reg_array_28_29_real;
  assign io_coef_out_payload_0_28_29_imag = int_reg_array_28_29_imag;
  assign io_coef_out_payload_0_28_30_real = int_reg_array_28_30_real;
  assign io_coef_out_payload_0_28_30_imag = int_reg_array_28_30_imag;
  assign io_coef_out_payload_0_28_31_real = int_reg_array_28_31_real;
  assign io_coef_out_payload_0_28_31_imag = int_reg_array_28_31_imag;
  assign io_coef_out_payload_0_28_32_real = int_reg_array_28_32_real;
  assign io_coef_out_payload_0_28_32_imag = int_reg_array_28_32_imag;
  assign io_coef_out_payload_0_28_33_real = int_reg_array_28_33_real;
  assign io_coef_out_payload_0_28_33_imag = int_reg_array_28_33_imag;
  assign io_coef_out_payload_0_28_34_real = int_reg_array_28_34_real;
  assign io_coef_out_payload_0_28_34_imag = int_reg_array_28_34_imag;
  assign io_coef_out_payload_0_28_35_real = int_reg_array_28_35_real;
  assign io_coef_out_payload_0_28_35_imag = int_reg_array_28_35_imag;
  assign io_coef_out_payload_0_28_36_real = int_reg_array_28_36_real;
  assign io_coef_out_payload_0_28_36_imag = int_reg_array_28_36_imag;
  assign io_coef_out_payload_0_28_37_real = int_reg_array_28_37_real;
  assign io_coef_out_payload_0_28_37_imag = int_reg_array_28_37_imag;
  assign io_coef_out_payload_0_28_38_real = int_reg_array_28_38_real;
  assign io_coef_out_payload_0_28_38_imag = int_reg_array_28_38_imag;
  assign io_coef_out_payload_0_28_39_real = int_reg_array_28_39_real;
  assign io_coef_out_payload_0_28_39_imag = int_reg_array_28_39_imag;
  assign io_coef_out_payload_0_28_40_real = int_reg_array_28_40_real;
  assign io_coef_out_payload_0_28_40_imag = int_reg_array_28_40_imag;
  assign io_coef_out_payload_0_28_41_real = int_reg_array_28_41_real;
  assign io_coef_out_payload_0_28_41_imag = int_reg_array_28_41_imag;
  assign io_coef_out_payload_0_28_42_real = int_reg_array_28_42_real;
  assign io_coef_out_payload_0_28_42_imag = int_reg_array_28_42_imag;
  assign io_coef_out_payload_0_28_43_real = int_reg_array_28_43_real;
  assign io_coef_out_payload_0_28_43_imag = int_reg_array_28_43_imag;
  assign io_coef_out_payload_0_28_44_real = int_reg_array_28_44_real;
  assign io_coef_out_payload_0_28_44_imag = int_reg_array_28_44_imag;
  assign io_coef_out_payload_0_28_45_real = int_reg_array_28_45_real;
  assign io_coef_out_payload_0_28_45_imag = int_reg_array_28_45_imag;
  assign io_coef_out_payload_0_28_46_real = int_reg_array_28_46_real;
  assign io_coef_out_payload_0_28_46_imag = int_reg_array_28_46_imag;
  assign io_coef_out_payload_0_28_47_real = int_reg_array_28_47_real;
  assign io_coef_out_payload_0_28_47_imag = int_reg_array_28_47_imag;
  assign io_coef_out_payload_0_28_48_real = int_reg_array_28_48_real;
  assign io_coef_out_payload_0_28_48_imag = int_reg_array_28_48_imag;
  assign io_coef_out_payload_0_28_49_real = int_reg_array_28_49_real;
  assign io_coef_out_payload_0_28_49_imag = int_reg_array_28_49_imag;
  assign io_coef_out_payload_0_29_0_real = int_reg_array_29_0_real;
  assign io_coef_out_payload_0_29_0_imag = int_reg_array_29_0_imag;
  assign io_coef_out_payload_0_29_1_real = int_reg_array_29_1_real;
  assign io_coef_out_payload_0_29_1_imag = int_reg_array_29_1_imag;
  assign io_coef_out_payload_0_29_2_real = int_reg_array_29_2_real;
  assign io_coef_out_payload_0_29_2_imag = int_reg_array_29_2_imag;
  assign io_coef_out_payload_0_29_3_real = int_reg_array_29_3_real;
  assign io_coef_out_payload_0_29_3_imag = int_reg_array_29_3_imag;
  assign io_coef_out_payload_0_29_4_real = int_reg_array_29_4_real;
  assign io_coef_out_payload_0_29_4_imag = int_reg_array_29_4_imag;
  assign io_coef_out_payload_0_29_5_real = int_reg_array_29_5_real;
  assign io_coef_out_payload_0_29_5_imag = int_reg_array_29_5_imag;
  assign io_coef_out_payload_0_29_6_real = int_reg_array_29_6_real;
  assign io_coef_out_payload_0_29_6_imag = int_reg_array_29_6_imag;
  assign io_coef_out_payload_0_29_7_real = int_reg_array_29_7_real;
  assign io_coef_out_payload_0_29_7_imag = int_reg_array_29_7_imag;
  assign io_coef_out_payload_0_29_8_real = int_reg_array_29_8_real;
  assign io_coef_out_payload_0_29_8_imag = int_reg_array_29_8_imag;
  assign io_coef_out_payload_0_29_9_real = int_reg_array_29_9_real;
  assign io_coef_out_payload_0_29_9_imag = int_reg_array_29_9_imag;
  assign io_coef_out_payload_0_29_10_real = int_reg_array_29_10_real;
  assign io_coef_out_payload_0_29_10_imag = int_reg_array_29_10_imag;
  assign io_coef_out_payload_0_29_11_real = int_reg_array_29_11_real;
  assign io_coef_out_payload_0_29_11_imag = int_reg_array_29_11_imag;
  assign io_coef_out_payload_0_29_12_real = int_reg_array_29_12_real;
  assign io_coef_out_payload_0_29_12_imag = int_reg_array_29_12_imag;
  assign io_coef_out_payload_0_29_13_real = int_reg_array_29_13_real;
  assign io_coef_out_payload_0_29_13_imag = int_reg_array_29_13_imag;
  assign io_coef_out_payload_0_29_14_real = int_reg_array_29_14_real;
  assign io_coef_out_payload_0_29_14_imag = int_reg_array_29_14_imag;
  assign io_coef_out_payload_0_29_15_real = int_reg_array_29_15_real;
  assign io_coef_out_payload_0_29_15_imag = int_reg_array_29_15_imag;
  assign io_coef_out_payload_0_29_16_real = int_reg_array_29_16_real;
  assign io_coef_out_payload_0_29_16_imag = int_reg_array_29_16_imag;
  assign io_coef_out_payload_0_29_17_real = int_reg_array_29_17_real;
  assign io_coef_out_payload_0_29_17_imag = int_reg_array_29_17_imag;
  assign io_coef_out_payload_0_29_18_real = int_reg_array_29_18_real;
  assign io_coef_out_payload_0_29_18_imag = int_reg_array_29_18_imag;
  assign io_coef_out_payload_0_29_19_real = int_reg_array_29_19_real;
  assign io_coef_out_payload_0_29_19_imag = int_reg_array_29_19_imag;
  assign io_coef_out_payload_0_29_20_real = int_reg_array_29_20_real;
  assign io_coef_out_payload_0_29_20_imag = int_reg_array_29_20_imag;
  assign io_coef_out_payload_0_29_21_real = int_reg_array_29_21_real;
  assign io_coef_out_payload_0_29_21_imag = int_reg_array_29_21_imag;
  assign io_coef_out_payload_0_29_22_real = int_reg_array_29_22_real;
  assign io_coef_out_payload_0_29_22_imag = int_reg_array_29_22_imag;
  assign io_coef_out_payload_0_29_23_real = int_reg_array_29_23_real;
  assign io_coef_out_payload_0_29_23_imag = int_reg_array_29_23_imag;
  assign io_coef_out_payload_0_29_24_real = int_reg_array_29_24_real;
  assign io_coef_out_payload_0_29_24_imag = int_reg_array_29_24_imag;
  assign io_coef_out_payload_0_29_25_real = int_reg_array_29_25_real;
  assign io_coef_out_payload_0_29_25_imag = int_reg_array_29_25_imag;
  assign io_coef_out_payload_0_29_26_real = int_reg_array_29_26_real;
  assign io_coef_out_payload_0_29_26_imag = int_reg_array_29_26_imag;
  assign io_coef_out_payload_0_29_27_real = int_reg_array_29_27_real;
  assign io_coef_out_payload_0_29_27_imag = int_reg_array_29_27_imag;
  assign io_coef_out_payload_0_29_28_real = int_reg_array_29_28_real;
  assign io_coef_out_payload_0_29_28_imag = int_reg_array_29_28_imag;
  assign io_coef_out_payload_0_29_29_real = int_reg_array_29_29_real;
  assign io_coef_out_payload_0_29_29_imag = int_reg_array_29_29_imag;
  assign io_coef_out_payload_0_29_30_real = int_reg_array_29_30_real;
  assign io_coef_out_payload_0_29_30_imag = int_reg_array_29_30_imag;
  assign io_coef_out_payload_0_29_31_real = int_reg_array_29_31_real;
  assign io_coef_out_payload_0_29_31_imag = int_reg_array_29_31_imag;
  assign io_coef_out_payload_0_29_32_real = int_reg_array_29_32_real;
  assign io_coef_out_payload_0_29_32_imag = int_reg_array_29_32_imag;
  assign io_coef_out_payload_0_29_33_real = int_reg_array_29_33_real;
  assign io_coef_out_payload_0_29_33_imag = int_reg_array_29_33_imag;
  assign io_coef_out_payload_0_29_34_real = int_reg_array_29_34_real;
  assign io_coef_out_payload_0_29_34_imag = int_reg_array_29_34_imag;
  assign io_coef_out_payload_0_29_35_real = int_reg_array_29_35_real;
  assign io_coef_out_payload_0_29_35_imag = int_reg_array_29_35_imag;
  assign io_coef_out_payload_0_29_36_real = int_reg_array_29_36_real;
  assign io_coef_out_payload_0_29_36_imag = int_reg_array_29_36_imag;
  assign io_coef_out_payload_0_29_37_real = int_reg_array_29_37_real;
  assign io_coef_out_payload_0_29_37_imag = int_reg_array_29_37_imag;
  assign io_coef_out_payload_0_29_38_real = int_reg_array_29_38_real;
  assign io_coef_out_payload_0_29_38_imag = int_reg_array_29_38_imag;
  assign io_coef_out_payload_0_29_39_real = int_reg_array_29_39_real;
  assign io_coef_out_payload_0_29_39_imag = int_reg_array_29_39_imag;
  assign io_coef_out_payload_0_29_40_real = int_reg_array_29_40_real;
  assign io_coef_out_payload_0_29_40_imag = int_reg_array_29_40_imag;
  assign io_coef_out_payload_0_29_41_real = int_reg_array_29_41_real;
  assign io_coef_out_payload_0_29_41_imag = int_reg_array_29_41_imag;
  assign io_coef_out_payload_0_29_42_real = int_reg_array_29_42_real;
  assign io_coef_out_payload_0_29_42_imag = int_reg_array_29_42_imag;
  assign io_coef_out_payload_0_29_43_real = int_reg_array_29_43_real;
  assign io_coef_out_payload_0_29_43_imag = int_reg_array_29_43_imag;
  assign io_coef_out_payload_0_29_44_real = int_reg_array_29_44_real;
  assign io_coef_out_payload_0_29_44_imag = int_reg_array_29_44_imag;
  assign io_coef_out_payload_0_29_45_real = int_reg_array_29_45_real;
  assign io_coef_out_payload_0_29_45_imag = int_reg_array_29_45_imag;
  assign io_coef_out_payload_0_29_46_real = int_reg_array_29_46_real;
  assign io_coef_out_payload_0_29_46_imag = int_reg_array_29_46_imag;
  assign io_coef_out_payload_0_29_47_real = int_reg_array_29_47_real;
  assign io_coef_out_payload_0_29_47_imag = int_reg_array_29_47_imag;
  assign io_coef_out_payload_0_29_48_real = int_reg_array_29_48_real;
  assign io_coef_out_payload_0_29_48_imag = int_reg_array_29_48_imag;
  assign io_coef_out_payload_0_29_49_real = int_reg_array_29_49_real;
  assign io_coef_out_payload_0_29_49_imag = int_reg_array_29_49_imag;
  assign io_coef_out_payload_0_30_0_real = int_reg_array_30_0_real;
  assign io_coef_out_payload_0_30_0_imag = int_reg_array_30_0_imag;
  assign io_coef_out_payload_0_30_1_real = int_reg_array_30_1_real;
  assign io_coef_out_payload_0_30_1_imag = int_reg_array_30_1_imag;
  assign io_coef_out_payload_0_30_2_real = int_reg_array_30_2_real;
  assign io_coef_out_payload_0_30_2_imag = int_reg_array_30_2_imag;
  assign io_coef_out_payload_0_30_3_real = int_reg_array_30_3_real;
  assign io_coef_out_payload_0_30_3_imag = int_reg_array_30_3_imag;
  assign io_coef_out_payload_0_30_4_real = int_reg_array_30_4_real;
  assign io_coef_out_payload_0_30_4_imag = int_reg_array_30_4_imag;
  assign io_coef_out_payload_0_30_5_real = int_reg_array_30_5_real;
  assign io_coef_out_payload_0_30_5_imag = int_reg_array_30_5_imag;
  assign io_coef_out_payload_0_30_6_real = int_reg_array_30_6_real;
  assign io_coef_out_payload_0_30_6_imag = int_reg_array_30_6_imag;
  assign io_coef_out_payload_0_30_7_real = int_reg_array_30_7_real;
  assign io_coef_out_payload_0_30_7_imag = int_reg_array_30_7_imag;
  assign io_coef_out_payload_0_30_8_real = int_reg_array_30_8_real;
  assign io_coef_out_payload_0_30_8_imag = int_reg_array_30_8_imag;
  assign io_coef_out_payload_0_30_9_real = int_reg_array_30_9_real;
  assign io_coef_out_payload_0_30_9_imag = int_reg_array_30_9_imag;
  assign io_coef_out_payload_0_30_10_real = int_reg_array_30_10_real;
  assign io_coef_out_payload_0_30_10_imag = int_reg_array_30_10_imag;
  assign io_coef_out_payload_0_30_11_real = int_reg_array_30_11_real;
  assign io_coef_out_payload_0_30_11_imag = int_reg_array_30_11_imag;
  assign io_coef_out_payload_0_30_12_real = int_reg_array_30_12_real;
  assign io_coef_out_payload_0_30_12_imag = int_reg_array_30_12_imag;
  assign io_coef_out_payload_0_30_13_real = int_reg_array_30_13_real;
  assign io_coef_out_payload_0_30_13_imag = int_reg_array_30_13_imag;
  assign io_coef_out_payload_0_30_14_real = int_reg_array_30_14_real;
  assign io_coef_out_payload_0_30_14_imag = int_reg_array_30_14_imag;
  assign io_coef_out_payload_0_30_15_real = int_reg_array_30_15_real;
  assign io_coef_out_payload_0_30_15_imag = int_reg_array_30_15_imag;
  assign io_coef_out_payload_0_30_16_real = int_reg_array_30_16_real;
  assign io_coef_out_payload_0_30_16_imag = int_reg_array_30_16_imag;
  assign io_coef_out_payload_0_30_17_real = int_reg_array_30_17_real;
  assign io_coef_out_payload_0_30_17_imag = int_reg_array_30_17_imag;
  assign io_coef_out_payload_0_30_18_real = int_reg_array_30_18_real;
  assign io_coef_out_payload_0_30_18_imag = int_reg_array_30_18_imag;
  assign io_coef_out_payload_0_30_19_real = int_reg_array_30_19_real;
  assign io_coef_out_payload_0_30_19_imag = int_reg_array_30_19_imag;
  assign io_coef_out_payload_0_30_20_real = int_reg_array_30_20_real;
  assign io_coef_out_payload_0_30_20_imag = int_reg_array_30_20_imag;
  assign io_coef_out_payload_0_30_21_real = int_reg_array_30_21_real;
  assign io_coef_out_payload_0_30_21_imag = int_reg_array_30_21_imag;
  assign io_coef_out_payload_0_30_22_real = int_reg_array_30_22_real;
  assign io_coef_out_payload_0_30_22_imag = int_reg_array_30_22_imag;
  assign io_coef_out_payload_0_30_23_real = int_reg_array_30_23_real;
  assign io_coef_out_payload_0_30_23_imag = int_reg_array_30_23_imag;
  assign io_coef_out_payload_0_30_24_real = int_reg_array_30_24_real;
  assign io_coef_out_payload_0_30_24_imag = int_reg_array_30_24_imag;
  assign io_coef_out_payload_0_30_25_real = int_reg_array_30_25_real;
  assign io_coef_out_payload_0_30_25_imag = int_reg_array_30_25_imag;
  assign io_coef_out_payload_0_30_26_real = int_reg_array_30_26_real;
  assign io_coef_out_payload_0_30_26_imag = int_reg_array_30_26_imag;
  assign io_coef_out_payload_0_30_27_real = int_reg_array_30_27_real;
  assign io_coef_out_payload_0_30_27_imag = int_reg_array_30_27_imag;
  assign io_coef_out_payload_0_30_28_real = int_reg_array_30_28_real;
  assign io_coef_out_payload_0_30_28_imag = int_reg_array_30_28_imag;
  assign io_coef_out_payload_0_30_29_real = int_reg_array_30_29_real;
  assign io_coef_out_payload_0_30_29_imag = int_reg_array_30_29_imag;
  assign io_coef_out_payload_0_30_30_real = int_reg_array_30_30_real;
  assign io_coef_out_payload_0_30_30_imag = int_reg_array_30_30_imag;
  assign io_coef_out_payload_0_30_31_real = int_reg_array_30_31_real;
  assign io_coef_out_payload_0_30_31_imag = int_reg_array_30_31_imag;
  assign io_coef_out_payload_0_30_32_real = int_reg_array_30_32_real;
  assign io_coef_out_payload_0_30_32_imag = int_reg_array_30_32_imag;
  assign io_coef_out_payload_0_30_33_real = int_reg_array_30_33_real;
  assign io_coef_out_payload_0_30_33_imag = int_reg_array_30_33_imag;
  assign io_coef_out_payload_0_30_34_real = int_reg_array_30_34_real;
  assign io_coef_out_payload_0_30_34_imag = int_reg_array_30_34_imag;
  assign io_coef_out_payload_0_30_35_real = int_reg_array_30_35_real;
  assign io_coef_out_payload_0_30_35_imag = int_reg_array_30_35_imag;
  assign io_coef_out_payload_0_30_36_real = int_reg_array_30_36_real;
  assign io_coef_out_payload_0_30_36_imag = int_reg_array_30_36_imag;
  assign io_coef_out_payload_0_30_37_real = int_reg_array_30_37_real;
  assign io_coef_out_payload_0_30_37_imag = int_reg_array_30_37_imag;
  assign io_coef_out_payload_0_30_38_real = int_reg_array_30_38_real;
  assign io_coef_out_payload_0_30_38_imag = int_reg_array_30_38_imag;
  assign io_coef_out_payload_0_30_39_real = int_reg_array_30_39_real;
  assign io_coef_out_payload_0_30_39_imag = int_reg_array_30_39_imag;
  assign io_coef_out_payload_0_30_40_real = int_reg_array_30_40_real;
  assign io_coef_out_payload_0_30_40_imag = int_reg_array_30_40_imag;
  assign io_coef_out_payload_0_30_41_real = int_reg_array_30_41_real;
  assign io_coef_out_payload_0_30_41_imag = int_reg_array_30_41_imag;
  assign io_coef_out_payload_0_30_42_real = int_reg_array_30_42_real;
  assign io_coef_out_payload_0_30_42_imag = int_reg_array_30_42_imag;
  assign io_coef_out_payload_0_30_43_real = int_reg_array_30_43_real;
  assign io_coef_out_payload_0_30_43_imag = int_reg_array_30_43_imag;
  assign io_coef_out_payload_0_30_44_real = int_reg_array_30_44_real;
  assign io_coef_out_payload_0_30_44_imag = int_reg_array_30_44_imag;
  assign io_coef_out_payload_0_30_45_real = int_reg_array_30_45_real;
  assign io_coef_out_payload_0_30_45_imag = int_reg_array_30_45_imag;
  assign io_coef_out_payload_0_30_46_real = int_reg_array_30_46_real;
  assign io_coef_out_payload_0_30_46_imag = int_reg_array_30_46_imag;
  assign io_coef_out_payload_0_30_47_real = int_reg_array_30_47_real;
  assign io_coef_out_payload_0_30_47_imag = int_reg_array_30_47_imag;
  assign io_coef_out_payload_0_30_48_real = int_reg_array_30_48_real;
  assign io_coef_out_payload_0_30_48_imag = int_reg_array_30_48_imag;
  assign io_coef_out_payload_0_30_49_real = int_reg_array_30_49_real;
  assign io_coef_out_payload_0_30_49_imag = int_reg_array_30_49_imag;
  assign io_coef_out_payload_0_31_0_real = int_reg_array_31_0_real;
  assign io_coef_out_payload_0_31_0_imag = int_reg_array_31_0_imag;
  assign io_coef_out_payload_0_31_1_real = int_reg_array_31_1_real;
  assign io_coef_out_payload_0_31_1_imag = int_reg_array_31_1_imag;
  assign io_coef_out_payload_0_31_2_real = int_reg_array_31_2_real;
  assign io_coef_out_payload_0_31_2_imag = int_reg_array_31_2_imag;
  assign io_coef_out_payload_0_31_3_real = int_reg_array_31_3_real;
  assign io_coef_out_payload_0_31_3_imag = int_reg_array_31_3_imag;
  assign io_coef_out_payload_0_31_4_real = int_reg_array_31_4_real;
  assign io_coef_out_payload_0_31_4_imag = int_reg_array_31_4_imag;
  assign io_coef_out_payload_0_31_5_real = int_reg_array_31_5_real;
  assign io_coef_out_payload_0_31_5_imag = int_reg_array_31_5_imag;
  assign io_coef_out_payload_0_31_6_real = int_reg_array_31_6_real;
  assign io_coef_out_payload_0_31_6_imag = int_reg_array_31_6_imag;
  assign io_coef_out_payload_0_31_7_real = int_reg_array_31_7_real;
  assign io_coef_out_payload_0_31_7_imag = int_reg_array_31_7_imag;
  assign io_coef_out_payload_0_31_8_real = int_reg_array_31_8_real;
  assign io_coef_out_payload_0_31_8_imag = int_reg_array_31_8_imag;
  assign io_coef_out_payload_0_31_9_real = int_reg_array_31_9_real;
  assign io_coef_out_payload_0_31_9_imag = int_reg_array_31_9_imag;
  assign io_coef_out_payload_0_31_10_real = int_reg_array_31_10_real;
  assign io_coef_out_payload_0_31_10_imag = int_reg_array_31_10_imag;
  assign io_coef_out_payload_0_31_11_real = int_reg_array_31_11_real;
  assign io_coef_out_payload_0_31_11_imag = int_reg_array_31_11_imag;
  assign io_coef_out_payload_0_31_12_real = int_reg_array_31_12_real;
  assign io_coef_out_payload_0_31_12_imag = int_reg_array_31_12_imag;
  assign io_coef_out_payload_0_31_13_real = int_reg_array_31_13_real;
  assign io_coef_out_payload_0_31_13_imag = int_reg_array_31_13_imag;
  assign io_coef_out_payload_0_31_14_real = int_reg_array_31_14_real;
  assign io_coef_out_payload_0_31_14_imag = int_reg_array_31_14_imag;
  assign io_coef_out_payload_0_31_15_real = int_reg_array_31_15_real;
  assign io_coef_out_payload_0_31_15_imag = int_reg_array_31_15_imag;
  assign io_coef_out_payload_0_31_16_real = int_reg_array_31_16_real;
  assign io_coef_out_payload_0_31_16_imag = int_reg_array_31_16_imag;
  assign io_coef_out_payload_0_31_17_real = int_reg_array_31_17_real;
  assign io_coef_out_payload_0_31_17_imag = int_reg_array_31_17_imag;
  assign io_coef_out_payload_0_31_18_real = int_reg_array_31_18_real;
  assign io_coef_out_payload_0_31_18_imag = int_reg_array_31_18_imag;
  assign io_coef_out_payload_0_31_19_real = int_reg_array_31_19_real;
  assign io_coef_out_payload_0_31_19_imag = int_reg_array_31_19_imag;
  assign io_coef_out_payload_0_31_20_real = int_reg_array_31_20_real;
  assign io_coef_out_payload_0_31_20_imag = int_reg_array_31_20_imag;
  assign io_coef_out_payload_0_31_21_real = int_reg_array_31_21_real;
  assign io_coef_out_payload_0_31_21_imag = int_reg_array_31_21_imag;
  assign io_coef_out_payload_0_31_22_real = int_reg_array_31_22_real;
  assign io_coef_out_payload_0_31_22_imag = int_reg_array_31_22_imag;
  assign io_coef_out_payload_0_31_23_real = int_reg_array_31_23_real;
  assign io_coef_out_payload_0_31_23_imag = int_reg_array_31_23_imag;
  assign io_coef_out_payload_0_31_24_real = int_reg_array_31_24_real;
  assign io_coef_out_payload_0_31_24_imag = int_reg_array_31_24_imag;
  assign io_coef_out_payload_0_31_25_real = int_reg_array_31_25_real;
  assign io_coef_out_payload_0_31_25_imag = int_reg_array_31_25_imag;
  assign io_coef_out_payload_0_31_26_real = int_reg_array_31_26_real;
  assign io_coef_out_payload_0_31_26_imag = int_reg_array_31_26_imag;
  assign io_coef_out_payload_0_31_27_real = int_reg_array_31_27_real;
  assign io_coef_out_payload_0_31_27_imag = int_reg_array_31_27_imag;
  assign io_coef_out_payload_0_31_28_real = int_reg_array_31_28_real;
  assign io_coef_out_payload_0_31_28_imag = int_reg_array_31_28_imag;
  assign io_coef_out_payload_0_31_29_real = int_reg_array_31_29_real;
  assign io_coef_out_payload_0_31_29_imag = int_reg_array_31_29_imag;
  assign io_coef_out_payload_0_31_30_real = int_reg_array_31_30_real;
  assign io_coef_out_payload_0_31_30_imag = int_reg_array_31_30_imag;
  assign io_coef_out_payload_0_31_31_real = int_reg_array_31_31_real;
  assign io_coef_out_payload_0_31_31_imag = int_reg_array_31_31_imag;
  assign io_coef_out_payload_0_31_32_real = int_reg_array_31_32_real;
  assign io_coef_out_payload_0_31_32_imag = int_reg_array_31_32_imag;
  assign io_coef_out_payload_0_31_33_real = int_reg_array_31_33_real;
  assign io_coef_out_payload_0_31_33_imag = int_reg_array_31_33_imag;
  assign io_coef_out_payload_0_31_34_real = int_reg_array_31_34_real;
  assign io_coef_out_payload_0_31_34_imag = int_reg_array_31_34_imag;
  assign io_coef_out_payload_0_31_35_real = int_reg_array_31_35_real;
  assign io_coef_out_payload_0_31_35_imag = int_reg_array_31_35_imag;
  assign io_coef_out_payload_0_31_36_real = int_reg_array_31_36_real;
  assign io_coef_out_payload_0_31_36_imag = int_reg_array_31_36_imag;
  assign io_coef_out_payload_0_31_37_real = int_reg_array_31_37_real;
  assign io_coef_out_payload_0_31_37_imag = int_reg_array_31_37_imag;
  assign io_coef_out_payload_0_31_38_real = int_reg_array_31_38_real;
  assign io_coef_out_payload_0_31_38_imag = int_reg_array_31_38_imag;
  assign io_coef_out_payload_0_31_39_real = int_reg_array_31_39_real;
  assign io_coef_out_payload_0_31_39_imag = int_reg_array_31_39_imag;
  assign io_coef_out_payload_0_31_40_real = int_reg_array_31_40_real;
  assign io_coef_out_payload_0_31_40_imag = int_reg_array_31_40_imag;
  assign io_coef_out_payload_0_31_41_real = int_reg_array_31_41_real;
  assign io_coef_out_payload_0_31_41_imag = int_reg_array_31_41_imag;
  assign io_coef_out_payload_0_31_42_real = int_reg_array_31_42_real;
  assign io_coef_out_payload_0_31_42_imag = int_reg_array_31_42_imag;
  assign io_coef_out_payload_0_31_43_real = int_reg_array_31_43_real;
  assign io_coef_out_payload_0_31_43_imag = int_reg_array_31_43_imag;
  assign io_coef_out_payload_0_31_44_real = int_reg_array_31_44_real;
  assign io_coef_out_payload_0_31_44_imag = int_reg_array_31_44_imag;
  assign io_coef_out_payload_0_31_45_real = int_reg_array_31_45_real;
  assign io_coef_out_payload_0_31_45_imag = int_reg_array_31_45_imag;
  assign io_coef_out_payload_0_31_46_real = int_reg_array_31_46_real;
  assign io_coef_out_payload_0_31_46_imag = int_reg_array_31_46_imag;
  assign io_coef_out_payload_0_31_47_real = int_reg_array_31_47_real;
  assign io_coef_out_payload_0_31_47_imag = int_reg_array_31_47_imag;
  assign io_coef_out_payload_0_31_48_real = int_reg_array_31_48_real;
  assign io_coef_out_payload_0_31_48_imag = int_reg_array_31_48_imag;
  assign io_coef_out_payload_0_31_49_real = int_reg_array_31_49_real;
  assign io_coef_out_payload_0_31_49_imag = int_reg_array_31_49_imag;
  assign io_coef_out_payload_0_32_0_real = int_reg_array_32_0_real;
  assign io_coef_out_payload_0_32_0_imag = int_reg_array_32_0_imag;
  assign io_coef_out_payload_0_32_1_real = int_reg_array_32_1_real;
  assign io_coef_out_payload_0_32_1_imag = int_reg_array_32_1_imag;
  assign io_coef_out_payload_0_32_2_real = int_reg_array_32_2_real;
  assign io_coef_out_payload_0_32_2_imag = int_reg_array_32_2_imag;
  assign io_coef_out_payload_0_32_3_real = int_reg_array_32_3_real;
  assign io_coef_out_payload_0_32_3_imag = int_reg_array_32_3_imag;
  assign io_coef_out_payload_0_32_4_real = int_reg_array_32_4_real;
  assign io_coef_out_payload_0_32_4_imag = int_reg_array_32_4_imag;
  assign io_coef_out_payload_0_32_5_real = int_reg_array_32_5_real;
  assign io_coef_out_payload_0_32_5_imag = int_reg_array_32_5_imag;
  assign io_coef_out_payload_0_32_6_real = int_reg_array_32_6_real;
  assign io_coef_out_payload_0_32_6_imag = int_reg_array_32_6_imag;
  assign io_coef_out_payload_0_32_7_real = int_reg_array_32_7_real;
  assign io_coef_out_payload_0_32_7_imag = int_reg_array_32_7_imag;
  assign io_coef_out_payload_0_32_8_real = int_reg_array_32_8_real;
  assign io_coef_out_payload_0_32_8_imag = int_reg_array_32_8_imag;
  assign io_coef_out_payload_0_32_9_real = int_reg_array_32_9_real;
  assign io_coef_out_payload_0_32_9_imag = int_reg_array_32_9_imag;
  assign io_coef_out_payload_0_32_10_real = int_reg_array_32_10_real;
  assign io_coef_out_payload_0_32_10_imag = int_reg_array_32_10_imag;
  assign io_coef_out_payload_0_32_11_real = int_reg_array_32_11_real;
  assign io_coef_out_payload_0_32_11_imag = int_reg_array_32_11_imag;
  assign io_coef_out_payload_0_32_12_real = int_reg_array_32_12_real;
  assign io_coef_out_payload_0_32_12_imag = int_reg_array_32_12_imag;
  assign io_coef_out_payload_0_32_13_real = int_reg_array_32_13_real;
  assign io_coef_out_payload_0_32_13_imag = int_reg_array_32_13_imag;
  assign io_coef_out_payload_0_32_14_real = int_reg_array_32_14_real;
  assign io_coef_out_payload_0_32_14_imag = int_reg_array_32_14_imag;
  assign io_coef_out_payload_0_32_15_real = int_reg_array_32_15_real;
  assign io_coef_out_payload_0_32_15_imag = int_reg_array_32_15_imag;
  assign io_coef_out_payload_0_32_16_real = int_reg_array_32_16_real;
  assign io_coef_out_payload_0_32_16_imag = int_reg_array_32_16_imag;
  assign io_coef_out_payload_0_32_17_real = int_reg_array_32_17_real;
  assign io_coef_out_payload_0_32_17_imag = int_reg_array_32_17_imag;
  assign io_coef_out_payload_0_32_18_real = int_reg_array_32_18_real;
  assign io_coef_out_payload_0_32_18_imag = int_reg_array_32_18_imag;
  assign io_coef_out_payload_0_32_19_real = int_reg_array_32_19_real;
  assign io_coef_out_payload_0_32_19_imag = int_reg_array_32_19_imag;
  assign io_coef_out_payload_0_32_20_real = int_reg_array_32_20_real;
  assign io_coef_out_payload_0_32_20_imag = int_reg_array_32_20_imag;
  assign io_coef_out_payload_0_32_21_real = int_reg_array_32_21_real;
  assign io_coef_out_payload_0_32_21_imag = int_reg_array_32_21_imag;
  assign io_coef_out_payload_0_32_22_real = int_reg_array_32_22_real;
  assign io_coef_out_payload_0_32_22_imag = int_reg_array_32_22_imag;
  assign io_coef_out_payload_0_32_23_real = int_reg_array_32_23_real;
  assign io_coef_out_payload_0_32_23_imag = int_reg_array_32_23_imag;
  assign io_coef_out_payload_0_32_24_real = int_reg_array_32_24_real;
  assign io_coef_out_payload_0_32_24_imag = int_reg_array_32_24_imag;
  assign io_coef_out_payload_0_32_25_real = int_reg_array_32_25_real;
  assign io_coef_out_payload_0_32_25_imag = int_reg_array_32_25_imag;
  assign io_coef_out_payload_0_32_26_real = int_reg_array_32_26_real;
  assign io_coef_out_payload_0_32_26_imag = int_reg_array_32_26_imag;
  assign io_coef_out_payload_0_32_27_real = int_reg_array_32_27_real;
  assign io_coef_out_payload_0_32_27_imag = int_reg_array_32_27_imag;
  assign io_coef_out_payload_0_32_28_real = int_reg_array_32_28_real;
  assign io_coef_out_payload_0_32_28_imag = int_reg_array_32_28_imag;
  assign io_coef_out_payload_0_32_29_real = int_reg_array_32_29_real;
  assign io_coef_out_payload_0_32_29_imag = int_reg_array_32_29_imag;
  assign io_coef_out_payload_0_32_30_real = int_reg_array_32_30_real;
  assign io_coef_out_payload_0_32_30_imag = int_reg_array_32_30_imag;
  assign io_coef_out_payload_0_32_31_real = int_reg_array_32_31_real;
  assign io_coef_out_payload_0_32_31_imag = int_reg_array_32_31_imag;
  assign io_coef_out_payload_0_32_32_real = int_reg_array_32_32_real;
  assign io_coef_out_payload_0_32_32_imag = int_reg_array_32_32_imag;
  assign io_coef_out_payload_0_32_33_real = int_reg_array_32_33_real;
  assign io_coef_out_payload_0_32_33_imag = int_reg_array_32_33_imag;
  assign io_coef_out_payload_0_32_34_real = int_reg_array_32_34_real;
  assign io_coef_out_payload_0_32_34_imag = int_reg_array_32_34_imag;
  assign io_coef_out_payload_0_32_35_real = int_reg_array_32_35_real;
  assign io_coef_out_payload_0_32_35_imag = int_reg_array_32_35_imag;
  assign io_coef_out_payload_0_32_36_real = int_reg_array_32_36_real;
  assign io_coef_out_payload_0_32_36_imag = int_reg_array_32_36_imag;
  assign io_coef_out_payload_0_32_37_real = int_reg_array_32_37_real;
  assign io_coef_out_payload_0_32_37_imag = int_reg_array_32_37_imag;
  assign io_coef_out_payload_0_32_38_real = int_reg_array_32_38_real;
  assign io_coef_out_payload_0_32_38_imag = int_reg_array_32_38_imag;
  assign io_coef_out_payload_0_32_39_real = int_reg_array_32_39_real;
  assign io_coef_out_payload_0_32_39_imag = int_reg_array_32_39_imag;
  assign io_coef_out_payload_0_32_40_real = int_reg_array_32_40_real;
  assign io_coef_out_payload_0_32_40_imag = int_reg_array_32_40_imag;
  assign io_coef_out_payload_0_32_41_real = int_reg_array_32_41_real;
  assign io_coef_out_payload_0_32_41_imag = int_reg_array_32_41_imag;
  assign io_coef_out_payload_0_32_42_real = int_reg_array_32_42_real;
  assign io_coef_out_payload_0_32_42_imag = int_reg_array_32_42_imag;
  assign io_coef_out_payload_0_32_43_real = int_reg_array_32_43_real;
  assign io_coef_out_payload_0_32_43_imag = int_reg_array_32_43_imag;
  assign io_coef_out_payload_0_32_44_real = int_reg_array_32_44_real;
  assign io_coef_out_payload_0_32_44_imag = int_reg_array_32_44_imag;
  assign io_coef_out_payload_0_32_45_real = int_reg_array_32_45_real;
  assign io_coef_out_payload_0_32_45_imag = int_reg_array_32_45_imag;
  assign io_coef_out_payload_0_32_46_real = int_reg_array_32_46_real;
  assign io_coef_out_payload_0_32_46_imag = int_reg_array_32_46_imag;
  assign io_coef_out_payload_0_32_47_real = int_reg_array_32_47_real;
  assign io_coef_out_payload_0_32_47_imag = int_reg_array_32_47_imag;
  assign io_coef_out_payload_0_32_48_real = int_reg_array_32_48_real;
  assign io_coef_out_payload_0_32_48_imag = int_reg_array_32_48_imag;
  assign io_coef_out_payload_0_32_49_real = int_reg_array_32_49_real;
  assign io_coef_out_payload_0_32_49_imag = int_reg_array_32_49_imag;
  assign io_coef_out_payload_0_33_0_real = int_reg_array_33_0_real;
  assign io_coef_out_payload_0_33_0_imag = int_reg_array_33_0_imag;
  assign io_coef_out_payload_0_33_1_real = int_reg_array_33_1_real;
  assign io_coef_out_payload_0_33_1_imag = int_reg_array_33_1_imag;
  assign io_coef_out_payload_0_33_2_real = int_reg_array_33_2_real;
  assign io_coef_out_payload_0_33_2_imag = int_reg_array_33_2_imag;
  assign io_coef_out_payload_0_33_3_real = int_reg_array_33_3_real;
  assign io_coef_out_payload_0_33_3_imag = int_reg_array_33_3_imag;
  assign io_coef_out_payload_0_33_4_real = int_reg_array_33_4_real;
  assign io_coef_out_payload_0_33_4_imag = int_reg_array_33_4_imag;
  assign io_coef_out_payload_0_33_5_real = int_reg_array_33_5_real;
  assign io_coef_out_payload_0_33_5_imag = int_reg_array_33_5_imag;
  assign io_coef_out_payload_0_33_6_real = int_reg_array_33_6_real;
  assign io_coef_out_payload_0_33_6_imag = int_reg_array_33_6_imag;
  assign io_coef_out_payload_0_33_7_real = int_reg_array_33_7_real;
  assign io_coef_out_payload_0_33_7_imag = int_reg_array_33_7_imag;
  assign io_coef_out_payload_0_33_8_real = int_reg_array_33_8_real;
  assign io_coef_out_payload_0_33_8_imag = int_reg_array_33_8_imag;
  assign io_coef_out_payload_0_33_9_real = int_reg_array_33_9_real;
  assign io_coef_out_payload_0_33_9_imag = int_reg_array_33_9_imag;
  assign io_coef_out_payload_0_33_10_real = int_reg_array_33_10_real;
  assign io_coef_out_payload_0_33_10_imag = int_reg_array_33_10_imag;
  assign io_coef_out_payload_0_33_11_real = int_reg_array_33_11_real;
  assign io_coef_out_payload_0_33_11_imag = int_reg_array_33_11_imag;
  assign io_coef_out_payload_0_33_12_real = int_reg_array_33_12_real;
  assign io_coef_out_payload_0_33_12_imag = int_reg_array_33_12_imag;
  assign io_coef_out_payload_0_33_13_real = int_reg_array_33_13_real;
  assign io_coef_out_payload_0_33_13_imag = int_reg_array_33_13_imag;
  assign io_coef_out_payload_0_33_14_real = int_reg_array_33_14_real;
  assign io_coef_out_payload_0_33_14_imag = int_reg_array_33_14_imag;
  assign io_coef_out_payload_0_33_15_real = int_reg_array_33_15_real;
  assign io_coef_out_payload_0_33_15_imag = int_reg_array_33_15_imag;
  assign io_coef_out_payload_0_33_16_real = int_reg_array_33_16_real;
  assign io_coef_out_payload_0_33_16_imag = int_reg_array_33_16_imag;
  assign io_coef_out_payload_0_33_17_real = int_reg_array_33_17_real;
  assign io_coef_out_payload_0_33_17_imag = int_reg_array_33_17_imag;
  assign io_coef_out_payload_0_33_18_real = int_reg_array_33_18_real;
  assign io_coef_out_payload_0_33_18_imag = int_reg_array_33_18_imag;
  assign io_coef_out_payload_0_33_19_real = int_reg_array_33_19_real;
  assign io_coef_out_payload_0_33_19_imag = int_reg_array_33_19_imag;
  assign io_coef_out_payload_0_33_20_real = int_reg_array_33_20_real;
  assign io_coef_out_payload_0_33_20_imag = int_reg_array_33_20_imag;
  assign io_coef_out_payload_0_33_21_real = int_reg_array_33_21_real;
  assign io_coef_out_payload_0_33_21_imag = int_reg_array_33_21_imag;
  assign io_coef_out_payload_0_33_22_real = int_reg_array_33_22_real;
  assign io_coef_out_payload_0_33_22_imag = int_reg_array_33_22_imag;
  assign io_coef_out_payload_0_33_23_real = int_reg_array_33_23_real;
  assign io_coef_out_payload_0_33_23_imag = int_reg_array_33_23_imag;
  assign io_coef_out_payload_0_33_24_real = int_reg_array_33_24_real;
  assign io_coef_out_payload_0_33_24_imag = int_reg_array_33_24_imag;
  assign io_coef_out_payload_0_33_25_real = int_reg_array_33_25_real;
  assign io_coef_out_payload_0_33_25_imag = int_reg_array_33_25_imag;
  assign io_coef_out_payload_0_33_26_real = int_reg_array_33_26_real;
  assign io_coef_out_payload_0_33_26_imag = int_reg_array_33_26_imag;
  assign io_coef_out_payload_0_33_27_real = int_reg_array_33_27_real;
  assign io_coef_out_payload_0_33_27_imag = int_reg_array_33_27_imag;
  assign io_coef_out_payload_0_33_28_real = int_reg_array_33_28_real;
  assign io_coef_out_payload_0_33_28_imag = int_reg_array_33_28_imag;
  assign io_coef_out_payload_0_33_29_real = int_reg_array_33_29_real;
  assign io_coef_out_payload_0_33_29_imag = int_reg_array_33_29_imag;
  assign io_coef_out_payload_0_33_30_real = int_reg_array_33_30_real;
  assign io_coef_out_payload_0_33_30_imag = int_reg_array_33_30_imag;
  assign io_coef_out_payload_0_33_31_real = int_reg_array_33_31_real;
  assign io_coef_out_payload_0_33_31_imag = int_reg_array_33_31_imag;
  assign io_coef_out_payload_0_33_32_real = int_reg_array_33_32_real;
  assign io_coef_out_payload_0_33_32_imag = int_reg_array_33_32_imag;
  assign io_coef_out_payload_0_33_33_real = int_reg_array_33_33_real;
  assign io_coef_out_payload_0_33_33_imag = int_reg_array_33_33_imag;
  assign io_coef_out_payload_0_33_34_real = int_reg_array_33_34_real;
  assign io_coef_out_payload_0_33_34_imag = int_reg_array_33_34_imag;
  assign io_coef_out_payload_0_33_35_real = int_reg_array_33_35_real;
  assign io_coef_out_payload_0_33_35_imag = int_reg_array_33_35_imag;
  assign io_coef_out_payload_0_33_36_real = int_reg_array_33_36_real;
  assign io_coef_out_payload_0_33_36_imag = int_reg_array_33_36_imag;
  assign io_coef_out_payload_0_33_37_real = int_reg_array_33_37_real;
  assign io_coef_out_payload_0_33_37_imag = int_reg_array_33_37_imag;
  assign io_coef_out_payload_0_33_38_real = int_reg_array_33_38_real;
  assign io_coef_out_payload_0_33_38_imag = int_reg_array_33_38_imag;
  assign io_coef_out_payload_0_33_39_real = int_reg_array_33_39_real;
  assign io_coef_out_payload_0_33_39_imag = int_reg_array_33_39_imag;
  assign io_coef_out_payload_0_33_40_real = int_reg_array_33_40_real;
  assign io_coef_out_payload_0_33_40_imag = int_reg_array_33_40_imag;
  assign io_coef_out_payload_0_33_41_real = int_reg_array_33_41_real;
  assign io_coef_out_payload_0_33_41_imag = int_reg_array_33_41_imag;
  assign io_coef_out_payload_0_33_42_real = int_reg_array_33_42_real;
  assign io_coef_out_payload_0_33_42_imag = int_reg_array_33_42_imag;
  assign io_coef_out_payload_0_33_43_real = int_reg_array_33_43_real;
  assign io_coef_out_payload_0_33_43_imag = int_reg_array_33_43_imag;
  assign io_coef_out_payload_0_33_44_real = int_reg_array_33_44_real;
  assign io_coef_out_payload_0_33_44_imag = int_reg_array_33_44_imag;
  assign io_coef_out_payload_0_33_45_real = int_reg_array_33_45_real;
  assign io_coef_out_payload_0_33_45_imag = int_reg_array_33_45_imag;
  assign io_coef_out_payload_0_33_46_real = int_reg_array_33_46_real;
  assign io_coef_out_payload_0_33_46_imag = int_reg_array_33_46_imag;
  assign io_coef_out_payload_0_33_47_real = int_reg_array_33_47_real;
  assign io_coef_out_payload_0_33_47_imag = int_reg_array_33_47_imag;
  assign io_coef_out_payload_0_33_48_real = int_reg_array_33_48_real;
  assign io_coef_out_payload_0_33_48_imag = int_reg_array_33_48_imag;
  assign io_coef_out_payload_0_33_49_real = int_reg_array_33_49_real;
  assign io_coef_out_payload_0_33_49_imag = int_reg_array_33_49_imag;
  assign io_coef_out_payload_0_34_0_real = int_reg_array_34_0_real;
  assign io_coef_out_payload_0_34_0_imag = int_reg_array_34_0_imag;
  assign io_coef_out_payload_0_34_1_real = int_reg_array_34_1_real;
  assign io_coef_out_payload_0_34_1_imag = int_reg_array_34_1_imag;
  assign io_coef_out_payload_0_34_2_real = int_reg_array_34_2_real;
  assign io_coef_out_payload_0_34_2_imag = int_reg_array_34_2_imag;
  assign io_coef_out_payload_0_34_3_real = int_reg_array_34_3_real;
  assign io_coef_out_payload_0_34_3_imag = int_reg_array_34_3_imag;
  assign io_coef_out_payload_0_34_4_real = int_reg_array_34_4_real;
  assign io_coef_out_payload_0_34_4_imag = int_reg_array_34_4_imag;
  assign io_coef_out_payload_0_34_5_real = int_reg_array_34_5_real;
  assign io_coef_out_payload_0_34_5_imag = int_reg_array_34_5_imag;
  assign io_coef_out_payload_0_34_6_real = int_reg_array_34_6_real;
  assign io_coef_out_payload_0_34_6_imag = int_reg_array_34_6_imag;
  assign io_coef_out_payload_0_34_7_real = int_reg_array_34_7_real;
  assign io_coef_out_payload_0_34_7_imag = int_reg_array_34_7_imag;
  assign io_coef_out_payload_0_34_8_real = int_reg_array_34_8_real;
  assign io_coef_out_payload_0_34_8_imag = int_reg_array_34_8_imag;
  assign io_coef_out_payload_0_34_9_real = int_reg_array_34_9_real;
  assign io_coef_out_payload_0_34_9_imag = int_reg_array_34_9_imag;
  assign io_coef_out_payload_0_34_10_real = int_reg_array_34_10_real;
  assign io_coef_out_payload_0_34_10_imag = int_reg_array_34_10_imag;
  assign io_coef_out_payload_0_34_11_real = int_reg_array_34_11_real;
  assign io_coef_out_payload_0_34_11_imag = int_reg_array_34_11_imag;
  assign io_coef_out_payload_0_34_12_real = int_reg_array_34_12_real;
  assign io_coef_out_payload_0_34_12_imag = int_reg_array_34_12_imag;
  assign io_coef_out_payload_0_34_13_real = int_reg_array_34_13_real;
  assign io_coef_out_payload_0_34_13_imag = int_reg_array_34_13_imag;
  assign io_coef_out_payload_0_34_14_real = int_reg_array_34_14_real;
  assign io_coef_out_payload_0_34_14_imag = int_reg_array_34_14_imag;
  assign io_coef_out_payload_0_34_15_real = int_reg_array_34_15_real;
  assign io_coef_out_payload_0_34_15_imag = int_reg_array_34_15_imag;
  assign io_coef_out_payload_0_34_16_real = int_reg_array_34_16_real;
  assign io_coef_out_payload_0_34_16_imag = int_reg_array_34_16_imag;
  assign io_coef_out_payload_0_34_17_real = int_reg_array_34_17_real;
  assign io_coef_out_payload_0_34_17_imag = int_reg_array_34_17_imag;
  assign io_coef_out_payload_0_34_18_real = int_reg_array_34_18_real;
  assign io_coef_out_payload_0_34_18_imag = int_reg_array_34_18_imag;
  assign io_coef_out_payload_0_34_19_real = int_reg_array_34_19_real;
  assign io_coef_out_payload_0_34_19_imag = int_reg_array_34_19_imag;
  assign io_coef_out_payload_0_34_20_real = int_reg_array_34_20_real;
  assign io_coef_out_payload_0_34_20_imag = int_reg_array_34_20_imag;
  assign io_coef_out_payload_0_34_21_real = int_reg_array_34_21_real;
  assign io_coef_out_payload_0_34_21_imag = int_reg_array_34_21_imag;
  assign io_coef_out_payload_0_34_22_real = int_reg_array_34_22_real;
  assign io_coef_out_payload_0_34_22_imag = int_reg_array_34_22_imag;
  assign io_coef_out_payload_0_34_23_real = int_reg_array_34_23_real;
  assign io_coef_out_payload_0_34_23_imag = int_reg_array_34_23_imag;
  assign io_coef_out_payload_0_34_24_real = int_reg_array_34_24_real;
  assign io_coef_out_payload_0_34_24_imag = int_reg_array_34_24_imag;
  assign io_coef_out_payload_0_34_25_real = int_reg_array_34_25_real;
  assign io_coef_out_payload_0_34_25_imag = int_reg_array_34_25_imag;
  assign io_coef_out_payload_0_34_26_real = int_reg_array_34_26_real;
  assign io_coef_out_payload_0_34_26_imag = int_reg_array_34_26_imag;
  assign io_coef_out_payload_0_34_27_real = int_reg_array_34_27_real;
  assign io_coef_out_payload_0_34_27_imag = int_reg_array_34_27_imag;
  assign io_coef_out_payload_0_34_28_real = int_reg_array_34_28_real;
  assign io_coef_out_payload_0_34_28_imag = int_reg_array_34_28_imag;
  assign io_coef_out_payload_0_34_29_real = int_reg_array_34_29_real;
  assign io_coef_out_payload_0_34_29_imag = int_reg_array_34_29_imag;
  assign io_coef_out_payload_0_34_30_real = int_reg_array_34_30_real;
  assign io_coef_out_payload_0_34_30_imag = int_reg_array_34_30_imag;
  assign io_coef_out_payload_0_34_31_real = int_reg_array_34_31_real;
  assign io_coef_out_payload_0_34_31_imag = int_reg_array_34_31_imag;
  assign io_coef_out_payload_0_34_32_real = int_reg_array_34_32_real;
  assign io_coef_out_payload_0_34_32_imag = int_reg_array_34_32_imag;
  assign io_coef_out_payload_0_34_33_real = int_reg_array_34_33_real;
  assign io_coef_out_payload_0_34_33_imag = int_reg_array_34_33_imag;
  assign io_coef_out_payload_0_34_34_real = int_reg_array_34_34_real;
  assign io_coef_out_payload_0_34_34_imag = int_reg_array_34_34_imag;
  assign io_coef_out_payload_0_34_35_real = int_reg_array_34_35_real;
  assign io_coef_out_payload_0_34_35_imag = int_reg_array_34_35_imag;
  assign io_coef_out_payload_0_34_36_real = int_reg_array_34_36_real;
  assign io_coef_out_payload_0_34_36_imag = int_reg_array_34_36_imag;
  assign io_coef_out_payload_0_34_37_real = int_reg_array_34_37_real;
  assign io_coef_out_payload_0_34_37_imag = int_reg_array_34_37_imag;
  assign io_coef_out_payload_0_34_38_real = int_reg_array_34_38_real;
  assign io_coef_out_payload_0_34_38_imag = int_reg_array_34_38_imag;
  assign io_coef_out_payload_0_34_39_real = int_reg_array_34_39_real;
  assign io_coef_out_payload_0_34_39_imag = int_reg_array_34_39_imag;
  assign io_coef_out_payload_0_34_40_real = int_reg_array_34_40_real;
  assign io_coef_out_payload_0_34_40_imag = int_reg_array_34_40_imag;
  assign io_coef_out_payload_0_34_41_real = int_reg_array_34_41_real;
  assign io_coef_out_payload_0_34_41_imag = int_reg_array_34_41_imag;
  assign io_coef_out_payload_0_34_42_real = int_reg_array_34_42_real;
  assign io_coef_out_payload_0_34_42_imag = int_reg_array_34_42_imag;
  assign io_coef_out_payload_0_34_43_real = int_reg_array_34_43_real;
  assign io_coef_out_payload_0_34_43_imag = int_reg_array_34_43_imag;
  assign io_coef_out_payload_0_34_44_real = int_reg_array_34_44_real;
  assign io_coef_out_payload_0_34_44_imag = int_reg_array_34_44_imag;
  assign io_coef_out_payload_0_34_45_real = int_reg_array_34_45_real;
  assign io_coef_out_payload_0_34_45_imag = int_reg_array_34_45_imag;
  assign io_coef_out_payload_0_34_46_real = int_reg_array_34_46_real;
  assign io_coef_out_payload_0_34_46_imag = int_reg_array_34_46_imag;
  assign io_coef_out_payload_0_34_47_real = int_reg_array_34_47_real;
  assign io_coef_out_payload_0_34_47_imag = int_reg_array_34_47_imag;
  assign io_coef_out_payload_0_34_48_real = int_reg_array_34_48_real;
  assign io_coef_out_payload_0_34_48_imag = int_reg_array_34_48_imag;
  assign io_coef_out_payload_0_34_49_real = int_reg_array_34_49_real;
  assign io_coef_out_payload_0_34_49_imag = int_reg_array_34_49_imag;
  assign io_coef_out_payload_0_35_0_real = int_reg_array_35_0_real;
  assign io_coef_out_payload_0_35_0_imag = int_reg_array_35_0_imag;
  assign io_coef_out_payload_0_35_1_real = int_reg_array_35_1_real;
  assign io_coef_out_payload_0_35_1_imag = int_reg_array_35_1_imag;
  assign io_coef_out_payload_0_35_2_real = int_reg_array_35_2_real;
  assign io_coef_out_payload_0_35_2_imag = int_reg_array_35_2_imag;
  assign io_coef_out_payload_0_35_3_real = int_reg_array_35_3_real;
  assign io_coef_out_payload_0_35_3_imag = int_reg_array_35_3_imag;
  assign io_coef_out_payload_0_35_4_real = int_reg_array_35_4_real;
  assign io_coef_out_payload_0_35_4_imag = int_reg_array_35_4_imag;
  assign io_coef_out_payload_0_35_5_real = int_reg_array_35_5_real;
  assign io_coef_out_payload_0_35_5_imag = int_reg_array_35_5_imag;
  assign io_coef_out_payload_0_35_6_real = int_reg_array_35_6_real;
  assign io_coef_out_payload_0_35_6_imag = int_reg_array_35_6_imag;
  assign io_coef_out_payload_0_35_7_real = int_reg_array_35_7_real;
  assign io_coef_out_payload_0_35_7_imag = int_reg_array_35_7_imag;
  assign io_coef_out_payload_0_35_8_real = int_reg_array_35_8_real;
  assign io_coef_out_payload_0_35_8_imag = int_reg_array_35_8_imag;
  assign io_coef_out_payload_0_35_9_real = int_reg_array_35_9_real;
  assign io_coef_out_payload_0_35_9_imag = int_reg_array_35_9_imag;
  assign io_coef_out_payload_0_35_10_real = int_reg_array_35_10_real;
  assign io_coef_out_payload_0_35_10_imag = int_reg_array_35_10_imag;
  assign io_coef_out_payload_0_35_11_real = int_reg_array_35_11_real;
  assign io_coef_out_payload_0_35_11_imag = int_reg_array_35_11_imag;
  assign io_coef_out_payload_0_35_12_real = int_reg_array_35_12_real;
  assign io_coef_out_payload_0_35_12_imag = int_reg_array_35_12_imag;
  assign io_coef_out_payload_0_35_13_real = int_reg_array_35_13_real;
  assign io_coef_out_payload_0_35_13_imag = int_reg_array_35_13_imag;
  assign io_coef_out_payload_0_35_14_real = int_reg_array_35_14_real;
  assign io_coef_out_payload_0_35_14_imag = int_reg_array_35_14_imag;
  assign io_coef_out_payload_0_35_15_real = int_reg_array_35_15_real;
  assign io_coef_out_payload_0_35_15_imag = int_reg_array_35_15_imag;
  assign io_coef_out_payload_0_35_16_real = int_reg_array_35_16_real;
  assign io_coef_out_payload_0_35_16_imag = int_reg_array_35_16_imag;
  assign io_coef_out_payload_0_35_17_real = int_reg_array_35_17_real;
  assign io_coef_out_payload_0_35_17_imag = int_reg_array_35_17_imag;
  assign io_coef_out_payload_0_35_18_real = int_reg_array_35_18_real;
  assign io_coef_out_payload_0_35_18_imag = int_reg_array_35_18_imag;
  assign io_coef_out_payload_0_35_19_real = int_reg_array_35_19_real;
  assign io_coef_out_payload_0_35_19_imag = int_reg_array_35_19_imag;
  assign io_coef_out_payload_0_35_20_real = int_reg_array_35_20_real;
  assign io_coef_out_payload_0_35_20_imag = int_reg_array_35_20_imag;
  assign io_coef_out_payload_0_35_21_real = int_reg_array_35_21_real;
  assign io_coef_out_payload_0_35_21_imag = int_reg_array_35_21_imag;
  assign io_coef_out_payload_0_35_22_real = int_reg_array_35_22_real;
  assign io_coef_out_payload_0_35_22_imag = int_reg_array_35_22_imag;
  assign io_coef_out_payload_0_35_23_real = int_reg_array_35_23_real;
  assign io_coef_out_payload_0_35_23_imag = int_reg_array_35_23_imag;
  assign io_coef_out_payload_0_35_24_real = int_reg_array_35_24_real;
  assign io_coef_out_payload_0_35_24_imag = int_reg_array_35_24_imag;
  assign io_coef_out_payload_0_35_25_real = int_reg_array_35_25_real;
  assign io_coef_out_payload_0_35_25_imag = int_reg_array_35_25_imag;
  assign io_coef_out_payload_0_35_26_real = int_reg_array_35_26_real;
  assign io_coef_out_payload_0_35_26_imag = int_reg_array_35_26_imag;
  assign io_coef_out_payload_0_35_27_real = int_reg_array_35_27_real;
  assign io_coef_out_payload_0_35_27_imag = int_reg_array_35_27_imag;
  assign io_coef_out_payload_0_35_28_real = int_reg_array_35_28_real;
  assign io_coef_out_payload_0_35_28_imag = int_reg_array_35_28_imag;
  assign io_coef_out_payload_0_35_29_real = int_reg_array_35_29_real;
  assign io_coef_out_payload_0_35_29_imag = int_reg_array_35_29_imag;
  assign io_coef_out_payload_0_35_30_real = int_reg_array_35_30_real;
  assign io_coef_out_payload_0_35_30_imag = int_reg_array_35_30_imag;
  assign io_coef_out_payload_0_35_31_real = int_reg_array_35_31_real;
  assign io_coef_out_payload_0_35_31_imag = int_reg_array_35_31_imag;
  assign io_coef_out_payload_0_35_32_real = int_reg_array_35_32_real;
  assign io_coef_out_payload_0_35_32_imag = int_reg_array_35_32_imag;
  assign io_coef_out_payload_0_35_33_real = int_reg_array_35_33_real;
  assign io_coef_out_payload_0_35_33_imag = int_reg_array_35_33_imag;
  assign io_coef_out_payload_0_35_34_real = int_reg_array_35_34_real;
  assign io_coef_out_payload_0_35_34_imag = int_reg_array_35_34_imag;
  assign io_coef_out_payload_0_35_35_real = int_reg_array_35_35_real;
  assign io_coef_out_payload_0_35_35_imag = int_reg_array_35_35_imag;
  assign io_coef_out_payload_0_35_36_real = int_reg_array_35_36_real;
  assign io_coef_out_payload_0_35_36_imag = int_reg_array_35_36_imag;
  assign io_coef_out_payload_0_35_37_real = int_reg_array_35_37_real;
  assign io_coef_out_payload_0_35_37_imag = int_reg_array_35_37_imag;
  assign io_coef_out_payload_0_35_38_real = int_reg_array_35_38_real;
  assign io_coef_out_payload_0_35_38_imag = int_reg_array_35_38_imag;
  assign io_coef_out_payload_0_35_39_real = int_reg_array_35_39_real;
  assign io_coef_out_payload_0_35_39_imag = int_reg_array_35_39_imag;
  assign io_coef_out_payload_0_35_40_real = int_reg_array_35_40_real;
  assign io_coef_out_payload_0_35_40_imag = int_reg_array_35_40_imag;
  assign io_coef_out_payload_0_35_41_real = int_reg_array_35_41_real;
  assign io_coef_out_payload_0_35_41_imag = int_reg_array_35_41_imag;
  assign io_coef_out_payload_0_35_42_real = int_reg_array_35_42_real;
  assign io_coef_out_payload_0_35_42_imag = int_reg_array_35_42_imag;
  assign io_coef_out_payload_0_35_43_real = int_reg_array_35_43_real;
  assign io_coef_out_payload_0_35_43_imag = int_reg_array_35_43_imag;
  assign io_coef_out_payload_0_35_44_real = int_reg_array_35_44_real;
  assign io_coef_out_payload_0_35_44_imag = int_reg_array_35_44_imag;
  assign io_coef_out_payload_0_35_45_real = int_reg_array_35_45_real;
  assign io_coef_out_payload_0_35_45_imag = int_reg_array_35_45_imag;
  assign io_coef_out_payload_0_35_46_real = int_reg_array_35_46_real;
  assign io_coef_out_payload_0_35_46_imag = int_reg_array_35_46_imag;
  assign io_coef_out_payload_0_35_47_real = int_reg_array_35_47_real;
  assign io_coef_out_payload_0_35_47_imag = int_reg_array_35_47_imag;
  assign io_coef_out_payload_0_35_48_real = int_reg_array_35_48_real;
  assign io_coef_out_payload_0_35_48_imag = int_reg_array_35_48_imag;
  assign io_coef_out_payload_0_35_49_real = int_reg_array_35_49_real;
  assign io_coef_out_payload_0_35_49_imag = int_reg_array_35_49_imag;
  assign io_coef_out_payload_0_36_0_real = int_reg_array_36_0_real;
  assign io_coef_out_payload_0_36_0_imag = int_reg_array_36_0_imag;
  assign io_coef_out_payload_0_36_1_real = int_reg_array_36_1_real;
  assign io_coef_out_payload_0_36_1_imag = int_reg_array_36_1_imag;
  assign io_coef_out_payload_0_36_2_real = int_reg_array_36_2_real;
  assign io_coef_out_payload_0_36_2_imag = int_reg_array_36_2_imag;
  assign io_coef_out_payload_0_36_3_real = int_reg_array_36_3_real;
  assign io_coef_out_payload_0_36_3_imag = int_reg_array_36_3_imag;
  assign io_coef_out_payload_0_36_4_real = int_reg_array_36_4_real;
  assign io_coef_out_payload_0_36_4_imag = int_reg_array_36_4_imag;
  assign io_coef_out_payload_0_36_5_real = int_reg_array_36_5_real;
  assign io_coef_out_payload_0_36_5_imag = int_reg_array_36_5_imag;
  assign io_coef_out_payload_0_36_6_real = int_reg_array_36_6_real;
  assign io_coef_out_payload_0_36_6_imag = int_reg_array_36_6_imag;
  assign io_coef_out_payload_0_36_7_real = int_reg_array_36_7_real;
  assign io_coef_out_payload_0_36_7_imag = int_reg_array_36_7_imag;
  assign io_coef_out_payload_0_36_8_real = int_reg_array_36_8_real;
  assign io_coef_out_payload_0_36_8_imag = int_reg_array_36_8_imag;
  assign io_coef_out_payload_0_36_9_real = int_reg_array_36_9_real;
  assign io_coef_out_payload_0_36_9_imag = int_reg_array_36_9_imag;
  assign io_coef_out_payload_0_36_10_real = int_reg_array_36_10_real;
  assign io_coef_out_payload_0_36_10_imag = int_reg_array_36_10_imag;
  assign io_coef_out_payload_0_36_11_real = int_reg_array_36_11_real;
  assign io_coef_out_payload_0_36_11_imag = int_reg_array_36_11_imag;
  assign io_coef_out_payload_0_36_12_real = int_reg_array_36_12_real;
  assign io_coef_out_payload_0_36_12_imag = int_reg_array_36_12_imag;
  assign io_coef_out_payload_0_36_13_real = int_reg_array_36_13_real;
  assign io_coef_out_payload_0_36_13_imag = int_reg_array_36_13_imag;
  assign io_coef_out_payload_0_36_14_real = int_reg_array_36_14_real;
  assign io_coef_out_payload_0_36_14_imag = int_reg_array_36_14_imag;
  assign io_coef_out_payload_0_36_15_real = int_reg_array_36_15_real;
  assign io_coef_out_payload_0_36_15_imag = int_reg_array_36_15_imag;
  assign io_coef_out_payload_0_36_16_real = int_reg_array_36_16_real;
  assign io_coef_out_payload_0_36_16_imag = int_reg_array_36_16_imag;
  assign io_coef_out_payload_0_36_17_real = int_reg_array_36_17_real;
  assign io_coef_out_payload_0_36_17_imag = int_reg_array_36_17_imag;
  assign io_coef_out_payload_0_36_18_real = int_reg_array_36_18_real;
  assign io_coef_out_payload_0_36_18_imag = int_reg_array_36_18_imag;
  assign io_coef_out_payload_0_36_19_real = int_reg_array_36_19_real;
  assign io_coef_out_payload_0_36_19_imag = int_reg_array_36_19_imag;
  assign io_coef_out_payload_0_36_20_real = int_reg_array_36_20_real;
  assign io_coef_out_payload_0_36_20_imag = int_reg_array_36_20_imag;
  assign io_coef_out_payload_0_36_21_real = int_reg_array_36_21_real;
  assign io_coef_out_payload_0_36_21_imag = int_reg_array_36_21_imag;
  assign io_coef_out_payload_0_36_22_real = int_reg_array_36_22_real;
  assign io_coef_out_payload_0_36_22_imag = int_reg_array_36_22_imag;
  assign io_coef_out_payload_0_36_23_real = int_reg_array_36_23_real;
  assign io_coef_out_payload_0_36_23_imag = int_reg_array_36_23_imag;
  assign io_coef_out_payload_0_36_24_real = int_reg_array_36_24_real;
  assign io_coef_out_payload_0_36_24_imag = int_reg_array_36_24_imag;
  assign io_coef_out_payload_0_36_25_real = int_reg_array_36_25_real;
  assign io_coef_out_payload_0_36_25_imag = int_reg_array_36_25_imag;
  assign io_coef_out_payload_0_36_26_real = int_reg_array_36_26_real;
  assign io_coef_out_payload_0_36_26_imag = int_reg_array_36_26_imag;
  assign io_coef_out_payload_0_36_27_real = int_reg_array_36_27_real;
  assign io_coef_out_payload_0_36_27_imag = int_reg_array_36_27_imag;
  assign io_coef_out_payload_0_36_28_real = int_reg_array_36_28_real;
  assign io_coef_out_payload_0_36_28_imag = int_reg_array_36_28_imag;
  assign io_coef_out_payload_0_36_29_real = int_reg_array_36_29_real;
  assign io_coef_out_payload_0_36_29_imag = int_reg_array_36_29_imag;
  assign io_coef_out_payload_0_36_30_real = int_reg_array_36_30_real;
  assign io_coef_out_payload_0_36_30_imag = int_reg_array_36_30_imag;
  assign io_coef_out_payload_0_36_31_real = int_reg_array_36_31_real;
  assign io_coef_out_payload_0_36_31_imag = int_reg_array_36_31_imag;
  assign io_coef_out_payload_0_36_32_real = int_reg_array_36_32_real;
  assign io_coef_out_payload_0_36_32_imag = int_reg_array_36_32_imag;
  assign io_coef_out_payload_0_36_33_real = int_reg_array_36_33_real;
  assign io_coef_out_payload_0_36_33_imag = int_reg_array_36_33_imag;
  assign io_coef_out_payload_0_36_34_real = int_reg_array_36_34_real;
  assign io_coef_out_payload_0_36_34_imag = int_reg_array_36_34_imag;
  assign io_coef_out_payload_0_36_35_real = int_reg_array_36_35_real;
  assign io_coef_out_payload_0_36_35_imag = int_reg_array_36_35_imag;
  assign io_coef_out_payload_0_36_36_real = int_reg_array_36_36_real;
  assign io_coef_out_payload_0_36_36_imag = int_reg_array_36_36_imag;
  assign io_coef_out_payload_0_36_37_real = int_reg_array_36_37_real;
  assign io_coef_out_payload_0_36_37_imag = int_reg_array_36_37_imag;
  assign io_coef_out_payload_0_36_38_real = int_reg_array_36_38_real;
  assign io_coef_out_payload_0_36_38_imag = int_reg_array_36_38_imag;
  assign io_coef_out_payload_0_36_39_real = int_reg_array_36_39_real;
  assign io_coef_out_payload_0_36_39_imag = int_reg_array_36_39_imag;
  assign io_coef_out_payload_0_36_40_real = int_reg_array_36_40_real;
  assign io_coef_out_payload_0_36_40_imag = int_reg_array_36_40_imag;
  assign io_coef_out_payload_0_36_41_real = int_reg_array_36_41_real;
  assign io_coef_out_payload_0_36_41_imag = int_reg_array_36_41_imag;
  assign io_coef_out_payload_0_36_42_real = int_reg_array_36_42_real;
  assign io_coef_out_payload_0_36_42_imag = int_reg_array_36_42_imag;
  assign io_coef_out_payload_0_36_43_real = int_reg_array_36_43_real;
  assign io_coef_out_payload_0_36_43_imag = int_reg_array_36_43_imag;
  assign io_coef_out_payload_0_36_44_real = int_reg_array_36_44_real;
  assign io_coef_out_payload_0_36_44_imag = int_reg_array_36_44_imag;
  assign io_coef_out_payload_0_36_45_real = int_reg_array_36_45_real;
  assign io_coef_out_payload_0_36_45_imag = int_reg_array_36_45_imag;
  assign io_coef_out_payload_0_36_46_real = int_reg_array_36_46_real;
  assign io_coef_out_payload_0_36_46_imag = int_reg_array_36_46_imag;
  assign io_coef_out_payload_0_36_47_real = int_reg_array_36_47_real;
  assign io_coef_out_payload_0_36_47_imag = int_reg_array_36_47_imag;
  assign io_coef_out_payload_0_36_48_real = int_reg_array_36_48_real;
  assign io_coef_out_payload_0_36_48_imag = int_reg_array_36_48_imag;
  assign io_coef_out_payload_0_36_49_real = int_reg_array_36_49_real;
  assign io_coef_out_payload_0_36_49_imag = int_reg_array_36_49_imag;
  assign io_coef_out_payload_0_37_0_real = int_reg_array_37_0_real;
  assign io_coef_out_payload_0_37_0_imag = int_reg_array_37_0_imag;
  assign io_coef_out_payload_0_37_1_real = int_reg_array_37_1_real;
  assign io_coef_out_payload_0_37_1_imag = int_reg_array_37_1_imag;
  assign io_coef_out_payload_0_37_2_real = int_reg_array_37_2_real;
  assign io_coef_out_payload_0_37_2_imag = int_reg_array_37_2_imag;
  assign io_coef_out_payload_0_37_3_real = int_reg_array_37_3_real;
  assign io_coef_out_payload_0_37_3_imag = int_reg_array_37_3_imag;
  assign io_coef_out_payload_0_37_4_real = int_reg_array_37_4_real;
  assign io_coef_out_payload_0_37_4_imag = int_reg_array_37_4_imag;
  assign io_coef_out_payload_0_37_5_real = int_reg_array_37_5_real;
  assign io_coef_out_payload_0_37_5_imag = int_reg_array_37_5_imag;
  assign io_coef_out_payload_0_37_6_real = int_reg_array_37_6_real;
  assign io_coef_out_payload_0_37_6_imag = int_reg_array_37_6_imag;
  assign io_coef_out_payload_0_37_7_real = int_reg_array_37_7_real;
  assign io_coef_out_payload_0_37_7_imag = int_reg_array_37_7_imag;
  assign io_coef_out_payload_0_37_8_real = int_reg_array_37_8_real;
  assign io_coef_out_payload_0_37_8_imag = int_reg_array_37_8_imag;
  assign io_coef_out_payload_0_37_9_real = int_reg_array_37_9_real;
  assign io_coef_out_payload_0_37_9_imag = int_reg_array_37_9_imag;
  assign io_coef_out_payload_0_37_10_real = int_reg_array_37_10_real;
  assign io_coef_out_payload_0_37_10_imag = int_reg_array_37_10_imag;
  assign io_coef_out_payload_0_37_11_real = int_reg_array_37_11_real;
  assign io_coef_out_payload_0_37_11_imag = int_reg_array_37_11_imag;
  assign io_coef_out_payload_0_37_12_real = int_reg_array_37_12_real;
  assign io_coef_out_payload_0_37_12_imag = int_reg_array_37_12_imag;
  assign io_coef_out_payload_0_37_13_real = int_reg_array_37_13_real;
  assign io_coef_out_payload_0_37_13_imag = int_reg_array_37_13_imag;
  assign io_coef_out_payload_0_37_14_real = int_reg_array_37_14_real;
  assign io_coef_out_payload_0_37_14_imag = int_reg_array_37_14_imag;
  assign io_coef_out_payload_0_37_15_real = int_reg_array_37_15_real;
  assign io_coef_out_payload_0_37_15_imag = int_reg_array_37_15_imag;
  assign io_coef_out_payload_0_37_16_real = int_reg_array_37_16_real;
  assign io_coef_out_payload_0_37_16_imag = int_reg_array_37_16_imag;
  assign io_coef_out_payload_0_37_17_real = int_reg_array_37_17_real;
  assign io_coef_out_payload_0_37_17_imag = int_reg_array_37_17_imag;
  assign io_coef_out_payload_0_37_18_real = int_reg_array_37_18_real;
  assign io_coef_out_payload_0_37_18_imag = int_reg_array_37_18_imag;
  assign io_coef_out_payload_0_37_19_real = int_reg_array_37_19_real;
  assign io_coef_out_payload_0_37_19_imag = int_reg_array_37_19_imag;
  assign io_coef_out_payload_0_37_20_real = int_reg_array_37_20_real;
  assign io_coef_out_payload_0_37_20_imag = int_reg_array_37_20_imag;
  assign io_coef_out_payload_0_37_21_real = int_reg_array_37_21_real;
  assign io_coef_out_payload_0_37_21_imag = int_reg_array_37_21_imag;
  assign io_coef_out_payload_0_37_22_real = int_reg_array_37_22_real;
  assign io_coef_out_payload_0_37_22_imag = int_reg_array_37_22_imag;
  assign io_coef_out_payload_0_37_23_real = int_reg_array_37_23_real;
  assign io_coef_out_payload_0_37_23_imag = int_reg_array_37_23_imag;
  assign io_coef_out_payload_0_37_24_real = int_reg_array_37_24_real;
  assign io_coef_out_payload_0_37_24_imag = int_reg_array_37_24_imag;
  assign io_coef_out_payload_0_37_25_real = int_reg_array_37_25_real;
  assign io_coef_out_payload_0_37_25_imag = int_reg_array_37_25_imag;
  assign io_coef_out_payload_0_37_26_real = int_reg_array_37_26_real;
  assign io_coef_out_payload_0_37_26_imag = int_reg_array_37_26_imag;
  assign io_coef_out_payload_0_37_27_real = int_reg_array_37_27_real;
  assign io_coef_out_payload_0_37_27_imag = int_reg_array_37_27_imag;
  assign io_coef_out_payload_0_37_28_real = int_reg_array_37_28_real;
  assign io_coef_out_payload_0_37_28_imag = int_reg_array_37_28_imag;
  assign io_coef_out_payload_0_37_29_real = int_reg_array_37_29_real;
  assign io_coef_out_payload_0_37_29_imag = int_reg_array_37_29_imag;
  assign io_coef_out_payload_0_37_30_real = int_reg_array_37_30_real;
  assign io_coef_out_payload_0_37_30_imag = int_reg_array_37_30_imag;
  assign io_coef_out_payload_0_37_31_real = int_reg_array_37_31_real;
  assign io_coef_out_payload_0_37_31_imag = int_reg_array_37_31_imag;
  assign io_coef_out_payload_0_37_32_real = int_reg_array_37_32_real;
  assign io_coef_out_payload_0_37_32_imag = int_reg_array_37_32_imag;
  assign io_coef_out_payload_0_37_33_real = int_reg_array_37_33_real;
  assign io_coef_out_payload_0_37_33_imag = int_reg_array_37_33_imag;
  assign io_coef_out_payload_0_37_34_real = int_reg_array_37_34_real;
  assign io_coef_out_payload_0_37_34_imag = int_reg_array_37_34_imag;
  assign io_coef_out_payload_0_37_35_real = int_reg_array_37_35_real;
  assign io_coef_out_payload_0_37_35_imag = int_reg_array_37_35_imag;
  assign io_coef_out_payload_0_37_36_real = int_reg_array_37_36_real;
  assign io_coef_out_payload_0_37_36_imag = int_reg_array_37_36_imag;
  assign io_coef_out_payload_0_37_37_real = int_reg_array_37_37_real;
  assign io_coef_out_payload_0_37_37_imag = int_reg_array_37_37_imag;
  assign io_coef_out_payload_0_37_38_real = int_reg_array_37_38_real;
  assign io_coef_out_payload_0_37_38_imag = int_reg_array_37_38_imag;
  assign io_coef_out_payload_0_37_39_real = int_reg_array_37_39_real;
  assign io_coef_out_payload_0_37_39_imag = int_reg_array_37_39_imag;
  assign io_coef_out_payload_0_37_40_real = int_reg_array_37_40_real;
  assign io_coef_out_payload_0_37_40_imag = int_reg_array_37_40_imag;
  assign io_coef_out_payload_0_37_41_real = int_reg_array_37_41_real;
  assign io_coef_out_payload_0_37_41_imag = int_reg_array_37_41_imag;
  assign io_coef_out_payload_0_37_42_real = int_reg_array_37_42_real;
  assign io_coef_out_payload_0_37_42_imag = int_reg_array_37_42_imag;
  assign io_coef_out_payload_0_37_43_real = int_reg_array_37_43_real;
  assign io_coef_out_payload_0_37_43_imag = int_reg_array_37_43_imag;
  assign io_coef_out_payload_0_37_44_real = int_reg_array_37_44_real;
  assign io_coef_out_payload_0_37_44_imag = int_reg_array_37_44_imag;
  assign io_coef_out_payload_0_37_45_real = int_reg_array_37_45_real;
  assign io_coef_out_payload_0_37_45_imag = int_reg_array_37_45_imag;
  assign io_coef_out_payload_0_37_46_real = int_reg_array_37_46_real;
  assign io_coef_out_payload_0_37_46_imag = int_reg_array_37_46_imag;
  assign io_coef_out_payload_0_37_47_real = int_reg_array_37_47_real;
  assign io_coef_out_payload_0_37_47_imag = int_reg_array_37_47_imag;
  assign io_coef_out_payload_0_37_48_real = int_reg_array_37_48_real;
  assign io_coef_out_payload_0_37_48_imag = int_reg_array_37_48_imag;
  assign io_coef_out_payload_0_37_49_real = int_reg_array_37_49_real;
  assign io_coef_out_payload_0_37_49_imag = int_reg_array_37_49_imag;
  assign io_coef_out_payload_0_38_0_real = int_reg_array_38_0_real;
  assign io_coef_out_payload_0_38_0_imag = int_reg_array_38_0_imag;
  assign io_coef_out_payload_0_38_1_real = int_reg_array_38_1_real;
  assign io_coef_out_payload_0_38_1_imag = int_reg_array_38_1_imag;
  assign io_coef_out_payload_0_38_2_real = int_reg_array_38_2_real;
  assign io_coef_out_payload_0_38_2_imag = int_reg_array_38_2_imag;
  assign io_coef_out_payload_0_38_3_real = int_reg_array_38_3_real;
  assign io_coef_out_payload_0_38_3_imag = int_reg_array_38_3_imag;
  assign io_coef_out_payload_0_38_4_real = int_reg_array_38_4_real;
  assign io_coef_out_payload_0_38_4_imag = int_reg_array_38_4_imag;
  assign io_coef_out_payload_0_38_5_real = int_reg_array_38_5_real;
  assign io_coef_out_payload_0_38_5_imag = int_reg_array_38_5_imag;
  assign io_coef_out_payload_0_38_6_real = int_reg_array_38_6_real;
  assign io_coef_out_payload_0_38_6_imag = int_reg_array_38_6_imag;
  assign io_coef_out_payload_0_38_7_real = int_reg_array_38_7_real;
  assign io_coef_out_payload_0_38_7_imag = int_reg_array_38_7_imag;
  assign io_coef_out_payload_0_38_8_real = int_reg_array_38_8_real;
  assign io_coef_out_payload_0_38_8_imag = int_reg_array_38_8_imag;
  assign io_coef_out_payload_0_38_9_real = int_reg_array_38_9_real;
  assign io_coef_out_payload_0_38_9_imag = int_reg_array_38_9_imag;
  assign io_coef_out_payload_0_38_10_real = int_reg_array_38_10_real;
  assign io_coef_out_payload_0_38_10_imag = int_reg_array_38_10_imag;
  assign io_coef_out_payload_0_38_11_real = int_reg_array_38_11_real;
  assign io_coef_out_payload_0_38_11_imag = int_reg_array_38_11_imag;
  assign io_coef_out_payload_0_38_12_real = int_reg_array_38_12_real;
  assign io_coef_out_payload_0_38_12_imag = int_reg_array_38_12_imag;
  assign io_coef_out_payload_0_38_13_real = int_reg_array_38_13_real;
  assign io_coef_out_payload_0_38_13_imag = int_reg_array_38_13_imag;
  assign io_coef_out_payload_0_38_14_real = int_reg_array_38_14_real;
  assign io_coef_out_payload_0_38_14_imag = int_reg_array_38_14_imag;
  assign io_coef_out_payload_0_38_15_real = int_reg_array_38_15_real;
  assign io_coef_out_payload_0_38_15_imag = int_reg_array_38_15_imag;
  assign io_coef_out_payload_0_38_16_real = int_reg_array_38_16_real;
  assign io_coef_out_payload_0_38_16_imag = int_reg_array_38_16_imag;
  assign io_coef_out_payload_0_38_17_real = int_reg_array_38_17_real;
  assign io_coef_out_payload_0_38_17_imag = int_reg_array_38_17_imag;
  assign io_coef_out_payload_0_38_18_real = int_reg_array_38_18_real;
  assign io_coef_out_payload_0_38_18_imag = int_reg_array_38_18_imag;
  assign io_coef_out_payload_0_38_19_real = int_reg_array_38_19_real;
  assign io_coef_out_payload_0_38_19_imag = int_reg_array_38_19_imag;
  assign io_coef_out_payload_0_38_20_real = int_reg_array_38_20_real;
  assign io_coef_out_payload_0_38_20_imag = int_reg_array_38_20_imag;
  assign io_coef_out_payload_0_38_21_real = int_reg_array_38_21_real;
  assign io_coef_out_payload_0_38_21_imag = int_reg_array_38_21_imag;
  assign io_coef_out_payload_0_38_22_real = int_reg_array_38_22_real;
  assign io_coef_out_payload_0_38_22_imag = int_reg_array_38_22_imag;
  assign io_coef_out_payload_0_38_23_real = int_reg_array_38_23_real;
  assign io_coef_out_payload_0_38_23_imag = int_reg_array_38_23_imag;
  assign io_coef_out_payload_0_38_24_real = int_reg_array_38_24_real;
  assign io_coef_out_payload_0_38_24_imag = int_reg_array_38_24_imag;
  assign io_coef_out_payload_0_38_25_real = int_reg_array_38_25_real;
  assign io_coef_out_payload_0_38_25_imag = int_reg_array_38_25_imag;
  assign io_coef_out_payload_0_38_26_real = int_reg_array_38_26_real;
  assign io_coef_out_payload_0_38_26_imag = int_reg_array_38_26_imag;
  assign io_coef_out_payload_0_38_27_real = int_reg_array_38_27_real;
  assign io_coef_out_payload_0_38_27_imag = int_reg_array_38_27_imag;
  assign io_coef_out_payload_0_38_28_real = int_reg_array_38_28_real;
  assign io_coef_out_payload_0_38_28_imag = int_reg_array_38_28_imag;
  assign io_coef_out_payload_0_38_29_real = int_reg_array_38_29_real;
  assign io_coef_out_payload_0_38_29_imag = int_reg_array_38_29_imag;
  assign io_coef_out_payload_0_38_30_real = int_reg_array_38_30_real;
  assign io_coef_out_payload_0_38_30_imag = int_reg_array_38_30_imag;
  assign io_coef_out_payload_0_38_31_real = int_reg_array_38_31_real;
  assign io_coef_out_payload_0_38_31_imag = int_reg_array_38_31_imag;
  assign io_coef_out_payload_0_38_32_real = int_reg_array_38_32_real;
  assign io_coef_out_payload_0_38_32_imag = int_reg_array_38_32_imag;
  assign io_coef_out_payload_0_38_33_real = int_reg_array_38_33_real;
  assign io_coef_out_payload_0_38_33_imag = int_reg_array_38_33_imag;
  assign io_coef_out_payload_0_38_34_real = int_reg_array_38_34_real;
  assign io_coef_out_payload_0_38_34_imag = int_reg_array_38_34_imag;
  assign io_coef_out_payload_0_38_35_real = int_reg_array_38_35_real;
  assign io_coef_out_payload_0_38_35_imag = int_reg_array_38_35_imag;
  assign io_coef_out_payload_0_38_36_real = int_reg_array_38_36_real;
  assign io_coef_out_payload_0_38_36_imag = int_reg_array_38_36_imag;
  assign io_coef_out_payload_0_38_37_real = int_reg_array_38_37_real;
  assign io_coef_out_payload_0_38_37_imag = int_reg_array_38_37_imag;
  assign io_coef_out_payload_0_38_38_real = int_reg_array_38_38_real;
  assign io_coef_out_payload_0_38_38_imag = int_reg_array_38_38_imag;
  assign io_coef_out_payload_0_38_39_real = int_reg_array_38_39_real;
  assign io_coef_out_payload_0_38_39_imag = int_reg_array_38_39_imag;
  assign io_coef_out_payload_0_38_40_real = int_reg_array_38_40_real;
  assign io_coef_out_payload_0_38_40_imag = int_reg_array_38_40_imag;
  assign io_coef_out_payload_0_38_41_real = int_reg_array_38_41_real;
  assign io_coef_out_payload_0_38_41_imag = int_reg_array_38_41_imag;
  assign io_coef_out_payload_0_38_42_real = int_reg_array_38_42_real;
  assign io_coef_out_payload_0_38_42_imag = int_reg_array_38_42_imag;
  assign io_coef_out_payload_0_38_43_real = int_reg_array_38_43_real;
  assign io_coef_out_payload_0_38_43_imag = int_reg_array_38_43_imag;
  assign io_coef_out_payload_0_38_44_real = int_reg_array_38_44_real;
  assign io_coef_out_payload_0_38_44_imag = int_reg_array_38_44_imag;
  assign io_coef_out_payload_0_38_45_real = int_reg_array_38_45_real;
  assign io_coef_out_payload_0_38_45_imag = int_reg_array_38_45_imag;
  assign io_coef_out_payload_0_38_46_real = int_reg_array_38_46_real;
  assign io_coef_out_payload_0_38_46_imag = int_reg_array_38_46_imag;
  assign io_coef_out_payload_0_38_47_real = int_reg_array_38_47_real;
  assign io_coef_out_payload_0_38_47_imag = int_reg_array_38_47_imag;
  assign io_coef_out_payload_0_38_48_real = int_reg_array_38_48_real;
  assign io_coef_out_payload_0_38_48_imag = int_reg_array_38_48_imag;
  assign io_coef_out_payload_0_38_49_real = int_reg_array_38_49_real;
  assign io_coef_out_payload_0_38_49_imag = int_reg_array_38_49_imag;
  assign io_coef_out_payload_0_39_0_real = int_reg_array_39_0_real;
  assign io_coef_out_payload_0_39_0_imag = int_reg_array_39_0_imag;
  assign io_coef_out_payload_0_39_1_real = int_reg_array_39_1_real;
  assign io_coef_out_payload_0_39_1_imag = int_reg_array_39_1_imag;
  assign io_coef_out_payload_0_39_2_real = int_reg_array_39_2_real;
  assign io_coef_out_payload_0_39_2_imag = int_reg_array_39_2_imag;
  assign io_coef_out_payload_0_39_3_real = int_reg_array_39_3_real;
  assign io_coef_out_payload_0_39_3_imag = int_reg_array_39_3_imag;
  assign io_coef_out_payload_0_39_4_real = int_reg_array_39_4_real;
  assign io_coef_out_payload_0_39_4_imag = int_reg_array_39_4_imag;
  assign io_coef_out_payload_0_39_5_real = int_reg_array_39_5_real;
  assign io_coef_out_payload_0_39_5_imag = int_reg_array_39_5_imag;
  assign io_coef_out_payload_0_39_6_real = int_reg_array_39_6_real;
  assign io_coef_out_payload_0_39_6_imag = int_reg_array_39_6_imag;
  assign io_coef_out_payload_0_39_7_real = int_reg_array_39_7_real;
  assign io_coef_out_payload_0_39_7_imag = int_reg_array_39_7_imag;
  assign io_coef_out_payload_0_39_8_real = int_reg_array_39_8_real;
  assign io_coef_out_payload_0_39_8_imag = int_reg_array_39_8_imag;
  assign io_coef_out_payload_0_39_9_real = int_reg_array_39_9_real;
  assign io_coef_out_payload_0_39_9_imag = int_reg_array_39_9_imag;
  assign io_coef_out_payload_0_39_10_real = int_reg_array_39_10_real;
  assign io_coef_out_payload_0_39_10_imag = int_reg_array_39_10_imag;
  assign io_coef_out_payload_0_39_11_real = int_reg_array_39_11_real;
  assign io_coef_out_payload_0_39_11_imag = int_reg_array_39_11_imag;
  assign io_coef_out_payload_0_39_12_real = int_reg_array_39_12_real;
  assign io_coef_out_payload_0_39_12_imag = int_reg_array_39_12_imag;
  assign io_coef_out_payload_0_39_13_real = int_reg_array_39_13_real;
  assign io_coef_out_payload_0_39_13_imag = int_reg_array_39_13_imag;
  assign io_coef_out_payload_0_39_14_real = int_reg_array_39_14_real;
  assign io_coef_out_payload_0_39_14_imag = int_reg_array_39_14_imag;
  assign io_coef_out_payload_0_39_15_real = int_reg_array_39_15_real;
  assign io_coef_out_payload_0_39_15_imag = int_reg_array_39_15_imag;
  assign io_coef_out_payload_0_39_16_real = int_reg_array_39_16_real;
  assign io_coef_out_payload_0_39_16_imag = int_reg_array_39_16_imag;
  assign io_coef_out_payload_0_39_17_real = int_reg_array_39_17_real;
  assign io_coef_out_payload_0_39_17_imag = int_reg_array_39_17_imag;
  assign io_coef_out_payload_0_39_18_real = int_reg_array_39_18_real;
  assign io_coef_out_payload_0_39_18_imag = int_reg_array_39_18_imag;
  assign io_coef_out_payload_0_39_19_real = int_reg_array_39_19_real;
  assign io_coef_out_payload_0_39_19_imag = int_reg_array_39_19_imag;
  assign io_coef_out_payload_0_39_20_real = int_reg_array_39_20_real;
  assign io_coef_out_payload_0_39_20_imag = int_reg_array_39_20_imag;
  assign io_coef_out_payload_0_39_21_real = int_reg_array_39_21_real;
  assign io_coef_out_payload_0_39_21_imag = int_reg_array_39_21_imag;
  assign io_coef_out_payload_0_39_22_real = int_reg_array_39_22_real;
  assign io_coef_out_payload_0_39_22_imag = int_reg_array_39_22_imag;
  assign io_coef_out_payload_0_39_23_real = int_reg_array_39_23_real;
  assign io_coef_out_payload_0_39_23_imag = int_reg_array_39_23_imag;
  assign io_coef_out_payload_0_39_24_real = int_reg_array_39_24_real;
  assign io_coef_out_payload_0_39_24_imag = int_reg_array_39_24_imag;
  assign io_coef_out_payload_0_39_25_real = int_reg_array_39_25_real;
  assign io_coef_out_payload_0_39_25_imag = int_reg_array_39_25_imag;
  assign io_coef_out_payload_0_39_26_real = int_reg_array_39_26_real;
  assign io_coef_out_payload_0_39_26_imag = int_reg_array_39_26_imag;
  assign io_coef_out_payload_0_39_27_real = int_reg_array_39_27_real;
  assign io_coef_out_payload_0_39_27_imag = int_reg_array_39_27_imag;
  assign io_coef_out_payload_0_39_28_real = int_reg_array_39_28_real;
  assign io_coef_out_payload_0_39_28_imag = int_reg_array_39_28_imag;
  assign io_coef_out_payload_0_39_29_real = int_reg_array_39_29_real;
  assign io_coef_out_payload_0_39_29_imag = int_reg_array_39_29_imag;
  assign io_coef_out_payload_0_39_30_real = int_reg_array_39_30_real;
  assign io_coef_out_payload_0_39_30_imag = int_reg_array_39_30_imag;
  assign io_coef_out_payload_0_39_31_real = int_reg_array_39_31_real;
  assign io_coef_out_payload_0_39_31_imag = int_reg_array_39_31_imag;
  assign io_coef_out_payload_0_39_32_real = int_reg_array_39_32_real;
  assign io_coef_out_payload_0_39_32_imag = int_reg_array_39_32_imag;
  assign io_coef_out_payload_0_39_33_real = int_reg_array_39_33_real;
  assign io_coef_out_payload_0_39_33_imag = int_reg_array_39_33_imag;
  assign io_coef_out_payload_0_39_34_real = int_reg_array_39_34_real;
  assign io_coef_out_payload_0_39_34_imag = int_reg_array_39_34_imag;
  assign io_coef_out_payload_0_39_35_real = int_reg_array_39_35_real;
  assign io_coef_out_payload_0_39_35_imag = int_reg_array_39_35_imag;
  assign io_coef_out_payload_0_39_36_real = int_reg_array_39_36_real;
  assign io_coef_out_payload_0_39_36_imag = int_reg_array_39_36_imag;
  assign io_coef_out_payload_0_39_37_real = int_reg_array_39_37_real;
  assign io_coef_out_payload_0_39_37_imag = int_reg_array_39_37_imag;
  assign io_coef_out_payload_0_39_38_real = int_reg_array_39_38_real;
  assign io_coef_out_payload_0_39_38_imag = int_reg_array_39_38_imag;
  assign io_coef_out_payload_0_39_39_real = int_reg_array_39_39_real;
  assign io_coef_out_payload_0_39_39_imag = int_reg_array_39_39_imag;
  assign io_coef_out_payload_0_39_40_real = int_reg_array_39_40_real;
  assign io_coef_out_payload_0_39_40_imag = int_reg_array_39_40_imag;
  assign io_coef_out_payload_0_39_41_real = int_reg_array_39_41_real;
  assign io_coef_out_payload_0_39_41_imag = int_reg_array_39_41_imag;
  assign io_coef_out_payload_0_39_42_real = int_reg_array_39_42_real;
  assign io_coef_out_payload_0_39_42_imag = int_reg_array_39_42_imag;
  assign io_coef_out_payload_0_39_43_real = int_reg_array_39_43_real;
  assign io_coef_out_payload_0_39_43_imag = int_reg_array_39_43_imag;
  assign io_coef_out_payload_0_39_44_real = int_reg_array_39_44_real;
  assign io_coef_out_payload_0_39_44_imag = int_reg_array_39_44_imag;
  assign io_coef_out_payload_0_39_45_real = int_reg_array_39_45_real;
  assign io_coef_out_payload_0_39_45_imag = int_reg_array_39_45_imag;
  assign io_coef_out_payload_0_39_46_real = int_reg_array_39_46_real;
  assign io_coef_out_payload_0_39_46_imag = int_reg_array_39_46_imag;
  assign io_coef_out_payload_0_39_47_real = int_reg_array_39_47_real;
  assign io_coef_out_payload_0_39_47_imag = int_reg_array_39_47_imag;
  assign io_coef_out_payload_0_39_48_real = int_reg_array_39_48_real;
  assign io_coef_out_payload_0_39_48_imag = int_reg_array_39_48_imag;
  assign io_coef_out_payload_0_39_49_real = int_reg_array_39_49_real;
  assign io_coef_out_payload_0_39_49_imag = int_reg_array_39_49_imag;
  assign io_coef_out_payload_0_40_0_real = int_reg_array_40_0_real;
  assign io_coef_out_payload_0_40_0_imag = int_reg_array_40_0_imag;
  assign io_coef_out_payload_0_40_1_real = int_reg_array_40_1_real;
  assign io_coef_out_payload_0_40_1_imag = int_reg_array_40_1_imag;
  assign io_coef_out_payload_0_40_2_real = int_reg_array_40_2_real;
  assign io_coef_out_payload_0_40_2_imag = int_reg_array_40_2_imag;
  assign io_coef_out_payload_0_40_3_real = int_reg_array_40_3_real;
  assign io_coef_out_payload_0_40_3_imag = int_reg_array_40_3_imag;
  assign io_coef_out_payload_0_40_4_real = int_reg_array_40_4_real;
  assign io_coef_out_payload_0_40_4_imag = int_reg_array_40_4_imag;
  assign io_coef_out_payload_0_40_5_real = int_reg_array_40_5_real;
  assign io_coef_out_payload_0_40_5_imag = int_reg_array_40_5_imag;
  assign io_coef_out_payload_0_40_6_real = int_reg_array_40_6_real;
  assign io_coef_out_payload_0_40_6_imag = int_reg_array_40_6_imag;
  assign io_coef_out_payload_0_40_7_real = int_reg_array_40_7_real;
  assign io_coef_out_payload_0_40_7_imag = int_reg_array_40_7_imag;
  assign io_coef_out_payload_0_40_8_real = int_reg_array_40_8_real;
  assign io_coef_out_payload_0_40_8_imag = int_reg_array_40_8_imag;
  assign io_coef_out_payload_0_40_9_real = int_reg_array_40_9_real;
  assign io_coef_out_payload_0_40_9_imag = int_reg_array_40_9_imag;
  assign io_coef_out_payload_0_40_10_real = int_reg_array_40_10_real;
  assign io_coef_out_payload_0_40_10_imag = int_reg_array_40_10_imag;
  assign io_coef_out_payload_0_40_11_real = int_reg_array_40_11_real;
  assign io_coef_out_payload_0_40_11_imag = int_reg_array_40_11_imag;
  assign io_coef_out_payload_0_40_12_real = int_reg_array_40_12_real;
  assign io_coef_out_payload_0_40_12_imag = int_reg_array_40_12_imag;
  assign io_coef_out_payload_0_40_13_real = int_reg_array_40_13_real;
  assign io_coef_out_payload_0_40_13_imag = int_reg_array_40_13_imag;
  assign io_coef_out_payload_0_40_14_real = int_reg_array_40_14_real;
  assign io_coef_out_payload_0_40_14_imag = int_reg_array_40_14_imag;
  assign io_coef_out_payload_0_40_15_real = int_reg_array_40_15_real;
  assign io_coef_out_payload_0_40_15_imag = int_reg_array_40_15_imag;
  assign io_coef_out_payload_0_40_16_real = int_reg_array_40_16_real;
  assign io_coef_out_payload_0_40_16_imag = int_reg_array_40_16_imag;
  assign io_coef_out_payload_0_40_17_real = int_reg_array_40_17_real;
  assign io_coef_out_payload_0_40_17_imag = int_reg_array_40_17_imag;
  assign io_coef_out_payload_0_40_18_real = int_reg_array_40_18_real;
  assign io_coef_out_payload_0_40_18_imag = int_reg_array_40_18_imag;
  assign io_coef_out_payload_0_40_19_real = int_reg_array_40_19_real;
  assign io_coef_out_payload_0_40_19_imag = int_reg_array_40_19_imag;
  assign io_coef_out_payload_0_40_20_real = int_reg_array_40_20_real;
  assign io_coef_out_payload_0_40_20_imag = int_reg_array_40_20_imag;
  assign io_coef_out_payload_0_40_21_real = int_reg_array_40_21_real;
  assign io_coef_out_payload_0_40_21_imag = int_reg_array_40_21_imag;
  assign io_coef_out_payload_0_40_22_real = int_reg_array_40_22_real;
  assign io_coef_out_payload_0_40_22_imag = int_reg_array_40_22_imag;
  assign io_coef_out_payload_0_40_23_real = int_reg_array_40_23_real;
  assign io_coef_out_payload_0_40_23_imag = int_reg_array_40_23_imag;
  assign io_coef_out_payload_0_40_24_real = int_reg_array_40_24_real;
  assign io_coef_out_payload_0_40_24_imag = int_reg_array_40_24_imag;
  assign io_coef_out_payload_0_40_25_real = int_reg_array_40_25_real;
  assign io_coef_out_payload_0_40_25_imag = int_reg_array_40_25_imag;
  assign io_coef_out_payload_0_40_26_real = int_reg_array_40_26_real;
  assign io_coef_out_payload_0_40_26_imag = int_reg_array_40_26_imag;
  assign io_coef_out_payload_0_40_27_real = int_reg_array_40_27_real;
  assign io_coef_out_payload_0_40_27_imag = int_reg_array_40_27_imag;
  assign io_coef_out_payload_0_40_28_real = int_reg_array_40_28_real;
  assign io_coef_out_payload_0_40_28_imag = int_reg_array_40_28_imag;
  assign io_coef_out_payload_0_40_29_real = int_reg_array_40_29_real;
  assign io_coef_out_payload_0_40_29_imag = int_reg_array_40_29_imag;
  assign io_coef_out_payload_0_40_30_real = int_reg_array_40_30_real;
  assign io_coef_out_payload_0_40_30_imag = int_reg_array_40_30_imag;
  assign io_coef_out_payload_0_40_31_real = int_reg_array_40_31_real;
  assign io_coef_out_payload_0_40_31_imag = int_reg_array_40_31_imag;
  assign io_coef_out_payload_0_40_32_real = int_reg_array_40_32_real;
  assign io_coef_out_payload_0_40_32_imag = int_reg_array_40_32_imag;
  assign io_coef_out_payload_0_40_33_real = int_reg_array_40_33_real;
  assign io_coef_out_payload_0_40_33_imag = int_reg_array_40_33_imag;
  assign io_coef_out_payload_0_40_34_real = int_reg_array_40_34_real;
  assign io_coef_out_payload_0_40_34_imag = int_reg_array_40_34_imag;
  assign io_coef_out_payload_0_40_35_real = int_reg_array_40_35_real;
  assign io_coef_out_payload_0_40_35_imag = int_reg_array_40_35_imag;
  assign io_coef_out_payload_0_40_36_real = int_reg_array_40_36_real;
  assign io_coef_out_payload_0_40_36_imag = int_reg_array_40_36_imag;
  assign io_coef_out_payload_0_40_37_real = int_reg_array_40_37_real;
  assign io_coef_out_payload_0_40_37_imag = int_reg_array_40_37_imag;
  assign io_coef_out_payload_0_40_38_real = int_reg_array_40_38_real;
  assign io_coef_out_payload_0_40_38_imag = int_reg_array_40_38_imag;
  assign io_coef_out_payload_0_40_39_real = int_reg_array_40_39_real;
  assign io_coef_out_payload_0_40_39_imag = int_reg_array_40_39_imag;
  assign io_coef_out_payload_0_40_40_real = int_reg_array_40_40_real;
  assign io_coef_out_payload_0_40_40_imag = int_reg_array_40_40_imag;
  assign io_coef_out_payload_0_40_41_real = int_reg_array_40_41_real;
  assign io_coef_out_payload_0_40_41_imag = int_reg_array_40_41_imag;
  assign io_coef_out_payload_0_40_42_real = int_reg_array_40_42_real;
  assign io_coef_out_payload_0_40_42_imag = int_reg_array_40_42_imag;
  assign io_coef_out_payload_0_40_43_real = int_reg_array_40_43_real;
  assign io_coef_out_payload_0_40_43_imag = int_reg_array_40_43_imag;
  assign io_coef_out_payload_0_40_44_real = int_reg_array_40_44_real;
  assign io_coef_out_payload_0_40_44_imag = int_reg_array_40_44_imag;
  assign io_coef_out_payload_0_40_45_real = int_reg_array_40_45_real;
  assign io_coef_out_payload_0_40_45_imag = int_reg_array_40_45_imag;
  assign io_coef_out_payload_0_40_46_real = int_reg_array_40_46_real;
  assign io_coef_out_payload_0_40_46_imag = int_reg_array_40_46_imag;
  assign io_coef_out_payload_0_40_47_real = int_reg_array_40_47_real;
  assign io_coef_out_payload_0_40_47_imag = int_reg_array_40_47_imag;
  assign io_coef_out_payload_0_40_48_real = int_reg_array_40_48_real;
  assign io_coef_out_payload_0_40_48_imag = int_reg_array_40_48_imag;
  assign io_coef_out_payload_0_40_49_real = int_reg_array_40_49_real;
  assign io_coef_out_payload_0_40_49_imag = int_reg_array_40_49_imag;
  assign io_coef_out_payload_0_41_0_real = int_reg_array_41_0_real;
  assign io_coef_out_payload_0_41_0_imag = int_reg_array_41_0_imag;
  assign io_coef_out_payload_0_41_1_real = int_reg_array_41_1_real;
  assign io_coef_out_payload_0_41_1_imag = int_reg_array_41_1_imag;
  assign io_coef_out_payload_0_41_2_real = int_reg_array_41_2_real;
  assign io_coef_out_payload_0_41_2_imag = int_reg_array_41_2_imag;
  assign io_coef_out_payload_0_41_3_real = int_reg_array_41_3_real;
  assign io_coef_out_payload_0_41_3_imag = int_reg_array_41_3_imag;
  assign io_coef_out_payload_0_41_4_real = int_reg_array_41_4_real;
  assign io_coef_out_payload_0_41_4_imag = int_reg_array_41_4_imag;
  assign io_coef_out_payload_0_41_5_real = int_reg_array_41_5_real;
  assign io_coef_out_payload_0_41_5_imag = int_reg_array_41_5_imag;
  assign io_coef_out_payload_0_41_6_real = int_reg_array_41_6_real;
  assign io_coef_out_payload_0_41_6_imag = int_reg_array_41_6_imag;
  assign io_coef_out_payload_0_41_7_real = int_reg_array_41_7_real;
  assign io_coef_out_payload_0_41_7_imag = int_reg_array_41_7_imag;
  assign io_coef_out_payload_0_41_8_real = int_reg_array_41_8_real;
  assign io_coef_out_payload_0_41_8_imag = int_reg_array_41_8_imag;
  assign io_coef_out_payload_0_41_9_real = int_reg_array_41_9_real;
  assign io_coef_out_payload_0_41_9_imag = int_reg_array_41_9_imag;
  assign io_coef_out_payload_0_41_10_real = int_reg_array_41_10_real;
  assign io_coef_out_payload_0_41_10_imag = int_reg_array_41_10_imag;
  assign io_coef_out_payload_0_41_11_real = int_reg_array_41_11_real;
  assign io_coef_out_payload_0_41_11_imag = int_reg_array_41_11_imag;
  assign io_coef_out_payload_0_41_12_real = int_reg_array_41_12_real;
  assign io_coef_out_payload_0_41_12_imag = int_reg_array_41_12_imag;
  assign io_coef_out_payload_0_41_13_real = int_reg_array_41_13_real;
  assign io_coef_out_payload_0_41_13_imag = int_reg_array_41_13_imag;
  assign io_coef_out_payload_0_41_14_real = int_reg_array_41_14_real;
  assign io_coef_out_payload_0_41_14_imag = int_reg_array_41_14_imag;
  assign io_coef_out_payload_0_41_15_real = int_reg_array_41_15_real;
  assign io_coef_out_payload_0_41_15_imag = int_reg_array_41_15_imag;
  assign io_coef_out_payload_0_41_16_real = int_reg_array_41_16_real;
  assign io_coef_out_payload_0_41_16_imag = int_reg_array_41_16_imag;
  assign io_coef_out_payload_0_41_17_real = int_reg_array_41_17_real;
  assign io_coef_out_payload_0_41_17_imag = int_reg_array_41_17_imag;
  assign io_coef_out_payload_0_41_18_real = int_reg_array_41_18_real;
  assign io_coef_out_payload_0_41_18_imag = int_reg_array_41_18_imag;
  assign io_coef_out_payload_0_41_19_real = int_reg_array_41_19_real;
  assign io_coef_out_payload_0_41_19_imag = int_reg_array_41_19_imag;
  assign io_coef_out_payload_0_41_20_real = int_reg_array_41_20_real;
  assign io_coef_out_payload_0_41_20_imag = int_reg_array_41_20_imag;
  assign io_coef_out_payload_0_41_21_real = int_reg_array_41_21_real;
  assign io_coef_out_payload_0_41_21_imag = int_reg_array_41_21_imag;
  assign io_coef_out_payload_0_41_22_real = int_reg_array_41_22_real;
  assign io_coef_out_payload_0_41_22_imag = int_reg_array_41_22_imag;
  assign io_coef_out_payload_0_41_23_real = int_reg_array_41_23_real;
  assign io_coef_out_payload_0_41_23_imag = int_reg_array_41_23_imag;
  assign io_coef_out_payload_0_41_24_real = int_reg_array_41_24_real;
  assign io_coef_out_payload_0_41_24_imag = int_reg_array_41_24_imag;
  assign io_coef_out_payload_0_41_25_real = int_reg_array_41_25_real;
  assign io_coef_out_payload_0_41_25_imag = int_reg_array_41_25_imag;
  assign io_coef_out_payload_0_41_26_real = int_reg_array_41_26_real;
  assign io_coef_out_payload_0_41_26_imag = int_reg_array_41_26_imag;
  assign io_coef_out_payload_0_41_27_real = int_reg_array_41_27_real;
  assign io_coef_out_payload_0_41_27_imag = int_reg_array_41_27_imag;
  assign io_coef_out_payload_0_41_28_real = int_reg_array_41_28_real;
  assign io_coef_out_payload_0_41_28_imag = int_reg_array_41_28_imag;
  assign io_coef_out_payload_0_41_29_real = int_reg_array_41_29_real;
  assign io_coef_out_payload_0_41_29_imag = int_reg_array_41_29_imag;
  assign io_coef_out_payload_0_41_30_real = int_reg_array_41_30_real;
  assign io_coef_out_payload_0_41_30_imag = int_reg_array_41_30_imag;
  assign io_coef_out_payload_0_41_31_real = int_reg_array_41_31_real;
  assign io_coef_out_payload_0_41_31_imag = int_reg_array_41_31_imag;
  assign io_coef_out_payload_0_41_32_real = int_reg_array_41_32_real;
  assign io_coef_out_payload_0_41_32_imag = int_reg_array_41_32_imag;
  assign io_coef_out_payload_0_41_33_real = int_reg_array_41_33_real;
  assign io_coef_out_payload_0_41_33_imag = int_reg_array_41_33_imag;
  assign io_coef_out_payload_0_41_34_real = int_reg_array_41_34_real;
  assign io_coef_out_payload_0_41_34_imag = int_reg_array_41_34_imag;
  assign io_coef_out_payload_0_41_35_real = int_reg_array_41_35_real;
  assign io_coef_out_payload_0_41_35_imag = int_reg_array_41_35_imag;
  assign io_coef_out_payload_0_41_36_real = int_reg_array_41_36_real;
  assign io_coef_out_payload_0_41_36_imag = int_reg_array_41_36_imag;
  assign io_coef_out_payload_0_41_37_real = int_reg_array_41_37_real;
  assign io_coef_out_payload_0_41_37_imag = int_reg_array_41_37_imag;
  assign io_coef_out_payload_0_41_38_real = int_reg_array_41_38_real;
  assign io_coef_out_payload_0_41_38_imag = int_reg_array_41_38_imag;
  assign io_coef_out_payload_0_41_39_real = int_reg_array_41_39_real;
  assign io_coef_out_payload_0_41_39_imag = int_reg_array_41_39_imag;
  assign io_coef_out_payload_0_41_40_real = int_reg_array_41_40_real;
  assign io_coef_out_payload_0_41_40_imag = int_reg_array_41_40_imag;
  assign io_coef_out_payload_0_41_41_real = int_reg_array_41_41_real;
  assign io_coef_out_payload_0_41_41_imag = int_reg_array_41_41_imag;
  assign io_coef_out_payload_0_41_42_real = int_reg_array_41_42_real;
  assign io_coef_out_payload_0_41_42_imag = int_reg_array_41_42_imag;
  assign io_coef_out_payload_0_41_43_real = int_reg_array_41_43_real;
  assign io_coef_out_payload_0_41_43_imag = int_reg_array_41_43_imag;
  assign io_coef_out_payload_0_41_44_real = int_reg_array_41_44_real;
  assign io_coef_out_payload_0_41_44_imag = int_reg_array_41_44_imag;
  assign io_coef_out_payload_0_41_45_real = int_reg_array_41_45_real;
  assign io_coef_out_payload_0_41_45_imag = int_reg_array_41_45_imag;
  assign io_coef_out_payload_0_41_46_real = int_reg_array_41_46_real;
  assign io_coef_out_payload_0_41_46_imag = int_reg_array_41_46_imag;
  assign io_coef_out_payload_0_41_47_real = int_reg_array_41_47_real;
  assign io_coef_out_payload_0_41_47_imag = int_reg_array_41_47_imag;
  assign io_coef_out_payload_0_41_48_real = int_reg_array_41_48_real;
  assign io_coef_out_payload_0_41_48_imag = int_reg_array_41_48_imag;
  assign io_coef_out_payload_0_41_49_real = int_reg_array_41_49_real;
  assign io_coef_out_payload_0_41_49_imag = int_reg_array_41_49_imag;
  assign io_coef_out_payload_0_42_0_real = int_reg_array_42_0_real;
  assign io_coef_out_payload_0_42_0_imag = int_reg_array_42_0_imag;
  assign io_coef_out_payload_0_42_1_real = int_reg_array_42_1_real;
  assign io_coef_out_payload_0_42_1_imag = int_reg_array_42_1_imag;
  assign io_coef_out_payload_0_42_2_real = int_reg_array_42_2_real;
  assign io_coef_out_payload_0_42_2_imag = int_reg_array_42_2_imag;
  assign io_coef_out_payload_0_42_3_real = int_reg_array_42_3_real;
  assign io_coef_out_payload_0_42_3_imag = int_reg_array_42_3_imag;
  assign io_coef_out_payload_0_42_4_real = int_reg_array_42_4_real;
  assign io_coef_out_payload_0_42_4_imag = int_reg_array_42_4_imag;
  assign io_coef_out_payload_0_42_5_real = int_reg_array_42_5_real;
  assign io_coef_out_payload_0_42_5_imag = int_reg_array_42_5_imag;
  assign io_coef_out_payload_0_42_6_real = int_reg_array_42_6_real;
  assign io_coef_out_payload_0_42_6_imag = int_reg_array_42_6_imag;
  assign io_coef_out_payload_0_42_7_real = int_reg_array_42_7_real;
  assign io_coef_out_payload_0_42_7_imag = int_reg_array_42_7_imag;
  assign io_coef_out_payload_0_42_8_real = int_reg_array_42_8_real;
  assign io_coef_out_payload_0_42_8_imag = int_reg_array_42_8_imag;
  assign io_coef_out_payload_0_42_9_real = int_reg_array_42_9_real;
  assign io_coef_out_payload_0_42_9_imag = int_reg_array_42_9_imag;
  assign io_coef_out_payload_0_42_10_real = int_reg_array_42_10_real;
  assign io_coef_out_payload_0_42_10_imag = int_reg_array_42_10_imag;
  assign io_coef_out_payload_0_42_11_real = int_reg_array_42_11_real;
  assign io_coef_out_payload_0_42_11_imag = int_reg_array_42_11_imag;
  assign io_coef_out_payload_0_42_12_real = int_reg_array_42_12_real;
  assign io_coef_out_payload_0_42_12_imag = int_reg_array_42_12_imag;
  assign io_coef_out_payload_0_42_13_real = int_reg_array_42_13_real;
  assign io_coef_out_payload_0_42_13_imag = int_reg_array_42_13_imag;
  assign io_coef_out_payload_0_42_14_real = int_reg_array_42_14_real;
  assign io_coef_out_payload_0_42_14_imag = int_reg_array_42_14_imag;
  assign io_coef_out_payload_0_42_15_real = int_reg_array_42_15_real;
  assign io_coef_out_payload_0_42_15_imag = int_reg_array_42_15_imag;
  assign io_coef_out_payload_0_42_16_real = int_reg_array_42_16_real;
  assign io_coef_out_payload_0_42_16_imag = int_reg_array_42_16_imag;
  assign io_coef_out_payload_0_42_17_real = int_reg_array_42_17_real;
  assign io_coef_out_payload_0_42_17_imag = int_reg_array_42_17_imag;
  assign io_coef_out_payload_0_42_18_real = int_reg_array_42_18_real;
  assign io_coef_out_payload_0_42_18_imag = int_reg_array_42_18_imag;
  assign io_coef_out_payload_0_42_19_real = int_reg_array_42_19_real;
  assign io_coef_out_payload_0_42_19_imag = int_reg_array_42_19_imag;
  assign io_coef_out_payload_0_42_20_real = int_reg_array_42_20_real;
  assign io_coef_out_payload_0_42_20_imag = int_reg_array_42_20_imag;
  assign io_coef_out_payload_0_42_21_real = int_reg_array_42_21_real;
  assign io_coef_out_payload_0_42_21_imag = int_reg_array_42_21_imag;
  assign io_coef_out_payload_0_42_22_real = int_reg_array_42_22_real;
  assign io_coef_out_payload_0_42_22_imag = int_reg_array_42_22_imag;
  assign io_coef_out_payload_0_42_23_real = int_reg_array_42_23_real;
  assign io_coef_out_payload_0_42_23_imag = int_reg_array_42_23_imag;
  assign io_coef_out_payload_0_42_24_real = int_reg_array_42_24_real;
  assign io_coef_out_payload_0_42_24_imag = int_reg_array_42_24_imag;
  assign io_coef_out_payload_0_42_25_real = int_reg_array_42_25_real;
  assign io_coef_out_payload_0_42_25_imag = int_reg_array_42_25_imag;
  assign io_coef_out_payload_0_42_26_real = int_reg_array_42_26_real;
  assign io_coef_out_payload_0_42_26_imag = int_reg_array_42_26_imag;
  assign io_coef_out_payload_0_42_27_real = int_reg_array_42_27_real;
  assign io_coef_out_payload_0_42_27_imag = int_reg_array_42_27_imag;
  assign io_coef_out_payload_0_42_28_real = int_reg_array_42_28_real;
  assign io_coef_out_payload_0_42_28_imag = int_reg_array_42_28_imag;
  assign io_coef_out_payload_0_42_29_real = int_reg_array_42_29_real;
  assign io_coef_out_payload_0_42_29_imag = int_reg_array_42_29_imag;
  assign io_coef_out_payload_0_42_30_real = int_reg_array_42_30_real;
  assign io_coef_out_payload_0_42_30_imag = int_reg_array_42_30_imag;
  assign io_coef_out_payload_0_42_31_real = int_reg_array_42_31_real;
  assign io_coef_out_payload_0_42_31_imag = int_reg_array_42_31_imag;
  assign io_coef_out_payload_0_42_32_real = int_reg_array_42_32_real;
  assign io_coef_out_payload_0_42_32_imag = int_reg_array_42_32_imag;
  assign io_coef_out_payload_0_42_33_real = int_reg_array_42_33_real;
  assign io_coef_out_payload_0_42_33_imag = int_reg_array_42_33_imag;
  assign io_coef_out_payload_0_42_34_real = int_reg_array_42_34_real;
  assign io_coef_out_payload_0_42_34_imag = int_reg_array_42_34_imag;
  assign io_coef_out_payload_0_42_35_real = int_reg_array_42_35_real;
  assign io_coef_out_payload_0_42_35_imag = int_reg_array_42_35_imag;
  assign io_coef_out_payload_0_42_36_real = int_reg_array_42_36_real;
  assign io_coef_out_payload_0_42_36_imag = int_reg_array_42_36_imag;
  assign io_coef_out_payload_0_42_37_real = int_reg_array_42_37_real;
  assign io_coef_out_payload_0_42_37_imag = int_reg_array_42_37_imag;
  assign io_coef_out_payload_0_42_38_real = int_reg_array_42_38_real;
  assign io_coef_out_payload_0_42_38_imag = int_reg_array_42_38_imag;
  assign io_coef_out_payload_0_42_39_real = int_reg_array_42_39_real;
  assign io_coef_out_payload_0_42_39_imag = int_reg_array_42_39_imag;
  assign io_coef_out_payload_0_42_40_real = int_reg_array_42_40_real;
  assign io_coef_out_payload_0_42_40_imag = int_reg_array_42_40_imag;
  assign io_coef_out_payload_0_42_41_real = int_reg_array_42_41_real;
  assign io_coef_out_payload_0_42_41_imag = int_reg_array_42_41_imag;
  assign io_coef_out_payload_0_42_42_real = int_reg_array_42_42_real;
  assign io_coef_out_payload_0_42_42_imag = int_reg_array_42_42_imag;
  assign io_coef_out_payload_0_42_43_real = int_reg_array_42_43_real;
  assign io_coef_out_payload_0_42_43_imag = int_reg_array_42_43_imag;
  assign io_coef_out_payload_0_42_44_real = int_reg_array_42_44_real;
  assign io_coef_out_payload_0_42_44_imag = int_reg_array_42_44_imag;
  assign io_coef_out_payload_0_42_45_real = int_reg_array_42_45_real;
  assign io_coef_out_payload_0_42_45_imag = int_reg_array_42_45_imag;
  assign io_coef_out_payload_0_42_46_real = int_reg_array_42_46_real;
  assign io_coef_out_payload_0_42_46_imag = int_reg_array_42_46_imag;
  assign io_coef_out_payload_0_42_47_real = int_reg_array_42_47_real;
  assign io_coef_out_payload_0_42_47_imag = int_reg_array_42_47_imag;
  assign io_coef_out_payload_0_42_48_real = int_reg_array_42_48_real;
  assign io_coef_out_payload_0_42_48_imag = int_reg_array_42_48_imag;
  assign io_coef_out_payload_0_42_49_real = int_reg_array_42_49_real;
  assign io_coef_out_payload_0_42_49_imag = int_reg_array_42_49_imag;
  assign io_coef_out_payload_0_43_0_real = int_reg_array_43_0_real;
  assign io_coef_out_payload_0_43_0_imag = int_reg_array_43_0_imag;
  assign io_coef_out_payload_0_43_1_real = int_reg_array_43_1_real;
  assign io_coef_out_payload_0_43_1_imag = int_reg_array_43_1_imag;
  assign io_coef_out_payload_0_43_2_real = int_reg_array_43_2_real;
  assign io_coef_out_payload_0_43_2_imag = int_reg_array_43_2_imag;
  assign io_coef_out_payload_0_43_3_real = int_reg_array_43_3_real;
  assign io_coef_out_payload_0_43_3_imag = int_reg_array_43_3_imag;
  assign io_coef_out_payload_0_43_4_real = int_reg_array_43_4_real;
  assign io_coef_out_payload_0_43_4_imag = int_reg_array_43_4_imag;
  assign io_coef_out_payload_0_43_5_real = int_reg_array_43_5_real;
  assign io_coef_out_payload_0_43_5_imag = int_reg_array_43_5_imag;
  assign io_coef_out_payload_0_43_6_real = int_reg_array_43_6_real;
  assign io_coef_out_payload_0_43_6_imag = int_reg_array_43_6_imag;
  assign io_coef_out_payload_0_43_7_real = int_reg_array_43_7_real;
  assign io_coef_out_payload_0_43_7_imag = int_reg_array_43_7_imag;
  assign io_coef_out_payload_0_43_8_real = int_reg_array_43_8_real;
  assign io_coef_out_payload_0_43_8_imag = int_reg_array_43_8_imag;
  assign io_coef_out_payload_0_43_9_real = int_reg_array_43_9_real;
  assign io_coef_out_payload_0_43_9_imag = int_reg_array_43_9_imag;
  assign io_coef_out_payload_0_43_10_real = int_reg_array_43_10_real;
  assign io_coef_out_payload_0_43_10_imag = int_reg_array_43_10_imag;
  assign io_coef_out_payload_0_43_11_real = int_reg_array_43_11_real;
  assign io_coef_out_payload_0_43_11_imag = int_reg_array_43_11_imag;
  assign io_coef_out_payload_0_43_12_real = int_reg_array_43_12_real;
  assign io_coef_out_payload_0_43_12_imag = int_reg_array_43_12_imag;
  assign io_coef_out_payload_0_43_13_real = int_reg_array_43_13_real;
  assign io_coef_out_payload_0_43_13_imag = int_reg_array_43_13_imag;
  assign io_coef_out_payload_0_43_14_real = int_reg_array_43_14_real;
  assign io_coef_out_payload_0_43_14_imag = int_reg_array_43_14_imag;
  assign io_coef_out_payload_0_43_15_real = int_reg_array_43_15_real;
  assign io_coef_out_payload_0_43_15_imag = int_reg_array_43_15_imag;
  assign io_coef_out_payload_0_43_16_real = int_reg_array_43_16_real;
  assign io_coef_out_payload_0_43_16_imag = int_reg_array_43_16_imag;
  assign io_coef_out_payload_0_43_17_real = int_reg_array_43_17_real;
  assign io_coef_out_payload_0_43_17_imag = int_reg_array_43_17_imag;
  assign io_coef_out_payload_0_43_18_real = int_reg_array_43_18_real;
  assign io_coef_out_payload_0_43_18_imag = int_reg_array_43_18_imag;
  assign io_coef_out_payload_0_43_19_real = int_reg_array_43_19_real;
  assign io_coef_out_payload_0_43_19_imag = int_reg_array_43_19_imag;
  assign io_coef_out_payload_0_43_20_real = int_reg_array_43_20_real;
  assign io_coef_out_payload_0_43_20_imag = int_reg_array_43_20_imag;
  assign io_coef_out_payload_0_43_21_real = int_reg_array_43_21_real;
  assign io_coef_out_payload_0_43_21_imag = int_reg_array_43_21_imag;
  assign io_coef_out_payload_0_43_22_real = int_reg_array_43_22_real;
  assign io_coef_out_payload_0_43_22_imag = int_reg_array_43_22_imag;
  assign io_coef_out_payload_0_43_23_real = int_reg_array_43_23_real;
  assign io_coef_out_payload_0_43_23_imag = int_reg_array_43_23_imag;
  assign io_coef_out_payload_0_43_24_real = int_reg_array_43_24_real;
  assign io_coef_out_payload_0_43_24_imag = int_reg_array_43_24_imag;
  assign io_coef_out_payload_0_43_25_real = int_reg_array_43_25_real;
  assign io_coef_out_payload_0_43_25_imag = int_reg_array_43_25_imag;
  assign io_coef_out_payload_0_43_26_real = int_reg_array_43_26_real;
  assign io_coef_out_payload_0_43_26_imag = int_reg_array_43_26_imag;
  assign io_coef_out_payload_0_43_27_real = int_reg_array_43_27_real;
  assign io_coef_out_payload_0_43_27_imag = int_reg_array_43_27_imag;
  assign io_coef_out_payload_0_43_28_real = int_reg_array_43_28_real;
  assign io_coef_out_payload_0_43_28_imag = int_reg_array_43_28_imag;
  assign io_coef_out_payload_0_43_29_real = int_reg_array_43_29_real;
  assign io_coef_out_payload_0_43_29_imag = int_reg_array_43_29_imag;
  assign io_coef_out_payload_0_43_30_real = int_reg_array_43_30_real;
  assign io_coef_out_payload_0_43_30_imag = int_reg_array_43_30_imag;
  assign io_coef_out_payload_0_43_31_real = int_reg_array_43_31_real;
  assign io_coef_out_payload_0_43_31_imag = int_reg_array_43_31_imag;
  assign io_coef_out_payload_0_43_32_real = int_reg_array_43_32_real;
  assign io_coef_out_payload_0_43_32_imag = int_reg_array_43_32_imag;
  assign io_coef_out_payload_0_43_33_real = int_reg_array_43_33_real;
  assign io_coef_out_payload_0_43_33_imag = int_reg_array_43_33_imag;
  assign io_coef_out_payload_0_43_34_real = int_reg_array_43_34_real;
  assign io_coef_out_payload_0_43_34_imag = int_reg_array_43_34_imag;
  assign io_coef_out_payload_0_43_35_real = int_reg_array_43_35_real;
  assign io_coef_out_payload_0_43_35_imag = int_reg_array_43_35_imag;
  assign io_coef_out_payload_0_43_36_real = int_reg_array_43_36_real;
  assign io_coef_out_payload_0_43_36_imag = int_reg_array_43_36_imag;
  assign io_coef_out_payload_0_43_37_real = int_reg_array_43_37_real;
  assign io_coef_out_payload_0_43_37_imag = int_reg_array_43_37_imag;
  assign io_coef_out_payload_0_43_38_real = int_reg_array_43_38_real;
  assign io_coef_out_payload_0_43_38_imag = int_reg_array_43_38_imag;
  assign io_coef_out_payload_0_43_39_real = int_reg_array_43_39_real;
  assign io_coef_out_payload_0_43_39_imag = int_reg_array_43_39_imag;
  assign io_coef_out_payload_0_43_40_real = int_reg_array_43_40_real;
  assign io_coef_out_payload_0_43_40_imag = int_reg_array_43_40_imag;
  assign io_coef_out_payload_0_43_41_real = int_reg_array_43_41_real;
  assign io_coef_out_payload_0_43_41_imag = int_reg_array_43_41_imag;
  assign io_coef_out_payload_0_43_42_real = int_reg_array_43_42_real;
  assign io_coef_out_payload_0_43_42_imag = int_reg_array_43_42_imag;
  assign io_coef_out_payload_0_43_43_real = int_reg_array_43_43_real;
  assign io_coef_out_payload_0_43_43_imag = int_reg_array_43_43_imag;
  assign io_coef_out_payload_0_43_44_real = int_reg_array_43_44_real;
  assign io_coef_out_payload_0_43_44_imag = int_reg_array_43_44_imag;
  assign io_coef_out_payload_0_43_45_real = int_reg_array_43_45_real;
  assign io_coef_out_payload_0_43_45_imag = int_reg_array_43_45_imag;
  assign io_coef_out_payload_0_43_46_real = int_reg_array_43_46_real;
  assign io_coef_out_payload_0_43_46_imag = int_reg_array_43_46_imag;
  assign io_coef_out_payload_0_43_47_real = int_reg_array_43_47_real;
  assign io_coef_out_payload_0_43_47_imag = int_reg_array_43_47_imag;
  assign io_coef_out_payload_0_43_48_real = int_reg_array_43_48_real;
  assign io_coef_out_payload_0_43_48_imag = int_reg_array_43_48_imag;
  assign io_coef_out_payload_0_43_49_real = int_reg_array_43_49_real;
  assign io_coef_out_payload_0_43_49_imag = int_reg_array_43_49_imag;
  assign io_coef_out_payload_0_44_0_real = int_reg_array_44_0_real;
  assign io_coef_out_payload_0_44_0_imag = int_reg_array_44_0_imag;
  assign io_coef_out_payload_0_44_1_real = int_reg_array_44_1_real;
  assign io_coef_out_payload_0_44_1_imag = int_reg_array_44_1_imag;
  assign io_coef_out_payload_0_44_2_real = int_reg_array_44_2_real;
  assign io_coef_out_payload_0_44_2_imag = int_reg_array_44_2_imag;
  assign io_coef_out_payload_0_44_3_real = int_reg_array_44_3_real;
  assign io_coef_out_payload_0_44_3_imag = int_reg_array_44_3_imag;
  assign io_coef_out_payload_0_44_4_real = int_reg_array_44_4_real;
  assign io_coef_out_payload_0_44_4_imag = int_reg_array_44_4_imag;
  assign io_coef_out_payload_0_44_5_real = int_reg_array_44_5_real;
  assign io_coef_out_payload_0_44_5_imag = int_reg_array_44_5_imag;
  assign io_coef_out_payload_0_44_6_real = int_reg_array_44_6_real;
  assign io_coef_out_payload_0_44_6_imag = int_reg_array_44_6_imag;
  assign io_coef_out_payload_0_44_7_real = int_reg_array_44_7_real;
  assign io_coef_out_payload_0_44_7_imag = int_reg_array_44_7_imag;
  assign io_coef_out_payload_0_44_8_real = int_reg_array_44_8_real;
  assign io_coef_out_payload_0_44_8_imag = int_reg_array_44_8_imag;
  assign io_coef_out_payload_0_44_9_real = int_reg_array_44_9_real;
  assign io_coef_out_payload_0_44_9_imag = int_reg_array_44_9_imag;
  assign io_coef_out_payload_0_44_10_real = int_reg_array_44_10_real;
  assign io_coef_out_payload_0_44_10_imag = int_reg_array_44_10_imag;
  assign io_coef_out_payload_0_44_11_real = int_reg_array_44_11_real;
  assign io_coef_out_payload_0_44_11_imag = int_reg_array_44_11_imag;
  assign io_coef_out_payload_0_44_12_real = int_reg_array_44_12_real;
  assign io_coef_out_payload_0_44_12_imag = int_reg_array_44_12_imag;
  assign io_coef_out_payload_0_44_13_real = int_reg_array_44_13_real;
  assign io_coef_out_payload_0_44_13_imag = int_reg_array_44_13_imag;
  assign io_coef_out_payload_0_44_14_real = int_reg_array_44_14_real;
  assign io_coef_out_payload_0_44_14_imag = int_reg_array_44_14_imag;
  assign io_coef_out_payload_0_44_15_real = int_reg_array_44_15_real;
  assign io_coef_out_payload_0_44_15_imag = int_reg_array_44_15_imag;
  assign io_coef_out_payload_0_44_16_real = int_reg_array_44_16_real;
  assign io_coef_out_payload_0_44_16_imag = int_reg_array_44_16_imag;
  assign io_coef_out_payload_0_44_17_real = int_reg_array_44_17_real;
  assign io_coef_out_payload_0_44_17_imag = int_reg_array_44_17_imag;
  assign io_coef_out_payload_0_44_18_real = int_reg_array_44_18_real;
  assign io_coef_out_payload_0_44_18_imag = int_reg_array_44_18_imag;
  assign io_coef_out_payload_0_44_19_real = int_reg_array_44_19_real;
  assign io_coef_out_payload_0_44_19_imag = int_reg_array_44_19_imag;
  assign io_coef_out_payload_0_44_20_real = int_reg_array_44_20_real;
  assign io_coef_out_payload_0_44_20_imag = int_reg_array_44_20_imag;
  assign io_coef_out_payload_0_44_21_real = int_reg_array_44_21_real;
  assign io_coef_out_payload_0_44_21_imag = int_reg_array_44_21_imag;
  assign io_coef_out_payload_0_44_22_real = int_reg_array_44_22_real;
  assign io_coef_out_payload_0_44_22_imag = int_reg_array_44_22_imag;
  assign io_coef_out_payload_0_44_23_real = int_reg_array_44_23_real;
  assign io_coef_out_payload_0_44_23_imag = int_reg_array_44_23_imag;
  assign io_coef_out_payload_0_44_24_real = int_reg_array_44_24_real;
  assign io_coef_out_payload_0_44_24_imag = int_reg_array_44_24_imag;
  assign io_coef_out_payload_0_44_25_real = int_reg_array_44_25_real;
  assign io_coef_out_payload_0_44_25_imag = int_reg_array_44_25_imag;
  assign io_coef_out_payload_0_44_26_real = int_reg_array_44_26_real;
  assign io_coef_out_payload_0_44_26_imag = int_reg_array_44_26_imag;
  assign io_coef_out_payload_0_44_27_real = int_reg_array_44_27_real;
  assign io_coef_out_payload_0_44_27_imag = int_reg_array_44_27_imag;
  assign io_coef_out_payload_0_44_28_real = int_reg_array_44_28_real;
  assign io_coef_out_payload_0_44_28_imag = int_reg_array_44_28_imag;
  assign io_coef_out_payload_0_44_29_real = int_reg_array_44_29_real;
  assign io_coef_out_payload_0_44_29_imag = int_reg_array_44_29_imag;
  assign io_coef_out_payload_0_44_30_real = int_reg_array_44_30_real;
  assign io_coef_out_payload_0_44_30_imag = int_reg_array_44_30_imag;
  assign io_coef_out_payload_0_44_31_real = int_reg_array_44_31_real;
  assign io_coef_out_payload_0_44_31_imag = int_reg_array_44_31_imag;
  assign io_coef_out_payload_0_44_32_real = int_reg_array_44_32_real;
  assign io_coef_out_payload_0_44_32_imag = int_reg_array_44_32_imag;
  assign io_coef_out_payload_0_44_33_real = int_reg_array_44_33_real;
  assign io_coef_out_payload_0_44_33_imag = int_reg_array_44_33_imag;
  assign io_coef_out_payload_0_44_34_real = int_reg_array_44_34_real;
  assign io_coef_out_payload_0_44_34_imag = int_reg_array_44_34_imag;
  assign io_coef_out_payload_0_44_35_real = int_reg_array_44_35_real;
  assign io_coef_out_payload_0_44_35_imag = int_reg_array_44_35_imag;
  assign io_coef_out_payload_0_44_36_real = int_reg_array_44_36_real;
  assign io_coef_out_payload_0_44_36_imag = int_reg_array_44_36_imag;
  assign io_coef_out_payload_0_44_37_real = int_reg_array_44_37_real;
  assign io_coef_out_payload_0_44_37_imag = int_reg_array_44_37_imag;
  assign io_coef_out_payload_0_44_38_real = int_reg_array_44_38_real;
  assign io_coef_out_payload_0_44_38_imag = int_reg_array_44_38_imag;
  assign io_coef_out_payload_0_44_39_real = int_reg_array_44_39_real;
  assign io_coef_out_payload_0_44_39_imag = int_reg_array_44_39_imag;
  assign io_coef_out_payload_0_44_40_real = int_reg_array_44_40_real;
  assign io_coef_out_payload_0_44_40_imag = int_reg_array_44_40_imag;
  assign io_coef_out_payload_0_44_41_real = int_reg_array_44_41_real;
  assign io_coef_out_payload_0_44_41_imag = int_reg_array_44_41_imag;
  assign io_coef_out_payload_0_44_42_real = int_reg_array_44_42_real;
  assign io_coef_out_payload_0_44_42_imag = int_reg_array_44_42_imag;
  assign io_coef_out_payload_0_44_43_real = int_reg_array_44_43_real;
  assign io_coef_out_payload_0_44_43_imag = int_reg_array_44_43_imag;
  assign io_coef_out_payload_0_44_44_real = int_reg_array_44_44_real;
  assign io_coef_out_payload_0_44_44_imag = int_reg_array_44_44_imag;
  assign io_coef_out_payload_0_44_45_real = int_reg_array_44_45_real;
  assign io_coef_out_payload_0_44_45_imag = int_reg_array_44_45_imag;
  assign io_coef_out_payload_0_44_46_real = int_reg_array_44_46_real;
  assign io_coef_out_payload_0_44_46_imag = int_reg_array_44_46_imag;
  assign io_coef_out_payload_0_44_47_real = int_reg_array_44_47_real;
  assign io_coef_out_payload_0_44_47_imag = int_reg_array_44_47_imag;
  assign io_coef_out_payload_0_44_48_real = int_reg_array_44_48_real;
  assign io_coef_out_payload_0_44_48_imag = int_reg_array_44_48_imag;
  assign io_coef_out_payload_0_44_49_real = int_reg_array_44_49_real;
  assign io_coef_out_payload_0_44_49_imag = int_reg_array_44_49_imag;
  assign io_coef_out_payload_0_45_0_real = int_reg_array_45_0_real;
  assign io_coef_out_payload_0_45_0_imag = int_reg_array_45_0_imag;
  assign io_coef_out_payload_0_45_1_real = int_reg_array_45_1_real;
  assign io_coef_out_payload_0_45_1_imag = int_reg_array_45_1_imag;
  assign io_coef_out_payload_0_45_2_real = int_reg_array_45_2_real;
  assign io_coef_out_payload_0_45_2_imag = int_reg_array_45_2_imag;
  assign io_coef_out_payload_0_45_3_real = int_reg_array_45_3_real;
  assign io_coef_out_payload_0_45_3_imag = int_reg_array_45_3_imag;
  assign io_coef_out_payload_0_45_4_real = int_reg_array_45_4_real;
  assign io_coef_out_payload_0_45_4_imag = int_reg_array_45_4_imag;
  assign io_coef_out_payload_0_45_5_real = int_reg_array_45_5_real;
  assign io_coef_out_payload_0_45_5_imag = int_reg_array_45_5_imag;
  assign io_coef_out_payload_0_45_6_real = int_reg_array_45_6_real;
  assign io_coef_out_payload_0_45_6_imag = int_reg_array_45_6_imag;
  assign io_coef_out_payload_0_45_7_real = int_reg_array_45_7_real;
  assign io_coef_out_payload_0_45_7_imag = int_reg_array_45_7_imag;
  assign io_coef_out_payload_0_45_8_real = int_reg_array_45_8_real;
  assign io_coef_out_payload_0_45_8_imag = int_reg_array_45_8_imag;
  assign io_coef_out_payload_0_45_9_real = int_reg_array_45_9_real;
  assign io_coef_out_payload_0_45_9_imag = int_reg_array_45_9_imag;
  assign io_coef_out_payload_0_45_10_real = int_reg_array_45_10_real;
  assign io_coef_out_payload_0_45_10_imag = int_reg_array_45_10_imag;
  assign io_coef_out_payload_0_45_11_real = int_reg_array_45_11_real;
  assign io_coef_out_payload_0_45_11_imag = int_reg_array_45_11_imag;
  assign io_coef_out_payload_0_45_12_real = int_reg_array_45_12_real;
  assign io_coef_out_payload_0_45_12_imag = int_reg_array_45_12_imag;
  assign io_coef_out_payload_0_45_13_real = int_reg_array_45_13_real;
  assign io_coef_out_payload_0_45_13_imag = int_reg_array_45_13_imag;
  assign io_coef_out_payload_0_45_14_real = int_reg_array_45_14_real;
  assign io_coef_out_payload_0_45_14_imag = int_reg_array_45_14_imag;
  assign io_coef_out_payload_0_45_15_real = int_reg_array_45_15_real;
  assign io_coef_out_payload_0_45_15_imag = int_reg_array_45_15_imag;
  assign io_coef_out_payload_0_45_16_real = int_reg_array_45_16_real;
  assign io_coef_out_payload_0_45_16_imag = int_reg_array_45_16_imag;
  assign io_coef_out_payload_0_45_17_real = int_reg_array_45_17_real;
  assign io_coef_out_payload_0_45_17_imag = int_reg_array_45_17_imag;
  assign io_coef_out_payload_0_45_18_real = int_reg_array_45_18_real;
  assign io_coef_out_payload_0_45_18_imag = int_reg_array_45_18_imag;
  assign io_coef_out_payload_0_45_19_real = int_reg_array_45_19_real;
  assign io_coef_out_payload_0_45_19_imag = int_reg_array_45_19_imag;
  assign io_coef_out_payload_0_45_20_real = int_reg_array_45_20_real;
  assign io_coef_out_payload_0_45_20_imag = int_reg_array_45_20_imag;
  assign io_coef_out_payload_0_45_21_real = int_reg_array_45_21_real;
  assign io_coef_out_payload_0_45_21_imag = int_reg_array_45_21_imag;
  assign io_coef_out_payload_0_45_22_real = int_reg_array_45_22_real;
  assign io_coef_out_payload_0_45_22_imag = int_reg_array_45_22_imag;
  assign io_coef_out_payload_0_45_23_real = int_reg_array_45_23_real;
  assign io_coef_out_payload_0_45_23_imag = int_reg_array_45_23_imag;
  assign io_coef_out_payload_0_45_24_real = int_reg_array_45_24_real;
  assign io_coef_out_payload_0_45_24_imag = int_reg_array_45_24_imag;
  assign io_coef_out_payload_0_45_25_real = int_reg_array_45_25_real;
  assign io_coef_out_payload_0_45_25_imag = int_reg_array_45_25_imag;
  assign io_coef_out_payload_0_45_26_real = int_reg_array_45_26_real;
  assign io_coef_out_payload_0_45_26_imag = int_reg_array_45_26_imag;
  assign io_coef_out_payload_0_45_27_real = int_reg_array_45_27_real;
  assign io_coef_out_payload_0_45_27_imag = int_reg_array_45_27_imag;
  assign io_coef_out_payload_0_45_28_real = int_reg_array_45_28_real;
  assign io_coef_out_payload_0_45_28_imag = int_reg_array_45_28_imag;
  assign io_coef_out_payload_0_45_29_real = int_reg_array_45_29_real;
  assign io_coef_out_payload_0_45_29_imag = int_reg_array_45_29_imag;
  assign io_coef_out_payload_0_45_30_real = int_reg_array_45_30_real;
  assign io_coef_out_payload_0_45_30_imag = int_reg_array_45_30_imag;
  assign io_coef_out_payload_0_45_31_real = int_reg_array_45_31_real;
  assign io_coef_out_payload_0_45_31_imag = int_reg_array_45_31_imag;
  assign io_coef_out_payload_0_45_32_real = int_reg_array_45_32_real;
  assign io_coef_out_payload_0_45_32_imag = int_reg_array_45_32_imag;
  assign io_coef_out_payload_0_45_33_real = int_reg_array_45_33_real;
  assign io_coef_out_payload_0_45_33_imag = int_reg_array_45_33_imag;
  assign io_coef_out_payload_0_45_34_real = int_reg_array_45_34_real;
  assign io_coef_out_payload_0_45_34_imag = int_reg_array_45_34_imag;
  assign io_coef_out_payload_0_45_35_real = int_reg_array_45_35_real;
  assign io_coef_out_payload_0_45_35_imag = int_reg_array_45_35_imag;
  assign io_coef_out_payload_0_45_36_real = int_reg_array_45_36_real;
  assign io_coef_out_payload_0_45_36_imag = int_reg_array_45_36_imag;
  assign io_coef_out_payload_0_45_37_real = int_reg_array_45_37_real;
  assign io_coef_out_payload_0_45_37_imag = int_reg_array_45_37_imag;
  assign io_coef_out_payload_0_45_38_real = int_reg_array_45_38_real;
  assign io_coef_out_payload_0_45_38_imag = int_reg_array_45_38_imag;
  assign io_coef_out_payload_0_45_39_real = int_reg_array_45_39_real;
  assign io_coef_out_payload_0_45_39_imag = int_reg_array_45_39_imag;
  assign io_coef_out_payload_0_45_40_real = int_reg_array_45_40_real;
  assign io_coef_out_payload_0_45_40_imag = int_reg_array_45_40_imag;
  assign io_coef_out_payload_0_45_41_real = int_reg_array_45_41_real;
  assign io_coef_out_payload_0_45_41_imag = int_reg_array_45_41_imag;
  assign io_coef_out_payload_0_45_42_real = int_reg_array_45_42_real;
  assign io_coef_out_payload_0_45_42_imag = int_reg_array_45_42_imag;
  assign io_coef_out_payload_0_45_43_real = int_reg_array_45_43_real;
  assign io_coef_out_payload_0_45_43_imag = int_reg_array_45_43_imag;
  assign io_coef_out_payload_0_45_44_real = int_reg_array_45_44_real;
  assign io_coef_out_payload_0_45_44_imag = int_reg_array_45_44_imag;
  assign io_coef_out_payload_0_45_45_real = int_reg_array_45_45_real;
  assign io_coef_out_payload_0_45_45_imag = int_reg_array_45_45_imag;
  assign io_coef_out_payload_0_45_46_real = int_reg_array_45_46_real;
  assign io_coef_out_payload_0_45_46_imag = int_reg_array_45_46_imag;
  assign io_coef_out_payload_0_45_47_real = int_reg_array_45_47_real;
  assign io_coef_out_payload_0_45_47_imag = int_reg_array_45_47_imag;
  assign io_coef_out_payload_0_45_48_real = int_reg_array_45_48_real;
  assign io_coef_out_payload_0_45_48_imag = int_reg_array_45_48_imag;
  assign io_coef_out_payload_0_45_49_real = int_reg_array_45_49_real;
  assign io_coef_out_payload_0_45_49_imag = int_reg_array_45_49_imag;
  assign io_coef_out_payload_0_46_0_real = int_reg_array_46_0_real;
  assign io_coef_out_payload_0_46_0_imag = int_reg_array_46_0_imag;
  assign io_coef_out_payload_0_46_1_real = int_reg_array_46_1_real;
  assign io_coef_out_payload_0_46_1_imag = int_reg_array_46_1_imag;
  assign io_coef_out_payload_0_46_2_real = int_reg_array_46_2_real;
  assign io_coef_out_payload_0_46_2_imag = int_reg_array_46_2_imag;
  assign io_coef_out_payload_0_46_3_real = int_reg_array_46_3_real;
  assign io_coef_out_payload_0_46_3_imag = int_reg_array_46_3_imag;
  assign io_coef_out_payload_0_46_4_real = int_reg_array_46_4_real;
  assign io_coef_out_payload_0_46_4_imag = int_reg_array_46_4_imag;
  assign io_coef_out_payload_0_46_5_real = int_reg_array_46_5_real;
  assign io_coef_out_payload_0_46_5_imag = int_reg_array_46_5_imag;
  assign io_coef_out_payload_0_46_6_real = int_reg_array_46_6_real;
  assign io_coef_out_payload_0_46_6_imag = int_reg_array_46_6_imag;
  assign io_coef_out_payload_0_46_7_real = int_reg_array_46_7_real;
  assign io_coef_out_payload_0_46_7_imag = int_reg_array_46_7_imag;
  assign io_coef_out_payload_0_46_8_real = int_reg_array_46_8_real;
  assign io_coef_out_payload_0_46_8_imag = int_reg_array_46_8_imag;
  assign io_coef_out_payload_0_46_9_real = int_reg_array_46_9_real;
  assign io_coef_out_payload_0_46_9_imag = int_reg_array_46_9_imag;
  assign io_coef_out_payload_0_46_10_real = int_reg_array_46_10_real;
  assign io_coef_out_payload_0_46_10_imag = int_reg_array_46_10_imag;
  assign io_coef_out_payload_0_46_11_real = int_reg_array_46_11_real;
  assign io_coef_out_payload_0_46_11_imag = int_reg_array_46_11_imag;
  assign io_coef_out_payload_0_46_12_real = int_reg_array_46_12_real;
  assign io_coef_out_payload_0_46_12_imag = int_reg_array_46_12_imag;
  assign io_coef_out_payload_0_46_13_real = int_reg_array_46_13_real;
  assign io_coef_out_payload_0_46_13_imag = int_reg_array_46_13_imag;
  assign io_coef_out_payload_0_46_14_real = int_reg_array_46_14_real;
  assign io_coef_out_payload_0_46_14_imag = int_reg_array_46_14_imag;
  assign io_coef_out_payload_0_46_15_real = int_reg_array_46_15_real;
  assign io_coef_out_payload_0_46_15_imag = int_reg_array_46_15_imag;
  assign io_coef_out_payload_0_46_16_real = int_reg_array_46_16_real;
  assign io_coef_out_payload_0_46_16_imag = int_reg_array_46_16_imag;
  assign io_coef_out_payload_0_46_17_real = int_reg_array_46_17_real;
  assign io_coef_out_payload_0_46_17_imag = int_reg_array_46_17_imag;
  assign io_coef_out_payload_0_46_18_real = int_reg_array_46_18_real;
  assign io_coef_out_payload_0_46_18_imag = int_reg_array_46_18_imag;
  assign io_coef_out_payload_0_46_19_real = int_reg_array_46_19_real;
  assign io_coef_out_payload_0_46_19_imag = int_reg_array_46_19_imag;
  assign io_coef_out_payload_0_46_20_real = int_reg_array_46_20_real;
  assign io_coef_out_payload_0_46_20_imag = int_reg_array_46_20_imag;
  assign io_coef_out_payload_0_46_21_real = int_reg_array_46_21_real;
  assign io_coef_out_payload_0_46_21_imag = int_reg_array_46_21_imag;
  assign io_coef_out_payload_0_46_22_real = int_reg_array_46_22_real;
  assign io_coef_out_payload_0_46_22_imag = int_reg_array_46_22_imag;
  assign io_coef_out_payload_0_46_23_real = int_reg_array_46_23_real;
  assign io_coef_out_payload_0_46_23_imag = int_reg_array_46_23_imag;
  assign io_coef_out_payload_0_46_24_real = int_reg_array_46_24_real;
  assign io_coef_out_payload_0_46_24_imag = int_reg_array_46_24_imag;
  assign io_coef_out_payload_0_46_25_real = int_reg_array_46_25_real;
  assign io_coef_out_payload_0_46_25_imag = int_reg_array_46_25_imag;
  assign io_coef_out_payload_0_46_26_real = int_reg_array_46_26_real;
  assign io_coef_out_payload_0_46_26_imag = int_reg_array_46_26_imag;
  assign io_coef_out_payload_0_46_27_real = int_reg_array_46_27_real;
  assign io_coef_out_payload_0_46_27_imag = int_reg_array_46_27_imag;
  assign io_coef_out_payload_0_46_28_real = int_reg_array_46_28_real;
  assign io_coef_out_payload_0_46_28_imag = int_reg_array_46_28_imag;
  assign io_coef_out_payload_0_46_29_real = int_reg_array_46_29_real;
  assign io_coef_out_payload_0_46_29_imag = int_reg_array_46_29_imag;
  assign io_coef_out_payload_0_46_30_real = int_reg_array_46_30_real;
  assign io_coef_out_payload_0_46_30_imag = int_reg_array_46_30_imag;
  assign io_coef_out_payload_0_46_31_real = int_reg_array_46_31_real;
  assign io_coef_out_payload_0_46_31_imag = int_reg_array_46_31_imag;
  assign io_coef_out_payload_0_46_32_real = int_reg_array_46_32_real;
  assign io_coef_out_payload_0_46_32_imag = int_reg_array_46_32_imag;
  assign io_coef_out_payload_0_46_33_real = int_reg_array_46_33_real;
  assign io_coef_out_payload_0_46_33_imag = int_reg_array_46_33_imag;
  assign io_coef_out_payload_0_46_34_real = int_reg_array_46_34_real;
  assign io_coef_out_payload_0_46_34_imag = int_reg_array_46_34_imag;
  assign io_coef_out_payload_0_46_35_real = int_reg_array_46_35_real;
  assign io_coef_out_payload_0_46_35_imag = int_reg_array_46_35_imag;
  assign io_coef_out_payload_0_46_36_real = int_reg_array_46_36_real;
  assign io_coef_out_payload_0_46_36_imag = int_reg_array_46_36_imag;
  assign io_coef_out_payload_0_46_37_real = int_reg_array_46_37_real;
  assign io_coef_out_payload_0_46_37_imag = int_reg_array_46_37_imag;
  assign io_coef_out_payload_0_46_38_real = int_reg_array_46_38_real;
  assign io_coef_out_payload_0_46_38_imag = int_reg_array_46_38_imag;
  assign io_coef_out_payload_0_46_39_real = int_reg_array_46_39_real;
  assign io_coef_out_payload_0_46_39_imag = int_reg_array_46_39_imag;
  assign io_coef_out_payload_0_46_40_real = int_reg_array_46_40_real;
  assign io_coef_out_payload_0_46_40_imag = int_reg_array_46_40_imag;
  assign io_coef_out_payload_0_46_41_real = int_reg_array_46_41_real;
  assign io_coef_out_payload_0_46_41_imag = int_reg_array_46_41_imag;
  assign io_coef_out_payload_0_46_42_real = int_reg_array_46_42_real;
  assign io_coef_out_payload_0_46_42_imag = int_reg_array_46_42_imag;
  assign io_coef_out_payload_0_46_43_real = int_reg_array_46_43_real;
  assign io_coef_out_payload_0_46_43_imag = int_reg_array_46_43_imag;
  assign io_coef_out_payload_0_46_44_real = int_reg_array_46_44_real;
  assign io_coef_out_payload_0_46_44_imag = int_reg_array_46_44_imag;
  assign io_coef_out_payload_0_46_45_real = int_reg_array_46_45_real;
  assign io_coef_out_payload_0_46_45_imag = int_reg_array_46_45_imag;
  assign io_coef_out_payload_0_46_46_real = int_reg_array_46_46_real;
  assign io_coef_out_payload_0_46_46_imag = int_reg_array_46_46_imag;
  assign io_coef_out_payload_0_46_47_real = int_reg_array_46_47_real;
  assign io_coef_out_payload_0_46_47_imag = int_reg_array_46_47_imag;
  assign io_coef_out_payload_0_46_48_real = int_reg_array_46_48_real;
  assign io_coef_out_payload_0_46_48_imag = int_reg_array_46_48_imag;
  assign io_coef_out_payload_0_46_49_real = int_reg_array_46_49_real;
  assign io_coef_out_payload_0_46_49_imag = int_reg_array_46_49_imag;
  assign io_coef_out_payload_0_47_0_real = int_reg_array_47_0_real;
  assign io_coef_out_payload_0_47_0_imag = int_reg_array_47_0_imag;
  assign io_coef_out_payload_0_47_1_real = int_reg_array_47_1_real;
  assign io_coef_out_payload_0_47_1_imag = int_reg_array_47_1_imag;
  assign io_coef_out_payload_0_47_2_real = int_reg_array_47_2_real;
  assign io_coef_out_payload_0_47_2_imag = int_reg_array_47_2_imag;
  assign io_coef_out_payload_0_47_3_real = int_reg_array_47_3_real;
  assign io_coef_out_payload_0_47_3_imag = int_reg_array_47_3_imag;
  assign io_coef_out_payload_0_47_4_real = int_reg_array_47_4_real;
  assign io_coef_out_payload_0_47_4_imag = int_reg_array_47_4_imag;
  assign io_coef_out_payload_0_47_5_real = int_reg_array_47_5_real;
  assign io_coef_out_payload_0_47_5_imag = int_reg_array_47_5_imag;
  assign io_coef_out_payload_0_47_6_real = int_reg_array_47_6_real;
  assign io_coef_out_payload_0_47_6_imag = int_reg_array_47_6_imag;
  assign io_coef_out_payload_0_47_7_real = int_reg_array_47_7_real;
  assign io_coef_out_payload_0_47_7_imag = int_reg_array_47_7_imag;
  assign io_coef_out_payload_0_47_8_real = int_reg_array_47_8_real;
  assign io_coef_out_payload_0_47_8_imag = int_reg_array_47_8_imag;
  assign io_coef_out_payload_0_47_9_real = int_reg_array_47_9_real;
  assign io_coef_out_payload_0_47_9_imag = int_reg_array_47_9_imag;
  assign io_coef_out_payload_0_47_10_real = int_reg_array_47_10_real;
  assign io_coef_out_payload_0_47_10_imag = int_reg_array_47_10_imag;
  assign io_coef_out_payload_0_47_11_real = int_reg_array_47_11_real;
  assign io_coef_out_payload_0_47_11_imag = int_reg_array_47_11_imag;
  assign io_coef_out_payload_0_47_12_real = int_reg_array_47_12_real;
  assign io_coef_out_payload_0_47_12_imag = int_reg_array_47_12_imag;
  assign io_coef_out_payload_0_47_13_real = int_reg_array_47_13_real;
  assign io_coef_out_payload_0_47_13_imag = int_reg_array_47_13_imag;
  assign io_coef_out_payload_0_47_14_real = int_reg_array_47_14_real;
  assign io_coef_out_payload_0_47_14_imag = int_reg_array_47_14_imag;
  assign io_coef_out_payload_0_47_15_real = int_reg_array_47_15_real;
  assign io_coef_out_payload_0_47_15_imag = int_reg_array_47_15_imag;
  assign io_coef_out_payload_0_47_16_real = int_reg_array_47_16_real;
  assign io_coef_out_payload_0_47_16_imag = int_reg_array_47_16_imag;
  assign io_coef_out_payload_0_47_17_real = int_reg_array_47_17_real;
  assign io_coef_out_payload_0_47_17_imag = int_reg_array_47_17_imag;
  assign io_coef_out_payload_0_47_18_real = int_reg_array_47_18_real;
  assign io_coef_out_payload_0_47_18_imag = int_reg_array_47_18_imag;
  assign io_coef_out_payload_0_47_19_real = int_reg_array_47_19_real;
  assign io_coef_out_payload_0_47_19_imag = int_reg_array_47_19_imag;
  assign io_coef_out_payload_0_47_20_real = int_reg_array_47_20_real;
  assign io_coef_out_payload_0_47_20_imag = int_reg_array_47_20_imag;
  assign io_coef_out_payload_0_47_21_real = int_reg_array_47_21_real;
  assign io_coef_out_payload_0_47_21_imag = int_reg_array_47_21_imag;
  assign io_coef_out_payload_0_47_22_real = int_reg_array_47_22_real;
  assign io_coef_out_payload_0_47_22_imag = int_reg_array_47_22_imag;
  assign io_coef_out_payload_0_47_23_real = int_reg_array_47_23_real;
  assign io_coef_out_payload_0_47_23_imag = int_reg_array_47_23_imag;
  assign io_coef_out_payload_0_47_24_real = int_reg_array_47_24_real;
  assign io_coef_out_payload_0_47_24_imag = int_reg_array_47_24_imag;
  assign io_coef_out_payload_0_47_25_real = int_reg_array_47_25_real;
  assign io_coef_out_payload_0_47_25_imag = int_reg_array_47_25_imag;
  assign io_coef_out_payload_0_47_26_real = int_reg_array_47_26_real;
  assign io_coef_out_payload_0_47_26_imag = int_reg_array_47_26_imag;
  assign io_coef_out_payload_0_47_27_real = int_reg_array_47_27_real;
  assign io_coef_out_payload_0_47_27_imag = int_reg_array_47_27_imag;
  assign io_coef_out_payload_0_47_28_real = int_reg_array_47_28_real;
  assign io_coef_out_payload_0_47_28_imag = int_reg_array_47_28_imag;
  assign io_coef_out_payload_0_47_29_real = int_reg_array_47_29_real;
  assign io_coef_out_payload_0_47_29_imag = int_reg_array_47_29_imag;
  assign io_coef_out_payload_0_47_30_real = int_reg_array_47_30_real;
  assign io_coef_out_payload_0_47_30_imag = int_reg_array_47_30_imag;
  assign io_coef_out_payload_0_47_31_real = int_reg_array_47_31_real;
  assign io_coef_out_payload_0_47_31_imag = int_reg_array_47_31_imag;
  assign io_coef_out_payload_0_47_32_real = int_reg_array_47_32_real;
  assign io_coef_out_payload_0_47_32_imag = int_reg_array_47_32_imag;
  assign io_coef_out_payload_0_47_33_real = int_reg_array_47_33_real;
  assign io_coef_out_payload_0_47_33_imag = int_reg_array_47_33_imag;
  assign io_coef_out_payload_0_47_34_real = int_reg_array_47_34_real;
  assign io_coef_out_payload_0_47_34_imag = int_reg_array_47_34_imag;
  assign io_coef_out_payload_0_47_35_real = int_reg_array_47_35_real;
  assign io_coef_out_payload_0_47_35_imag = int_reg_array_47_35_imag;
  assign io_coef_out_payload_0_47_36_real = int_reg_array_47_36_real;
  assign io_coef_out_payload_0_47_36_imag = int_reg_array_47_36_imag;
  assign io_coef_out_payload_0_47_37_real = int_reg_array_47_37_real;
  assign io_coef_out_payload_0_47_37_imag = int_reg_array_47_37_imag;
  assign io_coef_out_payload_0_47_38_real = int_reg_array_47_38_real;
  assign io_coef_out_payload_0_47_38_imag = int_reg_array_47_38_imag;
  assign io_coef_out_payload_0_47_39_real = int_reg_array_47_39_real;
  assign io_coef_out_payload_0_47_39_imag = int_reg_array_47_39_imag;
  assign io_coef_out_payload_0_47_40_real = int_reg_array_47_40_real;
  assign io_coef_out_payload_0_47_40_imag = int_reg_array_47_40_imag;
  assign io_coef_out_payload_0_47_41_real = int_reg_array_47_41_real;
  assign io_coef_out_payload_0_47_41_imag = int_reg_array_47_41_imag;
  assign io_coef_out_payload_0_47_42_real = int_reg_array_47_42_real;
  assign io_coef_out_payload_0_47_42_imag = int_reg_array_47_42_imag;
  assign io_coef_out_payload_0_47_43_real = int_reg_array_47_43_real;
  assign io_coef_out_payload_0_47_43_imag = int_reg_array_47_43_imag;
  assign io_coef_out_payload_0_47_44_real = int_reg_array_47_44_real;
  assign io_coef_out_payload_0_47_44_imag = int_reg_array_47_44_imag;
  assign io_coef_out_payload_0_47_45_real = int_reg_array_47_45_real;
  assign io_coef_out_payload_0_47_45_imag = int_reg_array_47_45_imag;
  assign io_coef_out_payload_0_47_46_real = int_reg_array_47_46_real;
  assign io_coef_out_payload_0_47_46_imag = int_reg_array_47_46_imag;
  assign io_coef_out_payload_0_47_47_real = int_reg_array_47_47_real;
  assign io_coef_out_payload_0_47_47_imag = int_reg_array_47_47_imag;
  assign io_coef_out_payload_0_47_48_real = int_reg_array_47_48_real;
  assign io_coef_out_payload_0_47_48_imag = int_reg_array_47_48_imag;
  assign io_coef_out_payload_0_47_49_real = int_reg_array_47_49_real;
  assign io_coef_out_payload_0_47_49_imag = int_reg_array_47_49_imag;
  assign io_coef_out_payload_0_48_0_real = int_reg_array_48_0_real;
  assign io_coef_out_payload_0_48_0_imag = int_reg_array_48_0_imag;
  assign io_coef_out_payload_0_48_1_real = int_reg_array_48_1_real;
  assign io_coef_out_payload_0_48_1_imag = int_reg_array_48_1_imag;
  assign io_coef_out_payload_0_48_2_real = int_reg_array_48_2_real;
  assign io_coef_out_payload_0_48_2_imag = int_reg_array_48_2_imag;
  assign io_coef_out_payload_0_48_3_real = int_reg_array_48_3_real;
  assign io_coef_out_payload_0_48_3_imag = int_reg_array_48_3_imag;
  assign io_coef_out_payload_0_48_4_real = int_reg_array_48_4_real;
  assign io_coef_out_payload_0_48_4_imag = int_reg_array_48_4_imag;
  assign io_coef_out_payload_0_48_5_real = int_reg_array_48_5_real;
  assign io_coef_out_payload_0_48_5_imag = int_reg_array_48_5_imag;
  assign io_coef_out_payload_0_48_6_real = int_reg_array_48_6_real;
  assign io_coef_out_payload_0_48_6_imag = int_reg_array_48_6_imag;
  assign io_coef_out_payload_0_48_7_real = int_reg_array_48_7_real;
  assign io_coef_out_payload_0_48_7_imag = int_reg_array_48_7_imag;
  assign io_coef_out_payload_0_48_8_real = int_reg_array_48_8_real;
  assign io_coef_out_payload_0_48_8_imag = int_reg_array_48_8_imag;
  assign io_coef_out_payload_0_48_9_real = int_reg_array_48_9_real;
  assign io_coef_out_payload_0_48_9_imag = int_reg_array_48_9_imag;
  assign io_coef_out_payload_0_48_10_real = int_reg_array_48_10_real;
  assign io_coef_out_payload_0_48_10_imag = int_reg_array_48_10_imag;
  assign io_coef_out_payload_0_48_11_real = int_reg_array_48_11_real;
  assign io_coef_out_payload_0_48_11_imag = int_reg_array_48_11_imag;
  assign io_coef_out_payload_0_48_12_real = int_reg_array_48_12_real;
  assign io_coef_out_payload_0_48_12_imag = int_reg_array_48_12_imag;
  assign io_coef_out_payload_0_48_13_real = int_reg_array_48_13_real;
  assign io_coef_out_payload_0_48_13_imag = int_reg_array_48_13_imag;
  assign io_coef_out_payload_0_48_14_real = int_reg_array_48_14_real;
  assign io_coef_out_payload_0_48_14_imag = int_reg_array_48_14_imag;
  assign io_coef_out_payload_0_48_15_real = int_reg_array_48_15_real;
  assign io_coef_out_payload_0_48_15_imag = int_reg_array_48_15_imag;
  assign io_coef_out_payload_0_48_16_real = int_reg_array_48_16_real;
  assign io_coef_out_payload_0_48_16_imag = int_reg_array_48_16_imag;
  assign io_coef_out_payload_0_48_17_real = int_reg_array_48_17_real;
  assign io_coef_out_payload_0_48_17_imag = int_reg_array_48_17_imag;
  assign io_coef_out_payload_0_48_18_real = int_reg_array_48_18_real;
  assign io_coef_out_payload_0_48_18_imag = int_reg_array_48_18_imag;
  assign io_coef_out_payload_0_48_19_real = int_reg_array_48_19_real;
  assign io_coef_out_payload_0_48_19_imag = int_reg_array_48_19_imag;
  assign io_coef_out_payload_0_48_20_real = int_reg_array_48_20_real;
  assign io_coef_out_payload_0_48_20_imag = int_reg_array_48_20_imag;
  assign io_coef_out_payload_0_48_21_real = int_reg_array_48_21_real;
  assign io_coef_out_payload_0_48_21_imag = int_reg_array_48_21_imag;
  assign io_coef_out_payload_0_48_22_real = int_reg_array_48_22_real;
  assign io_coef_out_payload_0_48_22_imag = int_reg_array_48_22_imag;
  assign io_coef_out_payload_0_48_23_real = int_reg_array_48_23_real;
  assign io_coef_out_payload_0_48_23_imag = int_reg_array_48_23_imag;
  assign io_coef_out_payload_0_48_24_real = int_reg_array_48_24_real;
  assign io_coef_out_payload_0_48_24_imag = int_reg_array_48_24_imag;
  assign io_coef_out_payload_0_48_25_real = int_reg_array_48_25_real;
  assign io_coef_out_payload_0_48_25_imag = int_reg_array_48_25_imag;
  assign io_coef_out_payload_0_48_26_real = int_reg_array_48_26_real;
  assign io_coef_out_payload_0_48_26_imag = int_reg_array_48_26_imag;
  assign io_coef_out_payload_0_48_27_real = int_reg_array_48_27_real;
  assign io_coef_out_payload_0_48_27_imag = int_reg_array_48_27_imag;
  assign io_coef_out_payload_0_48_28_real = int_reg_array_48_28_real;
  assign io_coef_out_payload_0_48_28_imag = int_reg_array_48_28_imag;
  assign io_coef_out_payload_0_48_29_real = int_reg_array_48_29_real;
  assign io_coef_out_payload_0_48_29_imag = int_reg_array_48_29_imag;
  assign io_coef_out_payload_0_48_30_real = int_reg_array_48_30_real;
  assign io_coef_out_payload_0_48_30_imag = int_reg_array_48_30_imag;
  assign io_coef_out_payload_0_48_31_real = int_reg_array_48_31_real;
  assign io_coef_out_payload_0_48_31_imag = int_reg_array_48_31_imag;
  assign io_coef_out_payload_0_48_32_real = int_reg_array_48_32_real;
  assign io_coef_out_payload_0_48_32_imag = int_reg_array_48_32_imag;
  assign io_coef_out_payload_0_48_33_real = int_reg_array_48_33_real;
  assign io_coef_out_payload_0_48_33_imag = int_reg_array_48_33_imag;
  assign io_coef_out_payload_0_48_34_real = int_reg_array_48_34_real;
  assign io_coef_out_payload_0_48_34_imag = int_reg_array_48_34_imag;
  assign io_coef_out_payload_0_48_35_real = int_reg_array_48_35_real;
  assign io_coef_out_payload_0_48_35_imag = int_reg_array_48_35_imag;
  assign io_coef_out_payload_0_48_36_real = int_reg_array_48_36_real;
  assign io_coef_out_payload_0_48_36_imag = int_reg_array_48_36_imag;
  assign io_coef_out_payload_0_48_37_real = int_reg_array_48_37_real;
  assign io_coef_out_payload_0_48_37_imag = int_reg_array_48_37_imag;
  assign io_coef_out_payload_0_48_38_real = int_reg_array_48_38_real;
  assign io_coef_out_payload_0_48_38_imag = int_reg_array_48_38_imag;
  assign io_coef_out_payload_0_48_39_real = int_reg_array_48_39_real;
  assign io_coef_out_payload_0_48_39_imag = int_reg_array_48_39_imag;
  assign io_coef_out_payload_0_48_40_real = int_reg_array_48_40_real;
  assign io_coef_out_payload_0_48_40_imag = int_reg_array_48_40_imag;
  assign io_coef_out_payload_0_48_41_real = int_reg_array_48_41_real;
  assign io_coef_out_payload_0_48_41_imag = int_reg_array_48_41_imag;
  assign io_coef_out_payload_0_48_42_real = int_reg_array_48_42_real;
  assign io_coef_out_payload_0_48_42_imag = int_reg_array_48_42_imag;
  assign io_coef_out_payload_0_48_43_real = int_reg_array_48_43_real;
  assign io_coef_out_payload_0_48_43_imag = int_reg_array_48_43_imag;
  assign io_coef_out_payload_0_48_44_real = int_reg_array_48_44_real;
  assign io_coef_out_payload_0_48_44_imag = int_reg_array_48_44_imag;
  assign io_coef_out_payload_0_48_45_real = int_reg_array_48_45_real;
  assign io_coef_out_payload_0_48_45_imag = int_reg_array_48_45_imag;
  assign io_coef_out_payload_0_48_46_real = int_reg_array_48_46_real;
  assign io_coef_out_payload_0_48_46_imag = int_reg_array_48_46_imag;
  assign io_coef_out_payload_0_48_47_real = int_reg_array_48_47_real;
  assign io_coef_out_payload_0_48_47_imag = int_reg_array_48_47_imag;
  assign io_coef_out_payload_0_48_48_real = int_reg_array_48_48_real;
  assign io_coef_out_payload_0_48_48_imag = int_reg_array_48_48_imag;
  assign io_coef_out_payload_0_48_49_real = int_reg_array_48_49_real;
  assign io_coef_out_payload_0_48_49_imag = int_reg_array_48_49_imag;
  assign io_coef_out_payload_0_49_0_real = int_reg_array_49_0_real;
  assign io_coef_out_payload_0_49_0_imag = int_reg_array_49_0_imag;
  assign io_coef_out_payload_0_49_1_real = int_reg_array_49_1_real;
  assign io_coef_out_payload_0_49_1_imag = int_reg_array_49_1_imag;
  assign io_coef_out_payload_0_49_2_real = int_reg_array_49_2_real;
  assign io_coef_out_payload_0_49_2_imag = int_reg_array_49_2_imag;
  assign io_coef_out_payload_0_49_3_real = int_reg_array_49_3_real;
  assign io_coef_out_payload_0_49_3_imag = int_reg_array_49_3_imag;
  assign io_coef_out_payload_0_49_4_real = int_reg_array_49_4_real;
  assign io_coef_out_payload_0_49_4_imag = int_reg_array_49_4_imag;
  assign io_coef_out_payload_0_49_5_real = int_reg_array_49_5_real;
  assign io_coef_out_payload_0_49_5_imag = int_reg_array_49_5_imag;
  assign io_coef_out_payload_0_49_6_real = int_reg_array_49_6_real;
  assign io_coef_out_payload_0_49_6_imag = int_reg_array_49_6_imag;
  assign io_coef_out_payload_0_49_7_real = int_reg_array_49_7_real;
  assign io_coef_out_payload_0_49_7_imag = int_reg_array_49_7_imag;
  assign io_coef_out_payload_0_49_8_real = int_reg_array_49_8_real;
  assign io_coef_out_payload_0_49_8_imag = int_reg_array_49_8_imag;
  assign io_coef_out_payload_0_49_9_real = int_reg_array_49_9_real;
  assign io_coef_out_payload_0_49_9_imag = int_reg_array_49_9_imag;
  assign io_coef_out_payload_0_49_10_real = int_reg_array_49_10_real;
  assign io_coef_out_payload_0_49_10_imag = int_reg_array_49_10_imag;
  assign io_coef_out_payload_0_49_11_real = int_reg_array_49_11_real;
  assign io_coef_out_payload_0_49_11_imag = int_reg_array_49_11_imag;
  assign io_coef_out_payload_0_49_12_real = int_reg_array_49_12_real;
  assign io_coef_out_payload_0_49_12_imag = int_reg_array_49_12_imag;
  assign io_coef_out_payload_0_49_13_real = int_reg_array_49_13_real;
  assign io_coef_out_payload_0_49_13_imag = int_reg_array_49_13_imag;
  assign io_coef_out_payload_0_49_14_real = int_reg_array_49_14_real;
  assign io_coef_out_payload_0_49_14_imag = int_reg_array_49_14_imag;
  assign io_coef_out_payload_0_49_15_real = int_reg_array_49_15_real;
  assign io_coef_out_payload_0_49_15_imag = int_reg_array_49_15_imag;
  assign io_coef_out_payload_0_49_16_real = int_reg_array_49_16_real;
  assign io_coef_out_payload_0_49_16_imag = int_reg_array_49_16_imag;
  assign io_coef_out_payload_0_49_17_real = int_reg_array_49_17_real;
  assign io_coef_out_payload_0_49_17_imag = int_reg_array_49_17_imag;
  assign io_coef_out_payload_0_49_18_real = int_reg_array_49_18_real;
  assign io_coef_out_payload_0_49_18_imag = int_reg_array_49_18_imag;
  assign io_coef_out_payload_0_49_19_real = int_reg_array_49_19_real;
  assign io_coef_out_payload_0_49_19_imag = int_reg_array_49_19_imag;
  assign io_coef_out_payload_0_49_20_real = int_reg_array_49_20_real;
  assign io_coef_out_payload_0_49_20_imag = int_reg_array_49_20_imag;
  assign io_coef_out_payload_0_49_21_real = int_reg_array_49_21_real;
  assign io_coef_out_payload_0_49_21_imag = int_reg_array_49_21_imag;
  assign io_coef_out_payload_0_49_22_real = int_reg_array_49_22_real;
  assign io_coef_out_payload_0_49_22_imag = int_reg_array_49_22_imag;
  assign io_coef_out_payload_0_49_23_real = int_reg_array_49_23_real;
  assign io_coef_out_payload_0_49_23_imag = int_reg_array_49_23_imag;
  assign io_coef_out_payload_0_49_24_real = int_reg_array_49_24_real;
  assign io_coef_out_payload_0_49_24_imag = int_reg_array_49_24_imag;
  assign io_coef_out_payload_0_49_25_real = int_reg_array_49_25_real;
  assign io_coef_out_payload_0_49_25_imag = int_reg_array_49_25_imag;
  assign io_coef_out_payload_0_49_26_real = int_reg_array_49_26_real;
  assign io_coef_out_payload_0_49_26_imag = int_reg_array_49_26_imag;
  assign io_coef_out_payload_0_49_27_real = int_reg_array_49_27_real;
  assign io_coef_out_payload_0_49_27_imag = int_reg_array_49_27_imag;
  assign io_coef_out_payload_0_49_28_real = int_reg_array_49_28_real;
  assign io_coef_out_payload_0_49_28_imag = int_reg_array_49_28_imag;
  assign io_coef_out_payload_0_49_29_real = int_reg_array_49_29_real;
  assign io_coef_out_payload_0_49_29_imag = int_reg_array_49_29_imag;
  assign io_coef_out_payload_0_49_30_real = int_reg_array_49_30_real;
  assign io_coef_out_payload_0_49_30_imag = int_reg_array_49_30_imag;
  assign io_coef_out_payload_0_49_31_real = int_reg_array_49_31_real;
  assign io_coef_out_payload_0_49_31_imag = int_reg_array_49_31_imag;
  assign io_coef_out_payload_0_49_32_real = int_reg_array_49_32_real;
  assign io_coef_out_payload_0_49_32_imag = int_reg_array_49_32_imag;
  assign io_coef_out_payload_0_49_33_real = int_reg_array_49_33_real;
  assign io_coef_out_payload_0_49_33_imag = int_reg_array_49_33_imag;
  assign io_coef_out_payload_0_49_34_real = int_reg_array_49_34_real;
  assign io_coef_out_payload_0_49_34_imag = int_reg_array_49_34_imag;
  assign io_coef_out_payload_0_49_35_real = int_reg_array_49_35_real;
  assign io_coef_out_payload_0_49_35_imag = int_reg_array_49_35_imag;
  assign io_coef_out_payload_0_49_36_real = int_reg_array_49_36_real;
  assign io_coef_out_payload_0_49_36_imag = int_reg_array_49_36_imag;
  assign io_coef_out_payload_0_49_37_real = int_reg_array_49_37_real;
  assign io_coef_out_payload_0_49_37_imag = int_reg_array_49_37_imag;
  assign io_coef_out_payload_0_49_38_real = int_reg_array_49_38_real;
  assign io_coef_out_payload_0_49_38_imag = int_reg_array_49_38_imag;
  assign io_coef_out_payload_0_49_39_real = int_reg_array_49_39_real;
  assign io_coef_out_payload_0_49_39_imag = int_reg_array_49_39_imag;
  assign io_coef_out_payload_0_49_40_real = int_reg_array_49_40_real;
  assign io_coef_out_payload_0_49_40_imag = int_reg_array_49_40_imag;
  assign io_coef_out_payload_0_49_41_real = int_reg_array_49_41_real;
  assign io_coef_out_payload_0_49_41_imag = int_reg_array_49_41_imag;
  assign io_coef_out_payload_0_49_42_real = int_reg_array_49_42_real;
  assign io_coef_out_payload_0_49_42_imag = int_reg_array_49_42_imag;
  assign io_coef_out_payload_0_49_43_real = int_reg_array_49_43_real;
  assign io_coef_out_payload_0_49_43_imag = int_reg_array_49_43_imag;
  assign io_coef_out_payload_0_49_44_real = int_reg_array_49_44_real;
  assign io_coef_out_payload_0_49_44_imag = int_reg_array_49_44_imag;
  assign io_coef_out_payload_0_49_45_real = int_reg_array_49_45_real;
  assign io_coef_out_payload_0_49_45_imag = int_reg_array_49_45_imag;
  assign io_coef_out_payload_0_49_46_real = int_reg_array_49_46_real;
  assign io_coef_out_payload_0_49_46_imag = int_reg_array_49_46_imag;
  assign io_coef_out_payload_0_49_47_real = int_reg_array_49_47_real;
  assign io_coef_out_payload_0_49_47_imag = int_reg_array_49_47_imag;
  assign io_coef_out_payload_0_49_48_real = int_reg_array_49_48_real;
  assign io_coef_out_payload_0_49_48_imag = int_reg_array_49_48_imag;
  assign io_coef_out_payload_0_49_49_real = int_reg_array_49_49_real;
  assign io_coef_out_payload_0_49_49_imag = int_reg_array_49_49_imag;
  always @ (posedge clk) begin
    if(_zz_1_)begin
      _zz_13_ <= _zz_3_;
      _zz_14_ <= _zz_5_;
      _zz_15_ <= _zz_4_;
    end
    if(_zz_7_)begin
      transfer_done <= (((32'h0 <= load_data_area_current_addr) && (load_data_area_current_addr < 32'h0)) ? _zz_9__regNext[0] : _zz_4565_[0]);
      if(_zz_19_)begin
        int_reg_array_0_0_real <= _zz_84_;
      end
      if(_zz_20_)begin
        int_reg_array_0_1_real <= _zz_84_;
      end
      if(_zz_21_)begin
        int_reg_array_0_2_real <= _zz_84_;
      end
      if(_zz_22_)begin
        int_reg_array_0_3_real <= _zz_84_;
      end
      if(_zz_23_)begin
        int_reg_array_0_4_real <= _zz_84_;
      end
      if(_zz_24_)begin
        int_reg_array_0_5_real <= _zz_84_;
      end
      if(_zz_25_)begin
        int_reg_array_0_6_real <= _zz_84_;
      end
      if(_zz_26_)begin
        int_reg_array_0_7_real <= _zz_84_;
      end
      if(_zz_27_)begin
        int_reg_array_0_8_real <= _zz_84_;
      end
      if(_zz_28_)begin
        int_reg_array_0_9_real <= _zz_84_;
      end
      if(_zz_29_)begin
        int_reg_array_0_10_real <= _zz_84_;
      end
      if(_zz_30_)begin
        int_reg_array_0_11_real <= _zz_84_;
      end
      if(_zz_31_)begin
        int_reg_array_0_12_real <= _zz_84_;
      end
      if(_zz_32_)begin
        int_reg_array_0_13_real <= _zz_84_;
      end
      if(_zz_33_)begin
        int_reg_array_0_14_real <= _zz_84_;
      end
      if(_zz_34_)begin
        int_reg_array_0_15_real <= _zz_84_;
      end
      if(_zz_35_)begin
        int_reg_array_0_16_real <= _zz_84_;
      end
      if(_zz_36_)begin
        int_reg_array_0_17_real <= _zz_84_;
      end
      if(_zz_37_)begin
        int_reg_array_0_18_real <= _zz_84_;
      end
      if(_zz_38_)begin
        int_reg_array_0_19_real <= _zz_84_;
      end
      if(_zz_39_)begin
        int_reg_array_0_20_real <= _zz_84_;
      end
      if(_zz_40_)begin
        int_reg_array_0_21_real <= _zz_84_;
      end
      if(_zz_41_)begin
        int_reg_array_0_22_real <= _zz_84_;
      end
      if(_zz_42_)begin
        int_reg_array_0_23_real <= _zz_84_;
      end
      if(_zz_43_)begin
        int_reg_array_0_24_real <= _zz_84_;
      end
      if(_zz_44_)begin
        int_reg_array_0_25_real <= _zz_84_;
      end
      if(_zz_45_)begin
        int_reg_array_0_26_real <= _zz_84_;
      end
      if(_zz_46_)begin
        int_reg_array_0_27_real <= _zz_84_;
      end
      if(_zz_47_)begin
        int_reg_array_0_28_real <= _zz_84_;
      end
      if(_zz_48_)begin
        int_reg_array_0_29_real <= _zz_84_;
      end
      if(_zz_49_)begin
        int_reg_array_0_30_real <= _zz_84_;
      end
      if(_zz_50_)begin
        int_reg_array_0_31_real <= _zz_84_;
      end
      if(_zz_51_)begin
        int_reg_array_0_32_real <= _zz_84_;
      end
      if(_zz_52_)begin
        int_reg_array_0_33_real <= _zz_84_;
      end
      if(_zz_53_)begin
        int_reg_array_0_34_real <= _zz_84_;
      end
      if(_zz_54_)begin
        int_reg_array_0_35_real <= _zz_84_;
      end
      if(_zz_55_)begin
        int_reg_array_0_36_real <= _zz_84_;
      end
      if(_zz_56_)begin
        int_reg_array_0_37_real <= _zz_84_;
      end
      if(_zz_57_)begin
        int_reg_array_0_38_real <= _zz_84_;
      end
      if(_zz_58_)begin
        int_reg_array_0_39_real <= _zz_84_;
      end
      if(_zz_59_)begin
        int_reg_array_0_40_real <= _zz_84_;
      end
      if(_zz_60_)begin
        int_reg_array_0_41_real <= _zz_84_;
      end
      if(_zz_61_)begin
        int_reg_array_0_42_real <= _zz_84_;
      end
      if(_zz_62_)begin
        int_reg_array_0_43_real <= _zz_84_;
      end
      if(_zz_63_)begin
        int_reg_array_0_44_real <= _zz_84_;
      end
      if(_zz_64_)begin
        int_reg_array_0_45_real <= _zz_84_;
      end
      if(_zz_65_)begin
        int_reg_array_0_46_real <= _zz_84_;
      end
      if(_zz_66_)begin
        int_reg_array_0_47_real <= _zz_84_;
      end
      if(_zz_67_)begin
        int_reg_array_0_48_real <= _zz_84_;
      end
      if(_zz_68_)begin
        int_reg_array_0_49_real <= _zz_84_;
      end
      if(_zz_69_)begin
        int_reg_array_0_50_real <= _zz_84_;
      end
      if(_zz_70_)begin
        int_reg_array_0_51_real <= _zz_84_;
      end
      if(_zz_71_)begin
        int_reg_array_0_52_real <= _zz_84_;
      end
      if(_zz_72_)begin
        int_reg_array_0_53_real <= _zz_84_;
      end
      if(_zz_73_)begin
        int_reg_array_0_54_real <= _zz_84_;
      end
      if(_zz_74_)begin
        int_reg_array_0_55_real <= _zz_84_;
      end
      if(_zz_75_)begin
        int_reg_array_0_56_real <= _zz_84_;
      end
      if(_zz_76_)begin
        int_reg_array_0_57_real <= _zz_84_;
      end
      if(_zz_77_)begin
        int_reg_array_0_58_real <= _zz_84_;
      end
      if(_zz_78_)begin
        int_reg_array_0_59_real <= _zz_84_;
      end
      if(_zz_79_)begin
        int_reg_array_0_60_real <= _zz_84_;
      end
      if(_zz_80_)begin
        int_reg_array_0_61_real <= _zz_84_;
      end
      if(_zz_81_)begin
        int_reg_array_0_62_real <= _zz_84_;
      end
      if(_zz_82_)begin
        int_reg_array_0_63_real <= _zz_84_;
      end
      if(_zz_19_)begin
        int_reg_array_0_0_imag <= _zz_85_;
      end
      if(_zz_20_)begin
        int_reg_array_0_1_imag <= _zz_85_;
      end
      if(_zz_21_)begin
        int_reg_array_0_2_imag <= _zz_85_;
      end
      if(_zz_22_)begin
        int_reg_array_0_3_imag <= _zz_85_;
      end
      if(_zz_23_)begin
        int_reg_array_0_4_imag <= _zz_85_;
      end
      if(_zz_24_)begin
        int_reg_array_0_5_imag <= _zz_85_;
      end
      if(_zz_25_)begin
        int_reg_array_0_6_imag <= _zz_85_;
      end
      if(_zz_26_)begin
        int_reg_array_0_7_imag <= _zz_85_;
      end
      if(_zz_27_)begin
        int_reg_array_0_8_imag <= _zz_85_;
      end
      if(_zz_28_)begin
        int_reg_array_0_9_imag <= _zz_85_;
      end
      if(_zz_29_)begin
        int_reg_array_0_10_imag <= _zz_85_;
      end
      if(_zz_30_)begin
        int_reg_array_0_11_imag <= _zz_85_;
      end
      if(_zz_31_)begin
        int_reg_array_0_12_imag <= _zz_85_;
      end
      if(_zz_32_)begin
        int_reg_array_0_13_imag <= _zz_85_;
      end
      if(_zz_33_)begin
        int_reg_array_0_14_imag <= _zz_85_;
      end
      if(_zz_34_)begin
        int_reg_array_0_15_imag <= _zz_85_;
      end
      if(_zz_35_)begin
        int_reg_array_0_16_imag <= _zz_85_;
      end
      if(_zz_36_)begin
        int_reg_array_0_17_imag <= _zz_85_;
      end
      if(_zz_37_)begin
        int_reg_array_0_18_imag <= _zz_85_;
      end
      if(_zz_38_)begin
        int_reg_array_0_19_imag <= _zz_85_;
      end
      if(_zz_39_)begin
        int_reg_array_0_20_imag <= _zz_85_;
      end
      if(_zz_40_)begin
        int_reg_array_0_21_imag <= _zz_85_;
      end
      if(_zz_41_)begin
        int_reg_array_0_22_imag <= _zz_85_;
      end
      if(_zz_42_)begin
        int_reg_array_0_23_imag <= _zz_85_;
      end
      if(_zz_43_)begin
        int_reg_array_0_24_imag <= _zz_85_;
      end
      if(_zz_44_)begin
        int_reg_array_0_25_imag <= _zz_85_;
      end
      if(_zz_45_)begin
        int_reg_array_0_26_imag <= _zz_85_;
      end
      if(_zz_46_)begin
        int_reg_array_0_27_imag <= _zz_85_;
      end
      if(_zz_47_)begin
        int_reg_array_0_28_imag <= _zz_85_;
      end
      if(_zz_48_)begin
        int_reg_array_0_29_imag <= _zz_85_;
      end
      if(_zz_49_)begin
        int_reg_array_0_30_imag <= _zz_85_;
      end
      if(_zz_50_)begin
        int_reg_array_0_31_imag <= _zz_85_;
      end
      if(_zz_51_)begin
        int_reg_array_0_32_imag <= _zz_85_;
      end
      if(_zz_52_)begin
        int_reg_array_0_33_imag <= _zz_85_;
      end
      if(_zz_53_)begin
        int_reg_array_0_34_imag <= _zz_85_;
      end
      if(_zz_54_)begin
        int_reg_array_0_35_imag <= _zz_85_;
      end
      if(_zz_55_)begin
        int_reg_array_0_36_imag <= _zz_85_;
      end
      if(_zz_56_)begin
        int_reg_array_0_37_imag <= _zz_85_;
      end
      if(_zz_57_)begin
        int_reg_array_0_38_imag <= _zz_85_;
      end
      if(_zz_58_)begin
        int_reg_array_0_39_imag <= _zz_85_;
      end
      if(_zz_59_)begin
        int_reg_array_0_40_imag <= _zz_85_;
      end
      if(_zz_60_)begin
        int_reg_array_0_41_imag <= _zz_85_;
      end
      if(_zz_61_)begin
        int_reg_array_0_42_imag <= _zz_85_;
      end
      if(_zz_62_)begin
        int_reg_array_0_43_imag <= _zz_85_;
      end
      if(_zz_63_)begin
        int_reg_array_0_44_imag <= _zz_85_;
      end
      if(_zz_64_)begin
        int_reg_array_0_45_imag <= _zz_85_;
      end
      if(_zz_65_)begin
        int_reg_array_0_46_imag <= _zz_85_;
      end
      if(_zz_66_)begin
        int_reg_array_0_47_imag <= _zz_85_;
      end
      if(_zz_67_)begin
        int_reg_array_0_48_imag <= _zz_85_;
      end
      if(_zz_68_)begin
        int_reg_array_0_49_imag <= _zz_85_;
      end
      if(_zz_69_)begin
        int_reg_array_0_50_imag <= _zz_85_;
      end
      if(_zz_70_)begin
        int_reg_array_0_51_imag <= _zz_85_;
      end
      if(_zz_71_)begin
        int_reg_array_0_52_imag <= _zz_85_;
      end
      if(_zz_72_)begin
        int_reg_array_0_53_imag <= _zz_85_;
      end
      if(_zz_73_)begin
        int_reg_array_0_54_imag <= _zz_85_;
      end
      if(_zz_74_)begin
        int_reg_array_0_55_imag <= _zz_85_;
      end
      if(_zz_75_)begin
        int_reg_array_0_56_imag <= _zz_85_;
      end
      if(_zz_76_)begin
        int_reg_array_0_57_imag <= _zz_85_;
      end
      if(_zz_77_)begin
        int_reg_array_0_58_imag <= _zz_85_;
      end
      if(_zz_78_)begin
        int_reg_array_0_59_imag <= _zz_85_;
      end
      if(_zz_79_)begin
        int_reg_array_0_60_imag <= _zz_85_;
      end
      if(_zz_80_)begin
        int_reg_array_0_61_imag <= _zz_85_;
      end
      if(_zz_81_)begin
        int_reg_array_0_62_imag <= _zz_85_;
      end
      if(_zz_82_)begin
        int_reg_array_0_63_imag <= _zz_85_;
      end
      if(_zz_88_)begin
        int_reg_array_1_0_real <= _zz_153_;
      end
      if(_zz_89_)begin
        int_reg_array_1_1_real <= _zz_153_;
      end
      if(_zz_90_)begin
        int_reg_array_1_2_real <= _zz_153_;
      end
      if(_zz_91_)begin
        int_reg_array_1_3_real <= _zz_153_;
      end
      if(_zz_92_)begin
        int_reg_array_1_4_real <= _zz_153_;
      end
      if(_zz_93_)begin
        int_reg_array_1_5_real <= _zz_153_;
      end
      if(_zz_94_)begin
        int_reg_array_1_6_real <= _zz_153_;
      end
      if(_zz_95_)begin
        int_reg_array_1_7_real <= _zz_153_;
      end
      if(_zz_96_)begin
        int_reg_array_1_8_real <= _zz_153_;
      end
      if(_zz_97_)begin
        int_reg_array_1_9_real <= _zz_153_;
      end
      if(_zz_98_)begin
        int_reg_array_1_10_real <= _zz_153_;
      end
      if(_zz_99_)begin
        int_reg_array_1_11_real <= _zz_153_;
      end
      if(_zz_100_)begin
        int_reg_array_1_12_real <= _zz_153_;
      end
      if(_zz_101_)begin
        int_reg_array_1_13_real <= _zz_153_;
      end
      if(_zz_102_)begin
        int_reg_array_1_14_real <= _zz_153_;
      end
      if(_zz_103_)begin
        int_reg_array_1_15_real <= _zz_153_;
      end
      if(_zz_104_)begin
        int_reg_array_1_16_real <= _zz_153_;
      end
      if(_zz_105_)begin
        int_reg_array_1_17_real <= _zz_153_;
      end
      if(_zz_106_)begin
        int_reg_array_1_18_real <= _zz_153_;
      end
      if(_zz_107_)begin
        int_reg_array_1_19_real <= _zz_153_;
      end
      if(_zz_108_)begin
        int_reg_array_1_20_real <= _zz_153_;
      end
      if(_zz_109_)begin
        int_reg_array_1_21_real <= _zz_153_;
      end
      if(_zz_110_)begin
        int_reg_array_1_22_real <= _zz_153_;
      end
      if(_zz_111_)begin
        int_reg_array_1_23_real <= _zz_153_;
      end
      if(_zz_112_)begin
        int_reg_array_1_24_real <= _zz_153_;
      end
      if(_zz_113_)begin
        int_reg_array_1_25_real <= _zz_153_;
      end
      if(_zz_114_)begin
        int_reg_array_1_26_real <= _zz_153_;
      end
      if(_zz_115_)begin
        int_reg_array_1_27_real <= _zz_153_;
      end
      if(_zz_116_)begin
        int_reg_array_1_28_real <= _zz_153_;
      end
      if(_zz_117_)begin
        int_reg_array_1_29_real <= _zz_153_;
      end
      if(_zz_118_)begin
        int_reg_array_1_30_real <= _zz_153_;
      end
      if(_zz_119_)begin
        int_reg_array_1_31_real <= _zz_153_;
      end
      if(_zz_120_)begin
        int_reg_array_1_32_real <= _zz_153_;
      end
      if(_zz_121_)begin
        int_reg_array_1_33_real <= _zz_153_;
      end
      if(_zz_122_)begin
        int_reg_array_1_34_real <= _zz_153_;
      end
      if(_zz_123_)begin
        int_reg_array_1_35_real <= _zz_153_;
      end
      if(_zz_124_)begin
        int_reg_array_1_36_real <= _zz_153_;
      end
      if(_zz_125_)begin
        int_reg_array_1_37_real <= _zz_153_;
      end
      if(_zz_126_)begin
        int_reg_array_1_38_real <= _zz_153_;
      end
      if(_zz_127_)begin
        int_reg_array_1_39_real <= _zz_153_;
      end
      if(_zz_128_)begin
        int_reg_array_1_40_real <= _zz_153_;
      end
      if(_zz_129_)begin
        int_reg_array_1_41_real <= _zz_153_;
      end
      if(_zz_130_)begin
        int_reg_array_1_42_real <= _zz_153_;
      end
      if(_zz_131_)begin
        int_reg_array_1_43_real <= _zz_153_;
      end
      if(_zz_132_)begin
        int_reg_array_1_44_real <= _zz_153_;
      end
      if(_zz_133_)begin
        int_reg_array_1_45_real <= _zz_153_;
      end
      if(_zz_134_)begin
        int_reg_array_1_46_real <= _zz_153_;
      end
      if(_zz_135_)begin
        int_reg_array_1_47_real <= _zz_153_;
      end
      if(_zz_136_)begin
        int_reg_array_1_48_real <= _zz_153_;
      end
      if(_zz_137_)begin
        int_reg_array_1_49_real <= _zz_153_;
      end
      if(_zz_138_)begin
        int_reg_array_1_50_real <= _zz_153_;
      end
      if(_zz_139_)begin
        int_reg_array_1_51_real <= _zz_153_;
      end
      if(_zz_140_)begin
        int_reg_array_1_52_real <= _zz_153_;
      end
      if(_zz_141_)begin
        int_reg_array_1_53_real <= _zz_153_;
      end
      if(_zz_142_)begin
        int_reg_array_1_54_real <= _zz_153_;
      end
      if(_zz_143_)begin
        int_reg_array_1_55_real <= _zz_153_;
      end
      if(_zz_144_)begin
        int_reg_array_1_56_real <= _zz_153_;
      end
      if(_zz_145_)begin
        int_reg_array_1_57_real <= _zz_153_;
      end
      if(_zz_146_)begin
        int_reg_array_1_58_real <= _zz_153_;
      end
      if(_zz_147_)begin
        int_reg_array_1_59_real <= _zz_153_;
      end
      if(_zz_148_)begin
        int_reg_array_1_60_real <= _zz_153_;
      end
      if(_zz_149_)begin
        int_reg_array_1_61_real <= _zz_153_;
      end
      if(_zz_150_)begin
        int_reg_array_1_62_real <= _zz_153_;
      end
      if(_zz_151_)begin
        int_reg_array_1_63_real <= _zz_153_;
      end
      if(_zz_88_)begin
        int_reg_array_1_0_imag <= _zz_154_;
      end
      if(_zz_89_)begin
        int_reg_array_1_1_imag <= _zz_154_;
      end
      if(_zz_90_)begin
        int_reg_array_1_2_imag <= _zz_154_;
      end
      if(_zz_91_)begin
        int_reg_array_1_3_imag <= _zz_154_;
      end
      if(_zz_92_)begin
        int_reg_array_1_4_imag <= _zz_154_;
      end
      if(_zz_93_)begin
        int_reg_array_1_5_imag <= _zz_154_;
      end
      if(_zz_94_)begin
        int_reg_array_1_6_imag <= _zz_154_;
      end
      if(_zz_95_)begin
        int_reg_array_1_7_imag <= _zz_154_;
      end
      if(_zz_96_)begin
        int_reg_array_1_8_imag <= _zz_154_;
      end
      if(_zz_97_)begin
        int_reg_array_1_9_imag <= _zz_154_;
      end
      if(_zz_98_)begin
        int_reg_array_1_10_imag <= _zz_154_;
      end
      if(_zz_99_)begin
        int_reg_array_1_11_imag <= _zz_154_;
      end
      if(_zz_100_)begin
        int_reg_array_1_12_imag <= _zz_154_;
      end
      if(_zz_101_)begin
        int_reg_array_1_13_imag <= _zz_154_;
      end
      if(_zz_102_)begin
        int_reg_array_1_14_imag <= _zz_154_;
      end
      if(_zz_103_)begin
        int_reg_array_1_15_imag <= _zz_154_;
      end
      if(_zz_104_)begin
        int_reg_array_1_16_imag <= _zz_154_;
      end
      if(_zz_105_)begin
        int_reg_array_1_17_imag <= _zz_154_;
      end
      if(_zz_106_)begin
        int_reg_array_1_18_imag <= _zz_154_;
      end
      if(_zz_107_)begin
        int_reg_array_1_19_imag <= _zz_154_;
      end
      if(_zz_108_)begin
        int_reg_array_1_20_imag <= _zz_154_;
      end
      if(_zz_109_)begin
        int_reg_array_1_21_imag <= _zz_154_;
      end
      if(_zz_110_)begin
        int_reg_array_1_22_imag <= _zz_154_;
      end
      if(_zz_111_)begin
        int_reg_array_1_23_imag <= _zz_154_;
      end
      if(_zz_112_)begin
        int_reg_array_1_24_imag <= _zz_154_;
      end
      if(_zz_113_)begin
        int_reg_array_1_25_imag <= _zz_154_;
      end
      if(_zz_114_)begin
        int_reg_array_1_26_imag <= _zz_154_;
      end
      if(_zz_115_)begin
        int_reg_array_1_27_imag <= _zz_154_;
      end
      if(_zz_116_)begin
        int_reg_array_1_28_imag <= _zz_154_;
      end
      if(_zz_117_)begin
        int_reg_array_1_29_imag <= _zz_154_;
      end
      if(_zz_118_)begin
        int_reg_array_1_30_imag <= _zz_154_;
      end
      if(_zz_119_)begin
        int_reg_array_1_31_imag <= _zz_154_;
      end
      if(_zz_120_)begin
        int_reg_array_1_32_imag <= _zz_154_;
      end
      if(_zz_121_)begin
        int_reg_array_1_33_imag <= _zz_154_;
      end
      if(_zz_122_)begin
        int_reg_array_1_34_imag <= _zz_154_;
      end
      if(_zz_123_)begin
        int_reg_array_1_35_imag <= _zz_154_;
      end
      if(_zz_124_)begin
        int_reg_array_1_36_imag <= _zz_154_;
      end
      if(_zz_125_)begin
        int_reg_array_1_37_imag <= _zz_154_;
      end
      if(_zz_126_)begin
        int_reg_array_1_38_imag <= _zz_154_;
      end
      if(_zz_127_)begin
        int_reg_array_1_39_imag <= _zz_154_;
      end
      if(_zz_128_)begin
        int_reg_array_1_40_imag <= _zz_154_;
      end
      if(_zz_129_)begin
        int_reg_array_1_41_imag <= _zz_154_;
      end
      if(_zz_130_)begin
        int_reg_array_1_42_imag <= _zz_154_;
      end
      if(_zz_131_)begin
        int_reg_array_1_43_imag <= _zz_154_;
      end
      if(_zz_132_)begin
        int_reg_array_1_44_imag <= _zz_154_;
      end
      if(_zz_133_)begin
        int_reg_array_1_45_imag <= _zz_154_;
      end
      if(_zz_134_)begin
        int_reg_array_1_46_imag <= _zz_154_;
      end
      if(_zz_135_)begin
        int_reg_array_1_47_imag <= _zz_154_;
      end
      if(_zz_136_)begin
        int_reg_array_1_48_imag <= _zz_154_;
      end
      if(_zz_137_)begin
        int_reg_array_1_49_imag <= _zz_154_;
      end
      if(_zz_138_)begin
        int_reg_array_1_50_imag <= _zz_154_;
      end
      if(_zz_139_)begin
        int_reg_array_1_51_imag <= _zz_154_;
      end
      if(_zz_140_)begin
        int_reg_array_1_52_imag <= _zz_154_;
      end
      if(_zz_141_)begin
        int_reg_array_1_53_imag <= _zz_154_;
      end
      if(_zz_142_)begin
        int_reg_array_1_54_imag <= _zz_154_;
      end
      if(_zz_143_)begin
        int_reg_array_1_55_imag <= _zz_154_;
      end
      if(_zz_144_)begin
        int_reg_array_1_56_imag <= _zz_154_;
      end
      if(_zz_145_)begin
        int_reg_array_1_57_imag <= _zz_154_;
      end
      if(_zz_146_)begin
        int_reg_array_1_58_imag <= _zz_154_;
      end
      if(_zz_147_)begin
        int_reg_array_1_59_imag <= _zz_154_;
      end
      if(_zz_148_)begin
        int_reg_array_1_60_imag <= _zz_154_;
      end
      if(_zz_149_)begin
        int_reg_array_1_61_imag <= _zz_154_;
      end
      if(_zz_150_)begin
        int_reg_array_1_62_imag <= _zz_154_;
      end
      if(_zz_151_)begin
        int_reg_array_1_63_imag <= _zz_154_;
      end
      if(_zz_157_)begin
        int_reg_array_2_0_real <= _zz_222_;
      end
      if(_zz_158_)begin
        int_reg_array_2_1_real <= _zz_222_;
      end
      if(_zz_159_)begin
        int_reg_array_2_2_real <= _zz_222_;
      end
      if(_zz_160_)begin
        int_reg_array_2_3_real <= _zz_222_;
      end
      if(_zz_161_)begin
        int_reg_array_2_4_real <= _zz_222_;
      end
      if(_zz_162_)begin
        int_reg_array_2_5_real <= _zz_222_;
      end
      if(_zz_163_)begin
        int_reg_array_2_6_real <= _zz_222_;
      end
      if(_zz_164_)begin
        int_reg_array_2_7_real <= _zz_222_;
      end
      if(_zz_165_)begin
        int_reg_array_2_8_real <= _zz_222_;
      end
      if(_zz_166_)begin
        int_reg_array_2_9_real <= _zz_222_;
      end
      if(_zz_167_)begin
        int_reg_array_2_10_real <= _zz_222_;
      end
      if(_zz_168_)begin
        int_reg_array_2_11_real <= _zz_222_;
      end
      if(_zz_169_)begin
        int_reg_array_2_12_real <= _zz_222_;
      end
      if(_zz_170_)begin
        int_reg_array_2_13_real <= _zz_222_;
      end
      if(_zz_171_)begin
        int_reg_array_2_14_real <= _zz_222_;
      end
      if(_zz_172_)begin
        int_reg_array_2_15_real <= _zz_222_;
      end
      if(_zz_173_)begin
        int_reg_array_2_16_real <= _zz_222_;
      end
      if(_zz_174_)begin
        int_reg_array_2_17_real <= _zz_222_;
      end
      if(_zz_175_)begin
        int_reg_array_2_18_real <= _zz_222_;
      end
      if(_zz_176_)begin
        int_reg_array_2_19_real <= _zz_222_;
      end
      if(_zz_177_)begin
        int_reg_array_2_20_real <= _zz_222_;
      end
      if(_zz_178_)begin
        int_reg_array_2_21_real <= _zz_222_;
      end
      if(_zz_179_)begin
        int_reg_array_2_22_real <= _zz_222_;
      end
      if(_zz_180_)begin
        int_reg_array_2_23_real <= _zz_222_;
      end
      if(_zz_181_)begin
        int_reg_array_2_24_real <= _zz_222_;
      end
      if(_zz_182_)begin
        int_reg_array_2_25_real <= _zz_222_;
      end
      if(_zz_183_)begin
        int_reg_array_2_26_real <= _zz_222_;
      end
      if(_zz_184_)begin
        int_reg_array_2_27_real <= _zz_222_;
      end
      if(_zz_185_)begin
        int_reg_array_2_28_real <= _zz_222_;
      end
      if(_zz_186_)begin
        int_reg_array_2_29_real <= _zz_222_;
      end
      if(_zz_187_)begin
        int_reg_array_2_30_real <= _zz_222_;
      end
      if(_zz_188_)begin
        int_reg_array_2_31_real <= _zz_222_;
      end
      if(_zz_189_)begin
        int_reg_array_2_32_real <= _zz_222_;
      end
      if(_zz_190_)begin
        int_reg_array_2_33_real <= _zz_222_;
      end
      if(_zz_191_)begin
        int_reg_array_2_34_real <= _zz_222_;
      end
      if(_zz_192_)begin
        int_reg_array_2_35_real <= _zz_222_;
      end
      if(_zz_193_)begin
        int_reg_array_2_36_real <= _zz_222_;
      end
      if(_zz_194_)begin
        int_reg_array_2_37_real <= _zz_222_;
      end
      if(_zz_195_)begin
        int_reg_array_2_38_real <= _zz_222_;
      end
      if(_zz_196_)begin
        int_reg_array_2_39_real <= _zz_222_;
      end
      if(_zz_197_)begin
        int_reg_array_2_40_real <= _zz_222_;
      end
      if(_zz_198_)begin
        int_reg_array_2_41_real <= _zz_222_;
      end
      if(_zz_199_)begin
        int_reg_array_2_42_real <= _zz_222_;
      end
      if(_zz_200_)begin
        int_reg_array_2_43_real <= _zz_222_;
      end
      if(_zz_201_)begin
        int_reg_array_2_44_real <= _zz_222_;
      end
      if(_zz_202_)begin
        int_reg_array_2_45_real <= _zz_222_;
      end
      if(_zz_203_)begin
        int_reg_array_2_46_real <= _zz_222_;
      end
      if(_zz_204_)begin
        int_reg_array_2_47_real <= _zz_222_;
      end
      if(_zz_205_)begin
        int_reg_array_2_48_real <= _zz_222_;
      end
      if(_zz_206_)begin
        int_reg_array_2_49_real <= _zz_222_;
      end
      if(_zz_207_)begin
        int_reg_array_2_50_real <= _zz_222_;
      end
      if(_zz_208_)begin
        int_reg_array_2_51_real <= _zz_222_;
      end
      if(_zz_209_)begin
        int_reg_array_2_52_real <= _zz_222_;
      end
      if(_zz_210_)begin
        int_reg_array_2_53_real <= _zz_222_;
      end
      if(_zz_211_)begin
        int_reg_array_2_54_real <= _zz_222_;
      end
      if(_zz_212_)begin
        int_reg_array_2_55_real <= _zz_222_;
      end
      if(_zz_213_)begin
        int_reg_array_2_56_real <= _zz_222_;
      end
      if(_zz_214_)begin
        int_reg_array_2_57_real <= _zz_222_;
      end
      if(_zz_215_)begin
        int_reg_array_2_58_real <= _zz_222_;
      end
      if(_zz_216_)begin
        int_reg_array_2_59_real <= _zz_222_;
      end
      if(_zz_217_)begin
        int_reg_array_2_60_real <= _zz_222_;
      end
      if(_zz_218_)begin
        int_reg_array_2_61_real <= _zz_222_;
      end
      if(_zz_219_)begin
        int_reg_array_2_62_real <= _zz_222_;
      end
      if(_zz_220_)begin
        int_reg_array_2_63_real <= _zz_222_;
      end
      if(_zz_157_)begin
        int_reg_array_2_0_imag <= _zz_223_;
      end
      if(_zz_158_)begin
        int_reg_array_2_1_imag <= _zz_223_;
      end
      if(_zz_159_)begin
        int_reg_array_2_2_imag <= _zz_223_;
      end
      if(_zz_160_)begin
        int_reg_array_2_3_imag <= _zz_223_;
      end
      if(_zz_161_)begin
        int_reg_array_2_4_imag <= _zz_223_;
      end
      if(_zz_162_)begin
        int_reg_array_2_5_imag <= _zz_223_;
      end
      if(_zz_163_)begin
        int_reg_array_2_6_imag <= _zz_223_;
      end
      if(_zz_164_)begin
        int_reg_array_2_7_imag <= _zz_223_;
      end
      if(_zz_165_)begin
        int_reg_array_2_8_imag <= _zz_223_;
      end
      if(_zz_166_)begin
        int_reg_array_2_9_imag <= _zz_223_;
      end
      if(_zz_167_)begin
        int_reg_array_2_10_imag <= _zz_223_;
      end
      if(_zz_168_)begin
        int_reg_array_2_11_imag <= _zz_223_;
      end
      if(_zz_169_)begin
        int_reg_array_2_12_imag <= _zz_223_;
      end
      if(_zz_170_)begin
        int_reg_array_2_13_imag <= _zz_223_;
      end
      if(_zz_171_)begin
        int_reg_array_2_14_imag <= _zz_223_;
      end
      if(_zz_172_)begin
        int_reg_array_2_15_imag <= _zz_223_;
      end
      if(_zz_173_)begin
        int_reg_array_2_16_imag <= _zz_223_;
      end
      if(_zz_174_)begin
        int_reg_array_2_17_imag <= _zz_223_;
      end
      if(_zz_175_)begin
        int_reg_array_2_18_imag <= _zz_223_;
      end
      if(_zz_176_)begin
        int_reg_array_2_19_imag <= _zz_223_;
      end
      if(_zz_177_)begin
        int_reg_array_2_20_imag <= _zz_223_;
      end
      if(_zz_178_)begin
        int_reg_array_2_21_imag <= _zz_223_;
      end
      if(_zz_179_)begin
        int_reg_array_2_22_imag <= _zz_223_;
      end
      if(_zz_180_)begin
        int_reg_array_2_23_imag <= _zz_223_;
      end
      if(_zz_181_)begin
        int_reg_array_2_24_imag <= _zz_223_;
      end
      if(_zz_182_)begin
        int_reg_array_2_25_imag <= _zz_223_;
      end
      if(_zz_183_)begin
        int_reg_array_2_26_imag <= _zz_223_;
      end
      if(_zz_184_)begin
        int_reg_array_2_27_imag <= _zz_223_;
      end
      if(_zz_185_)begin
        int_reg_array_2_28_imag <= _zz_223_;
      end
      if(_zz_186_)begin
        int_reg_array_2_29_imag <= _zz_223_;
      end
      if(_zz_187_)begin
        int_reg_array_2_30_imag <= _zz_223_;
      end
      if(_zz_188_)begin
        int_reg_array_2_31_imag <= _zz_223_;
      end
      if(_zz_189_)begin
        int_reg_array_2_32_imag <= _zz_223_;
      end
      if(_zz_190_)begin
        int_reg_array_2_33_imag <= _zz_223_;
      end
      if(_zz_191_)begin
        int_reg_array_2_34_imag <= _zz_223_;
      end
      if(_zz_192_)begin
        int_reg_array_2_35_imag <= _zz_223_;
      end
      if(_zz_193_)begin
        int_reg_array_2_36_imag <= _zz_223_;
      end
      if(_zz_194_)begin
        int_reg_array_2_37_imag <= _zz_223_;
      end
      if(_zz_195_)begin
        int_reg_array_2_38_imag <= _zz_223_;
      end
      if(_zz_196_)begin
        int_reg_array_2_39_imag <= _zz_223_;
      end
      if(_zz_197_)begin
        int_reg_array_2_40_imag <= _zz_223_;
      end
      if(_zz_198_)begin
        int_reg_array_2_41_imag <= _zz_223_;
      end
      if(_zz_199_)begin
        int_reg_array_2_42_imag <= _zz_223_;
      end
      if(_zz_200_)begin
        int_reg_array_2_43_imag <= _zz_223_;
      end
      if(_zz_201_)begin
        int_reg_array_2_44_imag <= _zz_223_;
      end
      if(_zz_202_)begin
        int_reg_array_2_45_imag <= _zz_223_;
      end
      if(_zz_203_)begin
        int_reg_array_2_46_imag <= _zz_223_;
      end
      if(_zz_204_)begin
        int_reg_array_2_47_imag <= _zz_223_;
      end
      if(_zz_205_)begin
        int_reg_array_2_48_imag <= _zz_223_;
      end
      if(_zz_206_)begin
        int_reg_array_2_49_imag <= _zz_223_;
      end
      if(_zz_207_)begin
        int_reg_array_2_50_imag <= _zz_223_;
      end
      if(_zz_208_)begin
        int_reg_array_2_51_imag <= _zz_223_;
      end
      if(_zz_209_)begin
        int_reg_array_2_52_imag <= _zz_223_;
      end
      if(_zz_210_)begin
        int_reg_array_2_53_imag <= _zz_223_;
      end
      if(_zz_211_)begin
        int_reg_array_2_54_imag <= _zz_223_;
      end
      if(_zz_212_)begin
        int_reg_array_2_55_imag <= _zz_223_;
      end
      if(_zz_213_)begin
        int_reg_array_2_56_imag <= _zz_223_;
      end
      if(_zz_214_)begin
        int_reg_array_2_57_imag <= _zz_223_;
      end
      if(_zz_215_)begin
        int_reg_array_2_58_imag <= _zz_223_;
      end
      if(_zz_216_)begin
        int_reg_array_2_59_imag <= _zz_223_;
      end
      if(_zz_217_)begin
        int_reg_array_2_60_imag <= _zz_223_;
      end
      if(_zz_218_)begin
        int_reg_array_2_61_imag <= _zz_223_;
      end
      if(_zz_219_)begin
        int_reg_array_2_62_imag <= _zz_223_;
      end
      if(_zz_220_)begin
        int_reg_array_2_63_imag <= _zz_223_;
      end
      if(_zz_226_)begin
        int_reg_array_3_0_real <= _zz_291_;
      end
      if(_zz_227_)begin
        int_reg_array_3_1_real <= _zz_291_;
      end
      if(_zz_228_)begin
        int_reg_array_3_2_real <= _zz_291_;
      end
      if(_zz_229_)begin
        int_reg_array_3_3_real <= _zz_291_;
      end
      if(_zz_230_)begin
        int_reg_array_3_4_real <= _zz_291_;
      end
      if(_zz_231_)begin
        int_reg_array_3_5_real <= _zz_291_;
      end
      if(_zz_232_)begin
        int_reg_array_3_6_real <= _zz_291_;
      end
      if(_zz_233_)begin
        int_reg_array_3_7_real <= _zz_291_;
      end
      if(_zz_234_)begin
        int_reg_array_3_8_real <= _zz_291_;
      end
      if(_zz_235_)begin
        int_reg_array_3_9_real <= _zz_291_;
      end
      if(_zz_236_)begin
        int_reg_array_3_10_real <= _zz_291_;
      end
      if(_zz_237_)begin
        int_reg_array_3_11_real <= _zz_291_;
      end
      if(_zz_238_)begin
        int_reg_array_3_12_real <= _zz_291_;
      end
      if(_zz_239_)begin
        int_reg_array_3_13_real <= _zz_291_;
      end
      if(_zz_240_)begin
        int_reg_array_3_14_real <= _zz_291_;
      end
      if(_zz_241_)begin
        int_reg_array_3_15_real <= _zz_291_;
      end
      if(_zz_242_)begin
        int_reg_array_3_16_real <= _zz_291_;
      end
      if(_zz_243_)begin
        int_reg_array_3_17_real <= _zz_291_;
      end
      if(_zz_244_)begin
        int_reg_array_3_18_real <= _zz_291_;
      end
      if(_zz_245_)begin
        int_reg_array_3_19_real <= _zz_291_;
      end
      if(_zz_246_)begin
        int_reg_array_3_20_real <= _zz_291_;
      end
      if(_zz_247_)begin
        int_reg_array_3_21_real <= _zz_291_;
      end
      if(_zz_248_)begin
        int_reg_array_3_22_real <= _zz_291_;
      end
      if(_zz_249_)begin
        int_reg_array_3_23_real <= _zz_291_;
      end
      if(_zz_250_)begin
        int_reg_array_3_24_real <= _zz_291_;
      end
      if(_zz_251_)begin
        int_reg_array_3_25_real <= _zz_291_;
      end
      if(_zz_252_)begin
        int_reg_array_3_26_real <= _zz_291_;
      end
      if(_zz_253_)begin
        int_reg_array_3_27_real <= _zz_291_;
      end
      if(_zz_254_)begin
        int_reg_array_3_28_real <= _zz_291_;
      end
      if(_zz_255_)begin
        int_reg_array_3_29_real <= _zz_291_;
      end
      if(_zz_256_)begin
        int_reg_array_3_30_real <= _zz_291_;
      end
      if(_zz_257_)begin
        int_reg_array_3_31_real <= _zz_291_;
      end
      if(_zz_258_)begin
        int_reg_array_3_32_real <= _zz_291_;
      end
      if(_zz_259_)begin
        int_reg_array_3_33_real <= _zz_291_;
      end
      if(_zz_260_)begin
        int_reg_array_3_34_real <= _zz_291_;
      end
      if(_zz_261_)begin
        int_reg_array_3_35_real <= _zz_291_;
      end
      if(_zz_262_)begin
        int_reg_array_3_36_real <= _zz_291_;
      end
      if(_zz_263_)begin
        int_reg_array_3_37_real <= _zz_291_;
      end
      if(_zz_264_)begin
        int_reg_array_3_38_real <= _zz_291_;
      end
      if(_zz_265_)begin
        int_reg_array_3_39_real <= _zz_291_;
      end
      if(_zz_266_)begin
        int_reg_array_3_40_real <= _zz_291_;
      end
      if(_zz_267_)begin
        int_reg_array_3_41_real <= _zz_291_;
      end
      if(_zz_268_)begin
        int_reg_array_3_42_real <= _zz_291_;
      end
      if(_zz_269_)begin
        int_reg_array_3_43_real <= _zz_291_;
      end
      if(_zz_270_)begin
        int_reg_array_3_44_real <= _zz_291_;
      end
      if(_zz_271_)begin
        int_reg_array_3_45_real <= _zz_291_;
      end
      if(_zz_272_)begin
        int_reg_array_3_46_real <= _zz_291_;
      end
      if(_zz_273_)begin
        int_reg_array_3_47_real <= _zz_291_;
      end
      if(_zz_274_)begin
        int_reg_array_3_48_real <= _zz_291_;
      end
      if(_zz_275_)begin
        int_reg_array_3_49_real <= _zz_291_;
      end
      if(_zz_276_)begin
        int_reg_array_3_50_real <= _zz_291_;
      end
      if(_zz_277_)begin
        int_reg_array_3_51_real <= _zz_291_;
      end
      if(_zz_278_)begin
        int_reg_array_3_52_real <= _zz_291_;
      end
      if(_zz_279_)begin
        int_reg_array_3_53_real <= _zz_291_;
      end
      if(_zz_280_)begin
        int_reg_array_3_54_real <= _zz_291_;
      end
      if(_zz_281_)begin
        int_reg_array_3_55_real <= _zz_291_;
      end
      if(_zz_282_)begin
        int_reg_array_3_56_real <= _zz_291_;
      end
      if(_zz_283_)begin
        int_reg_array_3_57_real <= _zz_291_;
      end
      if(_zz_284_)begin
        int_reg_array_3_58_real <= _zz_291_;
      end
      if(_zz_285_)begin
        int_reg_array_3_59_real <= _zz_291_;
      end
      if(_zz_286_)begin
        int_reg_array_3_60_real <= _zz_291_;
      end
      if(_zz_287_)begin
        int_reg_array_3_61_real <= _zz_291_;
      end
      if(_zz_288_)begin
        int_reg_array_3_62_real <= _zz_291_;
      end
      if(_zz_289_)begin
        int_reg_array_3_63_real <= _zz_291_;
      end
      if(_zz_226_)begin
        int_reg_array_3_0_imag <= _zz_292_;
      end
      if(_zz_227_)begin
        int_reg_array_3_1_imag <= _zz_292_;
      end
      if(_zz_228_)begin
        int_reg_array_3_2_imag <= _zz_292_;
      end
      if(_zz_229_)begin
        int_reg_array_3_3_imag <= _zz_292_;
      end
      if(_zz_230_)begin
        int_reg_array_3_4_imag <= _zz_292_;
      end
      if(_zz_231_)begin
        int_reg_array_3_5_imag <= _zz_292_;
      end
      if(_zz_232_)begin
        int_reg_array_3_6_imag <= _zz_292_;
      end
      if(_zz_233_)begin
        int_reg_array_3_7_imag <= _zz_292_;
      end
      if(_zz_234_)begin
        int_reg_array_3_8_imag <= _zz_292_;
      end
      if(_zz_235_)begin
        int_reg_array_3_9_imag <= _zz_292_;
      end
      if(_zz_236_)begin
        int_reg_array_3_10_imag <= _zz_292_;
      end
      if(_zz_237_)begin
        int_reg_array_3_11_imag <= _zz_292_;
      end
      if(_zz_238_)begin
        int_reg_array_3_12_imag <= _zz_292_;
      end
      if(_zz_239_)begin
        int_reg_array_3_13_imag <= _zz_292_;
      end
      if(_zz_240_)begin
        int_reg_array_3_14_imag <= _zz_292_;
      end
      if(_zz_241_)begin
        int_reg_array_3_15_imag <= _zz_292_;
      end
      if(_zz_242_)begin
        int_reg_array_3_16_imag <= _zz_292_;
      end
      if(_zz_243_)begin
        int_reg_array_3_17_imag <= _zz_292_;
      end
      if(_zz_244_)begin
        int_reg_array_3_18_imag <= _zz_292_;
      end
      if(_zz_245_)begin
        int_reg_array_3_19_imag <= _zz_292_;
      end
      if(_zz_246_)begin
        int_reg_array_3_20_imag <= _zz_292_;
      end
      if(_zz_247_)begin
        int_reg_array_3_21_imag <= _zz_292_;
      end
      if(_zz_248_)begin
        int_reg_array_3_22_imag <= _zz_292_;
      end
      if(_zz_249_)begin
        int_reg_array_3_23_imag <= _zz_292_;
      end
      if(_zz_250_)begin
        int_reg_array_3_24_imag <= _zz_292_;
      end
      if(_zz_251_)begin
        int_reg_array_3_25_imag <= _zz_292_;
      end
      if(_zz_252_)begin
        int_reg_array_3_26_imag <= _zz_292_;
      end
      if(_zz_253_)begin
        int_reg_array_3_27_imag <= _zz_292_;
      end
      if(_zz_254_)begin
        int_reg_array_3_28_imag <= _zz_292_;
      end
      if(_zz_255_)begin
        int_reg_array_3_29_imag <= _zz_292_;
      end
      if(_zz_256_)begin
        int_reg_array_3_30_imag <= _zz_292_;
      end
      if(_zz_257_)begin
        int_reg_array_3_31_imag <= _zz_292_;
      end
      if(_zz_258_)begin
        int_reg_array_3_32_imag <= _zz_292_;
      end
      if(_zz_259_)begin
        int_reg_array_3_33_imag <= _zz_292_;
      end
      if(_zz_260_)begin
        int_reg_array_3_34_imag <= _zz_292_;
      end
      if(_zz_261_)begin
        int_reg_array_3_35_imag <= _zz_292_;
      end
      if(_zz_262_)begin
        int_reg_array_3_36_imag <= _zz_292_;
      end
      if(_zz_263_)begin
        int_reg_array_3_37_imag <= _zz_292_;
      end
      if(_zz_264_)begin
        int_reg_array_3_38_imag <= _zz_292_;
      end
      if(_zz_265_)begin
        int_reg_array_3_39_imag <= _zz_292_;
      end
      if(_zz_266_)begin
        int_reg_array_3_40_imag <= _zz_292_;
      end
      if(_zz_267_)begin
        int_reg_array_3_41_imag <= _zz_292_;
      end
      if(_zz_268_)begin
        int_reg_array_3_42_imag <= _zz_292_;
      end
      if(_zz_269_)begin
        int_reg_array_3_43_imag <= _zz_292_;
      end
      if(_zz_270_)begin
        int_reg_array_3_44_imag <= _zz_292_;
      end
      if(_zz_271_)begin
        int_reg_array_3_45_imag <= _zz_292_;
      end
      if(_zz_272_)begin
        int_reg_array_3_46_imag <= _zz_292_;
      end
      if(_zz_273_)begin
        int_reg_array_3_47_imag <= _zz_292_;
      end
      if(_zz_274_)begin
        int_reg_array_3_48_imag <= _zz_292_;
      end
      if(_zz_275_)begin
        int_reg_array_3_49_imag <= _zz_292_;
      end
      if(_zz_276_)begin
        int_reg_array_3_50_imag <= _zz_292_;
      end
      if(_zz_277_)begin
        int_reg_array_3_51_imag <= _zz_292_;
      end
      if(_zz_278_)begin
        int_reg_array_3_52_imag <= _zz_292_;
      end
      if(_zz_279_)begin
        int_reg_array_3_53_imag <= _zz_292_;
      end
      if(_zz_280_)begin
        int_reg_array_3_54_imag <= _zz_292_;
      end
      if(_zz_281_)begin
        int_reg_array_3_55_imag <= _zz_292_;
      end
      if(_zz_282_)begin
        int_reg_array_3_56_imag <= _zz_292_;
      end
      if(_zz_283_)begin
        int_reg_array_3_57_imag <= _zz_292_;
      end
      if(_zz_284_)begin
        int_reg_array_3_58_imag <= _zz_292_;
      end
      if(_zz_285_)begin
        int_reg_array_3_59_imag <= _zz_292_;
      end
      if(_zz_286_)begin
        int_reg_array_3_60_imag <= _zz_292_;
      end
      if(_zz_287_)begin
        int_reg_array_3_61_imag <= _zz_292_;
      end
      if(_zz_288_)begin
        int_reg_array_3_62_imag <= _zz_292_;
      end
      if(_zz_289_)begin
        int_reg_array_3_63_imag <= _zz_292_;
      end
      if(_zz_295_)begin
        int_reg_array_4_0_real <= _zz_360_;
      end
      if(_zz_296_)begin
        int_reg_array_4_1_real <= _zz_360_;
      end
      if(_zz_297_)begin
        int_reg_array_4_2_real <= _zz_360_;
      end
      if(_zz_298_)begin
        int_reg_array_4_3_real <= _zz_360_;
      end
      if(_zz_299_)begin
        int_reg_array_4_4_real <= _zz_360_;
      end
      if(_zz_300_)begin
        int_reg_array_4_5_real <= _zz_360_;
      end
      if(_zz_301_)begin
        int_reg_array_4_6_real <= _zz_360_;
      end
      if(_zz_302_)begin
        int_reg_array_4_7_real <= _zz_360_;
      end
      if(_zz_303_)begin
        int_reg_array_4_8_real <= _zz_360_;
      end
      if(_zz_304_)begin
        int_reg_array_4_9_real <= _zz_360_;
      end
      if(_zz_305_)begin
        int_reg_array_4_10_real <= _zz_360_;
      end
      if(_zz_306_)begin
        int_reg_array_4_11_real <= _zz_360_;
      end
      if(_zz_307_)begin
        int_reg_array_4_12_real <= _zz_360_;
      end
      if(_zz_308_)begin
        int_reg_array_4_13_real <= _zz_360_;
      end
      if(_zz_309_)begin
        int_reg_array_4_14_real <= _zz_360_;
      end
      if(_zz_310_)begin
        int_reg_array_4_15_real <= _zz_360_;
      end
      if(_zz_311_)begin
        int_reg_array_4_16_real <= _zz_360_;
      end
      if(_zz_312_)begin
        int_reg_array_4_17_real <= _zz_360_;
      end
      if(_zz_313_)begin
        int_reg_array_4_18_real <= _zz_360_;
      end
      if(_zz_314_)begin
        int_reg_array_4_19_real <= _zz_360_;
      end
      if(_zz_315_)begin
        int_reg_array_4_20_real <= _zz_360_;
      end
      if(_zz_316_)begin
        int_reg_array_4_21_real <= _zz_360_;
      end
      if(_zz_317_)begin
        int_reg_array_4_22_real <= _zz_360_;
      end
      if(_zz_318_)begin
        int_reg_array_4_23_real <= _zz_360_;
      end
      if(_zz_319_)begin
        int_reg_array_4_24_real <= _zz_360_;
      end
      if(_zz_320_)begin
        int_reg_array_4_25_real <= _zz_360_;
      end
      if(_zz_321_)begin
        int_reg_array_4_26_real <= _zz_360_;
      end
      if(_zz_322_)begin
        int_reg_array_4_27_real <= _zz_360_;
      end
      if(_zz_323_)begin
        int_reg_array_4_28_real <= _zz_360_;
      end
      if(_zz_324_)begin
        int_reg_array_4_29_real <= _zz_360_;
      end
      if(_zz_325_)begin
        int_reg_array_4_30_real <= _zz_360_;
      end
      if(_zz_326_)begin
        int_reg_array_4_31_real <= _zz_360_;
      end
      if(_zz_327_)begin
        int_reg_array_4_32_real <= _zz_360_;
      end
      if(_zz_328_)begin
        int_reg_array_4_33_real <= _zz_360_;
      end
      if(_zz_329_)begin
        int_reg_array_4_34_real <= _zz_360_;
      end
      if(_zz_330_)begin
        int_reg_array_4_35_real <= _zz_360_;
      end
      if(_zz_331_)begin
        int_reg_array_4_36_real <= _zz_360_;
      end
      if(_zz_332_)begin
        int_reg_array_4_37_real <= _zz_360_;
      end
      if(_zz_333_)begin
        int_reg_array_4_38_real <= _zz_360_;
      end
      if(_zz_334_)begin
        int_reg_array_4_39_real <= _zz_360_;
      end
      if(_zz_335_)begin
        int_reg_array_4_40_real <= _zz_360_;
      end
      if(_zz_336_)begin
        int_reg_array_4_41_real <= _zz_360_;
      end
      if(_zz_337_)begin
        int_reg_array_4_42_real <= _zz_360_;
      end
      if(_zz_338_)begin
        int_reg_array_4_43_real <= _zz_360_;
      end
      if(_zz_339_)begin
        int_reg_array_4_44_real <= _zz_360_;
      end
      if(_zz_340_)begin
        int_reg_array_4_45_real <= _zz_360_;
      end
      if(_zz_341_)begin
        int_reg_array_4_46_real <= _zz_360_;
      end
      if(_zz_342_)begin
        int_reg_array_4_47_real <= _zz_360_;
      end
      if(_zz_343_)begin
        int_reg_array_4_48_real <= _zz_360_;
      end
      if(_zz_344_)begin
        int_reg_array_4_49_real <= _zz_360_;
      end
      if(_zz_345_)begin
        int_reg_array_4_50_real <= _zz_360_;
      end
      if(_zz_346_)begin
        int_reg_array_4_51_real <= _zz_360_;
      end
      if(_zz_347_)begin
        int_reg_array_4_52_real <= _zz_360_;
      end
      if(_zz_348_)begin
        int_reg_array_4_53_real <= _zz_360_;
      end
      if(_zz_349_)begin
        int_reg_array_4_54_real <= _zz_360_;
      end
      if(_zz_350_)begin
        int_reg_array_4_55_real <= _zz_360_;
      end
      if(_zz_351_)begin
        int_reg_array_4_56_real <= _zz_360_;
      end
      if(_zz_352_)begin
        int_reg_array_4_57_real <= _zz_360_;
      end
      if(_zz_353_)begin
        int_reg_array_4_58_real <= _zz_360_;
      end
      if(_zz_354_)begin
        int_reg_array_4_59_real <= _zz_360_;
      end
      if(_zz_355_)begin
        int_reg_array_4_60_real <= _zz_360_;
      end
      if(_zz_356_)begin
        int_reg_array_4_61_real <= _zz_360_;
      end
      if(_zz_357_)begin
        int_reg_array_4_62_real <= _zz_360_;
      end
      if(_zz_358_)begin
        int_reg_array_4_63_real <= _zz_360_;
      end
      if(_zz_295_)begin
        int_reg_array_4_0_imag <= _zz_361_;
      end
      if(_zz_296_)begin
        int_reg_array_4_1_imag <= _zz_361_;
      end
      if(_zz_297_)begin
        int_reg_array_4_2_imag <= _zz_361_;
      end
      if(_zz_298_)begin
        int_reg_array_4_3_imag <= _zz_361_;
      end
      if(_zz_299_)begin
        int_reg_array_4_4_imag <= _zz_361_;
      end
      if(_zz_300_)begin
        int_reg_array_4_5_imag <= _zz_361_;
      end
      if(_zz_301_)begin
        int_reg_array_4_6_imag <= _zz_361_;
      end
      if(_zz_302_)begin
        int_reg_array_4_7_imag <= _zz_361_;
      end
      if(_zz_303_)begin
        int_reg_array_4_8_imag <= _zz_361_;
      end
      if(_zz_304_)begin
        int_reg_array_4_9_imag <= _zz_361_;
      end
      if(_zz_305_)begin
        int_reg_array_4_10_imag <= _zz_361_;
      end
      if(_zz_306_)begin
        int_reg_array_4_11_imag <= _zz_361_;
      end
      if(_zz_307_)begin
        int_reg_array_4_12_imag <= _zz_361_;
      end
      if(_zz_308_)begin
        int_reg_array_4_13_imag <= _zz_361_;
      end
      if(_zz_309_)begin
        int_reg_array_4_14_imag <= _zz_361_;
      end
      if(_zz_310_)begin
        int_reg_array_4_15_imag <= _zz_361_;
      end
      if(_zz_311_)begin
        int_reg_array_4_16_imag <= _zz_361_;
      end
      if(_zz_312_)begin
        int_reg_array_4_17_imag <= _zz_361_;
      end
      if(_zz_313_)begin
        int_reg_array_4_18_imag <= _zz_361_;
      end
      if(_zz_314_)begin
        int_reg_array_4_19_imag <= _zz_361_;
      end
      if(_zz_315_)begin
        int_reg_array_4_20_imag <= _zz_361_;
      end
      if(_zz_316_)begin
        int_reg_array_4_21_imag <= _zz_361_;
      end
      if(_zz_317_)begin
        int_reg_array_4_22_imag <= _zz_361_;
      end
      if(_zz_318_)begin
        int_reg_array_4_23_imag <= _zz_361_;
      end
      if(_zz_319_)begin
        int_reg_array_4_24_imag <= _zz_361_;
      end
      if(_zz_320_)begin
        int_reg_array_4_25_imag <= _zz_361_;
      end
      if(_zz_321_)begin
        int_reg_array_4_26_imag <= _zz_361_;
      end
      if(_zz_322_)begin
        int_reg_array_4_27_imag <= _zz_361_;
      end
      if(_zz_323_)begin
        int_reg_array_4_28_imag <= _zz_361_;
      end
      if(_zz_324_)begin
        int_reg_array_4_29_imag <= _zz_361_;
      end
      if(_zz_325_)begin
        int_reg_array_4_30_imag <= _zz_361_;
      end
      if(_zz_326_)begin
        int_reg_array_4_31_imag <= _zz_361_;
      end
      if(_zz_327_)begin
        int_reg_array_4_32_imag <= _zz_361_;
      end
      if(_zz_328_)begin
        int_reg_array_4_33_imag <= _zz_361_;
      end
      if(_zz_329_)begin
        int_reg_array_4_34_imag <= _zz_361_;
      end
      if(_zz_330_)begin
        int_reg_array_4_35_imag <= _zz_361_;
      end
      if(_zz_331_)begin
        int_reg_array_4_36_imag <= _zz_361_;
      end
      if(_zz_332_)begin
        int_reg_array_4_37_imag <= _zz_361_;
      end
      if(_zz_333_)begin
        int_reg_array_4_38_imag <= _zz_361_;
      end
      if(_zz_334_)begin
        int_reg_array_4_39_imag <= _zz_361_;
      end
      if(_zz_335_)begin
        int_reg_array_4_40_imag <= _zz_361_;
      end
      if(_zz_336_)begin
        int_reg_array_4_41_imag <= _zz_361_;
      end
      if(_zz_337_)begin
        int_reg_array_4_42_imag <= _zz_361_;
      end
      if(_zz_338_)begin
        int_reg_array_4_43_imag <= _zz_361_;
      end
      if(_zz_339_)begin
        int_reg_array_4_44_imag <= _zz_361_;
      end
      if(_zz_340_)begin
        int_reg_array_4_45_imag <= _zz_361_;
      end
      if(_zz_341_)begin
        int_reg_array_4_46_imag <= _zz_361_;
      end
      if(_zz_342_)begin
        int_reg_array_4_47_imag <= _zz_361_;
      end
      if(_zz_343_)begin
        int_reg_array_4_48_imag <= _zz_361_;
      end
      if(_zz_344_)begin
        int_reg_array_4_49_imag <= _zz_361_;
      end
      if(_zz_345_)begin
        int_reg_array_4_50_imag <= _zz_361_;
      end
      if(_zz_346_)begin
        int_reg_array_4_51_imag <= _zz_361_;
      end
      if(_zz_347_)begin
        int_reg_array_4_52_imag <= _zz_361_;
      end
      if(_zz_348_)begin
        int_reg_array_4_53_imag <= _zz_361_;
      end
      if(_zz_349_)begin
        int_reg_array_4_54_imag <= _zz_361_;
      end
      if(_zz_350_)begin
        int_reg_array_4_55_imag <= _zz_361_;
      end
      if(_zz_351_)begin
        int_reg_array_4_56_imag <= _zz_361_;
      end
      if(_zz_352_)begin
        int_reg_array_4_57_imag <= _zz_361_;
      end
      if(_zz_353_)begin
        int_reg_array_4_58_imag <= _zz_361_;
      end
      if(_zz_354_)begin
        int_reg_array_4_59_imag <= _zz_361_;
      end
      if(_zz_355_)begin
        int_reg_array_4_60_imag <= _zz_361_;
      end
      if(_zz_356_)begin
        int_reg_array_4_61_imag <= _zz_361_;
      end
      if(_zz_357_)begin
        int_reg_array_4_62_imag <= _zz_361_;
      end
      if(_zz_358_)begin
        int_reg_array_4_63_imag <= _zz_361_;
      end
      if(_zz_364_)begin
        int_reg_array_5_0_real <= _zz_429_;
      end
      if(_zz_365_)begin
        int_reg_array_5_1_real <= _zz_429_;
      end
      if(_zz_366_)begin
        int_reg_array_5_2_real <= _zz_429_;
      end
      if(_zz_367_)begin
        int_reg_array_5_3_real <= _zz_429_;
      end
      if(_zz_368_)begin
        int_reg_array_5_4_real <= _zz_429_;
      end
      if(_zz_369_)begin
        int_reg_array_5_5_real <= _zz_429_;
      end
      if(_zz_370_)begin
        int_reg_array_5_6_real <= _zz_429_;
      end
      if(_zz_371_)begin
        int_reg_array_5_7_real <= _zz_429_;
      end
      if(_zz_372_)begin
        int_reg_array_5_8_real <= _zz_429_;
      end
      if(_zz_373_)begin
        int_reg_array_5_9_real <= _zz_429_;
      end
      if(_zz_374_)begin
        int_reg_array_5_10_real <= _zz_429_;
      end
      if(_zz_375_)begin
        int_reg_array_5_11_real <= _zz_429_;
      end
      if(_zz_376_)begin
        int_reg_array_5_12_real <= _zz_429_;
      end
      if(_zz_377_)begin
        int_reg_array_5_13_real <= _zz_429_;
      end
      if(_zz_378_)begin
        int_reg_array_5_14_real <= _zz_429_;
      end
      if(_zz_379_)begin
        int_reg_array_5_15_real <= _zz_429_;
      end
      if(_zz_380_)begin
        int_reg_array_5_16_real <= _zz_429_;
      end
      if(_zz_381_)begin
        int_reg_array_5_17_real <= _zz_429_;
      end
      if(_zz_382_)begin
        int_reg_array_5_18_real <= _zz_429_;
      end
      if(_zz_383_)begin
        int_reg_array_5_19_real <= _zz_429_;
      end
      if(_zz_384_)begin
        int_reg_array_5_20_real <= _zz_429_;
      end
      if(_zz_385_)begin
        int_reg_array_5_21_real <= _zz_429_;
      end
      if(_zz_386_)begin
        int_reg_array_5_22_real <= _zz_429_;
      end
      if(_zz_387_)begin
        int_reg_array_5_23_real <= _zz_429_;
      end
      if(_zz_388_)begin
        int_reg_array_5_24_real <= _zz_429_;
      end
      if(_zz_389_)begin
        int_reg_array_5_25_real <= _zz_429_;
      end
      if(_zz_390_)begin
        int_reg_array_5_26_real <= _zz_429_;
      end
      if(_zz_391_)begin
        int_reg_array_5_27_real <= _zz_429_;
      end
      if(_zz_392_)begin
        int_reg_array_5_28_real <= _zz_429_;
      end
      if(_zz_393_)begin
        int_reg_array_5_29_real <= _zz_429_;
      end
      if(_zz_394_)begin
        int_reg_array_5_30_real <= _zz_429_;
      end
      if(_zz_395_)begin
        int_reg_array_5_31_real <= _zz_429_;
      end
      if(_zz_396_)begin
        int_reg_array_5_32_real <= _zz_429_;
      end
      if(_zz_397_)begin
        int_reg_array_5_33_real <= _zz_429_;
      end
      if(_zz_398_)begin
        int_reg_array_5_34_real <= _zz_429_;
      end
      if(_zz_399_)begin
        int_reg_array_5_35_real <= _zz_429_;
      end
      if(_zz_400_)begin
        int_reg_array_5_36_real <= _zz_429_;
      end
      if(_zz_401_)begin
        int_reg_array_5_37_real <= _zz_429_;
      end
      if(_zz_402_)begin
        int_reg_array_5_38_real <= _zz_429_;
      end
      if(_zz_403_)begin
        int_reg_array_5_39_real <= _zz_429_;
      end
      if(_zz_404_)begin
        int_reg_array_5_40_real <= _zz_429_;
      end
      if(_zz_405_)begin
        int_reg_array_5_41_real <= _zz_429_;
      end
      if(_zz_406_)begin
        int_reg_array_5_42_real <= _zz_429_;
      end
      if(_zz_407_)begin
        int_reg_array_5_43_real <= _zz_429_;
      end
      if(_zz_408_)begin
        int_reg_array_5_44_real <= _zz_429_;
      end
      if(_zz_409_)begin
        int_reg_array_5_45_real <= _zz_429_;
      end
      if(_zz_410_)begin
        int_reg_array_5_46_real <= _zz_429_;
      end
      if(_zz_411_)begin
        int_reg_array_5_47_real <= _zz_429_;
      end
      if(_zz_412_)begin
        int_reg_array_5_48_real <= _zz_429_;
      end
      if(_zz_413_)begin
        int_reg_array_5_49_real <= _zz_429_;
      end
      if(_zz_414_)begin
        int_reg_array_5_50_real <= _zz_429_;
      end
      if(_zz_415_)begin
        int_reg_array_5_51_real <= _zz_429_;
      end
      if(_zz_416_)begin
        int_reg_array_5_52_real <= _zz_429_;
      end
      if(_zz_417_)begin
        int_reg_array_5_53_real <= _zz_429_;
      end
      if(_zz_418_)begin
        int_reg_array_5_54_real <= _zz_429_;
      end
      if(_zz_419_)begin
        int_reg_array_5_55_real <= _zz_429_;
      end
      if(_zz_420_)begin
        int_reg_array_5_56_real <= _zz_429_;
      end
      if(_zz_421_)begin
        int_reg_array_5_57_real <= _zz_429_;
      end
      if(_zz_422_)begin
        int_reg_array_5_58_real <= _zz_429_;
      end
      if(_zz_423_)begin
        int_reg_array_5_59_real <= _zz_429_;
      end
      if(_zz_424_)begin
        int_reg_array_5_60_real <= _zz_429_;
      end
      if(_zz_425_)begin
        int_reg_array_5_61_real <= _zz_429_;
      end
      if(_zz_426_)begin
        int_reg_array_5_62_real <= _zz_429_;
      end
      if(_zz_427_)begin
        int_reg_array_5_63_real <= _zz_429_;
      end
      if(_zz_364_)begin
        int_reg_array_5_0_imag <= _zz_430_;
      end
      if(_zz_365_)begin
        int_reg_array_5_1_imag <= _zz_430_;
      end
      if(_zz_366_)begin
        int_reg_array_5_2_imag <= _zz_430_;
      end
      if(_zz_367_)begin
        int_reg_array_5_3_imag <= _zz_430_;
      end
      if(_zz_368_)begin
        int_reg_array_5_4_imag <= _zz_430_;
      end
      if(_zz_369_)begin
        int_reg_array_5_5_imag <= _zz_430_;
      end
      if(_zz_370_)begin
        int_reg_array_5_6_imag <= _zz_430_;
      end
      if(_zz_371_)begin
        int_reg_array_5_7_imag <= _zz_430_;
      end
      if(_zz_372_)begin
        int_reg_array_5_8_imag <= _zz_430_;
      end
      if(_zz_373_)begin
        int_reg_array_5_9_imag <= _zz_430_;
      end
      if(_zz_374_)begin
        int_reg_array_5_10_imag <= _zz_430_;
      end
      if(_zz_375_)begin
        int_reg_array_5_11_imag <= _zz_430_;
      end
      if(_zz_376_)begin
        int_reg_array_5_12_imag <= _zz_430_;
      end
      if(_zz_377_)begin
        int_reg_array_5_13_imag <= _zz_430_;
      end
      if(_zz_378_)begin
        int_reg_array_5_14_imag <= _zz_430_;
      end
      if(_zz_379_)begin
        int_reg_array_5_15_imag <= _zz_430_;
      end
      if(_zz_380_)begin
        int_reg_array_5_16_imag <= _zz_430_;
      end
      if(_zz_381_)begin
        int_reg_array_5_17_imag <= _zz_430_;
      end
      if(_zz_382_)begin
        int_reg_array_5_18_imag <= _zz_430_;
      end
      if(_zz_383_)begin
        int_reg_array_5_19_imag <= _zz_430_;
      end
      if(_zz_384_)begin
        int_reg_array_5_20_imag <= _zz_430_;
      end
      if(_zz_385_)begin
        int_reg_array_5_21_imag <= _zz_430_;
      end
      if(_zz_386_)begin
        int_reg_array_5_22_imag <= _zz_430_;
      end
      if(_zz_387_)begin
        int_reg_array_5_23_imag <= _zz_430_;
      end
      if(_zz_388_)begin
        int_reg_array_5_24_imag <= _zz_430_;
      end
      if(_zz_389_)begin
        int_reg_array_5_25_imag <= _zz_430_;
      end
      if(_zz_390_)begin
        int_reg_array_5_26_imag <= _zz_430_;
      end
      if(_zz_391_)begin
        int_reg_array_5_27_imag <= _zz_430_;
      end
      if(_zz_392_)begin
        int_reg_array_5_28_imag <= _zz_430_;
      end
      if(_zz_393_)begin
        int_reg_array_5_29_imag <= _zz_430_;
      end
      if(_zz_394_)begin
        int_reg_array_5_30_imag <= _zz_430_;
      end
      if(_zz_395_)begin
        int_reg_array_5_31_imag <= _zz_430_;
      end
      if(_zz_396_)begin
        int_reg_array_5_32_imag <= _zz_430_;
      end
      if(_zz_397_)begin
        int_reg_array_5_33_imag <= _zz_430_;
      end
      if(_zz_398_)begin
        int_reg_array_5_34_imag <= _zz_430_;
      end
      if(_zz_399_)begin
        int_reg_array_5_35_imag <= _zz_430_;
      end
      if(_zz_400_)begin
        int_reg_array_5_36_imag <= _zz_430_;
      end
      if(_zz_401_)begin
        int_reg_array_5_37_imag <= _zz_430_;
      end
      if(_zz_402_)begin
        int_reg_array_5_38_imag <= _zz_430_;
      end
      if(_zz_403_)begin
        int_reg_array_5_39_imag <= _zz_430_;
      end
      if(_zz_404_)begin
        int_reg_array_5_40_imag <= _zz_430_;
      end
      if(_zz_405_)begin
        int_reg_array_5_41_imag <= _zz_430_;
      end
      if(_zz_406_)begin
        int_reg_array_5_42_imag <= _zz_430_;
      end
      if(_zz_407_)begin
        int_reg_array_5_43_imag <= _zz_430_;
      end
      if(_zz_408_)begin
        int_reg_array_5_44_imag <= _zz_430_;
      end
      if(_zz_409_)begin
        int_reg_array_5_45_imag <= _zz_430_;
      end
      if(_zz_410_)begin
        int_reg_array_5_46_imag <= _zz_430_;
      end
      if(_zz_411_)begin
        int_reg_array_5_47_imag <= _zz_430_;
      end
      if(_zz_412_)begin
        int_reg_array_5_48_imag <= _zz_430_;
      end
      if(_zz_413_)begin
        int_reg_array_5_49_imag <= _zz_430_;
      end
      if(_zz_414_)begin
        int_reg_array_5_50_imag <= _zz_430_;
      end
      if(_zz_415_)begin
        int_reg_array_5_51_imag <= _zz_430_;
      end
      if(_zz_416_)begin
        int_reg_array_5_52_imag <= _zz_430_;
      end
      if(_zz_417_)begin
        int_reg_array_5_53_imag <= _zz_430_;
      end
      if(_zz_418_)begin
        int_reg_array_5_54_imag <= _zz_430_;
      end
      if(_zz_419_)begin
        int_reg_array_5_55_imag <= _zz_430_;
      end
      if(_zz_420_)begin
        int_reg_array_5_56_imag <= _zz_430_;
      end
      if(_zz_421_)begin
        int_reg_array_5_57_imag <= _zz_430_;
      end
      if(_zz_422_)begin
        int_reg_array_5_58_imag <= _zz_430_;
      end
      if(_zz_423_)begin
        int_reg_array_5_59_imag <= _zz_430_;
      end
      if(_zz_424_)begin
        int_reg_array_5_60_imag <= _zz_430_;
      end
      if(_zz_425_)begin
        int_reg_array_5_61_imag <= _zz_430_;
      end
      if(_zz_426_)begin
        int_reg_array_5_62_imag <= _zz_430_;
      end
      if(_zz_427_)begin
        int_reg_array_5_63_imag <= _zz_430_;
      end
      if(_zz_433_)begin
        int_reg_array_6_0_real <= _zz_498_;
      end
      if(_zz_434_)begin
        int_reg_array_6_1_real <= _zz_498_;
      end
      if(_zz_435_)begin
        int_reg_array_6_2_real <= _zz_498_;
      end
      if(_zz_436_)begin
        int_reg_array_6_3_real <= _zz_498_;
      end
      if(_zz_437_)begin
        int_reg_array_6_4_real <= _zz_498_;
      end
      if(_zz_438_)begin
        int_reg_array_6_5_real <= _zz_498_;
      end
      if(_zz_439_)begin
        int_reg_array_6_6_real <= _zz_498_;
      end
      if(_zz_440_)begin
        int_reg_array_6_7_real <= _zz_498_;
      end
      if(_zz_441_)begin
        int_reg_array_6_8_real <= _zz_498_;
      end
      if(_zz_442_)begin
        int_reg_array_6_9_real <= _zz_498_;
      end
      if(_zz_443_)begin
        int_reg_array_6_10_real <= _zz_498_;
      end
      if(_zz_444_)begin
        int_reg_array_6_11_real <= _zz_498_;
      end
      if(_zz_445_)begin
        int_reg_array_6_12_real <= _zz_498_;
      end
      if(_zz_446_)begin
        int_reg_array_6_13_real <= _zz_498_;
      end
      if(_zz_447_)begin
        int_reg_array_6_14_real <= _zz_498_;
      end
      if(_zz_448_)begin
        int_reg_array_6_15_real <= _zz_498_;
      end
      if(_zz_449_)begin
        int_reg_array_6_16_real <= _zz_498_;
      end
      if(_zz_450_)begin
        int_reg_array_6_17_real <= _zz_498_;
      end
      if(_zz_451_)begin
        int_reg_array_6_18_real <= _zz_498_;
      end
      if(_zz_452_)begin
        int_reg_array_6_19_real <= _zz_498_;
      end
      if(_zz_453_)begin
        int_reg_array_6_20_real <= _zz_498_;
      end
      if(_zz_454_)begin
        int_reg_array_6_21_real <= _zz_498_;
      end
      if(_zz_455_)begin
        int_reg_array_6_22_real <= _zz_498_;
      end
      if(_zz_456_)begin
        int_reg_array_6_23_real <= _zz_498_;
      end
      if(_zz_457_)begin
        int_reg_array_6_24_real <= _zz_498_;
      end
      if(_zz_458_)begin
        int_reg_array_6_25_real <= _zz_498_;
      end
      if(_zz_459_)begin
        int_reg_array_6_26_real <= _zz_498_;
      end
      if(_zz_460_)begin
        int_reg_array_6_27_real <= _zz_498_;
      end
      if(_zz_461_)begin
        int_reg_array_6_28_real <= _zz_498_;
      end
      if(_zz_462_)begin
        int_reg_array_6_29_real <= _zz_498_;
      end
      if(_zz_463_)begin
        int_reg_array_6_30_real <= _zz_498_;
      end
      if(_zz_464_)begin
        int_reg_array_6_31_real <= _zz_498_;
      end
      if(_zz_465_)begin
        int_reg_array_6_32_real <= _zz_498_;
      end
      if(_zz_466_)begin
        int_reg_array_6_33_real <= _zz_498_;
      end
      if(_zz_467_)begin
        int_reg_array_6_34_real <= _zz_498_;
      end
      if(_zz_468_)begin
        int_reg_array_6_35_real <= _zz_498_;
      end
      if(_zz_469_)begin
        int_reg_array_6_36_real <= _zz_498_;
      end
      if(_zz_470_)begin
        int_reg_array_6_37_real <= _zz_498_;
      end
      if(_zz_471_)begin
        int_reg_array_6_38_real <= _zz_498_;
      end
      if(_zz_472_)begin
        int_reg_array_6_39_real <= _zz_498_;
      end
      if(_zz_473_)begin
        int_reg_array_6_40_real <= _zz_498_;
      end
      if(_zz_474_)begin
        int_reg_array_6_41_real <= _zz_498_;
      end
      if(_zz_475_)begin
        int_reg_array_6_42_real <= _zz_498_;
      end
      if(_zz_476_)begin
        int_reg_array_6_43_real <= _zz_498_;
      end
      if(_zz_477_)begin
        int_reg_array_6_44_real <= _zz_498_;
      end
      if(_zz_478_)begin
        int_reg_array_6_45_real <= _zz_498_;
      end
      if(_zz_479_)begin
        int_reg_array_6_46_real <= _zz_498_;
      end
      if(_zz_480_)begin
        int_reg_array_6_47_real <= _zz_498_;
      end
      if(_zz_481_)begin
        int_reg_array_6_48_real <= _zz_498_;
      end
      if(_zz_482_)begin
        int_reg_array_6_49_real <= _zz_498_;
      end
      if(_zz_483_)begin
        int_reg_array_6_50_real <= _zz_498_;
      end
      if(_zz_484_)begin
        int_reg_array_6_51_real <= _zz_498_;
      end
      if(_zz_485_)begin
        int_reg_array_6_52_real <= _zz_498_;
      end
      if(_zz_486_)begin
        int_reg_array_6_53_real <= _zz_498_;
      end
      if(_zz_487_)begin
        int_reg_array_6_54_real <= _zz_498_;
      end
      if(_zz_488_)begin
        int_reg_array_6_55_real <= _zz_498_;
      end
      if(_zz_489_)begin
        int_reg_array_6_56_real <= _zz_498_;
      end
      if(_zz_490_)begin
        int_reg_array_6_57_real <= _zz_498_;
      end
      if(_zz_491_)begin
        int_reg_array_6_58_real <= _zz_498_;
      end
      if(_zz_492_)begin
        int_reg_array_6_59_real <= _zz_498_;
      end
      if(_zz_493_)begin
        int_reg_array_6_60_real <= _zz_498_;
      end
      if(_zz_494_)begin
        int_reg_array_6_61_real <= _zz_498_;
      end
      if(_zz_495_)begin
        int_reg_array_6_62_real <= _zz_498_;
      end
      if(_zz_496_)begin
        int_reg_array_6_63_real <= _zz_498_;
      end
      if(_zz_433_)begin
        int_reg_array_6_0_imag <= _zz_499_;
      end
      if(_zz_434_)begin
        int_reg_array_6_1_imag <= _zz_499_;
      end
      if(_zz_435_)begin
        int_reg_array_6_2_imag <= _zz_499_;
      end
      if(_zz_436_)begin
        int_reg_array_6_3_imag <= _zz_499_;
      end
      if(_zz_437_)begin
        int_reg_array_6_4_imag <= _zz_499_;
      end
      if(_zz_438_)begin
        int_reg_array_6_5_imag <= _zz_499_;
      end
      if(_zz_439_)begin
        int_reg_array_6_6_imag <= _zz_499_;
      end
      if(_zz_440_)begin
        int_reg_array_6_7_imag <= _zz_499_;
      end
      if(_zz_441_)begin
        int_reg_array_6_8_imag <= _zz_499_;
      end
      if(_zz_442_)begin
        int_reg_array_6_9_imag <= _zz_499_;
      end
      if(_zz_443_)begin
        int_reg_array_6_10_imag <= _zz_499_;
      end
      if(_zz_444_)begin
        int_reg_array_6_11_imag <= _zz_499_;
      end
      if(_zz_445_)begin
        int_reg_array_6_12_imag <= _zz_499_;
      end
      if(_zz_446_)begin
        int_reg_array_6_13_imag <= _zz_499_;
      end
      if(_zz_447_)begin
        int_reg_array_6_14_imag <= _zz_499_;
      end
      if(_zz_448_)begin
        int_reg_array_6_15_imag <= _zz_499_;
      end
      if(_zz_449_)begin
        int_reg_array_6_16_imag <= _zz_499_;
      end
      if(_zz_450_)begin
        int_reg_array_6_17_imag <= _zz_499_;
      end
      if(_zz_451_)begin
        int_reg_array_6_18_imag <= _zz_499_;
      end
      if(_zz_452_)begin
        int_reg_array_6_19_imag <= _zz_499_;
      end
      if(_zz_453_)begin
        int_reg_array_6_20_imag <= _zz_499_;
      end
      if(_zz_454_)begin
        int_reg_array_6_21_imag <= _zz_499_;
      end
      if(_zz_455_)begin
        int_reg_array_6_22_imag <= _zz_499_;
      end
      if(_zz_456_)begin
        int_reg_array_6_23_imag <= _zz_499_;
      end
      if(_zz_457_)begin
        int_reg_array_6_24_imag <= _zz_499_;
      end
      if(_zz_458_)begin
        int_reg_array_6_25_imag <= _zz_499_;
      end
      if(_zz_459_)begin
        int_reg_array_6_26_imag <= _zz_499_;
      end
      if(_zz_460_)begin
        int_reg_array_6_27_imag <= _zz_499_;
      end
      if(_zz_461_)begin
        int_reg_array_6_28_imag <= _zz_499_;
      end
      if(_zz_462_)begin
        int_reg_array_6_29_imag <= _zz_499_;
      end
      if(_zz_463_)begin
        int_reg_array_6_30_imag <= _zz_499_;
      end
      if(_zz_464_)begin
        int_reg_array_6_31_imag <= _zz_499_;
      end
      if(_zz_465_)begin
        int_reg_array_6_32_imag <= _zz_499_;
      end
      if(_zz_466_)begin
        int_reg_array_6_33_imag <= _zz_499_;
      end
      if(_zz_467_)begin
        int_reg_array_6_34_imag <= _zz_499_;
      end
      if(_zz_468_)begin
        int_reg_array_6_35_imag <= _zz_499_;
      end
      if(_zz_469_)begin
        int_reg_array_6_36_imag <= _zz_499_;
      end
      if(_zz_470_)begin
        int_reg_array_6_37_imag <= _zz_499_;
      end
      if(_zz_471_)begin
        int_reg_array_6_38_imag <= _zz_499_;
      end
      if(_zz_472_)begin
        int_reg_array_6_39_imag <= _zz_499_;
      end
      if(_zz_473_)begin
        int_reg_array_6_40_imag <= _zz_499_;
      end
      if(_zz_474_)begin
        int_reg_array_6_41_imag <= _zz_499_;
      end
      if(_zz_475_)begin
        int_reg_array_6_42_imag <= _zz_499_;
      end
      if(_zz_476_)begin
        int_reg_array_6_43_imag <= _zz_499_;
      end
      if(_zz_477_)begin
        int_reg_array_6_44_imag <= _zz_499_;
      end
      if(_zz_478_)begin
        int_reg_array_6_45_imag <= _zz_499_;
      end
      if(_zz_479_)begin
        int_reg_array_6_46_imag <= _zz_499_;
      end
      if(_zz_480_)begin
        int_reg_array_6_47_imag <= _zz_499_;
      end
      if(_zz_481_)begin
        int_reg_array_6_48_imag <= _zz_499_;
      end
      if(_zz_482_)begin
        int_reg_array_6_49_imag <= _zz_499_;
      end
      if(_zz_483_)begin
        int_reg_array_6_50_imag <= _zz_499_;
      end
      if(_zz_484_)begin
        int_reg_array_6_51_imag <= _zz_499_;
      end
      if(_zz_485_)begin
        int_reg_array_6_52_imag <= _zz_499_;
      end
      if(_zz_486_)begin
        int_reg_array_6_53_imag <= _zz_499_;
      end
      if(_zz_487_)begin
        int_reg_array_6_54_imag <= _zz_499_;
      end
      if(_zz_488_)begin
        int_reg_array_6_55_imag <= _zz_499_;
      end
      if(_zz_489_)begin
        int_reg_array_6_56_imag <= _zz_499_;
      end
      if(_zz_490_)begin
        int_reg_array_6_57_imag <= _zz_499_;
      end
      if(_zz_491_)begin
        int_reg_array_6_58_imag <= _zz_499_;
      end
      if(_zz_492_)begin
        int_reg_array_6_59_imag <= _zz_499_;
      end
      if(_zz_493_)begin
        int_reg_array_6_60_imag <= _zz_499_;
      end
      if(_zz_494_)begin
        int_reg_array_6_61_imag <= _zz_499_;
      end
      if(_zz_495_)begin
        int_reg_array_6_62_imag <= _zz_499_;
      end
      if(_zz_496_)begin
        int_reg_array_6_63_imag <= _zz_499_;
      end
      if(_zz_502_)begin
        int_reg_array_7_0_real <= _zz_567_;
      end
      if(_zz_503_)begin
        int_reg_array_7_1_real <= _zz_567_;
      end
      if(_zz_504_)begin
        int_reg_array_7_2_real <= _zz_567_;
      end
      if(_zz_505_)begin
        int_reg_array_7_3_real <= _zz_567_;
      end
      if(_zz_506_)begin
        int_reg_array_7_4_real <= _zz_567_;
      end
      if(_zz_507_)begin
        int_reg_array_7_5_real <= _zz_567_;
      end
      if(_zz_508_)begin
        int_reg_array_7_6_real <= _zz_567_;
      end
      if(_zz_509_)begin
        int_reg_array_7_7_real <= _zz_567_;
      end
      if(_zz_510_)begin
        int_reg_array_7_8_real <= _zz_567_;
      end
      if(_zz_511_)begin
        int_reg_array_7_9_real <= _zz_567_;
      end
      if(_zz_512_)begin
        int_reg_array_7_10_real <= _zz_567_;
      end
      if(_zz_513_)begin
        int_reg_array_7_11_real <= _zz_567_;
      end
      if(_zz_514_)begin
        int_reg_array_7_12_real <= _zz_567_;
      end
      if(_zz_515_)begin
        int_reg_array_7_13_real <= _zz_567_;
      end
      if(_zz_516_)begin
        int_reg_array_7_14_real <= _zz_567_;
      end
      if(_zz_517_)begin
        int_reg_array_7_15_real <= _zz_567_;
      end
      if(_zz_518_)begin
        int_reg_array_7_16_real <= _zz_567_;
      end
      if(_zz_519_)begin
        int_reg_array_7_17_real <= _zz_567_;
      end
      if(_zz_520_)begin
        int_reg_array_7_18_real <= _zz_567_;
      end
      if(_zz_521_)begin
        int_reg_array_7_19_real <= _zz_567_;
      end
      if(_zz_522_)begin
        int_reg_array_7_20_real <= _zz_567_;
      end
      if(_zz_523_)begin
        int_reg_array_7_21_real <= _zz_567_;
      end
      if(_zz_524_)begin
        int_reg_array_7_22_real <= _zz_567_;
      end
      if(_zz_525_)begin
        int_reg_array_7_23_real <= _zz_567_;
      end
      if(_zz_526_)begin
        int_reg_array_7_24_real <= _zz_567_;
      end
      if(_zz_527_)begin
        int_reg_array_7_25_real <= _zz_567_;
      end
      if(_zz_528_)begin
        int_reg_array_7_26_real <= _zz_567_;
      end
      if(_zz_529_)begin
        int_reg_array_7_27_real <= _zz_567_;
      end
      if(_zz_530_)begin
        int_reg_array_7_28_real <= _zz_567_;
      end
      if(_zz_531_)begin
        int_reg_array_7_29_real <= _zz_567_;
      end
      if(_zz_532_)begin
        int_reg_array_7_30_real <= _zz_567_;
      end
      if(_zz_533_)begin
        int_reg_array_7_31_real <= _zz_567_;
      end
      if(_zz_534_)begin
        int_reg_array_7_32_real <= _zz_567_;
      end
      if(_zz_535_)begin
        int_reg_array_7_33_real <= _zz_567_;
      end
      if(_zz_536_)begin
        int_reg_array_7_34_real <= _zz_567_;
      end
      if(_zz_537_)begin
        int_reg_array_7_35_real <= _zz_567_;
      end
      if(_zz_538_)begin
        int_reg_array_7_36_real <= _zz_567_;
      end
      if(_zz_539_)begin
        int_reg_array_7_37_real <= _zz_567_;
      end
      if(_zz_540_)begin
        int_reg_array_7_38_real <= _zz_567_;
      end
      if(_zz_541_)begin
        int_reg_array_7_39_real <= _zz_567_;
      end
      if(_zz_542_)begin
        int_reg_array_7_40_real <= _zz_567_;
      end
      if(_zz_543_)begin
        int_reg_array_7_41_real <= _zz_567_;
      end
      if(_zz_544_)begin
        int_reg_array_7_42_real <= _zz_567_;
      end
      if(_zz_545_)begin
        int_reg_array_7_43_real <= _zz_567_;
      end
      if(_zz_546_)begin
        int_reg_array_7_44_real <= _zz_567_;
      end
      if(_zz_547_)begin
        int_reg_array_7_45_real <= _zz_567_;
      end
      if(_zz_548_)begin
        int_reg_array_7_46_real <= _zz_567_;
      end
      if(_zz_549_)begin
        int_reg_array_7_47_real <= _zz_567_;
      end
      if(_zz_550_)begin
        int_reg_array_7_48_real <= _zz_567_;
      end
      if(_zz_551_)begin
        int_reg_array_7_49_real <= _zz_567_;
      end
      if(_zz_552_)begin
        int_reg_array_7_50_real <= _zz_567_;
      end
      if(_zz_553_)begin
        int_reg_array_7_51_real <= _zz_567_;
      end
      if(_zz_554_)begin
        int_reg_array_7_52_real <= _zz_567_;
      end
      if(_zz_555_)begin
        int_reg_array_7_53_real <= _zz_567_;
      end
      if(_zz_556_)begin
        int_reg_array_7_54_real <= _zz_567_;
      end
      if(_zz_557_)begin
        int_reg_array_7_55_real <= _zz_567_;
      end
      if(_zz_558_)begin
        int_reg_array_7_56_real <= _zz_567_;
      end
      if(_zz_559_)begin
        int_reg_array_7_57_real <= _zz_567_;
      end
      if(_zz_560_)begin
        int_reg_array_7_58_real <= _zz_567_;
      end
      if(_zz_561_)begin
        int_reg_array_7_59_real <= _zz_567_;
      end
      if(_zz_562_)begin
        int_reg_array_7_60_real <= _zz_567_;
      end
      if(_zz_563_)begin
        int_reg_array_7_61_real <= _zz_567_;
      end
      if(_zz_564_)begin
        int_reg_array_7_62_real <= _zz_567_;
      end
      if(_zz_565_)begin
        int_reg_array_7_63_real <= _zz_567_;
      end
      if(_zz_502_)begin
        int_reg_array_7_0_imag <= _zz_568_;
      end
      if(_zz_503_)begin
        int_reg_array_7_1_imag <= _zz_568_;
      end
      if(_zz_504_)begin
        int_reg_array_7_2_imag <= _zz_568_;
      end
      if(_zz_505_)begin
        int_reg_array_7_3_imag <= _zz_568_;
      end
      if(_zz_506_)begin
        int_reg_array_7_4_imag <= _zz_568_;
      end
      if(_zz_507_)begin
        int_reg_array_7_5_imag <= _zz_568_;
      end
      if(_zz_508_)begin
        int_reg_array_7_6_imag <= _zz_568_;
      end
      if(_zz_509_)begin
        int_reg_array_7_7_imag <= _zz_568_;
      end
      if(_zz_510_)begin
        int_reg_array_7_8_imag <= _zz_568_;
      end
      if(_zz_511_)begin
        int_reg_array_7_9_imag <= _zz_568_;
      end
      if(_zz_512_)begin
        int_reg_array_7_10_imag <= _zz_568_;
      end
      if(_zz_513_)begin
        int_reg_array_7_11_imag <= _zz_568_;
      end
      if(_zz_514_)begin
        int_reg_array_7_12_imag <= _zz_568_;
      end
      if(_zz_515_)begin
        int_reg_array_7_13_imag <= _zz_568_;
      end
      if(_zz_516_)begin
        int_reg_array_7_14_imag <= _zz_568_;
      end
      if(_zz_517_)begin
        int_reg_array_7_15_imag <= _zz_568_;
      end
      if(_zz_518_)begin
        int_reg_array_7_16_imag <= _zz_568_;
      end
      if(_zz_519_)begin
        int_reg_array_7_17_imag <= _zz_568_;
      end
      if(_zz_520_)begin
        int_reg_array_7_18_imag <= _zz_568_;
      end
      if(_zz_521_)begin
        int_reg_array_7_19_imag <= _zz_568_;
      end
      if(_zz_522_)begin
        int_reg_array_7_20_imag <= _zz_568_;
      end
      if(_zz_523_)begin
        int_reg_array_7_21_imag <= _zz_568_;
      end
      if(_zz_524_)begin
        int_reg_array_7_22_imag <= _zz_568_;
      end
      if(_zz_525_)begin
        int_reg_array_7_23_imag <= _zz_568_;
      end
      if(_zz_526_)begin
        int_reg_array_7_24_imag <= _zz_568_;
      end
      if(_zz_527_)begin
        int_reg_array_7_25_imag <= _zz_568_;
      end
      if(_zz_528_)begin
        int_reg_array_7_26_imag <= _zz_568_;
      end
      if(_zz_529_)begin
        int_reg_array_7_27_imag <= _zz_568_;
      end
      if(_zz_530_)begin
        int_reg_array_7_28_imag <= _zz_568_;
      end
      if(_zz_531_)begin
        int_reg_array_7_29_imag <= _zz_568_;
      end
      if(_zz_532_)begin
        int_reg_array_7_30_imag <= _zz_568_;
      end
      if(_zz_533_)begin
        int_reg_array_7_31_imag <= _zz_568_;
      end
      if(_zz_534_)begin
        int_reg_array_7_32_imag <= _zz_568_;
      end
      if(_zz_535_)begin
        int_reg_array_7_33_imag <= _zz_568_;
      end
      if(_zz_536_)begin
        int_reg_array_7_34_imag <= _zz_568_;
      end
      if(_zz_537_)begin
        int_reg_array_7_35_imag <= _zz_568_;
      end
      if(_zz_538_)begin
        int_reg_array_7_36_imag <= _zz_568_;
      end
      if(_zz_539_)begin
        int_reg_array_7_37_imag <= _zz_568_;
      end
      if(_zz_540_)begin
        int_reg_array_7_38_imag <= _zz_568_;
      end
      if(_zz_541_)begin
        int_reg_array_7_39_imag <= _zz_568_;
      end
      if(_zz_542_)begin
        int_reg_array_7_40_imag <= _zz_568_;
      end
      if(_zz_543_)begin
        int_reg_array_7_41_imag <= _zz_568_;
      end
      if(_zz_544_)begin
        int_reg_array_7_42_imag <= _zz_568_;
      end
      if(_zz_545_)begin
        int_reg_array_7_43_imag <= _zz_568_;
      end
      if(_zz_546_)begin
        int_reg_array_7_44_imag <= _zz_568_;
      end
      if(_zz_547_)begin
        int_reg_array_7_45_imag <= _zz_568_;
      end
      if(_zz_548_)begin
        int_reg_array_7_46_imag <= _zz_568_;
      end
      if(_zz_549_)begin
        int_reg_array_7_47_imag <= _zz_568_;
      end
      if(_zz_550_)begin
        int_reg_array_7_48_imag <= _zz_568_;
      end
      if(_zz_551_)begin
        int_reg_array_7_49_imag <= _zz_568_;
      end
      if(_zz_552_)begin
        int_reg_array_7_50_imag <= _zz_568_;
      end
      if(_zz_553_)begin
        int_reg_array_7_51_imag <= _zz_568_;
      end
      if(_zz_554_)begin
        int_reg_array_7_52_imag <= _zz_568_;
      end
      if(_zz_555_)begin
        int_reg_array_7_53_imag <= _zz_568_;
      end
      if(_zz_556_)begin
        int_reg_array_7_54_imag <= _zz_568_;
      end
      if(_zz_557_)begin
        int_reg_array_7_55_imag <= _zz_568_;
      end
      if(_zz_558_)begin
        int_reg_array_7_56_imag <= _zz_568_;
      end
      if(_zz_559_)begin
        int_reg_array_7_57_imag <= _zz_568_;
      end
      if(_zz_560_)begin
        int_reg_array_7_58_imag <= _zz_568_;
      end
      if(_zz_561_)begin
        int_reg_array_7_59_imag <= _zz_568_;
      end
      if(_zz_562_)begin
        int_reg_array_7_60_imag <= _zz_568_;
      end
      if(_zz_563_)begin
        int_reg_array_7_61_imag <= _zz_568_;
      end
      if(_zz_564_)begin
        int_reg_array_7_62_imag <= _zz_568_;
      end
      if(_zz_565_)begin
        int_reg_array_7_63_imag <= _zz_568_;
      end
      if(_zz_571_)begin
        int_reg_array_8_0_real <= _zz_636_;
      end
      if(_zz_572_)begin
        int_reg_array_8_1_real <= _zz_636_;
      end
      if(_zz_573_)begin
        int_reg_array_8_2_real <= _zz_636_;
      end
      if(_zz_574_)begin
        int_reg_array_8_3_real <= _zz_636_;
      end
      if(_zz_575_)begin
        int_reg_array_8_4_real <= _zz_636_;
      end
      if(_zz_576_)begin
        int_reg_array_8_5_real <= _zz_636_;
      end
      if(_zz_577_)begin
        int_reg_array_8_6_real <= _zz_636_;
      end
      if(_zz_578_)begin
        int_reg_array_8_7_real <= _zz_636_;
      end
      if(_zz_579_)begin
        int_reg_array_8_8_real <= _zz_636_;
      end
      if(_zz_580_)begin
        int_reg_array_8_9_real <= _zz_636_;
      end
      if(_zz_581_)begin
        int_reg_array_8_10_real <= _zz_636_;
      end
      if(_zz_582_)begin
        int_reg_array_8_11_real <= _zz_636_;
      end
      if(_zz_583_)begin
        int_reg_array_8_12_real <= _zz_636_;
      end
      if(_zz_584_)begin
        int_reg_array_8_13_real <= _zz_636_;
      end
      if(_zz_585_)begin
        int_reg_array_8_14_real <= _zz_636_;
      end
      if(_zz_586_)begin
        int_reg_array_8_15_real <= _zz_636_;
      end
      if(_zz_587_)begin
        int_reg_array_8_16_real <= _zz_636_;
      end
      if(_zz_588_)begin
        int_reg_array_8_17_real <= _zz_636_;
      end
      if(_zz_589_)begin
        int_reg_array_8_18_real <= _zz_636_;
      end
      if(_zz_590_)begin
        int_reg_array_8_19_real <= _zz_636_;
      end
      if(_zz_591_)begin
        int_reg_array_8_20_real <= _zz_636_;
      end
      if(_zz_592_)begin
        int_reg_array_8_21_real <= _zz_636_;
      end
      if(_zz_593_)begin
        int_reg_array_8_22_real <= _zz_636_;
      end
      if(_zz_594_)begin
        int_reg_array_8_23_real <= _zz_636_;
      end
      if(_zz_595_)begin
        int_reg_array_8_24_real <= _zz_636_;
      end
      if(_zz_596_)begin
        int_reg_array_8_25_real <= _zz_636_;
      end
      if(_zz_597_)begin
        int_reg_array_8_26_real <= _zz_636_;
      end
      if(_zz_598_)begin
        int_reg_array_8_27_real <= _zz_636_;
      end
      if(_zz_599_)begin
        int_reg_array_8_28_real <= _zz_636_;
      end
      if(_zz_600_)begin
        int_reg_array_8_29_real <= _zz_636_;
      end
      if(_zz_601_)begin
        int_reg_array_8_30_real <= _zz_636_;
      end
      if(_zz_602_)begin
        int_reg_array_8_31_real <= _zz_636_;
      end
      if(_zz_603_)begin
        int_reg_array_8_32_real <= _zz_636_;
      end
      if(_zz_604_)begin
        int_reg_array_8_33_real <= _zz_636_;
      end
      if(_zz_605_)begin
        int_reg_array_8_34_real <= _zz_636_;
      end
      if(_zz_606_)begin
        int_reg_array_8_35_real <= _zz_636_;
      end
      if(_zz_607_)begin
        int_reg_array_8_36_real <= _zz_636_;
      end
      if(_zz_608_)begin
        int_reg_array_8_37_real <= _zz_636_;
      end
      if(_zz_609_)begin
        int_reg_array_8_38_real <= _zz_636_;
      end
      if(_zz_610_)begin
        int_reg_array_8_39_real <= _zz_636_;
      end
      if(_zz_611_)begin
        int_reg_array_8_40_real <= _zz_636_;
      end
      if(_zz_612_)begin
        int_reg_array_8_41_real <= _zz_636_;
      end
      if(_zz_613_)begin
        int_reg_array_8_42_real <= _zz_636_;
      end
      if(_zz_614_)begin
        int_reg_array_8_43_real <= _zz_636_;
      end
      if(_zz_615_)begin
        int_reg_array_8_44_real <= _zz_636_;
      end
      if(_zz_616_)begin
        int_reg_array_8_45_real <= _zz_636_;
      end
      if(_zz_617_)begin
        int_reg_array_8_46_real <= _zz_636_;
      end
      if(_zz_618_)begin
        int_reg_array_8_47_real <= _zz_636_;
      end
      if(_zz_619_)begin
        int_reg_array_8_48_real <= _zz_636_;
      end
      if(_zz_620_)begin
        int_reg_array_8_49_real <= _zz_636_;
      end
      if(_zz_621_)begin
        int_reg_array_8_50_real <= _zz_636_;
      end
      if(_zz_622_)begin
        int_reg_array_8_51_real <= _zz_636_;
      end
      if(_zz_623_)begin
        int_reg_array_8_52_real <= _zz_636_;
      end
      if(_zz_624_)begin
        int_reg_array_8_53_real <= _zz_636_;
      end
      if(_zz_625_)begin
        int_reg_array_8_54_real <= _zz_636_;
      end
      if(_zz_626_)begin
        int_reg_array_8_55_real <= _zz_636_;
      end
      if(_zz_627_)begin
        int_reg_array_8_56_real <= _zz_636_;
      end
      if(_zz_628_)begin
        int_reg_array_8_57_real <= _zz_636_;
      end
      if(_zz_629_)begin
        int_reg_array_8_58_real <= _zz_636_;
      end
      if(_zz_630_)begin
        int_reg_array_8_59_real <= _zz_636_;
      end
      if(_zz_631_)begin
        int_reg_array_8_60_real <= _zz_636_;
      end
      if(_zz_632_)begin
        int_reg_array_8_61_real <= _zz_636_;
      end
      if(_zz_633_)begin
        int_reg_array_8_62_real <= _zz_636_;
      end
      if(_zz_634_)begin
        int_reg_array_8_63_real <= _zz_636_;
      end
      if(_zz_571_)begin
        int_reg_array_8_0_imag <= _zz_637_;
      end
      if(_zz_572_)begin
        int_reg_array_8_1_imag <= _zz_637_;
      end
      if(_zz_573_)begin
        int_reg_array_8_2_imag <= _zz_637_;
      end
      if(_zz_574_)begin
        int_reg_array_8_3_imag <= _zz_637_;
      end
      if(_zz_575_)begin
        int_reg_array_8_4_imag <= _zz_637_;
      end
      if(_zz_576_)begin
        int_reg_array_8_5_imag <= _zz_637_;
      end
      if(_zz_577_)begin
        int_reg_array_8_6_imag <= _zz_637_;
      end
      if(_zz_578_)begin
        int_reg_array_8_7_imag <= _zz_637_;
      end
      if(_zz_579_)begin
        int_reg_array_8_8_imag <= _zz_637_;
      end
      if(_zz_580_)begin
        int_reg_array_8_9_imag <= _zz_637_;
      end
      if(_zz_581_)begin
        int_reg_array_8_10_imag <= _zz_637_;
      end
      if(_zz_582_)begin
        int_reg_array_8_11_imag <= _zz_637_;
      end
      if(_zz_583_)begin
        int_reg_array_8_12_imag <= _zz_637_;
      end
      if(_zz_584_)begin
        int_reg_array_8_13_imag <= _zz_637_;
      end
      if(_zz_585_)begin
        int_reg_array_8_14_imag <= _zz_637_;
      end
      if(_zz_586_)begin
        int_reg_array_8_15_imag <= _zz_637_;
      end
      if(_zz_587_)begin
        int_reg_array_8_16_imag <= _zz_637_;
      end
      if(_zz_588_)begin
        int_reg_array_8_17_imag <= _zz_637_;
      end
      if(_zz_589_)begin
        int_reg_array_8_18_imag <= _zz_637_;
      end
      if(_zz_590_)begin
        int_reg_array_8_19_imag <= _zz_637_;
      end
      if(_zz_591_)begin
        int_reg_array_8_20_imag <= _zz_637_;
      end
      if(_zz_592_)begin
        int_reg_array_8_21_imag <= _zz_637_;
      end
      if(_zz_593_)begin
        int_reg_array_8_22_imag <= _zz_637_;
      end
      if(_zz_594_)begin
        int_reg_array_8_23_imag <= _zz_637_;
      end
      if(_zz_595_)begin
        int_reg_array_8_24_imag <= _zz_637_;
      end
      if(_zz_596_)begin
        int_reg_array_8_25_imag <= _zz_637_;
      end
      if(_zz_597_)begin
        int_reg_array_8_26_imag <= _zz_637_;
      end
      if(_zz_598_)begin
        int_reg_array_8_27_imag <= _zz_637_;
      end
      if(_zz_599_)begin
        int_reg_array_8_28_imag <= _zz_637_;
      end
      if(_zz_600_)begin
        int_reg_array_8_29_imag <= _zz_637_;
      end
      if(_zz_601_)begin
        int_reg_array_8_30_imag <= _zz_637_;
      end
      if(_zz_602_)begin
        int_reg_array_8_31_imag <= _zz_637_;
      end
      if(_zz_603_)begin
        int_reg_array_8_32_imag <= _zz_637_;
      end
      if(_zz_604_)begin
        int_reg_array_8_33_imag <= _zz_637_;
      end
      if(_zz_605_)begin
        int_reg_array_8_34_imag <= _zz_637_;
      end
      if(_zz_606_)begin
        int_reg_array_8_35_imag <= _zz_637_;
      end
      if(_zz_607_)begin
        int_reg_array_8_36_imag <= _zz_637_;
      end
      if(_zz_608_)begin
        int_reg_array_8_37_imag <= _zz_637_;
      end
      if(_zz_609_)begin
        int_reg_array_8_38_imag <= _zz_637_;
      end
      if(_zz_610_)begin
        int_reg_array_8_39_imag <= _zz_637_;
      end
      if(_zz_611_)begin
        int_reg_array_8_40_imag <= _zz_637_;
      end
      if(_zz_612_)begin
        int_reg_array_8_41_imag <= _zz_637_;
      end
      if(_zz_613_)begin
        int_reg_array_8_42_imag <= _zz_637_;
      end
      if(_zz_614_)begin
        int_reg_array_8_43_imag <= _zz_637_;
      end
      if(_zz_615_)begin
        int_reg_array_8_44_imag <= _zz_637_;
      end
      if(_zz_616_)begin
        int_reg_array_8_45_imag <= _zz_637_;
      end
      if(_zz_617_)begin
        int_reg_array_8_46_imag <= _zz_637_;
      end
      if(_zz_618_)begin
        int_reg_array_8_47_imag <= _zz_637_;
      end
      if(_zz_619_)begin
        int_reg_array_8_48_imag <= _zz_637_;
      end
      if(_zz_620_)begin
        int_reg_array_8_49_imag <= _zz_637_;
      end
      if(_zz_621_)begin
        int_reg_array_8_50_imag <= _zz_637_;
      end
      if(_zz_622_)begin
        int_reg_array_8_51_imag <= _zz_637_;
      end
      if(_zz_623_)begin
        int_reg_array_8_52_imag <= _zz_637_;
      end
      if(_zz_624_)begin
        int_reg_array_8_53_imag <= _zz_637_;
      end
      if(_zz_625_)begin
        int_reg_array_8_54_imag <= _zz_637_;
      end
      if(_zz_626_)begin
        int_reg_array_8_55_imag <= _zz_637_;
      end
      if(_zz_627_)begin
        int_reg_array_8_56_imag <= _zz_637_;
      end
      if(_zz_628_)begin
        int_reg_array_8_57_imag <= _zz_637_;
      end
      if(_zz_629_)begin
        int_reg_array_8_58_imag <= _zz_637_;
      end
      if(_zz_630_)begin
        int_reg_array_8_59_imag <= _zz_637_;
      end
      if(_zz_631_)begin
        int_reg_array_8_60_imag <= _zz_637_;
      end
      if(_zz_632_)begin
        int_reg_array_8_61_imag <= _zz_637_;
      end
      if(_zz_633_)begin
        int_reg_array_8_62_imag <= _zz_637_;
      end
      if(_zz_634_)begin
        int_reg_array_8_63_imag <= _zz_637_;
      end
      if(_zz_640_)begin
        int_reg_array_9_0_real <= _zz_705_;
      end
      if(_zz_641_)begin
        int_reg_array_9_1_real <= _zz_705_;
      end
      if(_zz_642_)begin
        int_reg_array_9_2_real <= _zz_705_;
      end
      if(_zz_643_)begin
        int_reg_array_9_3_real <= _zz_705_;
      end
      if(_zz_644_)begin
        int_reg_array_9_4_real <= _zz_705_;
      end
      if(_zz_645_)begin
        int_reg_array_9_5_real <= _zz_705_;
      end
      if(_zz_646_)begin
        int_reg_array_9_6_real <= _zz_705_;
      end
      if(_zz_647_)begin
        int_reg_array_9_7_real <= _zz_705_;
      end
      if(_zz_648_)begin
        int_reg_array_9_8_real <= _zz_705_;
      end
      if(_zz_649_)begin
        int_reg_array_9_9_real <= _zz_705_;
      end
      if(_zz_650_)begin
        int_reg_array_9_10_real <= _zz_705_;
      end
      if(_zz_651_)begin
        int_reg_array_9_11_real <= _zz_705_;
      end
      if(_zz_652_)begin
        int_reg_array_9_12_real <= _zz_705_;
      end
      if(_zz_653_)begin
        int_reg_array_9_13_real <= _zz_705_;
      end
      if(_zz_654_)begin
        int_reg_array_9_14_real <= _zz_705_;
      end
      if(_zz_655_)begin
        int_reg_array_9_15_real <= _zz_705_;
      end
      if(_zz_656_)begin
        int_reg_array_9_16_real <= _zz_705_;
      end
      if(_zz_657_)begin
        int_reg_array_9_17_real <= _zz_705_;
      end
      if(_zz_658_)begin
        int_reg_array_9_18_real <= _zz_705_;
      end
      if(_zz_659_)begin
        int_reg_array_9_19_real <= _zz_705_;
      end
      if(_zz_660_)begin
        int_reg_array_9_20_real <= _zz_705_;
      end
      if(_zz_661_)begin
        int_reg_array_9_21_real <= _zz_705_;
      end
      if(_zz_662_)begin
        int_reg_array_9_22_real <= _zz_705_;
      end
      if(_zz_663_)begin
        int_reg_array_9_23_real <= _zz_705_;
      end
      if(_zz_664_)begin
        int_reg_array_9_24_real <= _zz_705_;
      end
      if(_zz_665_)begin
        int_reg_array_9_25_real <= _zz_705_;
      end
      if(_zz_666_)begin
        int_reg_array_9_26_real <= _zz_705_;
      end
      if(_zz_667_)begin
        int_reg_array_9_27_real <= _zz_705_;
      end
      if(_zz_668_)begin
        int_reg_array_9_28_real <= _zz_705_;
      end
      if(_zz_669_)begin
        int_reg_array_9_29_real <= _zz_705_;
      end
      if(_zz_670_)begin
        int_reg_array_9_30_real <= _zz_705_;
      end
      if(_zz_671_)begin
        int_reg_array_9_31_real <= _zz_705_;
      end
      if(_zz_672_)begin
        int_reg_array_9_32_real <= _zz_705_;
      end
      if(_zz_673_)begin
        int_reg_array_9_33_real <= _zz_705_;
      end
      if(_zz_674_)begin
        int_reg_array_9_34_real <= _zz_705_;
      end
      if(_zz_675_)begin
        int_reg_array_9_35_real <= _zz_705_;
      end
      if(_zz_676_)begin
        int_reg_array_9_36_real <= _zz_705_;
      end
      if(_zz_677_)begin
        int_reg_array_9_37_real <= _zz_705_;
      end
      if(_zz_678_)begin
        int_reg_array_9_38_real <= _zz_705_;
      end
      if(_zz_679_)begin
        int_reg_array_9_39_real <= _zz_705_;
      end
      if(_zz_680_)begin
        int_reg_array_9_40_real <= _zz_705_;
      end
      if(_zz_681_)begin
        int_reg_array_9_41_real <= _zz_705_;
      end
      if(_zz_682_)begin
        int_reg_array_9_42_real <= _zz_705_;
      end
      if(_zz_683_)begin
        int_reg_array_9_43_real <= _zz_705_;
      end
      if(_zz_684_)begin
        int_reg_array_9_44_real <= _zz_705_;
      end
      if(_zz_685_)begin
        int_reg_array_9_45_real <= _zz_705_;
      end
      if(_zz_686_)begin
        int_reg_array_9_46_real <= _zz_705_;
      end
      if(_zz_687_)begin
        int_reg_array_9_47_real <= _zz_705_;
      end
      if(_zz_688_)begin
        int_reg_array_9_48_real <= _zz_705_;
      end
      if(_zz_689_)begin
        int_reg_array_9_49_real <= _zz_705_;
      end
      if(_zz_690_)begin
        int_reg_array_9_50_real <= _zz_705_;
      end
      if(_zz_691_)begin
        int_reg_array_9_51_real <= _zz_705_;
      end
      if(_zz_692_)begin
        int_reg_array_9_52_real <= _zz_705_;
      end
      if(_zz_693_)begin
        int_reg_array_9_53_real <= _zz_705_;
      end
      if(_zz_694_)begin
        int_reg_array_9_54_real <= _zz_705_;
      end
      if(_zz_695_)begin
        int_reg_array_9_55_real <= _zz_705_;
      end
      if(_zz_696_)begin
        int_reg_array_9_56_real <= _zz_705_;
      end
      if(_zz_697_)begin
        int_reg_array_9_57_real <= _zz_705_;
      end
      if(_zz_698_)begin
        int_reg_array_9_58_real <= _zz_705_;
      end
      if(_zz_699_)begin
        int_reg_array_9_59_real <= _zz_705_;
      end
      if(_zz_700_)begin
        int_reg_array_9_60_real <= _zz_705_;
      end
      if(_zz_701_)begin
        int_reg_array_9_61_real <= _zz_705_;
      end
      if(_zz_702_)begin
        int_reg_array_9_62_real <= _zz_705_;
      end
      if(_zz_703_)begin
        int_reg_array_9_63_real <= _zz_705_;
      end
      if(_zz_640_)begin
        int_reg_array_9_0_imag <= _zz_706_;
      end
      if(_zz_641_)begin
        int_reg_array_9_1_imag <= _zz_706_;
      end
      if(_zz_642_)begin
        int_reg_array_9_2_imag <= _zz_706_;
      end
      if(_zz_643_)begin
        int_reg_array_9_3_imag <= _zz_706_;
      end
      if(_zz_644_)begin
        int_reg_array_9_4_imag <= _zz_706_;
      end
      if(_zz_645_)begin
        int_reg_array_9_5_imag <= _zz_706_;
      end
      if(_zz_646_)begin
        int_reg_array_9_6_imag <= _zz_706_;
      end
      if(_zz_647_)begin
        int_reg_array_9_7_imag <= _zz_706_;
      end
      if(_zz_648_)begin
        int_reg_array_9_8_imag <= _zz_706_;
      end
      if(_zz_649_)begin
        int_reg_array_9_9_imag <= _zz_706_;
      end
      if(_zz_650_)begin
        int_reg_array_9_10_imag <= _zz_706_;
      end
      if(_zz_651_)begin
        int_reg_array_9_11_imag <= _zz_706_;
      end
      if(_zz_652_)begin
        int_reg_array_9_12_imag <= _zz_706_;
      end
      if(_zz_653_)begin
        int_reg_array_9_13_imag <= _zz_706_;
      end
      if(_zz_654_)begin
        int_reg_array_9_14_imag <= _zz_706_;
      end
      if(_zz_655_)begin
        int_reg_array_9_15_imag <= _zz_706_;
      end
      if(_zz_656_)begin
        int_reg_array_9_16_imag <= _zz_706_;
      end
      if(_zz_657_)begin
        int_reg_array_9_17_imag <= _zz_706_;
      end
      if(_zz_658_)begin
        int_reg_array_9_18_imag <= _zz_706_;
      end
      if(_zz_659_)begin
        int_reg_array_9_19_imag <= _zz_706_;
      end
      if(_zz_660_)begin
        int_reg_array_9_20_imag <= _zz_706_;
      end
      if(_zz_661_)begin
        int_reg_array_9_21_imag <= _zz_706_;
      end
      if(_zz_662_)begin
        int_reg_array_9_22_imag <= _zz_706_;
      end
      if(_zz_663_)begin
        int_reg_array_9_23_imag <= _zz_706_;
      end
      if(_zz_664_)begin
        int_reg_array_9_24_imag <= _zz_706_;
      end
      if(_zz_665_)begin
        int_reg_array_9_25_imag <= _zz_706_;
      end
      if(_zz_666_)begin
        int_reg_array_9_26_imag <= _zz_706_;
      end
      if(_zz_667_)begin
        int_reg_array_9_27_imag <= _zz_706_;
      end
      if(_zz_668_)begin
        int_reg_array_9_28_imag <= _zz_706_;
      end
      if(_zz_669_)begin
        int_reg_array_9_29_imag <= _zz_706_;
      end
      if(_zz_670_)begin
        int_reg_array_9_30_imag <= _zz_706_;
      end
      if(_zz_671_)begin
        int_reg_array_9_31_imag <= _zz_706_;
      end
      if(_zz_672_)begin
        int_reg_array_9_32_imag <= _zz_706_;
      end
      if(_zz_673_)begin
        int_reg_array_9_33_imag <= _zz_706_;
      end
      if(_zz_674_)begin
        int_reg_array_9_34_imag <= _zz_706_;
      end
      if(_zz_675_)begin
        int_reg_array_9_35_imag <= _zz_706_;
      end
      if(_zz_676_)begin
        int_reg_array_9_36_imag <= _zz_706_;
      end
      if(_zz_677_)begin
        int_reg_array_9_37_imag <= _zz_706_;
      end
      if(_zz_678_)begin
        int_reg_array_9_38_imag <= _zz_706_;
      end
      if(_zz_679_)begin
        int_reg_array_9_39_imag <= _zz_706_;
      end
      if(_zz_680_)begin
        int_reg_array_9_40_imag <= _zz_706_;
      end
      if(_zz_681_)begin
        int_reg_array_9_41_imag <= _zz_706_;
      end
      if(_zz_682_)begin
        int_reg_array_9_42_imag <= _zz_706_;
      end
      if(_zz_683_)begin
        int_reg_array_9_43_imag <= _zz_706_;
      end
      if(_zz_684_)begin
        int_reg_array_9_44_imag <= _zz_706_;
      end
      if(_zz_685_)begin
        int_reg_array_9_45_imag <= _zz_706_;
      end
      if(_zz_686_)begin
        int_reg_array_9_46_imag <= _zz_706_;
      end
      if(_zz_687_)begin
        int_reg_array_9_47_imag <= _zz_706_;
      end
      if(_zz_688_)begin
        int_reg_array_9_48_imag <= _zz_706_;
      end
      if(_zz_689_)begin
        int_reg_array_9_49_imag <= _zz_706_;
      end
      if(_zz_690_)begin
        int_reg_array_9_50_imag <= _zz_706_;
      end
      if(_zz_691_)begin
        int_reg_array_9_51_imag <= _zz_706_;
      end
      if(_zz_692_)begin
        int_reg_array_9_52_imag <= _zz_706_;
      end
      if(_zz_693_)begin
        int_reg_array_9_53_imag <= _zz_706_;
      end
      if(_zz_694_)begin
        int_reg_array_9_54_imag <= _zz_706_;
      end
      if(_zz_695_)begin
        int_reg_array_9_55_imag <= _zz_706_;
      end
      if(_zz_696_)begin
        int_reg_array_9_56_imag <= _zz_706_;
      end
      if(_zz_697_)begin
        int_reg_array_9_57_imag <= _zz_706_;
      end
      if(_zz_698_)begin
        int_reg_array_9_58_imag <= _zz_706_;
      end
      if(_zz_699_)begin
        int_reg_array_9_59_imag <= _zz_706_;
      end
      if(_zz_700_)begin
        int_reg_array_9_60_imag <= _zz_706_;
      end
      if(_zz_701_)begin
        int_reg_array_9_61_imag <= _zz_706_;
      end
      if(_zz_702_)begin
        int_reg_array_9_62_imag <= _zz_706_;
      end
      if(_zz_703_)begin
        int_reg_array_9_63_imag <= _zz_706_;
      end
      if(_zz_709_)begin
        int_reg_array_10_0_real <= _zz_774_;
      end
      if(_zz_710_)begin
        int_reg_array_10_1_real <= _zz_774_;
      end
      if(_zz_711_)begin
        int_reg_array_10_2_real <= _zz_774_;
      end
      if(_zz_712_)begin
        int_reg_array_10_3_real <= _zz_774_;
      end
      if(_zz_713_)begin
        int_reg_array_10_4_real <= _zz_774_;
      end
      if(_zz_714_)begin
        int_reg_array_10_5_real <= _zz_774_;
      end
      if(_zz_715_)begin
        int_reg_array_10_6_real <= _zz_774_;
      end
      if(_zz_716_)begin
        int_reg_array_10_7_real <= _zz_774_;
      end
      if(_zz_717_)begin
        int_reg_array_10_8_real <= _zz_774_;
      end
      if(_zz_718_)begin
        int_reg_array_10_9_real <= _zz_774_;
      end
      if(_zz_719_)begin
        int_reg_array_10_10_real <= _zz_774_;
      end
      if(_zz_720_)begin
        int_reg_array_10_11_real <= _zz_774_;
      end
      if(_zz_721_)begin
        int_reg_array_10_12_real <= _zz_774_;
      end
      if(_zz_722_)begin
        int_reg_array_10_13_real <= _zz_774_;
      end
      if(_zz_723_)begin
        int_reg_array_10_14_real <= _zz_774_;
      end
      if(_zz_724_)begin
        int_reg_array_10_15_real <= _zz_774_;
      end
      if(_zz_725_)begin
        int_reg_array_10_16_real <= _zz_774_;
      end
      if(_zz_726_)begin
        int_reg_array_10_17_real <= _zz_774_;
      end
      if(_zz_727_)begin
        int_reg_array_10_18_real <= _zz_774_;
      end
      if(_zz_728_)begin
        int_reg_array_10_19_real <= _zz_774_;
      end
      if(_zz_729_)begin
        int_reg_array_10_20_real <= _zz_774_;
      end
      if(_zz_730_)begin
        int_reg_array_10_21_real <= _zz_774_;
      end
      if(_zz_731_)begin
        int_reg_array_10_22_real <= _zz_774_;
      end
      if(_zz_732_)begin
        int_reg_array_10_23_real <= _zz_774_;
      end
      if(_zz_733_)begin
        int_reg_array_10_24_real <= _zz_774_;
      end
      if(_zz_734_)begin
        int_reg_array_10_25_real <= _zz_774_;
      end
      if(_zz_735_)begin
        int_reg_array_10_26_real <= _zz_774_;
      end
      if(_zz_736_)begin
        int_reg_array_10_27_real <= _zz_774_;
      end
      if(_zz_737_)begin
        int_reg_array_10_28_real <= _zz_774_;
      end
      if(_zz_738_)begin
        int_reg_array_10_29_real <= _zz_774_;
      end
      if(_zz_739_)begin
        int_reg_array_10_30_real <= _zz_774_;
      end
      if(_zz_740_)begin
        int_reg_array_10_31_real <= _zz_774_;
      end
      if(_zz_741_)begin
        int_reg_array_10_32_real <= _zz_774_;
      end
      if(_zz_742_)begin
        int_reg_array_10_33_real <= _zz_774_;
      end
      if(_zz_743_)begin
        int_reg_array_10_34_real <= _zz_774_;
      end
      if(_zz_744_)begin
        int_reg_array_10_35_real <= _zz_774_;
      end
      if(_zz_745_)begin
        int_reg_array_10_36_real <= _zz_774_;
      end
      if(_zz_746_)begin
        int_reg_array_10_37_real <= _zz_774_;
      end
      if(_zz_747_)begin
        int_reg_array_10_38_real <= _zz_774_;
      end
      if(_zz_748_)begin
        int_reg_array_10_39_real <= _zz_774_;
      end
      if(_zz_749_)begin
        int_reg_array_10_40_real <= _zz_774_;
      end
      if(_zz_750_)begin
        int_reg_array_10_41_real <= _zz_774_;
      end
      if(_zz_751_)begin
        int_reg_array_10_42_real <= _zz_774_;
      end
      if(_zz_752_)begin
        int_reg_array_10_43_real <= _zz_774_;
      end
      if(_zz_753_)begin
        int_reg_array_10_44_real <= _zz_774_;
      end
      if(_zz_754_)begin
        int_reg_array_10_45_real <= _zz_774_;
      end
      if(_zz_755_)begin
        int_reg_array_10_46_real <= _zz_774_;
      end
      if(_zz_756_)begin
        int_reg_array_10_47_real <= _zz_774_;
      end
      if(_zz_757_)begin
        int_reg_array_10_48_real <= _zz_774_;
      end
      if(_zz_758_)begin
        int_reg_array_10_49_real <= _zz_774_;
      end
      if(_zz_759_)begin
        int_reg_array_10_50_real <= _zz_774_;
      end
      if(_zz_760_)begin
        int_reg_array_10_51_real <= _zz_774_;
      end
      if(_zz_761_)begin
        int_reg_array_10_52_real <= _zz_774_;
      end
      if(_zz_762_)begin
        int_reg_array_10_53_real <= _zz_774_;
      end
      if(_zz_763_)begin
        int_reg_array_10_54_real <= _zz_774_;
      end
      if(_zz_764_)begin
        int_reg_array_10_55_real <= _zz_774_;
      end
      if(_zz_765_)begin
        int_reg_array_10_56_real <= _zz_774_;
      end
      if(_zz_766_)begin
        int_reg_array_10_57_real <= _zz_774_;
      end
      if(_zz_767_)begin
        int_reg_array_10_58_real <= _zz_774_;
      end
      if(_zz_768_)begin
        int_reg_array_10_59_real <= _zz_774_;
      end
      if(_zz_769_)begin
        int_reg_array_10_60_real <= _zz_774_;
      end
      if(_zz_770_)begin
        int_reg_array_10_61_real <= _zz_774_;
      end
      if(_zz_771_)begin
        int_reg_array_10_62_real <= _zz_774_;
      end
      if(_zz_772_)begin
        int_reg_array_10_63_real <= _zz_774_;
      end
      if(_zz_709_)begin
        int_reg_array_10_0_imag <= _zz_775_;
      end
      if(_zz_710_)begin
        int_reg_array_10_1_imag <= _zz_775_;
      end
      if(_zz_711_)begin
        int_reg_array_10_2_imag <= _zz_775_;
      end
      if(_zz_712_)begin
        int_reg_array_10_3_imag <= _zz_775_;
      end
      if(_zz_713_)begin
        int_reg_array_10_4_imag <= _zz_775_;
      end
      if(_zz_714_)begin
        int_reg_array_10_5_imag <= _zz_775_;
      end
      if(_zz_715_)begin
        int_reg_array_10_6_imag <= _zz_775_;
      end
      if(_zz_716_)begin
        int_reg_array_10_7_imag <= _zz_775_;
      end
      if(_zz_717_)begin
        int_reg_array_10_8_imag <= _zz_775_;
      end
      if(_zz_718_)begin
        int_reg_array_10_9_imag <= _zz_775_;
      end
      if(_zz_719_)begin
        int_reg_array_10_10_imag <= _zz_775_;
      end
      if(_zz_720_)begin
        int_reg_array_10_11_imag <= _zz_775_;
      end
      if(_zz_721_)begin
        int_reg_array_10_12_imag <= _zz_775_;
      end
      if(_zz_722_)begin
        int_reg_array_10_13_imag <= _zz_775_;
      end
      if(_zz_723_)begin
        int_reg_array_10_14_imag <= _zz_775_;
      end
      if(_zz_724_)begin
        int_reg_array_10_15_imag <= _zz_775_;
      end
      if(_zz_725_)begin
        int_reg_array_10_16_imag <= _zz_775_;
      end
      if(_zz_726_)begin
        int_reg_array_10_17_imag <= _zz_775_;
      end
      if(_zz_727_)begin
        int_reg_array_10_18_imag <= _zz_775_;
      end
      if(_zz_728_)begin
        int_reg_array_10_19_imag <= _zz_775_;
      end
      if(_zz_729_)begin
        int_reg_array_10_20_imag <= _zz_775_;
      end
      if(_zz_730_)begin
        int_reg_array_10_21_imag <= _zz_775_;
      end
      if(_zz_731_)begin
        int_reg_array_10_22_imag <= _zz_775_;
      end
      if(_zz_732_)begin
        int_reg_array_10_23_imag <= _zz_775_;
      end
      if(_zz_733_)begin
        int_reg_array_10_24_imag <= _zz_775_;
      end
      if(_zz_734_)begin
        int_reg_array_10_25_imag <= _zz_775_;
      end
      if(_zz_735_)begin
        int_reg_array_10_26_imag <= _zz_775_;
      end
      if(_zz_736_)begin
        int_reg_array_10_27_imag <= _zz_775_;
      end
      if(_zz_737_)begin
        int_reg_array_10_28_imag <= _zz_775_;
      end
      if(_zz_738_)begin
        int_reg_array_10_29_imag <= _zz_775_;
      end
      if(_zz_739_)begin
        int_reg_array_10_30_imag <= _zz_775_;
      end
      if(_zz_740_)begin
        int_reg_array_10_31_imag <= _zz_775_;
      end
      if(_zz_741_)begin
        int_reg_array_10_32_imag <= _zz_775_;
      end
      if(_zz_742_)begin
        int_reg_array_10_33_imag <= _zz_775_;
      end
      if(_zz_743_)begin
        int_reg_array_10_34_imag <= _zz_775_;
      end
      if(_zz_744_)begin
        int_reg_array_10_35_imag <= _zz_775_;
      end
      if(_zz_745_)begin
        int_reg_array_10_36_imag <= _zz_775_;
      end
      if(_zz_746_)begin
        int_reg_array_10_37_imag <= _zz_775_;
      end
      if(_zz_747_)begin
        int_reg_array_10_38_imag <= _zz_775_;
      end
      if(_zz_748_)begin
        int_reg_array_10_39_imag <= _zz_775_;
      end
      if(_zz_749_)begin
        int_reg_array_10_40_imag <= _zz_775_;
      end
      if(_zz_750_)begin
        int_reg_array_10_41_imag <= _zz_775_;
      end
      if(_zz_751_)begin
        int_reg_array_10_42_imag <= _zz_775_;
      end
      if(_zz_752_)begin
        int_reg_array_10_43_imag <= _zz_775_;
      end
      if(_zz_753_)begin
        int_reg_array_10_44_imag <= _zz_775_;
      end
      if(_zz_754_)begin
        int_reg_array_10_45_imag <= _zz_775_;
      end
      if(_zz_755_)begin
        int_reg_array_10_46_imag <= _zz_775_;
      end
      if(_zz_756_)begin
        int_reg_array_10_47_imag <= _zz_775_;
      end
      if(_zz_757_)begin
        int_reg_array_10_48_imag <= _zz_775_;
      end
      if(_zz_758_)begin
        int_reg_array_10_49_imag <= _zz_775_;
      end
      if(_zz_759_)begin
        int_reg_array_10_50_imag <= _zz_775_;
      end
      if(_zz_760_)begin
        int_reg_array_10_51_imag <= _zz_775_;
      end
      if(_zz_761_)begin
        int_reg_array_10_52_imag <= _zz_775_;
      end
      if(_zz_762_)begin
        int_reg_array_10_53_imag <= _zz_775_;
      end
      if(_zz_763_)begin
        int_reg_array_10_54_imag <= _zz_775_;
      end
      if(_zz_764_)begin
        int_reg_array_10_55_imag <= _zz_775_;
      end
      if(_zz_765_)begin
        int_reg_array_10_56_imag <= _zz_775_;
      end
      if(_zz_766_)begin
        int_reg_array_10_57_imag <= _zz_775_;
      end
      if(_zz_767_)begin
        int_reg_array_10_58_imag <= _zz_775_;
      end
      if(_zz_768_)begin
        int_reg_array_10_59_imag <= _zz_775_;
      end
      if(_zz_769_)begin
        int_reg_array_10_60_imag <= _zz_775_;
      end
      if(_zz_770_)begin
        int_reg_array_10_61_imag <= _zz_775_;
      end
      if(_zz_771_)begin
        int_reg_array_10_62_imag <= _zz_775_;
      end
      if(_zz_772_)begin
        int_reg_array_10_63_imag <= _zz_775_;
      end
      if(_zz_778_)begin
        int_reg_array_11_0_real <= _zz_843_;
      end
      if(_zz_779_)begin
        int_reg_array_11_1_real <= _zz_843_;
      end
      if(_zz_780_)begin
        int_reg_array_11_2_real <= _zz_843_;
      end
      if(_zz_781_)begin
        int_reg_array_11_3_real <= _zz_843_;
      end
      if(_zz_782_)begin
        int_reg_array_11_4_real <= _zz_843_;
      end
      if(_zz_783_)begin
        int_reg_array_11_5_real <= _zz_843_;
      end
      if(_zz_784_)begin
        int_reg_array_11_6_real <= _zz_843_;
      end
      if(_zz_785_)begin
        int_reg_array_11_7_real <= _zz_843_;
      end
      if(_zz_786_)begin
        int_reg_array_11_8_real <= _zz_843_;
      end
      if(_zz_787_)begin
        int_reg_array_11_9_real <= _zz_843_;
      end
      if(_zz_788_)begin
        int_reg_array_11_10_real <= _zz_843_;
      end
      if(_zz_789_)begin
        int_reg_array_11_11_real <= _zz_843_;
      end
      if(_zz_790_)begin
        int_reg_array_11_12_real <= _zz_843_;
      end
      if(_zz_791_)begin
        int_reg_array_11_13_real <= _zz_843_;
      end
      if(_zz_792_)begin
        int_reg_array_11_14_real <= _zz_843_;
      end
      if(_zz_793_)begin
        int_reg_array_11_15_real <= _zz_843_;
      end
      if(_zz_794_)begin
        int_reg_array_11_16_real <= _zz_843_;
      end
      if(_zz_795_)begin
        int_reg_array_11_17_real <= _zz_843_;
      end
      if(_zz_796_)begin
        int_reg_array_11_18_real <= _zz_843_;
      end
      if(_zz_797_)begin
        int_reg_array_11_19_real <= _zz_843_;
      end
      if(_zz_798_)begin
        int_reg_array_11_20_real <= _zz_843_;
      end
      if(_zz_799_)begin
        int_reg_array_11_21_real <= _zz_843_;
      end
      if(_zz_800_)begin
        int_reg_array_11_22_real <= _zz_843_;
      end
      if(_zz_801_)begin
        int_reg_array_11_23_real <= _zz_843_;
      end
      if(_zz_802_)begin
        int_reg_array_11_24_real <= _zz_843_;
      end
      if(_zz_803_)begin
        int_reg_array_11_25_real <= _zz_843_;
      end
      if(_zz_804_)begin
        int_reg_array_11_26_real <= _zz_843_;
      end
      if(_zz_805_)begin
        int_reg_array_11_27_real <= _zz_843_;
      end
      if(_zz_806_)begin
        int_reg_array_11_28_real <= _zz_843_;
      end
      if(_zz_807_)begin
        int_reg_array_11_29_real <= _zz_843_;
      end
      if(_zz_808_)begin
        int_reg_array_11_30_real <= _zz_843_;
      end
      if(_zz_809_)begin
        int_reg_array_11_31_real <= _zz_843_;
      end
      if(_zz_810_)begin
        int_reg_array_11_32_real <= _zz_843_;
      end
      if(_zz_811_)begin
        int_reg_array_11_33_real <= _zz_843_;
      end
      if(_zz_812_)begin
        int_reg_array_11_34_real <= _zz_843_;
      end
      if(_zz_813_)begin
        int_reg_array_11_35_real <= _zz_843_;
      end
      if(_zz_814_)begin
        int_reg_array_11_36_real <= _zz_843_;
      end
      if(_zz_815_)begin
        int_reg_array_11_37_real <= _zz_843_;
      end
      if(_zz_816_)begin
        int_reg_array_11_38_real <= _zz_843_;
      end
      if(_zz_817_)begin
        int_reg_array_11_39_real <= _zz_843_;
      end
      if(_zz_818_)begin
        int_reg_array_11_40_real <= _zz_843_;
      end
      if(_zz_819_)begin
        int_reg_array_11_41_real <= _zz_843_;
      end
      if(_zz_820_)begin
        int_reg_array_11_42_real <= _zz_843_;
      end
      if(_zz_821_)begin
        int_reg_array_11_43_real <= _zz_843_;
      end
      if(_zz_822_)begin
        int_reg_array_11_44_real <= _zz_843_;
      end
      if(_zz_823_)begin
        int_reg_array_11_45_real <= _zz_843_;
      end
      if(_zz_824_)begin
        int_reg_array_11_46_real <= _zz_843_;
      end
      if(_zz_825_)begin
        int_reg_array_11_47_real <= _zz_843_;
      end
      if(_zz_826_)begin
        int_reg_array_11_48_real <= _zz_843_;
      end
      if(_zz_827_)begin
        int_reg_array_11_49_real <= _zz_843_;
      end
      if(_zz_828_)begin
        int_reg_array_11_50_real <= _zz_843_;
      end
      if(_zz_829_)begin
        int_reg_array_11_51_real <= _zz_843_;
      end
      if(_zz_830_)begin
        int_reg_array_11_52_real <= _zz_843_;
      end
      if(_zz_831_)begin
        int_reg_array_11_53_real <= _zz_843_;
      end
      if(_zz_832_)begin
        int_reg_array_11_54_real <= _zz_843_;
      end
      if(_zz_833_)begin
        int_reg_array_11_55_real <= _zz_843_;
      end
      if(_zz_834_)begin
        int_reg_array_11_56_real <= _zz_843_;
      end
      if(_zz_835_)begin
        int_reg_array_11_57_real <= _zz_843_;
      end
      if(_zz_836_)begin
        int_reg_array_11_58_real <= _zz_843_;
      end
      if(_zz_837_)begin
        int_reg_array_11_59_real <= _zz_843_;
      end
      if(_zz_838_)begin
        int_reg_array_11_60_real <= _zz_843_;
      end
      if(_zz_839_)begin
        int_reg_array_11_61_real <= _zz_843_;
      end
      if(_zz_840_)begin
        int_reg_array_11_62_real <= _zz_843_;
      end
      if(_zz_841_)begin
        int_reg_array_11_63_real <= _zz_843_;
      end
      if(_zz_778_)begin
        int_reg_array_11_0_imag <= _zz_844_;
      end
      if(_zz_779_)begin
        int_reg_array_11_1_imag <= _zz_844_;
      end
      if(_zz_780_)begin
        int_reg_array_11_2_imag <= _zz_844_;
      end
      if(_zz_781_)begin
        int_reg_array_11_3_imag <= _zz_844_;
      end
      if(_zz_782_)begin
        int_reg_array_11_4_imag <= _zz_844_;
      end
      if(_zz_783_)begin
        int_reg_array_11_5_imag <= _zz_844_;
      end
      if(_zz_784_)begin
        int_reg_array_11_6_imag <= _zz_844_;
      end
      if(_zz_785_)begin
        int_reg_array_11_7_imag <= _zz_844_;
      end
      if(_zz_786_)begin
        int_reg_array_11_8_imag <= _zz_844_;
      end
      if(_zz_787_)begin
        int_reg_array_11_9_imag <= _zz_844_;
      end
      if(_zz_788_)begin
        int_reg_array_11_10_imag <= _zz_844_;
      end
      if(_zz_789_)begin
        int_reg_array_11_11_imag <= _zz_844_;
      end
      if(_zz_790_)begin
        int_reg_array_11_12_imag <= _zz_844_;
      end
      if(_zz_791_)begin
        int_reg_array_11_13_imag <= _zz_844_;
      end
      if(_zz_792_)begin
        int_reg_array_11_14_imag <= _zz_844_;
      end
      if(_zz_793_)begin
        int_reg_array_11_15_imag <= _zz_844_;
      end
      if(_zz_794_)begin
        int_reg_array_11_16_imag <= _zz_844_;
      end
      if(_zz_795_)begin
        int_reg_array_11_17_imag <= _zz_844_;
      end
      if(_zz_796_)begin
        int_reg_array_11_18_imag <= _zz_844_;
      end
      if(_zz_797_)begin
        int_reg_array_11_19_imag <= _zz_844_;
      end
      if(_zz_798_)begin
        int_reg_array_11_20_imag <= _zz_844_;
      end
      if(_zz_799_)begin
        int_reg_array_11_21_imag <= _zz_844_;
      end
      if(_zz_800_)begin
        int_reg_array_11_22_imag <= _zz_844_;
      end
      if(_zz_801_)begin
        int_reg_array_11_23_imag <= _zz_844_;
      end
      if(_zz_802_)begin
        int_reg_array_11_24_imag <= _zz_844_;
      end
      if(_zz_803_)begin
        int_reg_array_11_25_imag <= _zz_844_;
      end
      if(_zz_804_)begin
        int_reg_array_11_26_imag <= _zz_844_;
      end
      if(_zz_805_)begin
        int_reg_array_11_27_imag <= _zz_844_;
      end
      if(_zz_806_)begin
        int_reg_array_11_28_imag <= _zz_844_;
      end
      if(_zz_807_)begin
        int_reg_array_11_29_imag <= _zz_844_;
      end
      if(_zz_808_)begin
        int_reg_array_11_30_imag <= _zz_844_;
      end
      if(_zz_809_)begin
        int_reg_array_11_31_imag <= _zz_844_;
      end
      if(_zz_810_)begin
        int_reg_array_11_32_imag <= _zz_844_;
      end
      if(_zz_811_)begin
        int_reg_array_11_33_imag <= _zz_844_;
      end
      if(_zz_812_)begin
        int_reg_array_11_34_imag <= _zz_844_;
      end
      if(_zz_813_)begin
        int_reg_array_11_35_imag <= _zz_844_;
      end
      if(_zz_814_)begin
        int_reg_array_11_36_imag <= _zz_844_;
      end
      if(_zz_815_)begin
        int_reg_array_11_37_imag <= _zz_844_;
      end
      if(_zz_816_)begin
        int_reg_array_11_38_imag <= _zz_844_;
      end
      if(_zz_817_)begin
        int_reg_array_11_39_imag <= _zz_844_;
      end
      if(_zz_818_)begin
        int_reg_array_11_40_imag <= _zz_844_;
      end
      if(_zz_819_)begin
        int_reg_array_11_41_imag <= _zz_844_;
      end
      if(_zz_820_)begin
        int_reg_array_11_42_imag <= _zz_844_;
      end
      if(_zz_821_)begin
        int_reg_array_11_43_imag <= _zz_844_;
      end
      if(_zz_822_)begin
        int_reg_array_11_44_imag <= _zz_844_;
      end
      if(_zz_823_)begin
        int_reg_array_11_45_imag <= _zz_844_;
      end
      if(_zz_824_)begin
        int_reg_array_11_46_imag <= _zz_844_;
      end
      if(_zz_825_)begin
        int_reg_array_11_47_imag <= _zz_844_;
      end
      if(_zz_826_)begin
        int_reg_array_11_48_imag <= _zz_844_;
      end
      if(_zz_827_)begin
        int_reg_array_11_49_imag <= _zz_844_;
      end
      if(_zz_828_)begin
        int_reg_array_11_50_imag <= _zz_844_;
      end
      if(_zz_829_)begin
        int_reg_array_11_51_imag <= _zz_844_;
      end
      if(_zz_830_)begin
        int_reg_array_11_52_imag <= _zz_844_;
      end
      if(_zz_831_)begin
        int_reg_array_11_53_imag <= _zz_844_;
      end
      if(_zz_832_)begin
        int_reg_array_11_54_imag <= _zz_844_;
      end
      if(_zz_833_)begin
        int_reg_array_11_55_imag <= _zz_844_;
      end
      if(_zz_834_)begin
        int_reg_array_11_56_imag <= _zz_844_;
      end
      if(_zz_835_)begin
        int_reg_array_11_57_imag <= _zz_844_;
      end
      if(_zz_836_)begin
        int_reg_array_11_58_imag <= _zz_844_;
      end
      if(_zz_837_)begin
        int_reg_array_11_59_imag <= _zz_844_;
      end
      if(_zz_838_)begin
        int_reg_array_11_60_imag <= _zz_844_;
      end
      if(_zz_839_)begin
        int_reg_array_11_61_imag <= _zz_844_;
      end
      if(_zz_840_)begin
        int_reg_array_11_62_imag <= _zz_844_;
      end
      if(_zz_841_)begin
        int_reg_array_11_63_imag <= _zz_844_;
      end
      if(_zz_847_)begin
        int_reg_array_12_0_real <= _zz_912_;
      end
      if(_zz_848_)begin
        int_reg_array_12_1_real <= _zz_912_;
      end
      if(_zz_849_)begin
        int_reg_array_12_2_real <= _zz_912_;
      end
      if(_zz_850_)begin
        int_reg_array_12_3_real <= _zz_912_;
      end
      if(_zz_851_)begin
        int_reg_array_12_4_real <= _zz_912_;
      end
      if(_zz_852_)begin
        int_reg_array_12_5_real <= _zz_912_;
      end
      if(_zz_853_)begin
        int_reg_array_12_6_real <= _zz_912_;
      end
      if(_zz_854_)begin
        int_reg_array_12_7_real <= _zz_912_;
      end
      if(_zz_855_)begin
        int_reg_array_12_8_real <= _zz_912_;
      end
      if(_zz_856_)begin
        int_reg_array_12_9_real <= _zz_912_;
      end
      if(_zz_857_)begin
        int_reg_array_12_10_real <= _zz_912_;
      end
      if(_zz_858_)begin
        int_reg_array_12_11_real <= _zz_912_;
      end
      if(_zz_859_)begin
        int_reg_array_12_12_real <= _zz_912_;
      end
      if(_zz_860_)begin
        int_reg_array_12_13_real <= _zz_912_;
      end
      if(_zz_861_)begin
        int_reg_array_12_14_real <= _zz_912_;
      end
      if(_zz_862_)begin
        int_reg_array_12_15_real <= _zz_912_;
      end
      if(_zz_863_)begin
        int_reg_array_12_16_real <= _zz_912_;
      end
      if(_zz_864_)begin
        int_reg_array_12_17_real <= _zz_912_;
      end
      if(_zz_865_)begin
        int_reg_array_12_18_real <= _zz_912_;
      end
      if(_zz_866_)begin
        int_reg_array_12_19_real <= _zz_912_;
      end
      if(_zz_867_)begin
        int_reg_array_12_20_real <= _zz_912_;
      end
      if(_zz_868_)begin
        int_reg_array_12_21_real <= _zz_912_;
      end
      if(_zz_869_)begin
        int_reg_array_12_22_real <= _zz_912_;
      end
      if(_zz_870_)begin
        int_reg_array_12_23_real <= _zz_912_;
      end
      if(_zz_871_)begin
        int_reg_array_12_24_real <= _zz_912_;
      end
      if(_zz_872_)begin
        int_reg_array_12_25_real <= _zz_912_;
      end
      if(_zz_873_)begin
        int_reg_array_12_26_real <= _zz_912_;
      end
      if(_zz_874_)begin
        int_reg_array_12_27_real <= _zz_912_;
      end
      if(_zz_875_)begin
        int_reg_array_12_28_real <= _zz_912_;
      end
      if(_zz_876_)begin
        int_reg_array_12_29_real <= _zz_912_;
      end
      if(_zz_877_)begin
        int_reg_array_12_30_real <= _zz_912_;
      end
      if(_zz_878_)begin
        int_reg_array_12_31_real <= _zz_912_;
      end
      if(_zz_879_)begin
        int_reg_array_12_32_real <= _zz_912_;
      end
      if(_zz_880_)begin
        int_reg_array_12_33_real <= _zz_912_;
      end
      if(_zz_881_)begin
        int_reg_array_12_34_real <= _zz_912_;
      end
      if(_zz_882_)begin
        int_reg_array_12_35_real <= _zz_912_;
      end
      if(_zz_883_)begin
        int_reg_array_12_36_real <= _zz_912_;
      end
      if(_zz_884_)begin
        int_reg_array_12_37_real <= _zz_912_;
      end
      if(_zz_885_)begin
        int_reg_array_12_38_real <= _zz_912_;
      end
      if(_zz_886_)begin
        int_reg_array_12_39_real <= _zz_912_;
      end
      if(_zz_887_)begin
        int_reg_array_12_40_real <= _zz_912_;
      end
      if(_zz_888_)begin
        int_reg_array_12_41_real <= _zz_912_;
      end
      if(_zz_889_)begin
        int_reg_array_12_42_real <= _zz_912_;
      end
      if(_zz_890_)begin
        int_reg_array_12_43_real <= _zz_912_;
      end
      if(_zz_891_)begin
        int_reg_array_12_44_real <= _zz_912_;
      end
      if(_zz_892_)begin
        int_reg_array_12_45_real <= _zz_912_;
      end
      if(_zz_893_)begin
        int_reg_array_12_46_real <= _zz_912_;
      end
      if(_zz_894_)begin
        int_reg_array_12_47_real <= _zz_912_;
      end
      if(_zz_895_)begin
        int_reg_array_12_48_real <= _zz_912_;
      end
      if(_zz_896_)begin
        int_reg_array_12_49_real <= _zz_912_;
      end
      if(_zz_897_)begin
        int_reg_array_12_50_real <= _zz_912_;
      end
      if(_zz_898_)begin
        int_reg_array_12_51_real <= _zz_912_;
      end
      if(_zz_899_)begin
        int_reg_array_12_52_real <= _zz_912_;
      end
      if(_zz_900_)begin
        int_reg_array_12_53_real <= _zz_912_;
      end
      if(_zz_901_)begin
        int_reg_array_12_54_real <= _zz_912_;
      end
      if(_zz_902_)begin
        int_reg_array_12_55_real <= _zz_912_;
      end
      if(_zz_903_)begin
        int_reg_array_12_56_real <= _zz_912_;
      end
      if(_zz_904_)begin
        int_reg_array_12_57_real <= _zz_912_;
      end
      if(_zz_905_)begin
        int_reg_array_12_58_real <= _zz_912_;
      end
      if(_zz_906_)begin
        int_reg_array_12_59_real <= _zz_912_;
      end
      if(_zz_907_)begin
        int_reg_array_12_60_real <= _zz_912_;
      end
      if(_zz_908_)begin
        int_reg_array_12_61_real <= _zz_912_;
      end
      if(_zz_909_)begin
        int_reg_array_12_62_real <= _zz_912_;
      end
      if(_zz_910_)begin
        int_reg_array_12_63_real <= _zz_912_;
      end
      if(_zz_847_)begin
        int_reg_array_12_0_imag <= _zz_913_;
      end
      if(_zz_848_)begin
        int_reg_array_12_1_imag <= _zz_913_;
      end
      if(_zz_849_)begin
        int_reg_array_12_2_imag <= _zz_913_;
      end
      if(_zz_850_)begin
        int_reg_array_12_3_imag <= _zz_913_;
      end
      if(_zz_851_)begin
        int_reg_array_12_4_imag <= _zz_913_;
      end
      if(_zz_852_)begin
        int_reg_array_12_5_imag <= _zz_913_;
      end
      if(_zz_853_)begin
        int_reg_array_12_6_imag <= _zz_913_;
      end
      if(_zz_854_)begin
        int_reg_array_12_7_imag <= _zz_913_;
      end
      if(_zz_855_)begin
        int_reg_array_12_8_imag <= _zz_913_;
      end
      if(_zz_856_)begin
        int_reg_array_12_9_imag <= _zz_913_;
      end
      if(_zz_857_)begin
        int_reg_array_12_10_imag <= _zz_913_;
      end
      if(_zz_858_)begin
        int_reg_array_12_11_imag <= _zz_913_;
      end
      if(_zz_859_)begin
        int_reg_array_12_12_imag <= _zz_913_;
      end
      if(_zz_860_)begin
        int_reg_array_12_13_imag <= _zz_913_;
      end
      if(_zz_861_)begin
        int_reg_array_12_14_imag <= _zz_913_;
      end
      if(_zz_862_)begin
        int_reg_array_12_15_imag <= _zz_913_;
      end
      if(_zz_863_)begin
        int_reg_array_12_16_imag <= _zz_913_;
      end
      if(_zz_864_)begin
        int_reg_array_12_17_imag <= _zz_913_;
      end
      if(_zz_865_)begin
        int_reg_array_12_18_imag <= _zz_913_;
      end
      if(_zz_866_)begin
        int_reg_array_12_19_imag <= _zz_913_;
      end
      if(_zz_867_)begin
        int_reg_array_12_20_imag <= _zz_913_;
      end
      if(_zz_868_)begin
        int_reg_array_12_21_imag <= _zz_913_;
      end
      if(_zz_869_)begin
        int_reg_array_12_22_imag <= _zz_913_;
      end
      if(_zz_870_)begin
        int_reg_array_12_23_imag <= _zz_913_;
      end
      if(_zz_871_)begin
        int_reg_array_12_24_imag <= _zz_913_;
      end
      if(_zz_872_)begin
        int_reg_array_12_25_imag <= _zz_913_;
      end
      if(_zz_873_)begin
        int_reg_array_12_26_imag <= _zz_913_;
      end
      if(_zz_874_)begin
        int_reg_array_12_27_imag <= _zz_913_;
      end
      if(_zz_875_)begin
        int_reg_array_12_28_imag <= _zz_913_;
      end
      if(_zz_876_)begin
        int_reg_array_12_29_imag <= _zz_913_;
      end
      if(_zz_877_)begin
        int_reg_array_12_30_imag <= _zz_913_;
      end
      if(_zz_878_)begin
        int_reg_array_12_31_imag <= _zz_913_;
      end
      if(_zz_879_)begin
        int_reg_array_12_32_imag <= _zz_913_;
      end
      if(_zz_880_)begin
        int_reg_array_12_33_imag <= _zz_913_;
      end
      if(_zz_881_)begin
        int_reg_array_12_34_imag <= _zz_913_;
      end
      if(_zz_882_)begin
        int_reg_array_12_35_imag <= _zz_913_;
      end
      if(_zz_883_)begin
        int_reg_array_12_36_imag <= _zz_913_;
      end
      if(_zz_884_)begin
        int_reg_array_12_37_imag <= _zz_913_;
      end
      if(_zz_885_)begin
        int_reg_array_12_38_imag <= _zz_913_;
      end
      if(_zz_886_)begin
        int_reg_array_12_39_imag <= _zz_913_;
      end
      if(_zz_887_)begin
        int_reg_array_12_40_imag <= _zz_913_;
      end
      if(_zz_888_)begin
        int_reg_array_12_41_imag <= _zz_913_;
      end
      if(_zz_889_)begin
        int_reg_array_12_42_imag <= _zz_913_;
      end
      if(_zz_890_)begin
        int_reg_array_12_43_imag <= _zz_913_;
      end
      if(_zz_891_)begin
        int_reg_array_12_44_imag <= _zz_913_;
      end
      if(_zz_892_)begin
        int_reg_array_12_45_imag <= _zz_913_;
      end
      if(_zz_893_)begin
        int_reg_array_12_46_imag <= _zz_913_;
      end
      if(_zz_894_)begin
        int_reg_array_12_47_imag <= _zz_913_;
      end
      if(_zz_895_)begin
        int_reg_array_12_48_imag <= _zz_913_;
      end
      if(_zz_896_)begin
        int_reg_array_12_49_imag <= _zz_913_;
      end
      if(_zz_897_)begin
        int_reg_array_12_50_imag <= _zz_913_;
      end
      if(_zz_898_)begin
        int_reg_array_12_51_imag <= _zz_913_;
      end
      if(_zz_899_)begin
        int_reg_array_12_52_imag <= _zz_913_;
      end
      if(_zz_900_)begin
        int_reg_array_12_53_imag <= _zz_913_;
      end
      if(_zz_901_)begin
        int_reg_array_12_54_imag <= _zz_913_;
      end
      if(_zz_902_)begin
        int_reg_array_12_55_imag <= _zz_913_;
      end
      if(_zz_903_)begin
        int_reg_array_12_56_imag <= _zz_913_;
      end
      if(_zz_904_)begin
        int_reg_array_12_57_imag <= _zz_913_;
      end
      if(_zz_905_)begin
        int_reg_array_12_58_imag <= _zz_913_;
      end
      if(_zz_906_)begin
        int_reg_array_12_59_imag <= _zz_913_;
      end
      if(_zz_907_)begin
        int_reg_array_12_60_imag <= _zz_913_;
      end
      if(_zz_908_)begin
        int_reg_array_12_61_imag <= _zz_913_;
      end
      if(_zz_909_)begin
        int_reg_array_12_62_imag <= _zz_913_;
      end
      if(_zz_910_)begin
        int_reg_array_12_63_imag <= _zz_913_;
      end
      if(_zz_916_)begin
        int_reg_array_13_0_real <= _zz_981_;
      end
      if(_zz_917_)begin
        int_reg_array_13_1_real <= _zz_981_;
      end
      if(_zz_918_)begin
        int_reg_array_13_2_real <= _zz_981_;
      end
      if(_zz_919_)begin
        int_reg_array_13_3_real <= _zz_981_;
      end
      if(_zz_920_)begin
        int_reg_array_13_4_real <= _zz_981_;
      end
      if(_zz_921_)begin
        int_reg_array_13_5_real <= _zz_981_;
      end
      if(_zz_922_)begin
        int_reg_array_13_6_real <= _zz_981_;
      end
      if(_zz_923_)begin
        int_reg_array_13_7_real <= _zz_981_;
      end
      if(_zz_924_)begin
        int_reg_array_13_8_real <= _zz_981_;
      end
      if(_zz_925_)begin
        int_reg_array_13_9_real <= _zz_981_;
      end
      if(_zz_926_)begin
        int_reg_array_13_10_real <= _zz_981_;
      end
      if(_zz_927_)begin
        int_reg_array_13_11_real <= _zz_981_;
      end
      if(_zz_928_)begin
        int_reg_array_13_12_real <= _zz_981_;
      end
      if(_zz_929_)begin
        int_reg_array_13_13_real <= _zz_981_;
      end
      if(_zz_930_)begin
        int_reg_array_13_14_real <= _zz_981_;
      end
      if(_zz_931_)begin
        int_reg_array_13_15_real <= _zz_981_;
      end
      if(_zz_932_)begin
        int_reg_array_13_16_real <= _zz_981_;
      end
      if(_zz_933_)begin
        int_reg_array_13_17_real <= _zz_981_;
      end
      if(_zz_934_)begin
        int_reg_array_13_18_real <= _zz_981_;
      end
      if(_zz_935_)begin
        int_reg_array_13_19_real <= _zz_981_;
      end
      if(_zz_936_)begin
        int_reg_array_13_20_real <= _zz_981_;
      end
      if(_zz_937_)begin
        int_reg_array_13_21_real <= _zz_981_;
      end
      if(_zz_938_)begin
        int_reg_array_13_22_real <= _zz_981_;
      end
      if(_zz_939_)begin
        int_reg_array_13_23_real <= _zz_981_;
      end
      if(_zz_940_)begin
        int_reg_array_13_24_real <= _zz_981_;
      end
      if(_zz_941_)begin
        int_reg_array_13_25_real <= _zz_981_;
      end
      if(_zz_942_)begin
        int_reg_array_13_26_real <= _zz_981_;
      end
      if(_zz_943_)begin
        int_reg_array_13_27_real <= _zz_981_;
      end
      if(_zz_944_)begin
        int_reg_array_13_28_real <= _zz_981_;
      end
      if(_zz_945_)begin
        int_reg_array_13_29_real <= _zz_981_;
      end
      if(_zz_946_)begin
        int_reg_array_13_30_real <= _zz_981_;
      end
      if(_zz_947_)begin
        int_reg_array_13_31_real <= _zz_981_;
      end
      if(_zz_948_)begin
        int_reg_array_13_32_real <= _zz_981_;
      end
      if(_zz_949_)begin
        int_reg_array_13_33_real <= _zz_981_;
      end
      if(_zz_950_)begin
        int_reg_array_13_34_real <= _zz_981_;
      end
      if(_zz_951_)begin
        int_reg_array_13_35_real <= _zz_981_;
      end
      if(_zz_952_)begin
        int_reg_array_13_36_real <= _zz_981_;
      end
      if(_zz_953_)begin
        int_reg_array_13_37_real <= _zz_981_;
      end
      if(_zz_954_)begin
        int_reg_array_13_38_real <= _zz_981_;
      end
      if(_zz_955_)begin
        int_reg_array_13_39_real <= _zz_981_;
      end
      if(_zz_956_)begin
        int_reg_array_13_40_real <= _zz_981_;
      end
      if(_zz_957_)begin
        int_reg_array_13_41_real <= _zz_981_;
      end
      if(_zz_958_)begin
        int_reg_array_13_42_real <= _zz_981_;
      end
      if(_zz_959_)begin
        int_reg_array_13_43_real <= _zz_981_;
      end
      if(_zz_960_)begin
        int_reg_array_13_44_real <= _zz_981_;
      end
      if(_zz_961_)begin
        int_reg_array_13_45_real <= _zz_981_;
      end
      if(_zz_962_)begin
        int_reg_array_13_46_real <= _zz_981_;
      end
      if(_zz_963_)begin
        int_reg_array_13_47_real <= _zz_981_;
      end
      if(_zz_964_)begin
        int_reg_array_13_48_real <= _zz_981_;
      end
      if(_zz_965_)begin
        int_reg_array_13_49_real <= _zz_981_;
      end
      if(_zz_966_)begin
        int_reg_array_13_50_real <= _zz_981_;
      end
      if(_zz_967_)begin
        int_reg_array_13_51_real <= _zz_981_;
      end
      if(_zz_968_)begin
        int_reg_array_13_52_real <= _zz_981_;
      end
      if(_zz_969_)begin
        int_reg_array_13_53_real <= _zz_981_;
      end
      if(_zz_970_)begin
        int_reg_array_13_54_real <= _zz_981_;
      end
      if(_zz_971_)begin
        int_reg_array_13_55_real <= _zz_981_;
      end
      if(_zz_972_)begin
        int_reg_array_13_56_real <= _zz_981_;
      end
      if(_zz_973_)begin
        int_reg_array_13_57_real <= _zz_981_;
      end
      if(_zz_974_)begin
        int_reg_array_13_58_real <= _zz_981_;
      end
      if(_zz_975_)begin
        int_reg_array_13_59_real <= _zz_981_;
      end
      if(_zz_976_)begin
        int_reg_array_13_60_real <= _zz_981_;
      end
      if(_zz_977_)begin
        int_reg_array_13_61_real <= _zz_981_;
      end
      if(_zz_978_)begin
        int_reg_array_13_62_real <= _zz_981_;
      end
      if(_zz_979_)begin
        int_reg_array_13_63_real <= _zz_981_;
      end
      if(_zz_916_)begin
        int_reg_array_13_0_imag <= _zz_982_;
      end
      if(_zz_917_)begin
        int_reg_array_13_1_imag <= _zz_982_;
      end
      if(_zz_918_)begin
        int_reg_array_13_2_imag <= _zz_982_;
      end
      if(_zz_919_)begin
        int_reg_array_13_3_imag <= _zz_982_;
      end
      if(_zz_920_)begin
        int_reg_array_13_4_imag <= _zz_982_;
      end
      if(_zz_921_)begin
        int_reg_array_13_5_imag <= _zz_982_;
      end
      if(_zz_922_)begin
        int_reg_array_13_6_imag <= _zz_982_;
      end
      if(_zz_923_)begin
        int_reg_array_13_7_imag <= _zz_982_;
      end
      if(_zz_924_)begin
        int_reg_array_13_8_imag <= _zz_982_;
      end
      if(_zz_925_)begin
        int_reg_array_13_9_imag <= _zz_982_;
      end
      if(_zz_926_)begin
        int_reg_array_13_10_imag <= _zz_982_;
      end
      if(_zz_927_)begin
        int_reg_array_13_11_imag <= _zz_982_;
      end
      if(_zz_928_)begin
        int_reg_array_13_12_imag <= _zz_982_;
      end
      if(_zz_929_)begin
        int_reg_array_13_13_imag <= _zz_982_;
      end
      if(_zz_930_)begin
        int_reg_array_13_14_imag <= _zz_982_;
      end
      if(_zz_931_)begin
        int_reg_array_13_15_imag <= _zz_982_;
      end
      if(_zz_932_)begin
        int_reg_array_13_16_imag <= _zz_982_;
      end
      if(_zz_933_)begin
        int_reg_array_13_17_imag <= _zz_982_;
      end
      if(_zz_934_)begin
        int_reg_array_13_18_imag <= _zz_982_;
      end
      if(_zz_935_)begin
        int_reg_array_13_19_imag <= _zz_982_;
      end
      if(_zz_936_)begin
        int_reg_array_13_20_imag <= _zz_982_;
      end
      if(_zz_937_)begin
        int_reg_array_13_21_imag <= _zz_982_;
      end
      if(_zz_938_)begin
        int_reg_array_13_22_imag <= _zz_982_;
      end
      if(_zz_939_)begin
        int_reg_array_13_23_imag <= _zz_982_;
      end
      if(_zz_940_)begin
        int_reg_array_13_24_imag <= _zz_982_;
      end
      if(_zz_941_)begin
        int_reg_array_13_25_imag <= _zz_982_;
      end
      if(_zz_942_)begin
        int_reg_array_13_26_imag <= _zz_982_;
      end
      if(_zz_943_)begin
        int_reg_array_13_27_imag <= _zz_982_;
      end
      if(_zz_944_)begin
        int_reg_array_13_28_imag <= _zz_982_;
      end
      if(_zz_945_)begin
        int_reg_array_13_29_imag <= _zz_982_;
      end
      if(_zz_946_)begin
        int_reg_array_13_30_imag <= _zz_982_;
      end
      if(_zz_947_)begin
        int_reg_array_13_31_imag <= _zz_982_;
      end
      if(_zz_948_)begin
        int_reg_array_13_32_imag <= _zz_982_;
      end
      if(_zz_949_)begin
        int_reg_array_13_33_imag <= _zz_982_;
      end
      if(_zz_950_)begin
        int_reg_array_13_34_imag <= _zz_982_;
      end
      if(_zz_951_)begin
        int_reg_array_13_35_imag <= _zz_982_;
      end
      if(_zz_952_)begin
        int_reg_array_13_36_imag <= _zz_982_;
      end
      if(_zz_953_)begin
        int_reg_array_13_37_imag <= _zz_982_;
      end
      if(_zz_954_)begin
        int_reg_array_13_38_imag <= _zz_982_;
      end
      if(_zz_955_)begin
        int_reg_array_13_39_imag <= _zz_982_;
      end
      if(_zz_956_)begin
        int_reg_array_13_40_imag <= _zz_982_;
      end
      if(_zz_957_)begin
        int_reg_array_13_41_imag <= _zz_982_;
      end
      if(_zz_958_)begin
        int_reg_array_13_42_imag <= _zz_982_;
      end
      if(_zz_959_)begin
        int_reg_array_13_43_imag <= _zz_982_;
      end
      if(_zz_960_)begin
        int_reg_array_13_44_imag <= _zz_982_;
      end
      if(_zz_961_)begin
        int_reg_array_13_45_imag <= _zz_982_;
      end
      if(_zz_962_)begin
        int_reg_array_13_46_imag <= _zz_982_;
      end
      if(_zz_963_)begin
        int_reg_array_13_47_imag <= _zz_982_;
      end
      if(_zz_964_)begin
        int_reg_array_13_48_imag <= _zz_982_;
      end
      if(_zz_965_)begin
        int_reg_array_13_49_imag <= _zz_982_;
      end
      if(_zz_966_)begin
        int_reg_array_13_50_imag <= _zz_982_;
      end
      if(_zz_967_)begin
        int_reg_array_13_51_imag <= _zz_982_;
      end
      if(_zz_968_)begin
        int_reg_array_13_52_imag <= _zz_982_;
      end
      if(_zz_969_)begin
        int_reg_array_13_53_imag <= _zz_982_;
      end
      if(_zz_970_)begin
        int_reg_array_13_54_imag <= _zz_982_;
      end
      if(_zz_971_)begin
        int_reg_array_13_55_imag <= _zz_982_;
      end
      if(_zz_972_)begin
        int_reg_array_13_56_imag <= _zz_982_;
      end
      if(_zz_973_)begin
        int_reg_array_13_57_imag <= _zz_982_;
      end
      if(_zz_974_)begin
        int_reg_array_13_58_imag <= _zz_982_;
      end
      if(_zz_975_)begin
        int_reg_array_13_59_imag <= _zz_982_;
      end
      if(_zz_976_)begin
        int_reg_array_13_60_imag <= _zz_982_;
      end
      if(_zz_977_)begin
        int_reg_array_13_61_imag <= _zz_982_;
      end
      if(_zz_978_)begin
        int_reg_array_13_62_imag <= _zz_982_;
      end
      if(_zz_979_)begin
        int_reg_array_13_63_imag <= _zz_982_;
      end
      if(_zz_985_)begin
        int_reg_array_14_0_real <= _zz_1050_;
      end
      if(_zz_986_)begin
        int_reg_array_14_1_real <= _zz_1050_;
      end
      if(_zz_987_)begin
        int_reg_array_14_2_real <= _zz_1050_;
      end
      if(_zz_988_)begin
        int_reg_array_14_3_real <= _zz_1050_;
      end
      if(_zz_989_)begin
        int_reg_array_14_4_real <= _zz_1050_;
      end
      if(_zz_990_)begin
        int_reg_array_14_5_real <= _zz_1050_;
      end
      if(_zz_991_)begin
        int_reg_array_14_6_real <= _zz_1050_;
      end
      if(_zz_992_)begin
        int_reg_array_14_7_real <= _zz_1050_;
      end
      if(_zz_993_)begin
        int_reg_array_14_8_real <= _zz_1050_;
      end
      if(_zz_994_)begin
        int_reg_array_14_9_real <= _zz_1050_;
      end
      if(_zz_995_)begin
        int_reg_array_14_10_real <= _zz_1050_;
      end
      if(_zz_996_)begin
        int_reg_array_14_11_real <= _zz_1050_;
      end
      if(_zz_997_)begin
        int_reg_array_14_12_real <= _zz_1050_;
      end
      if(_zz_998_)begin
        int_reg_array_14_13_real <= _zz_1050_;
      end
      if(_zz_999_)begin
        int_reg_array_14_14_real <= _zz_1050_;
      end
      if(_zz_1000_)begin
        int_reg_array_14_15_real <= _zz_1050_;
      end
      if(_zz_1001_)begin
        int_reg_array_14_16_real <= _zz_1050_;
      end
      if(_zz_1002_)begin
        int_reg_array_14_17_real <= _zz_1050_;
      end
      if(_zz_1003_)begin
        int_reg_array_14_18_real <= _zz_1050_;
      end
      if(_zz_1004_)begin
        int_reg_array_14_19_real <= _zz_1050_;
      end
      if(_zz_1005_)begin
        int_reg_array_14_20_real <= _zz_1050_;
      end
      if(_zz_1006_)begin
        int_reg_array_14_21_real <= _zz_1050_;
      end
      if(_zz_1007_)begin
        int_reg_array_14_22_real <= _zz_1050_;
      end
      if(_zz_1008_)begin
        int_reg_array_14_23_real <= _zz_1050_;
      end
      if(_zz_1009_)begin
        int_reg_array_14_24_real <= _zz_1050_;
      end
      if(_zz_1010_)begin
        int_reg_array_14_25_real <= _zz_1050_;
      end
      if(_zz_1011_)begin
        int_reg_array_14_26_real <= _zz_1050_;
      end
      if(_zz_1012_)begin
        int_reg_array_14_27_real <= _zz_1050_;
      end
      if(_zz_1013_)begin
        int_reg_array_14_28_real <= _zz_1050_;
      end
      if(_zz_1014_)begin
        int_reg_array_14_29_real <= _zz_1050_;
      end
      if(_zz_1015_)begin
        int_reg_array_14_30_real <= _zz_1050_;
      end
      if(_zz_1016_)begin
        int_reg_array_14_31_real <= _zz_1050_;
      end
      if(_zz_1017_)begin
        int_reg_array_14_32_real <= _zz_1050_;
      end
      if(_zz_1018_)begin
        int_reg_array_14_33_real <= _zz_1050_;
      end
      if(_zz_1019_)begin
        int_reg_array_14_34_real <= _zz_1050_;
      end
      if(_zz_1020_)begin
        int_reg_array_14_35_real <= _zz_1050_;
      end
      if(_zz_1021_)begin
        int_reg_array_14_36_real <= _zz_1050_;
      end
      if(_zz_1022_)begin
        int_reg_array_14_37_real <= _zz_1050_;
      end
      if(_zz_1023_)begin
        int_reg_array_14_38_real <= _zz_1050_;
      end
      if(_zz_1024_)begin
        int_reg_array_14_39_real <= _zz_1050_;
      end
      if(_zz_1025_)begin
        int_reg_array_14_40_real <= _zz_1050_;
      end
      if(_zz_1026_)begin
        int_reg_array_14_41_real <= _zz_1050_;
      end
      if(_zz_1027_)begin
        int_reg_array_14_42_real <= _zz_1050_;
      end
      if(_zz_1028_)begin
        int_reg_array_14_43_real <= _zz_1050_;
      end
      if(_zz_1029_)begin
        int_reg_array_14_44_real <= _zz_1050_;
      end
      if(_zz_1030_)begin
        int_reg_array_14_45_real <= _zz_1050_;
      end
      if(_zz_1031_)begin
        int_reg_array_14_46_real <= _zz_1050_;
      end
      if(_zz_1032_)begin
        int_reg_array_14_47_real <= _zz_1050_;
      end
      if(_zz_1033_)begin
        int_reg_array_14_48_real <= _zz_1050_;
      end
      if(_zz_1034_)begin
        int_reg_array_14_49_real <= _zz_1050_;
      end
      if(_zz_1035_)begin
        int_reg_array_14_50_real <= _zz_1050_;
      end
      if(_zz_1036_)begin
        int_reg_array_14_51_real <= _zz_1050_;
      end
      if(_zz_1037_)begin
        int_reg_array_14_52_real <= _zz_1050_;
      end
      if(_zz_1038_)begin
        int_reg_array_14_53_real <= _zz_1050_;
      end
      if(_zz_1039_)begin
        int_reg_array_14_54_real <= _zz_1050_;
      end
      if(_zz_1040_)begin
        int_reg_array_14_55_real <= _zz_1050_;
      end
      if(_zz_1041_)begin
        int_reg_array_14_56_real <= _zz_1050_;
      end
      if(_zz_1042_)begin
        int_reg_array_14_57_real <= _zz_1050_;
      end
      if(_zz_1043_)begin
        int_reg_array_14_58_real <= _zz_1050_;
      end
      if(_zz_1044_)begin
        int_reg_array_14_59_real <= _zz_1050_;
      end
      if(_zz_1045_)begin
        int_reg_array_14_60_real <= _zz_1050_;
      end
      if(_zz_1046_)begin
        int_reg_array_14_61_real <= _zz_1050_;
      end
      if(_zz_1047_)begin
        int_reg_array_14_62_real <= _zz_1050_;
      end
      if(_zz_1048_)begin
        int_reg_array_14_63_real <= _zz_1050_;
      end
      if(_zz_985_)begin
        int_reg_array_14_0_imag <= _zz_1051_;
      end
      if(_zz_986_)begin
        int_reg_array_14_1_imag <= _zz_1051_;
      end
      if(_zz_987_)begin
        int_reg_array_14_2_imag <= _zz_1051_;
      end
      if(_zz_988_)begin
        int_reg_array_14_3_imag <= _zz_1051_;
      end
      if(_zz_989_)begin
        int_reg_array_14_4_imag <= _zz_1051_;
      end
      if(_zz_990_)begin
        int_reg_array_14_5_imag <= _zz_1051_;
      end
      if(_zz_991_)begin
        int_reg_array_14_6_imag <= _zz_1051_;
      end
      if(_zz_992_)begin
        int_reg_array_14_7_imag <= _zz_1051_;
      end
      if(_zz_993_)begin
        int_reg_array_14_8_imag <= _zz_1051_;
      end
      if(_zz_994_)begin
        int_reg_array_14_9_imag <= _zz_1051_;
      end
      if(_zz_995_)begin
        int_reg_array_14_10_imag <= _zz_1051_;
      end
      if(_zz_996_)begin
        int_reg_array_14_11_imag <= _zz_1051_;
      end
      if(_zz_997_)begin
        int_reg_array_14_12_imag <= _zz_1051_;
      end
      if(_zz_998_)begin
        int_reg_array_14_13_imag <= _zz_1051_;
      end
      if(_zz_999_)begin
        int_reg_array_14_14_imag <= _zz_1051_;
      end
      if(_zz_1000_)begin
        int_reg_array_14_15_imag <= _zz_1051_;
      end
      if(_zz_1001_)begin
        int_reg_array_14_16_imag <= _zz_1051_;
      end
      if(_zz_1002_)begin
        int_reg_array_14_17_imag <= _zz_1051_;
      end
      if(_zz_1003_)begin
        int_reg_array_14_18_imag <= _zz_1051_;
      end
      if(_zz_1004_)begin
        int_reg_array_14_19_imag <= _zz_1051_;
      end
      if(_zz_1005_)begin
        int_reg_array_14_20_imag <= _zz_1051_;
      end
      if(_zz_1006_)begin
        int_reg_array_14_21_imag <= _zz_1051_;
      end
      if(_zz_1007_)begin
        int_reg_array_14_22_imag <= _zz_1051_;
      end
      if(_zz_1008_)begin
        int_reg_array_14_23_imag <= _zz_1051_;
      end
      if(_zz_1009_)begin
        int_reg_array_14_24_imag <= _zz_1051_;
      end
      if(_zz_1010_)begin
        int_reg_array_14_25_imag <= _zz_1051_;
      end
      if(_zz_1011_)begin
        int_reg_array_14_26_imag <= _zz_1051_;
      end
      if(_zz_1012_)begin
        int_reg_array_14_27_imag <= _zz_1051_;
      end
      if(_zz_1013_)begin
        int_reg_array_14_28_imag <= _zz_1051_;
      end
      if(_zz_1014_)begin
        int_reg_array_14_29_imag <= _zz_1051_;
      end
      if(_zz_1015_)begin
        int_reg_array_14_30_imag <= _zz_1051_;
      end
      if(_zz_1016_)begin
        int_reg_array_14_31_imag <= _zz_1051_;
      end
      if(_zz_1017_)begin
        int_reg_array_14_32_imag <= _zz_1051_;
      end
      if(_zz_1018_)begin
        int_reg_array_14_33_imag <= _zz_1051_;
      end
      if(_zz_1019_)begin
        int_reg_array_14_34_imag <= _zz_1051_;
      end
      if(_zz_1020_)begin
        int_reg_array_14_35_imag <= _zz_1051_;
      end
      if(_zz_1021_)begin
        int_reg_array_14_36_imag <= _zz_1051_;
      end
      if(_zz_1022_)begin
        int_reg_array_14_37_imag <= _zz_1051_;
      end
      if(_zz_1023_)begin
        int_reg_array_14_38_imag <= _zz_1051_;
      end
      if(_zz_1024_)begin
        int_reg_array_14_39_imag <= _zz_1051_;
      end
      if(_zz_1025_)begin
        int_reg_array_14_40_imag <= _zz_1051_;
      end
      if(_zz_1026_)begin
        int_reg_array_14_41_imag <= _zz_1051_;
      end
      if(_zz_1027_)begin
        int_reg_array_14_42_imag <= _zz_1051_;
      end
      if(_zz_1028_)begin
        int_reg_array_14_43_imag <= _zz_1051_;
      end
      if(_zz_1029_)begin
        int_reg_array_14_44_imag <= _zz_1051_;
      end
      if(_zz_1030_)begin
        int_reg_array_14_45_imag <= _zz_1051_;
      end
      if(_zz_1031_)begin
        int_reg_array_14_46_imag <= _zz_1051_;
      end
      if(_zz_1032_)begin
        int_reg_array_14_47_imag <= _zz_1051_;
      end
      if(_zz_1033_)begin
        int_reg_array_14_48_imag <= _zz_1051_;
      end
      if(_zz_1034_)begin
        int_reg_array_14_49_imag <= _zz_1051_;
      end
      if(_zz_1035_)begin
        int_reg_array_14_50_imag <= _zz_1051_;
      end
      if(_zz_1036_)begin
        int_reg_array_14_51_imag <= _zz_1051_;
      end
      if(_zz_1037_)begin
        int_reg_array_14_52_imag <= _zz_1051_;
      end
      if(_zz_1038_)begin
        int_reg_array_14_53_imag <= _zz_1051_;
      end
      if(_zz_1039_)begin
        int_reg_array_14_54_imag <= _zz_1051_;
      end
      if(_zz_1040_)begin
        int_reg_array_14_55_imag <= _zz_1051_;
      end
      if(_zz_1041_)begin
        int_reg_array_14_56_imag <= _zz_1051_;
      end
      if(_zz_1042_)begin
        int_reg_array_14_57_imag <= _zz_1051_;
      end
      if(_zz_1043_)begin
        int_reg_array_14_58_imag <= _zz_1051_;
      end
      if(_zz_1044_)begin
        int_reg_array_14_59_imag <= _zz_1051_;
      end
      if(_zz_1045_)begin
        int_reg_array_14_60_imag <= _zz_1051_;
      end
      if(_zz_1046_)begin
        int_reg_array_14_61_imag <= _zz_1051_;
      end
      if(_zz_1047_)begin
        int_reg_array_14_62_imag <= _zz_1051_;
      end
      if(_zz_1048_)begin
        int_reg_array_14_63_imag <= _zz_1051_;
      end
      if(_zz_1054_)begin
        int_reg_array_15_0_real <= _zz_1119_;
      end
      if(_zz_1055_)begin
        int_reg_array_15_1_real <= _zz_1119_;
      end
      if(_zz_1056_)begin
        int_reg_array_15_2_real <= _zz_1119_;
      end
      if(_zz_1057_)begin
        int_reg_array_15_3_real <= _zz_1119_;
      end
      if(_zz_1058_)begin
        int_reg_array_15_4_real <= _zz_1119_;
      end
      if(_zz_1059_)begin
        int_reg_array_15_5_real <= _zz_1119_;
      end
      if(_zz_1060_)begin
        int_reg_array_15_6_real <= _zz_1119_;
      end
      if(_zz_1061_)begin
        int_reg_array_15_7_real <= _zz_1119_;
      end
      if(_zz_1062_)begin
        int_reg_array_15_8_real <= _zz_1119_;
      end
      if(_zz_1063_)begin
        int_reg_array_15_9_real <= _zz_1119_;
      end
      if(_zz_1064_)begin
        int_reg_array_15_10_real <= _zz_1119_;
      end
      if(_zz_1065_)begin
        int_reg_array_15_11_real <= _zz_1119_;
      end
      if(_zz_1066_)begin
        int_reg_array_15_12_real <= _zz_1119_;
      end
      if(_zz_1067_)begin
        int_reg_array_15_13_real <= _zz_1119_;
      end
      if(_zz_1068_)begin
        int_reg_array_15_14_real <= _zz_1119_;
      end
      if(_zz_1069_)begin
        int_reg_array_15_15_real <= _zz_1119_;
      end
      if(_zz_1070_)begin
        int_reg_array_15_16_real <= _zz_1119_;
      end
      if(_zz_1071_)begin
        int_reg_array_15_17_real <= _zz_1119_;
      end
      if(_zz_1072_)begin
        int_reg_array_15_18_real <= _zz_1119_;
      end
      if(_zz_1073_)begin
        int_reg_array_15_19_real <= _zz_1119_;
      end
      if(_zz_1074_)begin
        int_reg_array_15_20_real <= _zz_1119_;
      end
      if(_zz_1075_)begin
        int_reg_array_15_21_real <= _zz_1119_;
      end
      if(_zz_1076_)begin
        int_reg_array_15_22_real <= _zz_1119_;
      end
      if(_zz_1077_)begin
        int_reg_array_15_23_real <= _zz_1119_;
      end
      if(_zz_1078_)begin
        int_reg_array_15_24_real <= _zz_1119_;
      end
      if(_zz_1079_)begin
        int_reg_array_15_25_real <= _zz_1119_;
      end
      if(_zz_1080_)begin
        int_reg_array_15_26_real <= _zz_1119_;
      end
      if(_zz_1081_)begin
        int_reg_array_15_27_real <= _zz_1119_;
      end
      if(_zz_1082_)begin
        int_reg_array_15_28_real <= _zz_1119_;
      end
      if(_zz_1083_)begin
        int_reg_array_15_29_real <= _zz_1119_;
      end
      if(_zz_1084_)begin
        int_reg_array_15_30_real <= _zz_1119_;
      end
      if(_zz_1085_)begin
        int_reg_array_15_31_real <= _zz_1119_;
      end
      if(_zz_1086_)begin
        int_reg_array_15_32_real <= _zz_1119_;
      end
      if(_zz_1087_)begin
        int_reg_array_15_33_real <= _zz_1119_;
      end
      if(_zz_1088_)begin
        int_reg_array_15_34_real <= _zz_1119_;
      end
      if(_zz_1089_)begin
        int_reg_array_15_35_real <= _zz_1119_;
      end
      if(_zz_1090_)begin
        int_reg_array_15_36_real <= _zz_1119_;
      end
      if(_zz_1091_)begin
        int_reg_array_15_37_real <= _zz_1119_;
      end
      if(_zz_1092_)begin
        int_reg_array_15_38_real <= _zz_1119_;
      end
      if(_zz_1093_)begin
        int_reg_array_15_39_real <= _zz_1119_;
      end
      if(_zz_1094_)begin
        int_reg_array_15_40_real <= _zz_1119_;
      end
      if(_zz_1095_)begin
        int_reg_array_15_41_real <= _zz_1119_;
      end
      if(_zz_1096_)begin
        int_reg_array_15_42_real <= _zz_1119_;
      end
      if(_zz_1097_)begin
        int_reg_array_15_43_real <= _zz_1119_;
      end
      if(_zz_1098_)begin
        int_reg_array_15_44_real <= _zz_1119_;
      end
      if(_zz_1099_)begin
        int_reg_array_15_45_real <= _zz_1119_;
      end
      if(_zz_1100_)begin
        int_reg_array_15_46_real <= _zz_1119_;
      end
      if(_zz_1101_)begin
        int_reg_array_15_47_real <= _zz_1119_;
      end
      if(_zz_1102_)begin
        int_reg_array_15_48_real <= _zz_1119_;
      end
      if(_zz_1103_)begin
        int_reg_array_15_49_real <= _zz_1119_;
      end
      if(_zz_1104_)begin
        int_reg_array_15_50_real <= _zz_1119_;
      end
      if(_zz_1105_)begin
        int_reg_array_15_51_real <= _zz_1119_;
      end
      if(_zz_1106_)begin
        int_reg_array_15_52_real <= _zz_1119_;
      end
      if(_zz_1107_)begin
        int_reg_array_15_53_real <= _zz_1119_;
      end
      if(_zz_1108_)begin
        int_reg_array_15_54_real <= _zz_1119_;
      end
      if(_zz_1109_)begin
        int_reg_array_15_55_real <= _zz_1119_;
      end
      if(_zz_1110_)begin
        int_reg_array_15_56_real <= _zz_1119_;
      end
      if(_zz_1111_)begin
        int_reg_array_15_57_real <= _zz_1119_;
      end
      if(_zz_1112_)begin
        int_reg_array_15_58_real <= _zz_1119_;
      end
      if(_zz_1113_)begin
        int_reg_array_15_59_real <= _zz_1119_;
      end
      if(_zz_1114_)begin
        int_reg_array_15_60_real <= _zz_1119_;
      end
      if(_zz_1115_)begin
        int_reg_array_15_61_real <= _zz_1119_;
      end
      if(_zz_1116_)begin
        int_reg_array_15_62_real <= _zz_1119_;
      end
      if(_zz_1117_)begin
        int_reg_array_15_63_real <= _zz_1119_;
      end
      if(_zz_1054_)begin
        int_reg_array_15_0_imag <= _zz_1120_;
      end
      if(_zz_1055_)begin
        int_reg_array_15_1_imag <= _zz_1120_;
      end
      if(_zz_1056_)begin
        int_reg_array_15_2_imag <= _zz_1120_;
      end
      if(_zz_1057_)begin
        int_reg_array_15_3_imag <= _zz_1120_;
      end
      if(_zz_1058_)begin
        int_reg_array_15_4_imag <= _zz_1120_;
      end
      if(_zz_1059_)begin
        int_reg_array_15_5_imag <= _zz_1120_;
      end
      if(_zz_1060_)begin
        int_reg_array_15_6_imag <= _zz_1120_;
      end
      if(_zz_1061_)begin
        int_reg_array_15_7_imag <= _zz_1120_;
      end
      if(_zz_1062_)begin
        int_reg_array_15_8_imag <= _zz_1120_;
      end
      if(_zz_1063_)begin
        int_reg_array_15_9_imag <= _zz_1120_;
      end
      if(_zz_1064_)begin
        int_reg_array_15_10_imag <= _zz_1120_;
      end
      if(_zz_1065_)begin
        int_reg_array_15_11_imag <= _zz_1120_;
      end
      if(_zz_1066_)begin
        int_reg_array_15_12_imag <= _zz_1120_;
      end
      if(_zz_1067_)begin
        int_reg_array_15_13_imag <= _zz_1120_;
      end
      if(_zz_1068_)begin
        int_reg_array_15_14_imag <= _zz_1120_;
      end
      if(_zz_1069_)begin
        int_reg_array_15_15_imag <= _zz_1120_;
      end
      if(_zz_1070_)begin
        int_reg_array_15_16_imag <= _zz_1120_;
      end
      if(_zz_1071_)begin
        int_reg_array_15_17_imag <= _zz_1120_;
      end
      if(_zz_1072_)begin
        int_reg_array_15_18_imag <= _zz_1120_;
      end
      if(_zz_1073_)begin
        int_reg_array_15_19_imag <= _zz_1120_;
      end
      if(_zz_1074_)begin
        int_reg_array_15_20_imag <= _zz_1120_;
      end
      if(_zz_1075_)begin
        int_reg_array_15_21_imag <= _zz_1120_;
      end
      if(_zz_1076_)begin
        int_reg_array_15_22_imag <= _zz_1120_;
      end
      if(_zz_1077_)begin
        int_reg_array_15_23_imag <= _zz_1120_;
      end
      if(_zz_1078_)begin
        int_reg_array_15_24_imag <= _zz_1120_;
      end
      if(_zz_1079_)begin
        int_reg_array_15_25_imag <= _zz_1120_;
      end
      if(_zz_1080_)begin
        int_reg_array_15_26_imag <= _zz_1120_;
      end
      if(_zz_1081_)begin
        int_reg_array_15_27_imag <= _zz_1120_;
      end
      if(_zz_1082_)begin
        int_reg_array_15_28_imag <= _zz_1120_;
      end
      if(_zz_1083_)begin
        int_reg_array_15_29_imag <= _zz_1120_;
      end
      if(_zz_1084_)begin
        int_reg_array_15_30_imag <= _zz_1120_;
      end
      if(_zz_1085_)begin
        int_reg_array_15_31_imag <= _zz_1120_;
      end
      if(_zz_1086_)begin
        int_reg_array_15_32_imag <= _zz_1120_;
      end
      if(_zz_1087_)begin
        int_reg_array_15_33_imag <= _zz_1120_;
      end
      if(_zz_1088_)begin
        int_reg_array_15_34_imag <= _zz_1120_;
      end
      if(_zz_1089_)begin
        int_reg_array_15_35_imag <= _zz_1120_;
      end
      if(_zz_1090_)begin
        int_reg_array_15_36_imag <= _zz_1120_;
      end
      if(_zz_1091_)begin
        int_reg_array_15_37_imag <= _zz_1120_;
      end
      if(_zz_1092_)begin
        int_reg_array_15_38_imag <= _zz_1120_;
      end
      if(_zz_1093_)begin
        int_reg_array_15_39_imag <= _zz_1120_;
      end
      if(_zz_1094_)begin
        int_reg_array_15_40_imag <= _zz_1120_;
      end
      if(_zz_1095_)begin
        int_reg_array_15_41_imag <= _zz_1120_;
      end
      if(_zz_1096_)begin
        int_reg_array_15_42_imag <= _zz_1120_;
      end
      if(_zz_1097_)begin
        int_reg_array_15_43_imag <= _zz_1120_;
      end
      if(_zz_1098_)begin
        int_reg_array_15_44_imag <= _zz_1120_;
      end
      if(_zz_1099_)begin
        int_reg_array_15_45_imag <= _zz_1120_;
      end
      if(_zz_1100_)begin
        int_reg_array_15_46_imag <= _zz_1120_;
      end
      if(_zz_1101_)begin
        int_reg_array_15_47_imag <= _zz_1120_;
      end
      if(_zz_1102_)begin
        int_reg_array_15_48_imag <= _zz_1120_;
      end
      if(_zz_1103_)begin
        int_reg_array_15_49_imag <= _zz_1120_;
      end
      if(_zz_1104_)begin
        int_reg_array_15_50_imag <= _zz_1120_;
      end
      if(_zz_1105_)begin
        int_reg_array_15_51_imag <= _zz_1120_;
      end
      if(_zz_1106_)begin
        int_reg_array_15_52_imag <= _zz_1120_;
      end
      if(_zz_1107_)begin
        int_reg_array_15_53_imag <= _zz_1120_;
      end
      if(_zz_1108_)begin
        int_reg_array_15_54_imag <= _zz_1120_;
      end
      if(_zz_1109_)begin
        int_reg_array_15_55_imag <= _zz_1120_;
      end
      if(_zz_1110_)begin
        int_reg_array_15_56_imag <= _zz_1120_;
      end
      if(_zz_1111_)begin
        int_reg_array_15_57_imag <= _zz_1120_;
      end
      if(_zz_1112_)begin
        int_reg_array_15_58_imag <= _zz_1120_;
      end
      if(_zz_1113_)begin
        int_reg_array_15_59_imag <= _zz_1120_;
      end
      if(_zz_1114_)begin
        int_reg_array_15_60_imag <= _zz_1120_;
      end
      if(_zz_1115_)begin
        int_reg_array_15_61_imag <= _zz_1120_;
      end
      if(_zz_1116_)begin
        int_reg_array_15_62_imag <= _zz_1120_;
      end
      if(_zz_1117_)begin
        int_reg_array_15_63_imag <= _zz_1120_;
      end
      if(_zz_1123_)begin
        int_reg_array_16_0_real <= _zz_1188_;
      end
      if(_zz_1124_)begin
        int_reg_array_16_1_real <= _zz_1188_;
      end
      if(_zz_1125_)begin
        int_reg_array_16_2_real <= _zz_1188_;
      end
      if(_zz_1126_)begin
        int_reg_array_16_3_real <= _zz_1188_;
      end
      if(_zz_1127_)begin
        int_reg_array_16_4_real <= _zz_1188_;
      end
      if(_zz_1128_)begin
        int_reg_array_16_5_real <= _zz_1188_;
      end
      if(_zz_1129_)begin
        int_reg_array_16_6_real <= _zz_1188_;
      end
      if(_zz_1130_)begin
        int_reg_array_16_7_real <= _zz_1188_;
      end
      if(_zz_1131_)begin
        int_reg_array_16_8_real <= _zz_1188_;
      end
      if(_zz_1132_)begin
        int_reg_array_16_9_real <= _zz_1188_;
      end
      if(_zz_1133_)begin
        int_reg_array_16_10_real <= _zz_1188_;
      end
      if(_zz_1134_)begin
        int_reg_array_16_11_real <= _zz_1188_;
      end
      if(_zz_1135_)begin
        int_reg_array_16_12_real <= _zz_1188_;
      end
      if(_zz_1136_)begin
        int_reg_array_16_13_real <= _zz_1188_;
      end
      if(_zz_1137_)begin
        int_reg_array_16_14_real <= _zz_1188_;
      end
      if(_zz_1138_)begin
        int_reg_array_16_15_real <= _zz_1188_;
      end
      if(_zz_1139_)begin
        int_reg_array_16_16_real <= _zz_1188_;
      end
      if(_zz_1140_)begin
        int_reg_array_16_17_real <= _zz_1188_;
      end
      if(_zz_1141_)begin
        int_reg_array_16_18_real <= _zz_1188_;
      end
      if(_zz_1142_)begin
        int_reg_array_16_19_real <= _zz_1188_;
      end
      if(_zz_1143_)begin
        int_reg_array_16_20_real <= _zz_1188_;
      end
      if(_zz_1144_)begin
        int_reg_array_16_21_real <= _zz_1188_;
      end
      if(_zz_1145_)begin
        int_reg_array_16_22_real <= _zz_1188_;
      end
      if(_zz_1146_)begin
        int_reg_array_16_23_real <= _zz_1188_;
      end
      if(_zz_1147_)begin
        int_reg_array_16_24_real <= _zz_1188_;
      end
      if(_zz_1148_)begin
        int_reg_array_16_25_real <= _zz_1188_;
      end
      if(_zz_1149_)begin
        int_reg_array_16_26_real <= _zz_1188_;
      end
      if(_zz_1150_)begin
        int_reg_array_16_27_real <= _zz_1188_;
      end
      if(_zz_1151_)begin
        int_reg_array_16_28_real <= _zz_1188_;
      end
      if(_zz_1152_)begin
        int_reg_array_16_29_real <= _zz_1188_;
      end
      if(_zz_1153_)begin
        int_reg_array_16_30_real <= _zz_1188_;
      end
      if(_zz_1154_)begin
        int_reg_array_16_31_real <= _zz_1188_;
      end
      if(_zz_1155_)begin
        int_reg_array_16_32_real <= _zz_1188_;
      end
      if(_zz_1156_)begin
        int_reg_array_16_33_real <= _zz_1188_;
      end
      if(_zz_1157_)begin
        int_reg_array_16_34_real <= _zz_1188_;
      end
      if(_zz_1158_)begin
        int_reg_array_16_35_real <= _zz_1188_;
      end
      if(_zz_1159_)begin
        int_reg_array_16_36_real <= _zz_1188_;
      end
      if(_zz_1160_)begin
        int_reg_array_16_37_real <= _zz_1188_;
      end
      if(_zz_1161_)begin
        int_reg_array_16_38_real <= _zz_1188_;
      end
      if(_zz_1162_)begin
        int_reg_array_16_39_real <= _zz_1188_;
      end
      if(_zz_1163_)begin
        int_reg_array_16_40_real <= _zz_1188_;
      end
      if(_zz_1164_)begin
        int_reg_array_16_41_real <= _zz_1188_;
      end
      if(_zz_1165_)begin
        int_reg_array_16_42_real <= _zz_1188_;
      end
      if(_zz_1166_)begin
        int_reg_array_16_43_real <= _zz_1188_;
      end
      if(_zz_1167_)begin
        int_reg_array_16_44_real <= _zz_1188_;
      end
      if(_zz_1168_)begin
        int_reg_array_16_45_real <= _zz_1188_;
      end
      if(_zz_1169_)begin
        int_reg_array_16_46_real <= _zz_1188_;
      end
      if(_zz_1170_)begin
        int_reg_array_16_47_real <= _zz_1188_;
      end
      if(_zz_1171_)begin
        int_reg_array_16_48_real <= _zz_1188_;
      end
      if(_zz_1172_)begin
        int_reg_array_16_49_real <= _zz_1188_;
      end
      if(_zz_1173_)begin
        int_reg_array_16_50_real <= _zz_1188_;
      end
      if(_zz_1174_)begin
        int_reg_array_16_51_real <= _zz_1188_;
      end
      if(_zz_1175_)begin
        int_reg_array_16_52_real <= _zz_1188_;
      end
      if(_zz_1176_)begin
        int_reg_array_16_53_real <= _zz_1188_;
      end
      if(_zz_1177_)begin
        int_reg_array_16_54_real <= _zz_1188_;
      end
      if(_zz_1178_)begin
        int_reg_array_16_55_real <= _zz_1188_;
      end
      if(_zz_1179_)begin
        int_reg_array_16_56_real <= _zz_1188_;
      end
      if(_zz_1180_)begin
        int_reg_array_16_57_real <= _zz_1188_;
      end
      if(_zz_1181_)begin
        int_reg_array_16_58_real <= _zz_1188_;
      end
      if(_zz_1182_)begin
        int_reg_array_16_59_real <= _zz_1188_;
      end
      if(_zz_1183_)begin
        int_reg_array_16_60_real <= _zz_1188_;
      end
      if(_zz_1184_)begin
        int_reg_array_16_61_real <= _zz_1188_;
      end
      if(_zz_1185_)begin
        int_reg_array_16_62_real <= _zz_1188_;
      end
      if(_zz_1186_)begin
        int_reg_array_16_63_real <= _zz_1188_;
      end
      if(_zz_1123_)begin
        int_reg_array_16_0_imag <= _zz_1189_;
      end
      if(_zz_1124_)begin
        int_reg_array_16_1_imag <= _zz_1189_;
      end
      if(_zz_1125_)begin
        int_reg_array_16_2_imag <= _zz_1189_;
      end
      if(_zz_1126_)begin
        int_reg_array_16_3_imag <= _zz_1189_;
      end
      if(_zz_1127_)begin
        int_reg_array_16_4_imag <= _zz_1189_;
      end
      if(_zz_1128_)begin
        int_reg_array_16_5_imag <= _zz_1189_;
      end
      if(_zz_1129_)begin
        int_reg_array_16_6_imag <= _zz_1189_;
      end
      if(_zz_1130_)begin
        int_reg_array_16_7_imag <= _zz_1189_;
      end
      if(_zz_1131_)begin
        int_reg_array_16_8_imag <= _zz_1189_;
      end
      if(_zz_1132_)begin
        int_reg_array_16_9_imag <= _zz_1189_;
      end
      if(_zz_1133_)begin
        int_reg_array_16_10_imag <= _zz_1189_;
      end
      if(_zz_1134_)begin
        int_reg_array_16_11_imag <= _zz_1189_;
      end
      if(_zz_1135_)begin
        int_reg_array_16_12_imag <= _zz_1189_;
      end
      if(_zz_1136_)begin
        int_reg_array_16_13_imag <= _zz_1189_;
      end
      if(_zz_1137_)begin
        int_reg_array_16_14_imag <= _zz_1189_;
      end
      if(_zz_1138_)begin
        int_reg_array_16_15_imag <= _zz_1189_;
      end
      if(_zz_1139_)begin
        int_reg_array_16_16_imag <= _zz_1189_;
      end
      if(_zz_1140_)begin
        int_reg_array_16_17_imag <= _zz_1189_;
      end
      if(_zz_1141_)begin
        int_reg_array_16_18_imag <= _zz_1189_;
      end
      if(_zz_1142_)begin
        int_reg_array_16_19_imag <= _zz_1189_;
      end
      if(_zz_1143_)begin
        int_reg_array_16_20_imag <= _zz_1189_;
      end
      if(_zz_1144_)begin
        int_reg_array_16_21_imag <= _zz_1189_;
      end
      if(_zz_1145_)begin
        int_reg_array_16_22_imag <= _zz_1189_;
      end
      if(_zz_1146_)begin
        int_reg_array_16_23_imag <= _zz_1189_;
      end
      if(_zz_1147_)begin
        int_reg_array_16_24_imag <= _zz_1189_;
      end
      if(_zz_1148_)begin
        int_reg_array_16_25_imag <= _zz_1189_;
      end
      if(_zz_1149_)begin
        int_reg_array_16_26_imag <= _zz_1189_;
      end
      if(_zz_1150_)begin
        int_reg_array_16_27_imag <= _zz_1189_;
      end
      if(_zz_1151_)begin
        int_reg_array_16_28_imag <= _zz_1189_;
      end
      if(_zz_1152_)begin
        int_reg_array_16_29_imag <= _zz_1189_;
      end
      if(_zz_1153_)begin
        int_reg_array_16_30_imag <= _zz_1189_;
      end
      if(_zz_1154_)begin
        int_reg_array_16_31_imag <= _zz_1189_;
      end
      if(_zz_1155_)begin
        int_reg_array_16_32_imag <= _zz_1189_;
      end
      if(_zz_1156_)begin
        int_reg_array_16_33_imag <= _zz_1189_;
      end
      if(_zz_1157_)begin
        int_reg_array_16_34_imag <= _zz_1189_;
      end
      if(_zz_1158_)begin
        int_reg_array_16_35_imag <= _zz_1189_;
      end
      if(_zz_1159_)begin
        int_reg_array_16_36_imag <= _zz_1189_;
      end
      if(_zz_1160_)begin
        int_reg_array_16_37_imag <= _zz_1189_;
      end
      if(_zz_1161_)begin
        int_reg_array_16_38_imag <= _zz_1189_;
      end
      if(_zz_1162_)begin
        int_reg_array_16_39_imag <= _zz_1189_;
      end
      if(_zz_1163_)begin
        int_reg_array_16_40_imag <= _zz_1189_;
      end
      if(_zz_1164_)begin
        int_reg_array_16_41_imag <= _zz_1189_;
      end
      if(_zz_1165_)begin
        int_reg_array_16_42_imag <= _zz_1189_;
      end
      if(_zz_1166_)begin
        int_reg_array_16_43_imag <= _zz_1189_;
      end
      if(_zz_1167_)begin
        int_reg_array_16_44_imag <= _zz_1189_;
      end
      if(_zz_1168_)begin
        int_reg_array_16_45_imag <= _zz_1189_;
      end
      if(_zz_1169_)begin
        int_reg_array_16_46_imag <= _zz_1189_;
      end
      if(_zz_1170_)begin
        int_reg_array_16_47_imag <= _zz_1189_;
      end
      if(_zz_1171_)begin
        int_reg_array_16_48_imag <= _zz_1189_;
      end
      if(_zz_1172_)begin
        int_reg_array_16_49_imag <= _zz_1189_;
      end
      if(_zz_1173_)begin
        int_reg_array_16_50_imag <= _zz_1189_;
      end
      if(_zz_1174_)begin
        int_reg_array_16_51_imag <= _zz_1189_;
      end
      if(_zz_1175_)begin
        int_reg_array_16_52_imag <= _zz_1189_;
      end
      if(_zz_1176_)begin
        int_reg_array_16_53_imag <= _zz_1189_;
      end
      if(_zz_1177_)begin
        int_reg_array_16_54_imag <= _zz_1189_;
      end
      if(_zz_1178_)begin
        int_reg_array_16_55_imag <= _zz_1189_;
      end
      if(_zz_1179_)begin
        int_reg_array_16_56_imag <= _zz_1189_;
      end
      if(_zz_1180_)begin
        int_reg_array_16_57_imag <= _zz_1189_;
      end
      if(_zz_1181_)begin
        int_reg_array_16_58_imag <= _zz_1189_;
      end
      if(_zz_1182_)begin
        int_reg_array_16_59_imag <= _zz_1189_;
      end
      if(_zz_1183_)begin
        int_reg_array_16_60_imag <= _zz_1189_;
      end
      if(_zz_1184_)begin
        int_reg_array_16_61_imag <= _zz_1189_;
      end
      if(_zz_1185_)begin
        int_reg_array_16_62_imag <= _zz_1189_;
      end
      if(_zz_1186_)begin
        int_reg_array_16_63_imag <= _zz_1189_;
      end
      if(_zz_1192_)begin
        int_reg_array_17_0_real <= _zz_1257_;
      end
      if(_zz_1193_)begin
        int_reg_array_17_1_real <= _zz_1257_;
      end
      if(_zz_1194_)begin
        int_reg_array_17_2_real <= _zz_1257_;
      end
      if(_zz_1195_)begin
        int_reg_array_17_3_real <= _zz_1257_;
      end
      if(_zz_1196_)begin
        int_reg_array_17_4_real <= _zz_1257_;
      end
      if(_zz_1197_)begin
        int_reg_array_17_5_real <= _zz_1257_;
      end
      if(_zz_1198_)begin
        int_reg_array_17_6_real <= _zz_1257_;
      end
      if(_zz_1199_)begin
        int_reg_array_17_7_real <= _zz_1257_;
      end
      if(_zz_1200_)begin
        int_reg_array_17_8_real <= _zz_1257_;
      end
      if(_zz_1201_)begin
        int_reg_array_17_9_real <= _zz_1257_;
      end
      if(_zz_1202_)begin
        int_reg_array_17_10_real <= _zz_1257_;
      end
      if(_zz_1203_)begin
        int_reg_array_17_11_real <= _zz_1257_;
      end
      if(_zz_1204_)begin
        int_reg_array_17_12_real <= _zz_1257_;
      end
      if(_zz_1205_)begin
        int_reg_array_17_13_real <= _zz_1257_;
      end
      if(_zz_1206_)begin
        int_reg_array_17_14_real <= _zz_1257_;
      end
      if(_zz_1207_)begin
        int_reg_array_17_15_real <= _zz_1257_;
      end
      if(_zz_1208_)begin
        int_reg_array_17_16_real <= _zz_1257_;
      end
      if(_zz_1209_)begin
        int_reg_array_17_17_real <= _zz_1257_;
      end
      if(_zz_1210_)begin
        int_reg_array_17_18_real <= _zz_1257_;
      end
      if(_zz_1211_)begin
        int_reg_array_17_19_real <= _zz_1257_;
      end
      if(_zz_1212_)begin
        int_reg_array_17_20_real <= _zz_1257_;
      end
      if(_zz_1213_)begin
        int_reg_array_17_21_real <= _zz_1257_;
      end
      if(_zz_1214_)begin
        int_reg_array_17_22_real <= _zz_1257_;
      end
      if(_zz_1215_)begin
        int_reg_array_17_23_real <= _zz_1257_;
      end
      if(_zz_1216_)begin
        int_reg_array_17_24_real <= _zz_1257_;
      end
      if(_zz_1217_)begin
        int_reg_array_17_25_real <= _zz_1257_;
      end
      if(_zz_1218_)begin
        int_reg_array_17_26_real <= _zz_1257_;
      end
      if(_zz_1219_)begin
        int_reg_array_17_27_real <= _zz_1257_;
      end
      if(_zz_1220_)begin
        int_reg_array_17_28_real <= _zz_1257_;
      end
      if(_zz_1221_)begin
        int_reg_array_17_29_real <= _zz_1257_;
      end
      if(_zz_1222_)begin
        int_reg_array_17_30_real <= _zz_1257_;
      end
      if(_zz_1223_)begin
        int_reg_array_17_31_real <= _zz_1257_;
      end
      if(_zz_1224_)begin
        int_reg_array_17_32_real <= _zz_1257_;
      end
      if(_zz_1225_)begin
        int_reg_array_17_33_real <= _zz_1257_;
      end
      if(_zz_1226_)begin
        int_reg_array_17_34_real <= _zz_1257_;
      end
      if(_zz_1227_)begin
        int_reg_array_17_35_real <= _zz_1257_;
      end
      if(_zz_1228_)begin
        int_reg_array_17_36_real <= _zz_1257_;
      end
      if(_zz_1229_)begin
        int_reg_array_17_37_real <= _zz_1257_;
      end
      if(_zz_1230_)begin
        int_reg_array_17_38_real <= _zz_1257_;
      end
      if(_zz_1231_)begin
        int_reg_array_17_39_real <= _zz_1257_;
      end
      if(_zz_1232_)begin
        int_reg_array_17_40_real <= _zz_1257_;
      end
      if(_zz_1233_)begin
        int_reg_array_17_41_real <= _zz_1257_;
      end
      if(_zz_1234_)begin
        int_reg_array_17_42_real <= _zz_1257_;
      end
      if(_zz_1235_)begin
        int_reg_array_17_43_real <= _zz_1257_;
      end
      if(_zz_1236_)begin
        int_reg_array_17_44_real <= _zz_1257_;
      end
      if(_zz_1237_)begin
        int_reg_array_17_45_real <= _zz_1257_;
      end
      if(_zz_1238_)begin
        int_reg_array_17_46_real <= _zz_1257_;
      end
      if(_zz_1239_)begin
        int_reg_array_17_47_real <= _zz_1257_;
      end
      if(_zz_1240_)begin
        int_reg_array_17_48_real <= _zz_1257_;
      end
      if(_zz_1241_)begin
        int_reg_array_17_49_real <= _zz_1257_;
      end
      if(_zz_1242_)begin
        int_reg_array_17_50_real <= _zz_1257_;
      end
      if(_zz_1243_)begin
        int_reg_array_17_51_real <= _zz_1257_;
      end
      if(_zz_1244_)begin
        int_reg_array_17_52_real <= _zz_1257_;
      end
      if(_zz_1245_)begin
        int_reg_array_17_53_real <= _zz_1257_;
      end
      if(_zz_1246_)begin
        int_reg_array_17_54_real <= _zz_1257_;
      end
      if(_zz_1247_)begin
        int_reg_array_17_55_real <= _zz_1257_;
      end
      if(_zz_1248_)begin
        int_reg_array_17_56_real <= _zz_1257_;
      end
      if(_zz_1249_)begin
        int_reg_array_17_57_real <= _zz_1257_;
      end
      if(_zz_1250_)begin
        int_reg_array_17_58_real <= _zz_1257_;
      end
      if(_zz_1251_)begin
        int_reg_array_17_59_real <= _zz_1257_;
      end
      if(_zz_1252_)begin
        int_reg_array_17_60_real <= _zz_1257_;
      end
      if(_zz_1253_)begin
        int_reg_array_17_61_real <= _zz_1257_;
      end
      if(_zz_1254_)begin
        int_reg_array_17_62_real <= _zz_1257_;
      end
      if(_zz_1255_)begin
        int_reg_array_17_63_real <= _zz_1257_;
      end
      if(_zz_1192_)begin
        int_reg_array_17_0_imag <= _zz_1258_;
      end
      if(_zz_1193_)begin
        int_reg_array_17_1_imag <= _zz_1258_;
      end
      if(_zz_1194_)begin
        int_reg_array_17_2_imag <= _zz_1258_;
      end
      if(_zz_1195_)begin
        int_reg_array_17_3_imag <= _zz_1258_;
      end
      if(_zz_1196_)begin
        int_reg_array_17_4_imag <= _zz_1258_;
      end
      if(_zz_1197_)begin
        int_reg_array_17_5_imag <= _zz_1258_;
      end
      if(_zz_1198_)begin
        int_reg_array_17_6_imag <= _zz_1258_;
      end
      if(_zz_1199_)begin
        int_reg_array_17_7_imag <= _zz_1258_;
      end
      if(_zz_1200_)begin
        int_reg_array_17_8_imag <= _zz_1258_;
      end
      if(_zz_1201_)begin
        int_reg_array_17_9_imag <= _zz_1258_;
      end
      if(_zz_1202_)begin
        int_reg_array_17_10_imag <= _zz_1258_;
      end
      if(_zz_1203_)begin
        int_reg_array_17_11_imag <= _zz_1258_;
      end
      if(_zz_1204_)begin
        int_reg_array_17_12_imag <= _zz_1258_;
      end
      if(_zz_1205_)begin
        int_reg_array_17_13_imag <= _zz_1258_;
      end
      if(_zz_1206_)begin
        int_reg_array_17_14_imag <= _zz_1258_;
      end
      if(_zz_1207_)begin
        int_reg_array_17_15_imag <= _zz_1258_;
      end
      if(_zz_1208_)begin
        int_reg_array_17_16_imag <= _zz_1258_;
      end
      if(_zz_1209_)begin
        int_reg_array_17_17_imag <= _zz_1258_;
      end
      if(_zz_1210_)begin
        int_reg_array_17_18_imag <= _zz_1258_;
      end
      if(_zz_1211_)begin
        int_reg_array_17_19_imag <= _zz_1258_;
      end
      if(_zz_1212_)begin
        int_reg_array_17_20_imag <= _zz_1258_;
      end
      if(_zz_1213_)begin
        int_reg_array_17_21_imag <= _zz_1258_;
      end
      if(_zz_1214_)begin
        int_reg_array_17_22_imag <= _zz_1258_;
      end
      if(_zz_1215_)begin
        int_reg_array_17_23_imag <= _zz_1258_;
      end
      if(_zz_1216_)begin
        int_reg_array_17_24_imag <= _zz_1258_;
      end
      if(_zz_1217_)begin
        int_reg_array_17_25_imag <= _zz_1258_;
      end
      if(_zz_1218_)begin
        int_reg_array_17_26_imag <= _zz_1258_;
      end
      if(_zz_1219_)begin
        int_reg_array_17_27_imag <= _zz_1258_;
      end
      if(_zz_1220_)begin
        int_reg_array_17_28_imag <= _zz_1258_;
      end
      if(_zz_1221_)begin
        int_reg_array_17_29_imag <= _zz_1258_;
      end
      if(_zz_1222_)begin
        int_reg_array_17_30_imag <= _zz_1258_;
      end
      if(_zz_1223_)begin
        int_reg_array_17_31_imag <= _zz_1258_;
      end
      if(_zz_1224_)begin
        int_reg_array_17_32_imag <= _zz_1258_;
      end
      if(_zz_1225_)begin
        int_reg_array_17_33_imag <= _zz_1258_;
      end
      if(_zz_1226_)begin
        int_reg_array_17_34_imag <= _zz_1258_;
      end
      if(_zz_1227_)begin
        int_reg_array_17_35_imag <= _zz_1258_;
      end
      if(_zz_1228_)begin
        int_reg_array_17_36_imag <= _zz_1258_;
      end
      if(_zz_1229_)begin
        int_reg_array_17_37_imag <= _zz_1258_;
      end
      if(_zz_1230_)begin
        int_reg_array_17_38_imag <= _zz_1258_;
      end
      if(_zz_1231_)begin
        int_reg_array_17_39_imag <= _zz_1258_;
      end
      if(_zz_1232_)begin
        int_reg_array_17_40_imag <= _zz_1258_;
      end
      if(_zz_1233_)begin
        int_reg_array_17_41_imag <= _zz_1258_;
      end
      if(_zz_1234_)begin
        int_reg_array_17_42_imag <= _zz_1258_;
      end
      if(_zz_1235_)begin
        int_reg_array_17_43_imag <= _zz_1258_;
      end
      if(_zz_1236_)begin
        int_reg_array_17_44_imag <= _zz_1258_;
      end
      if(_zz_1237_)begin
        int_reg_array_17_45_imag <= _zz_1258_;
      end
      if(_zz_1238_)begin
        int_reg_array_17_46_imag <= _zz_1258_;
      end
      if(_zz_1239_)begin
        int_reg_array_17_47_imag <= _zz_1258_;
      end
      if(_zz_1240_)begin
        int_reg_array_17_48_imag <= _zz_1258_;
      end
      if(_zz_1241_)begin
        int_reg_array_17_49_imag <= _zz_1258_;
      end
      if(_zz_1242_)begin
        int_reg_array_17_50_imag <= _zz_1258_;
      end
      if(_zz_1243_)begin
        int_reg_array_17_51_imag <= _zz_1258_;
      end
      if(_zz_1244_)begin
        int_reg_array_17_52_imag <= _zz_1258_;
      end
      if(_zz_1245_)begin
        int_reg_array_17_53_imag <= _zz_1258_;
      end
      if(_zz_1246_)begin
        int_reg_array_17_54_imag <= _zz_1258_;
      end
      if(_zz_1247_)begin
        int_reg_array_17_55_imag <= _zz_1258_;
      end
      if(_zz_1248_)begin
        int_reg_array_17_56_imag <= _zz_1258_;
      end
      if(_zz_1249_)begin
        int_reg_array_17_57_imag <= _zz_1258_;
      end
      if(_zz_1250_)begin
        int_reg_array_17_58_imag <= _zz_1258_;
      end
      if(_zz_1251_)begin
        int_reg_array_17_59_imag <= _zz_1258_;
      end
      if(_zz_1252_)begin
        int_reg_array_17_60_imag <= _zz_1258_;
      end
      if(_zz_1253_)begin
        int_reg_array_17_61_imag <= _zz_1258_;
      end
      if(_zz_1254_)begin
        int_reg_array_17_62_imag <= _zz_1258_;
      end
      if(_zz_1255_)begin
        int_reg_array_17_63_imag <= _zz_1258_;
      end
      if(_zz_1261_)begin
        int_reg_array_18_0_real <= _zz_1326_;
      end
      if(_zz_1262_)begin
        int_reg_array_18_1_real <= _zz_1326_;
      end
      if(_zz_1263_)begin
        int_reg_array_18_2_real <= _zz_1326_;
      end
      if(_zz_1264_)begin
        int_reg_array_18_3_real <= _zz_1326_;
      end
      if(_zz_1265_)begin
        int_reg_array_18_4_real <= _zz_1326_;
      end
      if(_zz_1266_)begin
        int_reg_array_18_5_real <= _zz_1326_;
      end
      if(_zz_1267_)begin
        int_reg_array_18_6_real <= _zz_1326_;
      end
      if(_zz_1268_)begin
        int_reg_array_18_7_real <= _zz_1326_;
      end
      if(_zz_1269_)begin
        int_reg_array_18_8_real <= _zz_1326_;
      end
      if(_zz_1270_)begin
        int_reg_array_18_9_real <= _zz_1326_;
      end
      if(_zz_1271_)begin
        int_reg_array_18_10_real <= _zz_1326_;
      end
      if(_zz_1272_)begin
        int_reg_array_18_11_real <= _zz_1326_;
      end
      if(_zz_1273_)begin
        int_reg_array_18_12_real <= _zz_1326_;
      end
      if(_zz_1274_)begin
        int_reg_array_18_13_real <= _zz_1326_;
      end
      if(_zz_1275_)begin
        int_reg_array_18_14_real <= _zz_1326_;
      end
      if(_zz_1276_)begin
        int_reg_array_18_15_real <= _zz_1326_;
      end
      if(_zz_1277_)begin
        int_reg_array_18_16_real <= _zz_1326_;
      end
      if(_zz_1278_)begin
        int_reg_array_18_17_real <= _zz_1326_;
      end
      if(_zz_1279_)begin
        int_reg_array_18_18_real <= _zz_1326_;
      end
      if(_zz_1280_)begin
        int_reg_array_18_19_real <= _zz_1326_;
      end
      if(_zz_1281_)begin
        int_reg_array_18_20_real <= _zz_1326_;
      end
      if(_zz_1282_)begin
        int_reg_array_18_21_real <= _zz_1326_;
      end
      if(_zz_1283_)begin
        int_reg_array_18_22_real <= _zz_1326_;
      end
      if(_zz_1284_)begin
        int_reg_array_18_23_real <= _zz_1326_;
      end
      if(_zz_1285_)begin
        int_reg_array_18_24_real <= _zz_1326_;
      end
      if(_zz_1286_)begin
        int_reg_array_18_25_real <= _zz_1326_;
      end
      if(_zz_1287_)begin
        int_reg_array_18_26_real <= _zz_1326_;
      end
      if(_zz_1288_)begin
        int_reg_array_18_27_real <= _zz_1326_;
      end
      if(_zz_1289_)begin
        int_reg_array_18_28_real <= _zz_1326_;
      end
      if(_zz_1290_)begin
        int_reg_array_18_29_real <= _zz_1326_;
      end
      if(_zz_1291_)begin
        int_reg_array_18_30_real <= _zz_1326_;
      end
      if(_zz_1292_)begin
        int_reg_array_18_31_real <= _zz_1326_;
      end
      if(_zz_1293_)begin
        int_reg_array_18_32_real <= _zz_1326_;
      end
      if(_zz_1294_)begin
        int_reg_array_18_33_real <= _zz_1326_;
      end
      if(_zz_1295_)begin
        int_reg_array_18_34_real <= _zz_1326_;
      end
      if(_zz_1296_)begin
        int_reg_array_18_35_real <= _zz_1326_;
      end
      if(_zz_1297_)begin
        int_reg_array_18_36_real <= _zz_1326_;
      end
      if(_zz_1298_)begin
        int_reg_array_18_37_real <= _zz_1326_;
      end
      if(_zz_1299_)begin
        int_reg_array_18_38_real <= _zz_1326_;
      end
      if(_zz_1300_)begin
        int_reg_array_18_39_real <= _zz_1326_;
      end
      if(_zz_1301_)begin
        int_reg_array_18_40_real <= _zz_1326_;
      end
      if(_zz_1302_)begin
        int_reg_array_18_41_real <= _zz_1326_;
      end
      if(_zz_1303_)begin
        int_reg_array_18_42_real <= _zz_1326_;
      end
      if(_zz_1304_)begin
        int_reg_array_18_43_real <= _zz_1326_;
      end
      if(_zz_1305_)begin
        int_reg_array_18_44_real <= _zz_1326_;
      end
      if(_zz_1306_)begin
        int_reg_array_18_45_real <= _zz_1326_;
      end
      if(_zz_1307_)begin
        int_reg_array_18_46_real <= _zz_1326_;
      end
      if(_zz_1308_)begin
        int_reg_array_18_47_real <= _zz_1326_;
      end
      if(_zz_1309_)begin
        int_reg_array_18_48_real <= _zz_1326_;
      end
      if(_zz_1310_)begin
        int_reg_array_18_49_real <= _zz_1326_;
      end
      if(_zz_1311_)begin
        int_reg_array_18_50_real <= _zz_1326_;
      end
      if(_zz_1312_)begin
        int_reg_array_18_51_real <= _zz_1326_;
      end
      if(_zz_1313_)begin
        int_reg_array_18_52_real <= _zz_1326_;
      end
      if(_zz_1314_)begin
        int_reg_array_18_53_real <= _zz_1326_;
      end
      if(_zz_1315_)begin
        int_reg_array_18_54_real <= _zz_1326_;
      end
      if(_zz_1316_)begin
        int_reg_array_18_55_real <= _zz_1326_;
      end
      if(_zz_1317_)begin
        int_reg_array_18_56_real <= _zz_1326_;
      end
      if(_zz_1318_)begin
        int_reg_array_18_57_real <= _zz_1326_;
      end
      if(_zz_1319_)begin
        int_reg_array_18_58_real <= _zz_1326_;
      end
      if(_zz_1320_)begin
        int_reg_array_18_59_real <= _zz_1326_;
      end
      if(_zz_1321_)begin
        int_reg_array_18_60_real <= _zz_1326_;
      end
      if(_zz_1322_)begin
        int_reg_array_18_61_real <= _zz_1326_;
      end
      if(_zz_1323_)begin
        int_reg_array_18_62_real <= _zz_1326_;
      end
      if(_zz_1324_)begin
        int_reg_array_18_63_real <= _zz_1326_;
      end
      if(_zz_1261_)begin
        int_reg_array_18_0_imag <= _zz_1327_;
      end
      if(_zz_1262_)begin
        int_reg_array_18_1_imag <= _zz_1327_;
      end
      if(_zz_1263_)begin
        int_reg_array_18_2_imag <= _zz_1327_;
      end
      if(_zz_1264_)begin
        int_reg_array_18_3_imag <= _zz_1327_;
      end
      if(_zz_1265_)begin
        int_reg_array_18_4_imag <= _zz_1327_;
      end
      if(_zz_1266_)begin
        int_reg_array_18_5_imag <= _zz_1327_;
      end
      if(_zz_1267_)begin
        int_reg_array_18_6_imag <= _zz_1327_;
      end
      if(_zz_1268_)begin
        int_reg_array_18_7_imag <= _zz_1327_;
      end
      if(_zz_1269_)begin
        int_reg_array_18_8_imag <= _zz_1327_;
      end
      if(_zz_1270_)begin
        int_reg_array_18_9_imag <= _zz_1327_;
      end
      if(_zz_1271_)begin
        int_reg_array_18_10_imag <= _zz_1327_;
      end
      if(_zz_1272_)begin
        int_reg_array_18_11_imag <= _zz_1327_;
      end
      if(_zz_1273_)begin
        int_reg_array_18_12_imag <= _zz_1327_;
      end
      if(_zz_1274_)begin
        int_reg_array_18_13_imag <= _zz_1327_;
      end
      if(_zz_1275_)begin
        int_reg_array_18_14_imag <= _zz_1327_;
      end
      if(_zz_1276_)begin
        int_reg_array_18_15_imag <= _zz_1327_;
      end
      if(_zz_1277_)begin
        int_reg_array_18_16_imag <= _zz_1327_;
      end
      if(_zz_1278_)begin
        int_reg_array_18_17_imag <= _zz_1327_;
      end
      if(_zz_1279_)begin
        int_reg_array_18_18_imag <= _zz_1327_;
      end
      if(_zz_1280_)begin
        int_reg_array_18_19_imag <= _zz_1327_;
      end
      if(_zz_1281_)begin
        int_reg_array_18_20_imag <= _zz_1327_;
      end
      if(_zz_1282_)begin
        int_reg_array_18_21_imag <= _zz_1327_;
      end
      if(_zz_1283_)begin
        int_reg_array_18_22_imag <= _zz_1327_;
      end
      if(_zz_1284_)begin
        int_reg_array_18_23_imag <= _zz_1327_;
      end
      if(_zz_1285_)begin
        int_reg_array_18_24_imag <= _zz_1327_;
      end
      if(_zz_1286_)begin
        int_reg_array_18_25_imag <= _zz_1327_;
      end
      if(_zz_1287_)begin
        int_reg_array_18_26_imag <= _zz_1327_;
      end
      if(_zz_1288_)begin
        int_reg_array_18_27_imag <= _zz_1327_;
      end
      if(_zz_1289_)begin
        int_reg_array_18_28_imag <= _zz_1327_;
      end
      if(_zz_1290_)begin
        int_reg_array_18_29_imag <= _zz_1327_;
      end
      if(_zz_1291_)begin
        int_reg_array_18_30_imag <= _zz_1327_;
      end
      if(_zz_1292_)begin
        int_reg_array_18_31_imag <= _zz_1327_;
      end
      if(_zz_1293_)begin
        int_reg_array_18_32_imag <= _zz_1327_;
      end
      if(_zz_1294_)begin
        int_reg_array_18_33_imag <= _zz_1327_;
      end
      if(_zz_1295_)begin
        int_reg_array_18_34_imag <= _zz_1327_;
      end
      if(_zz_1296_)begin
        int_reg_array_18_35_imag <= _zz_1327_;
      end
      if(_zz_1297_)begin
        int_reg_array_18_36_imag <= _zz_1327_;
      end
      if(_zz_1298_)begin
        int_reg_array_18_37_imag <= _zz_1327_;
      end
      if(_zz_1299_)begin
        int_reg_array_18_38_imag <= _zz_1327_;
      end
      if(_zz_1300_)begin
        int_reg_array_18_39_imag <= _zz_1327_;
      end
      if(_zz_1301_)begin
        int_reg_array_18_40_imag <= _zz_1327_;
      end
      if(_zz_1302_)begin
        int_reg_array_18_41_imag <= _zz_1327_;
      end
      if(_zz_1303_)begin
        int_reg_array_18_42_imag <= _zz_1327_;
      end
      if(_zz_1304_)begin
        int_reg_array_18_43_imag <= _zz_1327_;
      end
      if(_zz_1305_)begin
        int_reg_array_18_44_imag <= _zz_1327_;
      end
      if(_zz_1306_)begin
        int_reg_array_18_45_imag <= _zz_1327_;
      end
      if(_zz_1307_)begin
        int_reg_array_18_46_imag <= _zz_1327_;
      end
      if(_zz_1308_)begin
        int_reg_array_18_47_imag <= _zz_1327_;
      end
      if(_zz_1309_)begin
        int_reg_array_18_48_imag <= _zz_1327_;
      end
      if(_zz_1310_)begin
        int_reg_array_18_49_imag <= _zz_1327_;
      end
      if(_zz_1311_)begin
        int_reg_array_18_50_imag <= _zz_1327_;
      end
      if(_zz_1312_)begin
        int_reg_array_18_51_imag <= _zz_1327_;
      end
      if(_zz_1313_)begin
        int_reg_array_18_52_imag <= _zz_1327_;
      end
      if(_zz_1314_)begin
        int_reg_array_18_53_imag <= _zz_1327_;
      end
      if(_zz_1315_)begin
        int_reg_array_18_54_imag <= _zz_1327_;
      end
      if(_zz_1316_)begin
        int_reg_array_18_55_imag <= _zz_1327_;
      end
      if(_zz_1317_)begin
        int_reg_array_18_56_imag <= _zz_1327_;
      end
      if(_zz_1318_)begin
        int_reg_array_18_57_imag <= _zz_1327_;
      end
      if(_zz_1319_)begin
        int_reg_array_18_58_imag <= _zz_1327_;
      end
      if(_zz_1320_)begin
        int_reg_array_18_59_imag <= _zz_1327_;
      end
      if(_zz_1321_)begin
        int_reg_array_18_60_imag <= _zz_1327_;
      end
      if(_zz_1322_)begin
        int_reg_array_18_61_imag <= _zz_1327_;
      end
      if(_zz_1323_)begin
        int_reg_array_18_62_imag <= _zz_1327_;
      end
      if(_zz_1324_)begin
        int_reg_array_18_63_imag <= _zz_1327_;
      end
      if(_zz_1330_)begin
        int_reg_array_19_0_real <= _zz_1395_;
      end
      if(_zz_1331_)begin
        int_reg_array_19_1_real <= _zz_1395_;
      end
      if(_zz_1332_)begin
        int_reg_array_19_2_real <= _zz_1395_;
      end
      if(_zz_1333_)begin
        int_reg_array_19_3_real <= _zz_1395_;
      end
      if(_zz_1334_)begin
        int_reg_array_19_4_real <= _zz_1395_;
      end
      if(_zz_1335_)begin
        int_reg_array_19_5_real <= _zz_1395_;
      end
      if(_zz_1336_)begin
        int_reg_array_19_6_real <= _zz_1395_;
      end
      if(_zz_1337_)begin
        int_reg_array_19_7_real <= _zz_1395_;
      end
      if(_zz_1338_)begin
        int_reg_array_19_8_real <= _zz_1395_;
      end
      if(_zz_1339_)begin
        int_reg_array_19_9_real <= _zz_1395_;
      end
      if(_zz_1340_)begin
        int_reg_array_19_10_real <= _zz_1395_;
      end
      if(_zz_1341_)begin
        int_reg_array_19_11_real <= _zz_1395_;
      end
      if(_zz_1342_)begin
        int_reg_array_19_12_real <= _zz_1395_;
      end
      if(_zz_1343_)begin
        int_reg_array_19_13_real <= _zz_1395_;
      end
      if(_zz_1344_)begin
        int_reg_array_19_14_real <= _zz_1395_;
      end
      if(_zz_1345_)begin
        int_reg_array_19_15_real <= _zz_1395_;
      end
      if(_zz_1346_)begin
        int_reg_array_19_16_real <= _zz_1395_;
      end
      if(_zz_1347_)begin
        int_reg_array_19_17_real <= _zz_1395_;
      end
      if(_zz_1348_)begin
        int_reg_array_19_18_real <= _zz_1395_;
      end
      if(_zz_1349_)begin
        int_reg_array_19_19_real <= _zz_1395_;
      end
      if(_zz_1350_)begin
        int_reg_array_19_20_real <= _zz_1395_;
      end
      if(_zz_1351_)begin
        int_reg_array_19_21_real <= _zz_1395_;
      end
      if(_zz_1352_)begin
        int_reg_array_19_22_real <= _zz_1395_;
      end
      if(_zz_1353_)begin
        int_reg_array_19_23_real <= _zz_1395_;
      end
      if(_zz_1354_)begin
        int_reg_array_19_24_real <= _zz_1395_;
      end
      if(_zz_1355_)begin
        int_reg_array_19_25_real <= _zz_1395_;
      end
      if(_zz_1356_)begin
        int_reg_array_19_26_real <= _zz_1395_;
      end
      if(_zz_1357_)begin
        int_reg_array_19_27_real <= _zz_1395_;
      end
      if(_zz_1358_)begin
        int_reg_array_19_28_real <= _zz_1395_;
      end
      if(_zz_1359_)begin
        int_reg_array_19_29_real <= _zz_1395_;
      end
      if(_zz_1360_)begin
        int_reg_array_19_30_real <= _zz_1395_;
      end
      if(_zz_1361_)begin
        int_reg_array_19_31_real <= _zz_1395_;
      end
      if(_zz_1362_)begin
        int_reg_array_19_32_real <= _zz_1395_;
      end
      if(_zz_1363_)begin
        int_reg_array_19_33_real <= _zz_1395_;
      end
      if(_zz_1364_)begin
        int_reg_array_19_34_real <= _zz_1395_;
      end
      if(_zz_1365_)begin
        int_reg_array_19_35_real <= _zz_1395_;
      end
      if(_zz_1366_)begin
        int_reg_array_19_36_real <= _zz_1395_;
      end
      if(_zz_1367_)begin
        int_reg_array_19_37_real <= _zz_1395_;
      end
      if(_zz_1368_)begin
        int_reg_array_19_38_real <= _zz_1395_;
      end
      if(_zz_1369_)begin
        int_reg_array_19_39_real <= _zz_1395_;
      end
      if(_zz_1370_)begin
        int_reg_array_19_40_real <= _zz_1395_;
      end
      if(_zz_1371_)begin
        int_reg_array_19_41_real <= _zz_1395_;
      end
      if(_zz_1372_)begin
        int_reg_array_19_42_real <= _zz_1395_;
      end
      if(_zz_1373_)begin
        int_reg_array_19_43_real <= _zz_1395_;
      end
      if(_zz_1374_)begin
        int_reg_array_19_44_real <= _zz_1395_;
      end
      if(_zz_1375_)begin
        int_reg_array_19_45_real <= _zz_1395_;
      end
      if(_zz_1376_)begin
        int_reg_array_19_46_real <= _zz_1395_;
      end
      if(_zz_1377_)begin
        int_reg_array_19_47_real <= _zz_1395_;
      end
      if(_zz_1378_)begin
        int_reg_array_19_48_real <= _zz_1395_;
      end
      if(_zz_1379_)begin
        int_reg_array_19_49_real <= _zz_1395_;
      end
      if(_zz_1380_)begin
        int_reg_array_19_50_real <= _zz_1395_;
      end
      if(_zz_1381_)begin
        int_reg_array_19_51_real <= _zz_1395_;
      end
      if(_zz_1382_)begin
        int_reg_array_19_52_real <= _zz_1395_;
      end
      if(_zz_1383_)begin
        int_reg_array_19_53_real <= _zz_1395_;
      end
      if(_zz_1384_)begin
        int_reg_array_19_54_real <= _zz_1395_;
      end
      if(_zz_1385_)begin
        int_reg_array_19_55_real <= _zz_1395_;
      end
      if(_zz_1386_)begin
        int_reg_array_19_56_real <= _zz_1395_;
      end
      if(_zz_1387_)begin
        int_reg_array_19_57_real <= _zz_1395_;
      end
      if(_zz_1388_)begin
        int_reg_array_19_58_real <= _zz_1395_;
      end
      if(_zz_1389_)begin
        int_reg_array_19_59_real <= _zz_1395_;
      end
      if(_zz_1390_)begin
        int_reg_array_19_60_real <= _zz_1395_;
      end
      if(_zz_1391_)begin
        int_reg_array_19_61_real <= _zz_1395_;
      end
      if(_zz_1392_)begin
        int_reg_array_19_62_real <= _zz_1395_;
      end
      if(_zz_1393_)begin
        int_reg_array_19_63_real <= _zz_1395_;
      end
      if(_zz_1330_)begin
        int_reg_array_19_0_imag <= _zz_1396_;
      end
      if(_zz_1331_)begin
        int_reg_array_19_1_imag <= _zz_1396_;
      end
      if(_zz_1332_)begin
        int_reg_array_19_2_imag <= _zz_1396_;
      end
      if(_zz_1333_)begin
        int_reg_array_19_3_imag <= _zz_1396_;
      end
      if(_zz_1334_)begin
        int_reg_array_19_4_imag <= _zz_1396_;
      end
      if(_zz_1335_)begin
        int_reg_array_19_5_imag <= _zz_1396_;
      end
      if(_zz_1336_)begin
        int_reg_array_19_6_imag <= _zz_1396_;
      end
      if(_zz_1337_)begin
        int_reg_array_19_7_imag <= _zz_1396_;
      end
      if(_zz_1338_)begin
        int_reg_array_19_8_imag <= _zz_1396_;
      end
      if(_zz_1339_)begin
        int_reg_array_19_9_imag <= _zz_1396_;
      end
      if(_zz_1340_)begin
        int_reg_array_19_10_imag <= _zz_1396_;
      end
      if(_zz_1341_)begin
        int_reg_array_19_11_imag <= _zz_1396_;
      end
      if(_zz_1342_)begin
        int_reg_array_19_12_imag <= _zz_1396_;
      end
      if(_zz_1343_)begin
        int_reg_array_19_13_imag <= _zz_1396_;
      end
      if(_zz_1344_)begin
        int_reg_array_19_14_imag <= _zz_1396_;
      end
      if(_zz_1345_)begin
        int_reg_array_19_15_imag <= _zz_1396_;
      end
      if(_zz_1346_)begin
        int_reg_array_19_16_imag <= _zz_1396_;
      end
      if(_zz_1347_)begin
        int_reg_array_19_17_imag <= _zz_1396_;
      end
      if(_zz_1348_)begin
        int_reg_array_19_18_imag <= _zz_1396_;
      end
      if(_zz_1349_)begin
        int_reg_array_19_19_imag <= _zz_1396_;
      end
      if(_zz_1350_)begin
        int_reg_array_19_20_imag <= _zz_1396_;
      end
      if(_zz_1351_)begin
        int_reg_array_19_21_imag <= _zz_1396_;
      end
      if(_zz_1352_)begin
        int_reg_array_19_22_imag <= _zz_1396_;
      end
      if(_zz_1353_)begin
        int_reg_array_19_23_imag <= _zz_1396_;
      end
      if(_zz_1354_)begin
        int_reg_array_19_24_imag <= _zz_1396_;
      end
      if(_zz_1355_)begin
        int_reg_array_19_25_imag <= _zz_1396_;
      end
      if(_zz_1356_)begin
        int_reg_array_19_26_imag <= _zz_1396_;
      end
      if(_zz_1357_)begin
        int_reg_array_19_27_imag <= _zz_1396_;
      end
      if(_zz_1358_)begin
        int_reg_array_19_28_imag <= _zz_1396_;
      end
      if(_zz_1359_)begin
        int_reg_array_19_29_imag <= _zz_1396_;
      end
      if(_zz_1360_)begin
        int_reg_array_19_30_imag <= _zz_1396_;
      end
      if(_zz_1361_)begin
        int_reg_array_19_31_imag <= _zz_1396_;
      end
      if(_zz_1362_)begin
        int_reg_array_19_32_imag <= _zz_1396_;
      end
      if(_zz_1363_)begin
        int_reg_array_19_33_imag <= _zz_1396_;
      end
      if(_zz_1364_)begin
        int_reg_array_19_34_imag <= _zz_1396_;
      end
      if(_zz_1365_)begin
        int_reg_array_19_35_imag <= _zz_1396_;
      end
      if(_zz_1366_)begin
        int_reg_array_19_36_imag <= _zz_1396_;
      end
      if(_zz_1367_)begin
        int_reg_array_19_37_imag <= _zz_1396_;
      end
      if(_zz_1368_)begin
        int_reg_array_19_38_imag <= _zz_1396_;
      end
      if(_zz_1369_)begin
        int_reg_array_19_39_imag <= _zz_1396_;
      end
      if(_zz_1370_)begin
        int_reg_array_19_40_imag <= _zz_1396_;
      end
      if(_zz_1371_)begin
        int_reg_array_19_41_imag <= _zz_1396_;
      end
      if(_zz_1372_)begin
        int_reg_array_19_42_imag <= _zz_1396_;
      end
      if(_zz_1373_)begin
        int_reg_array_19_43_imag <= _zz_1396_;
      end
      if(_zz_1374_)begin
        int_reg_array_19_44_imag <= _zz_1396_;
      end
      if(_zz_1375_)begin
        int_reg_array_19_45_imag <= _zz_1396_;
      end
      if(_zz_1376_)begin
        int_reg_array_19_46_imag <= _zz_1396_;
      end
      if(_zz_1377_)begin
        int_reg_array_19_47_imag <= _zz_1396_;
      end
      if(_zz_1378_)begin
        int_reg_array_19_48_imag <= _zz_1396_;
      end
      if(_zz_1379_)begin
        int_reg_array_19_49_imag <= _zz_1396_;
      end
      if(_zz_1380_)begin
        int_reg_array_19_50_imag <= _zz_1396_;
      end
      if(_zz_1381_)begin
        int_reg_array_19_51_imag <= _zz_1396_;
      end
      if(_zz_1382_)begin
        int_reg_array_19_52_imag <= _zz_1396_;
      end
      if(_zz_1383_)begin
        int_reg_array_19_53_imag <= _zz_1396_;
      end
      if(_zz_1384_)begin
        int_reg_array_19_54_imag <= _zz_1396_;
      end
      if(_zz_1385_)begin
        int_reg_array_19_55_imag <= _zz_1396_;
      end
      if(_zz_1386_)begin
        int_reg_array_19_56_imag <= _zz_1396_;
      end
      if(_zz_1387_)begin
        int_reg_array_19_57_imag <= _zz_1396_;
      end
      if(_zz_1388_)begin
        int_reg_array_19_58_imag <= _zz_1396_;
      end
      if(_zz_1389_)begin
        int_reg_array_19_59_imag <= _zz_1396_;
      end
      if(_zz_1390_)begin
        int_reg_array_19_60_imag <= _zz_1396_;
      end
      if(_zz_1391_)begin
        int_reg_array_19_61_imag <= _zz_1396_;
      end
      if(_zz_1392_)begin
        int_reg_array_19_62_imag <= _zz_1396_;
      end
      if(_zz_1393_)begin
        int_reg_array_19_63_imag <= _zz_1396_;
      end
      if(_zz_1399_)begin
        int_reg_array_20_0_real <= _zz_1464_;
      end
      if(_zz_1400_)begin
        int_reg_array_20_1_real <= _zz_1464_;
      end
      if(_zz_1401_)begin
        int_reg_array_20_2_real <= _zz_1464_;
      end
      if(_zz_1402_)begin
        int_reg_array_20_3_real <= _zz_1464_;
      end
      if(_zz_1403_)begin
        int_reg_array_20_4_real <= _zz_1464_;
      end
      if(_zz_1404_)begin
        int_reg_array_20_5_real <= _zz_1464_;
      end
      if(_zz_1405_)begin
        int_reg_array_20_6_real <= _zz_1464_;
      end
      if(_zz_1406_)begin
        int_reg_array_20_7_real <= _zz_1464_;
      end
      if(_zz_1407_)begin
        int_reg_array_20_8_real <= _zz_1464_;
      end
      if(_zz_1408_)begin
        int_reg_array_20_9_real <= _zz_1464_;
      end
      if(_zz_1409_)begin
        int_reg_array_20_10_real <= _zz_1464_;
      end
      if(_zz_1410_)begin
        int_reg_array_20_11_real <= _zz_1464_;
      end
      if(_zz_1411_)begin
        int_reg_array_20_12_real <= _zz_1464_;
      end
      if(_zz_1412_)begin
        int_reg_array_20_13_real <= _zz_1464_;
      end
      if(_zz_1413_)begin
        int_reg_array_20_14_real <= _zz_1464_;
      end
      if(_zz_1414_)begin
        int_reg_array_20_15_real <= _zz_1464_;
      end
      if(_zz_1415_)begin
        int_reg_array_20_16_real <= _zz_1464_;
      end
      if(_zz_1416_)begin
        int_reg_array_20_17_real <= _zz_1464_;
      end
      if(_zz_1417_)begin
        int_reg_array_20_18_real <= _zz_1464_;
      end
      if(_zz_1418_)begin
        int_reg_array_20_19_real <= _zz_1464_;
      end
      if(_zz_1419_)begin
        int_reg_array_20_20_real <= _zz_1464_;
      end
      if(_zz_1420_)begin
        int_reg_array_20_21_real <= _zz_1464_;
      end
      if(_zz_1421_)begin
        int_reg_array_20_22_real <= _zz_1464_;
      end
      if(_zz_1422_)begin
        int_reg_array_20_23_real <= _zz_1464_;
      end
      if(_zz_1423_)begin
        int_reg_array_20_24_real <= _zz_1464_;
      end
      if(_zz_1424_)begin
        int_reg_array_20_25_real <= _zz_1464_;
      end
      if(_zz_1425_)begin
        int_reg_array_20_26_real <= _zz_1464_;
      end
      if(_zz_1426_)begin
        int_reg_array_20_27_real <= _zz_1464_;
      end
      if(_zz_1427_)begin
        int_reg_array_20_28_real <= _zz_1464_;
      end
      if(_zz_1428_)begin
        int_reg_array_20_29_real <= _zz_1464_;
      end
      if(_zz_1429_)begin
        int_reg_array_20_30_real <= _zz_1464_;
      end
      if(_zz_1430_)begin
        int_reg_array_20_31_real <= _zz_1464_;
      end
      if(_zz_1431_)begin
        int_reg_array_20_32_real <= _zz_1464_;
      end
      if(_zz_1432_)begin
        int_reg_array_20_33_real <= _zz_1464_;
      end
      if(_zz_1433_)begin
        int_reg_array_20_34_real <= _zz_1464_;
      end
      if(_zz_1434_)begin
        int_reg_array_20_35_real <= _zz_1464_;
      end
      if(_zz_1435_)begin
        int_reg_array_20_36_real <= _zz_1464_;
      end
      if(_zz_1436_)begin
        int_reg_array_20_37_real <= _zz_1464_;
      end
      if(_zz_1437_)begin
        int_reg_array_20_38_real <= _zz_1464_;
      end
      if(_zz_1438_)begin
        int_reg_array_20_39_real <= _zz_1464_;
      end
      if(_zz_1439_)begin
        int_reg_array_20_40_real <= _zz_1464_;
      end
      if(_zz_1440_)begin
        int_reg_array_20_41_real <= _zz_1464_;
      end
      if(_zz_1441_)begin
        int_reg_array_20_42_real <= _zz_1464_;
      end
      if(_zz_1442_)begin
        int_reg_array_20_43_real <= _zz_1464_;
      end
      if(_zz_1443_)begin
        int_reg_array_20_44_real <= _zz_1464_;
      end
      if(_zz_1444_)begin
        int_reg_array_20_45_real <= _zz_1464_;
      end
      if(_zz_1445_)begin
        int_reg_array_20_46_real <= _zz_1464_;
      end
      if(_zz_1446_)begin
        int_reg_array_20_47_real <= _zz_1464_;
      end
      if(_zz_1447_)begin
        int_reg_array_20_48_real <= _zz_1464_;
      end
      if(_zz_1448_)begin
        int_reg_array_20_49_real <= _zz_1464_;
      end
      if(_zz_1449_)begin
        int_reg_array_20_50_real <= _zz_1464_;
      end
      if(_zz_1450_)begin
        int_reg_array_20_51_real <= _zz_1464_;
      end
      if(_zz_1451_)begin
        int_reg_array_20_52_real <= _zz_1464_;
      end
      if(_zz_1452_)begin
        int_reg_array_20_53_real <= _zz_1464_;
      end
      if(_zz_1453_)begin
        int_reg_array_20_54_real <= _zz_1464_;
      end
      if(_zz_1454_)begin
        int_reg_array_20_55_real <= _zz_1464_;
      end
      if(_zz_1455_)begin
        int_reg_array_20_56_real <= _zz_1464_;
      end
      if(_zz_1456_)begin
        int_reg_array_20_57_real <= _zz_1464_;
      end
      if(_zz_1457_)begin
        int_reg_array_20_58_real <= _zz_1464_;
      end
      if(_zz_1458_)begin
        int_reg_array_20_59_real <= _zz_1464_;
      end
      if(_zz_1459_)begin
        int_reg_array_20_60_real <= _zz_1464_;
      end
      if(_zz_1460_)begin
        int_reg_array_20_61_real <= _zz_1464_;
      end
      if(_zz_1461_)begin
        int_reg_array_20_62_real <= _zz_1464_;
      end
      if(_zz_1462_)begin
        int_reg_array_20_63_real <= _zz_1464_;
      end
      if(_zz_1399_)begin
        int_reg_array_20_0_imag <= _zz_1465_;
      end
      if(_zz_1400_)begin
        int_reg_array_20_1_imag <= _zz_1465_;
      end
      if(_zz_1401_)begin
        int_reg_array_20_2_imag <= _zz_1465_;
      end
      if(_zz_1402_)begin
        int_reg_array_20_3_imag <= _zz_1465_;
      end
      if(_zz_1403_)begin
        int_reg_array_20_4_imag <= _zz_1465_;
      end
      if(_zz_1404_)begin
        int_reg_array_20_5_imag <= _zz_1465_;
      end
      if(_zz_1405_)begin
        int_reg_array_20_6_imag <= _zz_1465_;
      end
      if(_zz_1406_)begin
        int_reg_array_20_7_imag <= _zz_1465_;
      end
      if(_zz_1407_)begin
        int_reg_array_20_8_imag <= _zz_1465_;
      end
      if(_zz_1408_)begin
        int_reg_array_20_9_imag <= _zz_1465_;
      end
      if(_zz_1409_)begin
        int_reg_array_20_10_imag <= _zz_1465_;
      end
      if(_zz_1410_)begin
        int_reg_array_20_11_imag <= _zz_1465_;
      end
      if(_zz_1411_)begin
        int_reg_array_20_12_imag <= _zz_1465_;
      end
      if(_zz_1412_)begin
        int_reg_array_20_13_imag <= _zz_1465_;
      end
      if(_zz_1413_)begin
        int_reg_array_20_14_imag <= _zz_1465_;
      end
      if(_zz_1414_)begin
        int_reg_array_20_15_imag <= _zz_1465_;
      end
      if(_zz_1415_)begin
        int_reg_array_20_16_imag <= _zz_1465_;
      end
      if(_zz_1416_)begin
        int_reg_array_20_17_imag <= _zz_1465_;
      end
      if(_zz_1417_)begin
        int_reg_array_20_18_imag <= _zz_1465_;
      end
      if(_zz_1418_)begin
        int_reg_array_20_19_imag <= _zz_1465_;
      end
      if(_zz_1419_)begin
        int_reg_array_20_20_imag <= _zz_1465_;
      end
      if(_zz_1420_)begin
        int_reg_array_20_21_imag <= _zz_1465_;
      end
      if(_zz_1421_)begin
        int_reg_array_20_22_imag <= _zz_1465_;
      end
      if(_zz_1422_)begin
        int_reg_array_20_23_imag <= _zz_1465_;
      end
      if(_zz_1423_)begin
        int_reg_array_20_24_imag <= _zz_1465_;
      end
      if(_zz_1424_)begin
        int_reg_array_20_25_imag <= _zz_1465_;
      end
      if(_zz_1425_)begin
        int_reg_array_20_26_imag <= _zz_1465_;
      end
      if(_zz_1426_)begin
        int_reg_array_20_27_imag <= _zz_1465_;
      end
      if(_zz_1427_)begin
        int_reg_array_20_28_imag <= _zz_1465_;
      end
      if(_zz_1428_)begin
        int_reg_array_20_29_imag <= _zz_1465_;
      end
      if(_zz_1429_)begin
        int_reg_array_20_30_imag <= _zz_1465_;
      end
      if(_zz_1430_)begin
        int_reg_array_20_31_imag <= _zz_1465_;
      end
      if(_zz_1431_)begin
        int_reg_array_20_32_imag <= _zz_1465_;
      end
      if(_zz_1432_)begin
        int_reg_array_20_33_imag <= _zz_1465_;
      end
      if(_zz_1433_)begin
        int_reg_array_20_34_imag <= _zz_1465_;
      end
      if(_zz_1434_)begin
        int_reg_array_20_35_imag <= _zz_1465_;
      end
      if(_zz_1435_)begin
        int_reg_array_20_36_imag <= _zz_1465_;
      end
      if(_zz_1436_)begin
        int_reg_array_20_37_imag <= _zz_1465_;
      end
      if(_zz_1437_)begin
        int_reg_array_20_38_imag <= _zz_1465_;
      end
      if(_zz_1438_)begin
        int_reg_array_20_39_imag <= _zz_1465_;
      end
      if(_zz_1439_)begin
        int_reg_array_20_40_imag <= _zz_1465_;
      end
      if(_zz_1440_)begin
        int_reg_array_20_41_imag <= _zz_1465_;
      end
      if(_zz_1441_)begin
        int_reg_array_20_42_imag <= _zz_1465_;
      end
      if(_zz_1442_)begin
        int_reg_array_20_43_imag <= _zz_1465_;
      end
      if(_zz_1443_)begin
        int_reg_array_20_44_imag <= _zz_1465_;
      end
      if(_zz_1444_)begin
        int_reg_array_20_45_imag <= _zz_1465_;
      end
      if(_zz_1445_)begin
        int_reg_array_20_46_imag <= _zz_1465_;
      end
      if(_zz_1446_)begin
        int_reg_array_20_47_imag <= _zz_1465_;
      end
      if(_zz_1447_)begin
        int_reg_array_20_48_imag <= _zz_1465_;
      end
      if(_zz_1448_)begin
        int_reg_array_20_49_imag <= _zz_1465_;
      end
      if(_zz_1449_)begin
        int_reg_array_20_50_imag <= _zz_1465_;
      end
      if(_zz_1450_)begin
        int_reg_array_20_51_imag <= _zz_1465_;
      end
      if(_zz_1451_)begin
        int_reg_array_20_52_imag <= _zz_1465_;
      end
      if(_zz_1452_)begin
        int_reg_array_20_53_imag <= _zz_1465_;
      end
      if(_zz_1453_)begin
        int_reg_array_20_54_imag <= _zz_1465_;
      end
      if(_zz_1454_)begin
        int_reg_array_20_55_imag <= _zz_1465_;
      end
      if(_zz_1455_)begin
        int_reg_array_20_56_imag <= _zz_1465_;
      end
      if(_zz_1456_)begin
        int_reg_array_20_57_imag <= _zz_1465_;
      end
      if(_zz_1457_)begin
        int_reg_array_20_58_imag <= _zz_1465_;
      end
      if(_zz_1458_)begin
        int_reg_array_20_59_imag <= _zz_1465_;
      end
      if(_zz_1459_)begin
        int_reg_array_20_60_imag <= _zz_1465_;
      end
      if(_zz_1460_)begin
        int_reg_array_20_61_imag <= _zz_1465_;
      end
      if(_zz_1461_)begin
        int_reg_array_20_62_imag <= _zz_1465_;
      end
      if(_zz_1462_)begin
        int_reg_array_20_63_imag <= _zz_1465_;
      end
      if(_zz_1468_)begin
        int_reg_array_21_0_real <= _zz_1533_;
      end
      if(_zz_1469_)begin
        int_reg_array_21_1_real <= _zz_1533_;
      end
      if(_zz_1470_)begin
        int_reg_array_21_2_real <= _zz_1533_;
      end
      if(_zz_1471_)begin
        int_reg_array_21_3_real <= _zz_1533_;
      end
      if(_zz_1472_)begin
        int_reg_array_21_4_real <= _zz_1533_;
      end
      if(_zz_1473_)begin
        int_reg_array_21_5_real <= _zz_1533_;
      end
      if(_zz_1474_)begin
        int_reg_array_21_6_real <= _zz_1533_;
      end
      if(_zz_1475_)begin
        int_reg_array_21_7_real <= _zz_1533_;
      end
      if(_zz_1476_)begin
        int_reg_array_21_8_real <= _zz_1533_;
      end
      if(_zz_1477_)begin
        int_reg_array_21_9_real <= _zz_1533_;
      end
      if(_zz_1478_)begin
        int_reg_array_21_10_real <= _zz_1533_;
      end
      if(_zz_1479_)begin
        int_reg_array_21_11_real <= _zz_1533_;
      end
      if(_zz_1480_)begin
        int_reg_array_21_12_real <= _zz_1533_;
      end
      if(_zz_1481_)begin
        int_reg_array_21_13_real <= _zz_1533_;
      end
      if(_zz_1482_)begin
        int_reg_array_21_14_real <= _zz_1533_;
      end
      if(_zz_1483_)begin
        int_reg_array_21_15_real <= _zz_1533_;
      end
      if(_zz_1484_)begin
        int_reg_array_21_16_real <= _zz_1533_;
      end
      if(_zz_1485_)begin
        int_reg_array_21_17_real <= _zz_1533_;
      end
      if(_zz_1486_)begin
        int_reg_array_21_18_real <= _zz_1533_;
      end
      if(_zz_1487_)begin
        int_reg_array_21_19_real <= _zz_1533_;
      end
      if(_zz_1488_)begin
        int_reg_array_21_20_real <= _zz_1533_;
      end
      if(_zz_1489_)begin
        int_reg_array_21_21_real <= _zz_1533_;
      end
      if(_zz_1490_)begin
        int_reg_array_21_22_real <= _zz_1533_;
      end
      if(_zz_1491_)begin
        int_reg_array_21_23_real <= _zz_1533_;
      end
      if(_zz_1492_)begin
        int_reg_array_21_24_real <= _zz_1533_;
      end
      if(_zz_1493_)begin
        int_reg_array_21_25_real <= _zz_1533_;
      end
      if(_zz_1494_)begin
        int_reg_array_21_26_real <= _zz_1533_;
      end
      if(_zz_1495_)begin
        int_reg_array_21_27_real <= _zz_1533_;
      end
      if(_zz_1496_)begin
        int_reg_array_21_28_real <= _zz_1533_;
      end
      if(_zz_1497_)begin
        int_reg_array_21_29_real <= _zz_1533_;
      end
      if(_zz_1498_)begin
        int_reg_array_21_30_real <= _zz_1533_;
      end
      if(_zz_1499_)begin
        int_reg_array_21_31_real <= _zz_1533_;
      end
      if(_zz_1500_)begin
        int_reg_array_21_32_real <= _zz_1533_;
      end
      if(_zz_1501_)begin
        int_reg_array_21_33_real <= _zz_1533_;
      end
      if(_zz_1502_)begin
        int_reg_array_21_34_real <= _zz_1533_;
      end
      if(_zz_1503_)begin
        int_reg_array_21_35_real <= _zz_1533_;
      end
      if(_zz_1504_)begin
        int_reg_array_21_36_real <= _zz_1533_;
      end
      if(_zz_1505_)begin
        int_reg_array_21_37_real <= _zz_1533_;
      end
      if(_zz_1506_)begin
        int_reg_array_21_38_real <= _zz_1533_;
      end
      if(_zz_1507_)begin
        int_reg_array_21_39_real <= _zz_1533_;
      end
      if(_zz_1508_)begin
        int_reg_array_21_40_real <= _zz_1533_;
      end
      if(_zz_1509_)begin
        int_reg_array_21_41_real <= _zz_1533_;
      end
      if(_zz_1510_)begin
        int_reg_array_21_42_real <= _zz_1533_;
      end
      if(_zz_1511_)begin
        int_reg_array_21_43_real <= _zz_1533_;
      end
      if(_zz_1512_)begin
        int_reg_array_21_44_real <= _zz_1533_;
      end
      if(_zz_1513_)begin
        int_reg_array_21_45_real <= _zz_1533_;
      end
      if(_zz_1514_)begin
        int_reg_array_21_46_real <= _zz_1533_;
      end
      if(_zz_1515_)begin
        int_reg_array_21_47_real <= _zz_1533_;
      end
      if(_zz_1516_)begin
        int_reg_array_21_48_real <= _zz_1533_;
      end
      if(_zz_1517_)begin
        int_reg_array_21_49_real <= _zz_1533_;
      end
      if(_zz_1518_)begin
        int_reg_array_21_50_real <= _zz_1533_;
      end
      if(_zz_1519_)begin
        int_reg_array_21_51_real <= _zz_1533_;
      end
      if(_zz_1520_)begin
        int_reg_array_21_52_real <= _zz_1533_;
      end
      if(_zz_1521_)begin
        int_reg_array_21_53_real <= _zz_1533_;
      end
      if(_zz_1522_)begin
        int_reg_array_21_54_real <= _zz_1533_;
      end
      if(_zz_1523_)begin
        int_reg_array_21_55_real <= _zz_1533_;
      end
      if(_zz_1524_)begin
        int_reg_array_21_56_real <= _zz_1533_;
      end
      if(_zz_1525_)begin
        int_reg_array_21_57_real <= _zz_1533_;
      end
      if(_zz_1526_)begin
        int_reg_array_21_58_real <= _zz_1533_;
      end
      if(_zz_1527_)begin
        int_reg_array_21_59_real <= _zz_1533_;
      end
      if(_zz_1528_)begin
        int_reg_array_21_60_real <= _zz_1533_;
      end
      if(_zz_1529_)begin
        int_reg_array_21_61_real <= _zz_1533_;
      end
      if(_zz_1530_)begin
        int_reg_array_21_62_real <= _zz_1533_;
      end
      if(_zz_1531_)begin
        int_reg_array_21_63_real <= _zz_1533_;
      end
      if(_zz_1468_)begin
        int_reg_array_21_0_imag <= _zz_1534_;
      end
      if(_zz_1469_)begin
        int_reg_array_21_1_imag <= _zz_1534_;
      end
      if(_zz_1470_)begin
        int_reg_array_21_2_imag <= _zz_1534_;
      end
      if(_zz_1471_)begin
        int_reg_array_21_3_imag <= _zz_1534_;
      end
      if(_zz_1472_)begin
        int_reg_array_21_4_imag <= _zz_1534_;
      end
      if(_zz_1473_)begin
        int_reg_array_21_5_imag <= _zz_1534_;
      end
      if(_zz_1474_)begin
        int_reg_array_21_6_imag <= _zz_1534_;
      end
      if(_zz_1475_)begin
        int_reg_array_21_7_imag <= _zz_1534_;
      end
      if(_zz_1476_)begin
        int_reg_array_21_8_imag <= _zz_1534_;
      end
      if(_zz_1477_)begin
        int_reg_array_21_9_imag <= _zz_1534_;
      end
      if(_zz_1478_)begin
        int_reg_array_21_10_imag <= _zz_1534_;
      end
      if(_zz_1479_)begin
        int_reg_array_21_11_imag <= _zz_1534_;
      end
      if(_zz_1480_)begin
        int_reg_array_21_12_imag <= _zz_1534_;
      end
      if(_zz_1481_)begin
        int_reg_array_21_13_imag <= _zz_1534_;
      end
      if(_zz_1482_)begin
        int_reg_array_21_14_imag <= _zz_1534_;
      end
      if(_zz_1483_)begin
        int_reg_array_21_15_imag <= _zz_1534_;
      end
      if(_zz_1484_)begin
        int_reg_array_21_16_imag <= _zz_1534_;
      end
      if(_zz_1485_)begin
        int_reg_array_21_17_imag <= _zz_1534_;
      end
      if(_zz_1486_)begin
        int_reg_array_21_18_imag <= _zz_1534_;
      end
      if(_zz_1487_)begin
        int_reg_array_21_19_imag <= _zz_1534_;
      end
      if(_zz_1488_)begin
        int_reg_array_21_20_imag <= _zz_1534_;
      end
      if(_zz_1489_)begin
        int_reg_array_21_21_imag <= _zz_1534_;
      end
      if(_zz_1490_)begin
        int_reg_array_21_22_imag <= _zz_1534_;
      end
      if(_zz_1491_)begin
        int_reg_array_21_23_imag <= _zz_1534_;
      end
      if(_zz_1492_)begin
        int_reg_array_21_24_imag <= _zz_1534_;
      end
      if(_zz_1493_)begin
        int_reg_array_21_25_imag <= _zz_1534_;
      end
      if(_zz_1494_)begin
        int_reg_array_21_26_imag <= _zz_1534_;
      end
      if(_zz_1495_)begin
        int_reg_array_21_27_imag <= _zz_1534_;
      end
      if(_zz_1496_)begin
        int_reg_array_21_28_imag <= _zz_1534_;
      end
      if(_zz_1497_)begin
        int_reg_array_21_29_imag <= _zz_1534_;
      end
      if(_zz_1498_)begin
        int_reg_array_21_30_imag <= _zz_1534_;
      end
      if(_zz_1499_)begin
        int_reg_array_21_31_imag <= _zz_1534_;
      end
      if(_zz_1500_)begin
        int_reg_array_21_32_imag <= _zz_1534_;
      end
      if(_zz_1501_)begin
        int_reg_array_21_33_imag <= _zz_1534_;
      end
      if(_zz_1502_)begin
        int_reg_array_21_34_imag <= _zz_1534_;
      end
      if(_zz_1503_)begin
        int_reg_array_21_35_imag <= _zz_1534_;
      end
      if(_zz_1504_)begin
        int_reg_array_21_36_imag <= _zz_1534_;
      end
      if(_zz_1505_)begin
        int_reg_array_21_37_imag <= _zz_1534_;
      end
      if(_zz_1506_)begin
        int_reg_array_21_38_imag <= _zz_1534_;
      end
      if(_zz_1507_)begin
        int_reg_array_21_39_imag <= _zz_1534_;
      end
      if(_zz_1508_)begin
        int_reg_array_21_40_imag <= _zz_1534_;
      end
      if(_zz_1509_)begin
        int_reg_array_21_41_imag <= _zz_1534_;
      end
      if(_zz_1510_)begin
        int_reg_array_21_42_imag <= _zz_1534_;
      end
      if(_zz_1511_)begin
        int_reg_array_21_43_imag <= _zz_1534_;
      end
      if(_zz_1512_)begin
        int_reg_array_21_44_imag <= _zz_1534_;
      end
      if(_zz_1513_)begin
        int_reg_array_21_45_imag <= _zz_1534_;
      end
      if(_zz_1514_)begin
        int_reg_array_21_46_imag <= _zz_1534_;
      end
      if(_zz_1515_)begin
        int_reg_array_21_47_imag <= _zz_1534_;
      end
      if(_zz_1516_)begin
        int_reg_array_21_48_imag <= _zz_1534_;
      end
      if(_zz_1517_)begin
        int_reg_array_21_49_imag <= _zz_1534_;
      end
      if(_zz_1518_)begin
        int_reg_array_21_50_imag <= _zz_1534_;
      end
      if(_zz_1519_)begin
        int_reg_array_21_51_imag <= _zz_1534_;
      end
      if(_zz_1520_)begin
        int_reg_array_21_52_imag <= _zz_1534_;
      end
      if(_zz_1521_)begin
        int_reg_array_21_53_imag <= _zz_1534_;
      end
      if(_zz_1522_)begin
        int_reg_array_21_54_imag <= _zz_1534_;
      end
      if(_zz_1523_)begin
        int_reg_array_21_55_imag <= _zz_1534_;
      end
      if(_zz_1524_)begin
        int_reg_array_21_56_imag <= _zz_1534_;
      end
      if(_zz_1525_)begin
        int_reg_array_21_57_imag <= _zz_1534_;
      end
      if(_zz_1526_)begin
        int_reg_array_21_58_imag <= _zz_1534_;
      end
      if(_zz_1527_)begin
        int_reg_array_21_59_imag <= _zz_1534_;
      end
      if(_zz_1528_)begin
        int_reg_array_21_60_imag <= _zz_1534_;
      end
      if(_zz_1529_)begin
        int_reg_array_21_61_imag <= _zz_1534_;
      end
      if(_zz_1530_)begin
        int_reg_array_21_62_imag <= _zz_1534_;
      end
      if(_zz_1531_)begin
        int_reg_array_21_63_imag <= _zz_1534_;
      end
      if(_zz_1537_)begin
        int_reg_array_22_0_real <= _zz_1602_;
      end
      if(_zz_1538_)begin
        int_reg_array_22_1_real <= _zz_1602_;
      end
      if(_zz_1539_)begin
        int_reg_array_22_2_real <= _zz_1602_;
      end
      if(_zz_1540_)begin
        int_reg_array_22_3_real <= _zz_1602_;
      end
      if(_zz_1541_)begin
        int_reg_array_22_4_real <= _zz_1602_;
      end
      if(_zz_1542_)begin
        int_reg_array_22_5_real <= _zz_1602_;
      end
      if(_zz_1543_)begin
        int_reg_array_22_6_real <= _zz_1602_;
      end
      if(_zz_1544_)begin
        int_reg_array_22_7_real <= _zz_1602_;
      end
      if(_zz_1545_)begin
        int_reg_array_22_8_real <= _zz_1602_;
      end
      if(_zz_1546_)begin
        int_reg_array_22_9_real <= _zz_1602_;
      end
      if(_zz_1547_)begin
        int_reg_array_22_10_real <= _zz_1602_;
      end
      if(_zz_1548_)begin
        int_reg_array_22_11_real <= _zz_1602_;
      end
      if(_zz_1549_)begin
        int_reg_array_22_12_real <= _zz_1602_;
      end
      if(_zz_1550_)begin
        int_reg_array_22_13_real <= _zz_1602_;
      end
      if(_zz_1551_)begin
        int_reg_array_22_14_real <= _zz_1602_;
      end
      if(_zz_1552_)begin
        int_reg_array_22_15_real <= _zz_1602_;
      end
      if(_zz_1553_)begin
        int_reg_array_22_16_real <= _zz_1602_;
      end
      if(_zz_1554_)begin
        int_reg_array_22_17_real <= _zz_1602_;
      end
      if(_zz_1555_)begin
        int_reg_array_22_18_real <= _zz_1602_;
      end
      if(_zz_1556_)begin
        int_reg_array_22_19_real <= _zz_1602_;
      end
      if(_zz_1557_)begin
        int_reg_array_22_20_real <= _zz_1602_;
      end
      if(_zz_1558_)begin
        int_reg_array_22_21_real <= _zz_1602_;
      end
      if(_zz_1559_)begin
        int_reg_array_22_22_real <= _zz_1602_;
      end
      if(_zz_1560_)begin
        int_reg_array_22_23_real <= _zz_1602_;
      end
      if(_zz_1561_)begin
        int_reg_array_22_24_real <= _zz_1602_;
      end
      if(_zz_1562_)begin
        int_reg_array_22_25_real <= _zz_1602_;
      end
      if(_zz_1563_)begin
        int_reg_array_22_26_real <= _zz_1602_;
      end
      if(_zz_1564_)begin
        int_reg_array_22_27_real <= _zz_1602_;
      end
      if(_zz_1565_)begin
        int_reg_array_22_28_real <= _zz_1602_;
      end
      if(_zz_1566_)begin
        int_reg_array_22_29_real <= _zz_1602_;
      end
      if(_zz_1567_)begin
        int_reg_array_22_30_real <= _zz_1602_;
      end
      if(_zz_1568_)begin
        int_reg_array_22_31_real <= _zz_1602_;
      end
      if(_zz_1569_)begin
        int_reg_array_22_32_real <= _zz_1602_;
      end
      if(_zz_1570_)begin
        int_reg_array_22_33_real <= _zz_1602_;
      end
      if(_zz_1571_)begin
        int_reg_array_22_34_real <= _zz_1602_;
      end
      if(_zz_1572_)begin
        int_reg_array_22_35_real <= _zz_1602_;
      end
      if(_zz_1573_)begin
        int_reg_array_22_36_real <= _zz_1602_;
      end
      if(_zz_1574_)begin
        int_reg_array_22_37_real <= _zz_1602_;
      end
      if(_zz_1575_)begin
        int_reg_array_22_38_real <= _zz_1602_;
      end
      if(_zz_1576_)begin
        int_reg_array_22_39_real <= _zz_1602_;
      end
      if(_zz_1577_)begin
        int_reg_array_22_40_real <= _zz_1602_;
      end
      if(_zz_1578_)begin
        int_reg_array_22_41_real <= _zz_1602_;
      end
      if(_zz_1579_)begin
        int_reg_array_22_42_real <= _zz_1602_;
      end
      if(_zz_1580_)begin
        int_reg_array_22_43_real <= _zz_1602_;
      end
      if(_zz_1581_)begin
        int_reg_array_22_44_real <= _zz_1602_;
      end
      if(_zz_1582_)begin
        int_reg_array_22_45_real <= _zz_1602_;
      end
      if(_zz_1583_)begin
        int_reg_array_22_46_real <= _zz_1602_;
      end
      if(_zz_1584_)begin
        int_reg_array_22_47_real <= _zz_1602_;
      end
      if(_zz_1585_)begin
        int_reg_array_22_48_real <= _zz_1602_;
      end
      if(_zz_1586_)begin
        int_reg_array_22_49_real <= _zz_1602_;
      end
      if(_zz_1587_)begin
        int_reg_array_22_50_real <= _zz_1602_;
      end
      if(_zz_1588_)begin
        int_reg_array_22_51_real <= _zz_1602_;
      end
      if(_zz_1589_)begin
        int_reg_array_22_52_real <= _zz_1602_;
      end
      if(_zz_1590_)begin
        int_reg_array_22_53_real <= _zz_1602_;
      end
      if(_zz_1591_)begin
        int_reg_array_22_54_real <= _zz_1602_;
      end
      if(_zz_1592_)begin
        int_reg_array_22_55_real <= _zz_1602_;
      end
      if(_zz_1593_)begin
        int_reg_array_22_56_real <= _zz_1602_;
      end
      if(_zz_1594_)begin
        int_reg_array_22_57_real <= _zz_1602_;
      end
      if(_zz_1595_)begin
        int_reg_array_22_58_real <= _zz_1602_;
      end
      if(_zz_1596_)begin
        int_reg_array_22_59_real <= _zz_1602_;
      end
      if(_zz_1597_)begin
        int_reg_array_22_60_real <= _zz_1602_;
      end
      if(_zz_1598_)begin
        int_reg_array_22_61_real <= _zz_1602_;
      end
      if(_zz_1599_)begin
        int_reg_array_22_62_real <= _zz_1602_;
      end
      if(_zz_1600_)begin
        int_reg_array_22_63_real <= _zz_1602_;
      end
      if(_zz_1537_)begin
        int_reg_array_22_0_imag <= _zz_1603_;
      end
      if(_zz_1538_)begin
        int_reg_array_22_1_imag <= _zz_1603_;
      end
      if(_zz_1539_)begin
        int_reg_array_22_2_imag <= _zz_1603_;
      end
      if(_zz_1540_)begin
        int_reg_array_22_3_imag <= _zz_1603_;
      end
      if(_zz_1541_)begin
        int_reg_array_22_4_imag <= _zz_1603_;
      end
      if(_zz_1542_)begin
        int_reg_array_22_5_imag <= _zz_1603_;
      end
      if(_zz_1543_)begin
        int_reg_array_22_6_imag <= _zz_1603_;
      end
      if(_zz_1544_)begin
        int_reg_array_22_7_imag <= _zz_1603_;
      end
      if(_zz_1545_)begin
        int_reg_array_22_8_imag <= _zz_1603_;
      end
      if(_zz_1546_)begin
        int_reg_array_22_9_imag <= _zz_1603_;
      end
      if(_zz_1547_)begin
        int_reg_array_22_10_imag <= _zz_1603_;
      end
      if(_zz_1548_)begin
        int_reg_array_22_11_imag <= _zz_1603_;
      end
      if(_zz_1549_)begin
        int_reg_array_22_12_imag <= _zz_1603_;
      end
      if(_zz_1550_)begin
        int_reg_array_22_13_imag <= _zz_1603_;
      end
      if(_zz_1551_)begin
        int_reg_array_22_14_imag <= _zz_1603_;
      end
      if(_zz_1552_)begin
        int_reg_array_22_15_imag <= _zz_1603_;
      end
      if(_zz_1553_)begin
        int_reg_array_22_16_imag <= _zz_1603_;
      end
      if(_zz_1554_)begin
        int_reg_array_22_17_imag <= _zz_1603_;
      end
      if(_zz_1555_)begin
        int_reg_array_22_18_imag <= _zz_1603_;
      end
      if(_zz_1556_)begin
        int_reg_array_22_19_imag <= _zz_1603_;
      end
      if(_zz_1557_)begin
        int_reg_array_22_20_imag <= _zz_1603_;
      end
      if(_zz_1558_)begin
        int_reg_array_22_21_imag <= _zz_1603_;
      end
      if(_zz_1559_)begin
        int_reg_array_22_22_imag <= _zz_1603_;
      end
      if(_zz_1560_)begin
        int_reg_array_22_23_imag <= _zz_1603_;
      end
      if(_zz_1561_)begin
        int_reg_array_22_24_imag <= _zz_1603_;
      end
      if(_zz_1562_)begin
        int_reg_array_22_25_imag <= _zz_1603_;
      end
      if(_zz_1563_)begin
        int_reg_array_22_26_imag <= _zz_1603_;
      end
      if(_zz_1564_)begin
        int_reg_array_22_27_imag <= _zz_1603_;
      end
      if(_zz_1565_)begin
        int_reg_array_22_28_imag <= _zz_1603_;
      end
      if(_zz_1566_)begin
        int_reg_array_22_29_imag <= _zz_1603_;
      end
      if(_zz_1567_)begin
        int_reg_array_22_30_imag <= _zz_1603_;
      end
      if(_zz_1568_)begin
        int_reg_array_22_31_imag <= _zz_1603_;
      end
      if(_zz_1569_)begin
        int_reg_array_22_32_imag <= _zz_1603_;
      end
      if(_zz_1570_)begin
        int_reg_array_22_33_imag <= _zz_1603_;
      end
      if(_zz_1571_)begin
        int_reg_array_22_34_imag <= _zz_1603_;
      end
      if(_zz_1572_)begin
        int_reg_array_22_35_imag <= _zz_1603_;
      end
      if(_zz_1573_)begin
        int_reg_array_22_36_imag <= _zz_1603_;
      end
      if(_zz_1574_)begin
        int_reg_array_22_37_imag <= _zz_1603_;
      end
      if(_zz_1575_)begin
        int_reg_array_22_38_imag <= _zz_1603_;
      end
      if(_zz_1576_)begin
        int_reg_array_22_39_imag <= _zz_1603_;
      end
      if(_zz_1577_)begin
        int_reg_array_22_40_imag <= _zz_1603_;
      end
      if(_zz_1578_)begin
        int_reg_array_22_41_imag <= _zz_1603_;
      end
      if(_zz_1579_)begin
        int_reg_array_22_42_imag <= _zz_1603_;
      end
      if(_zz_1580_)begin
        int_reg_array_22_43_imag <= _zz_1603_;
      end
      if(_zz_1581_)begin
        int_reg_array_22_44_imag <= _zz_1603_;
      end
      if(_zz_1582_)begin
        int_reg_array_22_45_imag <= _zz_1603_;
      end
      if(_zz_1583_)begin
        int_reg_array_22_46_imag <= _zz_1603_;
      end
      if(_zz_1584_)begin
        int_reg_array_22_47_imag <= _zz_1603_;
      end
      if(_zz_1585_)begin
        int_reg_array_22_48_imag <= _zz_1603_;
      end
      if(_zz_1586_)begin
        int_reg_array_22_49_imag <= _zz_1603_;
      end
      if(_zz_1587_)begin
        int_reg_array_22_50_imag <= _zz_1603_;
      end
      if(_zz_1588_)begin
        int_reg_array_22_51_imag <= _zz_1603_;
      end
      if(_zz_1589_)begin
        int_reg_array_22_52_imag <= _zz_1603_;
      end
      if(_zz_1590_)begin
        int_reg_array_22_53_imag <= _zz_1603_;
      end
      if(_zz_1591_)begin
        int_reg_array_22_54_imag <= _zz_1603_;
      end
      if(_zz_1592_)begin
        int_reg_array_22_55_imag <= _zz_1603_;
      end
      if(_zz_1593_)begin
        int_reg_array_22_56_imag <= _zz_1603_;
      end
      if(_zz_1594_)begin
        int_reg_array_22_57_imag <= _zz_1603_;
      end
      if(_zz_1595_)begin
        int_reg_array_22_58_imag <= _zz_1603_;
      end
      if(_zz_1596_)begin
        int_reg_array_22_59_imag <= _zz_1603_;
      end
      if(_zz_1597_)begin
        int_reg_array_22_60_imag <= _zz_1603_;
      end
      if(_zz_1598_)begin
        int_reg_array_22_61_imag <= _zz_1603_;
      end
      if(_zz_1599_)begin
        int_reg_array_22_62_imag <= _zz_1603_;
      end
      if(_zz_1600_)begin
        int_reg_array_22_63_imag <= _zz_1603_;
      end
      if(_zz_1606_)begin
        int_reg_array_23_0_real <= _zz_1671_;
      end
      if(_zz_1607_)begin
        int_reg_array_23_1_real <= _zz_1671_;
      end
      if(_zz_1608_)begin
        int_reg_array_23_2_real <= _zz_1671_;
      end
      if(_zz_1609_)begin
        int_reg_array_23_3_real <= _zz_1671_;
      end
      if(_zz_1610_)begin
        int_reg_array_23_4_real <= _zz_1671_;
      end
      if(_zz_1611_)begin
        int_reg_array_23_5_real <= _zz_1671_;
      end
      if(_zz_1612_)begin
        int_reg_array_23_6_real <= _zz_1671_;
      end
      if(_zz_1613_)begin
        int_reg_array_23_7_real <= _zz_1671_;
      end
      if(_zz_1614_)begin
        int_reg_array_23_8_real <= _zz_1671_;
      end
      if(_zz_1615_)begin
        int_reg_array_23_9_real <= _zz_1671_;
      end
      if(_zz_1616_)begin
        int_reg_array_23_10_real <= _zz_1671_;
      end
      if(_zz_1617_)begin
        int_reg_array_23_11_real <= _zz_1671_;
      end
      if(_zz_1618_)begin
        int_reg_array_23_12_real <= _zz_1671_;
      end
      if(_zz_1619_)begin
        int_reg_array_23_13_real <= _zz_1671_;
      end
      if(_zz_1620_)begin
        int_reg_array_23_14_real <= _zz_1671_;
      end
      if(_zz_1621_)begin
        int_reg_array_23_15_real <= _zz_1671_;
      end
      if(_zz_1622_)begin
        int_reg_array_23_16_real <= _zz_1671_;
      end
      if(_zz_1623_)begin
        int_reg_array_23_17_real <= _zz_1671_;
      end
      if(_zz_1624_)begin
        int_reg_array_23_18_real <= _zz_1671_;
      end
      if(_zz_1625_)begin
        int_reg_array_23_19_real <= _zz_1671_;
      end
      if(_zz_1626_)begin
        int_reg_array_23_20_real <= _zz_1671_;
      end
      if(_zz_1627_)begin
        int_reg_array_23_21_real <= _zz_1671_;
      end
      if(_zz_1628_)begin
        int_reg_array_23_22_real <= _zz_1671_;
      end
      if(_zz_1629_)begin
        int_reg_array_23_23_real <= _zz_1671_;
      end
      if(_zz_1630_)begin
        int_reg_array_23_24_real <= _zz_1671_;
      end
      if(_zz_1631_)begin
        int_reg_array_23_25_real <= _zz_1671_;
      end
      if(_zz_1632_)begin
        int_reg_array_23_26_real <= _zz_1671_;
      end
      if(_zz_1633_)begin
        int_reg_array_23_27_real <= _zz_1671_;
      end
      if(_zz_1634_)begin
        int_reg_array_23_28_real <= _zz_1671_;
      end
      if(_zz_1635_)begin
        int_reg_array_23_29_real <= _zz_1671_;
      end
      if(_zz_1636_)begin
        int_reg_array_23_30_real <= _zz_1671_;
      end
      if(_zz_1637_)begin
        int_reg_array_23_31_real <= _zz_1671_;
      end
      if(_zz_1638_)begin
        int_reg_array_23_32_real <= _zz_1671_;
      end
      if(_zz_1639_)begin
        int_reg_array_23_33_real <= _zz_1671_;
      end
      if(_zz_1640_)begin
        int_reg_array_23_34_real <= _zz_1671_;
      end
      if(_zz_1641_)begin
        int_reg_array_23_35_real <= _zz_1671_;
      end
      if(_zz_1642_)begin
        int_reg_array_23_36_real <= _zz_1671_;
      end
      if(_zz_1643_)begin
        int_reg_array_23_37_real <= _zz_1671_;
      end
      if(_zz_1644_)begin
        int_reg_array_23_38_real <= _zz_1671_;
      end
      if(_zz_1645_)begin
        int_reg_array_23_39_real <= _zz_1671_;
      end
      if(_zz_1646_)begin
        int_reg_array_23_40_real <= _zz_1671_;
      end
      if(_zz_1647_)begin
        int_reg_array_23_41_real <= _zz_1671_;
      end
      if(_zz_1648_)begin
        int_reg_array_23_42_real <= _zz_1671_;
      end
      if(_zz_1649_)begin
        int_reg_array_23_43_real <= _zz_1671_;
      end
      if(_zz_1650_)begin
        int_reg_array_23_44_real <= _zz_1671_;
      end
      if(_zz_1651_)begin
        int_reg_array_23_45_real <= _zz_1671_;
      end
      if(_zz_1652_)begin
        int_reg_array_23_46_real <= _zz_1671_;
      end
      if(_zz_1653_)begin
        int_reg_array_23_47_real <= _zz_1671_;
      end
      if(_zz_1654_)begin
        int_reg_array_23_48_real <= _zz_1671_;
      end
      if(_zz_1655_)begin
        int_reg_array_23_49_real <= _zz_1671_;
      end
      if(_zz_1656_)begin
        int_reg_array_23_50_real <= _zz_1671_;
      end
      if(_zz_1657_)begin
        int_reg_array_23_51_real <= _zz_1671_;
      end
      if(_zz_1658_)begin
        int_reg_array_23_52_real <= _zz_1671_;
      end
      if(_zz_1659_)begin
        int_reg_array_23_53_real <= _zz_1671_;
      end
      if(_zz_1660_)begin
        int_reg_array_23_54_real <= _zz_1671_;
      end
      if(_zz_1661_)begin
        int_reg_array_23_55_real <= _zz_1671_;
      end
      if(_zz_1662_)begin
        int_reg_array_23_56_real <= _zz_1671_;
      end
      if(_zz_1663_)begin
        int_reg_array_23_57_real <= _zz_1671_;
      end
      if(_zz_1664_)begin
        int_reg_array_23_58_real <= _zz_1671_;
      end
      if(_zz_1665_)begin
        int_reg_array_23_59_real <= _zz_1671_;
      end
      if(_zz_1666_)begin
        int_reg_array_23_60_real <= _zz_1671_;
      end
      if(_zz_1667_)begin
        int_reg_array_23_61_real <= _zz_1671_;
      end
      if(_zz_1668_)begin
        int_reg_array_23_62_real <= _zz_1671_;
      end
      if(_zz_1669_)begin
        int_reg_array_23_63_real <= _zz_1671_;
      end
      if(_zz_1606_)begin
        int_reg_array_23_0_imag <= _zz_1672_;
      end
      if(_zz_1607_)begin
        int_reg_array_23_1_imag <= _zz_1672_;
      end
      if(_zz_1608_)begin
        int_reg_array_23_2_imag <= _zz_1672_;
      end
      if(_zz_1609_)begin
        int_reg_array_23_3_imag <= _zz_1672_;
      end
      if(_zz_1610_)begin
        int_reg_array_23_4_imag <= _zz_1672_;
      end
      if(_zz_1611_)begin
        int_reg_array_23_5_imag <= _zz_1672_;
      end
      if(_zz_1612_)begin
        int_reg_array_23_6_imag <= _zz_1672_;
      end
      if(_zz_1613_)begin
        int_reg_array_23_7_imag <= _zz_1672_;
      end
      if(_zz_1614_)begin
        int_reg_array_23_8_imag <= _zz_1672_;
      end
      if(_zz_1615_)begin
        int_reg_array_23_9_imag <= _zz_1672_;
      end
      if(_zz_1616_)begin
        int_reg_array_23_10_imag <= _zz_1672_;
      end
      if(_zz_1617_)begin
        int_reg_array_23_11_imag <= _zz_1672_;
      end
      if(_zz_1618_)begin
        int_reg_array_23_12_imag <= _zz_1672_;
      end
      if(_zz_1619_)begin
        int_reg_array_23_13_imag <= _zz_1672_;
      end
      if(_zz_1620_)begin
        int_reg_array_23_14_imag <= _zz_1672_;
      end
      if(_zz_1621_)begin
        int_reg_array_23_15_imag <= _zz_1672_;
      end
      if(_zz_1622_)begin
        int_reg_array_23_16_imag <= _zz_1672_;
      end
      if(_zz_1623_)begin
        int_reg_array_23_17_imag <= _zz_1672_;
      end
      if(_zz_1624_)begin
        int_reg_array_23_18_imag <= _zz_1672_;
      end
      if(_zz_1625_)begin
        int_reg_array_23_19_imag <= _zz_1672_;
      end
      if(_zz_1626_)begin
        int_reg_array_23_20_imag <= _zz_1672_;
      end
      if(_zz_1627_)begin
        int_reg_array_23_21_imag <= _zz_1672_;
      end
      if(_zz_1628_)begin
        int_reg_array_23_22_imag <= _zz_1672_;
      end
      if(_zz_1629_)begin
        int_reg_array_23_23_imag <= _zz_1672_;
      end
      if(_zz_1630_)begin
        int_reg_array_23_24_imag <= _zz_1672_;
      end
      if(_zz_1631_)begin
        int_reg_array_23_25_imag <= _zz_1672_;
      end
      if(_zz_1632_)begin
        int_reg_array_23_26_imag <= _zz_1672_;
      end
      if(_zz_1633_)begin
        int_reg_array_23_27_imag <= _zz_1672_;
      end
      if(_zz_1634_)begin
        int_reg_array_23_28_imag <= _zz_1672_;
      end
      if(_zz_1635_)begin
        int_reg_array_23_29_imag <= _zz_1672_;
      end
      if(_zz_1636_)begin
        int_reg_array_23_30_imag <= _zz_1672_;
      end
      if(_zz_1637_)begin
        int_reg_array_23_31_imag <= _zz_1672_;
      end
      if(_zz_1638_)begin
        int_reg_array_23_32_imag <= _zz_1672_;
      end
      if(_zz_1639_)begin
        int_reg_array_23_33_imag <= _zz_1672_;
      end
      if(_zz_1640_)begin
        int_reg_array_23_34_imag <= _zz_1672_;
      end
      if(_zz_1641_)begin
        int_reg_array_23_35_imag <= _zz_1672_;
      end
      if(_zz_1642_)begin
        int_reg_array_23_36_imag <= _zz_1672_;
      end
      if(_zz_1643_)begin
        int_reg_array_23_37_imag <= _zz_1672_;
      end
      if(_zz_1644_)begin
        int_reg_array_23_38_imag <= _zz_1672_;
      end
      if(_zz_1645_)begin
        int_reg_array_23_39_imag <= _zz_1672_;
      end
      if(_zz_1646_)begin
        int_reg_array_23_40_imag <= _zz_1672_;
      end
      if(_zz_1647_)begin
        int_reg_array_23_41_imag <= _zz_1672_;
      end
      if(_zz_1648_)begin
        int_reg_array_23_42_imag <= _zz_1672_;
      end
      if(_zz_1649_)begin
        int_reg_array_23_43_imag <= _zz_1672_;
      end
      if(_zz_1650_)begin
        int_reg_array_23_44_imag <= _zz_1672_;
      end
      if(_zz_1651_)begin
        int_reg_array_23_45_imag <= _zz_1672_;
      end
      if(_zz_1652_)begin
        int_reg_array_23_46_imag <= _zz_1672_;
      end
      if(_zz_1653_)begin
        int_reg_array_23_47_imag <= _zz_1672_;
      end
      if(_zz_1654_)begin
        int_reg_array_23_48_imag <= _zz_1672_;
      end
      if(_zz_1655_)begin
        int_reg_array_23_49_imag <= _zz_1672_;
      end
      if(_zz_1656_)begin
        int_reg_array_23_50_imag <= _zz_1672_;
      end
      if(_zz_1657_)begin
        int_reg_array_23_51_imag <= _zz_1672_;
      end
      if(_zz_1658_)begin
        int_reg_array_23_52_imag <= _zz_1672_;
      end
      if(_zz_1659_)begin
        int_reg_array_23_53_imag <= _zz_1672_;
      end
      if(_zz_1660_)begin
        int_reg_array_23_54_imag <= _zz_1672_;
      end
      if(_zz_1661_)begin
        int_reg_array_23_55_imag <= _zz_1672_;
      end
      if(_zz_1662_)begin
        int_reg_array_23_56_imag <= _zz_1672_;
      end
      if(_zz_1663_)begin
        int_reg_array_23_57_imag <= _zz_1672_;
      end
      if(_zz_1664_)begin
        int_reg_array_23_58_imag <= _zz_1672_;
      end
      if(_zz_1665_)begin
        int_reg_array_23_59_imag <= _zz_1672_;
      end
      if(_zz_1666_)begin
        int_reg_array_23_60_imag <= _zz_1672_;
      end
      if(_zz_1667_)begin
        int_reg_array_23_61_imag <= _zz_1672_;
      end
      if(_zz_1668_)begin
        int_reg_array_23_62_imag <= _zz_1672_;
      end
      if(_zz_1669_)begin
        int_reg_array_23_63_imag <= _zz_1672_;
      end
      if(_zz_1675_)begin
        int_reg_array_24_0_real <= _zz_1740_;
      end
      if(_zz_1676_)begin
        int_reg_array_24_1_real <= _zz_1740_;
      end
      if(_zz_1677_)begin
        int_reg_array_24_2_real <= _zz_1740_;
      end
      if(_zz_1678_)begin
        int_reg_array_24_3_real <= _zz_1740_;
      end
      if(_zz_1679_)begin
        int_reg_array_24_4_real <= _zz_1740_;
      end
      if(_zz_1680_)begin
        int_reg_array_24_5_real <= _zz_1740_;
      end
      if(_zz_1681_)begin
        int_reg_array_24_6_real <= _zz_1740_;
      end
      if(_zz_1682_)begin
        int_reg_array_24_7_real <= _zz_1740_;
      end
      if(_zz_1683_)begin
        int_reg_array_24_8_real <= _zz_1740_;
      end
      if(_zz_1684_)begin
        int_reg_array_24_9_real <= _zz_1740_;
      end
      if(_zz_1685_)begin
        int_reg_array_24_10_real <= _zz_1740_;
      end
      if(_zz_1686_)begin
        int_reg_array_24_11_real <= _zz_1740_;
      end
      if(_zz_1687_)begin
        int_reg_array_24_12_real <= _zz_1740_;
      end
      if(_zz_1688_)begin
        int_reg_array_24_13_real <= _zz_1740_;
      end
      if(_zz_1689_)begin
        int_reg_array_24_14_real <= _zz_1740_;
      end
      if(_zz_1690_)begin
        int_reg_array_24_15_real <= _zz_1740_;
      end
      if(_zz_1691_)begin
        int_reg_array_24_16_real <= _zz_1740_;
      end
      if(_zz_1692_)begin
        int_reg_array_24_17_real <= _zz_1740_;
      end
      if(_zz_1693_)begin
        int_reg_array_24_18_real <= _zz_1740_;
      end
      if(_zz_1694_)begin
        int_reg_array_24_19_real <= _zz_1740_;
      end
      if(_zz_1695_)begin
        int_reg_array_24_20_real <= _zz_1740_;
      end
      if(_zz_1696_)begin
        int_reg_array_24_21_real <= _zz_1740_;
      end
      if(_zz_1697_)begin
        int_reg_array_24_22_real <= _zz_1740_;
      end
      if(_zz_1698_)begin
        int_reg_array_24_23_real <= _zz_1740_;
      end
      if(_zz_1699_)begin
        int_reg_array_24_24_real <= _zz_1740_;
      end
      if(_zz_1700_)begin
        int_reg_array_24_25_real <= _zz_1740_;
      end
      if(_zz_1701_)begin
        int_reg_array_24_26_real <= _zz_1740_;
      end
      if(_zz_1702_)begin
        int_reg_array_24_27_real <= _zz_1740_;
      end
      if(_zz_1703_)begin
        int_reg_array_24_28_real <= _zz_1740_;
      end
      if(_zz_1704_)begin
        int_reg_array_24_29_real <= _zz_1740_;
      end
      if(_zz_1705_)begin
        int_reg_array_24_30_real <= _zz_1740_;
      end
      if(_zz_1706_)begin
        int_reg_array_24_31_real <= _zz_1740_;
      end
      if(_zz_1707_)begin
        int_reg_array_24_32_real <= _zz_1740_;
      end
      if(_zz_1708_)begin
        int_reg_array_24_33_real <= _zz_1740_;
      end
      if(_zz_1709_)begin
        int_reg_array_24_34_real <= _zz_1740_;
      end
      if(_zz_1710_)begin
        int_reg_array_24_35_real <= _zz_1740_;
      end
      if(_zz_1711_)begin
        int_reg_array_24_36_real <= _zz_1740_;
      end
      if(_zz_1712_)begin
        int_reg_array_24_37_real <= _zz_1740_;
      end
      if(_zz_1713_)begin
        int_reg_array_24_38_real <= _zz_1740_;
      end
      if(_zz_1714_)begin
        int_reg_array_24_39_real <= _zz_1740_;
      end
      if(_zz_1715_)begin
        int_reg_array_24_40_real <= _zz_1740_;
      end
      if(_zz_1716_)begin
        int_reg_array_24_41_real <= _zz_1740_;
      end
      if(_zz_1717_)begin
        int_reg_array_24_42_real <= _zz_1740_;
      end
      if(_zz_1718_)begin
        int_reg_array_24_43_real <= _zz_1740_;
      end
      if(_zz_1719_)begin
        int_reg_array_24_44_real <= _zz_1740_;
      end
      if(_zz_1720_)begin
        int_reg_array_24_45_real <= _zz_1740_;
      end
      if(_zz_1721_)begin
        int_reg_array_24_46_real <= _zz_1740_;
      end
      if(_zz_1722_)begin
        int_reg_array_24_47_real <= _zz_1740_;
      end
      if(_zz_1723_)begin
        int_reg_array_24_48_real <= _zz_1740_;
      end
      if(_zz_1724_)begin
        int_reg_array_24_49_real <= _zz_1740_;
      end
      if(_zz_1725_)begin
        int_reg_array_24_50_real <= _zz_1740_;
      end
      if(_zz_1726_)begin
        int_reg_array_24_51_real <= _zz_1740_;
      end
      if(_zz_1727_)begin
        int_reg_array_24_52_real <= _zz_1740_;
      end
      if(_zz_1728_)begin
        int_reg_array_24_53_real <= _zz_1740_;
      end
      if(_zz_1729_)begin
        int_reg_array_24_54_real <= _zz_1740_;
      end
      if(_zz_1730_)begin
        int_reg_array_24_55_real <= _zz_1740_;
      end
      if(_zz_1731_)begin
        int_reg_array_24_56_real <= _zz_1740_;
      end
      if(_zz_1732_)begin
        int_reg_array_24_57_real <= _zz_1740_;
      end
      if(_zz_1733_)begin
        int_reg_array_24_58_real <= _zz_1740_;
      end
      if(_zz_1734_)begin
        int_reg_array_24_59_real <= _zz_1740_;
      end
      if(_zz_1735_)begin
        int_reg_array_24_60_real <= _zz_1740_;
      end
      if(_zz_1736_)begin
        int_reg_array_24_61_real <= _zz_1740_;
      end
      if(_zz_1737_)begin
        int_reg_array_24_62_real <= _zz_1740_;
      end
      if(_zz_1738_)begin
        int_reg_array_24_63_real <= _zz_1740_;
      end
      if(_zz_1675_)begin
        int_reg_array_24_0_imag <= _zz_1741_;
      end
      if(_zz_1676_)begin
        int_reg_array_24_1_imag <= _zz_1741_;
      end
      if(_zz_1677_)begin
        int_reg_array_24_2_imag <= _zz_1741_;
      end
      if(_zz_1678_)begin
        int_reg_array_24_3_imag <= _zz_1741_;
      end
      if(_zz_1679_)begin
        int_reg_array_24_4_imag <= _zz_1741_;
      end
      if(_zz_1680_)begin
        int_reg_array_24_5_imag <= _zz_1741_;
      end
      if(_zz_1681_)begin
        int_reg_array_24_6_imag <= _zz_1741_;
      end
      if(_zz_1682_)begin
        int_reg_array_24_7_imag <= _zz_1741_;
      end
      if(_zz_1683_)begin
        int_reg_array_24_8_imag <= _zz_1741_;
      end
      if(_zz_1684_)begin
        int_reg_array_24_9_imag <= _zz_1741_;
      end
      if(_zz_1685_)begin
        int_reg_array_24_10_imag <= _zz_1741_;
      end
      if(_zz_1686_)begin
        int_reg_array_24_11_imag <= _zz_1741_;
      end
      if(_zz_1687_)begin
        int_reg_array_24_12_imag <= _zz_1741_;
      end
      if(_zz_1688_)begin
        int_reg_array_24_13_imag <= _zz_1741_;
      end
      if(_zz_1689_)begin
        int_reg_array_24_14_imag <= _zz_1741_;
      end
      if(_zz_1690_)begin
        int_reg_array_24_15_imag <= _zz_1741_;
      end
      if(_zz_1691_)begin
        int_reg_array_24_16_imag <= _zz_1741_;
      end
      if(_zz_1692_)begin
        int_reg_array_24_17_imag <= _zz_1741_;
      end
      if(_zz_1693_)begin
        int_reg_array_24_18_imag <= _zz_1741_;
      end
      if(_zz_1694_)begin
        int_reg_array_24_19_imag <= _zz_1741_;
      end
      if(_zz_1695_)begin
        int_reg_array_24_20_imag <= _zz_1741_;
      end
      if(_zz_1696_)begin
        int_reg_array_24_21_imag <= _zz_1741_;
      end
      if(_zz_1697_)begin
        int_reg_array_24_22_imag <= _zz_1741_;
      end
      if(_zz_1698_)begin
        int_reg_array_24_23_imag <= _zz_1741_;
      end
      if(_zz_1699_)begin
        int_reg_array_24_24_imag <= _zz_1741_;
      end
      if(_zz_1700_)begin
        int_reg_array_24_25_imag <= _zz_1741_;
      end
      if(_zz_1701_)begin
        int_reg_array_24_26_imag <= _zz_1741_;
      end
      if(_zz_1702_)begin
        int_reg_array_24_27_imag <= _zz_1741_;
      end
      if(_zz_1703_)begin
        int_reg_array_24_28_imag <= _zz_1741_;
      end
      if(_zz_1704_)begin
        int_reg_array_24_29_imag <= _zz_1741_;
      end
      if(_zz_1705_)begin
        int_reg_array_24_30_imag <= _zz_1741_;
      end
      if(_zz_1706_)begin
        int_reg_array_24_31_imag <= _zz_1741_;
      end
      if(_zz_1707_)begin
        int_reg_array_24_32_imag <= _zz_1741_;
      end
      if(_zz_1708_)begin
        int_reg_array_24_33_imag <= _zz_1741_;
      end
      if(_zz_1709_)begin
        int_reg_array_24_34_imag <= _zz_1741_;
      end
      if(_zz_1710_)begin
        int_reg_array_24_35_imag <= _zz_1741_;
      end
      if(_zz_1711_)begin
        int_reg_array_24_36_imag <= _zz_1741_;
      end
      if(_zz_1712_)begin
        int_reg_array_24_37_imag <= _zz_1741_;
      end
      if(_zz_1713_)begin
        int_reg_array_24_38_imag <= _zz_1741_;
      end
      if(_zz_1714_)begin
        int_reg_array_24_39_imag <= _zz_1741_;
      end
      if(_zz_1715_)begin
        int_reg_array_24_40_imag <= _zz_1741_;
      end
      if(_zz_1716_)begin
        int_reg_array_24_41_imag <= _zz_1741_;
      end
      if(_zz_1717_)begin
        int_reg_array_24_42_imag <= _zz_1741_;
      end
      if(_zz_1718_)begin
        int_reg_array_24_43_imag <= _zz_1741_;
      end
      if(_zz_1719_)begin
        int_reg_array_24_44_imag <= _zz_1741_;
      end
      if(_zz_1720_)begin
        int_reg_array_24_45_imag <= _zz_1741_;
      end
      if(_zz_1721_)begin
        int_reg_array_24_46_imag <= _zz_1741_;
      end
      if(_zz_1722_)begin
        int_reg_array_24_47_imag <= _zz_1741_;
      end
      if(_zz_1723_)begin
        int_reg_array_24_48_imag <= _zz_1741_;
      end
      if(_zz_1724_)begin
        int_reg_array_24_49_imag <= _zz_1741_;
      end
      if(_zz_1725_)begin
        int_reg_array_24_50_imag <= _zz_1741_;
      end
      if(_zz_1726_)begin
        int_reg_array_24_51_imag <= _zz_1741_;
      end
      if(_zz_1727_)begin
        int_reg_array_24_52_imag <= _zz_1741_;
      end
      if(_zz_1728_)begin
        int_reg_array_24_53_imag <= _zz_1741_;
      end
      if(_zz_1729_)begin
        int_reg_array_24_54_imag <= _zz_1741_;
      end
      if(_zz_1730_)begin
        int_reg_array_24_55_imag <= _zz_1741_;
      end
      if(_zz_1731_)begin
        int_reg_array_24_56_imag <= _zz_1741_;
      end
      if(_zz_1732_)begin
        int_reg_array_24_57_imag <= _zz_1741_;
      end
      if(_zz_1733_)begin
        int_reg_array_24_58_imag <= _zz_1741_;
      end
      if(_zz_1734_)begin
        int_reg_array_24_59_imag <= _zz_1741_;
      end
      if(_zz_1735_)begin
        int_reg_array_24_60_imag <= _zz_1741_;
      end
      if(_zz_1736_)begin
        int_reg_array_24_61_imag <= _zz_1741_;
      end
      if(_zz_1737_)begin
        int_reg_array_24_62_imag <= _zz_1741_;
      end
      if(_zz_1738_)begin
        int_reg_array_24_63_imag <= _zz_1741_;
      end
      if(_zz_1744_)begin
        int_reg_array_25_0_real <= _zz_1809_;
      end
      if(_zz_1745_)begin
        int_reg_array_25_1_real <= _zz_1809_;
      end
      if(_zz_1746_)begin
        int_reg_array_25_2_real <= _zz_1809_;
      end
      if(_zz_1747_)begin
        int_reg_array_25_3_real <= _zz_1809_;
      end
      if(_zz_1748_)begin
        int_reg_array_25_4_real <= _zz_1809_;
      end
      if(_zz_1749_)begin
        int_reg_array_25_5_real <= _zz_1809_;
      end
      if(_zz_1750_)begin
        int_reg_array_25_6_real <= _zz_1809_;
      end
      if(_zz_1751_)begin
        int_reg_array_25_7_real <= _zz_1809_;
      end
      if(_zz_1752_)begin
        int_reg_array_25_8_real <= _zz_1809_;
      end
      if(_zz_1753_)begin
        int_reg_array_25_9_real <= _zz_1809_;
      end
      if(_zz_1754_)begin
        int_reg_array_25_10_real <= _zz_1809_;
      end
      if(_zz_1755_)begin
        int_reg_array_25_11_real <= _zz_1809_;
      end
      if(_zz_1756_)begin
        int_reg_array_25_12_real <= _zz_1809_;
      end
      if(_zz_1757_)begin
        int_reg_array_25_13_real <= _zz_1809_;
      end
      if(_zz_1758_)begin
        int_reg_array_25_14_real <= _zz_1809_;
      end
      if(_zz_1759_)begin
        int_reg_array_25_15_real <= _zz_1809_;
      end
      if(_zz_1760_)begin
        int_reg_array_25_16_real <= _zz_1809_;
      end
      if(_zz_1761_)begin
        int_reg_array_25_17_real <= _zz_1809_;
      end
      if(_zz_1762_)begin
        int_reg_array_25_18_real <= _zz_1809_;
      end
      if(_zz_1763_)begin
        int_reg_array_25_19_real <= _zz_1809_;
      end
      if(_zz_1764_)begin
        int_reg_array_25_20_real <= _zz_1809_;
      end
      if(_zz_1765_)begin
        int_reg_array_25_21_real <= _zz_1809_;
      end
      if(_zz_1766_)begin
        int_reg_array_25_22_real <= _zz_1809_;
      end
      if(_zz_1767_)begin
        int_reg_array_25_23_real <= _zz_1809_;
      end
      if(_zz_1768_)begin
        int_reg_array_25_24_real <= _zz_1809_;
      end
      if(_zz_1769_)begin
        int_reg_array_25_25_real <= _zz_1809_;
      end
      if(_zz_1770_)begin
        int_reg_array_25_26_real <= _zz_1809_;
      end
      if(_zz_1771_)begin
        int_reg_array_25_27_real <= _zz_1809_;
      end
      if(_zz_1772_)begin
        int_reg_array_25_28_real <= _zz_1809_;
      end
      if(_zz_1773_)begin
        int_reg_array_25_29_real <= _zz_1809_;
      end
      if(_zz_1774_)begin
        int_reg_array_25_30_real <= _zz_1809_;
      end
      if(_zz_1775_)begin
        int_reg_array_25_31_real <= _zz_1809_;
      end
      if(_zz_1776_)begin
        int_reg_array_25_32_real <= _zz_1809_;
      end
      if(_zz_1777_)begin
        int_reg_array_25_33_real <= _zz_1809_;
      end
      if(_zz_1778_)begin
        int_reg_array_25_34_real <= _zz_1809_;
      end
      if(_zz_1779_)begin
        int_reg_array_25_35_real <= _zz_1809_;
      end
      if(_zz_1780_)begin
        int_reg_array_25_36_real <= _zz_1809_;
      end
      if(_zz_1781_)begin
        int_reg_array_25_37_real <= _zz_1809_;
      end
      if(_zz_1782_)begin
        int_reg_array_25_38_real <= _zz_1809_;
      end
      if(_zz_1783_)begin
        int_reg_array_25_39_real <= _zz_1809_;
      end
      if(_zz_1784_)begin
        int_reg_array_25_40_real <= _zz_1809_;
      end
      if(_zz_1785_)begin
        int_reg_array_25_41_real <= _zz_1809_;
      end
      if(_zz_1786_)begin
        int_reg_array_25_42_real <= _zz_1809_;
      end
      if(_zz_1787_)begin
        int_reg_array_25_43_real <= _zz_1809_;
      end
      if(_zz_1788_)begin
        int_reg_array_25_44_real <= _zz_1809_;
      end
      if(_zz_1789_)begin
        int_reg_array_25_45_real <= _zz_1809_;
      end
      if(_zz_1790_)begin
        int_reg_array_25_46_real <= _zz_1809_;
      end
      if(_zz_1791_)begin
        int_reg_array_25_47_real <= _zz_1809_;
      end
      if(_zz_1792_)begin
        int_reg_array_25_48_real <= _zz_1809_;
      end
      if(_zz_1793_)begin
        int_reg_array_25_49_real <= _zz_1809_;
      end
      if(_zz_1794_)begin
        int_reg_array_25_50_real <= _zz_1809_;
      end
      if(_zz_1795_)begin
        int_reg_array_25_51_real <= _zz_1809_;
      end
      if(_zz_1796_)begin
        int_reg_array_25_52_real <= _zz_1809_;
      end
      if(_zz_1797_)begin
        int_reg_array_25_53_real <= _zz_1809_;
      end
      if(_zz_1798_)begin
        int_reg_array_25_54_real <= _zz_1809_;
      end
      if(_zz_1799_)begin
        int_reg_array_25_55_real <= _zz_1809_;
      end
      if(_zz_1800_)begin
        int_reg_array_25_56_real <= _zz_1809_;
      end
      if(_zz_1801_)begin
        int_reg_array_25_57_real <= _zz_1809_;
      end
      if(_zz_1802_)begin
        int_reg_array_25_58_real <= _zz_1809_;
      end
      if(_zz_1803_)begin
        int_reg_array_25_59_real <= _zz_1809_;
      end
      if(_zz_1804_)begin
        int_reg_array_25_60_real <= _zz_1809_;
      end
      if(_zz_1805_)begin
        int_reg_array_25_61_real <= _zz_1809_;
      end
      if(_zz_1806_)begin
        int_reg_array_25_62_real <= _zz_1809_;
      end
      if(_zz_1807_)begin
        int_reg_array_25_63_real <= _zz_1809_;
      end
      if(_zz_1744_)begin
        int_reg_array_25_0_imag <= _zz_1810_;
      end
      if(_zz_1745_)begin
        int_reg_array_25_1_imag <= _zz_1810_;
      end
      if(_zz_1746_)begin
        int_reg_array_25_2_imag <= _zz_1810_;
      end
      if(_zz_1747_)begin
        int_reg_array_25_3_imag <= _zz_1810_;
      end
      if(_zz_1748_)begin
        int_reg_array_25_4_imag <= _zz_1810_;
      end
      if(_zz_1749_)begin
        int_reg_array_25_5_imag <= _zz_1810_;
      end
      if(_zz_1750_)begin
        int_reg_array_25_6_imag <= _zz_1810_;
      end
      if(_zz_1751_)begin
        int_reg_array_25_7_imag <= _zz_1810_;
      end
      if(_zz_1752_)begin
        int_reg_array_25_8_imag <= _zz_1810_;
      end
      if(_zz_1753_)begin
        int_reg_array_25_9_imag <= _zz_1810_;
      end
      if(_zz_1754_)begin
        int_reg_array_25_10_imag <= _zz_1810_;
      end
      if(_zz_1755_)begin
        int_reg_array_25_11_imag <= _zz_1810_;
      end
      if(_zz_1756_)begin
        int_reg_array_25_12_imag <= _zz_1810_;
      end
      if(_zz_1757_)begin
        int_reg_array_25_13_imag <= _zz_1810_;
      end
      if(_zz_1758_)begin
        int_reg_array_25_14_imag <= _zz_1810_;
      end
      if(_zz_1759_)begin
        int_reg_array_25_15_imag <= _zz_1810_;
      end
      if(_zz_1760_)begin
        int_reg_array_25_16_imag <= _zz_1810_;
      end
      if(_zz_1761_)begin
        int_reg_array_25_17_imag <= _zz_1810_;
      end
      if(_zz_1762_)begin
        int_reg_array_25_18_imag <= _zz_1810_;
      end
      if(_zz_1763_)begin
        int_reg_array_25_19_imag <= _zz_1810_;
      end
      if(_zz_1764_)begin
        int_reg_array_25_20_imag <= _zz_1810_;
      end
      if(_zz_1765_)begin
        int_reg_array_25_21_imag <= _zz_1810_;
      end
      if(_zz_1766_)begin
        int_reg_array_25_22_imag <= _zz_1810_;
      end
      if(_zz_1767_)begin
        int_reg_array_25_23_imag <= _zz_1810_;
      end
      if(_zz_1768_)begin
        int_reg_array_25_24_imag <= _zz_1810_;
      end
      if(_zz_1769_)begin
        int_reg_array_25_25_imag <= _zz_1810_;
      end
      if(_zz_1770_)begin
        int_reg_array_25_26_imag <= _zz_1810_;
      end
      if(_zz_1771_)begin
        int_reg_array_25_27_imag <= _zz_1810_;
      end
      if(_zz_1772_)begin
        int_reg_array_25_28_imag <= _zz_1810_;
      end
      if(_zz_1773_)begin
        int_reg_array_25_29_imag <= _zz_1810_;
      end
      if(_zz_1774_)begin
        int_reg_array_25_30_imag <= _zz_1810_;
      end
      if(_zz_1775_)begin
        int_reg_array_25_31_imag <= _zz_1810_;
      end
      if(_zz_1776_)begin
        int_reg_array_25_32_imag <= _zz_1810_;
      end
      if(_zz_1777_)begin
        int_reg_array_25_33_imag <= _zz_1810_;
      end
      if(_zz_1778_)begin
        int_reg_array_25_34_imag <= _zz_1810_;
      end
      if(_zz_1779_)begin
        int_reg_array_25_35_imag <= _zz_1810_;
      end
      if(_zz_1780_)begin
        int_reg_array_25_36_imag <= _zz_1810_;
      end
      if(_zz_1781_)begin
        int_reg_array_25_37_imag <= _zz_1810_;
      end
      if(_zz_1782_)begin
        int_reg_array_25_38_imag <= _zz_1810_;
      end
      if(_zz_1783_)begin
        int_reg_array_25_39_imag <= _zz_1810_;
      end
      if(_zz_1784_)begin
        int_reg_array_25_40_imag <= _zz_1810_;
      end
      if(_zz_1785_)begin
        int_reg_array_25_41_imag <= _zz_1810_;
      end
      if(_zz_1786_)begin
        int_reg_array_25_42_imag <= _zz_1810_;
      end
      if(_zz_1787_)begin
        int_reg_array_25_43_imag <= _zz_1810_;
      end
      if(_zz_1788_)begin
        int_reg_array_25_44_imag <= _zz_1810_;
      end
      if(_zz_1789_)begin
        int_reg_array_25_45_imag <= _zz_1810_;
      end
      if(_zz_1790_)begin
        int_reg_array_25_46_imag <= _zz_1810_;
      end
      if(_zz_1791_)begin
        int_reg_array_25_47_imag <= _zz_1810_;
      end
      if(_zz_1792_)begin
        int_reg_array_25_48_imag <= _zz_1810_;
      end
      if(_zz_1793_)begin
        int_reg_array_25_49_imag <= _zz_1810_;
      end
      if(_zz_1794_)begin
        int_reg_array_25_50_imag <= _zz_1810_;
      end
      if(_zz_1795_)begin
        int_reg_array_25_51_imag <= _zz_1810_;
      end
      if(_zz_1796_)begin
        int_reg_array_25_52_imag <= _zz_1810_;
      end
      if(_zz_1797_)begin
        int_reg_array_25_53_imag <= _zz_1810_;
      end
      if(_zz_1798_)begin
        int_reg_array_25_54_imag <= _zz_1810_;
      end
      if(_zz_1799_)begin
        int_reg_array_25_55_imag <= _zz_1810_;
      end
      if(_zz_1800_)begin
        int_reg_array_25_56_imag <= _zz_1810_;
      end
      if(_zz_1801_)begin
        int_reg_array_25_57_imag <= _zz_1810_;
      end
      if(_zz_1802_)begin
        int_reg_array_25_58_imag <= _zz_1810_;
      end
      if(_zz_1803_)begin
        int_reg_array_25_59_imag <= _zz_1810_;
      end
      if(_zz_1804_)begin
        int_reg_array_25_60_imag <= _zz_1810_;
      end
      if(_zz_1805_)begin
        int_reg_array_25_61_imag <= _zz_1810_;
      end
      if(_zz_1806_)begin
        int_reg_array_25_62_imag <= _zz_1810_;
      end
      if(_zz_1807_)begin
        int_reg_array_25_63_imag <= _zz_1810_;
      end
      if(_zz_1813_)begin
        int_reg_array_26_0_real <= _zz_1878_;
      end
      if(_zz_1814_)begin
        int_reg_array_26_1_real <= _zz_1878_;
      end
      if(_zz_1815_)begin
        int_reg_array_26_2_real <= _zz_1878_;
      end
      if(_zz_1816_)begin
        int_reg_array_26_3_real <= _zz_1878_;
      end
      if(_zz_1817_)begin
        int_reg_array_26_4_real <= _zz_1878_;
      end
      if(_zz_1818_)begin
        int_reg_array_26_5_real <= _zz_1878_;
      end
      if(_zz_1819_)begin
        int_reg_array_26_6_real <= _zz_1878_;
      end
      if(_zz_1820_)begin
        int_reg_array_26_7_real <= _zz_1878_;
      end
      if(_zz_1821_)begin
        int_reg_array_26_8_real <= _zz_1878_;
      end
      if(_zz_1822_)begin
        int_reg_array_26_9_real <= _zz_1878_;
      end
      if(_zz_1823_)begin
        int_reg_array_26_10_real <= _zz_1878_;
      end
      if(_zz_1824_)begin
        int_reg_array_26_11_real <= _zz_1878_;
      end
      if(_zz_1825_)begin
        int_reg_array_26_12_real <= _zz_1878_;
      end
      if(_zz_1826_)begin
        int_reg_array_26_13_real <= _zz_1878_;
      end
      if(_zz_1827_)begin
        int_reg_array_26_14_real <= _zz_1878_;
      end
      if(_zz_1828_)begin
        int_reg_array_26_15_real <= _zz_1878_;
      end
      if(_zz_1829_)begin
        int_reg_array_26_16_real <= _zz_1878_;
      end
      if(_zz_1830_)begin
        int_reg_array_26_17_real <= _zz_1878_;
      end
      if(_zz_1831_)begin
        int_reg_array_26_18_real <= _zz_1878_;
      end
      if(_zz_1832_)begin
        int_reg_array_26_19_real <= _zz_1878_;
      end
      if(_zz_1833_)begin
        int_reg_array_26_20_real <= _zz_1878_;
      end
      if(_zz_1834_)begin
        int_reg_array_26_21_real <= _zz_1878_;
      end
      if(_zz_1835_)begin
        int_reg_array_26_22_real <= _zz_1878_;
      end
      if(_zz_1836_)begin
        int_reg_array_26_23_real <= _zz_1878_;
      end
      if(_zz_1837_)begin
        int_reg_array_26_24_real <= _zz_1878_;
      end
      if(_zz_1838_)begin
        int_reg_array_26_25_real <= _zz_1878_;
      end
      if(_zz_1839_)begin
        int_reg_array_26_26_real <= _zz_1878_;
      end
      if(_zz_1840_)begin
        int_reg_array_26_27_real <= _zz_1878_;
      end
      if(_zz_1841_)begin
        int_reg_array_26_28_real <= _zz_1878_;
      end
      if(_zz_1842_)begin
        int_reg_array_26_29_real <= _zz_1878_;
      end
      if(_zz_1843_)begin
        int_reg_array_26_30_real <= _zz_1878_;
      end
      if(_zz_1844_)begin
        int_reg_array_26_31_real <= _zz_1878_;
      end
      if(_zz_1845_)begin
        int_reg_array_26_32_real <= _zz_1878_;
      end
      if(_zz_1846_)begin
        int_reg_array_26_33_real <= _zz_1878_;
      end
      if(_zz_1847_)begin
        int_reg_array_26_34_real <= _zz_1878_;
      end
      if(_zz_1848_)begin
        int_reg_array_26_35_real <= _zz_1878_;
      end
      if(_zz_1849_)begin
        int_reg_array_26_36_real <= _zz_1878_;
      end
      if(_zz_1850_)begin
        int_reg_array_26_37_real <= _zz_1878_;
      end
      if(_zz_1851_)begin
        int_reg_array_26_38_real <= _zz_1878_;
      end
      if(_zz_1852_)begin
        int_reg_array_26_39_real <= _zz_1878_;
      end
      if(_zz_1853_)begin
        int_reg_array_26_40_real <= _zz_1878_;
      end
      if(_zz_1854_)begin
        int_reg_array_26_41_real <= _zz_1878_;
      end
      if(_zz_1855_)begin
        int_reg_array_26_42_real <= _zz_1878_;
      end
      if(_zz_1856_)begin
        int_reg_array_26_43_real <= _zz_1878_;
      end
      if(_zz_1857_)begin
        int_reg_array_26_44_real <= _zz_1878_;
      end
      if(_zz_1858_)begin
        int_reg_array_26_45_real <= _zz_1878_;
      end
      if(_zz_1859_)begin
        int_reg_array_26_46_real <= _zz_1878_;
      end
      if(_zz_1860_)begin
        int_reg_array_26_47_real <= _zz_1878_;
      end
      if(_zz_1861_)begin
        int_reg_array_26_48_real <= _zz_1878_;
      end
      if(_zz_1862_)begin
        int_reg_array_26_49_real <= _zz_1878_;
      end
      if(_zz_1863_)begin
        int_reg_array_26_50_real <= _zz_1878_;
      end
      if(_zz_1864_)begin
        int_reg_array_26_51_real <= _zz_1878_;
      end
      if(_zz_1865_)begin
        int_reg_array_26_52_real <= _zz_1878_;
      end
      if(_zz_1866_)begin
        int_reg_array_26_53_real <= _zz_1878_;
      end
      if(_zz_1867_)begin
        int_reg_array_26_54_real <= _zz_1878_;
      end
      if(_zz_1868_)begin
        int_reg_array_26_55_real <= _zz_1878_;
      end
      if(_zz_1869_)begin
        int_reg_array_26_56_real <= _zz_1878_;
      end
      if(_zz_1870_)begin
        int_reg_array_26_57_real <= _zz_1878_;
      end
      if(_zz_1871_)begin
        int_reg_array_26_58_real <= _zz_1878_;
      end
      if(_zz_1872_)begin
        int_reg_array_26_59_real <= _zz_1878_;
      end
      if(_zz_1873_)begin
        int_reg_array_26_60_real <= _zz_1878_;
      end
      if(_zz_1874_)begin
        int_reg_array_26_61_real <= _zz_1878_;
      end
      if(_zz_1875_)begin
        int_reg_array_26_62_real <= _zz_1878_;
      end
      if(_zz_1876_)begin
        int_reg_array_26_63_real <= _zz_1878_;
      end
      if(_zz_1813_)begin
        int_reg_array_26_0_imag <= _zz_1879_;
      end
      if(_zz_1814_)begin
        int_reg_array_26_1_imag <= _zz_1879_;
      end
      if(_zz_1815_)begin
        int_reg_array_26_2_imag <= _zz_1879_;
      end
      if(_zz_1816_)begin
        int_reg_array_26_3_imag <= _zz_1879_;
      end
      if(_zz_1817_)begin
        int_reg_array_26_4_imag <= _zz_1879_;
      end
      if(_zz_1818_)begin
        int_reg_array_26_5_imag <= _zz_1879_;
      end
      if(_zz_1819_)begin
        int_reg_array_26_6_imag <= _zz_1879_;
      end
      if(_zz_1820_)begin
        int_reg_array_26_7_imag <= _zz_1879_;
      end
      if(_zz_1821_)begin
        int_reg_array_26_8_imag <= _zz_1879_;
      end
      if(_zz_1822_)begin
        int_reg_array_26_9_imag <= _zz_1879_;
      end
      if(_zz_1823_)begin
        int_reg_array_26_10_imag <= _zz_1879_;
      end
      if(_zz_1824_)begin
        int_reg_array_26_11_imag <= _zz_1879_;
      end
      if(_zz_1825_)begin
        int_reg_array_26_12_imag <= _zz_1879_;
      end
      if(_zz_1826_)begin
        int_reg_array_26_13_imag <= _zz_1879_;
      end
      if(_zz_1827_)begin
        int_reg_array_26_14_imag <= _zz_1879_;
      end
      if(_zz_1828_)begin
        int_reg_array_26_15_imag <= _zz_1879_;
      end
      if(_zz_1829_)begin
        int_reg_array_26_16_imag <= _zz_1879_;
      end
      if(_zz_1830_)begin
        int_reg_array_26_17_imag <= _zz_1879_;
      end
      if(_zz_1831_)begin
        int_reg_array_26_18_imag <= _zz_1879_;
      end
      if(_zz_1832_)begin
        int_reg_array_26_19_imag <= _zz_1879_;
      end
      if(_zz_1833_)begin
        int_reg_array_26_20_imag <= _zz_1879_;
      end
      if(_zz_1834_)begin
        int_reg_array_26_21_imag <= _zz_1879_;
      end
      if(_zz_1835_)begin
        int_reg_array_26_22_imag <= _zz_1879_;
      end
      if(_zz_1836_)begin
        int_reg_array_26_23_imag <= _zz_1879_;
      end
      if(_zz_1837_)begin
        int_reg_array_26_24_imag <= _zz_1879_;
      end
      if(_zz_1838_)begin
        int_reg_array_26_25_imag <= _zz_1879_;
      end
      if(_zz_1839_)begin
        int_reg_array_26_26_imag <= _zz_1879_;
      end
      if(_zz_1840_)begin
        int_reg_array_26_27_imag <= _zz_1879_;
      end
      if(_zz_1841_)begin
        int_reg_array_26_28_imag <= _zz_1879_;
      end
      if(_zz_1842_)begin
        int_reg_array_26_29_imag <= _zz_1879_;
      end
      if(_zz_1843_)begin
        int_reg_array_26_30_imag <= _zz_1879_;
      end
      if(_zz_1844_)begin
        int_reg_array_26_31_imag <= _zz_1879_;
      end
      if(_zz_1845_)begin
        int_reg_array_26_32_imag <= _zz_1879_;
      end
      if(_zz_1846_)begin
        int_reg_array_26_33_imag <= _zz_1879_;
      end
      if(_zz_1847_)begin
        int_reg_array_26_34_imag <= _zz_1879_;
      end
      if(_zz_1848_)begin
        int_reg_array_26_35_imag <= _zz_1879_;
      end
      if(_zz_1849_)begin
        int_reg_array_26_36_imag <= _zz_1879_;
      end
      if(_zz_1850_)begin
        int_reg_array_26_37_imag <= _zz_1879_;
      end
      if(_zz_1851_)begin
        int_reg_array_26_38_imag <= _zz_1879_;
      end
      if(_zz_1852_)begin
        int_reg_array_26_39_imag <= _zz_1879_;
      end
      if(_zz_1853_)begin
        int_reg_array_26_40_imag <= _zz_1879_;
      end
      if(_zz_1854_)begin
        int_reg_array_26_41_imag <= _zz_1879_;
      end
      if(_zz_1855_)begin
        int_reg_array_26_42_imag <= _zz_1879_;
      end
      if(_zz_1856_)begin
        int_reg_array_26_43_imag <= _zz_1879_;
      end
      if(_zz_1857_)begin
        int_reg_array_26_44_imag <= _zz_1879_;
      end
      if(_zz_1858_)begin
        int_reg_array_26_45_imag <= _zz_1879_;
      end
      if(_zz_1859_)begin
        int_reg_array_26_46_imag <= _zz_1879_;
      end
      if(_zz_1860_)begin
        int_reg_array_26_47_imag <= _zz_1879_;
      end
      if(_zz_1861_)begin
        int_reg_array_26_48_imag <= _zz_1879_;
      end
      if(_zz_1862_)begin
        int_reg_array_26_49_imag <= _zz_1879_;
      end
      if(_zz_1863_)begin
        int_reg_array_26_50_imag <= _zz_1879_;
      end
      if(_zz_1864_)begin
        int_reg_array_26_51_imag <= _zz_1879_;
      end
      if(_zz_1865_)begin
        int_reg_array_26_52_imag <= _zz_1879_;
      end
      if(_zz_1866_)begin
        int_reg_array_26_53_imag <= _zz_1879_;
      end
      if(_zz_1867_)begin
        int_reg_array_26_54_imag <= _zz_1879_;
      end
      if(_zz_1868_)begin
        int_reg_array_26_55_imag <= _zz_1879_;
      end
      if(_zz_1869_)begin
        int_reg_array_26_56_imag <= _zz_1879_;
      end
      if(_zz_1870_)begin
        int_reg_array_26_57_imag <= _zz_1879_;
      end
      if(_zz_1871_)begin
        int_reg_array_26_58_imag <= _zz_1879_;
      end
      if(_zz_1872_)begin
        int_reg_array_26_59_imag <= _zz_1879_;
      end
      if(_zz_1873_)begin
        int_reg_array_26_60_imag <= _zz_1879_;
      end
      if(_zz_1874_)begin
        int_reg_array_26_61_imag <= _zz_1879_;
      end
      if(_zz_1875_)begin
        int_reg_array_26_62_imag <= _zz_1879_;
      end
      if(_zz_1876_)begin
        int_reg_array_26_63_imag <= _zz_1879_;
      end
      if(_zz_1882_)begin
        int_reg_array_27_0_real <= _zz_1947_;
      end
      if(_zz_1883_)begin
        int_reg_array_27_1_real <= _zz_1947_;
      end
      if(_zz_1884_)begin
        int_reg_array_27_2_real <= _zz_1947_;
      end
      if(_zz_1885_)begin
        int_reg_array_27_3_real <= _zz_1947_;
      end
      if(_zz_1886_)begin
        int_reg_array_27_4_real <= _zz_1947_;
      end
      if(_zz_1887_)begin
        int_reg_array_27_5_real <= _zz_1947_;
      end
      if(_zz_1888_)begin
        int_reg_array_27_6_real <= _zz_1947_;
      end
      if(_zz_1889_)begin
        int_reg_array_27_7_real <= _zz_1947_;
      end
      if(_zz_1890_)begin
        int_reg_array_27_8_real <= _zz_1947_;
      end
      if(_zz_1891_)begin
        int_reg_array_27_9_real <= _zz_1947_;
      end
      if(_zz_1892_)begin
        int_reg_array_27_10_real <= _zz_1947_;
      end
      if(_zz_1893_)begin
        int_reg_array_27_11_real <= _zz_1947_;
      end
      if(_zz_1894_)begin
        int_reg_array_27_12_real <= _zz_1947_;
      end
      if(_zz_1895_)begin
        int_reg_array_27_13_real <= _zz_1947_;
      end
      if(_zz_1896_)begin
        int_reg_array_27_14_real <= _zz_1947_;
      end
      if(_zz_1897_)begin
        int_reg_array_27_15_real <= _zz_1947_;
      end
      if(_zz_1898_)begin
        int_reg_array_27_16_real <= _zz_1947_;
      end
      if(_zz_1899_)begin
        int_reg_array_27_17_real <= _zz_1947_;
      end
      if(_zz_1900_)begin
        int_reg_array_27_18_real <= _zz_1947_;
      end
      if(_zz_1901_)begin
        int_reg_array_27_19_real <= _zz_1947_;
      end
      if(_zz_1902_)begin
        int_reg_array_27_20_real <= _zz_1947_;
      end
      if(_zz_1903_)begin
        int_reg_array_27_21_real <= _zz_1947_;
      end
      if(_zz_1904_)begin
        int_reg_array_27_22_real <= _zz_1947_;
      end
      if(_zz_1905_)begin
        int_reg_array_27_23_real <= _zz_1947_;
      end
      if(_zz_1906_)begin
        int_reg_array_27_24_real <= _zz_1947_;
      end
      if(_zz_1907_)begin
        int_reg_array_27_25_real <= _zz_1947_;
      end
      if(_zz_1908_)begin
        int_reg_array_27_26_real <= _zz_1947_;
      end
      if(_zz_1909_)begin
        int_reg_array_27_27_real <= _zz_1947_;
      end
      if(_zz_1910_)begin
        int_reg_array_27_28_real <= _zz_1947_;
      end
      if(_zz_1911_)begin
        int_reg_array_27_29_real <= _zz_1947_;
      end
      if(_zz_1912_)begin
        int_reg_array_27_30_real <= _zz_1947_;
      end
      if(_zz_1913_)begin
        int_reg_array_27_31_real <= _zz_1947_;
      end
      if(_zz_1914_)begin
        int_reg_array_27_32_real <= _zz_1947_;
      end
      if(_zz_1915_)begin
        int_reg_array_27_33_real <= _zz_1947_;
      end
      if(_zz_1916_)begin
        int_reg_array_27_34_real <= _zz_1947_;
      end
      if(_zz_1917_)begin
        int_reg_array_27_35_real <= _zz_1947_;
      end
      if(_zz_1918_)begin
        int_reg_array_27_36_real <= _zz_1947_;
      end
      if(_zz_1919_)begin
        int_reg_array_27_37_real <= _zz_1947_;
      end
      if(_zz_1920_)begin
        int_reg_array_27_38_real <= _zz_1947_;
      end
      if(_zz_1921_)begin
        int_reg_array_27_39_real <= _zz_1947_;
      end
      if(_zz_1922_)begin
        int_reg_array_27_40_real <= _zz_1947_;
      end
      if(_zz_1923_)begin
        int_reg_array_27_41_real <= _zz_1947_;
      end
      if(_zz_1924_)begin
        int_reg_array_27_42_real <= _zz_1947_;
      end
      if(_zz_1925_)begin
        int_reg_array_27_43_real <= _zz_1947_;
      end
      if(_zz_1926_)begin
        int_reg_array_27_44_real <= _zz_1947_;
      end
      if(_zz_1927_)begin
        int_reg_array_27_45_real <= _zz_1947_;
      end
      if(_zz_1928_)begin
        int_reg_array_27_46_real <= _zz_1947_;
      end
      if(_zz_1929_)begin
        int_reg_array_27_47_real <= _zz_1947_;
      end
      if(_zz_1930_)begin
        int_reg_array_27_48_real <= _zz_1947_;
      end
      if(_zz_1931_)begin
        int_reg_array_27_49_real <= _zz_1947_;
      end
      if(_zz_1932_)begin
        int_reg_array_27_50_real <= _zz_1947_;
      end
      if(_zz_1933_)begin
        int_reg_array_27_51_real <= _zz_1947_;
      end
      if(_zz_1934_)begin
        int_reg_array_27_52_real <= _zz_1947_;
      end
      if(_zz_1935_)begin
        int_reg_array_27_53_real <= _zz_1947_;
      end
      if(_zz_1936_)begin
        int_reg_array_27_54_real <= _zz_1947_;
      end
      if(_zz_1937_)begin
        int_reg_array_27_55_real <= _zz_1947_;
      end
      if(_zz_1938_)begin
        int_reg_array_27_56_real <= _zz_1947_;
      end
      if(_zz_1939_)begin
        int_reg_array_27_57_real <= _zz_1947_;
      end
      if(_zz_1940_)begin
        int_reg_array_27_58_real <= _zz_1947_;
      end
      if(_zz_1941_)begin
        int_reg_array_27_59_real <= _zz_1947_;
      end
      if(_zz_1942_)begin
        int_reg_array_27_60_real <= _zz_1947_;
      end
      if(_zz_1943_)begin
        int_reg_array_27_61_real <= _zz_1947_;
      end
      if(_zz_1944_)begin
        int_reg_array_27_62_real <= _zz_1947_;
      end
      if(_zz_1945_)begin
        int_reg_array_27_63_real <= _zz_1947_;
      end
      if(_zz_1882_)begin
        int_reg_array_27_0_imag <= _zz_1948_;
      end
      if(_zz_1883_)begin
        int_reg_array_27_1_imag <= _zz_1948_;
      end
      if(_zz_1884_)begin
        int_reg_array_27_2_imag <= _zz_1948_;
      end
      if(_zz_1885_)begin
        int_reg_array_27_3_imag <= _zz_1948_;
      end
      if(_zz_1886_)begin
        int_reg_array_27_4_imag <= _zz_1948_;
      end
      if(_zz_1887_)begin
        int_reg_array_27_5_imag <= _zz_1948_;
      end
      if(_zz_1888_)begin
        int_reg_array_27_6_imag <= _zz_1948_;
      end
      if(_zz_1889_)begin
        int_reg_array_27_7_imag <= _zz_1948_;
      end
      if(_zz_1890_)begin
        int_reg_array_27_8_imag <= _zz_1948_;
      end
      if(_zz_1891_)begin
        int_reg_array_27_9_imag <= _zz_1948_;
      end
      if(_zz_1892_)begin
        int_reg_array_27_10_imag <= _zz_1948_;
      end
      if(_zz_1893_)begin
        int_reg_array_27_11_imag <= _zz_1948_;
      end
      if(_zz_1894_)begin
        int_reg_array_27_12_imag <= _zz_1948_;
      end
      if(_zz_1895_)begin
        int_reg_array_27_13_imag <= _zz_1948_;
      end
      if(_zz_1896_)begin
        int_reg_array_27_14_imag <= _zz_1948_;
      end
      if(_zz_1897_)begin
        int_reg_array_27_15_imag <= _zz_1948_;
      end
      if(_zz_1898_)begin
        int_reg_array_27_16_imag <= _zz_1948_;
      end
      if(_zz_1899_)begin
        int_reg_array_27_17_imag <= _zz_1948_;
      end
      if(_zz_1900_)begin
        int_reg_array_27_18_imag <= _zz_1948_;
      end
      if(_zz_1901_)begin
        int_reg_array_27_19_imag <= _zz_1948_;
      end
      if(_zz_1902_)begin
        int_reg_array_27_20_imag <= _zz_1948_;
      end
      if(_zz_1903_)begin
        int_reg_array_27_21_imag <= _zz_1948_;
      end
      if(_zz_1904_)begin
        int_reg_array_27_22_imag <= _zz_1948_;
      end
      if(_zz_1905_)begin
        int_reg_array_27_23_imag <= _zz_1948_;
      end
      if(_zz_1906_)begin
        int_reg_array_27_24_imag <= _zz_1948_;
      end
      if(_zz_1907_)begin
        int_reg_array_27_25_imag <= _zz_1948_;
      end
      if(_zz_1908_)begin
        int_reg_array_27_26_imag <= _zz_1948_;
      end
      if(_zz_1909_)begin
        int_reg_array_27_27_imag <= _zz_1948_;
      end
      if(_zz_1910_)begin
        int_reg_array_27_28_imag <= _zz_1948_;
      end
      if(_zz_1911_)begin
        int_reg_array_27_29_imag <= _zz_1948_;
      end
      if(_zz_1912_)begin
        int_reg_array_27_30_imag <= _zz_1948_;
      end
      if(_zz_1913_)begin
        int_reg_array_27_31_imag <= _zz_1948_;
      end
      if(_zz_1914_)begin
        int_reg_array_27_32_imag <= _zz_1948_;
      end
      if(_zz_1915_)begin
        int_reg_array_27_33_imag <= _zz_1948_;
      end
      if(_zz_1916_)begin
        int_reg_array_27_34_imag <= _zz_1948_;
      end
      if(_zz_1917_)begin
        int_reg_array_27_35_imag <= _zz_1948_;
      end
      if(_zz_1918_)begin
        int_reg_array_27_36_imag <= _zz_1948_;
      end
      if(_zz_1919_)begin
        int_reg_array_27_37_imag <= _zz_1948_;
      end
      if(_zz_1920_)begin
        int_reg_array_27_38_imag <= _zz_1948_;
      end
      if(_zz_1921_)begin
        int_reg_array_27_39_imag <= _zz_1948_;
      end
      if(_zz_1922_)begin
        int_reg_array_27_40_imag <= _zz_1948_;
      end
      if(_zz_1923_)begin
        int_reg_array_27_41_imag <= _zz_1948_;
      end
      if(_zz_1924_)begin
        int_reg_array_27_42_imag <= _zz_1948_;
      end
      if(_zz_1925_)begin
        int_reg_array_27_43_imag <= _zz_1948_;
      end
      if(_zz_1926_)begin
        int_reg_array_27_44_imag <= _zz_1948_;
      end
      if(_zz_1927_)begin
        int_reg_array_27_45_imag <= _zz_1948_;
      end
      if(_zz_1928_)begin
        int_reg_array_27_46_imag <= _zz_1948_;
      end
      if(_zz_1929_)begin
        int_reg_array_27_47_imag <= _zz_1948_;
      end
      if(_zz_1930_)begin
        int_reg_array_27_48_imag <= _zz_1948_;
      end
      if(_zz_1931_)begin
        int_reg_array_27_49_imag <= _zz_1948_;
      end
      if(_zz_1932_)begin
        int_reg_array_27_50_imag <= _zz_1948_;
      end
      if(_zz_1933_)begin
        int_reg_array_27_51_imag <= _zz_1948_;
      end
      if(_zz_1934_)begin
        int_reg_array_27_52_imag <= _zz_1948_;
      end
      if(_zz_1935_)begin
        int_reg_array_27_53_imag <= _zz_1948_;
      end
      if(_zz_1936_)begin
        int_reg_array_27_54_imag <= _zz_1948_;
      end
      if(_zz_1937_)begin
        int_reg_array_27_55_imag <= _zz_1948_;
      end
      if(_zz_1938_)begin
        int_reg_array_27_56_imag <= _zz_1948_;
      end
      if(_zz_1939_)begin
        int_reg_array_27_57_imag <= _zz_1948_;
      end
      if(_zz_1940_)begin
        int_reg_array_27_58_imag <= _zz_1948_;
      end
      if(_zz_1941_)begin
        int_reg_array_27_59_imag <= _zz_1948_;
      end
      if(_zz_1942_)begin
        int_reg_array_27_60_imag <= _zz_1948_;
      end
      if(_zz_1943_)begin
        int_reg_array_27_61_imag <= _zz_1948_;
      end
      if(_zz_1944_)begin
        int_reg_array_27_62_imag <= _zz_1948_;
      end
      if(_zz_1945_)begin
        int_reg_array_27_63_imag <= _zz_1948_;
      end
      if(_zz_1951_)begin
        int_reg_array_28_0_real <= _zz_2016_;
      end
      if(_zz_1952_)begin
        int_reg_array_28_1_real <= _zz_2016_;
      end
      if(_zz_1953_)begin
        int_reg_array_28_2_real <= _zz_2016_;
      end
      if(_zz_1954_)begin
        int_reg_array_28_3_real <= _zz_2016_;
      end
      if(_zz_1955_)begin
        int_reg_array_28_4_real <= _zz_2016_;
      end
      if(_zz_1956_)begin
        int_reg_array_28_5_real <= _zz_2016_;
      end
      if(_zz_1957_)begin
        int_reg_array_28_6_real <= _zz_2016_;
      end
      if(_zz_1958_)begin
        int_reg_array_28_7_real <= _zz_2016_;
      end
      if(_zz_1959_)begin
        int_reg_array_28_8_real <= _zz_2016_;
      end
      if(_zz_1960_)begin
        int_reg_array_28_9_real <= _zz_2016_;
      end
      if(_zz_1961_)begin
        int_reg_array_28_10_real <= _zz_2016_;
      end
      if(_zz_1962_)begin
        int_reg_array_28_11_real <= _zz_2016_;
      end
      if(_zz_1963_)begin
        int_reg_array_28_12_real <= _zz_2016_;
      end
      if(_zz_1964_)begin
        int_reg_array_28_13_real <= _zz_2016_;
      end
      if(_zz_1965_)begin
        int_reg_array_28_14_real <= _zz_2016_;
      end
      if(_zz_1966_)begin
        int_reg_array_28_15_real <= _zz_2016_;
      end
      if(_zz_1967_)begin
        int_reg_array_28_16_real <= _zz_2016_;
      end
      if(_zz_1968_)begin
        int_reg_array_28_17_real <= _zz_2016_;
      end
      if(_zz_1969_)begin
        int_reg_array_28_18_real <= _zz_2016_;
      end
      if(_zz_1970_)begin
        int_reg_array_28_19_real <= _zz_2016_;
      end
      if(_zz_1971_)begin
        int_reg_array_28_20_real <= _zz_2016_;
      end
      if(_zz_1972_)begin
        int_reg_array_28_21_real <= _zz_2016_;
      end
      if(_zz_1973_)begin
        int_reg_array_28_22_real <= _zz_2016_;
      end
      if(_zz_1974_)begin
        int_reg_array_28_23_real <= _zz_2016_;
      end
      if(_zz_1975_)begin
        int_reg_array_28_24_real <= _zz_2016_;
      end
      if(_zz_1976_)begin
        int_reg_array_28_25_real <= _zz_2016_;
      end
      if(_zz_1977_)begin
        int_reg_array_28_26_real <= _zz_2016_;
      end
      if(_zz_1978_)begin
        int_reg_array_28_27_real <= _zz_2016_;
      end
      if(_zz_1979_)begin
        int_reg_array_28_28_real <= _zz_2016_;
      end
      if(_zz_1980_)begin
        int_reg_array_28_29_real <= _zz_2016_;
      end
      if(_zz_1981_)begin
        int_reg_array_28_30_real <= _zz_2016_;
      end
      if(_zz_1982_)begin
        int_reg_array_28_31_real <= _zz_2016_;
      end
      if(_zz_1983_)begin
        int_reg_array_28_32_real <= _zz_2016_;
      end
      if(_zz_1984_)begin
        int_reg_array_28_33_real <= _zz_2016_;
      end
      if(_zz_1985_)begin
        int_reg_array_28_34_real <= _zz_2016_;
      end
      if(_zz_1986_)begin
        int_reg_array_28_35_real <= _zz_2016_;
      end
      if(_zz_1987_)begin
        int_reg_array_28_36_real <= _zz_2016_;
      end
      if(_zz_1988_)begin
        int_reg_array_28_37_real <= _zz_2016_;
      end
      if(_zz_1989_)begin
        int_reg_array_28_38_real <= _zz_2016_;
      end
      if(_zz_1990_)begin
        int_reg_array_28_39_real <= _zz_2016_;
      end
      if(_zz_1991_)begin
        int_reg_array_28_40_real <= _zz_2016_;
      end
      if(_zz_1992_)begin
        int_reg_array_28_41_real <= _zz_2016_;
      end
      if(_zz_1993_)begin
        int_reg_array_28_42_real <= _zz_2016_;
      end
      if(_zz_1994_)begin
        int_reg_array_28_43_real <= _zz_2016_;
      end
      if(_zz_1995_)begin
        int_reg_array_28_44_real <= _zz_2016_;
      end
      if(_zz_1996_)begin
        int_reg_array_28_45_real <= _zz_2016_;
      end
      if(_zz_1997_)begin
        int_reg_array_28_46_real <= _zz_2016_;
      end
      if(_zz_1998_)begin
        int_reg_array_28_47_real <= _zz_2016_;
      end
      if(_zz_1999_)begin
        int_reg_array_28_48_real <= _zz_2016_;
      end
      if(_zz_2000_)begin
        int_reg_array_28_49_real <= _zz_2016_;
      end
      if(_zz_2001_)begin
        int_reg_array_28_50_real <= _zz_2016_;
      end
      if(_zz_2002_)begin
        int_reg_array_28_51_real <= _zz_2016_;
      end
      if(_zz_2003_)begin
        int_reg_array_28_52_real <= _zz_2016_;
      end
      if(_zz_2004_)begin
        int_reg_array_28_53_real <= _zz_2016_;
      end
      if(_zz_2005_)begin
        int_reg_array_28_54_real <= _zz_2016_;
      end
      if(_zz_2006_)begin
        int_reg_array_28_55_real <= _zz_2016_;
      end
      if(_zz_2007_)begin
        int_reg_array_28_56_real <= _zz_2016_;
      end
      if(_zz_2008_)begin
        int_reg_array_28_57_real <= _zz_2016_;
      end
      if(_zz_2009_)begin
        int_reg_array_28_58_real <= _zz_2016_;
      end
      if(_zz_2010_)begin
        int_reg_array_28_59_real <= _zz_2016_;
      end
      if(_zz_2011_)begin
        int_reg_array_28_60_real <= _zz_2016_;
      end
      if(_zz_2012_)begin
        int_reg_array_28_61_real <= _zz_2016_;
      end
      if(_zz_2013_)begin
        int_reg_array_28_62_real <= _zz_2016_;
      end
      if(_zz_2014_)begin
        int_reg_array_28_63_real <= _zz_2016_;
      end
      if(_zz_1951_)begin
        int_reg_array_28_0_imag <= _zz_2017_;
      end
      if(_zz_1952_)begin
        int_reg_array_28_1_imag <= _zz_2017_;
      end
      if(_zz_1953_)begin
        int_reg_array_28_2_imag <= _zz_2017_;
      end
      if(_zz_1954_)begin
        int_reg_array_28_3_imag <= _zz_2017_;
      end
      if(_zz_1955_)begin
        int_reg_array_28_4_imag <= _zz_2017_;
      end
      if(_zz_1956_)begin
        int_reg_array_28_5_imag <= _zz_2017_;
      end
      if(_zz_1957_)begin
        int_reg_array_28_6_imag <= _zz_2017_;
      end
      if(_zz_1958_)begin
        int_reg_array_28_7_imag <= _zz_2017_;
      end
      if(_zz_1959_)begin
        int_reg_array_28_8_imag <= _zz_2017_;
      end
      if(_zz_1960_)begin
        int_reg_array_28_9_imag <= _zz_2017_;
      end
      if(_zz_1961_)begin
        int_reg_array_28_10_imag <= _zz_2017_;
      end
      if(_zz_1962_)begin
        int_reg_array_28_11_imag <= _zz_2017_;
      end
      if(_zz_1963_)begin
        int_reg_array_28_12_imag <= _zz_2017_;
      end
      if(_zz_1964_)begin
        int_reg_array_28_13_imag <= _zz_2017_;
      end
      if(_zz_1965_)begin
        int_reg_array_28_14_imag <= _zz_2017_;
      end
      if(_zz_1966_)begin
        int_reg_array_28_15_imag <= _zz_2017_;
      end
      if(_zz_1967_)begin
        int_reg_array_28_16_imag <= _zz_2017_;
      end
      if(_zz_1968_)begin
        int_reg_array_28_17_imag <= _zz_2017_;
      end
      if(_zz_1969_)begin
        int_reg_array_28_18_imag <= _zz_2017_;
      end
      if(_zz_1970_)begin
        int_reg_array_28_19_imag <= _zz_2017_;
      end
      if(_zz_1971_)begin
        int_reg_array_28_20_imag <= _zz_2017_;
      end
      if(_zz_1972_)begin
        int_reg_array_28_21_imag <= _zz_2017_;
      end
      if(_zz_1973_)begin
        int_reg_array_28_22_imag <= _zz_2017_;
      end
      if(_zz_1974_)begin
        int_reg_array_28_23_imag <= _zz_2017_;
      end
      if(_zz_1975_)begin
        int_reg_array_28_24_imag <= _zz_2017_;
      end
      if(_zz_1976_)begin
        int_reg_array_28_25_imag <= _zz_2017_;
      end
      if(_zz_1977_)begin
        int_reg_array_28_26_imag <= _zz_2017_;
      end
      if(_zz_1978_)begin
        int_reg_array_28_27_imag <= _zz_2017_;
      end
      if(_zz_1979_)begin
        int_reg_array_28_28_imag <= _zz_2017_;
      end
      if(_zz_1980_)begin
        int_reg_array_28_29_imag <= _zz_2017_;
      end
      if(_zz_1981_)begin
        int_reg_array_28_30_imag <= _zz_2017_;
      end
      if(_zz_1982_)begin
        int_reg_array_28_31_imag <= _zz_2017_;
      end
      if(_zz_1983_)begin
        int_reg_array_28_32_imag <= _zz_2017_;
      end
      if(_zz_1984_)begin
        int_reg_array_28_33_imag <= _zz_2017_;
      end
      if(_zz_1985_)begin
        int_reg_array_28_34_imag <= _zz_2017_;
      end
      if(_zz_1986_)begin
        int_reg_array_28_35_imag <= _zz_2017_;
      end
      if(_zz_1987_)begin
        int_reg_array_28_36_imag <= _zz_2017_;
      end
      if(_zz_1988_)begin
        int_reg_array_28_37_imag <= _zz_2017_;
      end
      if(_zz_1989_)begin
        int_reg_array_28_38_imag <= _zz_2017_;
      end
      if(_zz_1990_)begin
        int_reg_array_28_39_imag <= _zz_2017_;
      end
      if(_zz_1991_)begin
        int_reg_array_28_40_imag <= _zz_2017_;
      end
      if(_zz_1992_)begin
        int_reg_array_28_41_imag <= _zz_2017_;
      end
      if(_zz_1993_)begin
        int_reg_array_28_42_imag <= _zz_2017_;
      end
      if(_zz_1994_)begin
        int_reg_array_28_43_imag <= _zz_2017_;
      end
      if(_zz_1995_)begin
        int_reg_array_28_44_imag <= _zz_2017_;
      end
      if(_zz_1996_)begin
        int_reg_array_28_45_imag <= _zz_2017_;
      end
      if(_zz_1997_)begin
        int_reg_array_28_46_imag <= _zz_2017_;
      end
      if(_zz_1998_)begin
        int_reg_array_28_47_imag <= _zz_2017_;
      end
      if(_zz_1999_)begin
        int_reg_array_28_48_imag <= _zz_2017_;
      end
      if(_zz_2000_)begin
        int_reg_array_28_49_imag <= _zz_2017_;
      end
      if(_zz_2001_)begin
        int_reg_array_28_50_imag <= _zz_2017_;
      end
      if(_zz_2002_)begin
        int_reg_array_28_51_imag <= _zz_2017_;
      end
      if(_zz_2003_)begin
        int_reg_array_28_52_imag <= _zz_2017_;
      end
      if(_zz_2004_)begin
        int_reg_array_28_53_imag <= _zz_2017_;
      end
      if(_zz_2005_)begin
        int_reg_array_28_54_imag <= _zz_2017_;
      end
      if(_zz_2006_)begin
        int_reg_array_28_55_imag <= _zz_2017_;
      end
      if(_zz_2007_)begin
        int_reg_array_28_56_imag <= _zz_2017_;
      end
      if(_zz_2008_)begin
        int_reg_array_28_57_imag <= _zz_2017_;
      end
      if(_zz_2009_)begin
        int_reg_array_28_58_imag <= _zz_2017_;
      end
      if(_zz_2010_)begin
        int_reg_array_28_59_imag <= _zz_2017_;
      end
      if(_zz_2011_)begin
        int_reg_array_28_60_imag <= _zz_2017_;
      end
      if(_zz_2012_)begin
        int_reg_array_28_61_imag <= _zz_2017_;
      end
      if(_zz_2013_)begin
        int_reg_array_28_62_imag <= _zz_2017_;
      end
      if(_zz_2014_)begin
        int_reg_array_28_63_imag <= _zz_2017_;
      end
      if(_zz_2020_)begin
        int_reg_array_29_0_real <= _zz_2085_;
      end
      if(_zz_2021_)begin
        int_reg_array_29_1_real <= _zz_2085_;
      end
      if(_zz_2022_)begin
        int_reg_array_29_2_real <= _zz_2085_;
      end
      if(_zz_2023_)begin
        int_reg_array_29_3_real <= _zz_2085_;
      end
      if(_zz_2024_)begin
        int_reg_array_29_4_real <= _zz_2085_;
      end
      if(_zz_2025_)begin
        int_reg_array_29_5_real <= _zz_2085_;
      end
      if(_zz_2026_)begin
        int_reg_array_29_6_real <= _zz_2085_;
      end
      if(_zz_2027_)begin
        int_reg_array_29_7_real <= _zz_2085_;
      end
      if(_zz_2028_)begin
        int_reg_array_29_8_real <= _zz_2085_;
      end
      if(_zz_2029_)begin
        int_reg_array_29_9_real <= _zz_2085_;
      end
      if(_zz_2030_)begin
        int_reg_array_29_10_real <= _zz_2085_;
      end
      if(_zz_2031_)begin
        int_reg_array_29_11_real <= _zz_2085_;
      end
      if(_zz_2032_)begin
        int_reg_array_29_12_real <= _zz_2085_;
      end
      if(_zz_2033_)begin
        int_reg_array_29_13_real <= _zz_2085_;
      end
      if(_zz_2034_)begin
        int_reg_array_29_14_real <= _zz_2085_;
      end
      if(_zz_2035_)begin
        int_reg_array_29_15_real <= _zz_2085_;
      end
      if(_zz_2036_)begin
        int_reg_array_29_16_real <= _zz_2085_;
      end
      if(_zz_2037_)begin
        int_reg_array_29_17_real <= _zz_2085_;
      end
      if(_zz_2038_)begin
        int_reg_array_29_18_real <= _zz_2085_;
      end
      if(_zz_2039_)begin
        int_reg_array_29_19_real <= _zz_2085_;
      end
      if(_zz_2040_)begin
        int_reg_array_29_20_real <= _zz_2085_;
      end
      if(_zz_2041_)begin
        int_reg_array_29_21_real <= _zz_2085_;
      end
      if(_zz_2042_)begin
        int_reg_array_29_22_real <= _zz_2085_;
      end
      if(_zz_2043_)begin
        int_reg_array_29_23_real <= _zz_2085_;
      end
      if(_zz_2044_)begin
        int_reg_array_29_24_real <= _zz_2085_;
      end
      if(_zz_2045_)begin
        int_reg_array_29_25_real <= _zz_2085_;
      end
      if(_zz_2046_)begin
        int_reg_array_29_26_real <= _zz_2085_;
      end
      if(_zz_2047_)begin
        int_reg_array_29_27_real <= _zz_2085_;
      end
      if(_zz_2048_)begin
        int_reg_array_29_28_real <= _zz_2085_;
      end
      if(_zz_2049_)begin
        int_reg_array_29_29_real <= _zz_2085_;
      end
      if(_zz_2050_)begin
        int_reg_array_29_30_real <= _zz_2085_;
      end
      if(_zz_2051_)begin
        int_reg_array_29_31_real <= _zz_2085_;
      end
      if(_zz_2052_)begin
        int_reg_array_29_32_real <= _zz_2085_;
      end
      if(_zz_2053_)begin
        int_reg_array_29_33_real <= _zz_2085_;
      end
      if(_zz_2054_)begin
        int_reg_array_29_34_real <= _zz_2085_;
      end
      if(_zz_2055_)begin
        int_reg_array_29_35_real <= _zz_2085_;
      end
      if(_zz_2056_)begin
        int_reg_array_29_36_real <= _zz_2085_;
      end
      if(_zz_2057_)begin
        int_reg_array_29_37_real <= _zz_2085_;
      end
      if(_zz_2058_)begin
        int_reg_array_29_38_real <= _zz_2085_;
      end
      if(_zz_2059_)begin
        int_reg_array_29_39_real <= _zz_2085_;
      end
      if(_zz_2060_)begin
        int_reg_array_29_40_real <= _zz_2085_;
      end
      if(_zz_2061_)begin
        int_reg_array_29_41_real <= _zz_2085_;
      end
      if(_zz_2062_)begin
        int_reg_array_29_42_real <= _zz_2085_;
      end
      if(_zz_2063_)begin
        int_reg_array_29_43_real <= _zz_2085_;
      end
      if(_zz_2064_)begin
        int_reg_array_29_44_real <= _zz_2085_;
      end
      if(_zz_2065_)begin
        int_reg_array_29_45_real <= _zz_2085_;
      end
      if(_zz_2066_)begin
        int_reg_array_29_46_real <= _zz_2085_;
      end
      if(_zz_2067_)begin
        int_reg_array_29_47_real <= _zz_2085_;
      end
      if(_zz_2068_)begin
        int_reg_array_29_48_real <= _zz_2085_;
      end
      if(_zz_2069_)begin
        int_reg_array_29_49_real <= _zz_2085_;
      end
      if(_zz_2070_)begin
        int_reg_array_29_50_real <= _zz_2085_;
      end
      if(_zz_2071_)begin
        int_reg_array_29_51_real <= _zz_2085_;
      end
      if(_zz_2072_)begin
        int_reg_array_29_52_real <= _zz_2085_;
      end
      if(_zz_2073_)begin
        int_reg_array_29_53_real <= _zz_2085_;
      end
      if(_zz_2074_)begin
        int_reg_array_29_54_real <= _zz_2085_;
      end
      if(_zz_2075_)begin
        int_reg_array_29_55_real <= _zz_2085_;
      end
      if(_zz_2076_)begin
        int_reg_array_29_56_real <= _zz_2085_;
      end
      if(_zz_2077_)begin
        int_reg_array_29_57_real <= _zz_2085_;
      end
      if(_zz_2078_)begin
        int_reg_array_29_58_real <= _zz_2085_;
      end
      if(_zz_2079_)begin
        int_reg_array_29_59_real <= _zz_2085_;
      end
      if(_zz_2080_)begin
        int_reg_array_29_60_real <= _zz_2085_;
      end
      if(_zz_2081_)begin
        int_reg_array_29_61_real <= _zz_2085_;
      end
      if(_zz_2082_)begin
        int_reg_array_29_62_real <= _zz_2085_;
      end
      if(_zz_2083_)begin
        int_reg_array_29_63_real <= _zz_2085_;
      end
      if(_zz_2020_)begin
        int_reg_array_29_0_imag <= _zz_2086_;
      end
      if(_zz_2021_)begin
        int_reg_array_29_1_imag <= _zz_2086_;
      end
      if(_zz_2022_)begin
        int_reg_array_29_2_imag <= _zz_2086_;
      end
      if(_zz_2023_)begin
        int_reg_array_29_3_imag <= _zz_2086_;
      end
      if(_zz_2024_)begin
        int_reg_array_29_4_imag <= _zz_2086_;
      end
      if(_zz_2025_)begin
        int_reg_array_29_5_imag <= _zz_2086_;
      end
      if(_zz_2026_)begin
        int_reg_array_29_6_imag <= _zz_2086_;
      end
      if(_zz_2027_)begin
        int_reg_array_29_7_imag <= _zz_2086_;
      end
      if(_zz_2028_)begin
        int_reg_array_29_8_imag <= _zz_2086_;
      end
      if(_zz_2029_)begin
        int_reg_array_29_9_imag <= _zz_2086_;
      end
      if(_zz_2030_)begin
        int_reg_array_29_10_imag <= _zz_2086_;
      end
      if(_zz_2031_)begin
        int_reg_array_29_11_imag <= _zz_2086_;
      end
      if(_zz_2032_)begin
        int_reg_array_29_12_imag <= _zz_2086_;
      end
      if(_zz_2033_)begin
        int_reg_array_29_13_imag <= _zz_2086_;
      end
      if(_zz_2034_)begin
        int_reg_array_29_14_imag <= _zz_2086_;
      end
      if(_zz_2035_)begin
        int_reg_array_29_15_imag <= _zz_2086_;
      end
      if(_zz_2036_)begin
        int_reg_array_29_16_imag <= _zz_2086_;
      end
      if(_zz_2037_)begin
        int_reg_array_29_17_imag <= _zz_2086_;
      end
      if(_zz_2038_)begin
        int_reg_array_29_18_imag <= _zz_2086_;
      end
      if(_zz_2039_)begin
        int_reg_array_29_19_imag <= _zz_2086_;
      end
      if(_zz_2040_)begin
        int_reg_array_29_20_imag <= _zz_2086_;
      end
      if(_zz_2041_)begin
        int_reg_array_29_21_imag <= _zz_2086_;
      end
      if(_zz_2042_)begin
        int_reg_array_29_22_imag <= _zz_2086_;
      end
      if(_zz_2043_)begin
        int_reg_array_29_23_imag <= _zz_2086_;
      end
      if(_zz_2044_)begin
        int_reg_array_29_24_imag <= _zz_2086_;
      end
      if(_zz_2045_)begin
        int_reg_array_29_25_imag <= _zz_2086_;
      end
      if(_zz_2046_)begin
        int_reg_array_29_26_imag <= _zz_2086_;
      end
      if(_zz_2047_)begin
        int_reg_array_29_27_imag <= _zz_2086_;
      end
      if(_zz_2048_)begin
        int_reg_array_29_28_imag <= _zz_2086_;
      end
      if(_zz_2049_)begin
        int_reg_array_29_29_imag <= _zz_2086_;
      end
      if(_zz_2050_)begin
        int_reg_array_29_30_imag <= _zz_2086_;
      end
      if(_zz_2051_)begin
        int_reg_array_29_31_imag <= _zz_2086_;
      end
      if(_zz_2052_)begin
        int_reg_array_29_32_imag <= _zz_2086_;
      end
      if(_zz_2053_)begin
        int_reg_array_29_33_imag <= _zz_2086_;
      end
      if(_zz_2054_)begin
        int_reg_array_29_34_imag <= _zz_2086_;
      end
      if(_zz_2055_)begin
        int_reg_array_29_35_imag <= _zz_2086_;
      end
      if(_zz_2056_)begin
        int_reg_array_29_36_imag <= _zz_2086_;
      end
      if(_zz_2057_)begin
        int_reg_array_29_37_imag <= _zz_2086_;
      end
      if(_zz_2058_)begin
        int_reg_array_29_38_imag <= _zz_2086_;
      end
      if(_zz_2059_)begin
        int_reg_array_29_39_imag <= _zz_2086_;
      end
      if(_zz_2060_)begin
        int_reg_array_29_40_imag <= _zz_2086_;
      end
      if(_zz_2061_)begin
        int_reg_array_29_41_imag <= _zz_2086_;
      end
      if(_zz_2062_)begin
        int_reg_array_29_42_imag <= _zz_2086_;
      end
      if(_zz_2063_)begin
        int_reg_array_29_43_imag <= _zz_2086_;
      end
      if(_zz_2064_)begin
        int_reg_array_29_44_imag <= _zz_2086_;
      end
      if(_zz_2065_)begin
        int_reg_array_29_45_imag <= _zz_2086_;
      end
      if(_zz_2066_)begin
        int_reg_array_29_46_imag <= _zz_2086_;
      end
      if(_zz_2067_)begin
        int_reg_array_29_47_imag <= _zz_2086_;
      end
      if(_zz_2068_)begin
        int_reg_array_29_48_imag <= _zz_2086_;
      end
      if(_zz_2069_)begin
        int_reg_array_29_49_imag <= _zz_2086_;
      end
      if(_zz_2070_)begin
        int_reg_array_29_50_imag <= _zz_2086_;
      end
      if(_zz_2071_)begin
        int_reg_array_29_51_imag <= _zz_2086_;
      end
      if(_zz_2072_)begin
        int_reg_array_29_52_imag <= _zz_2086_;
      end
      if(_zz_2073_)begin
        int_reg_array_29_53_imag <= _zz_2086_;
      end
      if(_zz_2074_)begin
        int_reg_array_29_54_imag <= _zz_2086_;
      end
      if(_zz_2075_)begin
        int_reg_array_29_55_imag <= _zz_2086_;
      end
      if(_zz_2076_)begin
        int_reg_array_29_56_imag <= _zz_2086_;
      end
      if(_zz_2077_)begin
        int_reg_array_29_57_imag <= _zz_2086_;
      end
      if(_zz_2078_)begin
        int_reg_array_29_58_imag <= _zz_2086_;
      end
      if(_zz_2079_)begin
        int_reg_array_29_59_imag <= _zz_2086_;
      end
      if(_zz_2080_)begin
        int_reg_array_29_60_imag <= _zz_2086_;
      end
      if(_zz_2081_)begin
        int_reg_array_29_61_imag <= _zz_2086_;
      end
      if(_zz_2082_)begin
        int_reg_array_29_62_imag <= _zz_2086_;
      end
      if(_zz_2083_)begin
        int_reg_array_29_63_imag <= _zz_2086_;
      end
      if(_zz_2089_)begin
        int_reg_array_30_0_real <= _zz_2154_;
      end
      if(_zz_2090_)begin
        int_reg_array_30_1_real <= _zz_2154_;
      end
      if(_zz_2091_)begin
        int_reg_array_30_2_real <= _zz_2154_;
      end
      if(_zz_2092_)begin
        int_reg_array_30_3_real <= _zz_2154_;
      end
      if(_zz_2093_)begin
        int_reg_array_30_4_real <= _zz_2154_;
      end
      if(_zz_2094_)begin
        int_reg_array_30_5_real <= _zz_2154_;
      end
      if(_zz_2095_)begin
        int_reg_array_30_6_real <= _zz_2154_;
      end
      if(_zz_2096_)begin
        int_reg_array_30_7_real <= _zz_2154_;
      end
      if(_zz_2097_)begin
        int_reg_array_30_8_real <= _zz_2154_;
      end
      if(_zz_2098_)begin
        int_reg_array_30_9_real <= _zz_2154_;
      end
      if(_zz_2099_)begin
        int_reg_array_30_10_real <= _zz_2154_;
      end
      if(_zz_2100_)begin
        int_reg_array_30_11_real <= _zz_2154_;
      end
      if(_zz_2101_)begin
        int_reg_array_30_12_real <= _zz_2154_;
      end
      if(_zz_2102_)begin
        int_reg_array_30_13_real <= _zz_2154_;
      end
      if(_zz_2103_)begin
        int_reg_array_30_14_real <= _zz_2154_;
      end
      if(_zz_2104_)begin
        int_reg_array_30_15_real <= _zz_2154_;
      end
      if(_zz_2105_)begin
        int_reg_array_30_16_real <= _zz_2154_;
      end
      if(_zz_2106_)begin
        int_reg_array_30_17_real <= _zz_2154_;
      end
      if(_zz_2107_)begin
        int_reg_array_30_18_real <= _zz_2154_;
      end
      if(_zz_2108_)begin
        int_reg_array_30_19_real <= _zz_2154_;
      end
      if(_zz_2109_)begin
        int_reg_array_30_20_real <= _zz_2154_;
      end
      if(_zz_2110_)begin
        int_reg_array_30_21_real <= _zz_2154_;
      end
      if(_zz_2111_)begin
        int_reg_array_30_22_real <= _zz_2154_;
      end
      if(_zz_2112_)begin
        int_reg_array_30_23_real <= _zz_2154_;
      end
      if(_zz_2113_)begin
        int_reg_array_30_24_real <= _zz_2154_;
      end
      if(_zz_2114_)begin
        int_reg_array_30_25_real <= _zz_2154_;
      end
      if(_zz_2115_)begin
        int_reg_array_30_26_real <= _zz_2154_;
      end
      if(_zz_2116_)begin
        int_reg_array_30_27_real <= _zz_2154_;
      end
      if(_zz_2117_)begin
        int_reg_array_30_28_real <= _zz_2154_;
      end
      if(_zz_2118_)begin
        int_reg_array_30_29_real <= _zz_2154_;
      end
      if(_zz_2119_)begin
        int_reg_array_30_30_real <= _zz_2154_;
      end
      if(_zz_2120_)begin
        int_reg_array_30_31_real <= _zz_2154_;
      end
      if(_zz_2121_)begin
        int_reg_array_30_32_real <= _zz_2154_;
      end
      if(_zz_2122_)begin
        int_reg_array_30_33_real <= _zz_2154_;
      end
      if(_zz_2123_)begin
        int_reg_array_30_34_real <= _zz_2154_;
      end
      if(_zz_2124_)begin
        int_reg_array_30_35_real <= _zz_2154_;
      end
      if(_zz_2125_)begin
        int_reg_array_30_36_real <= _zz_2154_;
      end
      if(_zz_2126_)begin
        int_reg_array_30_37_real <= _zz_2154_;
      end
      if(_zz_2127_)begin
        int_reg_array_30_38_real <= _zz_2154_;
      end
      if(_zz_2128_)begin
        int_reg_array_30_39_real <= _zz_2154_;
      end
      if(_zz_2129_)begin
        int_reg_array_30_40_real <= _zz_2154_;
      end
      if(_zz_2130_)begin
        int_reg_array_30_41_real <= _zz_2154_;
      end
      if(_zz_2131_)begin
        int_reg_array_30_42_real <= _zz_2154_;
      end
      if(_zz_2132_)begin
        int_reg_array_30_43_real <= _zz_2154_;
      end
      if(_zz_2133_)begin
        int_reg_array_30_44_real <= _zz_2154_;
      end
      if(_zz_2134_)begin
        int_reg_array_30_45_real <= _zz_2154_;
      end
      if(_zz_2135_)begin
        int_reg_array_30_46_real <= _zz_2154_;
      end
      if(_zz_2136_)begin
        int_reg_array_30_47_real <= _zz_2154_;
      end
      if(_zz_2137_)begin
        int_reg_array_30_48_real <= _zz_2154_;
      end
      if(_zz_2138_)begin
        int_reg_array_30_49_real <= _zz_2154_;
      end
      if(_zz_2139_)begin
        int_reg_array_30_50_real <= _zz_2154_;
      end
      if(_zz_2140_)begin
        int_reg_array_30_51_real <= _zz_2154_;
      end
      if(_zz_2141_)begin
        int_reg_array_30_52_real <= _zz_2154_;
      end
      if(_zz_2142_)begin
        int_reg_array_30_53_real <= _zz_2154_;
      end
      if(_zz_2143_)begin
        int_reg_array_30_54_real <= _zz_2154_;
      end
      if(_zz_2144_)begin
        int_reg_array_30_55_real <= _zz_2154_;
      end
      if(_zz_2145_)begin
        int_reg_array_30_56_real <= _zz_2154_;
      end
      if(_zz_2146_)begin
        int_reg_array_30_57_real <= _zz_2154_;
      end
      if(_zz_2147_)begin
        int_reg_array_30_58_real <= _zz_2154_;
      end
      if(_zz_2148_)begin
        int_reg_array_30_59_real <= _zz_2154_;
      end
      if(_zz_2149_)begin
        int_reg_array_30_60_real <= _zz_2154_;
      end
      if(_zz_2150_)begin
        int_reg_array_30_61_real <= _zz_2154_;
      end
      if(_zz_2151_)begin
        int_reg_array_30_62_real <= _zz_2154_;
      end
      if(_zz_2152_)begin
        int_reg_array_30_63_real <= _zz_2154_;
      end
      if(_zz_2089_)begin
        int_reg_array_30_0_imag <= _zz_2155_;
      end
      if(_zz_2090_)begin
        int_reg_array_30_1_imag <= _zz_2155_;
      end
      if(_zz_2091_)begin
        int_reg_array_30_2_imag <= _zz_2155_;
      end
      if(_zz_2092_)begin
        int_reg_array_30_3_imag <= _zz_2155_;
      end
      if(_zz_2093_)begin
        int_reg_array_30_4_imag <= _zz_2155_;
      end
      if(_zz_2094_)begin
        int_reg_array_30_5_imag <= _zz_2155_;
      end
      if(_zz_2095_)begin
        int_reg_array_30_6_imag <= _zz_2155_;
      end
      if(_zz_2096_)begin
        int_reg_array_30_7_imag <= _zz_2155_;
      end
      if(_zz_2097_)begin
        int_reg_array_30_8_imag <= _zz_2155_;
      end
      if(_zz_2098_)begin
        int_reg_array_30_9_imag <= _zz_2155_;
      end
      if(_zz_2099_)begin
        int_reg_array_30_10_imag <= _zz_2155_;
      end
      if(_zz_2100_)begin
        int_reg_array_30_11_imag <= _zz_2155_;
      end
      if(_zz_2101_)begin
        int_reg_array_30_12_imag <= _zz_2155_;
      end
      if(_zz_2102_)begin
        int_reg_array_30_13_imag <= _zz_2155_;
      end
      if(_zz_2103_)begin
        int_reg_array_30_14_imag <= _zz_2155_;
      end
      if(_zz_2104_)begin
        int_reg_array_30_15_imag <= _zz_2155_;
      end
      if(_zz_2105_)begin
        int_reg_array_30_16_imag <= _zz_2155_;
      end
      if(_zz_2106_)begin
        int_reg_array_30_17_imag <= _zz_2155_;
      end
      if(_zz_2107_)begin
        int_reg_array_30_18_imag <= _zz_2155_;
      end
      if(_zz_2108_)begin
        int_reg_array_30_19_imag <= _zz_2155_;
      end
      if(_zz_2109_)begin
        int_reg_array_30_20_imag <= _zz_2155_;
      end
      if(_zz_2110_)begin
        int_reg_array_30_21_imag <= _zz_2155_;
      end
      if(_zz_2111_)begin
        int_reg_array_30_22_imag <= _zz_2155_;
      end
      if(_zz_2112_)begin
        int_reg_array_30_23_imag <= _zz_2155_;
      end
      if(_zz_2113_)begin
        int_reg_array_30_24_imag <= _zz_2155_;
      end
      if(_zz_2114_)begin
        int_reg_array_30_25_imag <= _zz_2155_;
      end
      if(_zz_2115_)begin
        int_reg_array_30_26_imag <= _zz_2155_;
      end
      if(_zz_2116_)begin
        int_reg_array_30_27_imag <= _zz_2155_;
      end
      if(_zz_2117_)begin
        int_reg_array_30_28_imag <= _zz_2155_;
      end
      if(_zz_2118_)begin
        int_reg_array_30_29_imag <= _zz_2155_;
      end
      if(_zz_2119_)begin
        int_reg_array_30_30_imag <= _zz_2155_;
      end
      if(_zz_2120_)begin
        int_reg_array_30_31_imag <= _zz_2155_;
      end
      if(_zz_2121_)begin
        int_reg_array_30_32_imag <= _zz_2155_;
      end
      if(_zz_2122_)begin
        int_reg_array_30_33_imag <= _zz_2155_;
      end
      if(_zz_2123_)begin
        int_reg_array_30_34_imag <= _zz_2155_;
      end
      if(_zz_2124_)begin
        int_reg_array_30_35_imag <= _zz_2155_;
      end
      if(_zz_2125_)begin
        int_reg_array_30_36_imag <= _zz_2155_;
      end
      if(_zz_2126_)begin
        int_reg_array_30_37_imag <= _zz_2155_;
      end
      if(_zz_2127_)begin
        int_reg_array_30_38_imag <= _zz_2155_;
      end
      if(_zz_2128_)begin
        int_reg_array_30_39_imag <= _zz_2155_;
      end
      if(_zz_2129_)begin
        int_reg_array_30_40_imag <= _zz_2155_;
      end
      if(_zz_2130_)begin
        int_reg_array_30_41_imag <= _zz_2155_;
      end
      if(_zz_2131_)begin
        int_reg_array_30_42_imag <= _zz_2155_;
      end
      if(_zz_2132_)begin
        int_reg_array_30_43_imag <= _zz_2155_;
      end
      if(_zz_2133_)begin
        int_reg_array_30_44_imag <= _zz_2155_;
      end
      if(_zz_2134_)begin
        int_reg_array_30_45_imag <= _zz_2155_;
      end
      if(_zz_2135_)begin
        int_reg_array_30_46_imag <= _zz_2155_;
      end
      if(_zz_2136_)begin
        int_reg_array_30_47_imag <= _zz_2155_;
      end
      if(_zz_2137_)begin
        int_reg_array_30_48_imag <= _zz_2155_;
      end
      if(_zz_2138_)begin
        int_reg_array_30_49_imag <= _zz_2155_;
      end
      if(_zz_2139_)begin
        int_reg_array_30_50_imag <= _zz_2155_;
      end
      if(_zz_2140_)begin
        int_reg_array_30_51_imag <= _zz_2155_;
      end
      if(_zz_2141_)begin
        int_reg_array_30_52_imag <= _zz_2155_;
      end
      if(_zz_2142_)begin
        int_reg_array_30_53_imag <= _zz_2155_;
      end
      if(_zz_2143_)begin
        int_reg_array_30_54_imag <= _zz_2155_;
      end
      if(_zz_2144_)begin
        int_reg_array_30_55_imag <= _zz_2155_;
      end
      if(_zz_2145_)begin
        int_reg_array_30_56_imag <= _zz_2155_;
      end
      if(_zz_2146_)begin
        int_reg_array_30_57_imag <= _zz_2155_;
      end
      if(_zz_2147_)begin
        int_reg_array_30_58_imag <= _zz_2155_;
      end
      if(_zz_2148_)begin
        int_reg_array_30_59_imag <= _zz_2155_;
      end
      if(_zz_2149_)begin
        int_reg_array_30_60_imag <= _zz_2155_;
      end
      if(_zz_2150_)begin
        int_reg_array_30_61_imag <= _zz_2155_;
      end
      if(_zz_2151_)begin
        int_reg_array_30_62_imag <= _zz_2155_;
      end
      if(_zz_2152_)begin
        int_reg_array_30_63_imag <= _zz_2155_;
      end
      if(_zz_2158_)begin
        int_reg_array_31_0_real <= _zz_2223_;
      end
      if(_zz_2159_)begin
        int_reg_array_31_1_real <= _zz_2223_;
      end
      if(_zz_2160_)begin
        int_reg_array_31_2_real <= _zz_2223_;
      end
      if(_zz_2161_)begin
        int_reg_array_31_3_real <= _zz_2223_;
      end
      if(_zz_2162_)begin
        int_reg_array_31_4_real <= _zz_2223_;
      end
      if(_zz_2163_)begin
        int_reg_array_31_5_real <= _zz_2223_;
      end
      if(_zz_2164_)begin
        int_reg_array_31_6_real <= _zz_2223_;
      end
      if(_zz_2165_)begin
        int_reg_array_31_7_real <= _zz_2223_;
      end
      if(_zz_2166_)begin
        int_reg_array_31_8_real <= _zz_2223_;
      end
      if(_zz_2167_)begin
        int_reg_array_31_9_real <= _zz_2223_;
      end
      if(_zz_2168_)begin
        int_reg_array_31_10_real <= _zz_2223_;
      end
      if(_zz_2169_)begin
        int_reg_array_31_11_real <= _zz_2223_;
      end
      if(_zz_2170_)begin
        int_reg_array_31_12_real <= _zz_2223_;
      end
      if(_zz_2171_)begin
        int_reg_array_31_13_real <= _zz_2223_;
      end
      if(_zz_2172_)begin
        int_reg_array_31_14_real <= _zz_2223_;
      end
      if(_zz_2173_)begin
        int_reg_array_31_15_real <= _zz_2223_;
      end
      if(_zz_2174_)begin
        int_reg_array_31_16_real <= _zz_2223_;
      end
      if(_zz_2175_)begin
        int_reg_array_31_17_real <= _zz_2223_;
      end
      if(_zz_2176_)begin
        int_reg_array_31_18_real <= _zz_2223_;
      end
      if(_zz_2177_)begin
        int_reg_array_31_19_real <= _zz_2223_;
      end
      if(_zz_2178_)begin
        int_reg_array_31_20_real <= _zz_2223_;
      end
      if(_zz_2179_)begin
        int_reg_array_31_21_real <= _zz_2223_;
      end
      if(_zz_2180_)begin
        int_reg_array_31_22_real <= _zz_2223_;
      end
      if(_zz_2181_)begin
        int_reg_array_31_23_real <= _zz_2223_;
      end
      if(_zz_2182_)begin
        int_reg_array_31_24_real <= _zz_2223_;
      end
      if(_zz_2183_)begin
        int_reg_array_31_25_real <= _zz_2223_;
      end
      if(_zz_2184_)begin
        int_reg_array_31_26_real <= _zz_2223_;
      end
      if(_zz_2185_)begin
        int_reg_array_31_27_real <= _zz_2223_;
      end
      if(_zz_2186_)begin
        int_reg_array_31_28_real <= _zz_2223_;
      end
      if(_zz_2187_)begin
        int_reg_array_31_29_real <= _zz_2223_;
      end
      if(_zz_2188_)begin
        int_reg_array_31_30_real <= _zz_2223_;
      end
      if(_zz_2189_)begin
        int_reg_array_31_31_real <= _zz_2223_;
      end
      if(_zz_2190_)begin
        int_reg_array_31_32_real <= _zz_2223_;
      end
      if(_zz_2191_)begin
        int_reg_array_31_33_real <= _zz_2223_;
      end
      if(_zz_2192_)begin
        int_reg_array_31_34_real <= _zz_2223_;
      end
      if(_zz_2193_)begin
        int_reg_array_31_35_real <= _zz_2223_;
      end
      if(_zz_2194_)begin
        int_reg_array_31_36_real <= _zz_2223_;
      end
      if(_zz_2195_)begin
        int_reg_array_31_37_real <= _zz_2223_;
      end
      if(_zz_2196_)begin
        int_reg_array_31_38_real <= _zz_2223_;
      end
      if(_zz_2197_)begin
        int_reg_array_31_39_real <= _zz_2223_;
      end
      if(_zz_2198_)begin
        int_reg_array_31_40_real <= _zz_2223_;
      end
      if(_zz_2199_)begin
        int_reg_array_31_41_real <= _zz_2223_;
      end
      if(_zz_2200_)begin
        int_reg_array_31_42_real <= _zz_2223_;
      end
      if(_zz_2201_)begin
        int_reg_array_31_43_real <= _zz_2223_;
      end
      if(_zz_2202_)begin
        int_reg_array_31_44_real <= _zz_2223_;
      end
      if(_zz_2203_)begin
        int_reg_array_31_45_real <= _zz_2223_;
      end
      if(_zz_2204_)begin
        int_reg_array_31_46_real <= _zz_2223_;
      end
      if(_zz_2205_)begin
        int_reg_array_31_47_real <= _zz_2223_;
      end
      if(_zz_2206_)begin
        int_reg_array_31_48_real <= _zz_2223_;
      end
      if(_zz_2207_)begin
        int_reg_array_31_49_real <= _zz_2223_;
      end
      if(_zz_2208_)begin
        int_reg_array_31_50_real <= _zz_2223_;
      end
      if(_zz_2209_)begin
        int_reg_array_31_51_real <= _zz_2223_;
      end
      if(_zz_2210_)begin
        int_reg_array_31_52_real <= _zz_2223_;
      end
      if(_zz_2211_)begin
        int_reg_array_31_53_real <= _zz_2223_;
      end
      if(_zz_2212_)begin
        int_reg_array_31_54_real <= _zz_2223_;
      end
      if(_zz_2213_)begin
        int_reg_array_31_55_real <= _zz_2223_;
      end
      if(_zz_2214_)begin
        int_reg_array_31_56_real <= _zz_2223_;
      end
      if(_zz_2215_)begin
        int_reg_array_31_57_real <= _zz_2223_;
      end
      if(_zz_2216_)begin
        int_reg_array_31_58_real <= _zz_2223_;
      end
      if(_zz_2217_)begin
        int_reg_array_31_59_real <= _zz_2223_;
      end
      if(_zz_2218_)begin
        int_reg_array_31_60_real <= _zz_2223_;
      end
      if(_zz_2219_)begin
        int_reg_array_31_61_real <= _zz_2223_;
      end
      if(_zz_2220_)begin
        int_reg_array_31_62_real <= _zz_2223_;
      end
      if(_zz_2221_)begin
        int_reg_array_31_63_real <= _zz_2223_;
      end
      if(_zz_2158_)begin
        int_reg_array_31_0_imag <= _zz_2224_;
      end
      if(_zz_2159_)begin
        int_reg_array_31_1_imag <= _zz_2224_;
      end
      if(_zz_2160_)begin
        int_reg_array_31_2_imag <= _zz_2224_;
      end
      if(_zz_2161_)begin
        int_reg_array_31_3_imag <= _zz_2224_;
      end
      if(_zz_2162_)begin
        int_reg_array_31_4_imag <= _zz_2224_;
      end
      if(_zz_2163_)begin
        int_reg_array_31_5_imag <= _zz_2224_;
      end
      if(_zz_2164_)begin
        int_reg_array_31_6_imag <= _zz_2224_;
      end
      if(_zz_2165_)begin
        int_reg_array_31_7_imag <= _zz_2224_;
      end
      if(_zz_2166_)begin
        int_reg_array_31_8_imag <= _zz_2224_;
      end
      if(_zz_2167_)begin
        int_reg_array_31_9_imag <= _zz_2224_;
      end
      if(_zz_2168_)begin
        int_reg_array_31_10_imag <= _zz_2224_;
      end
      if(_zz_2169_)begin
        int_reg_array_31_11_imag <= _zz_2224_;
      end
      if(_zz_2170_)begin
        int_reg_array_31_12_imag <= _zz_2224_;
      end
      if(_zz_2171_)begin
        int_reg_array_31_13_imag <= _zz_2224_;
      end
      if(_zz_2172_)begin
        int_reg_array_31_14_imag <= _zz_2224_;
      end
      if(_zz_2173_)begin
        int_reg_array_31_15_imag <= _zz_2224_;
      end
      if(_zz_2174_)begin
        int_reg_array_31_16_imag <= _zz_2224_;
      end
      if(_zz_2175_)begin
        int_reg_array_31_17_imag <= _zz_2224_;
      end
      if(_zz_2176_)begin
        int_reg_array_31_18_imag <= _zz_2224_;
      end
      if(_zz_2177_)begin
        int_reg_array_31_19_imag <= _zz_2224_;
      end
      if(_zz_2178_)begin
        int_reg_array_31_20_imag <= _zz_2224_;
      end
      if(_zz_2179_)begin
        int_reg_array_31_21_imag <= _zz_2224_;
      end
      if(_zz_2180_)begin
        int_reg_array_31_22_imag <= _zz_2224_;
      end
      if(_zz_2181_)begin
        int_reg_array_31_23_imag <= _zz_2224_;
      end
      if(_zz_2182_)begin
        int_reg_array_31_24_imag <= _zz_2224_;
      end
      if(_zz_2183_)begin
        int_reg_array_31_25_imag <= _zz_2224_;
      end
      if(_zz_2184_)begin
        int_reg_array_31_26_imag <= _zz_2224_;
      end
      if(_zz_2185_)begin
        int_reg_array_31_27_imag <= _zz_2224_;
      end
      if(_zz_2186_)begin
        int_reg_array_31_28_imag <= _zz_2224_;
      end
      if(_zz_2187_)begin
        int_reg_array_31_29_imag <= _zz_2224_;
      end
      if(_zz_2188_)begin
        int_reg_array_31_30_imag <= _zz_2224_;
      end
      if(_zz_2189_)begin
        int_reg_array_31_31_imag <= _zz_2224_;
      end
      if(_zz_2190_)begin
        int_reg_array_31_32_imag <= _zz_2224_;
      end
      if(_zz_2191_)begin
        int_reg_array_31_33_imag <= _zz_2224_;
      end
      if(_zz_2192_)begin
        int_reg_array_31_34_imag <= _zz_2224_;
      end
      if(_zz_2193_)begin
        int_reg_array_31_35_imag <= _zz_2224_;
      end
      if(_zz_2194_)begin
        int_reg_array_31_36_imag <= _zz_2224_;
      end
      if(_zz_2195_)begin
        int_reg_array_31_37_imag <= _zz_2224_;
      end
      if(_zz_2196_)begin
        int_reg_array_31_38_imag <= _zz_2224_;
      end
      if(_zz_2197_)begin
        int_reg_array_31_39_imag <= _zz_2224_;
      end
      if(_zz_2198_)begin
        int_reg_array_31_40_imag <= _zz_2224_;
      end
      if(_zz_2199_)begin
        int_reg_array_31_41_imag <= _zz_2224_;
      end
      if(_zz_2200_)begin
        int_reg_array_31_42_imag <= _zz_2224_;
      end
      if(_zz_2201_)begin
        int_reg_array_31_43_imag <= _zz_2224_;
      end
      if(_zz_2202_)begin
        int_reg_array_31_44_imag <= _zz_2224_;
      end
      if(_zz_2203_)begin
        int_reg_array_31_45_imag <= _zz_2224_;
      end
      if(_zz_2204_)begin
        int_reg_array_31_46_imag <= _zz_2224_;
      end
      if(_zz_2205_)begin
        int_reg_array_31_47_imag <= _zz_2224_;
      end
      if(_zz_2206_)begin
        int_reg_array_31_48_imag <= _zz_2224_;
      end
      if(_zz_2207_)begin
        int_reg_array_31_49_imag <= _zz_2224_;
      end
      if(_zz_2208_)begin
        int_reg_array_31_50_imag <= _zz_2224_;
      end
      if(_zz_2209_)begin
        int_reg_array_31_51_imag <= _zz_2224_;
      end
      if(_zz_2210_)begin
        int_reg_array_31_52_imag <= _zz_2224_;
      end
      if(_zz_2211_)begin
        int_reg_array_31_53_imag <= _zz_2224_;
      end
      if(_zz_2212_)begin
        int_reg_array_31_54_imag <= _zz_2224_;
      end
      if(_zz_2213_)begin
        int_reg_array_31_55_imag <= _zz_2224_;
      end
      if(_zz_2214_)begin
        int_reg_array_31_56_imag <= _zz_2224_;
      end
      if(_zz_2215_)begin
        int_reg_array_31_57_imag <= _zz_2224_;
      end
      if(_zz_2216_)begin
        int_reg_array_31_58_imag <= _zz_2224_;
      end
      if(_zz_2217_)begin
        int_reg_array_31_59_imag <= _zz_2224_;
      end
      if(_zz_2218_)begin
        int_reg_array_31_60_imag <= _zz_2224_;
      end
      if(_zz_2219_)begin
        int_reg_array_31_61_imag <= _zz_2224_;
      end
      if(_zz_2220_)begin
        int_reg_array_31_62_imag <= _zz_2224_;
      end
      if(_zz_2221_)begin
        int_reg_array_31_63_imag <= _zz_2224_;
      end
      if(_zz_2227_)begin
        int_reg_array_32_0_real <= _zz_2292_;
      end
      if(_zz_2228_)begin
        int_reg_array_32_1_real <= _zz_2292_;
      end
      if(_zz_2229_)begin
        int_reg_array_32_2_real <= _zz_2292_;
      end
      if(_zz_2230_)begin
        int_reg_array_32_3_real <= _zz_2292_;
      end
      if(_zz_2231_)begin
        int_reg_array_32_4_real <= _zz_2292_;
      end
      if(_zz_2232_)begin
        int_reg_array_32_5_real <= _zz_2292_;
      end
      if(_zz_2233_)begin
        int_reg_array_32_6_real <= _zz_2292_;
      end
      if(_zz_2234_)begin
        int_reg_array_32_7_real <= _zz_2292_;
      end
      if(_zz_2235_)begin
        int_reg_array_32_8_real <= _zz_2292_;
      end
      if(_zz_2236_)begin
        int_reg_array_32_9_real <= _zz_2292_;
      end
      if(_zz_2237_)begin
        int_reg_array_32_10_real <= _zz_2292_;
      end
      if(_zz_2238_)begin
        int_reg_array_32_11_real <= _zz_2292_;
      end
      if(_zz_2239_)begin
        int_reg_array_32_12_real <= _zz_2292_;
      end
      if(_zz_2240_)begin
        int_reg_array_32_13_real <= _zz_2292_;
      end
      if(_zz_2241_)begin
        int_reg_array_32_14_real <= _zz_2292_;
      end
      if(_zz_2242_)begin
        int_reg_array_32_15_real <= _zz_2292_;
      end
      if(_zz_2243_)begin
        int_reg_array_32_16_real <= _zz_2292_;
      end
      if(_zz_2244_)begin
        int_reg_array_32_17_real <= _zz_2292_;
      end
      if(_zz_2245_)begin
        int_reg_array_32_18_real <= _zz_2292_;
      end
      if(_zz_2246_)begin
        int_reg_array_32_19_real <= _zz_2292_;
      end
      if(_zz_2247_)begin
        int_reg_array_32_20_real <= _zz_2292_;
      end
      if(_zz_2248_)begin
        int_reg_array_32_21_real <= _zz_2292_;
      end
      if(_zz_2249_)begin
        int_reg_array_32_22_real <= _zz_2292_;
      end
      if(_zz_2250_)begin
        int_reg_array_32_23_real <= _zz_2292_;
      end
      if(_zz_2251_)begin
        int_reg_array_32_24_real <= _zz_2292_;
      end
      if(_zz_2252_)begin
        int_reg_array_32_25_real <= _zz_2292_;
      end
      if(_zz_2253_)begin
        int_reg_array_32_26_real <= _zz_2292_;
      end
      if(_zz_2254_)begin
        int_reg_array_32_27_real <= _zz_2292_;
      end
      if(_zz_2255_)begin
        int_reg_array_32_28_real <= _zz_2292_;
      end
      if(_zz_2256_)begin
        int_reg_array_32_29_real <= _zz_2292_;
      end
      if(_zz_2257_)begin
        int_reg_array_32_30_real <= _zz_2292_;
      end
      if(_zz_2258_)begin
        int_reg_array_32_31_real <= _zz_2292_;
      end
      if(_zz_2259_)begin
        int_reg_array_32_32_real <= _zz_2292_;
      end
      if(_zz_2260_)begin
        int_reg_array_32_33_real <= _zz_2292_;
      end
      if(_zz_2261_)begin
        int_reg_array_32_34_real <= _zz_2292_;
      end
      if(_zz_2262_)begin
        int_reg_array_32_35_real <= _zz_2292_;
      end
      if(_zz_2263_)begin
        int_reg_array_32_36_real <= _zz_2292_;
      end
      if(_zz_2264_)begin
        int_reg_array_32_37_real <= _zz_2292_;
      end
      if(_zz_2265_)begin
        int_reg_array_32_38_real <= _zz_2292_;
      end
      if(_zz_2266_)begin
        int_reg_array_32_39_real <= _zz_2292_;
      end
      if(_zz_2267_)begin
        int_reg_array_32_40_real <= _zz_2292_;
      end
      if(_zz_2268_)begin
        int_reg_array_32_41_real <= _zz_2292_;
      end
      if(_zz_2269_)begin
        int_reg_array_32_42_real <= _zz_2292_;
      end
      if(_zz_2270_)begin
        int_reg_array_32_43_real <= _zz_2292_;
      end
      if(_zz_2271_)begin
        int_reg_array_32_44_real <= _zz_2292_;
      end
      if(_zz_2272_)begin
        int_reg_array_32_45_real <= _zz_2292_;
      end
      if(_zz_2273_)begin
        int_reg_array_32_46_real <= _zz_2292_;
      end
      if(_zz_2274_)begin
        int_reg_array_32_47_real <= _zz_2292_;
      end
      if(_zz_2275_)begin
        int_reg_array_32_48_real <= _zz_2292_;
      end
      if(_zz_2276_)begin
        int_reg_array_32_49_real <= _zz_2292_;
      end
      if(_zz_2277_)begin
        int_reg_array_32_50_real <= _zz_2292_;
      end
      if(_zz_2278_)begin
        int_reg_array_32_51_real <= _zz_2292_;
      end
      if(_zz_2279_)begin
        int_reg_array_32_52_real <= _zz_2292_;
      end
      if(_zz_2280_)begin
        int_reg_array_32_53_real <= _zz_2292_;
      end
      if(_zz_2281_)begin
        int_reg_array_32_54_real <= _zz_2292_;
      end
      if(_zz_2282_)begin
        int_reg_array_32_55_real <= _zz_2292_;
      end
      if(_zz_2283_)begin
        int_reg_array_32_56_real <= _zz_2292_;
      end
      if(_zz_2284_)begin
        int_reg_array_32_57_real <= _zz_2292_;
      end
      if(_zz_2285_)begin
        int_reg_array_32_58_real <= _zz_2292_;
      end
      if(_zz_2286_)begin
        int_reg_array_32_59_real <= _zz_2292_;
      end
      if(_zz_2287_)begin
        int_reg_array_32_60_real <= _zz_2292_;
      end
      if(_zz_2288_)begin
        int_reg_array_32_61_real <= _zz_2292_;
      end
      if(_zz_2289_)begin
        int_reg_array_32_62_real <= _zz_2292_;
      end
      if(_zz_2290_)begin
        int_reg_array_32_63_real <= _zz_2292_;
      end
      if(_zz_2227_)begin
        int_reg_array_32_0_imag <= _zz_2293_;
      end
      if(_zz_2228_)begin
        int_reg_array_32_1_imag <= _zz_2293_;
      end
      if(_zz_2229_)begin
        int_reg_array_32_2_imag <= _zz_2293_;
      end
      if(_zz_2230_)begin
        int_reg_array_32_3_imag <= _zz_2293_;
      end
      if(_zz_2231_)begin
        int_reg_array_32_4_imag <= _zz_2293_;
      end
      if(_zz_2232_)begin
        int_reg_array_32_5_imag <= _zz_2293_;
      end
      if(_zz_2233_)begin
        int_reg_array_32_6_imag <= _zz_2293_;
      end
      if(_zz_2234_)begin
        int_reg_array_32_7_imag <= _zz_2293_;
      end
      if(_zz_2235_)begin
        int_reg_array_32_8_imag <= _zz_2293_;
      end
      if(_zz_2236_)begin
        int_reg_array_32_9_imag <= _zz_2293_;
      end
      if(_zz_2237_)begin
        int_reg_array_32_10_imag <= _zz_2293_;
      end
      if(_zz_2238_)begin
        int_reg_array_32_11_imag <= _zz_2293_;
      end
      if(_zz_2239_)begin
        int_reg_array_32_12_imag <= _zz_2293_;
      end
      if(_zz_2240_)begin
        int_reg_array_32_13_imag <= _zz_2293_;
      end
      if(_zz_2241_)begin
        int_reg_array_32_14_imag <= _zz_2293_;
      end
      if(_zz_2242_)begin
        int_reg_array_32_15_imag <= _zz_2293_;
      end
      if(_zz_2243_)begin
        int_reg_array_32_16_imag <= _zz_2293_;
      end
      if(_zz_2244_)begin
        int_reg_array_32_17_imag <= _zz_2293_;
      end
      if(_zz_2245_)begin
        int_reg_array_32_18_imag <= _zz_2293_;
      end
      if(_zz_2246_)begin
        int_reg_array_32_19_imag <= _zz_2293_;
      end
      if(_zz_2247_)begin
        int_reg_array_32_20_imag <= _zz_2293_;
      end
      if(_zz_2248_)begin
        int_reg_array_32_21_imag <= _zz_2293_;
      end
      if(_zz_2249_)begin
        int_reg_array_32_22_imag <= _zz_2293_;
      end
      if(_zz_2250_)begin
        int_reg_array_32_23_imag <= _zz_2293_;
      end
      if(_zz_2251_)begin
        int_reg_array_32_24_imag <= _zz_2293_;
      end
      if(_zz_2252_)begin
        int_reg_array_32_25_imag <= _zz_2293_;
      end
      if(_zz_2253_)begin
        int_reg_array_32_26_imag <= _zz_2293_;
      end
      if(_zz_2254_)begin
        int_reg_array_32_27_imag <= _zz_2293_;
      end
      if(_zz_2255_)begin
        int_reg_array_32_28_imag <= _zz_2293_;
      end
      if(_zz_2256_)begin
        int_reg_array_32_29_imag <= _zz_2293_;
      end
      if(_zz_2257_)begin
        int_reg_array_32_30_imag <= _zz_2293_;
      end
      if(_zz_2258_)begin
        int_reg_array_32_31_imag <= _zz_2293_;
      end
      if(_zz_2259_)begin
        int_reg_array_32_32_imag <= _zz_2293_;
      end
      if(_zz_2260_)begin
        int_reg_array_32_33_imag <= _zz_2293_;
      end
      if(_zz_2261_)begin
        int_reg_array_32_34_imag <= _zz_2293_;
      end
      if(_zz_2262_)begin
        int_reg_array_32_35_imag <= _zz_2293_;
      end
      if(_zz_2263_)begin
        int_reg_array_32_36_imag <= _zz_2293_;
      end
      if(_zz_2264_)begin
        int_reg_array_32_37_imag <= _zz_2293_;
      end
      if(_zz_2265_)begin
        int_reg_array_32_38_imag <= _zz_2293_;
      end
      if(_zz_2266_)begin
        int_reg_array_32_39_imag <= _zz_2293_;
      end
      if(_zz_2267_)begin
        int_reg_array_32_40_imag <= _zz_2293_;
      end
      if(_zz_2268_)begin
        int_reg_array_32_41_imag <= _zz_2293_;
      end
      if(_zz_2269_)begin
        int_reg_array_32_42_imag <= _zz_2293_;
      end
      if(_zz_2270_)begin
        int_reg_array_32_43_imag <= _zz_2293_;
      end
      if(_zz_2271_)begin
        int_reg_array_32_44_imag <= _zz_2293_;
      end
      if(_zz_2272_)begin
        int_reg_array_32_45_imag <= _zz_2293_;
      end
      if(_zz_2273_)begin
        int_reg_array_32_46_imag <= _zz_2293_;
      end
      if(_zz_2274_)begin
        int_reg_array_32_47_imag <= _zz_2293_;
      end
      if(_zz_2275_)begin
        int_reg_array_32_48_imag <= _zz_2293_;
      end
      if(_zz_2276_)begin
        int_reg_array_32_49_imag <= _zz_2293_;
      end
      if(_zz_2277_)begin
        int_reg_array_32_50_imag <= _zz_2293_;
      end
      if(_zz_2278_)begin
        int_reg_array_32_51_imag <= _zz_2293_;
      end
      if(_zz_2279_)begin
        int_reg_array_32_52_imag <= _zz_2293_;
      end
      if(_zz_2280_)begin
        int_reg_array_32_53_imag <= _zz_2293_;
      end
      if(_zz_2281_)begin
        int_reg_array_32_54_imag <= _zz_2293_;
      end
      if(_zz_2282_)begin
        int_reg_array_32_55_imag <= _zz_2293_;
      end
      if(_zz_2283_)begin
        int_reg_array_32_56_imag <= _zz_2293_;
      end
      if(_zz_2284_)begin
        int_reg_array_32_57_imag <= _zz_2293_;
      end
      if(_zz_2285_)begin
        int_reg_array_32_58_imag <= _zz_2293_;
      end
      if(_zz_2286_)begin
        int_reg_array_32_59_imag <= _zz_2293_;
      end
      if(_zz_2287_)begin
        int_reg_array_32_60_imag <= _zz_2293_;
      end
      if(_zz_2288_)begin
        int_reg_array_32_61_imag <= _zz_2293_;
      end
      if(_zz_2289_)begin
        int_reg_array_32_62_imag <= _zz_2293_;
      end
      if(_zz_2290_)begin
        int_reg_array_32_63_imag <= _zz_2293_;
      end
      if(_zz_2296_)begin
        int_reg_array_33_0_real <= _zz_2361_;
      end
      if(_zz_2297_)begin
        int_reg_array_33_1_real <= _zz_2361_;
      end
      if(_zz_2298_)begin
        int_reg_array_33_2_real <= _zz_2361_;
      end
      if(_zz_2299_)begin
        int_reg_array_33_3_real <= _zz_2361_;
      end
      if(_zz_2300_)begin
        int_reg_array_33_4_real <= _zz_2361_;
      end
      if(_zz_2301_)begin
        int_reg_array_33_5_real <= _zz_2361_;
      end
      if(_zz_2302_)begin
        int_reg_array_33_6_real <= _zz_2361_;
      end
      if(_zz_2303_)begin
        int_reg_array_33_7_real <= _zz_2361_;
      end
      if(_zz_2304_)begin
        int_reg_array_33_8_real <= _zz_2361_;
      end
      if(_zz_2305_)begin
        int_reg_array_33_9_real <= _zz_2361_;
      end
      if(_zz_2306_)begin
        int_reg_array_33_10_real <= _zz_2361_;
      end
      if(_zz_2307_)begin
        int_reg_array_33_11_real <= _zz_2361_;
      end
      if(_zz_2308_)begin
        int_reg_array_33_12_real <= _zz_2361_;
      end
      if(_zz_2309_)begin
        int_reg_array_33_13_real <= _zz_2361_;
      end
      if(_zz_2310_)begin
        int_reg_array_33_14_real <= _zz_2361_;
      end
      if(_zz_2311_)begin
        int_reg_array_33_15_real <= _zz_2361_;
      end
      if(_zz_2312_)begin
        int_reg_array_33_16_real <= _zz_2361_;
      end
      if(_zz_2313_)begin
        int_reg_array_33_17_real <= _zz_2361_;
      end
      if(_zz_2314_)begin
        int_reg_array_33_18_real <= _zz_2361_;
      end
      if(_zz_2315_)begin
        int_reg_array_33_19_real <= _zz_2361_;
      end
      if(_zz_2316_)begin
        int_reg_array_33_20_real <= _zz_2361_;
      end
      if(_zz_2317_)begin
        int_reg_array_33_21_real <= _zz_2361_;
      end
      if(_zz_2318_)begin
        int_reg_array_33_22_real <= _zz_2361_;
      end
      if(_zz_2319_)begin
        int_reg_array_33_23_real <= _zz_2361_;
      end
      if(_zz_2320_)begin
        int_reg_array_33_24_real <= _zz_2361_;
      end
      if(_zz_2321_)begin
        int_reg_array_33_25_real <= _zz_2361_;
      end
      if(_zz_2322_)begin
        int_reg_array_33_26_real <= _zz_2361_;
      end
      if(_zz_2323_)begin
        int_reg_array_33_27_real <= _zz_2361_;
      end
      if(_zz_2324_)begin
        int_reg_array_33_28_real <= _zz_2361_;
      end
      if(_zz_2325_)begin
        int_reg_array_33_29_real <= _zz_2361_;
      end
      if(_zz_2326_)begin
        int_reg_array_33_30_real <= _zz_2361_;
      end
      if(_zz_2327_)begin
        int_reg_array_33_31_real <= _zz_2361_;
      end
      if(_zz_2328_)begin
        int_reg_array_33_32_real <= _zz_2361_;
      end
      if(_zz_2329_)begin
        int_reg_array_33_33_real <= _zz_2361_;
      end
      if(_zz_2330_)begin
        int_reg_array_33_34_real <= _zz_2361_;
      end
      if(_zz_2331_)begin
        int_reg_array_33_35_real <= _zz_2361_;
      end
      if(_zz_2332_)begin
        int_reg_array_33_36_real <= _zz_2361_;
      end
      if(_zz_2333_)begin
        int_reg_array_33_37_real <= _zz_2361_;
      end
      if(_zz_2334_)begin
        int_reg_array_33_38_real <= _zz_2361_;
      end
      if(_zz_2335_)begin
        int_reg_array_33_39_real <= _zz_2361_;
      end
      if(_zz_2336_)begin
        int_reg_array_33_40_real <= _zz_2361_;
      end
      if(_zz_2337_)begin
        int_reg_array_33_41_real <= _zz_2361_;
      end
      if(_zz_2338_)begin
        int_reg_array_33_42_real <= _zz_2361_;
      end
      if(_zz_2339_)begin
        int_reg_array_33_43_real <= _zz_2361_;
      end
      if(_zz_2340_)begin
        int_reg_array_33_44_real <= _zz_2361_;
      end
      if(_zz_2341_)begin
        int_reg_array_33_45_real <= _zz_2361_;
      end
      if(_zz_2342_)begin
        int_reg_array_33_46_real <= _zz_2361_;
      end
      if(_zz_2343_)begin
        int_reg_array_33_47_real <= _zz_2361_;
      end
      if(_zz_2344_)begin
        int_reg_array_33_48_real <= _zz_2361_;
      end
      if(_zz_2345_)begin
        int_reg_array_33_49_real <= _zz_2361_;
      end
      if(_zz_2346_)begin
        int_reg_array_33_50_real <= _zz_2361_;
      end
      if(_zz_2347_)begin
        int_reg_array_33_51_real <= _zz_2361_;
      end
      if(_zz_2348_)begin
        int_reg_array_33_52_real <= _zz_2361_;
      end
      if(_zz_2349_)begin
        int_reg_array_33_53_real <= _zz_2361_;
      end
      if(_zz_2350_)begin
        int_reg_array_33_54_real <= _zz_2361_;
      end
      if(_zz_2351_)begin
        int_reg_array_33_55_real <= _zz_2361_;
      end
      if(_zz_2352_)begin
        int_reg_array_33_56_real <= _zz_2361_;
      end
      if(_zz_2353_)begin
        int_reg_array_33_57_real <= _zz_2361_;
      end
      if(_zz_2354_)begin
        int_reg_array_33_58_real <= _zz_2361_;
      end
      if(_zz_2355_)begin
        int_reg_array_33_59_real <= _zz_2361_;
      end
      if(_zz_2356_)begin
        int_reg_array_33_60_real <= _zz_2361_;
      end
      if(_zz_2357_)begin
        int_reg_array_33_61_real <= _zz_2361_;
      end
      if(_zz_2358_)begin
        int_reg_array_33_62_real <= _zz_2361_;
      end
      if(_zz_2359_)begin
        int_reg_array_33_63_real <= _zz_2361_;
      end
      if(_zz_2296_)begin
        int_reg_array_33_0_imag <= _zz_2362_;
      end
      if(_zz_2297_)begin
        int_reg_array_33_1_imag <= _zz_2362_;
      end
      if(_zz_2298_)begin
        int_reg_array_33_2_imag <= _zz_2362_;
      end
      if(_zz_2299_)begin
        int_reg_array_33_3_imag <= _zz_2362_;
      end
      if(_zz_2300_)begin
        int_reg_array_33_4_imag <= _zz_2362_;
      end
      if(_zz_2301_)begin
        int_reg_array_33_5_imag <= _zz_2362_;
      end
      if(_zz_2302_)begin
        int_reg_array_33_6_imag <= _zz_2362_;
      end
      if(_zz_2303_)begin
        int_reg_array_33_7_imag <= _zz_2362_;
      end
      if(_zz_2304_)begin
        int_reg_array_33_8_imag <= _zz_2362_;
      end
      if(_zz_2305_)begin
        int_reg_array_33_9_imag <= _zz_2362_;
      end
      if(_zz_2306_)begin
        int_reg_array_33_10_imag <= _zz_2362_;
      end
      if(_zz_2307_)begin
        int_reg_array_33_11_imag <= _zz_2362_;
      end
      if(_zz_2308_)begin
        int_reg_array_33_12_imag <= _zz_2362_;
      end
      if(_zz_2309_)begin
        int_reg_array_33_13_imag <= _zz_2362_;
      end
      if(_zz_2310_)begin
        int_reg_array_33_14_imag <= _zz_2362_;
      end
      if(_zz_2311_)begin
        int_reg_array_33_15_imag <= _zz_2362_;
      end
      if(_zz_2312_)begin
        int_reg_array_33_16_imag <= _zz_2362_;
      end
      if(_zz_2313_)begin
        int_reg_array_33_17_imag <= _zz_2362_;
      end
      if(_zz_2314_)begin
        int_reg_array_33_18_imag <= _zz_2362_;
      end
      if(_zz_2315_)begin
        int_reg_array_33_19_imag <= _zz_2362_;
      end
      if(_zz_2316_)begin
        int_reg_array_33_20_imag <= _zz_2362_;
      end
      if(_zz_2317_)begin
        int_reg_array_33_21_imag <= _zz_2362_;
      end
      if(_zz_2318_)begin
        int_reg_array_33_22_imag <= _zz_2362_;
      end
      if(_zz_2319_)begin
        int_reg_array_33_23_imag <= _zz_2362_;
      end
      if(_zz_2320_)begin
        int_reg_array_33_24_imag <= _zz_2362_;
      end
      if(_zz_2321_)begin
        int_reg_array_33_25_imag <= _zz_2362_;
      end
      if(_zz_2322_)begin
        int_reg_array_33_26_imag <= _zz_2362_;
      end
      if(_zz_2323_)begin
        int_reg_array_33_27_imag <= _zz_2362_;
      end
      if(_zz_2324_)begin
        int_reg_array_33_28_imag <= _zz_2362_;
      end
      if(_zz_2325_)begin
        int_reg_array_33_29_imag <= _zz_2362_;
      end
      if(_zz_2326_)begin
        int_reg_array_33_30_imag <= _zz_2362_;
      end
      if(_zz_2327_)begin
        int_reg_array_33_31_imag <= _zz_2362_;
      end
      if(_zz_2328_)begin
        int_reg_array_33_32_imag <= _zz_2362_;
      end
      if(_zz_2329_)begin
        int_reg_array_33_33_imag <= _zz_2362_;
      end
      if(_zz_2330_)begin
        int_reg_array_33_34_imag <= _zz_2362_;
      end
      if(_zz_2331_)begin
        int_reg_array_33_35_imag <= _zz_2362_;
      end
      if(_zz_2332_)begin
        int_reg_array_33_36_imag <= _zz_2362_;
      end
      if(_zz_2333_)begin
        int_reg_array_33_37_imag <= _zz_2362_;
      end
      if(_zz_2334_)begin
        int_reg_array_33_38_imag <= _zz_2362_;
      end
      if(_zz_2335_)begin
        int_reg_array_33_39_imag <= _zz_2362_;
      end
      if(_zz_2336_)begin
        int_reg_array_33_40_imag <= _zz_2362_;
      end
      if(_zz_2337_)begin
        int_reg_array_33_41_imag <= _zz_2362_;
      end
      if(_zz_2338_)begin
        int_reg_array_33_42_imag <= _zz_2362_;
      end
      if(_zz_2339_)begin
        int_reg_array_33_43_imag <= _zz_2362_;
      end
      if(_zz_2340_)begin
        int_reg_array_33_44_imag <= _zz_2362_;
      end
      if(_zz_2341_)begin
        int_reg_array_33_45_imag <= _zz_2362_;
      end
      if(_zz_2342_)begin
        int_reg_array_33_46_imag <= _zz_2362_;
      end
      if(_zz_2343_)begin
        int_reg_array_33_47_imag <= _zz_2362_;
      end
      if(_zz_2344_)begin
        int_reg_array_33_48_imag <= _zz_2362_;
      end
      if(_zz_2345_)begin
        int_reg_array_33_49_imag <= _zz_2362_;
      end
      if(_zz_2346_)begin
        int_reg_array_33_50_imag <= _zz_2362_;
      end
      if(_zz_2347_)begin
        int_reg_array_33_51_imag <= _zz_2362_;
      end
      if(_zz_2348_)begin
        int_reg_array_33_52_imag <= _zz_2362_;
      end
      if(_zz_2349_)begin
        int_reg_array_33_53_imag <= _zz_2362_;
      end
      if(_zz_2350_)begin
        int_reg_array_33_54_imag <= _zz_2362_;
      end
      if(_zz_2351_)begin
        int_reg_array_33_55_imag <= _zz_2362_;
      end
      if(_zz_2352_)begin
        int_reg_array_33_56_imag <= _zz_2362_;
      end
      if(_zz_2353_)begin
        int_reg_array_33_57_imag <= _zz_2362_;
      end
      if(_zz_2354_)begin
        int_reg_array_33_58_imag <= _zz_2362_;
      end
      if(_zz_2355_)begin
        int_reg_array_33_59_imag <= _zz_2362_;
      end
      if(_zz_2356_)begin
        int_reg_array_33_60_imag <= _zz_2362_;
      end
      if(_zz_2357_)begin
        int_reg_array_33_61_imag <= _zz_2362_;
      end
      if(_zz_2358_)begin
        int_reg_array_33_62_imag <= _zz_2362_;
      end
      if(_zz_2359_)begin
        int_reg_array_33_63_imag <= _zz_2362_;
      end
      if(_zz_2365_)begin
        int_reg_array_34_0_real <= _zz_2430_;
      end
      if(_zz_2366_)begin
        int_reg_array_34_1_real <= _zz_2430_;
      end
      if(_zz_2367_)begin
        int_reg_array_34_2_real <= _zz_2430_;
      end
      if(_zz_2368_)begin
        int_reg_array_34_3_real <= _zz_2430_;
      end
      if(_zz_2369_)begin
        int_reg_array_34_4_real <= _zz_2430_;
      end
      if(_zz_2370_)begin
        int_reg_array_34_5_real <= _zz_2430_;
      end
      if(_zz_2371_)begin
        int_reg_array_34_6_real <= _zz_2430_;
      end
      if(_zz_2372_)begin
        int_reg_array_34_7_real <= _zz_2430_;
      end
      if(_zz_2373_)begin
        int_reg_array_34_8_real <= _zz_2430_;
      end
      if(_zz_2374_)begin
        int_reg_array_34_9_real <= _zz_2430_;
      end
      if(_zz_2375_)begin
        int_reg_array_34_10_real <= _zz_2430_;
      end
      if(_zz_2376_)begin
        int_reg_array_34_11_real <= _zz_2430_;
      end
      if(_zz_2377_)begin
        int_reg_array_34_12_real <= _zz_2430_;
      end
      if(_zz_2378_)begin
        int_reg_array_34_13_real <= _zz_2430_;
      end
      if(_zz_2379_)begin
        int_reg_array_34_14_real <= _zz_2430_;
      end
      if(_zz_2380_)begin
        int_reg_array_34_15_real <= _zz_2430_;
      end
      if(_zz_2381_)begin
        int_reg_array_34_16_real <= _zz_2430_;
      end
      if(_zz_2382_)begin
        int_reg_array_34_17_real <= _zz_2430_;
      end
      if(_zz_2383_)begin
        int_reg_array_34_18_real <= _zz_2430_;
      end
      if(_zz_2384_)begin
        int_reg_array_34_19_real <= _zz_2430_;
      end
      if(_zz_2385_)begin
        int_reg_array_34_20_real <= _zz_2430_;
      end
      if(_zz_2386_)begin
        int_reg_array_34_21_real <= _zz_2430_;
      end
      if(_zz_2387_)begin
        int_reg_array_34_22_real <= _zz_2430_;
      end
      if(_zz_2388_)begin
        int_reg_array_34_23_real <= _zz_2430_;
      end
      if(_zz_2389_)begin
        int_reg_array_34_24_real <= _zz_2430_;
      end
      if(_zz_2390_)begin
        int_reg_array_34_25_real <= _zz_2430_;
      end
      if(_zz_2391_)begin
        int_reg_array_34_26_real <= _zz_2430_;
      end
      if(_zz_2392_)begin
        int_reg_array_34_27_real <= _zz_2430_;
      end
      if(_zz_2393_)begin
        int_reg_array_34_28_real <= _zz_2430_;
      end
      if(_zz_2394_)begin
        int_reg_array_34_29_real <= _zz_2430_;
      end
      if(_zz_2395_)begin
        int_reg_array_34_30_real <= _zz_2430_;
      end
      if(_zz_2396_)begin
        int_reg_array_34_31_real <= _zz_2430_;
      end
      if(_zz_2397_)begin
        int_reg_array_34_32_real <= _zz_2430_;
      end
      if(_zz_2398_)begin
        int_reg_array_34_33_real <= _zz_2430_;
      end
      if(_zz_2399_)begin
        int_reg_array_34_34_real <= _zz_2430_;
      end
      if(_zz_2400_)begin
        int_reg_array_34_35_real <= _zz_2430_;
      end
      if(_zz_2401_)begin
        int_reg_array_34_36_real <= _zz_2430_;
      end
      if(_zz_2402_)begin
        int_reg_array_34_37_real <= _zz_2430_;
      end
      if(_zz_2403_)begin
        int_reg_array_34_38_real <= _zz_2430_;
      end
      if(_zz_2404_)begin
        int_reg_array_34_39_real <= _zz_2430_;
      end
      if(_zz_2405_)begin
        int_reg_array_34_40_real <= _zz_2430_;
      end
      if(_zz_2406_)begin
        int_reg_array_34_41_real <= _zz_2430_;
      end
      if(_zz_2407_)begin
        int_reg_array_34_42_real <= _zz_2430_;
      end
      if(_zz_2408_)begin
        int_reg_array_34_43_real <= _zz_2430_;
      end
      if(_zz_2409_)begin
        int_reg_array_34_44_real <= _zz_2430_;
      end
      if(_zz_2410_)begin
        int_reg_array_34_45_real <= _zz_2430_;
      end
      if(_zz_2411_)begin
        int_reg_array_34_46_real <= _zz_2430_;
      end
      if(_zz_2412_)begin
        int_reg_array_34_47_real <= _zz_2430_;
      end
      if(_zz_2413_)begin
        int_reg_array_34_48_real <= _zz_2430_;
      end
      if(_zz_2414_)begin
        int_reg_array_34_49_real <= _zz_2430_;
      end
      if(_zz_2415_)begin
        int_reg_array_34_50_real <= _zz_2430_;
      end
      if(_zz_2416_)begin
        int_reg_array_34_51_real <= _zz_2430_;
      end
      if(_zz_2417_)begin
        int_reg_array_34_52_real <= _zz_2430_;
      end
      if(_zz_2418_)begin
        int_reg_array_34_53_real <= _zz_2430_;
      end
      if(_zz_2419_)begin
        int_reg_array_34_54_real <= _zz_2430_;
      end
      if(_zz_2420_)begin
        int_reg_array_34_55_real <= _zz_2430_;
      end
      if(_zz_2421_)begin
        int_reg_array_34_56_real <= _zz_2430_;
      end
      if(_zz_2422_)begin
        int_reg_array_34_57_real <= _zz_2430_;
      end
      if(_zz_2423_)begin
        int_reg_array_34_58_real <= _zz_2430_;
      end
      if(_zz_2424_)begin
        int_reg_array_34_59_real <= _zz_2430_;
      end
      if(_zz_2425_)begin
        int_reg_array_34_60_real <= _zz_2430_;
      end
      if(_zz_2426_)begin
        int_reg_array_34_61_real <= _zz_2430_;
      end
      if(_zz_2427_)begin
        int_reg_array_34_62_real <= _zz_2430_;
      end
      if(_zz_2428_)begin
        int_reg_array_34_63_real <= _zz_2430_;
      end
      if(_zz_2365_)begin
        int_reg_array_34_0_imag <= _zz_2431_;
      end
      if(_zz_2366_)begin
        int_reg_array_34_1_imag <= _zz_2431_;
      end
      if(_zz_2367_)begin
        int_reg_array_34_2_imag <= _zz_2431_;
      end
      if(_zz_2368_)begin
        int_reg_array_34_3_imag <= _zz_2431_;
      end
      if(_zz_2369_)begin
        int_reg_array_34_4_imag <= _zz_2431_;
      end
      if(_zz_2370_)begin
        int_reg_array_34_5_imag <= _zz_2431_;
      end
      if(_zz_2371_)begin
        int_reg_array_34_6_imag <= _zz_2431_;
      end
      if(_zz_2372_)begin
        int_reg_array_34_7_imag <= _zz_2431_;
      end
      if(_zz_2373_)begin
        int_reg_array_34_8_imag <= _zz_2431_;
      end
      if(_zz_2374_)begin
        int_reg_array_34_9_imag <= _zz_2431_;
      end
      if(_zz_2375_)begin
        int_reg_array_34_10_imag <= _zz_2431_;
      end
      if(_zz_2376_)begin
        int_reg_array_34_11_imag <= _zz_2431_;
      end
      if(_zz_2377_)begin
        int_reg_array_34_12_imag <= _zz_2431_;
      end
      if(_zz_2378_)begin
        int_reg_array_34_13_imag <= _zz_2431_;
      end
      if(_zz_2379_)begin
        int_reg_array_34_14_imag <= _zz_2431_;
      end
      if(_zz_2380_)begin
        int_reg_array_34_15_imag <= _zz_2431_;
      end
      if(_zz_2381_)begin
        int_reg_array_34_16_imag <= _zz_2431_;
      end
      if(_zz_2382_)begin
        int_reg_array_34_17_imag <= _zz_2431_;
      end
      if(_zz_2383_)begin
        int_reg_array_34_18_imag <= _zz_2431_;
      end
      if(_zz_2384_)begin
        int_reg_array_34_19_imag <= _zz_2431_;
      end
      if(_zz_2385_)begin
        int_reg_array_34_20_imag <= _zz_2431_;
      end
      if(_zz_2386_)begin
        int_reg_array_34_21_imag <= _zz_2431_;
      end
      if(_zz_2387_)begin
        int_reg_array_34_22_imag <= _zz_2431_;
      end
      if(_zz_2388_)begin
        int_reg_array_34_23_imag <= _zz_2431_;
      end
      if(_zz_2389_)begin
        int_reg_array_34_24_imag <= _zz_2431_;
      end
      if(_zz_2390_)begin
        int_reg_array_34_25_imag <= _zz_2431_;
      end
      if(_zz_2391_)begin
        int_reg_array_34_26_imag <= _zz_2431_;
      end
      if(_zz_2392_)begin
        int_reg_array_34_27_imag <= _zz_2431_;
      end
      if(_zz_2393_)begin
        int_reg_array_34_28_imag <= _zz_2431_;
      end
      if(_zz_2394_)begin
        int_reg_array_34_29_imag <= _zz_2431_;
      end
      if(_zz_2395_)begin
        int_reg_array_34_30_imag <= _zz_2431_;
      end
      if(_zz_2396_)begin
        int_reg_array_34_31_imag <= _zz_2431_;
      end
      if(_zz_2397_)begin
        int_reg_array_34_32_imag <= _zz_2431_;
      end
      if(_zz_2398_)begin
        int_reg_array_34_33_imag <= _zz_2431_;
      end
      if(_zz_2399_)begin
        int_reg_array_34_34_imag <= _zz_2431_;
      end
      if(_zz_2400_)begin
        int_reg_array_34_35_imag <= _zz_2431_;
      end
      if(_zz_2401_)begin
        int_reg_array_34_36_imag <= _zz_2431_;
      end
      if(_zz_2402_)begin
        int_reg_array_34_37_imag <= _zz_2431_;
      end
      if(_zz_2403_)begin
        int_reg_array_34_38_imag <= _zz_2431_;
      end
      if(_zz_2404_)begin
        int_reg_array_34_39_imag <= _zz_2431_;
      end
      if(_zz_2405_)begin
        int_reg_array_34_40_imag <= _zz_2431_;
      end
      if(_zz_2406_)begin
        int_reg_array_34_41_imag <= _zz_2431_;
      end
      if(_zz_2407_)begin
        int_reg_array_34_42_imag <= _zz_2431_;
      end
      if(_zz_2408_)begin
        int_reg_array_34_43_imag <= _zz_2431_;
      end
      if(_zz_2409_)begin
        int_reg_array_34_44_imag <= _zz_2431_;
      end
      if(_zz_2410_)begin
        int_reg_array_34_45_imag <= _zz_2431_;
      end
      if(_zz_2411_)begin
        int_reg_array_34_46_imag <= _zz_2431_;
      end
      if(_zz_2412_)begin
        int_reg_array_34_47_imag <= _zz_2431_;
      end
      if(_zz_2413_)begin
        int_reg_array_34_48_imag <= _zz_2431_;
      end
      if(_zz_2414_)begin
        int_reg_array_34_49_imag <= _zz_2431_;
      end
      if(_zz_2415_)begin
        int_reg_array_34_50_imag <= _zz_2431_;
      end
      if(_zz_2416_)begin
        int_reg_array_34_51_imag <= _zz_2431_;
      end
      if(_zz_2417_)begin
        int_reg_array_34_52_imag <= _zz_2431_;
      end
      if(_zz_2418_)begin
        int_reg_array_34_53_imag <= _zz_2431_;
      end
      if(_zz_2419_)begin
        int_reg_array_34_54_imag <= _zz_2431_;
      end
      if(_zz_2420_)begin
        int_reg_array_34_55_imag <= _zz_2431_;
      end
      if(_zz_2421_)begin
        int_reg_array_34_56_imag <= _zz_2431_;
      end
      if(_zz_2422_)begin
        int_reg_array_34_57_imag <= _zz_2431_;
      end
      if(_zz_2423_)begin
        int_reg_array_34_58_imag <= _zz_2431_;
      end
      if(_zz_2424_)begin
        int_reg_array_34_59_imag <= _zz_2431_;
      end
      if(_zz_2425_)begin
        int_reg_array_34_60_imag <= _zz_2431_;
      end
      if(_zz_2426_)begin
        int_reg_array_34_61_imag <= _zz_2431_;
      end
      if(_zz_2427_)begin
        int_reg_array_34_62_imag <= _zz_2431_;
      end
      if(_zz_2428_)begin
        int_reg_array_34_63_imag <= _zz_2431_;
      end
      if(_zz_2434_)begin
        int_reg_array_35_0_real <= _zz_2499_;
      end
      if(_zz_2435_)begin
        int_reg_array_35_1_real <= _zz_2499_;
      end
      if(_zz_2436_)begin
        int_reg_array_35_2_real <= _zz_2499_;
      end
      if(_zz_2437_)begin
        int_reg_array_35_3_real <= _zz_2499_;
      end
      if(_zz_2438_)begin
        int_reg_array_35_4_real <= _zz_2499_;
      end
      if(_zz_2439_)begin
        int_reg_array_35_5_real <= _zz_2499_;
      end
      if(_zz_2440_)begin
        int_reg_array_35_6_real <= _zz_2499_;
      end
      if(_zz_2441_)begin
        int_reg_array_35_7_real <= _zz_2499_;
      end
      if(_zz_2442_)begin
        int_reg_array_35_8_real <= _zz_2499_;
      end
      if(_zz_2443_)begin
        int_reg_array_35_9_real <= _zz_2499_;
      end
      if(_zz_2444_)begin
        int_reg_array_35_10_real <= _zz_2499_;
      end
      if(_zz_2445_)begin
        int_reg_array_35_11_real <= _zz_2499_;
      end
      if(_zz_2446_)begin
        int_reg_array_35_12_real <= _zz_2499_;
      end
      if(_zz_2447_)begin
        int_reg_array_35_13_real <= _zz_2499_;
      end
      if(_zz_2448_)begin
        int_reg_array_35_14_real <= _zz_2499_;
      end
      if(_zz_2449_)begin
        int_reg_array_35_15_real <= _zz_2499_;
      end
      if(_zz_2450_)begin
        int_reg_array_35_16_real <= _zz_2499_;
      end
      if(_zz_2451_)begin
        int_reg_array_35_17_real <= _zz_2499_;
      end
      if(_zz_2452_)begin
        int_reg_array_35_18_real <= _zz_2499_;
      end
      if(_zz_2453_)begin
        int_reg_array_35_19_real <= _zz_2499_;
      end
      if(_zz_2454_)begin
        int_reg_array_35_20_real <= _zz_2499_;
      end
      if(_zz_2455_)begin
        int_reg_array_35_21_real <= _zz_2499_;
      end
      if(_zz_2456_)begin
        int_reg_array_35_22_real <= _zz_2499_;
      end
      if(_zz_2457_)begin
        int_reg_array_35_23_real <= _zz_2499_;
      end
      if(_zz_2458_)begin
        int_reg_array_35_24_real <= _zz_2499_;
      end
      if(_zz_2459_)begin
        int_reg_array_35_25_real <= _zz_2499_;
      end
      if(_zz_2460_)begin
        int_reg_array_35_26_real <= _zz_2499_;
      end
      if(_zz_2461_)begin
        int_reg_array_35_27_real <= _zz_2499_;
      end
      if(_zz_2462_)begin
        int_reg_array_35_28_real <= _zz_2499_;
      end
      if(_zz_2463_)begin
        int_reg_array_35_29_real <= _zz_2499_;
      end
      if(_zz_2464_)begin
        int_reg_array_35_30_real <= _zz_2499_;
      end
      if(_zz_2465_)begin
        int_reg_array_35_31_real <= _zz_2499_;
      end
      if(_zz_2466_)begin
        int_reg_array_35_32_real <= _zz_2499_;
      end
      if(_zz_2467_)begin
        int_reg_array_35_33_real <= _zz_2499_;
      end
      if(_zz_2468_)begin
        int_reg_array_35_34_real <= _zz_2499_;
      end
      if(_zz_2469_)begin
        int_reg_array_35_35_real <= _zz_2499_;
      end
      if(_zz_2470_)begin
        int_reg_array_35_36_real <= _zz_2499_;
      end
      if(_zz_2471_)begin
        int_reg_array_35_37_real <= _zz_2499_;
      end
      if(_zz_2472_)begin
        int_reg_array_35_38_real <= _zz_2499_;
      end
      if(_zz_2473_)begin
        int_reg_array_35_39_real <= _zz_2499_;
      end
      if(_zz_2474_)begin
        int_reg_array_35_40_real <= _zz_2499_;
      end
      if(_zz_2475_)begin
        int_reg_array_35_41_real <= _zz_2499_;
      end
      if(_zz_2476_)begin
        int_reg_array_35_42_real <= _zz_2499_;
      end
      if(_zz_2477_)begin
        int_reg_array_35_43_real <= _zz_2499_;
      end
      if(_zz_2478_)begin
        int_reg_array_35_44_real <= _zz_2499_;
      end
      if(_zz_2479_)begin
        int_reg_array_35_45_real <= _zz_2499_;
      end
      if(_zz_2480_)begin
        int_reg_array_35_46_real <= _zz_2499_;
      end
      if(_zz_2481_)begin
        int_reg_array_35_47_real <= _zz_2499_;
      end
      if(_zz_2482_)begin
        int_reg_array_35_48_real <= _zz_2499_;
      end
      if(_zz_2483_)begin
        int_reg_array_35_49_real <= _zz_2499_;
      end
      if(_zz_2484_)begin
        int_reg_array_35_50_real <= _zz_2499_;
      end
      if(_zz_2485_)begin
        int_reg_array_35_51_real <= _zz_2499_;
      end
      if(_zz_2486_)begin
        int_reg_array_35_52_real <= _zz_2499_;
      end
      if(_zz_2487_)begin
        int_reg_array_35_53_real <= _zz_2499_;
      end
      if(_zz_2488_)begin
        int_reg_array_35_54_real <= _zz_2499_;
      end
      if(_zz_2489_)begin
        int_reg_array_35_55_real <= _zz_2499_;
      end
      if(_zz_2490_)begin
        int_reg_array_35_56_real <= _zz_2499_;
      end
      if(_zz_2491_)begin
        int_reg_array_35_57_real <= _zz_2499_;
      end
      if(_zz_2492_)begin
        int_reg_array_35_58_real <= _zz_2499_;
      end
      if(_zz_2493_)begin
        int_reg_array_35_59_real <= _zz_2499_;
      end
      if(_zz_2494_)begin
        int_reg_array_35_60_real <= _zz_2499_;
      end
      if(_zz_2495_)begin
        int_reg_array_35_61_real <= _zz_2499_;
      end
      if(_zz_2496_)begin
        int_reg_array_35_62_real <= _zz_2499_;
      end
      if(_zz_2497_)begin
        int_reg_array_35_63_real <= _zz_2499_;
      end
      if(_zz_2434_)begin
        int_reg_array_35_0_imag <= _zz_2500_;
      end
      if(_zz_2435_)begin
        int_reg_array_35_1_imag <= _zz_2500_;
      end
      if(_zz_2436_)begin
        int_reg_array_35_2_imag <= _zz_2500_;
      end
      if(_zz_2437_)begin
        int_reg_array_35_3_imag <= _zz_2500_;
      end
      if(_zz_2438_)begin
        int_reg_array_35_4_imag <= _zz_2500_;
      end
      if(_zz_2439_)begin
        int_reg_array_35_5_imag <= _zz_2500_;
      end
      if(_zz_2440_)begin
        int_reg_array_35_6_imag <= _zz_2500_;
      end
      if(_zz_2441_)begin
        int_reg_array_35_7_imag <= _zz_2500_;
      end
      if(_zz_2442_)begin
        int_reg_array_35_8_imag <= _zz_2500_;
      end
      if(_zz_2443_)begin
        int_reg_array_35_9_imag <= _zz_2500_;
      end
      if(_zz_2444_)begin
        int_reg_array_35_10_imag <= _zz_2500_;
      end
      if(_zz_2445_)begin
        int_reg_array_35_11_imag <= _zz_2500_;
      end
      if(_zz_2446_)begin
        int_reg_array_35_12_imag <= _zz_2500_;
      end
      if(_zz_2447_)begin
        int_reg_array_35_13_imag <= _zz_2500_;
      end
      if(_zz_2448_)begin
        int_reg_array_35_14_imag <= _zz_2500_;
      end
      if(_zz_2449_)begin
        int_reg_array_35_15_imag <= _zz_2500_;
      end
      if(_zz_2450_)begin
        int_reg_array_35_16_imag <= _zz_2500_;
      end
      if(_zz_2451_)begin
        int_reg_array_35_17_imag <= _zz_2500_;
      end
      if(_zz_2452_)begin
        int_reg_array_35_18_imag <= _zz_2500_;
      end
      if(_zz_2453_)begin
        int_reg_array_35_19_imag <= _zz_2500_;
      end
      if(_zz_2454_)begin
        int_reg_array_35_20_imag <= _zz_2500_;
      end
      if(_zz_2455_)begin
        int_reg_array_35_21_imag <= _zz_2500_;
      end
      if(_zz_2456_)begin
        int_reg_array_35_22_imag <= _zz_2500_;
      end
      if(_zz_2457_)begin
        int_reg_array_35_23_imag <= _zz_2500_;
      end
      if(_zz_2458_)begin
        int_reg_array_35_24_imag <= _zz_2500_;
      end
      if(_zz_2459_)begin
        int_reg_array_35_25_imag <= _zz_2500_;
      end
      if(_zz_2460_)begin
        int_reg_array_35_26_imag <= _zz_2500_;
      end
      if(_zz_2461_)begin
        int_reg_array_35_27_imag <= _zz_2500_;
      end
      if(_zz_2462_)begin
        int_reg_array_35_28_imag <= _zz_2500_;
      end
      if(_zz_2463_)begin
        int_reg_array_35_29_imag <= _zz_2500_;
      end
      if(_zz_2464_)begin
        int_reg_array_35_30_imag <= _zz_2500_;
      end
      if(_zz_2465_)begin
        int_reg_array_35_31_imag <= _zz_2500_;
      end
      if(_zz_2466_)begin
        int_reg_array_35_32_imag <= _zz_2500_;
      end
      if(_zz_2467_)begin
        int_reg_array_35_33_imag <= _zz_2500_;
      end
      if(_zz_2468_)begin
        int_reg_array_35_34_imag <= _zz_2500_;
      end
      if(_zz_2469_)begin
        int_reg_array_35_35_imag <= _zz_2500_;
      end
      if(_zz_2470_)begin
        int_reg_array_35_36_imag <= _zz_2500_;
      end
      if(_zz_2471_)begin
        int_reg_array_35_37_imag <= _zz_2500_;
      end
      if(_zz_2472_)begin
        int_reg_array_35_38_imag <= _zz_2500_;
      end
      if(_zz_2473_)begin
        int_reg_array_35_39_imag <= _zz_2500_;
      end
      if(_zz_2474_)begin
        int_reg_array_35_40_imag <= _zz_2500_;
      end
      if(_zz_2475_)begin
        int_reg_array_35_41_imag <= _zz_2500_;
      end
      if(_zz_2476_)begin
        int_reg_array_35_42_imag <= _zz_2500_;
      end
      if(_zz_2477_)begin
        int_reg_array_35_43_imag <= _zz_2500_;
      end
      if(_zz_2478_)begin
        int_reg_array_35_44_imag <= _zz_2500_;
      end
      if(_zz_2479_)begin
        int_reg_array_35_45_imag <= _zz_2500_;
      end
      if(_zz_2480_)begin
        int_reg_array_35_46_imag <= _zz_2500_;
      end
      if(_zz_2481_)begin
        int_reg_array_35_47_imag <= _zz_2500_;
      end
      if(_zz_2482_)begin
        int_reg_array_35_48_imag <= _zz_2500_;
      end
      if(_zz_2483_)begin
        int_reg_array_35_49_imag <= _zz_2500_;
      end
      if(_zz_2484_)begin
        int_reg_array_35_50_imag <= _zz_2500_;
      end
      if(_zz_2485_)begin
        int_reg_array_35_51_imag <= _zz_2500_;
      end
      if(_zz_2486_)begin
        int_reg_array_35_52_imag <= _zz_2500_;
      end
      if(_zz_2487_)begin
        int_reg_array_35_53_imag <= _zz_2500_;
      end
      if(_zz_2488_)begin
        int_reg_array_35_54_imag <= _zz_2500_;
      end
      if(_zz_2489_)begin
        int_reg_array_35_55_imag <= _zz_2500_;
      end
      if(_zz_2490_)begin
        int_reg_array_35_56_imag <= _zz_2500_;
      end
      if(_zz_2491_)begin
        int_reg_array_35_57_imag <= _zz_2500_;
      end
      if(_zz_2492_)begin
        int_reg_array_35_58_imag <= _zz_2500_;
      end
      if(_zz_2493_)begin
        int_reg_array_35_59_imag <= _zz_2500_;
      end
      if(_zz_2494_)begin
        int_reg_array_35_60_imag <= _zz_2500_;
      end
      if(_zz_2495_)begin
        int_reg_array_35_61_imag <= _zz_2500_;
      end
      if(_zz_2496_)begin
        int_reg_array_35_62_imag <= _zz_2500_;
      end
      if(_zz_2497_)begin
        int_reg_array_35_63_imag <= _zz_2500_;
      end
      if(_zz_2503_)begin
        int_reg_array_36_0_real <= _zz_2568_;
      end
      if(_zz_2504_)begin
        int_reg_array_36_1_real <= _zz_2568_;
      end
      if(_zz_2505_)begin
        int_reg_array_36_2_real <= _zz_2568_;
      end
      if(_zz_2506_)begin
        int_reg_array_36_3_real <= _zz_2568_;
      end
      if(_zz_2507_)begin
        int_reg_array_36_4_real <= _zz_2568_;
      end
      if(_zz_2508_)begin
        int_reg_array_36_5_real <= _zz_2568_;
      end
      if(_zz_2509_)begin
        int_reg_array_36_6_real <= _zz_2568_;
      end
      if(_zz_2510_)begin
        int_reg_array_36_7_real <= _zz_2568_;
      end
      if(_zz_2511_)begin
        int_reg_array_36_8_real <= _zz_2568_;
      end
      if(_zz_2512_)begin
        int_reg_array_36_9_real <= _zz_2568_;
      end
      if(_zz_2513_)begin
        int_reg_array_36_10_real <= _zz_2568_;
      end
      if(_zz_2514_)begin
        int_reg_array_36_11_real <= _zz_2568_;
      end
      if(_zz_2515_)begin
        int_reg_array_36_12_real <= _zz_2568_;
      end
      if(_zz_2516_)begin
        int_reg_array_36_13_real <= _zz_2568_;
      end
      if(_zz_2517_)begin
        int_reg_array_36_14_real <= _zz_2568_;
      end
      if(_zz_2518_)begin
        int_reg_array_36_15_real <= _zz_2568_;
      end
      if(_zz_2519_)begin
        int_reg_array_36_16_real <= _zz_2568_;
      end
      if(_zz_2520_)begin
        int_reg_array_36_17_real <= _zz_2568_;
      end
      if(_zz_2521_)begin
        int_reg_array_36_18_real <= _zz_2568_;
      end
      if(_zz_2522_)begin
        int_reg_array_36_19_real <= _zz_2568_;
      end
      if(_zz_2523_)begin
        int_reg_array_36_20_real <= _zz_2568_;
      end
      if(_zz_2524_)begin
        int_reg_array_36_21_real <= _zz_2568_;
      end
      if(_zz_2525_)begin
        int_reg_array_36_22_real <= _zz_2568_;
      end
      if(_zz_2526_)begin
        int_reg_array_36_23_real <= _zz_2568_;
      end
      if(_zz_2527_)begin
        int_reg_array_36_24_real <= _zz_2568_;
      end
      if(_zz_2528_)begin
        int_reg_array_36_25_real <= _zz_2568_;
      end
      if(_zz_2529_)begin
        int_reg_array_36_26_real <= _zz_2568_;
      end
      if(_zz_2530_)begin
        int_reg_array_36_27_real <= _zz_2568_;
      end
      if(_zz_2531_)begin
        int_reg_array_36_28_real <= _zz_2568_;
      end
      if(_zz_2532_)begin
        int_reg_array_36_29_real <= _zz_2568_;
      end
      if(_zz_2533_)begin
        int_reg_array_36_30_real <= _zz_2568_;
      end
      if(_zz_2534_)begin
        int_reg_array_36_31_real <= _zz_2568_;
      end
      if(_zz_2535_)begin
        int_reg_array_36_32_real <= _zz_2568_;
      end
      if(_zz_2536_)begin
        int_reg_array_36_33_real <= _zz_2568_;
      end
      if(_zz_2537_)begin
        int_reg_array_36_34_real <= _zz_2568_;
      end
      if(_zz_2538_)begin
        int_reg_array_36_35_real <= _zz_2568_;
      end
      if(_zz_2539_)begin
        int_reg_array_36_36_real <= _zz_2568_;
      end
      if(_zz_2540_)begin
        int_reg_array_36_37_real <= _zz_2568_;
      end
      if(_zz_2541_)begin
        int_reg_array_36_38_real <= _zz_2568_;
      end
      if(_zz_2542_)begin
        int_reg_array_36_39_real <= _zz_2568_;
      end
      if(_zz_2543_)begin
        int_reg_array_36_40_real <= _zz_2568_;
      end
      if(_zz_2544_)begin
        int_reg_array_36_41_real <= _zz_2568_;
      end
      if(_zz_2545_)begin
        int_reg_array_36_42_real <= _zz_2568_;
      end
      if(_zz_2546_)begin
        int_reg_array_36_43_real <= _zz_2568_;
      end
      if(_zz_2547_)begin
        int_reg_array_36_44_real <= _zz_2568_;
      end
      if(_zz_2548_)begin
        int_reg_array_36_45_real <= _zz_2568_;
      end
      if(_zz_2549_)begin
        int_reg_array_36_46_real <= _zz_2568_;
      end
      if(_zz_2550_)begin
        int_reg_array_36_47_real <= _zz_2568_;
      end
      if(_zz_2551_)begin
        int_reg_array_36_48_real <= _zz_2568_;
      end
      if(_zz_2552_)begin
        int_reg_array_36_49_real <= _zz_2568_;
      end
      if(_zz_2553_)begin
        int_reg_array_36_50_real <= _zz_2568_;
      end
      if(_zz_2554_)begin
        int_reg_array_36_51_real <= _zz_2568_;
      end
      if(_zz_2555_)begin
        int_reg_array_36_52_real <= _zz_2568_;
      end
      if(_zz_2556_)begin
        int_reg_array_36_53_real <= _zz_2568_;
      end
      if(_zz_2557_)begin
        int_reg_array_36_54_real <= _zz_2568_;
      end
      if(_zz_2558_)begin
        int_reg_array_36_55_real <= _zz_2568_;
      end
      if(_zz_2559_)begin
        int_reg_array_36_56_real <= _zz_2568_;
      end
      if(_zz_2560_)begin
        int_reg_array_36_57_real <= _zz_2568_;
      end
      if(_zz_2561_)begin
        int_reg_array_36_58_real <= _zz_2568_;
      end
      if(_zz_2562_)begin
        int_reg_array_36_59_real <= _zz_2568_;
      end
      if(_zz_2563_)begin
        int_reg_array_36_60_real <= _zz_2568_;
      end
      if(_zz_2564_)begin
        int_reg_array_36_61_real <= _zz_2568_;
      end
      if(_zz_2565_)begin
        int_reg_array_36_62_real <= _zz_2568_;
      end
      if(_zz_2566_)begin
        int_reg_array_36_63_real <= _zz_2568_;
      end
      if(_zz_2503_)begin
        int_reg_array_36_0_imag <= _zz_2569_;
      end
      if(_zz_2504_)begin
        int_reg_array_36_1_imag <= _zz_2569_;
      end
      if(_zz_2505_)begin
        int_reg_array_36_2_imag <= _zz_2569_;
      end
      if(_zz_2506_)begin
        int_reg_array_36_3_imag <= _zz_2569_;
      end
      if(_zz_2507_)begin
        int_reg_array_36_4_imag <= _zz_2569_;
      end
      if(_zz_2508_)begin
        int_reg_array_36_5_imag <= _zz_2569_;
      end
      if(_zz_2509_)begin
        int_reg_array_36_6_imag <= _zz_2569_;
      end
      if(_zz_2510_)begin
        int_reg_array_36_7_imag <= _zz_2569_;
      end
      if(_zz_2511_)begin
        int_reg_array_36_8_imag <= _zz_2569_;
      end
      if(_zz_2512_)begin
        int_reg_array_36_9_imag <= _zz_2569_;
      end
      if(_zz_2513_)begin
        int_reg_array_36_10_imag <= _zz_2569_;
      end
      if(_zz_2514_)begin
        int_reg_array_36_11_imag <= _zz_2569_;
      end
      if(_zz_2515_)begin
        int_reg_array_36_12_imag <= _zz_2569_;
      end
      if(_zz_2516_)begin
        int_reg_array_36_13_imag <= _zz_2569_;
      end
      if(_zz_2517_)begin
        int_reg_array_36_14_imag <= _zz_2569_;
      end
      if(_zz_2518_)begin
        int_reg_array_36_15_imag <= _zz_2569_;
      end
      if(_zz_2519_)begin
        int_reg_array_36_16_imag <= _zz_2569_;
      end
      if(_zz_2520_)begin
        int_reg_array_36_17_imag <= _zz_2569_;
      end
      if(_zz_2521_)begin
        int_reg_array_36_18_imag <= _zz_2569_;
      end
      if(_zz_2522_)begin
        int_reg_array_36_19_imag <= _zz_2569_;
      end
      if(_zz_2523_)begin
        int_reg_array_36_20_imag <= _zz_2569_;
      end
      if(_zz_2524_)begin
        int_reg_array_36_21_imag <= _zz_2569_;
      end
      if(_zz_2525_)begin
        int_reg_array_36_22_imag <= _zz_2569_;
      end
      if(_zz_2526_)begin
        int_reg_array_36_23_imag <= _zz_2569_;
      end
      if(_zz_2527_)begin
        int_reg_array_36_24_imag <= _zz_2569_;
      end
      if(_zz_2528_)begin
        int_reg_array_36_25_imag <= _zz_2569_;
      end
      if(_zz_2529_)begin
        int_reg_array_36_26_imag <= _zz_2569_;
      end
      if(_zz_2530_)begin
        int_reg_array_36_27_imag <= _zz_2569_;
      end
      if(_zz_2531_)begin
        int_reg_array_36_28_imag <= _zz_2569_;
      end
      if(_zz_2532_)begin
        int_reg_array_36_29_imag <= _zz_2569_;
      end
      if(_zz_2533_)begin
        int_reg_array_36_30_imag <= _zz_2569_;
      end
      if(_zz_2534_)begin
        int_reg_array_36_31_imag <= _zz_2569_;
      end
      if(_zz_2535_)begin
        int_reg_array_36_32_imag <= _zz_2569_;
      end
      if(_zz_2536_)begin
        int_reg_array_36_33_imag <= _zz_2569_;
      end
      if(_zz_2537_)begin
        int_reg_array_36_34_imag <= _zz_2569_;
      end
      if(_zz_2538_)begin
        int_reg_array_36_35_imag <= _zz_2569_;
      end
      if(_zz_2539_)begin
        int_reg_array_36_36_imag <= _zz_2569_;
      end
      if(_zz_2540_)begin
        int_reg_array_36_37_imag <= _zz_2569_;
      end
      if(_zz_2541_)begin
        int_reg_array_36_38_imag <= _zz_2569_;
      end
      if(_zz_2542_)begin
        int_reg_array_36_39_imag <= _zz_2569_;
      end
      if(_zz_2543_)begin
        int_reg_array_36_40_imag <= _zz_2569_;
      end
      if(_zz_2544_)begin
        int_reg_array_36_41_imag <= _zz_2569_;
      end
      if(_zz_2545_)begin
        int_reg_array_36_42_imag <= _zz_2569_;
      end
      if(_zz_2546_)begin
        int_reg_array_36_43_imag <= _zz_2569_;
      end
      if(_zz_2547_)begin
        int_reg_array_36_44_imag <= _zz_2569_;
      end
      if(_zz_2548_)begin
        int_reg_array_36_45_imag <= _zz_2569_;
      end
      if(_zz_2549_)begin
        int_reg_array_36_46_imag <= _zz_2569_;
      end
      if(_zz_2550_)begin
        int_reg_array_36_47_imag <= _zz_2569_;
      end
      if(_zz_2551_)begin
        int_reg_array_36_48_imag <= _zz_2569_;
      end
      if(_zz_2552_)begin
        int_reg_array_36_49_imag <= _zz_2569_;
      end
      if(_zz_2553_)begin
        int_reg_array_36_50_imag <= _zz_2569_;
      end
      if(_zz_2554_)begin
        int_reg_array_36_51_imag <= _zz_2569_;
      end
      if(_zz_2555_)begin
        int_reg_array_36_52_imag <= _zz_2569_;
      end
      if(_zz_2556_)begin
        int_reg_array_36_53_imag <= _zz_2569_;
      end
      if(_zz_2557_)begin
        int_reg_array_36_54_imag <= _zz_2569_;
      end
      if(_zz_2558_)begin
        int_reg_array_36_55_imag <= _zz_2569_;
      end
      if(_zz_2559_)begin
        int_reg_array_36_56_imag <= _zz_2569_;
      end
      if(_zz_2560_)begin
        int_reg_array_36_57_imag <= _zz_2569_;
      end
      if(_zz_2561_)begin
        int_reg_array_36_58_imag <= _zz_2569_;
      end
      if(_zz_2562_)begin
        int_reg_array_36_59_imag <= _zz_2569_;
      end
      if(_zz_2563_)begin
        int_reg_array_36_60_imag <= _zz_2569_;
      end
      if(_zz_2564_)begin
        int_reg_array_36_61_imag <= _zz_2569_;
      end
      if(_zz_2565_)begin
        int_reg_array_36_62_imag <= _zz_2569_;
      end
      if(_zz_2566_)begin
        int_reg_array_36_63_imag <= _zz_2569_;
      end
      if(_zz_2572_)begin
        int_reg_array_37_0_real <= _zz_2637_;
      end
      if(_zz_2573_)begin
        int_reg_array_37_1_real <= _zz_2637_;
      end
      if(_zz_2574_)begin
        int_reg_array_37_2_real <= _zz_2637_;
      end
      if(_zz_2575_)begin
        int_reg_array_37_3_real <= _zz_2637_;
      end
      if(_zz_2576_)begin
        int_reg_array_37_4_real <= _zz_2637_;
      end
      if(_zz_2577_)begin
        int_reg_array_37_5_real <= _zz_2637_;
      end
      if(_zz_2578_)begin
        int_reg_array_37_6_real <= _zz_2637_;
      end
      if(_zz_2579_)begin
        int_reg_array_37_7_real <= _zz_2637_;
      end
      if(_zz_2580_)begin
        int_reg_array_37_8_real <= _zz_2637_;
      end
      if(_zz_2581_)begin
        int_reg_array_37_9_real <= _zz_2637_;
      end
      if(_zz_2582_)begin
        int_reg_array_37_10_real <= _zz_2637_;
      end
      if(_zz_2583_)begin
        int_reg_array_37_11_real <= _zz_2637_;
      end
      if(_zz_2584_)begin
        int_reg_array_37_12_real <= _zz_2637_;
      end
      if(_zz_2585_)begin
        int_reg_array_37_13_real <= _zz_2637_;
      end
      if(_zz_2586_)begin
        int_reg_array_37_14_real <= _zz_2637_;
      end
      if(_zz_2587_)begin
        int_reg_array_37_15_real <= _zz_2637_;
      end
      if(_zz_2588_)begin
        int_reg_array_37_16_real <= _zz_2637_;
      end
      if(_zz_2589_)begin
        int_reg_array_37_17_real <= _zz_2637_;
      end
      if(_zz_2590_)begin
        int_reg_array_37_18_real <= _zz_2637_;
      end
      if(_zz_2591_)begin
        int_reg_array_37_19_real <= _zz_2637_;
      end
      if(_zz_2592_)begin
        int_reg_array_37_20_real <= _zz_2637_;
      end
      if(_zz_2593_)begin
        int_reg_array_37_21_real <= _zz_2637_;
      end
      if(_zz_2594_)begin
        int_reg_array_37_22_real <= _zz_2637_;
      end
      if(_zz_2595_)begin
        int_reg_array_37_23_real <= _zz_2637_;
      end
      if(_zz_2596_)begin
        int_reg_array_37_24_real <= _zz_2637_;
      end
      if(_zz_2597_)begin
        int_reg_array_37_25_real <= _zz_2637_;
      end
      if(_zz_2598_)begin
        int_reg_array_37_26_real <= _zz_2637_;
      end
      if(_zz_2599_)begin
        int_reg_array_37_27_real <= _zz_2637_;
      end
      if(_zz_2600_)begin
        int_reg_array_37_28_real <= _zz_2637_;
      end
      if(_zz_2601_)begin
        int_reg_array_37_29_real <= _zz_2637_;
      end
      if(_zz_2602_)begin
        int_reg_array_37_30_real <= _zz_2637_;
      end
      if(_zz_2603_)begin
        int_reg_array_37_31_real <= _zz_2637_;
      end
      if(_zz_2604_)begin
        int_reg_array_37_32_real <= _zz_2637_;
      end
      if(_zz_2605_)begin
        int_reg_array_37_33_real <= _zz_2637_;
      end
      if(_zz_2606_)begin
        int_reg_array_37_34_real <= _zz_2637_;
      end
      if(_zz_2607_)begin
        int_reg_array_37_35_real <= _zz_2637_;
      end
      if(_zz_2608_)begin
        int_reg_array_37_36_real <= _zz_2637_;
      end
      if(_zz_2609_)begin
        int_reg_array_37_37_real <= _zz_2637_;
      end
      if(_zz_2610_)begin
        int_reg_array_37_38_real <= _zz_2637_;
      end
      if(_zz_2611_)begin
        int_reg_array_37_39_real <= _zz_2637_;
      end
      if(_zz_2612_)begin
        int_reg_array_37_40_real <= _zz_2637_;
      end
      if(_zz_2613_)begin
        int_reg_array_37_41_real <= _zz_2637_;
      end
      if(_zz_2614_)begin
        int_reg_array_37_42_real <= _zz_2637_;
      end
      if(_zz_2615_)begin
        int_reg_array_37_43_real <= _zz_2637_;
      end
      if(_zz_2616_)begin
        int_reg_array_37_44_real <= _zz_2637_;
      end
      if(_zz_2617_)begin
        int_reg_array_37_45_real <= _zz_2637_;
      end
      if(_zz_2618_)begin
        int_reg_array_37_46_real <= _zz_2637_;
      end
      if(_zz_2619_)begin
        int_reg_array_37_47_real <= _zz_2637_;
      end
      if(_zz_2620_)begin
        int_reg_array_37_48_real <= _zz_2637_;
      end
      if(_zz_2621_)begin
        int_reg_array_37_49_real <= _zz_2637_;
      end
      if(_zz_2622_)begin
        int_reg_array_37_50_real <= _zz_2637_;
      end
      if(_zz_2623_)begin
        int_reg_array_37_51_real <= _zz_2637_;
      end
      if(_zz_2624_)begin
        int_reg_array_37_52_real <= _zz_2637_;
      end
      if(_zz_2625_)begin
        int_reg_array_37_53_real <= _zz_2637_;
      end
      if(_zz_2626_)begin
        int_reg_array_37_54_real <= _zz_2637_;
      end
      if(_zz_2627_)begin
        int_reg_array_37_55_real <= _zz_2637_;
      end
      if(_zz_2628_)begin
        int_reg_array_37_56_real <= _zz_2637_;
      end
      if(_zz_2629_)begin
        int_reg_array_37_57_real <= _zz_2637_;
      end
      if(_zz_2630_)begin
        int_reg_array_37_58_real <= _zz_2637_;
      end
      if(_zz_2631_)begin
        int_reg_array_37_59_real <= _zz_2637_;
      end
      if(_zz_2632_)begin
        int_reg_array_37_60_real <= _zz_2637_;
      end
      if(_zz_2633_)begin
        int_reg_array_37_61_real <= _zz_2637_;
      end
      if(_zz_2634_)begin
        int_reg_array_37_62_real <= _zz_2637_;
      end
      if(_zz_2635_)begin
        int_reg_array_37_63_real <= _zz_2637_;
      end
      if(_zz_2572_)begin
        int_reg_array_37_0_imag <= _zz_2638_;
      end
      if(_zz_2573_)begin
        int_reg_array_37_1_imag <= _zz_2638_;
      end
      if(_zz_2574_)begin
        int_reg_array_37_2_imag <= _zz_2638_;
      end
      if(_zz_2575_)begin
        int_reg_array_37_3_imag <= _zz_2638_;
      end
      if(_zz_2576_)begin
        int_reg_array_37_4_imag <= _zz_2638_;
      end
      if(_zz_2577_)begin
        int_reg_array_37_5_imag <= _zz_2638_;
      end
      if(_zz_2578_)begin
        int_reg_array_37_6_imag <= _zz_2638_;
      end
      if(_zz_2579_)begin
        int_reg_array_37_7_imag <= _zz_2638_;
      end
      if(_zz_2580_)begin
        int_reg_array_37_8_imag <= _zz_2638_;
      end
      if(_zz_2581_)begin
        int_reg_array_37_9_imag <= _zz_2638_;
      end
      if(_zz_2582_)begin
        int_reg_array_37_10_imag <= _zz_2638_;
      end
      if(_zz_2583_)begin
        int_reg_array_37_11_imag <= _zz_2638_;
      end
      if(_zz_2584_)begin
        int_reg_array_37_12_imag <= _zz_2638_;
      end
      if(_zz_2585_)begin
        int_reg_array_37_13_imag <= _zz_2638_;
      end
      if(_zz_2586_)begin
        int_reg_array_37_14_imag <= _zz_2638_;
      end
      if(_zz_2587_)begin
        int_reg_array_37_15_imag <= _zz_2638_;
      end
      if(_zz_2588_)begin
        int_reg_array_37_16_imag <= _zz_2638_;
      end
      if(_zz_2589_)begin
        int_reg_array_37_17_imag <= _zz_2638_;
      end
      if(_zz_2590_)begin
        int_reg_array_37_18_imag <= _zz_2638_;
      end
      if(_zz_2591_)begin
        int_reg_array_37_19_imag <= _zz_2638_;
      end
      if(_zz_2592_)begin
        int_reg_array_37_20_imag <= _zz_2638_;
      end
      if(_zz_2593_)begin
        int_reg_array_37_21_imag <= _zz_2638_;
      end
      if(_zz_2594_)begin
        int_reg_array_37_22_imag <= _zz_2638_;
      end
      if(_zz_2595_)begin
        int_reg_array_37_23_imag <= _zz_2638_;
      end
      if(_zz_2596_)begin
        int_reg_array_37_24_imag <= _zz_2638_;
      end
      if(_zz_2597_)begin
        int_reg_array_37_25_imag <= _zz_2638_;
      end
      if(_zz_2598_)begin
        int_reg_array_37_26_imag <= _zz_2638_;
      end
      if(_zz_2599_)begin
        int_reg_array_37_27_imag <= _zz_2638_;
      end
      if(_zz_2600_)begin
        int_reg_array_37_28_imag <= _zz_2638_;
      end
      if(_zz_2601_)begin
        int_reg_array_37_29_imag <= _zz_2638_;
      end
      if(_zz_2602_)begin
        int_reg_array_37_30_imag <= _zz_2638_;
      end
      if(_zz_2603_)begin
        int_reg_array_37_31_imag <= _zz_2638_;
      end
      if(_zz_2604_)begin
        int_reg_array_37_32_imag <= _zz_2638_;
      end
      if(_zz_2605_)begin
        int_reg_array_37_33_imag <= _zz_2638_;
      end
      if(_zz_2606_)begin
        int_reg_array_37_34_imag <= _zz_2638_;
      end
      if(_zz_2607_)begin
        int_reg_array_37_35_imag <= _zz_2638_;
      end
      if(_zz_2608_)begin
        int_reg_array_37_36_imag <= _zz_2638_;
      end
      if(_zz_2609_)begin
        int_reg_array_37_37_imag <= _zz_2638_;
      end
      if(_zz_2610_)begin
        int_reg_array_37_38_imag <= _zz_2638_;
      end
      if(_zz_2611_)begin
        int_reg_array_37_39_imag <= _zz_2638_;
      end
      if(_zz_2612_)begin
        int_reg_array_37_40_imag <= _zz_2638_;
      end
      if(_zz_2613_)begin
        int_reg_array_37_41_imag <= _zz_2638_;
      end
      if(_zz_2614_)begin
        int_reg_array_37_42_imag <= _zz_2638_;
      end
      if(_zz_2615_)begin
        int_reg_array_37_43_imag <= _zz_2638_;
      end
      if(_zz_2616_)begin
        int_reg_array_37_44_imag <= _zz_2638_;
      end
      if(_zz_2617_)begin
        int_reg_array_37_45_imag <= _zz_2638_;
      end
      if(_zz_2618_)begin
        int_reg_array_37_46_imag <= _zz_2638_;
      end
      if(_zz_2619_)begin
        int_reg_array_37_47_imag <= _zz_2638_;
      end
      if(_zz_2620_)begin
        int_reg_array_37_48_imag <= _zz_2638_;
      end
      if(_zz_2621_)begin
        int_reg_array_37_49_imag <= _zz_2638_;
      end
      if(_zz_2622_)begin
        int_reg_array_37_50_imag <= _zz_2638_;
      end
      if(_zz_2623_)begin
        int_reg_array_37_51_imag <= _zz_2638_;
      end
      if(_zz_2624_)begin
        int_reg_array_37_52_imag <= _zz_2638_;
      end
      if(_zz_2625_)begin
        int_reg_array_37_53_imag <= _zz_2638_;
      end
      if(_zz_2626_)begin
        int_reg_array_37_54_imag <= _zz_2638_;
      end
      if(_zz_2627_)begin
        int_reg_array_37_55_imag <= _zz_2638_;
      end
      if(_zz_2628_)begin
        int_reg_array_37_56_imag <= _zz_2638_;
      end
      if(_zz_2629_)begin
        int_reg_array_37_57_imag <= _zz_2638_;
      end
      if(_zz_2630_)begin
        int_reg_array_37_58_imag <= _zz_2638_;
      end
      if(_zz_2631_)begin
        int_reg_array_37_59_imag <= _zz_2638_;
      end
      if(_zz_2632_)begin
        int_reg_array_37_60_imag <= _zz_2638_;
      end
      if(_zz_2633_)begin
        int_reg_array_37_61_imag <= _zz_2638_;
      end
      if(_zz_2634_)begin
        int_reg_array_37_62_imag <= _zz_2638_;
      end
      if(_zz_2635_)begin
        int_reg_array_37_63_imag <= _zz_2638_;
      end
      if(_zz_2641_)begin
        int_reg_array_38_0_real <= _zz_2706_;
      end
      if(_zz_2642_)begin
        int_reg_array_38_1_real <= _zz_2706_;
      end
      if(_zz_2643_)begin
        int_reg_array_38_2_real <= _zz_2706_;
      end
      if(_zz_2644_)begin
        int_reg_array_38_3_real <= _zz_2706_;
      end
      if(_zz_2645_)begin
        int_reg_array_38_4_real <= _zz_2706_;
      end
      if(_zz_2646_)begin
        int_reg_array_38_5_real <= _zz_2706_;
      end
      if(_zz_2647_)begin
        int_reg_array_38_6_real <= _zz_2706_;
      end
      if(_zz_2648_)begin
        int_reg_array_38_7_real <= _zz_2706_;
      end
      if(_zz_2649_)begin
        int_reg_array_38_8_real <= _zz_2706_;
      end
      if(_zz_2650_)begin
        int_reg_array_38_9_real <= _zz_2706_;
      end
      if(_zz_2651_)begin
        int_reg_array_38_10_real <= _zz_2706_;
      end
      if(_zz_2652_)begin
        int_reg_array_38_11_real <= _zz_2706_;
      end
      if(_zz_2653_)begin
        int_reg_array_38_12_real <= _zz_2706_;
      end
      if(_zz_2654_)begin
        int_reg_array_38_13_real <= _zz_2706_;
      end
      if(_zz_2655_)begin
        int_reg_array_38_14_real <= _zz_2706_;
      end
      if(_zz_2656_)begin
        int_reg_array_38_15_real <= _zz_2706_;
      end
      if(_zz_2657_)begin
        int_reg_array_38_16_real <= _zz_2706_;
      end
      if(_zz_2658_)begin
        int_reg_array_38_17_real <= _zz_2706_;
      end
      if(_zz_2659_)begin
        int_reg_array_38_18_real <= _zz_2706_;
      end
      if(_zz_2660_)begin
        int_reg_array_38_19_real <= _zz_2706_;
      end
      if(_zz_2661_)begin
        int_reg_array_38_20_real <= _zz_2706_;
      end
      if(_zz_2662_)begin
        int_reg_array_38_21_real <= _zz_2706_;
      end
      if(_zz_2663_)begin
        int_reg_array_38_22_real <= _zz_2706_;
      end
      if(_zz_2664_)begin
        int_reg_array_38_23_real <= _zz_2706_;
      end
      if(_zz_2665_)begin
        int_reg_array_38_24_real <= _zz_2706_;
      end
      if(_zz_2666_)begin
        int_reg_array_38_25_real <= _zz_2706_;
      end
      if(_zz_2667_)begin
        int_reg_array_38_26_real <= _zz_2706_;
      end
      if(_zz_2668_)begin
        int_reg_array_38_27_real <= _zz_2706_;
      end
      if(_zz_2669_)begin
        int_reg_array_38_28_real <= _zz_2706_;
      end
      if(_zz_2670_)begin
        int_reg_array_38_29_real <= _zz_2706_;
      end
      if(_zz_2671_)begin
        int_reg_array_38_30_real <= _zz_2706_;
      end
      if(_zz_2672_)begin
        int_reg_array_38_31_real <= _zz_2706_;
      end
      if(_zz_2673_)begin
        int_reg_array_38_32_real <= _zz_2706_;
      end
      if(_zz_2674_)begin
        int_reg_array_38_33_real <= _zz_2706_;
      end
      if(_zz_2675_)begin
        int_reg_array_38_34_real <= _zz_2706_;
      end
      if(_zz_2676_)begin
        int_reg_array_38_35_real <= _zz_2706_;
      end
      if(_zz_2677_)begin
        int_reg_array_38_36_real <= _zz_2706_;
      end
      if(_zz_2678_)begin
        int_reg_array_38_37_real <= _zz_2706_;
      end
      if(_zz_2679_)begin
        int_reg_array_38_38_real <= _zz_2706_;
      end
      if(_zz_2680_)begin
        int_reg_array_38_39_real <= _zz_2706_;
      end
      if(_zz_2681_)begin
        int_reg_array_38_40_real <= _zz_2706_;
      end
      if(_zz_2682_)begin
        int_reg_array_38_41_real <= _zz_2706_;
      end
      if(_zz_2683_)begin
        int_reg_array_38_42_real <= _zz_2706_;
      end
      if(_zz_2684_)begin
        int_reg_array_38_43_real <= _zz_2706_;
      end
      if(_zz_2685_)begin
        int_reg_array_38_44_real <= _zz_2706_;
      end
      if(_zz_2686_)begin
        int_reg_array_38_45_real <= _zz_2706_;
      end
      if(_zz_2687_)begin
        int_reg_array_38_46_real <= _zz_2706_;
      end
      if(_zz_2688_)begin
        int_reg_array_38_47_real <= _zz_2706_;
      end
      if(_zz_2689_)begin
        int_reg_array_38_48_real <= _zz_2706_;
      end
      if(_zz_2690_)begin
        int_reg_array_38_49_real <= _zz_2706_;
      end
      if(_zz_2691_)begin
        int_reg_array_38_50_real <= _zz_2706_;
      end
      if(_zz_2692_)begin
        int_reg_array_38_51_real <= _zz_2706_;
      end
      if(_zz_2693_)begin
        int_reg_array_38_52_real <= _zz_2706_;
      end
      if(_zz_2694_)begin
        int_reg_array_38_53_real <= _zz_2706_;
      end
      if(_zz_2695_)begin
        int_reg_array_38_54_real <= _zz_2706_;
      end
      if(_zz_2696_)begin
        int_reg_array_38_55_real <= _zz_2706_;
      end
      if(_zz_2697_)begin
        int_reg_array_38_56_real <= _zz_2706_;
      end
      if(_zz_2698_)begin
        int_reg_array_38_57_real <= _zz_2706_;
      end
      if(_zz_2699_)begin
        int_reg_array_38_58_real <= _zz_2706_;
      end
      if(_zz_2700_)begin
        int_reg_array_38_59_real <= _zz_2706_;
      end
      if(_zz_2701_)begin
        int_reg_array_38_60_real <= _zz_2706_;
      end
      if(_zz_2702_)begin
        int_reg_array_38_61_real <= _zz_2706_;
      end
      if(_zz_2703_)begin
        int_reg_array_38_62_real <= _zz_2706_;
      end
      if(_zz_2704_)begin
        int_reg_array_38_63_real <= _zz_2706_;
      end
      if(_zz_2641_)begin
        int_reg_array_38_0_imag <= _zz_2707_;
      end
      if(_zz_2642_)begin
        int_reg_array_38_1_imag <= _zz_2707_;
      end
      if(_zz_2643_)begin
        int_reg_array_38_2_imag <= _zz_2707_;
      end
      if(_zz_2644_)begin
        int_reg_array_38_3_imag <= _zz_2707_;
      end
      if(_zz_2645_)begin
        int_reg_array_38_4_imag <= _zz_2707_;
      end
      if(_zz_2646_)begin
        int_reg_array_38_5_imag <= _zz_2707_;
      end
      if(_zz_2647_)begin
        int_reg_array_38_6_imag <= _zz_2707_;
      end
      if(_zz_2648_)begin
        int_reg_array_38_7_imag <= _zz_2707_;
      end
      if(_zz_2649_)begin
        int_reg_array_38_8_imag <= _zz_2707_;
      end
      if(_zz_2650_)begin
        int_reg_array_38_9_imag <= _zz_2707_;
      end
      if(_zz_2651_)begin
        int_reg_array_38_10_imag <= _zz_2707_;
      end
      if(_zz_2652_)begin
        int_reg_array_38_11_imag <= _zz_2707_;
      end
      if(_zz_2653_)begin
        int_reg_array_38_12_imag <= _zz_2707_;
      end
      if(_zz_2654_)begin
        int_reg_array_38_13_imag <= _zz_2707_;
      end
      if(_zz_2655_)begin
        int_reg_array_38_14_imag <= _zz_2707_;
      end
      if(_zz_2656_)begin
        int_reg_array_38_15_imag <= _zz_2707_;
      end
      if(_zz_2657_)begin
        int_reg_array_38_16_imag <= _zz_2707_;
      end
      if(_zz_2658_)begin
        int_reg_array_38_17_imag <= _zz_2707_;
      end
      if(_zz_2659_)begin
        int_reg_array_38_18_imag <= _zz_2707_;
      end
      if(_zz_2660_)begin
        int_reg_array_38_19_imag <= _zz_2707_;
      end
      if(_zz_2661_)begin
        int_reg_array_38_20_imag <= _zz_2707_;
      end
      if(_zz_2662_)begin
        int_reg_array_38_21_imag <= _zz_2707_;
      end
      if(_zz_2663_)begin
        int_reg_array_38_22_imag <= _zz_2707_;
      end
      if(_zz_2664_)begin
        int_reg_array_38_23_imag <= _zz_2707_;
      end
      if(_zz_2665_)begin
        int_reg_array_38_24_imag <= _zz_2707_;
      end
      if(_zz_2666_)begin
        int_reg_array_38_25_imag <= _zz_2707_;
      end
      if(_zz_2667_)begin
        int_reg_array_38_26_imag <= _zz_2707_;
      end
      if(_zz_2668_)begin
        int_reg_array_38_27_imag <= _zz_2707_;
      end
      if(_zz_2669_)begin
        int_reg_array_38_28_imag <= _zz_2707_;
      end
      if(_zz_2670_)begin
        int_reg_array_38_29_imag <= _zz_2707_;
      end
      if(_zz_2671_)begin
        int_reg_array_38_30_imag <= _zz_2707_;
      end
      if(_zz_2672_)begin
        int_reg_array_38_31_imag <= _zz_2707_;
      end
      if(_zz_2673_)begin
        int_reg_array_38_32_imag <= _zz_2707_;
      end
      if(_zz_2674_)begin
        int_reg_array_38_33_imag <= _zz_2707_;
      end
      if(_zz_2675_)begin
        int_reg_array_38_34_imag <= _zz_2707_;
      end
      if(_zz_2676_)begin
        int_reg_array_38_35_imag <= _zz_2707_;
      end
      if(_zz_2677_)begin
        int_reg_array_38_36_imag <= _zz_2707_;
      end
      if(_zz_2678_)begin
        int_reg_array_38_37_imag <= _zz_2707_;
      end
      if(_zz_2679_)begin
        int_reg_array_38_38_imag <= _zz_2707_;
      end
      if(_zz_2680_)begin
        int_reg_array_38_39_imag <= _zz_2707_;
      end
      if(_zz_2681_)begin
        int_reg_array_38_40_imag <= _zz_2707_;
      end
      if(_zz_2682_)begin
        int_reg_array_38_41_imag <= _zz_2707_;
      end
      if(_zz_2683_)begin
        int_reg_array_38_42_imag <= _zz_2707_;
      end
      if(_zz_2684_)begin
        int_reg_array_38_43_imag <= _zz_2707_;
      end
      if(_zz_2685_)begin
        int_reg_array_38_44_imag <= _zz_2707_;
      end
      if(_zz_2686_)begin
        int_reg_array_38_45_imag <= _zz_2707_;
      end
      if(_zz_2687_)begin
        int_reg_array_38_46_imag <= _zz_2707_;
      end
      if(_zz_2688_)begin
        int_reg_array_38_47_imag <= _zz_2707_;
      end
      if(_zz_2689_)begin
        int_reg_array_38_48_imag <= _zz_2707_;
      end
      if(_zz_2690_)begin
        int_reg_array_38_49_imag <= _zz_2707_;
      end
      if(_zz_2691_)begin
        int_reg_array_38_50_imag <= _zz_2707_;
      end
      if(_zz_2692_)begin
        int_reg_array_38_51_imag <= _zz_2707_;
      end
      if(_zz_2693_)begin
        int_reg_array_38_52_imag <= _zz_2707_;
      end
      if(_zz_2694_)begin
        int_reg_array_38_53_imag <= _zz_2707_;
      end
      if(_zz_2695_)begin
        int_reg_array_38_54_imag <= _zz_2707_;
      end
      if(_zz_2696_)begin
        int_reg_array_38_55_imag <= _zz_2707_;
      end
      if(_zz_2697_)begin
        int_reg_array_38_56_imag <= _zz_2707_;
      end
      if(_zz_2698_)begin
        int_reg_array_38_57_imag <= _zz_2707_;
      end
      if(_zz_2699_)begin
        int_reg_array_38_58_imag <= _zz_2707_;
      end
      if(_zz_2700_)begin
        int_reg_array_38_59_imag <= _zz_2707_;
      end
      if(_zz_2701_)begin
        int_reg_array_38_60_imag <= _zz_2707_;
      end
      if(_zz_2702_)begin
        int_reg_array_38_61_imag <= _zz_2707_;
      end
      if(_zz_2703_)begin
        int_reg_array_38_62_imag <= _zz_2707_;
      end
      if(_zz_2704_)begin
        int_reg_array_38_63_imag <= _zz_2707_;
      end
      if(_zz_2710_)begin
        int_reg_array_39_0_real <= _zz_2775_;
      end
      if(_zz_2711_)begin
        int_reg_array_39_1_real <= _zz_2775_;
      end
      if(_zz_2712_)begin
        int_reg_array_39_2_real <= _zz_2775_;
      end
      if(_zz_2713_)begin
        int_reg_array_39_3_real <= _zz_2775_;
      end
      if(_zz_2714_)begin
        int_reg_array_39_4_real <= _zz_2775_;
      end
      if(_zz_2715_)begin
        int_reg_array_39_5_real <= _zz_2775_;
      end
      if(_zz_2716_)begin
        int_reg_array_39_6_real <= _zz_2775_;
      end
      if(_zz_2717_)begin
        int_reg_array_39_7_real <= _zz_2775_;
      end
      if(_zz_2718_)begin
        int_reg_array_39_8_real <= _zz_2775_;
      end
      if(_zz_2719_)begin
        int_reg_array_39_9_real <= _zz_2775_;
      end
      if(_zz_2720_)begin
        int_reg_array_39_10_real <= _zz_2775_;
      end
      if(_zz_2721_)begin
        int_reg_array_39_11_real <= _zz_2775_;
      end
      if(_zz_2722_)begin
        int_reg_array_39_12_real <= _zz_2775_;
      end
      if(_zz_2723_)begin
        int_reg_array_39_13_real <= _zz_2775_;
      end
      if(_zz_2724_)begin
        int_reg_array_39_14_real <= _zz_2775_;
      end
      if(_zz_2725_)begin
        int_reg_array_39_15_real <= _zz_2775_;
      end
      if(_zz_2726_)begin
        int_reg_array_39_16_real <= _zz_2775_;
      end
      if(_zz_2727_)begin
        int_reg_array_39_17_real <= _zz_2775_;
      end
      if(_zz_2728_)begin
        int_reg_array_39_18_real <= _zz_2775_;
      end
      if(_zz_2729_)begin
        int_reg_array_39_19_real <= _zz_2775_;
      end
      if(_zz_2730_)begin
        int_reg_array_39_20_real <= _zz_2775_;
      end
      if(_zz_2731_)begin
        int_reg_array_39_21_real <= _zz_2775_;
      end
      if(_zz_2732_)begin
        int_reg_array_39_22_real <= _zz_2775_;
      end
      if(_zz_2733_)begin
        int_reg_array_39_23_real <= _zz_2775_;
      end
      if(_zz_2734_)begin
        int_reg_array_39_24_real <= _zz_2775_;
      end
      if(_zz_2735_)begin
        int_reg_array_39_25_real <= _zz_2775_;
      end
      if(_zz_2736_)begin
        int_reg_array_39_26_real <= _zz_2775_;
      end
      if(_zz_2737_)begin
        int_reg_array_39_27_real <= _zz_2775_;
      end
      if(_zz_2738_)begin
        int_reg_array_39_28_real <= _zz_2775_;
      end
      if(_zz_2739_)begin
        int_reg_array_39_29_real <= _zz_2775_;
      end
      if(_zz_2740_)begin
        int_reg_array_39_30_real <= _zz_2775_;
      end
      if(_zz_2741_)begin
        int_reg_array_39_31_real <= _zz_2775_;
      end
      if(_zz_2742_)begin
        int_reg_array_39_32_real <= _zz_2775_;
      end
      if(_zz_2743_)begin
        int_reg_array_39_33_real <= _zz_2775_;
      end
      if(_zz_2744_)begin
        int_reg_array_39_34_real <= _zz_2775_;
      end
      if(_zz_2745_)begin
        int_reg_array_39_35_real <= _zz_2775_;
      end
      if(_zz_2746_)begin
        int_reg_array_39_36_real <= _zz_2775_;
      end
      if(_zz_2747_)begin
        int_reg_array_39_37_real <= _zz_2775_;
      end
      if(_zz_2748_)begin
        int_reg_array_39_38_real <= _zz_2775_;
      end
      if(_zz_2749_)begin
        int_reg_array_39_39_real <= _zz_2775_;
      end
      if(_zz_2750_)begin
        int_reg_array_39_40_real <= _zz_2775_;
      end
      if(_zz_2751_)begin
        int_reg_array_39_41_real <= _zz_2775_;
      end
      if(_zz_2752_)begin
        int_reg_array_39_42_real <= _zz_2775_;
      end
      if(_zz_2753_)begin
        int_reg_array_39_43_real <= _zz_2775_;
      end
      if(_zz_2754_)begin
        int_reg_array_39_44_real <= _zz_2775_;
      end
      if(_zz_2755_)begin
        int_reg_array_39_45_real <= _zz_2775_;
      end
      if(_zz_2756_)begin
        int_reg_array_39_46_real <= _zz_2775_;
      end
      if(_zz_2757_)begin
        int_reg_array_39_47_real <= _zz_2775_;
      end
      if(_zz_2758_)begin
        int_reg_array_39_48_real <= _zz_2775_;
      end
      if(_zz_2759_)begin
        int_reg_array_39_49_real <= _zz_2775_;
      end
      if(_zz_2760_)begin
        int_reg_array_39_50_real <= _zz_2775_;
      end
      if(_zz_2761_)begin
        int_reg_array_39_51_real <= _zz_2775_;
      end
      if(_zz_2762_)begin
        int_reg_array_39_52_real <= _zz_2775_;
      end
      if(_zz_2763_)begin
        int_reg_array_39_53_real <= _zz_2775_;
      end
      if(_zz_2764_)begin
        int_reg_array_39_54_real <= _zz_2775_;
      end
      if(_zz_2765_)begin
        int_reg_array_39_55_real <= _zz_2775_;
      end
      if(_zz_2766_)begin
        int_reg_array_39_56_real <= _zz_2775_;
      end
      if(_zz_2767_)begin
        int_reg_array_39_57_real <= _zz_2775_;
      end
      if(_zz_2768_)begin
        int_reg_array_39_58_real <= _zz_2775_;
      end
      if(_zz_2769_)begin
        int_reg_array_39_59_real <= _zz_2775_;
      end
      if(_zz_2770_)begin
        int_reg_array_39_60_real <= _zz_2775_;
      end
      if(_zz_2771_)begin
        int_reg_array_39_61_real <= _zz_2775_;
      end
      if(_zz_2772_)begin
        int_reg_array_39_62_real <= _zz_2775_;
      end
      if(_zz_2773_)begin
        int_reg_array_39_63_real <= _zz_2775_;
      end
      if(_zz_2710_)begin
        int_reg_array_39_0_imag <= _zz_2776_;
      end
      if(_zz_2711_)begin
        int_reg_array_39_1_imag <= _zz_2776_;
      end
      if(_zz_2712_)begin
        int_reg_array_39_2_imag <= _zz_2776_;
      end
      if(_zz_2713_)begin
        int_reg_array_39_3_imag <= _zz_2776_;
      end
      if(_zz_2714_)begin
        int_reg_array_39_4_imag <= _zz_2776_;
      end
      if(_zz_2715_)begin
        int_reg_array_39_5_imag <= _zz_2776_;
      end
      if(_zz_2716_)begin
        int_reg_array_39_6_imag <= _zz_2776_;
      end
      if(_zz_2717_)begin
        int_reg_array_39_7_imag <= _zz_2776_;
      end
      if(_zz_2718_)begin
        int_reg_array_39_8_imag <= _zz_2776_;
      end
      if(_zz_2719_)begin
        int_reg_array_39_9_imag <= _zz_2776_;
      end
      if(_zz_2720_)begin
        int_reg_array_39_10_imag <= _zz_2776_;
      end
      if(_zz_2721_)begin
        int_reg_array_39_11_imag <= _zz_2776_;
      end
      if(_zz_2722_)begin
        int_reg_array_39_12_imag <= _zz_2776_;
      end
      if(_zz_2723_)begin
        int_reg_array_39_13_imag <= _zz_2776_;
      end
      if(_zz_2724_)begin
        int_reg_array_39_14_imag <= _zz_2776_;
      end
      if(_zz_2725_)begin
        int_reg_array_39_15_imag <= _zz_2776_;
      end
      if(_zz_2726_)begin
        int_reg_array_39_16_imag <= _zz_2776_;
      end
      if(_zz_2727_)begin
        int_reg_array_39_17_imag <= _zz_2776_;
      end
      if(_zz_2728_)begin
        int_reg_array_39_18_imag <= _zz_2776_;
      end
      if(_zz_2729_)begin
        int_reg_array_39_19_imag <= _zz_2776_;
      end
      if(_zz_2730_)begin
        int_reg_array_39_20_imag <= _zz_2776_;
      end
      if(_zz_2731_)begin
        int_reg_array_39_21_imag <= _zz_2776_;
      end
      if(_zz_2732_)begin
        int_reg_array_39_22_imag <= _zz_2776_;
      end
      if(_zz_2733_)begin
        int_reg_array_39_23_imag <= _zz_2776_;
      end
      if(_zz_2734_)begin
        int_reg_array_39_24_imag <= _zz_2776_;
      end
      if(_zz_2735_)begin
        int_reg_array_39_25_imag <= _zz_2776_;
      end
      if(_zz_2736_)begin
        int_reg_array_39_26_imag <= _zz_2776_;
      end
      if(_zz_2737_)begin
        int_reg_array_39_27_imag <= _zz_2776_;
      end
      if(_zz_2738_)begin
        int_reg_array_39_28_imag <= _zz_2776_;
      end
      if(_zz_2739_)begin
        int_reg_array_39_29_imag <= _zz_2776_;
      end
      if(_zz_2740_)begin
        int_reg_array_39_30_imag <= _zz_2776_;
      end
      if(_zz_2741_)begin
        int_reg_array_39_31_imag <= _zz_2776_;
      end
      if(_zz_2742_)begin
        int_reg_array_39_32_imag <= _zz_2776_;
      end
      if(_zz_2743_)begin
        int_reg_array_39_33_imag <= _zz_2776_;
      end
      if(_zz_2744_)begin
        int_reg_array_39_34_imag <= _zz_2776_;
      end
      if(_zz_2745_)begin
        int_reg_array_39_35_imag <= _zz_2776_;
      end
      if(_zz_2746_)begin
        int_reg_array_39_36_imag <= _zz_2776_;
      end
      if(_zz_2747_)begin
        int_reg_array_39_37_imag <= _zz_2776_;
      end
      if(_zz_2748_)begin
        int_reg_array_39_38_imag <= _zz_2776_;
      end
      if(_zz_2749_)begin
        int_reg_array_39_39_imag <= _zz_2776_;
      end
      if(_zz_2750_)begin
        int_reg_array_39_40_imag <= _zz_2776_;
      end
      if(_zz_2751_)begin
        int_reg_array_39_41_imag <= _zz_2776_;
      end
      if(_zz_2752_)begin
        int_reg_array_39_42_imag <= _zz_2776_;
      end
      if(_zz_2753_)begin
        int_reg_array_39_43_imag <= _zz_2776_;
      end
      if(_zz_2754_)begin
        int_reg_array_39_44_imag <= _zz_2776_;
      end
      if(_zz_2755_)begin
        int_reg_array_39_45_imag <= _zz_2776_;
      end
      if(_zz_2756_)begin
        int_reg_array_39_46_imag <= _zz_2776_;
      end
      if(_zz_2757_)begin
        int_reg_array_39_47_imag <= _zz_2776_;
      end
      if(_zz_2758_)begin
        int_reg_array_39_48_imag <= _zz_2776_;
      end
      if(_zz_2759_)begin
        int_reg_array_39_49_imag <= _zz_2776_;
      end
      if(_zz_2760_)begin
        int_reg_array_39_50_imag <= _zz_2776_;
      end
      if(_zz_2761_)begin
        int_reg_array_39_51_imag <= _zz_2776_;
      end
      if(_zz_2762_)begin
        int_reg_array_39_52_imag <= _zz_2776_;
      end
      if(_zz_2763_)begin
        int_reg_array_39_53_imag <= _zz_2776_;
      end
      if(_zz_2764_)begin
        int_reg_array_39_54_imag <= _zz_2776_;
      end
      if(_zz_2765_)begin
        int_reg_array_39_55_imag <= _zz_2776_;
      end
      if(_zz_2766_)begin
        int_reg_array_39_56_imag <= _zz_2776_;
      end
      if(_zz_2767_)begin
        int_reg_array_39_57_imag <= _zz_2776_;
      end
      if(_zz_2768_)begin
        int_reg_array_39_58_imag <= _zz_2776_;
      end
      if(_zz_2769_)begin
        int_reg_array_39_59_imag <= _zz_2776_;
      end
      if(_zz_2770_)begin
        int_reg_array_39_60_imag <= _zz_2776_;
      end
      if(_zz_2771_)begin
        int_reg_array_39_61_imag <= _zz_2776_;
      end
      if(_zz_2772_)begin
        int_reg_array_39_62_imag <= _zz_2776_;
      end
      if(_zz_2773_)begin
        int_reg_array_39_63_imag <= _zz_2776_;
      end
      if(_zz_2779_)begin
        int_reg_array_40_0_real <= _zz_2844_;
      end
      if(_zz_2780_)begin
        int_reg_array_40_1_real <= _zz_2844_;
      end
      if(_zz_2781_)begin
        int_reg_array_40_2_real <= _zz_2844_;
      end
      if(_zz_2782_)begin
        int_reg_array_40_3_real <= _zz_2844_;
      end
      if(_zz_2783_)begin
        int_reg_array_40_4_real <= _zz_2844_;
      end
      if(_zz_2784_)begin
        int_reg_array_40_5_real <= _zz_2844_;
      end
      if(_zz_2785_)begin
        int_reg_array_40_6_real <= _zz_2844_;
      end
      if(_zz_2786_)begin
        int_reg_array_40_7_real <= _zz_2844_;
      end
      if(_zz_2787_)begin
        int_reg_array_40_8_real <= _zz_2844_;
      end
      if(_zz_2788_)begin
        int_reg_array_40_9_real <= _zz_2844_;
      end
      if(_zz_2789_)begin
        int_reg_array_40_10_real <= _zz_2844_;
      end
      if(_zz_2790_)begin
        int_reg_array_40_11_real <= _zz_2844_;
      end
      if(_zz_2791_)begin
        int_reg_array_40_12_real <= _zz_2844_;
      end
      if(_zz_2792_)begin
        int_reg_array_40_13_real <= _zz_2844_;
      end
      if(_zz_2793_)begin
        int_reg_array_40_14_real <= _zz_2844_;
      end
      if(_zz_2794_)begin
        int_reg_array_40_15_real <= _zz_2844_;
      end
      if(_zz_2795_)begin
        int_reg_array_40_16_real <= _zz_2844_;
      end
      if(_zz_2796_)begin
        int_reg_array_40_17_real <= _zz_2844_;
      end
      if(_zz_2797_)begin
        int_reg_array_40_18_real <= _zz_2844_;
      end
      if(_zz_2798_)begin
        int_reg_array_40_19_real <= _zz_2844_;
      end
      if(_zz_2799_)begin
        int_reg_array_40_20_real <= _zz_2844_;
      end
      if(_zz_2800_)begin
        int_reg_array_40_21_real <= _zz_2844_;
      end
      if(_zz_2801_)begin
        int_reg_array_40_22_real <= _zz_2844_;
      end
      if(_zz_2802_)begin
        int_reg_array_40_23_real <= _zz_2844_;
      end
      if(_zz_2803_)begin
        int_reg_array_40_24_real <= _zz_2844_;
      end
      if(_zz_2804_)begin
        int_reg_array_40_25_real <= _zz_2844_;
      end
      if(_zz_2805_)begin
        int_reg_array_40_26_real <= _zz_2844_;
      end
      if(_zz_2806_)begin
        int_reg_array_40_27_real <= _zz_2844_;
      end
      if(_zz_2807_)begin
        int_reg_array_40_28_real <= _zz_2844_;
      end
      if(_zz_2808_)begin
        int_reg_array_40_29_real <= _zz_2844_;
      end
      if(_zz_2809_)begin
        int_reg_array_40_30_real <= _zz_2844_;
      end
      if(_zz_2810_)begin
        int_reg_array_40_31_real <= _zz_2844_;
      end
      if(_zz_2811_)begin
        int_reg_array_40_32_real <= _zz_2844_;
      end
      if(_zz_2812_)begin
        int_reg_array_40_33_real <= _zz_2844_;
      end
      if(_zz_2813_)begin
        int_reg_array_40_34_real <= _zz_2844_;
      end
      if(_zz_2814_)begin
        int_reg_array_40_35_real <= _zz_2844_;
      end
      if(_zz_2815_)begin
        int_reg_array_40_36_real <= _zz_2844_;
      end
      if(_zz_2816_)begin
        int_reg_array_40_37_real <= _zz_2844_;
      end
      if(_zz_2817_)begin
        int_reg_array_40_38_real <= _zz_2844_;
      end
      if(_zz_2818_)begin
        int_reg_array_40_39_real <= _zz_2844_;
      end
      if(_zz_2819_)begin
        int_reg_array_40_40_real <= _zz_2844_;
      end
      if(_zz_2820_)begin
        int_reg_array_40_41_real <= _zz_2844_;
      end
      if(_zz_2821_)begin
        int_reg_array_40_42_real <= _zz_2844_;
      end
      if(_zz_2822_)begin
        int_reg_array_40_43_real <= _zz_2844_;
      end
      if(_zz_2823_)begin
        int_reg_array_40_44_real <= _zz_2844_;
      end
      if(_zz_2824_)begin
        int_reg_array_40_45_real <= _zz_2844_;
      end
      if(_zz_2825_)begin
        int_reg_array_40_46_real <= _zz_2844_;
      end
      if(_zz_2826_)begin
        int_reg_array_40_47_real <= _zz_2844_;
      end
      if(_zz_2827_)begin
        int_reg_array_40_48_real <= _zz_2844_;
      end
      if(_zz_2828_)begin
        int_reg_array_40_49_real <= _zz_2844_;
      end
      if(_zz_2829_)begin
        int_reg_array_40_50_real <= _zz_2844_;
      end
      if(_zz_2830_)begin
        int_reg_array_40_51_real <= _zz_2844_;
      end
      if(_zz_2831_)begin
        int_reg_array_40_52_real <= _zz_2844_;
      end
      if(_zz_2832_)begin
        int_reg_array_40_53_real <= _zz_2844_;
      end
      if(_zz_2833_)begin
        int_reg_array_40_54_real <= _zz_2844_;
      end
      if(_zz_2834_)begin
        int_reg_array_40_55_real <= _zz_2844_;
      end
      if(_zz_2835_)begin
        int_reg_array_40_56_real <= _zz_2844_;
      end
      if(_zz_2836_)begin
        int_reg_array_40_57_real <= _zz_2844_;
      end
      if(_zz_2837_)begin
        int_reg_array_40_58_real <= _zz_2844_;
      end
      if(_zz_2838_)begin
        int_reg_array_40_59_real <= _zz_2844_;
      end
      if(_zz_2839_)begin
        int_reg_array_40_60_real <= _zz_2844_;
      end
      if(_zz_2840_)begin
        int_reg_array_40_61_real <= _zz_2844_;
      end
      if(_zz_2841_)begin
        int_reg_array_40_62_real <= _zz_2844_;
      end
      if(_zz_2842_)begin
        int_reg_array_40_63_real <= _zz_2844_;
      end
      if(_zz_2779_)begin
        int_reg_array_40_0_imag <= _zz_2845_;
      end
      if(_zz_2780_)begin
        int_reg_array_40_1_imag <= _zz_2845_;
      end
      if(_zz_2781_)begin
        int_reg_array_40_2_imag <= _zz_2845_;
      end
      if(_zz_2782_)begin
        int_reg_array_40_3_imag <= _zz_2845_;
      end
      if(_zz_2783_)begin
        int_reg_array_40_4_imag <= _zz_2845_;
      end
      if(_zz_2784_)begin
        int_reg_array_40_5_imag <= _zz_2845_;
      end
      if(_zz_2785_)begin
        int_reg_array_40_6_imag <= _zz_2845_;
      end
      if(_zz_2786_)begin
        int_reg_array_40_7_imag <= _zz_2845_;
      end
      if(_zz_2787_)begin
        int_reg_array_40_8_imag <= _zz_2845_;
      end
      if(_zz_2788_)begin
        int_reg_array_40_9_imag <= _zz_2845_;
      end
      if(_zz_2789_)begin
        int_reg_array_40_10_imag <= _zz_2845_;
      end
      if(_zz_2790_)begin
        int_reg_array_40_11_imag <= _zz_2845_;
      end
      if(_zz_2791_)begin
        int_reg_array_40_12_imag <= _zz_2845_;
      end
      if(_zz_2792_)begin
        int_reg_array_40_13_imag <= _zz_2845_;
      end
      if(_zz_2793_)begin
        int_reg_array_40_14_imag <= _zz_2845_;
      end
      if(_zz_2794_)begin
        int_reg_array_40_15_imag <= _zz_2845_;
      end
      if(_zz_2795_)begin
        int_reg_array_40_16_imag <= _zz_2845_;
      end
      if(_zz_2796_)begin
        int_reg_array_40_17_imag <= _zz_2845_;
      end
      if(_zz_2797_)begin
        int_reg_array_40_18_imag <= _zz_2845_;
      end
      if(_zz_2798_)begin
        int_reg_array_40_19_imag <= _zz_2845_;
      end
      if(_zz_2799_)begin
        int_reg_array_40_20_imag <= _zz_2845_;
      end
      if(_zz_2800_)begin
        int_reg_array_40_21_imag <= _zz_2845_;
      end
      if(_zz_2801_)begin
        int_reg_array_40_22_imag <= _zz_2845_;
      end
      if(_zz_2802_)begin
        int_reg_array_40_23_imag <= _zz_2845_;
      end
      if(_zz_2803_)begin
        int_reg_array_40_24_imag <= _zz_2845_;
      end
      if(_zz_2804_)begin
        int_reg_array_40_25_imag <= _zz_2845_;
      end
      if(_zz_2805_)begin
        int_reg_array_40_26_imag <= _zz_2845_;
      end
      if(_zz_2806_)begin
        int_reg_array_40_27_imag <= _zz_2845_;
      end
      if(_zz_2807_)begin
        int_reg_array_40_28_imag <= _zz_2845_;
      end
      if(_zz_2808_)begin
        int_reg_array_40_29_imag <= _zz_2845_;
      end
      if(_zz_2809_)begin
        int_reg_array_40_30_imag <= _zz_2845_;
      end
      if(_zz_2810_)begin
        int_reg_array_40_31_imag <= _zz_2845_;
      end
      if(_zz_2811_)begin
        int_reg_array_40_32_imag <= _zz_2845_;
      end
      if(_zz_2812_)begin
        int_reg_array_40_33_imag <= _zz_2845_;
      end
      if(_zz_2813_)begin
        int_reg_array_40_34_imag <= _zz_2845_;
      end
      if(_zz_2814_)begin
        int_reg_array_40_35_imag <= _zz_2845_;
      end
      if(_zz_2815_)begin
        int_reg_array_40_36_imag <= _zz_2845_;
      end
      if(_zz_2816_)begin
        int_reg_array_40_37_imag <= _zz_2845_;
      end
      if(_zz_2817_)begin
        int_reg_array_40_38_imag <= _zz_2845_;
      end
      if(_zz_2818_)begin
        int_reg_array_40_39_imag <= _zz_2845_;
      end
      if(_zz_2819_)begin
        int_reg_array_40_40_imag <= _zz_2845_;
      end
      if(_zz_2820_)begin
        int_reg_array_40_41_imag <= _zz_2845_;
      end
      if(_zz_2821_)begin
        int_reg_array_40_42_imag <= _zz_2845_;
      end
      if(_zz_2822_)begin
        int_reg_array_40_43_imag <= _zz_2845_;
      end
      if(_zz_2823_)begin
        int_reg_array_40_44_imag <= _zz_2845_;
      end
      if(_zz_2824_)begin
        int_reg_array_40_45_imag <= _zz_2845_;
      end
      if(_zz_2825_)begin
        int_reg_array_40_46_imag <= _zz_2845_;
      end
      if(_zz_2826_)begin
        int_reg_array_40_47_imag <= _zz_2845_;
      end
      if(_zz_2827_)begin
        int_reg_array_40_48_imag <= _zz_2845_;
      end
      if(_zz_2828_)begin
        int_reg_array_40_49_imag <= _zz_2845_;
      end
      if(_zz_2829_)begin
        int_reg_array_40_50_imag <= _zz_2845_;
      end
      if(_zz_2830_)begin
        int_reg_array_40_51_imag <= _zz_2845_;
      end
      if(_zz_2831_)begin
        int_reg_array_40_52_imag <= _zz_2845_;
      end
      if(_zz_2832_)begin
        int_reg_array_40_53_imag <= _zz_2845_;
      end
      if(_zz_2833_)begin
        int_reg_array_40_54_imag <= _zz_2845_;
      end
      if(_zz_2834_)begin
        int_reg_array_40_55_imag <= _zz_2845_;
      end
      if(_zz_2835_)begin
        int_reg_array_40_56_imag <= _zz_2845_;
      end
      if(_zz_2836_)begin
        int_reg_array_40_57_imag <= _zz_2845_;
      end
      if(_zz_2837_)begin
        int_reg_array_40_58_imag <= _zz_2845_;
      end
      if(_zz_2838_)begin
        int_reg_array_40_59_imag <= _zz_2845_;
      end
      if(_zz_2839_)begin
        int_reg_array_40_60_imag <= _zz_2845_;
      end
      if(_zz_2840_)begin
        int_reg_array_40_61_imag <= _zz_2845_;
      end
      if(_zz_2841_)begin
        int_reg_array_40_62_imag <= _zz_2845_;
      end
      if(_zz_2842_)begin
        int_reg_array_40_63_imag <= _zz_2845_;
      end
      if(_zz_2848_)begin
        int_reg_array_41_0_real <= _zz_2913_;
      end
      if(_zz_2849_)begin
        int_reg_array_41_1_real <= _zz_2913_;
      end
      if(_zz_2850_)begin
        int_reg_array_41_2_real <= _zz_2913_;
      end
      if(_zz_2851_)begin
        int_reg_array_41_3_real <= _zz_2913_;
      end
      if(_zz_2852_)begin
        int_reg_array_41_4_real <= _zz_2913_;
      end
      if(_zz_2853_)begin
        int_reg_array_41_5_real <= _zz_2913_;
      end
      if(_zz_2854_)begin
        int_reg_array_41_6_real <= _zz_2913_;
      end
      if(_zz_2855_)begin
        int_reg_array_41_7_real <= _zz_2913_;
      end
      if(_zz_2856_)begin
        int_reg_array_41_8_real <= _zz_2913_;
      end
      if(_zz_2857_)begin
        int_reg_array_41_9_real <= _zz_2913_;
      end
      if(_zz_2858_)begin
        int_reg_array_41_10_real <= _zz_2913_;
      end
      if(_zz_2859_)begin
        int_reg_array_41_11_real <= _zz_2913_;
      end
      if(_zz_2860_)begin
        int_reg_array_41_12_real <= _zz_2913_;
      end
      if(_zz_2861_)begin
        int_reg_array_41_13_real <= _zz_2913_;
      end
      if(_zz_2862_)begin
        int_reg_array_41_14_real <= _zz_2913_;
      end
      if(_zz_2863_)begin
        int_reg_array_41_15_real <= _zz_2913_;
      end
      if(_zz_2864_)begin
        int_reg_array_41_16_real <= _zz_2913_;
      end
      if(_zz_2865_)begin
        int_reg_array_41_17_real <= _zz_2913_;
      end
      if(_zz_2866_)begin
        int_reg_array_41_18_real <= _zz_2913_;
      end
      if(_zz_2867_)begin
        int_reg_array_41_19_real <= _zz_2913_;
      end
      if(_zz_2868_)begin
        int_reg_array_41_20_real <= _zz_2913_;
      end
      if(_zz_2869_)begin
        int_reg_array_41_21_real <= _zz_2913_;
      end
      if(_zz_2870_)begin
        int_reg_array_41_22_real <= _zz_2913_;
      end
      if(_zz_2871_)begin
        int_reg_array_41_23_real <= _zz_2913_;
      end
      if(_zz_2872_)begin
        int_reg_array_41_24_real <= _zz_2913_;
      end
      if(_zz_2873_)begin
        int_reg_array_41_25_real <= _zz_2913_;
      end
      if(_zz_2874_)begin
        int_reg_array_41_26_real <= _zz_2913_;
      end
      if(_zz_2875_)begin
        int_reg_array_41_27_real <= _zz_2913_;
      end
      if(_zz_2876_)begin
        int_reg_array_41_28_real <= _zz_2913_;
      end
      if(_zz_2877_)begin
        int_reg_array_41_29_real <= _zz_2913_;
      end
      if(_zz_2878_)begin
        int_reg_array_41_30_real <= _zz_2913_;
      end
      if(_zz_2879_)begin
        int_reg_array_41_31_real <= _zz_2913_;
      end
      if(_zz_2880_)begin
        int_reg_array_41_32_real <= _zz_2913_;
      end
      if(_zz_2881_)begin
        int_reg_array_41_33_real <= _zz_2913_;
      end
      if(_zz_2882_)begin
        int_reg_array_41_34_real <= _zz_2913_;
      end
      if(_zz_2883_)begin
        int_reg_array_41_35_real <= _zz_2913_;
      end
      if(_zz_2884_)begin
        int_reg_array_41_36_real <= _zz_2913_;
      end
      if(_zz_2885_)begin
        int_reg_array_41_37_real <= _zz_2913_;
      end
      if(_zz_2886_)begin
        int_reg_array_41_38_real <= _zz_2913_;
      end
      if(_zz_2887_)begin
        int_reg_array_41_39_real <= _zz_2913_;
      end
      if(_zz_2888_)begin
        int_reg_array_41_40_real <= _zz_2913_;
      end
      if(_zz_2889_)begin
        int_reg_array_41_41_real <= _zz_2913_;
      end
      if(_zz_2890_)begin
        int_reg_array_41_42_real <= _zz_2913_;
      end
      if(_zz_2891_)begin
        int_reg_array_41_43_real <= _zz_2913_;
      end
      if(_zz_2892_)begin
        int_reg_array_41_44_real <= _zz_2913_;
      end
      if(_zz_2893_)begin
        int_reg_array_41_45_real <= _zz_2913_;
      end
      if(_zz_2894_)begin
        int_reg_array_41_46_real <= _zz_2913_;
      end
      if(_zz_2895_)begin
        int_reg_array_41_47_real <= _zz_2913_;
      end
      if(_zz_2896_)begin
        int_reg_array_41_48_real <= _zz_2913_;
      end
      if(_zz_2897_)begin
        int_reg_array_41_49_real <= _zz_2913_;
      end
      if(_zz_2898_)begin
        int_reg_array_41_50_real <= _zz_2913_;
      end
      if(_zz_2899_)begin
        int_reg_array_41_51_real <= _zz_2913_;
      end
      if(_zz_2900_)begin
        int_reg_array_41_52_real <= _zz_2913_;
      end
      if(_zz_2901_)begin
        int_reg_array_41_53_real <= _zz_2913_;
      end
      if(_zz_2902_)begin
        int_reg_array_41_54_real <= _zz_2913_;
      end
      if(_zz_2903_)begin
        int_reg_array_41_55_real <= _zz_2913_;
      end
      if(_zz_2904_)begin
        int_reg_array_41_56_real <= _zz_2913_;
      end
      if(_zz_2905_)begin
        int_reg_array_41_57_real <= _zz_2913_;
      end
      if(_zz_2906_)begin
        int_reg_array_41_58_real <= _zz_2913_;
      end
      if(_zz_2907_)begin
        int_reg_array_41_59_real <= _zz_2913_;
      end
      if(_zz_2908_)begin
        int_reg_array_41_60_real <= _zz_2913_;
      end
      if(_zz_2909_)begin
        int_reg_array_41_61_real <= _zz_2913_;
      end
      if(_zz_2910_)begin
        int_reg_array_41_62_real <= _zz_2913_;
      end
      if(_zz_2911_)begin
        int_reg_array_41_63_real <= _zz_2913_;
      end
      if(_zz_2848_)begin
        int_reg_array_41_0_imag <= _zz_2914_;
      end
      if(_zz_2849_)begin
        int_reg_array_41_1_imag <= _zz_2914_;
      end
      if(_zz_2850_)begin
        int_reg_array_41_2_imag <= _zz_2914_;
      end
      if(_zz_2851_)begin
        int_reg_array_41_3_imag <= _zz_2914_;
      end
      if(_zz_2852_)begin
        int_reg_array_41_4_imag <= _zz_2914_;
      end
      if(_zz_2853_)begin
        int_reg_array_41_5_imag <= _zz_2914_;
      end
      if(_zz_2854_)begin
        int_reg_array_41_6_imag <= _zz_2914_;
      end
      if(_zz_2855_)begin
        int_reg_array_41_7_imag <= _zz_2914_;
      end
      if(_zz_2856_)begin
        int_reg_array_41_8_imag <= _zz_2914_;
      end
      if(_zz_2857_)begin
        int_reg_array_41_9_imag <= _zz_2914_;
      end
      if(_zz_2858_)begin
        int_reg_array_41_10_imag <= _zz_2914_;
      end
      if(_zz_2859_)begin
        int_reg_array_41_11_imag <= _zz_2914_;
      end
      if(_zz_2860_)begin
        int_reg_array_41_12_imag <= _zz_2914_;
      end
      if(_zz_2861_)begin
        int_reg_array_41_13_imag <= _zz_2914_;
      end
      if(_zz_2862_)begin
        int_reg_array_41_14_imag <= _zz_2914_;
      end
      if(_zz_2863_)begin
        int_reg_array_41_15_imag <= _zz_2914_;
      end
      if(_zz_2864_)begin
        int_reg_array_41_16_imag <= _zz_2914_;
      end
      if(_zz_2865_)begin
        int_reg_array_41_17_imag <= _zz_2914_;
      end
      if(_zz_2866_)begin
        int_reg_array_41_18_imag <= _zz_2914_;
      end
      if(_zz_2867_)begin
        int_reg_array_41_19_imag <= _zz_2914_;
      end
      if(_zz_2868_)begin
        int_reg_array_41_20_imag <= _zz_2914_;
      end
      if(_zz_2869_)begin
        int_reg_array_41_21_imag <= _zz_2914_;
      end
      if(_zz_2870_)begin
        int_reg_array_41_22_imag <= _zz_2914_;
      end
      if(_zz_2871_)begin
        int_reg_array_41_23_imag <= _zz_2914_;
      end
      if(_zz_2872_)begin
        int_reg_array_41_24_imag <= _zz_2914_;
      end
      if(_zz_2873_)begin
        int_reg_array_41_25_imag <= _zz_2914_;
      end
      if(_zz_2874_)begin
        int_reg_array_41_26_imag <= _zz_2914_;
      end
      if(_zz_2875_)begin
        int_reg_array_41_27_imag <= _zz_2914_;
      end
      if(_zz_2876_)begin
        int_reg_array_41_28_imag <= _zz_2914_;
      end
      if(_zz_2877_)begin
        int_reg_array_41_29_imag <= _zz_2914_;
      end
      if(_zz_2878_)begin
        int_reg_array_41_30_imag <= _zz_2914_;
      end
      if(_zz_2879_)begin
        int_reg_array_41_31_imag <= _zz_2914_;
      end
      if(_zz_2880_)begin
        int_reg_array_41_32_imag <= _zz_2914_;
      end
      if(_zz_2881_)begin
        int_reg_array_41_33_imag <= _zz_2914_;
      end
      if(_zz_2882_)begin
        int_reg_array_41_34_imag <= _zz_2914_;
      end
      if(_zz_2883_)begin
        int_reg_array_41_35_imag <= _zz_2914_;
      end
      if(_zz_2884_)begin
        int_reg_array_41_36_imag <= _zz_2914_;
      end
      if(_zz_2885_)begin
        int_reg_array_41_37_imag <= _zz_2914_;
      end
      if(_zz_2886_)begin
        int_reg_array_41_38_imag <= _zz_2914_;
      end
      if(_zz_2887_)begin
        int_reg_array_41_39_imag <= _zz_2914_;
      end
      if(_zz_2888_)begin
        int_reg_array_41_40_imag <= _zz_2914_;
      end
      if(_zz_2889_)begin
        int_reg_array_41_41_imag <= _zz_2914_;
      end
      if(_zz_2890_)begin
        int_reg_array_41_42_imag <= _zz_2914_;
      end
      if(_zz_2891_)begin
        int_reg_array_41_43_imag <= _zz_2914_;
      end
      if(_zz_2892_)begin
        int_reg_array_41_44_imag <= _zz_2914_;
      end
      if(_zz_2893_)begin
        int_reg_array_41_45_imag <= _zz_2914_;
      end
      if(_zz_2894_)begin
        int_reg_array_41_46_imag <= _zz_2914_;
      end
      if(_zz_2895_)begin
        int_reg_array_41_47_imag <= _zz_2914_;
      end
      if(_zz_2896_)begin
        int_reg_array_41_48_imag <= _zz_2914_;
      end
      if(_zz_2897_)begin
        int_reg_array_41_49_imag <= _zz_2914_;
      end
      if(_zz_2898_)begin
        int_reg_array_41_50_imag <= _zz_2914_;
      end
      if(_zz_2899_)begin
        int_reg_array_41_51_imag <= _zz_2914_;
      end
      if(_zz_2900_)begin
        int_reg_array_41_52_imag <= _zz_2914_;
      end
      if(_zz_2901_)begin
        int_reg_array_41_53_imag <= _zz_2914_;
      end
      if(_zz_2902_)begin
        int_reg_array_41_54_imag <= _zz_2914_;
      end
      if(_zz_2903_)begin
        int_reg_array_41_55_imag <= _zz_2914_;
      end
      if(_zz_2904_)begin
        int_reg_array_41_56_imag <= _zz_2914_;
      end
      if(_zz_2905_)begin
        int_reg_array_41_57_imag <= _zz_2914_;
      end
      if(_zz_2906_)begin
        int_reg_array_41_58_imag <= _zz_2914_;
      end
      if(_zz_2907_)begin
        int_reg_array_41_59_imag <= _zz_2914_;
      end
      if(_zz_2908_)begin
        int_reg_array_41_60_imag <= _zz_2914_;
      end
      if(_zz_2909_)begin
        int_reg_array_41_61_imag <= _zz_2914_;
      end
      if(_zz_2910_)begin
        int_reg_array_41_62_imag <= _zz_2914_;
      end
      if(_zz_2911_)begin
        int_reg_array_41_63_imag <= _zz_2914_;
      end
      if(_zz_2917_)begin
        int_reg_array_42_0_real <= _zz_2982_;
      end
      if(_zz_2918_)begin
        int_reg_array_42_1_real <= _zz_2982_;
      end
      if(_zz_2919_)begin
        int_reg_array_42_2_real <= _zz_2982_;
      end
      if(_zz_2920_)begin
        int_reg_array_42_3_real <= _zz_2982_;
      end
      if(_zz_2921_)begin
        int_reg_array_42_4_real <= _zz_2982_;
      end
      if(_zz_2922_)begin
        int_reg_array_42_5_real <= _zz_2982_;
      end
      if(_zz_2923_)begin
        int_reg_array_42_6_real <= _zz_2982_;
      end
      if(_zz_2924_)begin
        int_reg_array_42_7_real <= _zz_2982_;
      end
      if(_zz_2925_)begin
        int_reg_array_42_8_real <= _zz_2982_;
      end
      if(_zz_2926_)begin
        int_reg_array_42_9_real <= _zz_2982_;
      end
      if(_zz_2927_)begin
        int_reg_array_42_10_real <= _zz_2982_;
      end
      if(_zz_2928_)begin
        int_reg_array_42_11_real <= _zz_2982_;
      end
      if(_zz_2929_)begin
        int_reg_array_42_12_real <= _zz_2982_;
      end
      if(_zz_2930_)begin
        int_reg_array_42_13_real <= _zz_2982_;
      end
      if(_zz_2931_)begin
        int_reg_array_42_14_real <= _zz_2982_;
      end
      if(_zz_2932_)begin
        int_reg_array_42_15_real <= _zz_2982_;
      end
      if(_zz_2933_)begin
        int_reg_array_42_16_real <= _zz_2982_;
      end
      if(_zz_2934_)begin
        int_reg_array_42_17_real <= _zz_2982_;
      end
      if(_zz_2935_)begin
        int_reg_array_42_18_real <= _zz_2982_;
      end
      if(_zz_2936_)begin
        int_reg_array_42_19_real <= _zz_2982_;
      end
      if(_zz_2937_)begin
        int_reg_array_42_20_real <= _zz_2982_;
      end
      if(_zz_2938_)begin
        int_reg_array_42_21_real <= _zz_2982_;
      end
      if(_zz_2939_)begin
        int_reg_array_42_22_real <= _zz_2982_;
      end
      if(_zz_2940_)begin
        int_reg_array_42_23_real <= _zz_2982_;
      end
      if(_zz_2941_)begin
        int_reg_array_42_24_real <= _zz_2982_;
      end
      if(_zz_2942_)begin
        int_reg_array_42_25_real <= _zz_2982_;
      end
      if(_zz_2943_)begin
        int_reg_array_42_26_real <= _zz_2982_;
      end
      if(_zz_2944_)begin
        int_reg_array_42_27_real <= _zz_2982_;
      end
      if(_zz_2945_)begin
        int_reg_array_42_28_real <= _zz_2982_;
      end
      if(_zz_2946_)begin
        int_reg_array_42_29_real <= _zz_2982_;
      end
      if(_zz_2947_)begin
        int_reg_array_42_30_real <= _zz_2982_;
      end
      if(_zz_2948_)begin
        int_reg_array_42_31_real <= _zz_2982_;
      end
      if(_zz_2949_)begin
        int_reg_array_42_32_real <= _zz_2982_;
      end
      if(_zz_2950_)begin
        int_reg_array_42_33_real <= _zz_2982_;
      end
      if(_zz_2951_)begin
        int_reg_array_42_34_real <= _zz_2982_;
      end
      if(_zz_2952_)begin
        int_reg_array_42_35_real <= _zz_2982_;
      end
      if(_zz_2953_)begin
        int_reg_array_42_36_real <= _zz_2982_;
      end
      if(_zz_2954_)begin
        int_reg_array_42_37_real <= _zz_2982_;
      end
      if(_zz_2955_)begin
        int_reg_array_42_38_real <= _zz_2982_;
      end
      if(_zz_2956_)begin
        int_reg_array_42_39_real <= _zz_2982_;
      end
      if(_zz_2957_)begin
        int_reg_array_42_40_real <= _zz_2982_;
      end
      if(_zz_2958_)begin
        int_reg_array_42_41_real <= _zz_2982_;
      end
      if(_zz_2959_)begin
        int_reg_array_42_42_real <= _zz_2982_;
      end
      if(_zz_2960_)begin
        int_reg_array_42_43_real <= _zz_2982_;
      end
      if(_zz_2961_)begin
        int_reg_array_42_44_real <= _zz_2982_;
      end
      if(_zz_2962_)begin
        int_reg_array_42_45_real <= _zz_2982_;
      end
      if(_zz_2963_)begin
        int_reg_array_42_46_real <= _zz_2982_;
      end
      if(_zz_2964_)begin
        int_reg_array_42_47_real <= _zz_2982_;
      end
      if(_zz_2965_)begin
        int_reg_array_42_48_real <= _zz_2982_;
      end
      if(_zz_2966_)begin
        int_reg_array_42_49_real <= _zz_2982_;
      end
      if(_zz_2967_)begin
        int_reg_array_42_50_real <= _zz_2982_;
      end
      if(_zz_2968_)begin
        int_reg_array_42_51_real <= _zz_2982_;
      end
      if(_zz_2969_)begin
        int_reg_array_42_52_real <= _zz_2982_;
      end
      if(_zz_2970_)begin
        int_reg_array_42_53_real <= _zz_2982_;
      end
      if(_zz_2971_)begin
        int_reg_array_42_54_real <= _zz_2982_;
      end
      if(_zz_2972_)begin
        int_reg_array_42_55_real <= _zz_2982_;
      end
      if(_zz_2973_)begin
        int_reg_array_42_56_real <= _zz_2982_;
      end
      if(_zz_2974_)begin
        int_reg_array_42_57_real <= _zz_2982_;
      end
      if(_zz_2975_)begin
        int_reg_array_42_58_real <= _zz_2982_;
      end
      if(_zz_2976_)begin
        int_reg_array_42_59_real <= _zz_2982_;
      end
      if(_zz_2977_)begin
        int_reg_array_42_60_real <= _zz_2982_;
      end
      if(_zz_2978_)begin
        int_reg_array_42_61_real <= _zz_2982_;
      end
      if(_zz_2979_)begin
        int_reg_array_42_62_real <= _zz_2982_;
      end
      if(_zz_2980_)begin
        int_reg_array_42_63_real <= _zz_2982_;
      end
      if(_zz_2917_)begin
        int_reg_array_42_0_imag <= _zz_2983_;
      end
      if(_zz_2918_)begin
        int_reg_array_42_1_imag <= _zz_2983_;
      end
      if(_zz_2919_)begin
        int_reg_array_42_2_imag <= _zz_2983_;
      end
      if(_zz_2920_)begin
        int_reg_array_42_3_imag <= _zz_2983_;
      end
      if(_zz_2921_)begin
        int_reg_array_42_4_imag <= _zz_2983_;
      end
      if(_zz_2922_)begin
        int_reg_array_42_5_imag <= _zz_2983_;
      end
      if(_zz_2923_)begin
        int_reg_array_42_6_imag <= _zz_2983_;
      end
      if(_zz_2924_)begin
        int_reg_array_42_7_imag <= _zz_2983_;
      end
      if(_zz_2925_)begin
        int_reg_array_42_8_imag <= _zz_2983_;
      end
      if(_zz_2926_)begin
        int_reg_array_42_9_imag <= _zz_2983_;
      end
      if(_zz_2927_)begin
        int_reg_array_42_10_imag <= _zz_2983_;
      end
      if(_zz_2928_)begin
        int_reg_array_42_11_imag <= _zz_2983_;
      end
      if(_zz_2929_)begin
        int_reg_array_42_12_imag <= _zz_2983_;
      end
      if(_zz_2930_)begin
        int_reg_array_42_13_imag <= _zz_2983_;
      end
      if(_zz_2931_)begin
        int_reg_array_42_14_imag <= _zz_2983_;
      end
      if(_zz_2932_)begin
        int_reg_array_42_15_imag <= _zz_2983_;
      end
      if(_zz_2933_)begin
        int_reg_array_42_16_imag <= _zz_2983_;
      end
      if(_zz_2934_)begin
        int_reg_array_42_17_imag <= _zz_2983_;
      end
      if(_zz_2935_)begin
        int_reg_array_42_18_imag <= _zz_2983_;
      end
      if(_zz_2936_)begin
        int_reg_array_42_19_imag <= _zz_2983_;
      end
      if(_zz_2937_)begin
        int_reg_array_42_20_imag <= _zz_2983_;
      end
      if(_zz_2938_)begin
        int_reg_array_42_21_imag <= _zz_2983_;
      end
      if(_zz_2939_)begin
        int_reg_array_42_22_imag <= _zz_2983_;
      end
      if(_zz_2940_)begin
        int_reg_array_42_23_imag <= _zz_2983_;
      end
      if(_zz_2941_)begin
        int_reg_array_42_24_imag <= _zz_2983_;
      end
      if(_zz_2942_)begin
        int_reg_array_42_25_imag <= _zz_2983_;
      end
      if(_zz_2943_)begin
        int_reg_array_42_26_imag <= _zz_2983_;
      end
      if(_zz_2944_)begin
        int_reg_array_42_27_imag <= _zz_2983_;
      end
      if(_zz_2945_)begin
        int_reg_array_42_28_imag <= _zz_2983_;
      end
      if(_zz_2946_)begin
        int_reg_array_42_29_imag <= _zz_2983_;
      end
      if(_zz_2947_)begin
        int_reg_array_42_30_imag <= _zz_2983_;
      end
      if(_zz_2948_)begin
        int_reg_array_42_31_imag <= _zz_2983_;
      end
      if(_zz_2949_)begin
        int_reg_array_42_32_imag <= _zz_2983_;
      end
      if(_zz_2950_)begin
        int_reg_array_42_33_imag <= _zz_2983_;
      end
      if(_zz_2951_)begin
        int_reg_array_42_34_imag <= _zz_2983_;
      end
      if(_zz_2952_)begin
        int_reg_array_42_35_imag <= _zz_2983_;
      end
      if(_zz_2953_)begin
        int_reg_array_42_36_imag <= _zz_2983_;
      end
      if(_zz_2954_)begin
        int_reg_array_42_37_imag <= _zz_2983_;
      end
      if(_zz_2955_)begin
        int_reg_array_42_38_imag <= _zz_2983_;
      end
      if(_zz_2956_)begin
        int_reg_array_42_39_imag <= _zz_2983_;
      end
      if(_zz_2957_)begin
        int_reg_array_42_40_imag <= _zz_2983_;
      end
      if(_zz_2958_)begin
        int_reg_array_42_41_imag <= _zz_2983_;
      end
      if(_zz_2959_)begin
        int_reg_array_42_42_imag <= _zz_2983_;
      end
      if(_zz_2960_)begin
        int_reg_array_42_43_imag <= _zz_2983_;
      end
      if(_zz_2961_)begin
        int_reg_array_42_44_imag <= _zz_2983_;
      end
      if(_zz_2962_)begin
        int_reg_array_42_45_imag <= _zz_2983_;
      end
      if(_zz_2963_)begin
        int_reg_array_42_46_imag <= _zz_2983_;
      end
      if(_zz_2964_)begin
        int_reg_array_42_47_imag <= _zz_2983_;
      end
      if(_zz_2965_)begin
        int_reg_array_42_48_imag <= _zz_2983_;
      end
      if(_zz_2966_)begin
        int_reg_array_42_49_imag <= _zz_2983_;
      end
      if(_zz_2967_)begin
        int_reg_array_42_50_imag <= _zz_2983_;
      end
      if(_zz_2968_)begin
        int_reg_array_42_51_imag <= _zz_2983_;
      end
      if(_zz_2969_)begin
        int_reg_array_42_52_imag <= _zz_2983_;
      end
      if(_zz_2970_)begin
        int_reg_array_42_53_imag <= _zz_2983_;
      end
      if(_zz_2971_)begin
        int_reg_array_42_54_imag <= _zz_2983_;
      end
      if(_zz_2972_)begin
        int_reg_array_42_55_imag <= _zz_2983_;
      end
      if(_zz_2973_)begin
        int_reg_array_42_56_imag <= _zz_2983_;
      end
      if(_zz_2974_)begin
        int_reg_array_42_57_imag <= _zz_2983_;
      end
      if(_zz_2975_)begin
        int_reg_array_42_58_imag <= _zz_2983_;
      end
      if(_zz_2976_)begin
        int_reg_array_42_59_imag <= _zz_2983_;
      end
      if(_zz_2977_)begin
        int_reg_array_42_60_imag <= _zz_2983_;
      end
      if(_zz_2978_)begin
        int_reg_array_42_61_imag <= _zz_2983_;
      end
      if(_zz_2979_)begin
        int_reg_array_42_62_imag <= _zz_2983_;
      end
      if(_zz_2980_)begin
        int_reg_array_42_63_imag <= _zz_2983_;
      end
      if(_zz_2986_)begin
        int_reg_array_43_0_real <= _zz_3051_;
      end
      if(_zz_2987_)begin
        int_reg_array_43_1_real <= _zz_3051_;
      end
      if(_zz_2988_)begin
        int_reg_array_43_2_real <= _zz_3051_;
      end
      if(_zz_2989_)begin
        int_reg_array_43_3_real <= _zz_3051_;
      end
      if(_zz_2990_)begin
        int_reg_array_43_4_real <= _zz_3051_;
      end
      if(_zz_2991_)begin
        int_reg_array_43_5_real <= _zz_3051_;
      end
      if(_zz_2992_)begin
        int_reg_array_43_6_real <= _zz_3051_;
      end
      if(_zz_2993_)begin
        int_reg_array_43_7_real <= _zz_3051_;
      end
      if(_zz_2994_)begin
        int_reg_array_43_8_real <= _zz_3051_;
      end
      if(_zz_2995_)begin
        int_reg_array_43_9_real <= _zz_3051_;
      end
      if(_zz_2996_)begin
        int_reg_array_43_10_real <= _zz_3051_;
      end
      if(_zz_2997_)begin
        int_reg_array_43_11_real <= _zz_3051_;
      end
      if(_zz_2998_)begin
        int_reg_array_43_12_real <= _zz_3051_;
      end
      if(_zz_2999_)begin
        int_reg_array_43_13_real <= _zz_3051_;
      end
      if(_zz_3000_)begin
        int_reg_array_43_14_real <= _zz_3051_;
      end
      if(_zz_3001_)begin
        int_reg_array_43_15_real <= _zz_3051_;
      end
      if(_zz_3002_)begin
        int_reg_array_43_16_real <= _zz_3051_;
      end
      if(_zz_3003_)begin
        int_reg_array_43_17_real <= _zz_3051_;
      end
      if(_zz_3004_)begin
        int_reg_array_43_18_real <= _zz_3051_;
      end
      if(_zz_3005_)begin
        int_reg_array_43_19_real <= _zz_3051_;
      end
      if(_zz_3006_)begin
        int_reg_array_43_20_real <= _zz_3051_;
      end
      if(_zz_3007_)begin
        int_reg_array_43_21_real <= _zz_3051_;
      end
      if(_zz_3008_)begin
        int_reg_array_43_22_real <= _zz_3051_;
      end
      if(_zz_3009_)begin
        int_reg_array_43_23_real <= _zz_3051_;
      end
      if(_zz_3010_)begin
        int_reg_array_43_24_real <= _zz_3051_;
      end
      if(_zz_3011_)begin
        int_reg_array_43_25_real <= _zz_3051_;
      end
      if(_zz_3012_)begin
        int_reg_array_43_26_real <= _zz_3051_;
      end
      if(_zz_3013_)begin
        int_reg_array_43_27_real <= _zz_3051_;
      end
      if(_zz_3014_)begin
        int_reg_array_43_28_real <= _zz_3051_;
      end
      if(_zz_3015_)begin
        int_reg_array_43_29_real <= _zz_3051_;
      end
      if(_zz_3016_)begin
        int_reg_array_43_30_real <= _zz_3051_;
      end
      if(_zz_3017_)begin
        int_reg_array_43_31_real <= _zz_3051_;
      end
      if(_zz_3018_)begin
        int_reg_array_43_32_real <= _zz_3051_;
      end
      if(_zz_3019_)begin
        int_reg_array_43_33_real <= _zz_3051_;
      end
      if(_zz_3020_)begin
        int_reg_array_43_34_real <= _zz_3051_;
      end
      if(_zz_3021_)begin
        int_reg_array_43_35_real <= _zz_3051_;
      end
      if(_zz_3022_)begin
        int_reg_array_43_36_real <= _zz_3051_;
      end
      if(_zz_3023_)begin
        int_reg_array_43_37_real <= _zz_3051_;
      end
      if(_zz_3024_)begin
        int_reg_array_43_38_real <= _zz_3051_;
      end
      if(_zz_3025_)begin
        int_reg_array_43_39_real <= _zz_3051_;
      end
      if(_zz_3026_)begin
        int_reg_array_43_40_real <= _zz_3051_;
      end
      if(_zz_3027_)begin
        int_reg_array_43_41_real <= _zz_3051_;
      end
      if(_zz_3028_)begin
        int_reg_array_43_42_real <= _zz_3051_;
      end
      if(_zz_3029_)begin
        int_reg_array_43_43_real <= _zz_3051_;
      end
      if(_zz_3030_)begin
        int_reg_array_43_44_real <= _zz_3051_;
      end
      if(_zz_3031_)begin
        int_reg_array_43_45_real <= _zz_3051_;
      end
      if(_zz_3032_)begin
        int_reg_array_43_46_real <= _zz_3051_;
      end
      if(_zz_3033_)begin
        int_reg_array_43_47_real <= _zz_3051_;
      end
      if(_zz_3034_)begin
        int_reg_array_43_48_real <= _zz_3051_;
      end
      if(_zz_3035_)begin
        int_reg_array_43_49_real <= _zz_3051_;
      end
      if(_zz_3036_)begin
        int_reg_array_43_50_real <= _zz_3051_;
      end
      if(_zz_3037_)begin
        int_reg_array_43_51_real <= _zz_3051_;
      end
      if(_zz_3038_)begin
        int_reg_array_43_52_real <= _zz_3051_;
      end
      if(_zz_3039_)begin
        int_reg_array_43_53_real <= _zz_3051_;
      end
      if(_zz_3040_)begin
        int_reg_array_43_54_real <= _zz_3051_;
      end
      if(_zz_3041_)begin
        int_reg_array_43_55_real <= _zz_3051_;
      end
      if(_zz_3042_)begin
        int_reg_array_43_56_real <= _zz_3051_;
      end
      if(_zz_3043_)begin
        int_reg_array_43_57_real <= _zz_3051_;
      end
      if(_zz_3044_)begin
        int_reg_array_43_58_real <= _zz_3051_;
      end
      if(_zz_3045_)begin
        int_reg_array_43_59_real <= _zz_3051_;
      end
      if(_zz_3046_)begin
        int_reg_array_43_60_real <= _zz_3051_;
      end
      if(_zz_3047_)begin
        int_reg_array_43_61_real <= _zz_3051_;
      end
      if(_zz_3048_)begin
        int_reg_array_43_62_real <= _zz_3051_;
      end
      if(_zz_3049_)begin
        int_reg_array_43_63_real <= _zz_3051_;
      end
      if(_zz_2986_)begin
        int_reg_array_43_0_imag <= _zz_3052_;
      end
      if(_zz_2987_)begin
        int_reg_array_43_1_imag <= _zz_3052_;
      end
      if(_zz_2988_)begin
        int_reg_array_43_2_imag <= _zz_3052_;
      end
      if(_zz_2989_)begin
        int_reg_array_43_3_imag <= _zz_3052_;
      end
      if(_zz_2990_)begin
        int_reg_array_43_4_imag <= _zz_3052_;
      end
      if(_zz_2991_)begin
        int_reg_array_43_5_imag <= _zz_3052_;
      end
      if(_zz_2992_)begin
        int_reg_array_43_6_imag <= _zz_3052_;
      end
      if(_zz_2993_)begin
        int_reg_array_43_7_imag <= _zz_3052_;
      end
      if(_zz_2994_)begin
        int_reg_array_43_8_imag <= _zz_3052_;
      end
      if(_zz_2995_)begin
        int_reg_array_43_9_imag <= _zz_3052_;
      end
      if(_zz_2996_)begin
        int_reg_array_43_10_imag <= _zz_3052_;
      end
      if(_zz_2997_)begin
        int_reg_array_43_11_imag <= _zz_3052_;
      end
      if(_zz_2998_)begin
        int_reg_array_43_12_imag <= _zz_3052_;
      end
      if(_zz_2999_)begin
        int_reg_array_43_13_imag <= _zz_3052_;
      end
      if(_zz_3000_)begin
        int_reg_array_43_14_imag <= _zz_3052_;
      end
      if(_zz_3001_)begin
        int_reg_array_43_15_imag <= _zz_3052_;
      end
      if(_zz_3002_)begin
        int_reg_array_43_16_imag <= _zz_3052_;
      end
      if(_zz_3003_)begin
        int_reg_array_43_17_imag <= _zz_3052_;
      end
      if(_zz_3004_)begin
        int_reg_array_43_18_imag <= _zz_3052_;
      end
      if(_zz_3005_)begin
        int_reg_array_43_19_imag <= _zz_3052_;
      end
      if(_zz_3006_)begin
        int_reg_array_43_20_imag <= _zz_3052_;
      end
      if(_zz_3007_)begin
        int_reg_array_43_21_imag <= _zz_3052_;
      end
      if(_zz_3008_)begin
        int_reg_array_43_22_imag <= _zz_3052_;
      end
      if(_zz_3009_)begin
        int_reg_array_43_23_imag <= _zz_3052_;
      end
      if(_zz_3010_)begin
        int_reg_array_43_24_imag <= _zz_3052_;
      end
      if(_zz_3011_)begin
        int_reg_array_43_25_imag <= _zz_3052_;
      end
      if(_zz_3012_)begin
        int_reg_array_43_26_imag <= _zz_3052_;
      end
      if(_zz_3013_)begin
        int_reg_array_43_27_imag <= _zz_3052_;
      end
      if(_zz_3014_)begin
        int_reg_array_43_28_imag <= _zz_3052_;
      end
      if(_zz_3015_)begin
        int_reg_array_43_29_imag <= _zz_3052_;
      end
      if(_zz_3016_)begin
        int_reg_array_43_30_imag <= _zz_3052_;
      end
      if(_zz_3017_)begin
        int_reg_array_43_31_imag <= _zz_3052_;
      end
      if(_zz_3018_)begin
        int_reg_array_43_32_imag <= _zz_3052_;
      end
      if(_zz_3019_)begin
        int_reg_array_43_33_imag <= _zz_3052_;
      end
      if(_zz_3020_)begin
        int_reg_array_43_34_imag <= _zz_3052_;
      end
      if(_zz_3021_)begin
        int_reg_array_43_35_imag <= _zz_3052_;
      end
      if(_zz_3022_)begin
        int_reg_array_43_36_imag <= _zz_3052_;
      end
      if(_zz_3023_)begin
        int_reg_array_43_37_imag <= _zz_3052_;
      end
      if(_zz_3024_)begin
        int_reg_array_43_38_imag <= _zz_3052_;
      end
      if(_zz_3025_)begin
        int_reg_array_43_39_imag <= _zz_3052_;
      end
      if(_zz_3026_)begin
        int_reg_array_43_40_imag <= _zz_3052_;
      end
      if(_zz_3027_)begin
        int_reg_array_43_41_imag <= _zz_3052_;
      end
      if(_zz_3028_)begin
        int_reg_array_43_42_imag <= _zz_3052_;
      end
      if(_zz_3029_)begin
        int_reg_array_43_43_imag <= _zz_3052_;
      end
      if(_zz_3030_)begin
        int_reg_array_43_44_imag <= _zz_3052_;
      end
      if(_zz_3031_)begin
        int_reg_array_43_45_imag <= _zz_3052_;
      end
      if(_zz_3032_)begin
        int_reg_array_43_46_imag <= _zz_3052_;
      end
      if(_zz_3033_)begin
        int_reg_array_43_47_imag <= _zz_3052_;
      end
      if(_zz_3034_)begin
        int_reg_array_43_48_imag <= _zz_3052_;
      end
      if(_zz_3035_)begin
        int_reg_array_43_49_imag <= _zz_3052_;
      end
      if(_zz_3036_)begin
        int_reg_array_43_50_imag <= _zz_3052_;
      end
      if(_zz_3037_)begin
        int_reg_array_43_51_imag <= _zz_3052_;
      end
      if(_zz_3038_)begin
        int_reg_array_43_52_imag <= _zz_3052_;
      end
      if(_zz_3039_)begin
        int_reg_array_43_53_imag <= _zz_3052_;
      end
      if(_zz_3040_)begin
        int_reg_array_43_54_imag <= _zz_3052_;
      end
      if(_zz_3041_)begin
        int_reg_array_43_55_imag <= _zz_3052_;
      end
      if(_zz_3042_)begin
        int_reg_array_43_56_imag <= _zz_3052_;
      end
      if(_zz_3043_)begin
        int_reg_array_43_57_imag <= _zz_3052_;
      end
      if(_zz_3044_)begin
        int_reg_array_43_58_imag <= _zz_3052_;
      end
      if(_zz_3045_)begin
        int_reg_array_43_59_imag <= _zz_3052_;
      end
      if(_zz_3046_)begin
        int_reg_array_43_60_imag <= _zz_3052_;
      end
      if(_zz_3047_)begin
        int_reg_array_43_61_imag <= _zz_3052_;
      end
      if(_zz_3048_)begin
        int_reg_array_43_62_imag <= _zz_3052_;
      end
      if(_zz_3049_)begin
        int_reg_array_43_63_imag <= _zz_3052_;
      end
      if(_zz_3055_)begin
        int_reg_array_44_0_real <= _zz_3120_;
      end
      if(_zz_3056_)begin
        int_reg_array_44_1_real <= _zz_3120_;
      end
      if(_zz_3057_)begin
        int_reg_array_44_2_real <= _zz_3120_;
      end
      if(_zz_3058_)begin
        int_reg_array_44_3_real <= _zz_3120_;
      end
      if(_zz_3059_)begin
        int_reg_array_44_4_real <= _zz_3120_;
      end
      if(_zz_3060_)begin
        int_reg_array_44_5_real <= _zz_3120_;
      end
      if(_zz_3061_)begin
        int_reg_array_44_6_real <= _zz_3120_;
      end
      if(_zz_3062_)begin
        int_reg_array_44_7_real <= _zz_3120_;
      end
      if(_zz_3063_)begin
        int_reg_array_44_8_real <= _zz_3120_;
      end
      if(_zz_3064_)begin
        int_reg_array_44_9_real <= _zz_3120_;
      end
      if(_zz_3065_)begin
        int_reg_array_44_10_real <= _zz_3120_;
      end
      if(_zz_3066_)begin
        int_reg_array_44_11_real <= _zz_3120_;
      end
      if(_zz_3067_)begin
        int_reg_array_44_12_real <= _zz_3120_;
      end
      if(_zz_3068_)begin
        int_reg_array_44_13_real <= _zz_3120_;
      end
      if(_zz_3069_)begin
        int_reg_array_44_14_real <= _zz_3120_;
      end
      if(_zz_3070_)begin
        int_reg_array_44_15_real <= _zz_3120_;
      end
      if(_zz_3071_)begin
        int_reg_array_44_16_real <= _zz_3120_;
      end
      if(_zz_3072_)begin
        int_reg_array_44_17_real <= _zz_3120_;
      end
      if(_zz_3073_)begin
        int_reg_array_44_18_real <= _zz_3120_;
      end
      if(_zz_3074_)begin
        int_reg_array_44_19_real <= _zz_3120_;
      end
      if(_zz_3075_)begin
        int_reg_array_44_20_real <= _zz_3120_;
      end
      if(_zz_3076_)begin
        int_reg_array_44_21_real <= _zz_3120_;
      end
      if(_zz_3077_)begin
        int_reg_array_44_22_real <= _zz_3120_;
      end
      if(_zz_3078_)begin
        int_reg_array_44_23_real <= _zz_3120_;
      end
      if(_zz_3079_)begin
        int_reg_array_44_24_real <= _zz_3120_;
      end
      if(_zz_3080_)begin
        int_reg_array_44_25_real <= _zz_3120_;
      end
      if(_zz_3081_)begin
        int_reg_array_44_26_real <= _zz_3120_;
      end
      if(_zz_3082_)begin
        int_reg_array_44_27_real <= _zz_3120_;
      end
      if(_zz_3083_)begin
        int_reg_array_44_28_real <= _zz_3120_;
      end
      if(_zz_3084_)begin
        int_reg_array_44_29_real <= _zz_3120_;
      end
      if(_zz_3085_)begin
        int_reg_array_44_30_real <= _zz_3120_;
      end
      if(_zz_3086_)begin
        int_reg_array_44_31_real <= _zz_3120_;
      end
      if(_zz_3087_)begin
        int_reg_array_44_32_real <= _zz_3120_;
      end
      if(_zz_3088_)begin
        int_reg_array_44_33_real <= _zz_3120_;
      end
      if(_zz_3089_)begin
        int_reg_array_44_34_real <= _zz_3120_;
      end
      if(_zz_3090_)begin
        int_reg_array_44_35_real <= _zz_3120_;
      end
      if(_zz_3091_)begin
        int_reg_array_44_36_real <= _zz_3120_;
      end
      if(_zz_3092_)begin
        int_reg_array_44_37_real <= _zz_3120_;
      end
      if(_zz_3093_)begin
        int_reg_array_44_38_real <= _zz_3120_;
      end
      if(_zz_3094_)begin
        int_reg_array_44_39_real <= _zz_3120_;
      end
      if(_zz_3095_)begin
        int_reg_array_44_40_real <= _zz_3120_;
      end
      if(_zz_3096_)begin
        int_reg_array_44_41_real <= _zz_3120_;
      end
      if(_zz_3097_)begin
        int_reg_array_44_42_real <= _zz_3120_;
      end
      if(_zz_3098_)begin
        int_reg_array_44_43_real <= _zz_3120_;
      end
      if(_zz_3099_)begin
        int_reg_array_44_44_real <= _zz_3120_;
      end
      if(_zz_3100_)begin
        int_reg_array_44_45_real <= _zz_3120_;
      end
      if(_zz_3101_)begin
        int_reg_array_44_46_real <= _zz_3120_;
      end
      if(_zz_3102_)begin
        int_reg_array_44_47_real <= _zz_3120_;
      end
      if(_zz_3103_)begin
        int_reg_array_44_48_real <= _zz_3120_;
      end
      if(_zz_3104_)begin
        int_reg_array_44_49_real <= _zz_3120_;
      end
      if(_zz_3105_)begin
        int_reg_array_44_50_real <= _zz_3120_;
      end
      if(_zz_3106_)begin
        int_reg_array_44_51_real <= _zz_3120_;
      end
      if(_zz_3107_)begin
        int_reg_array_44_52_real <= _zz_3120_;
      end
      if(_zz_3108_)begin
        int_reg_array_44_53_real <= _zz_3120_;
      end
      if(_zz_3109_)begin
        int_reg_array_44_54_real <= _zz_3120_;
      end
      if(_zz_3110_)begin
        int_reg_array_44_55_real <= _zz_3120_;
      end
      if(_zz_3111_)begin
        int_reg_array_44_56_real <= _zz_3120_;
      end
      if(_zz_3112_)begin
        int_reg_array_44_57_real <= _zz_3120_;
      end
      if(_zz_3113_)begin
        int_reg_array_44_58_real <= _zz_3120_;
      end
      if(_zz_3114_)begin
        int_reg_array_44_59_real <= _zz_3120_;
      end
      if(_zz_3115_)begin
        int_reg_array_44_60_real <= _zz_3120_;
      end
      if(_zz_3116_)begin
        int_reg_array_44_61_real <= _zz_3120_;
      end
      if(_zz_3117_)begin
        int_reg_array_44_62_real <= _zz_3120_;
      end
      if(_zz_3118_)begin
        int_reg_array_44_63_real <= _zz_3120_;
      end
      if(_zz_3055_)begin
        int_reg_array_44_0_imag <= _zz_3121_;
      end
      if(_zz_3056_)begin
        int_reg_array_44_1_imag <= _zz_3121_;
      end
      if(_zz_3057_)begin
        int_reg_array_44_2_imag <= _zz_3121_;
      end
      if(_zz_3058_)begin
        int_reg_array_44_3_imag <= _zz_3121_;
      end
      if(_zz_3059_)begin
        int_reg_array_44_4_imag <= _zz_3121_;
      end
      if(_zz_3060_)begin
        int_reg_array_44_5_imag <= _zz_3121_;
      end
      if(_zz_3061_)begin
        int_reg_array_44_6_imag <= _zz_3121_;
      end
      if(_zz_3062_)begin
        int_reg_array_44_7_imag <= _zz_3121_;
      end
      if(_zz_3063_)begin
        int_reg_array_44_8_imag <= _zz_3121_;
      end
      if(_zz_3064_)begin
        int_reg_array_44_9_imag <= _zz_3121_;
      end
      if(_zz_3065_)begin
        int_reg_array_44_10_imag <= _zz_3121_;
      end
      if(_zz_3066_)begin
        int_reg_array_44_11_imag <= _zz_3121_;
      end
      if(_zz_3067_)begin
        int_reg_array_44_12_imag <= _zz_3121_;
      end
      if(_zz_3068_)begin
        int_reg_array_44_13_imag <= _zz_3121_;
      end
      if(_zz_3069_)begin
        int_reg_array_44_14_imag <= _zz_3121_;
      end
      if(_zz_3070_)begin
        int_reg_array_44_15_imag <= _zz_3121_;
      end
      if(_zz_3071_)begin
        int_reg_array_44_16_imag <= _zz_3121_;
      end
      if(_zz_3072_)begin
        int_reg_array_44_17_imag <= _zz_3121_;
      end
      if(_zz_3073_)begin
        int_reg_array_44_18_imag <= _zz_3121_;
      end
      if(_zz_3074_)begin
        int_reg_array_44_19_imag <= _zz_3121_;
      end
      if(_zz_3075_)begin
        int_reg_array_44_20_imag <= _zz_3121_;
      end
      if(_zz_3076_)begin
        int_reg_array_44_21_imag <= _zz_3121_;
      end
      if(_zz_3077_)begin
        int_reg_array_44_22_imag <= _zz_3121_;
      end
      if(_zz_3078_)begin
        int_reg_array_44_23_imag <= _zz_3121_;
      end
      if(_zz_3079_)begin
        int_reg_array_44_24_imag <= _zz_3121_;
      end
      if(_zz_3080_)begin
        int_reg_array_44_25_imag <= _zz_3121_;
      end
      if(_zz_3081_)begin
        int_reg_array_44_26_imag <= _zz_3121_;
      end
      if(_zz_3082_)begin
        int_reg_array_44_27_imag <= _zz_3121_;
      end
      if(_zz_3083_)begin
        int_reg_array_44_28_imag <= _zz_3121_;
      end
      if(_zz_3084_)begin
        int_reg_array_44_29_imag <= _zz_3121_;
      end
      if(_zz_3085_)begin
        int_reg_array_44_30_imag <= _zz_3121_;
      end
      if(_zz_3086_)begin
        int_reg_array_44_31_imag <= _zz_3121_;
      end
      if(_zz_3087_)begin
        int_reg_array_44_32_imag <= _zz_3121_;
      end
      if(_zz_3088_)begin
        int_reg_array_44_33_imag <= _zz_3121_;
      end
      if(_zz_3089_)begin
        int_reg_array_44_34_imag <= _zz_3121_;
      end
      if(_zz_3090_)begin
        int_reg_array_44_35_imag <= _zz_3121_;
      end
      if(_zz_3091_)begin
        int_reg_array_44_36_imag <= _zz_3121_;
      end
      if(_zz_3092_)begin
        int_reg_array_44_37_imag <= _zz_3121_;
      end
      if(_zz_3093_)begin
        int_reg_array_44_38_imag <= _zz_3121_;
      end
      if(_zz_3094_)begin
        int_reg_array_44_39_imag <= _zz_3121_;
      end
      if(_zz_3095_)begin
        int_reg_array_44_40_imag <= _zz_3121_;
      end
      if(_zz_3096_)begin
        int_reg_array_44_41_imag <= _zz_3121_;
      end
      if(_zz_3097_)begin
        int_reg_array_44_42_imag <= _zz_3121_;
      end
      if(_zz_3098_)begin
        int_reg_array_44_43_imag <= _zz_3121_;
      end
      if(_zz_3099_)begin
        int_reg_array_44_44_imag <= _zz_3121_;
      end
      if(_zz_3100_)begin
        int_reg_array_44_45_imag <= _zz_3121_;
      end
      if(_zz_3101_)begin
        int_reg_array_44_46_imag <= _zz_3121_;
      end
      if(_zz_3102_)begin
        int_reg_array_44_47_imag <= _zz_3121_;
      end
      if(_zz_3103_)begin
        int_reg_array_44_48_imag <= _zz_3121_;
      end
      if(_zz_3104_)begin
        int_reg_array_44_49_imag <= _zz_3121_;
      end
      if(_zz_3105_)begin
        int_reg_array_44_50_imag <= _zz_3121_;
      end
      if(_zz_3106_)begin
        int_reg_array_44_51_imag <= _zz_3121_;
      end
      if(_zz_3107_)begin
        int_reg_array_44_52_imag <= _zz_3121_;
      end
      if(_zz_3108_)begin
        int_reg_array_44_53_imag <= _zz_3121_;
      end
      if(_zz_3109_)begin
        int_reg_array_44_54_imag <= _zz_3121_;
      end
      if(_zz_3110_)begin
        int_reg_array_44_55_imag <= _zz_3121_;
      end
      if(_zz_3111_)begin
        int_reg_array_44_56_imag <= _zz_3121_;
      end
      if(_zz_3112_)begin
        int_reg_array_44_57_imag <= _zz_3121_;
      end
      if(_zz_3113_)begin
        int_reg_array_44_58_imag <= _zz_3121_;
      end
      if(_zz_3114_)begin
        int_reg_array_44_59_imag <= _zz_3121_;
      end
      if(_zz_3115_)begin
        int_reg_array_44_60_imag <= _zz_3121_;
      end
      if(_zz_3116_)begin
        int_reg_array_44_61_imag <= _zz_3121_;
      end
      if(_zz_3117_)begin
        int_reg_array_44_62_imag <= _zz_3121_;
      end
      if(_zz_3118_)begin
        int_reg_array_44_63_imag <= _zz_3121_;
      end
      if(_zz_3124_)begin
        int_reg_array_45_0_real <= _zz_3189_;
      end
      if(_zz_3125_)begin
        int_reg_array_45_1_real <= _zz_3189_;
      end
      if(_zz_3126_)begin
        int_reg_array_45_2_real <= _zz_3189_;
      end
      if(_zz_3127_)begin
        int_reg_array_45_3_real <= _zz_3189_;
      end
      if(_zz_3128_)begin
        int_reg_array_45_4_real <= _zz_3189_;
      end
      if(_zz_3129_)begin
        int_reg_array_45_5_real <= _zz_3189_;
      end
      if(_zz_3130_)begin
        int_reg_array_45_6_real <= _zz_3189_;
      end
      if(_zz_3131_)begin
        int_reg_array_45_7_real <= _zz_3189_;
      end
      if(_zz_3132_)begin
        int_reg_array_45_8_real <= _zz_3189_;
      end
      if(_zz_3133_)begin
        int_reg_array_45_9_real <= _zz_3189_;
      end
      if(_zz_3134_)begin
        int_reg_array_45_10_real <= _zz_3189_;
      end
      if(_zz_3135_)begin
        int_reg_array_45_11_real <= _zz_3189_;
      end
      if(_zz_3136_)begin
        int_reg_array_45_12_real <= _zz_3189_;
      end
      if(_zz_3137_)begin
        int_reg_array_45_13_real <= _zz_3189_;
      end
      if(_zz_3138_)begin
        int_reg_array_45_14_real <= _zz_3189_;
      end
      if(_zz_3139_)begin
        int_reg_array_45_15_real <= _zz_3189_;
      end
      if(_zz_3140_)begin
        int_reg_array_45_16_real <= _zz_3189_;
      end
      if(_zz_3141_)begin
        int_reg_array_45_17_real <= _zz_3189_;
      end
      if(_zz_3142_)begin
        int_reg_array_45_18_real <= _zz_3189_;
      end
      if(_zz_3143_)begin
        int_reg_array_45_19_real <= _zz_3189_;
      end
      if(_zz_3144_)begin
        int_reg_array_45_20_real <= _zz_3189_;
      end
      if(_zz_3145_)begin
        int_reg_array_45_21_real <= _zz_3189_;
      end
      if(_zz_3146_)begin
        int_reg_array_45_22_real <= _zz_3189_;
      end
      if(_zz_3147_)begin
        int_reg_array_45_23_real <= _zz_3189_;
      end
      if(_zz_3148_)begin
        int_reg_array_45_24_real <= _zz_3189_;
      end
      if(_zz_3149_)begin
        int_reg_array_45_25_real <= _zz_3189_;
      end
      if(_zz_3150_)begin
        int_reg_array_45_26_real <= _zz_3189_;
      end
      if(_zz_3151_)begin
        int_reg_array_45_27_real <= _zz_3189_;
      end
      if(_zz_3152_)begin
        int_reg_array_45_28_real <= _zz_3189_;
      end
      if(_zz_3153_)begin
        int_reg_array_45_29_real <= _zz_3189_;
      end
      if(_zz_3154_)begin
        int_reg_array_45_30_real <= _zz_3189_;
      end
      if(_zz_3155_)begin
        int_reg_array_45_31_real <= _zz_3189_;
      end
      if(_zz_3156_)begin
        int_reg_array_45_32_real <= _zz_3189_;
      end
      if(_zz_3157_)begin
        int_reg_array_45_33_real <= _zz_3189_;
      end
      if(_zz_3158_)begin
        int_reg_array_45_34_real <= _zz_3189_;
      end
      if(_zz_3159_)begin
        int_reg_array_45_35_real <= _zz_3189_;
      end
      if(_zz_3160_)begin
        int_reg_array_45_36_real <= _zz_3189_;
      end
      if(_zz_3161_)begin
        int_reg_array_45_37_real <= _zz_3189_;
      end
      if(_zz_3162_)begin
        int_reg_array_45_38_real <= _zz_3189_;
      end
      if(_zz_3163_)begin
        int_reg_array_45_39_real <= _zz_3189_;
      end
      if(_zz_3164_)begin
        int_reg_array_45_40_real <= _zz_3189_;
      end
      if(_zz_3165_)begin
        int_reg_array_45_41_real <= _zz_3189_;
      end
      if(_zz_3166_)begin
        int_reg_array_45_42_real <= _zz_3189_;
      end
      if(_zz_3167_)begin
        int_reg_array_45_43_real <= _zz_3189_;
      end
      if(_zz_3168_)begin
        int_reg_array_45_44_real <= _zz_3189_;
      end
      if(_zz_3169_)begin
        int_reg_array_45_45_real <= _zz_3189_;
      end
      if(_zz_3170_)begin
        int_reg_array_45_46_real <= _zz_3189_;
      end
      if(_zz_3171_)begin
        int_reg_array_45_47_real <= _zz_3189_;
      end
      if(_zz_3172_)begin
        int_reg_array_45_48_real <= _zz_3189_;
      end
      if(_zz_3173_)begin
        int_reg_array_45_49_real <= _zz_3189_;
      end
      if(_zz_3174_)begin
        int_reg_array_45_50_real <= _zz_3189_;
      end
      if(_zz_3175_)begin
        int_reg_array_45_51_real <= _zz_3189_;
      end
      if(_zz_3176_)begin
        int_reg_array_45_52_real <= _zz_3189_;
      end
      if(_zz_3177_)begin
        int_reg_array_45_53_real <= _zz_3189_;
      end
      if(_zz_3178_)begin
        int_reg_array_45_54_real <= _zz_3189_;
      end
      if(_zz_3179_)begin
        int_reg_array_45_55_real <= _zz_3189_;
      end
      if(_zz_3180_)begin
        int_reg_array_45_56_real <= _zz_3189_;
      end
      if(_zz_3181_)begin
        int_reg_array_45_57_real <= _zz_3189_;
      end
      if(_zz_3182_)begin
        int_reg_array_45_58_real <= _zz_3189_;
      end
      if(_zz_3183_)begin
        int_reg_array_45_59_real <= _zz_3189_;
      end
      if(_zz_3184_)begin
        int_reg_array_45_60_real <= _zz_3189_;
      end
      if(_zz_3185_)begin
        int_reg_array_45_61_real <= _zz_3189_;
      end
      if(_zz_3186_)begin
        int_reg_array_45_62_real <= _zz_3189_;
      end
      if(_zz_3187_)begin
        int_reg_array_45_63_real <= _zz_3189_;
      end
      if(_zz_3124_)begin
        int_reg_array_45_0_imag <= _zz_3190_;
      end
      if(_zz_3125_)begin
        int_reg_array_45_1_imag <= _zz_3190_;
      end
      if(_zz_3126_)begin
        int_reg_array_45_2_imag <= _zz_3190_;
      end
      if(_zz_3127_)begin
        int_reg_array_45_3_imag <= _zz_3190_;
      end
      if(_zz_3128_)begin
        int_reg_array_45_4_imag <= _zz_3190_;
      end
      if(_zz_3129_)begin
        int_reg_array_45_5_imag <= _zz_3190_;
      end
      if(_zz_3130_)begin
        int_reg_array_45_6_imag <= _zz_3190_;
      end
      if(_zz_3131_)begin
        int_reg_array_45_7_imag <= _zz_3190_;
      end
      if(_zz_3132_)begin
        int_reg_array_45_8_imag <= _zz_3190_;
      end
      if(_zz_3133_)begin
        int_reg_array_45_9_imag <= _zz_3190_;
      end
      if(_zz_3134_)begin
        int_reg_array_45_10_imag <= _zz_3190_;
      end
      if(_zz_3135_)begin
        int_reg_array_45_11_imag <= _zz_3190_;
      end
      if(_zz_3136_)begin
        int_reg_array_45_12_imag <= _zz_3190_;
      end
      if(_zz_3137_)begin
        int_reg_array_45_13_imag <= _zz_3190_;
      end
      if(_zz_3138_)begin
        int_reg_array_45_14_imag <= _zz_3190_;
      end
      if(_zz_3139_)begin
        int_reg_array_45_15_imag <= _zz_3190_;
      end
      if(_zz_3140_)begin
        int_reg_array_45_16_imag <= _zz_3190_;
      end
      if(_zz_3141_)begin
        int_reg_array_45_17_imag <= _zz_3190_;
      end
      if(_zz_3142_)begin
        int_reg_array_45_18_imag <= _zz_3190_;
      end
      if(_zz_3143_)begin
        int_reg_array_45_19_imag <= _zz_3190_;
      end
      if(_zz_3144_)begin
        int_reg_array_45_20_imag <= _zz_3190_;
      end
      if(_zz_3145_)begin
        int_reg_array_45_21_imag <= _zz_3190_;
      end
      if(_zz_3146_)begin
        int_reg_array_45_22_imag <= _zz_3190_;
      end
      if(_zz_3147_)begin
        int_reg_array_45_23_imag <= _zz_3190_;
      end
      if(_zz_3148_)begin
        int_reg_array_45_24_imag <= _zz_3190_;
      end
      if(_zz_3149_)begin
        int_reg_array_45_25_imag <= _zz_3190_;
      end
      if(_zz_3150_)begin
        int_reg_array_45_26_imag <= _zz_3190_;
      end
      if(_zz_3151_)begin
        int_reg_array_45_27_imag <= _zz_3190_;
      end
      if(_zz_3152_)begin
        int_reg_array_45_28_imag <= _zz_3190_;
      end
      if(_zz_3153_)begin
        int_reg_array_45_29_imag <= _zz_3190_;
      end
      if(_zz_3154_)begin
        int_reg_array_45_30_imag <= _zz_3190_;
      end
      if(_zz_3155_)begin
        int_reg_array_45_31_imag <= _zz_3190_;
      end
      if(_zz_3156_)begin
        int_reg_array_45_32_imag <= _zz_3190_;
      end
      if(_zz_3157_)begin
        int_reg_array_45_33_imag <= _zz_3190_;
      end
      if(_zz_3158_)begin
        int_reg_array_45_34_imag <= _zz_3190_;
      end
      if(_zz_3159_)begin
        int_reg_array_45_35_imag <= _zz_3190_;
      end
      if(_zz_3160_)begin
        int_reg_array_45_36_imag <= _zz_3190_;
      end
      if(_zz_3161_)begin
        int_reg_array_45_37_imag <= _zz_3190_;
      end
      if(_zz_3162_)begin
        int_reg_array_45_38_imag <= _zz_3190_;
      end
      if(_zz_3163_)begin
        int_reg_array_45_39_imag <= _zz_3190_;
      end
      if(_zz_3164_)begin
        int_reg_array_45_40_imag <= _zz_3190_;
      end
      if(_zz_3165_)begin
        int_reg_array_45_41_imag <= _zz_3190_;
      end
      if(_zz_3166_)begin
        int_reg_array_45_42_imag <= _zz_3190_;
      end
      if(_zz_3167_)begin
        int_reg_array_45_43_imag <= _zz_3190_;
      end
      if(_zz_3168_)begin
        int_reg_array_45_44_imag <= _zz_3190_;
      end
      if(_zz_3169_)begin
        int_reg_array_45_45_imag <= _zz_3190_;
      end
      if(_zz_3170_)begin
        int_reg_array_45_46_imag <= _zz_3190_;
      end
      if(_zz_3171_)begin
        int_reg_array_45_47_imag <= _zz_3190_;
      end
      if(_zz_3172_)begin
        int_reg_array_45_48_imag <= _zz_3190_;
      end
      if(_zz_3173_)begin
        int_reg_array_45_49_imag <= _zz_3190_;
      end
      if(_zz_3174_)begin
        int_reg_array_45_50_imag <= _zz_3190_;
      end
      if(_zz_3175_)begin
        int_reg_array_45_51_imag <= _zz_3190_;
      end
      if(_zz_3176_)begin
        int_reg_array_45_52_imag <= _zz_3190_;
      end
      if(_zz_3177_)begin
        int_reg_array_45_53_imag <= _zz_3190_;
      end
      if(_zz_3178_)begin
        int_reg_array_45_54_imag <= _zz_3190_;
      end
      if(_zz_3179_)begin
        int_reg_array_45_55_imag <= _zz_3190_;
      end
      if(_zz_3180_)begin
        int_reg_array_45_56_imag <= _zz_3190_;
      end
      if(_zz_3181_)begin
        int_reg_array_45_57_imag <= _zz_3190_;
      end
      if(_zz_3182_)begin
        int_reg_array_45_58_imag <= _zz_3190_;
      end
      if(_zz_3183_)begin
        int_reg_array_45_59_imag <= _zz_3190_;
      end
      if(_zz_3184_)begin
        int_reg_array_45_60_imag <= _zz_3190_;
      end
      if(_zz_3185_)begin
        int_reg_array_45_61_imag <= _zz_3190_;
      end
      if(_zz_3186_)begin
        int_reg_array_45_62_imag <= _zz_3190_;
      end
      if(_zz_3187_)begin
        int_reg_array_45_63_imag <= _zz_3190_;
      end
      if(_zz_3193_)begin
        int_reg_array_46_0_real <= _zz_3258_;
      end
      if(_zz_3194_)begin
        int_reg_array_46_1_real <= _zz_3258_;
      end
      if(_zz_3195_)begin
        int_reg_array_46_2_real <= _zz_3258_;
      end
      if(_zz_3196_)begin
        int_reg_array_46_3_real <= _zz_3258_;
      end
      if(_zz_3197_)begin
        int_reg_array_46_4_real <= _zz_3258_;
      end
      if(_zz_3198_)begin
        int_reg_array_46_5_real <= _zz_3258_;
      end
      if(_zz_3199_)begin
        int_reg_array_46_6_real <= _zz_3258_;
      end
      if(_zz_3200_)begin
        int_reg_array_46_7_real <= _zz_3258_;
      end
      if(_zz_3201_)begin
        int_reg_array_46_8_real <= _zz_3258_;
      end
      if(_zz_3202_)begin
        int_reg_array_46_9_real <= _zz_3258_;
      end
      if(_zz_3203_)begin
        int_reg_array_46_10_real <= _zz_3258_;
      end
      if(_zz_3204_)begin
        int_reg_array_46_11_real <= _zz_3258_;
      end
      if(_zz_3205_)begin
        int_reg_array_46_12_real <= _zz_3258_;
      end
      if(_zz_3206_)begin
        int_reg_array_46_13_real <= _zz_3258_;
      end
      if(_zz_3207_)begin
        int_reg_array_46_14_real <= _zz_3258_;
      end
      if(_zz_3208_)begin
        int_reg_array_46_15_real <= _zz_3258_;
      end
      if(_zz_3209_)begin
        int_reg_array_46_16_real <= _zz_3258_;
      end
      if(_zz_3210_)begin
        int_reg_array_46_17_real <= _zz_3258_;
      end
      if(_zz_3211_)begin
        int_reg_array_46_18_real <= _zz_3258_;
      end
      if(_zz_3212_)begin
        int_reg_array_46_19_real <= _zz_3258_;
      end
      if(_zz_3213_)begin
        int_reg_array_46_20_real <= _zz_3258_;
      end
      if(_zz_3214_)begin
        int_reg_array_46_21_real <= _zz_3258_;
      end
      if(_zz_3215_)begin
        int_reg_array_46_22_real <= _zz_3258_;
      end
      if(_zz_3216_)begin
        int_reg_array_46_23_real <= _zz_3258_;
      end
      if(_zz_3217_)begin
        int_reg_array_46_24_real <= _zz_3258_;
      end
      if(_zz_3218_)begin
        int_reg_array_46_25_real <= _zz_3258_;
      end
      if(_zz_3219_)begin
        int_reg_array_46_26_real <= _zz_3258_;
      end
      if(_zz_3220_)begin
        int_reg_array_46_27_real <= _zz_3258_;
      end
      if(_zz_3221_)begin
        int_reg_array_46_28_real <= _zz_3258_;
      end
      if(_zz_3222_)begin
        int_reg_array_46_29_real <= _zz_3258_;
      end
      if(_zz_3223_)begin
        int_reg_array_46_30_real <= _zz_3258_;
      end
      if(_zz_3224_)begin
        int_reg_array_46_31_real <= _zz_3258_;
      end
      if(_zz_3225_)begin
        int_reg_array_46_32_real <= _zz_3258_;
      end
      if(_zz_3226_)begin
        int_reg_array_46_33_real <= _zz_3258_;
      end
      if(_zz_3227_)begin
        int_reg_array_46_34_real <= _zz_3258_;
      end
      if(_zz_3228_)begin
        int_reg_array_46_35_real <= _zz_3258_;
      end
      if(_zz_3229_)begin
        int_reg_array_46_36_real <= _zz_3258_;
      end
      if(_zz_3230_)begin
        int_reg_array_46_37_real <= _zz_3258_;
      end
      if(_zz_3231_)begin
        int_reg_array_46_38_real <= _zz_3258_;
      end
      if(_zz_3232_)begin
        int_reg_array_46_39_real <= _zz_3258_;
      end
      if(_zz_3233_)begin
        int_reg_array_46_40_real <= _zz_3258_;
      end
      if(_zz_3234_)begin
        int_reg_array_46_41_real <= _zz_3258_;
      end
      if(_zz_3235_)begin
        int_reg_array_46_42_real <= _zz_3258_;
      end
      if(_zz_3236_)begin
        int_reg_array_46_43_real <= _zz_3258_;
      end
      if(_zz_3237_)begin
        int_reg_array_46_44_real <= _zz_3258_;
      end
      if(_zz_3238_)begin
        int_reg_array_46_45_real <= _zz_3258_;
      end
      if(_zz_3239_)begin
        int_reg_array_46_46_real <= _zz_3258_;
      end
      if(_zz_3240_)begin
        int_reg_array_46_47_real <= _zz_3258_;
      end
      if(_zz_3241_)begin
        int_reg_array_46_48_real <= _zz_3258_;
      end
      if(_zz_3242_)begin
        int_reg_array_46_49_real <= _zz_3258_;
      end
      if(_zz_3243_)begin
        int_reg_array_46_50_real <= _zz_3258_;
      end
      if(_zz_3244_)begin
        int_reg_array_46_51_real <= _zz_3258_;
      end
      if(_zz_3245_)begin
        int_reg_array_46_52_real <= _zz_3258_;
      end
      if(_zz_3246_)begin
        int_reg_array_46_53_real <= _zz_3258_;
      end
      if(_zz_3247_)begin
        int_reg_array_46_54_real <= _zz_3258_;
      end
      if(_zz_3248_)begin
        int_reg_array_46_55_real <= _zz_3258_;
      end
      if(_zz_3249_)begin
        int_reg_array_46_56_real <= _zz_3258_;
      end
      if(_zz_3250_)begin
        int_reg_array_46_57_real <= _zz_3258_;
      end
      if(_zz_3251_)begin
        int_reg_array_46_58_real <= _zz_3258_;
      end
      if(_zz_3252_)begin
        int_reg_array_46_59_real <= _zz_3258_;
      end
      if(_zz_3253_)begin
        int_reg_array_46_60_real <= _zz_3258_;
      end
      if(_zz_3254_)begin
        int_reg_array_46_61_real <= _zz_3258_;
      end
      if(_zz_3255_)begin
        int_reg_array_46_62_real <= _zz_3258_;
      end
      if(_zz_3256_)begin
        int_reg_array_46_63_real <= _zz_3258_;
      end
      if(_zz_3193_)begin
        int_reg_array_46_0_imag <= _zz_3259_;
      end
      if(_zz_3194_)begin
        int_reg_array_46_1_imag <= _zz_3259_;
      end
      if(_zz_3195_)begin
        int_reg_array_46_2_imag <= _zz_3259_;
      end
      if(_zz_3196_)begin
        int_reg_array_46_3_imag <= _zz_3259_;
      end
      if(_zz_3197_)begin
        int_reg_array_46_4_imag <= _zz_3259_;
      end
      if(_zz_3198_)begin
        int_reg_array_46_5_imag <= _zz_3259_;
      end
      if(_zz_3199_)begin
        int_reg_array_46_6_imag <= _zz_3259_;
      end
      if(_zz_3200_)begin
        int_reg_array_46_7_imag <= _zz_3259_;
      end
      if(_zz_3201_)begin
        int_reg_array_46_8_imag <= _zz_3259_;
      end
      if(_zz_3202_)begin
        int_reg_array_46_9_imag <= _zz_3259_;
      end
      if(_zz_3203_)begin
        int_reg_array_46_10_imag <= _zz_3259_;
      end
      if(_zz_3204_)begin
        int_reg_array_46_11_imag <= _zz_3259_;
      end
      if(_zz_3205_)begin
        int_reg_array_46_12_imag <= _zz_3259_;
      end
      if(_zz_3206_)begin
        int_reg_array_46_13_imag <= _zz_3259_;
      end
      if(_zz_3207_)begin
        int_reg_array_46_14_imag <= _zz_3259_;
      end
      if(_zz_3208_)begin
        int_reg_array_46_15_imag <= _zz_3259_;
      end
      if(_zz_3209_)begin
        int_reg_array_46_16_imag <= _zz_3259_;
      end
      if(_zz_3210_)begin
        int_reg_array_46_17_imag <= _zz_3259_;
      end
      if(_zz_3211_)begin
        int_reg_array_46_18_imag <= _zz_3259_;
      end
      if(_zz_3212_)begin
        int_reg_array_46_19_imag <= _zz_3259_;
      end
      if(_zz_3213_)begin
        int_reg_array_46_20_imag <= _zz_3259_;
      end
      if(_zz_3214_)begin
        int_reg_array_46_21_imag <= _zz_3259_;
      end
      if(_zz_3215_)begin
        int_reg_array_46_22_imag <= _zz_3259_;
      end
      if(_zz_3216_)begin
        int_reg_array_46_23_imag <= _zz_3259_;
      end
      if(_zz_3217_)begin
        int_reg_array_46_24_imag <= _zz_3259_;
      end
      if(_zz_3218_)begin
        int_reg_array_46_25_imag <= _zz_3259_;
      end
      if(_zz_3219_)begin
        int_reg_array_46_26_imag <= _zz_3259_;
      end
      if(_zz_3220_)begin
        int_reg_array_46_27_imag <= _zz_3259_;
      end
      if(_zz_3221_)begin
        int_reg_array_46_28_imag <= _zz_3259_;
      end
      if(_zz_3222_)begin
        int_reg_array_46_29_imag <= _zz_3259_;
      end
      if(_zz_3223_)begin
        int_reg_array_46_30_imag <= _zz_3259_;
      end
      if(_zz_3224_)begin
        int_reg_array_46_31_imag <= _zz_3259_;
      end
      if(_zz_3225_)begin
        int_reg_array_46_32_imag <= _zz_3259_;
      end
      if(_zz_3226_)begin
        int_reg_array_46_33_imag <= _zz_3259_;
      end
      if(_zz_3227_)begin
        int_reg_array_46_34_imag <= _zz_3259_;
      end
      if(_zz_3228_)begin
        int_reg_array_46_35_imag <= _zz_3259_;
      end
      if(_zz_3229_)begin
        int_reg_array_46_36_imag <= _zz_3259_;
      end
      if(_zz_3230_)begin
        int_reg_array_46_37_imag <= _zz_3259_;
      end
      if(_zz_3231_)begin
        int_reg_array_46_38_imag <= _zz_3259_;
      end
      if(_zz_3232_)begin
        int_reg_array_46_39_imag <= _zz_3259_;
      end
      if(_zz_3233_)begin
        int_reg_array_46_40_imag <= _zz_3259_;
      end
      if(_zz_3234_)begin
        int_reg_array_46_41_imag <= _zz_3259_;
      end
      if(_zz_3235_)begin
        int_reg_array_46_42_imag <= _zz_3259_;
      end
      if(_zz_3236_)begin
        int_reg_array_46_43_imag <= _zz_3259_;
      end
      if(_zz_3237_)begin
        int_reg_array_46_44_imag <= _zz_3259_;
      end
      if(_zz_3238_)begin
        int_reg_array_46_45_imag <= _zz_3259_;
      end
      if(_zz_3239_)begin
        int_reg_array_46_46_imag <= _zz_3259_;
      end
      if(_zz_3240_)begin
        int_reg_array_46_47_imag <= _zz_3259_;
      end
      if(_zz_3241_)begin
        int_reg_array_46_48_imag <= _zz_3259_;
      end
      if(_zz_3242_)begin
        int_reg_array_46_49_imag <= _zz_3259_;
      end
      if(_zz_3243_)begin
        int_reg_array_46_50_imag <= _zz_3259_;
      end
      if(_zz_3244_)begin
        int_reg_array_46_51_imag <= _zz_3259_;
      end
      if(_zz_3245_)begin
        int_reg_array_46_52_imag <= _zz_3259_;
      end
      if(_zz_3246_)begin
        int_reg_array_46_53_imag <= _zz_3259_;
      end
      if(_zz_3247_)begin
        int_reg_array_46_54_imag <= _zz_3259_;
      end
      if(_zz_3248_)begin
        int_reg_array_46_55_imag <= _zz_3259_;
      end
      if(_zz_3249_)begin
        int_reg_array_46_56_imag <= _zz_3259_;
      end
      if(_zz_3250_)begin
        int_reg_array_46_57_imag <= _zz_3259_;
      end
      if(_zz_3251_)begin
        int_reg_array_46_58_imag <= _zz_3259_;
      end
      if(_zz_3252_)begin
        int_reg_array_46_59_imag <= _zz_3259_;
      end
      if(_zz_3253_)begin
        int_reg_array_46_60_imag <= _zz_3259_;
      end
      if(_zz_3254_)begin
        int_reg_array_46_61_imag <= _zz_3259_;
      end
      if(_zz_3255_)begin
        int_reg_array_46_62_imag <= _zz_3259_;
      end
      if(_zz_3256_)begin
        int_reg_array_46_63_imag <= _zz_3259_;
      end
      if(_zz_3262_)begin
        int_reg_array_47_0_real <= _zz_3327_;
      end
      if(_zz_3263_)begin
        int_reg_array_47_1_real <= _zz_3327_;
      end
      if(_zz_3264_)begin
        int_reg_array_47_2_real <= _zz_3327_;
      end
      if(_zz_3265_)begin
        int_reg_array_47_3_real <= _zz_3327_;
      end
      if(_zz_3266_)begin
        int_reg_array_47_4_real <= _zz_3327_;
      end
      if(_zz_3267_)begin
        int_reg_array_47_5_real <= _zz_3327_;
      end
      if(_zz_3268_)begin
        int_reg_array_47_6_real <= _zz_3327_;
      end
      if(_zz_3269_)begin
        int_reg_array_47_7_real <= _zz_3327_;
      end
      if(_zz_3270_)begin
        int_reg_array_47_8_real <= _zz_3327_;
      end
      if(_zz_3271_)begin
        int_reg_array_47_9_real <= _zz_3327_;
      end
      if(_zz_3272_)begin
        int_reg_array_47_10_real <= _zz_3327_;
      end
      if(_zz_3273_)begin
        int_reg_array_47_11_real <= _zz_3327_;
      end
      if(_zz_3274_)begin
        int_reg_array_47_12_real <= _zz_3327_;
      end
      if(_zz_3275_)begin
        int_reg_array_47_13_real <= _zz_3327_;
      end
      if(_zz_3276_)begin
        int_reg_array_47_14_real <= _zz_3327_;
      end
      if(_zz_3277_)begin
        int_reg_array_47_15_real <= _zz_3327_;
      end
      if(_zz_3278_)begin
        int_reg_array_47_16_real <= _zz_3327_;
      end
      if(_zz_3279_)begin
        int_reg_array_47_17_real <= _zz_3327_;
      end
      if(_zz_3280_)begin
        int_reg_array_47_18_real <= _zz_3327_;
      end
      if(_zz_3281_)begin
        int_reg_array_47_19_real <= _zz_3327_;
      end
      if(_zz_3282_)begin
        int_reg_array_47_20_real <= _zz_3327_;
      end
      if(_zz_3283_)begin
        int_reg_array_47_21_real <= _zz_3327_;
      end
      if(_zz_3284_)begin
        int_reg_array_47_22_real <= _zz_3327_;
      end
      if(_zz_3285_)begin
        int_reg_array_47_23_real <= _zz_3327_;
      end
      if(_zz_3286_)begin
        int_reg_array_47_24_real <= _zz_3327_;
      end
      if(_zz_3287_)begin
        int_reg_array_47_25_real <= _zz_3327_;
      end
      if(_zz_3288_)begin
        int_reg_array_47_26_real <= _zz_3327_;
      end
      if(_zz_3289_)begin
        int_reg_array_47_27_real <= _zz_3327_;
      end
      if(_zz_3290_)begin
        int_reg_array_47_28_real <= _zz_3327_;
      end
      if(_zz_3291_)begin
        int_reg_array_47_29_real <= _zz_3327_;
      end
      if(_zz_3292_)begin
        int_reg_array_47_30_real <= _zz_3327_;
      end
      if(_zz_3293_)begin
        int_reg_array_47_31_real <= _zz_3327_;
      end
      if(_zz_3294_)begin
        int_reg_array_47_32_real <= _zz_3327_;
      end
      if(_zz_3295_)begin
        int_reg_array_47_33_real <= _zz_3327_;
      end
      if(_zz_3296_)begin
        int_reg_array_47_34_real <= _zz_3327_;
      end
      if(_zz_3297_)begin
        int_reg_array_47_35_real <= _zz_3327_;
      end
      if(_zz_3298_)begin
        int_reg_array_47_36_real <= _zz_3327_;
      end
      if(_zz_3299_)begin
        int_reg_array_47_37_real <= _zz_3327_;
      end
      if(_zz_3300_)begin
        int_reg_array_47_38_real <= _zz_3327_;
      end
      if(_zz_3301_)begin
        int_reg_array_47_39_real <= _zz_3327_;
      end
      if(_zz_3302_)begin
        int_reg_array_47_40_real <= _zz_3327_;
      end
      if(_zz_3303_)begin
        int_reg_array_47_41_real <= _zz_3327_;
      end
      if(_zz_3304_)begin
        int_reg_array_47_42_real <= _zz_3327_;
      end
      if(_zz_3305_)begin
        int_reg_array_47_43_real <= _zz_3327_;
      end
      if(_zz_3306_)begin
        int_reg_array_47_44_real <= _zz_3327_;
      end
      if(_zz_3307_)begin
        int_reg_array_47_45_real <= _zz_3327_;
      end
      if(_zz_3308_)begin
        int_reg_array_47_46_real <= _zz_3327_;
      end
      if(_zz_3309_)begin
        int_reg_array_47_47_real <= _zz_3327_;
      end
      if(_zz_3310_)begin
        int_reg_array_47_48_real <= _zz_3327_;
      end
      if(_zz_3311_)begin
        int_reg_array_47_49_real <= _zz_3327_;
      end
      if(_zz_3312_)begin
        int_reg_array_47_50_real <= _zz_3327_;
      end
      if(_zz_3313_)begin
        int_reg_array_47_51_real <= _zz_3327_;
      end
      if(_zz_3314_)begin
        int_reg_array_47_52_real <= _zz_3327_;
      end
      if(_zz_3315_)begin
        int_reg_array_47_53_real <= _zz_3327_;
      end
      if(_zz_3316_)begin
        int_reg_array_47_54_real <= _zz_3327_;
      end
      if(_zz_3317_)begin
        int_reg_array_47_55_real <= _zz_3327_;
      end
      if(_zz_3318_)begin
        int_reg_array_47_56_real <= _zz_3327_;
      end
      if(_zz_3319_)begin
        int_reg_array_47_57_real <= _zz_3327_;
      end
      if(_zz_3320_)begin
        int_reg_array_47_58_real <= _zz_3327_;
      end
      if(_zz_3321_)begin
        int_reg_array_47_59_real <= _zz_3327_;
      end
      if(_zz_3322_)begin
        int_reg_array_47_60_real <= _zz_3327_;
      end
      if(_zz_3323_)begin
        int_reg_array_47_61_real <= _zz_3327_;
      end
      if(_zz_3324_)begin
        int_reg_array_47_62_real <= _zz_3327_;
      end
      if(_zz_3325_)begin
        int_reg_array_47_63_real <= _zz_3327_;
      end
      if(_zz_3262_)begin
        int_reg_array_47_0_imag <= _zz_3328_;
      end
      if(_zz_3263_)begin
        int_reg_array_47_1_imag <= _zz_3328_;
      end
      if(_zz_3264_)begin
        int_reg_array_47_2_imag <= _zz_3328_;
      end
      if(_zz_3265_)begin
        int_reg_array_47_3_imag <= _zz_3328_;
      end
      if(_zz_3266_)begin
        int_reg_array_47_4_imag <= _zz_3328_;
      end
      if(_zz_3267_)begin
        int_reg_array_47_5_imag <= _zz_3328_;
      end
      if(_zz_3268_)begin
        int_reg_array_47_6_imag <= _zz_3328_;
      end
      if(_zz_3269_)begin
        int_reg_array_47_7_imag <= _zz_3328_;
      end
      if(_zz_3270_)begin
        int_reg_array_47_8_imag <= _zz_3328_;
      end
      if(_zz_3271_)begin
        int_reg_array_47_9_imag <= _zz_3328_;
      end
      if(_zz_3272_)begin
        int_reg_array_47_10_imag <= _zz_3328_;
      end
      if(_zz_3273_)begin
        int_reg_array_47_11_imag <= _zz_3328_;
      end
      if(_zz_3274_)begin
        int_reg_array_47_12_imag <= _zz_3328_;
      end
      if(_zz_3275_)begin
        int_reg_array_47_13_imag <= _zz_3328_;
      end
      if(_zz_3276_)begin
        int_reg_array_47_14_imag <= _zz_3328_;
      end
      if(_zz_3277_)begin
        int_reg_array_47_15_imag <= _zz_3328_;
      end
      if(_zz_3278_)begin
        int_reg_array_47_16_imag <= _zz_3328_;
      end
      if(_zz_3279_)begin
        int_reg_array_47_17_imag <= _zz_3328_;
      end
      if(_zz_3280_)begin
        int_reg_array_47_18_imag <= _zz_3328_;
      end
      if(_zz_3281_)begin
        int_reg_array_47_19_imag <= _zz_3328_;
      end
      if(_zz_3282_)begin
        int_reg_array_47_20_imag <= _zz_3328_;
      end
      if(_zz_3283_)begin
        int_reg_array_47_21_imag <= _zz_3328_;
      end
      if(_zz_3284_)begin
        int_reg_array_47_22_imag <= _zz_3328_;
      end
      if(_zz_3285_)begin
        int_reg_array_47_23_imag <= _zz_3328_;
      end
      if(_zz_3286_)begin
        int_reg_array_47_24_imag <= _zz_3328_;
      end
      if(_zz_3287_)begin
        int_reg_array_47_25_imag <= _zz_3328_;
      end
      if(_zz_3288_)begin
        int_reg_array_47_26_imag <= _zz_3328_;
      end
      if(_zz_3289_)begin
        int_reg_array_47_27_imag <= _zz_3328_;
      end
      if(_zz_3290_)begin
        int_reg_array_47_28_imag <= _zz_3328_;
      end
      if(_zz_3291_)begin
        int_reg_array_47_29_imag <= _zz_3328_;
      end
      if(_zz_3292_)begin
        int_reg_array_47_30_imag <= _zz_3328_;
      end
      if(_zz_3293_)begin
        int_reg_array_47_31_imag <= _zz_3328_;
      end
      if(_zz_3294_)begin
        int_reg_array_47_32_imag <= _zz_3328_;
      end
      if(_zz_3295_)begin
        int_reg_array_47_33_imag <= _zz_3328_;
      end
      if(_zz_3296_)begin
        int_reg_array_47_34_imag <= _zz_3328_;
      end
      if(_zz_3297_)begin
        int_reg_array_47_35_imag <= _zz_3328_;
      end
      if(_zz_3298_)begin
        int_reg_array_47_36_imag <= _zz_3328_;
      end
      if(_zz_3299_)begin
        int_reg_array_47_37_imag <= _zz_3328_;
      end
      if(_zz_3300_)begin
        int_reg_array_47_38_imag <= _zz_3328_;
      end
      if(_zz_3301_)begin
        int_reg_array_47_39_imag <= _zz_3328_;
      end
      if(_zz_3302_)begin
        int_reg_array_47_40_imag <= _zz_3328_;
      end
      if(_zz_3303_)begin
        int_reg_array_47_41_imag <= _zz_3328_;
      end
      if(_zz_3304_)begin
        int_reg_array_47_42_imag <= _zz_3328_;
      end
      if(_zz_3305_)begin
        int_reg_array_47_43_imag <= _zz_3328_;
      end
      if(_zz_3306_)begin
        int_reg_array_47_44_imag <= _zz_3328_;
      end
      if(_zz_3307_)begin
        int_reg_array_47_45_imag <= _zz_3328_;
      end
      if(_zz_3308_)begin
        int_reg_array_47_46_imag <= _zz_3328_;
      end
      if(_zz_3309_)begin
        int_reg_array_47_47_imag <= _zz_3328_;
      end
      if(_zz_3310_)begin
        int_reg_array_47_48_imag <= _zz_3328_;
      end
      if(_zz_3311_)begin
        int_reg_array_47_49_imag <= _zz_3328_;
      end
      if(_zz_3312_)begin
        int_reg_array_47_50_imag <= _zz_3328_;
      end
      if(_zz_3313_)begin
        int_reg_array_47_51_imag <= _zz_3328_;
      end
      if(_zz_3314_)begin
        int_reg_array_47_52_imag <= _zz_3328_;
      end
      if(_zz_3315_)begin
        int_reg_array_47_53_imag <= _zz_3328_;
      end
      if(_zz_3316_)begin
        int_reg_array_47_54_imag <= _zz_3328_;
      end
      if(_zz_3317_)begin
        int_reg_array_47_55_imag <= _zz_3328_;
      end
      if(_zz_3318_)begin
        int_reg_array_47_56_imag <= _zz_3328_;
      end
      if(_zz_3319_)begin
        int_reg_array_47_57_imag <= _zz_3328_;
      end
      if(_zz_3320_)begin
        int_reg_array_47_58_imag <= _zz_3328_;
      end
      if(_zz_3321_)begin
        int_reg_array_47_59_imag <= _zz_3328_;
      end
      if(_zz_3322_)begin
        int_reg_array_47_60_imag <= _zz_3328_;
      end
      if(_zz_3323_)begin
        int_reg_array_47_61_imag <= _zz_3328_;
      end
      if(_zz_3324_)begin
        int_reg_array_47_62_imag <= _zz_3328_;
      end
      if(_zz_3325_)begin
        int_reg_array_47_63_imag <= _zz_3328_;
      end
      if(_zz_3331_)begin
        int_reg_array_48_0_real <= _zz_3396_;
      end
      if(_zz_3332_)begin
        int_reg_array_48_1_real <= _zz_3396_;
      end
      if(_zz_3333_)begin
        int_reg_array_48_2_real <= _zz_3396_;
      end
      if(_zz_3334_)begin
        int_reg_array_48_3_real <= _zz_3396_;
      end
      if(_zz_3335_)begin
        int_reg_array_48_4_real <= _zz_3396_;
      end
      if(_zz_3336_)begin
        int_reg_array_48_5_real <= _zz_3396_;
      end
      if(_zz_3337_)begin
        int_reg_array_48_6_real <= _zz_3396_;
      end
      if(_zz_3338_)begin
        int_reg_array_48_7_real <= _zz_3396_;
      end
      if(_zz_3339_)begin
        int_reg_array_48_8_real <= _zz_3396_;
      end
      if(_zz_3340_)begin
        int_reg_array_48_9_real <= _zz_3396_;
      end
      if(_zz_3341_)begin
        int_reg_array_48_10_real <= _zz_3396_;
      end
      if(_zz_3342_)begin
        int_reg_array_48_11_real <= _zz_3396_;
      end
      if(_zz_3343_)begin
        int_reg_array_48_12_real <= _zz_3396_;
      end
      if(_zz_3344_)begin
        int_reg_array_48_13_real <= _zz_3396_;
      end
      if(_zz_3345_)begin
        int_reg_array_48_14_real <= _zz_3396_;
      end
      if(_zz_3346_)begin
        int_reg_array_48_15_real <= _zz_3396_;
      end
      if(_zz_3347_)begin
        int_reg_array_48_16_real <= _zz_3396_;
      end
      if(_zz_3348_)begin
        int_reg_array_48_17_real <= _zz_3396_;
      end
      if(_zz_3349_)begin
        int_reg_array_48_18_real <= _zz_3396_;
      end
      if(_zz_3350_)begin
        int_reg_array_48_19_real <= _zz_3396_;
      end
      if(_zz_3351_)begin
        int_reg_array_48_20_real <= _zz_3396_;
      end
      if(_zz_3352_)begin
        int_reg_array_48_21_real <= _zz_3396_;
      end
      if(_zz_3353_)begin
        int_reg_array_48_22_real <= _zz_3396_;
      end
      if(_zz_3354_)begin
        int_reg_array_48_23_real <= _zz_3396_;
      end
      if(_zz_3355_)begin
        int_reg_array_48_24_real <= _zz_3396_;
      end
      if(_zz_3356_)begin
        int_reg_array_48_25_real <= _zz_3396_;
      end
      if(_zz_3357_)begin
        int_reg_array_48_26_real <= _zz_3396_;
      end
      if(_zz_3358_)begin
        int_reg_array_48_27_real <= _zz_3396_;
      end
      if(_zz_3359_)begin
        int_reg_array_48_28_real <= _zz_3396_;
      end
      if(_zz_3360_)begin
        int_reg_array_48_29_real <= _zz_3396_;
      end
      if(_zz_3361_)begin
        int_reg_array_48_30_real <= _zz_3396_;
      end
      if(_zz_3362_)begin
        int_reg_array_48_31_real <= _zz_3396_;
      end
      if(_zz_3363_)begin
        int_reg_array_48_32_real <= _zz_3396_;
      end
      if(_zz_3364_)begin
        int_reg_array_48_33_real <= _zz_3396_;
      end
      if(_zz_3365_)begin
        int_reg_array_48_34_real <= _zz_3396_;
      end
      if(_zz_3366_)begin
        int_reg_array_48_35_real <= _zz_3396_;
      end
      if(_zz_3367_)begin
        int_reg_array_48_36_real <= _zz_3396_;
      end
      if(_zz_3368_)begin
        int_reg_array_48_37_real <= _zz_3396_;
      end
      if(_zz_3369_)begin
        int_reg_array_48_38_real <= _zz_3396_;
      end
      if(_zz_3370_)begin
        int_reg_array_48_39_real <= _zz_3396_;
      end
      if(_zz_3371_)begin
        int_reg_array_48_40_real <= _zz_3396_;
      end
      if(_zz_3372_)begin
        int_reg_array_48_41_real <= _zz_3396_;
      end
      if(_zz_3373_)begin
        int_reg_array_48_42_real <= _zz_3396_;
      end
      if(_zz_3374_)begin
        int_reg_array_48_43_real <= _zz_3396_;
      end
      if(_zz_3375_)begin
        int_reg_array_48_44_real <= _zz_3396_;
      end
      if(_zz_3376_)begin
        int_reg_array_48_45_real <= _zz_3396_;
      end
      if(_zz_3377_)begin
        int_reg_array_48_46_real <= _zz_3396_;
      end
      if(_zz_3378_)begin
        int_reg_array_48_47_real <= _zz_3396_;
      end
      if(_zz_3379_)begin
        int_reg_array_48_48_real <= _zz_3396_;
      end
      if(_zz_3380_)begin
        int_reg_array_48_49_real <= _zz_3396_;
      end
      if(_zz_3381_)begin
        int_reg_array_48_50_real <= _zz_3396_;
      end
      if(_zz_3382_)begin
        int_reg_array_48_51_real <= _zz_3396_;
      end
      if(_zz_3383_)begin
        int_reg_array_48_52_real <= _zz_3396_;
      end
      if(_zz_3384_)begin
        int_reg_array_48_53_real <= _zz_3396_;
      end
      if(_zz_3385_)begin
        int_reg_array_48_54_real <= _zz_3396_;
      end
      if(_zz_3386_)begin
        int_reg_array_48_55_real <= _zz_3396_;
      end
      if(_zz_3387_)begin
        int_reg_array_48_56_real <= _zz_3396_;
      end
      if(_zz_3388_)begin
        int_reg_array_48_57_real <= _zz_3396_;
      end
      if(_zz_3389_)begin
        int_reg_array_48_58_real <= _zz_3396_;
      end
      if(_zz_3390_)begin
        int_reg_array_48_59_real <= _zz_3396_;
      end
      if(_zz_3391_)begin
        int_reg_array_48_60_real <= _zz_3396_;
      end
      if(_zz_3392_)begin
        int_reg_array_48_61_real <= _zz_3396_;
      end
      if(_zz_3393_)begin
        int_reg_array_48_62_real <= _zz_3396_;
      end
      if(_zz_3394_)begin
        int_reg_array_48_63_real <= _zz_3396_;
      end
      if(_zz_3331_)begin
        int_reg_array_48_0_imag <= _zz_3397_;
      end
      if(_zz_3332_)begin
        int_reg_array_48_1_imag <= _zz_3397_;
      end
      if(_zz_3333_)begin
        int_reg_array_48_2_imag <= _zz_3397_;
      end
      if(_zz_3334_)begin
        int_reg_array_48_3_imag <= _zz_3397_;
      end
      if(_zz_3335_)begin
        int_reg_array_48_4_imag <= _zz_3397_;
      end
      if(_zz_3336_)begin
        int_reg_array_48_5_imag <= _zz_3397_;
      end
      if(_zz_3337_)begin
        int_reg_array_48_6_imag <= _zz_3397_;
      end
      if(_zz_3338_)begin
        int_reg_array_48_7_imag <= _zz_3397_;
      end
      if(_zz_3339_)begin
        int_reg_array_48_8_imag <= _zz_3397_;
      end
      if(_zz_3340_)begin
        int_reg_array_48_9_imag <= _zz_3397_;
      end
      if(_zz_3341_)begin
        int_reg_array_48_10_imag <= _zz_3397_;
      end
      if(_zz_3342_)begin
        int_reg_array_48_11_imag <= _zz_3397_;
      end
      if(_zz_3343_)begin
        int_reg_array_48_12_imag <= _zz_3397_;
      end
      if(_zz_3344_)begin
        int_reg_array_48_13_imag <= _zz_3397_;
      end
      if(_zz_3345_)begin
        int_reg_array_48_14_imag <= _zz_3397_;
      end
      if(_zz_3346_)begin
        int_reg_array_48_15_imag <= _zz_3397_;
      end
      if(_zz_3347_)begin
        int_reg_array_48_16_imag <= _zz_3397_;
      end
      if(_zz_3348_)begin
        int_reg_array_48_17_imag <= _zz_3397_;
      end
      if(_zz_3349_)begin
        int_reg_array_48_18_imag <= _zz_3397_;
      end
      if(_zz_3350_)begin
        int_reg_array_48_19_imag <= _zz_3397_;
      end
      if(_zz_3351_)begin
        int_reg_array_48_20_imag <= _zz_3397_;
      end
      if(_zz_3352_)begin
        int_reg_array_48_21_imag <= _zz_3397_;
      end
      if(_zz_3353_)begin
        int_reg_array_48_22_imag <= _zz_3397_;
      end
      if(_zz_3354_)begin
        int_reg_array_48_23_imag <= _zz_3397_;
      end
      if(_zz_3355_)begin
        int_reg_array_48_24_imag <= _zz_3397_;
      end
      if(_zz_3356_)begin
        int_reg_array_48_25_imag <= _zz_3397_;
      end
      if(_zz_3357_)begin
        int_reg_array_48_26_imag <= _zz_3397_;
      end
      if(_zz_3358_)begin
        int_reg_array_48_27_imag <= _zz_3397_;
      end
      if(_zz_3359_)begin
        int_reg_array_48_28_imag <= _zz_3397_;
      end
      if(_zz_3360_)begin
        int_reg_array_48_29_imag <= _zz_3397_;
      end
      if(_zz_3361_)begin
        int_reg_array_48_30_imag <= _zz_3397_;
      end
      if(_zz_3362_)begin
        int_reg_array_48_31_imag <= _zz_3397_;
      end
      if(_zz_3363_)begin
        int_reg_array_48_32_imag <= _zz_3397_;
      end
      if(_zz_3364_)begin
        int_reg_array_48_33_imag <= _zz_3397_;
      end
      if(_zz_3365_)begin
        int_reg_array_48_34_imag <= _zz_3397_;
      end
      if(_zz_3366_)begin
        int_reg_array_48_35_imag <= _zz_3397_;
      end
      if(_zz_3367_)begin
        int_reg_array_48_36_imag <= _zz_3397_;
      end
      if(_zz_3368_)begin
        int_reg_array_48_37_imag <= _zz_3397_;
      end
      if(_zz_3369_)begin
        int_reg_array_48_38_imag <= _zz_3397_;
      end
      if(_zz_3370_)begin
        int_reg_array_48_39_imag <= _zz_3397_;
      end
      if(_zz_3371_)begin
        int_reg_array_48_40_imag <= _zz_3397_;
      end
      if(_zz_3372_)begin
        int_reg_array_48_41_imag <= _zz_3397_;
      end
      if(_zz_3373_)begin
        int_reg_array_48_42_imag <= _zz_3397_;
      end
      if(_zz_3374_)begin
        int_reg_array_48_43_imag <= _zz_3397_;
      end
      if(_zz_3375_)begin
        int_reg_array_48_44_imag <= _zz_3397_;
      end
      if(_zz_3376_)begin
        int_reg_array_48_45_imag <= _zz_3397_;
      end
      if(_zz_3377_)begin
        int_reg_array_48_46_imag <= _zz_3397_;
      end
      if(_zz_3378_)begin
        int_reg_array_48_47_imag <= _zz_3397_;
      end
      if(_zz_3379_)begin
        int_reg_array_48_48_imag <= _zz_3397_;
      end
      if(_zz_3380_)begin
        int_reg_array_48_49_imag <= _zz_3397_;
      end
      if(_zz_3381_)begin
        int_reg_array_48_50_imag <= _zz_3397_;
      end
      if(_zz_3382_)begin
        int_reg_array_48_51_imag <= _zz_3397_;
      end
      if(_zz_3383_)begin
        int_reg_array_48_52_imag <= _zz_3397_;
      end
      if(_zz_3384_)begin
        int_reg_array_48_53_imag <= _zz_3397_;
      end
      if(_zz_3385_)begin
        int_reg_array_48_54_imag <= _zz_3397_;
      end
      if(_zz_3386_)begin
        int_reg_array_48_55_imag <= _zz_3397_;
      end
      if(_zz_3387_)begin
        int_reg_array_48_56_imag <= _zz_3397_;
      end
      if(_zz_3388_)begin
        int_reg_array_48_57_imag <= _zz_3397_;
      end
      if(_zz_3389_)begin
        int_reg_array_48_58_imag <= _zz_3397_;
      end
      if(_zz_3390_)begin
        int_reg_array_48_59_imag <= _zz_3397_;
      end
      if(_zz_3391_)begin
        int_reg_array_48_60_imag <= _zz_3397_;
      end
      if(_zz_3392_)begin
        int_reg_array_48_61_imag <= _zz_3397_;
      end
      if(_zz_3393_)begin
        int_reg_array_48_62_imag <= _zz_3397_;
      end
      if(_zz_3394_)begin
        int_reg_array_48_63_imag <= _zz_3397_;
      end
      if(_zz_3400_)begin
        int_reg_array_49_0_real <= _zz_3465_;
      end
      if(_zz_3401_)begin
        int_reg_array_49_1_real <= _zz_3465_;
      end
      if(_zz_3402_)begin
        int_reg_array_49_2_real <= _zz_3465_;
      end
      if(_zz_3403_)begin
        int_reg_array_49_3_real <= _zz_3465_;
      end
      if(_zz_3404_)begin
        int_reg_array_49_4_real <= _zz_3465_;
      end
      if(_zz_3405_)begin
        int_reg_array_49_5_real <= _zz_3465_;
      end
      if(_zz_3406_)begin
        int_reg_array_49_6_real <= _zz_3465_;
      end
      if(_zz_3407_)begin
        int_reg_array_49_7_real <= _zz_3465_;
      end
      if(_zz_3408_)begin
        int_reg_array_49_8_real <= _zz_3465_;
      end
      if(_zz_3409_)begin
        int_reg_array_49_9_real <= _zz_3465_;
      end
      if(_zz_3410_)begin
        int_reg_array_49_10_real <= _zz_3465_;
      end
      if(_zz_3411_)begin
        int_reg_array_49_11_real <= _zz_3465_;
      end
      if(_zz_3412_)begin
        int_reg_array_49_12_real <= _zz_3465_;
      end
      if(_zz_3413_)begin
        int_reg_array_49_13_real <= _zz_3465_;
      end
      if(_zz_3414_)begin
        int_reg_array_49_14_real <= _zz_3465_;
      end
      if(_zz_3415_)begin
        int_reg_array_49_15_real <= _zz_3465_;
      end
      if(_zz_3416_)begin
        int_reg_array_49_16_real <= _zz_3465_;
      end
      if(_zz_3417_)begin
        int_reg_array_49_17_real <= _zz_3465_;
      end
      if(_zz_3418_)begin
        int_reg_array_49_18_real <= _zz_3465_;
      end
      if(_zz_3419_)begin
        int_reg_array_49_19_real <= _zz_3465_;
      end
      if(_zz_3420_)begin
        int_reg_array_49_20_real <= _zz_3465_;
      end
      if(_zz_3421_)begin
        int_reg_array_49_21_real <= _zz_3465_;
      end
      if(_zz_3422_)begin
        int_reg_array_49_22_real <= _zz_3465_;
      end
      if(_zz_3423_)begin
        int_reg_array_49_23_real <= _zz_3465_;
      end
      if(_zz_3424_)begin
        int_reg_array_49_24_real <= _zz_3465_;
      end
      if(_zz_3425_)begin
        int_reg_array_49_25_real <= _zz_3465_;
      end
      if(_zz_3426_)begin
        int_reg_array_49_26_real <= _zz_3465_;
      end
      if(_zz_3427_)begin
        int_reg_array_49_27_real <= _zz_3465_;
      end
      if(_zz_3428_)begin
        int_reg_array_49_28_real <= _zz_3465_;
      end
      if(_zz_3429_)begin
        int_reg_array_49_29_real <= _zz_3465_;
      end
      if(_zz_3430_)begin
        int_reg_array_49_30_real <= _zz_3465_;
      end
      if(_zz_3431_)begin
        int_reg_array_49_31_real <= _zz_3465_;
      end
      if(_zz_3432_)begin
        int_reg_array_49_32_real <= _zz_3465_;
      end
      if(_zz_3433_)begin
        int_reg_array_49_33_real <= _zz_3465_;
      end
      if(_zz_3434_)begin
        int_reg_array_49_34_real <= _zz_3465_;
      end
      if(_zz_3435_)begin
        int_reg_array_49_35_real <= _zz_3465_;
      end
      if(_zz_3436_)begin
        int_reg_array_49_36_real <= _zz_3465_;
      end
      if(_zz_3437_)begin
        int_reg_array_49_37_real <= _zz_3465_;
      end
      if(_zz_3438_)begin
        int_reg_array_49_38_real <= _zz_3465_;
      end
      if(_zz_3439_)begin
        int_reg_array_49_39_real <= _zz_3465_;
      end
      if(_zz_3440_)begin
        int_reg_array_49_40_real <= _zz_3465_;
      end
      if(_zz_3441_)begin
        int_reg_array_49_41_real <= _zz_3465_;
      end
      if(_zz_3442_)begin
        int_reg_array_49_42_real <= _zz_3465_;
      end
      if(_zz_3443_)begin
        int_reg_array_49_43_real <= _zz_3465_;
      end
      if(_zz_3444_)begin
        int_reg_array_49_44_real <= _zz_3465_;
      end
      if(_zz_3445_)begin
        int_reg_array_49_45_real <= _zz_3465_;
      end
      if(_zz_3446_)begin
        int_reg_array_49_46_real <= _zz_3465_;
      end
      if(_zz_3447_)begin
        int_reg_array_49_47_real <= _zz_3465_;
      end
      if(_zz_3448_)begin
        int_reg_array_49_48_real <= _zz_3465_;
      end
      if(_zz_3449_)begin
        int_reg_array_49_49_real <= _zz_3465_;
      end
      if(_zz_3450_)begin
        int_reg_array_49_50_real <= _zz_3465_;
      end
      if(_zz_3451_)begin
        int_reg_array_49_51_real <= _zz_3465_;
      end
      if(_zz_3452_)begin
        int_reg_array_49_52_real <= _zz_3465_;
      end
      if(_zz_3453_)begin
        int_reg_array_49_53_real <= _zz_3465_;
      end
      if(_zz_3454_)begin
        int_reg_array_49_54_real <= _zz_3465_;
      end
      if(_zz_3455_)begin
        int_reg_array_49_55_real <= _zz_3465_;
      end
      if(_zz_3456_)begin
        int_reg_array_49_56_real <= _zz_3465_;
      end
      if(_zz_3457_)begin
        int_reg_array_49_57_real <= _zz_3465_;
      end
      if(_zz_3458_)begin
        int_reg_array_49_58_real <= _zz_3465_;
      end
      if(_zz_3459_)begin
        int_reg_array_49_59_real <= _zz_3465_;
      end
      if(_zz_3460_)begin
        int_reg_array_49_60_real <= _zz_3465_;
      end
      if(_zz_3461_)begin
        int_reg_array_49_61_real <= _zz_3465_;
      end
      if(_zz_3462_)begin
        int_reg_array_49_62_real <= _zz_3465_;
      end
      if(_zz_3463_)begin
        int_reg_array_49_63_real <= _zz_3465_;
      end
      if(_zz_3400_)begin
        int_reg_array_49_0_imag <= _zz_3466_;
      end
      if(_zz_3401_)begin
        int_reg_array_49_1_imag <= _zz_3466_;
      end
      if(_zz_3402_)begin
        int_reg_array_49_2_imag <= _zz_3466_;
      end
      if(_zz_3403_)begin
        int_reg_array_49_3_imag <= _zz_3466_;
      end
      if(_zz_3404_)begin
        int_reg_array_49_4_imag <= _zz_3466_;
      end
      if(_zz_3405_)begin
        int_reg_array_49_5_imag <= _zz_3466_;
      end
      if(_zz_3406_)begin
        int_reg_array_49_6_imag <= _zz_3466_;
      end
      if(_zz_3407_)begin
        int_reg_array_49_7_imag <= _zz_3466_;
      end
      if(_zz_3408_)begin
        int_reg_array_49_8_imag <= _zz_3466_;
      end
      if(_zz_3409_)begin
        int_reg_array_49_9_imag <= _zz_3466_;
      end
      if(_zz_3410_)begin
        int_reg_array_49_10_imag <= _zz_3466_;
      end
      if(_zz_3411_)begin
        int_reg_array_49_11_imag <= _zz_3466_;
      end
      if(_zz_3412_)begin
        int_reg_array_49_12_imag <= _zz_3466_;
      end
      if(_zz_3413_)begin
        int_reg_array_49_13_imag <= _zz_3466_;
      end
      if(_zz_3414_)begin
        int_reg_array_49_14_imag <= _zz_3466_;
      end
      if(_zz_3415_)begin
        int_reg_array_49_15_imag <= _zz_3466_;
      end
      if(_zz_3416_)begin
        int_reg_array_49_16_imag <= _zz_3466_;
      end
      if(_zz_3417_)begin
        int_reg_array_49_17_imag <= _zz_3466_;
      end
      if(_zz_3418_)begin
        int_reg_array_49_18_imag <= _zz_3466_;
      end
      if(_zz_3419_)begin
        int_reg_array_49_19_imag <= _zz_3466_;
      end
      if(_zz_3420_)begin
        int_reg_array_49_20_imag <= _zz_3466_;
      end
      if(_zz_3421_)begin
        int_reg_array_49_21_imag <= _zz_3466_;
      end
      if(_zz_3422_)begin
        int_reg_array_49_22_imag <= _zz_3466_;
      end
      if(_zz_3423_)begin
        int_reg_array_49_23_imag <= _zz_3466_;
      end
      if(_zz_3424_)begin
        int_reg_array_49_24_imag <= _zz_3466_;
      end
      if(_zz_3425_)begin
        int_reg_array_49_25_imag <= _zz_3466_;
      end
      if(_zz_3426_)begin
        int_reg_array_49_26_imag <= _zz_3466_;
      end
      if(_zz_3427_)begin
        int_reg_array_49_27_imag <= _zz_3466_;
      end
      if(_zz_3428_)begin
        int_reg_array_49_28_imag <= _zz_3466_;
      end
      if(_zz_3429_)begin
        int_reg_array_49_29_imag <= _zz_3466_;
      end
      if(_zz_3430_)begin
        int_reg_array_49_30_imag <= _zz_3466_;
      end
      if(_zz_3431_)begin
        int_reg_array_49_31_imag <= _zz_3466_;
      end
      if(_zz_3432_)begin
        int_reg_array_49_32_imag <= _zz_3466_;
      end
      if(_zz_3433_)begin
        int_reg_array_49_33_imag <= _zz_3466_;
      end
      if(_zz_3434_)begin
        int_reg_array_49_34_imag <= _zz_3466_;
      end
      if(_zz_3435_)begin
        int_reg_array_49_35_imag <= _zz_3466_;
      end
      if(_zz_3436_)begin
        int_reg_array_49_36_imag <= _zz_3466_;
      end
      if(_zz_3437_)begin
        int_reg_array_49_37_imag <= _zz_3466_;
      end
      if(_zz_3438_)begin
        int_reg_array_49_38_imag <= _zz_3466_;
      end
      if(_zz_3439_)begin
        int_reg_array_49_39_imag <= _zz_3466_;
      end
      if(_zz_3440_)begin
        int_reg_array_49_40_imag <= _zz_3466_;
      end
      if(_zz_3441_)begin
        int_reg_array_49_41_imag <= _zz_3466_;
      end
      if(_zz_3442_)begin
        int_reg_array_49_42_imag <= _zz_3466_;
      end
      if(_zz_3443_)begin
        int_reg_array_49_43_imag <= _zz_3466_;
      end
      if(_zz_3444_)begin
        int_reg_array_49_44_imag <= _zz_3466_;
      end
      if(_zz_3445_)begin
        int_reg_array_49_45_imag <= _zz_3466_;
      end
      if(_zz_3446_)begin
        int_reg_array_49_46_imag <= _zz_3466_;
      end
      if(_zz_3447_)begin
        int_reg_array_49_47_imag <= _zz_3466_;
      end
      if(_zz_3448_)begin
        int_reg_array_49_48_imag <= _zz_3466_;
      end
      if(_zz_3449_)begin
        int_reg_array_49_49_imag <= _zz_3466_;
      end
      if(_zz_3450_)begin
        int_reg_array_49_50_imag <= _zz_3466_;
      end
      if(_zz_3451_)begin
        int_reg_array_49_51_imag <= _zz_3466_;
      end
      if(_zz_3452_)begin
        int_reg_array_49_52_imag <= _zz_3466_;
      end
      if(_zz_3453_)begin
        int_reg_array_49_53_imag <= _zz_3466_;
      end
      if(_zz_3454_)begin
        int_reg_array_49_54_imag <= _zz_3466_;
      end
      if(_zz_3455_)begin
        int_reg_array_49_55_imag <= _zz_3466_;
      end
      if(_zz_3456_)begin
        int_reg_array_49_56_imag <= _zz_3466_;
      end
      if(_zz_3457_)begin
        int_reg_array_49_57_imag <= _zz_3466_;
      end
      if(_zz_3458_)begin
        int_reg_array_49_58_imag <= _zz_3466_;
      end
      if(_zz_3459_)begin
        int_reg_array_49_59_imag <= _zz_3466_;
      end
      if(_zz_3460_)begin
        int_reg_array_49_60_imag <= _zz_3466_;
      end
      if(_zz_3461_)begin
        int_reg_array_49_61_imag <= _zz_3466_;
      end
      if(_zz_3462_)begin
        int_reg_array_49_62_imag <= _zz_3466_;
      end
      if(_zz_3463_)begin
        int_reg_array_49_63_imag <= _zz_3466_;
      end
      if(_zz_3469_)begin
        int_reg_array_50_0_real <= _zz_3534_;
      end
      if(_zz_3470_)begin
        int_reg_array_50_1_real <= _zz_3534_;
      end
      if(_zz_3471_)begin
        int_reg_array_50_2_real <= _zz_3534_;
      end
      if(_zz_3472_)begin
        int_reg_array_50_3_real <= _zz_3534_;
      end
      if(_zz_3473_)begin
        int_reg_array_50_4_real <= _zz_3534_;
      end
      if(_zz_3474_)begin
        int_reg_array_50_5_real <= _zz_3534_;
      end
      if(_zz_3475_)begin
        int_reg_array_50_6_real <= _zz_3534_;
      end
      if(_zz_3476_)begin
        int_reg_array_50_7_real <= _zz_3534_;
      end
      if(_zz_3477_)begin
        int_reg_array_50_8_real <= _zz_3534_;
      end
      if(_zz_3478_)begin
        int_reg_array_50_9_real <= _zz_3534_;
      end
      if(_zz_3479_)begin
        int_reg_array_50_10_real <= _zz_3534_;
      end
      if(_zz_3480_)begin
        int_reg_array_50_11_real <= _zz_3534_;
      end
      if(_zz_3481_)begin
        int_reg_array_50_12_real <= _zz_3534_;
      end
      if(_zz_3482_)begin
        int_reg_array_50_13_real <= _zz_3534_;
      end
      if(_zz_3483_)begin
        int_reg_array_50_14_real <= _zz_3534_;
      end
      if(_zz_3484_)begin
        int_reg_array_50_15_real <= _zz_3534_;
      end
      if(_zz_3485_)begin
        int_reg_array_50_16_real <= _zz_3534_;
      end
      if(_zz_3486_)begin
        int_reg_array_50_17_real <= _zz_3534_;
      end
      if(_zz_3487_)begin
        int_reg_array_50_18_real <= _zz_3534_;
      end
      if(_zz_3488_)begin
        int_reg_array_50_19_real <= _zz_3534_;
      end
      if(_zz_3489_)begin
        int_reg_array_50_20_real <= _zz_3534_;
      end
      if(_zz_3490_)begin
        int_reg_array_50_21_real <= _zz_3534_;
      end
      if(_zz_3491_)begin
        int_reg_array_50_22_real <= _zz_3534_;
      end
      if(_zz_3492_)begin
        int_reg_array_50_23_real <= _zz_3534_;
      end
      if(_zz_3493_)begin
        int_reg_array_50_24_real <= _zz_3534_;
      end
      if(_zz_3494_)begin
        int_reg_array_50_25_real <= _zz_3534_;
      end
      if(_zz_3495_)begin
        int_reg_array_50_26_real <= _zz_3534_;
      end
      if(_zz_3496_)begin
        int_reg_array_50_27_real <= _zz_3534_;
      end
      if(_zz_3497_)begin
        int_reg_array_50_28_real <= _zz_3534_;
      end
      if(_zz_3498_)begin
        int_reg_array_50_29_real <= _zz_3534_;
      end
      if(_zz_3499_)begin
        int_reg_array_50_30_real <= _zz_3534_;
      end
      if(_zz_3500_)begin
        int_reg_array_50_31_real <= _zz_3534_;
      end
      if(_zz_3501_)begin
        int_reg_array_50_32_real <= _zz_3534_;
      end
      if(_zz_3502_)begin
        int_reg_array_50_33_real <= _zz_3534_;
      end
      if(_zz_3503_)begin
        int_reg_array_50_34_real <= _zz_3534_;
      end
      if(_zz_3504_)begin
        int_reg_array_50_35_real <= _zz_3534_;
      end
      if(_zz_3505_)begin
        int_reg_array_50_36_real <= _zz_3534_;
      end
      if(_zz_3506_)begin
        int_reg_array_50_37_real <= _zz_3534_;
      end
      if(_zz_3507_)begin
        int_reg_array_50_38_real <= _zz_3534_;
      end
      if(_zz_3508_)begin
        int_reg_array_50_39_real <= _zz_3534_;
      end
      if(_zz_3509_)begin
        int_reg_array_50_40_real <= _zz_3534_;
      end
      if(_zz_3510_)begin
        int_reg_array_50_41_real <= _zz_3534_;
      end
      if(_zz_3511_)begin
        int_reg_array_50_42_real <= _zz_3534_;
      end
      if(_zz_3512_)begin
        int_reg_array_50_43_real <= _zz_3534_;
      end
      if(_zz_3513_)begin
        int_reg_array_50_44_real <= _zz_3534_;
      end
      if(_zz_3514_)begin
        int_reg_array_50_45_real <= _zz_3534_;
      end
      if(_zz_3515_)begin
        int_reg_array_50_46_real <= _zz_3534_;
      end
      if(_zz_3516_)begin
        int_reg_array_50_47_real <= _zz_3534_;
      end
      if(_zz_3517_)begin
        int_reg_array_50_48_real <= _zz_3534_;
      end
      if(_zz_3518_)begin
        int_reg_array_50_49_real <= _zz_3534_;
      end
      if(_zz_3519_)begin
        int_reg_array_50_50_real <= _zz_3534_;
      end
      if(_zz_3520_)begin
        int_reg_array_50_51_real <= _zz_3534_;
      end
      if(_zz_3521_)begin
        int_reg_array_50_52_real <= _zz_3534_;
      end
      if(_zz_3522_)begin
        int_reg_array_50_53_real <= _zz_3534_;
      end
      if(_zz_3523_)begin
        int_reg_array_50_54_real <= _zz_3534_;
      end
      if(_zz_3524_)begin
        int_reg_array_50_55_real <= _zz_3534_;
      end
      if(_zz_3525_)begin
        int_reg_array_50_56_real <= _zz_3534_;
      end
      if(_zz_3526_)begin
        int_reg_array_50_57_real <= _zz_3534_;
      end
      if(_zz_3527_)begin
        int_reg_array_50_58_real <= _zz_3534_;
      end
      if(_zz_3528_)begin
        int_reg_array_50_59_real <= _zz_3534_;
      end
      if(_zz_3529_)begin
        int_reg_array_50_60_real <= _zz_3534_;
      end
      if(_zz_3530_)begin
        int_reg_array_50_61_real <= _zz_3534_;
      end
      if(_zz_3531_)begin
        int_reg_array_50_62_real <= _zz_3534_;
      end
      if(_zz_3532_)begin
        int_reg_array_50_63_real <= _zz_3534_;
      end
      if(_zz_3469_)begin
        int_reg_array_50_0_imag <= _zz_3535_;
      end
      if(_zz_3470_)begin
        int_reg_array_50_1_imag <= _zz_3535_;
      end
      if(_zz_3471_)begin
        int_reg_array_50_2_imag <= _zz_3535_;
      end
      if(_zz_3472_)begin
        int_reg_array_50_3_imag <= _zz_3535_;
      end
      if(_zz_3473_)begin
        int_reg_array_50_4_imag <= _zz_3535_;
      end
      if(_zz_3474_)begin
        int_reg_array_50_5_imag <= _zz_3535_;
      end
      if(_zz_3475_)begin
        int_reg_array_50_6_imag <= _zz_3535_;
      end
      if(_zz_3476_)begin
        int_reg_array_50_7_imag <= _zz_3535_;
      end
      if(_zz_3477_)begin
        int_reg_array_50_8_imag <= _zz_3535_;
      end
      if(_zz_3478_)begin
        int_reg_array_50_9_imag <= _zz_3535_;
      end
      if(_zz_3479_)begin
        int_reg_array_50_10_imag <= _zz_3535_;
      end
      if(_zz_3480_)begin
        int_reg_array_50_11_imag <= _zz_3535_;
      end
      if(_zz_3481_)begin
        int_reg_array_50_12_imag <= _zz_3535_;
      end
      if(_zz_3482_)begin
        int_reg_array_50_13_imag <= _zz_3535_;
      end
      if(_zz_3483_)begin
        int_reg_array_50_14_imag <= _zz_3535_;
      end
      if(_zz_3484_)begin
        int_reg_array_50_15_imag <= _zz_3535_;
      end
      if(_zz_3485_)begin
        int_reg_array_50_16_imag <= _zz_3535_;
      end
      if(_zz_3486_)begin
        int_reg_array_50_17_imag <= _zz_3535_;
      end
      if(_zz_3487_)begin
        int_reg_array_50_18_imag <= _zz_3535_;
      end
      if(_zz_3488_)begin
        int_reg_array_50_19_imag <= _zz_3535_;
      end
      if(_zz_3489_)begin
        int_reg_array_50_20_imag <= _zz_3535_;
      end
      if(_zz_3490_)begin
        int_reg_array_50_21_imag <= _zz_3535_;
      end
      if(_zz_3491_)begin
        int_reg_array_50_22_imag <= _zz_3535_;
      end
      if(_zz_3492_)begin
        int_reg_array_50_23_imag <= _zz_3535_;
      end
      if(_zz_3493_)begin
        int_reg_array_50_24_imag <= _zz_3535_;
      end
      if(_zz_3494_)begin
        int_reg_array_50_25_imag <= _zz_3535_;
      end
      if(_zz_3495_)begin
        int_reg_array_50_26_imag <= _zz_3535_;
      end
      if(_zz_3496_)begin
        int_reg_array_50_27_imag <= _zz_3535_;
      end
      if(_zz_3497_)begin
        int_reg_array_50_28_imag <= _zz_3535_;
      end
      if(_zz_3498_)begin
        int_reg_array_50_29_imag <= _zz_3535_;
      end
      if(_zz_3499_)begin
        int_reg_array_50_30_imag <= _zz_3535_;
      end
      if(_zz_3500_)begin
        int_reg_array_50_31_imag <= _zz_3535_;
      end
      if(_zz_3501_)begin
        int_reg_array_50_32_imag <= _zz_3535_;
      end
      if(_zz_3502_)begin
        int_reg_array_50_33_imag <= _zz_3535_;
      end
      if(_zz_3503_)begin
        int_reg_array_50_34_imag <= _zz_3535_;
      end
      if(_zz_3504_)begin
        int_reg_array_50_35_imag <= _zz_3535_;
      end
      if(_zz_3505_)begin
        int_reg_array_50_36_imag <= _zz_3535_;
      end
      if(_zz_3506_)begin
        int_reg_array_50_37_imag <= _zz_3535_;
      end
      if(_zz_3507_)begin
        int_reg_array_50_38_imag <= _zz_3535_;
      end
      if(_zz_3508_)begin
        int_reg_array_50_39_imag <= _zz_3535_;
      end
      if(_zz_3509_)begin
        int_reg_array_50_40_imag <= _zz_3535_;
      end
      if(_zz_3510_)begin
        int_reg_array_50_41_imag <= _zz_3535_;
      end
      if(_zz_3511_)begin
        int_reg_array_50_42_imag <= _zz_3535_;
      end
      if(_zz_3512_)begin
        int_reg_array_50_43_imag <= _zz_3535_;
      end
      if(_zz_3513_)begin
        int_reg_array_50_44_imag <= _zz_3535_;
      end
      if(_zz_3514_)begin
        int_reg_array_50_45_imag <= _zz_3535_;
      end
      if(_zz_3515_)begin
        int_reg_array_50_46_imag <= _zz_3535_;
      end
      if(_zz_3516_)begin
        int_reg_array_50_47_imag <= _zz_3535_;
      end
      if(_zz_3517_)begin
        int_reg_array_50_48_imag <= _zz_3535_;
      end
      if(_zz_3518_)begin
        int_reg_array_50_49_imag <= _zz_3535_;
      end
      if(_zz_3519_)begin
        int_reg_array_50_50_imag <= _zz_3535_;
      end
      if(_zz_3520_)begin
        int_reg_array_50_51_imag <= _zz_3535_;
      end
      if(_zz_3521_)begin
        int_reg_array_50_52_imag <= _zz_3535_;
      end
      if(_zz_3522_)begin
        int_reg_array_50_53_imag <= _zz_3535_;
      end
      if(_zz_3523_)begin
        int_reg_array_50_54_imag <= _zz_3535_;
      end
      if(_zz_3524_)begin
        int_reg_array_50_55_imag <= _zz_3535_;
      end
      if(_zz_3525_)begin
        int_reg_array_50_56_imag <= _zz_3535_;
      end
      if(_zz_3526_)begin
        int_reg_array_50_57_imag <= _zz_3535_;
      end
      if(_zz_3527_)begin
        int_reg_array_50_58_imag <= _zz_3535_;
      end
      if(_zz_3528_)begin
        int_reg_array_50_59_imag <= _zz_3535_;
      end
      if(_zz_3529_)begin
        int_reg_array_50_60_imag <= _zz_3535_;
      end
      if(_zz_3530_)begin
        int_reg_array_50_61_imag <= _zz_3535_;
      end
      if(_zz_3531_)begin
        int_reg_array_50_62_imag <= _zz_3535_;
      end
      if(_zz_3532_)begin
        int_reg_array_50_63_imag <= _zz_3535_;
      end
      if(_zz_3538_)begin
        int_reg_array_51_0_real <= _zz_3603_;
      end
      if(_zz_3539_)begin
        int_reg_array_51_1_real <= _zz_3603_;
      end
      if(_zz_3540_)begin
        int_reg_array_51_2_real <= _zz_3603_;
      end
      if(_zz_3541_)begin
        int_reg_array_51_3_real <= _zz_3603_;
      end
      if(_zz_3542_)begin
        int_reg_array_51_4_real <= _zz_3603_;
      end
      if(_zz_3543_)begin
        int_reg_array_51_5_real <= _zz_3603_;
      end
      if(_zz_3544_)begin
        int_reg_array_51_6_real <= _zz_3603_;
      end
      if(_zz_3545_)begin
        int_reg_array_51_7_real <= _zz_3603_;
      end
      if(_zz_3546_)begin
        int_reg_array_51_8_real <= _zz_3603_;
      end
      if(_zz_3547_)begin
        int_reg_array_51_9_real <= _zz_3603_;
      end
      if(_zz_3548_)begin
        int_reg_array_51_10_real <= _zz_3603_;
      end
      if(_zz_3549_)begin
        int_reg_array_51_11_real <= _zz_3603_;
      end
      if(_zz_3550_)begin
        int_reg_array_51_12_real <= _zz_3603_;
      end
      if(_zz_3551_)begin
        int_reg_array_51_13_real <= _zz_3603_;
      end
      if(_zz_3552_)begin
        int_reg_array_51_14_real <= _zz_3603_;
      end
      if(_zz_3553_)begin
        int_reg_array_51_15_real <= _zz_3603_;
      end
      if(_zz_3554_)begin
        int_reg_array_51_16_real <= _zz_3603_;
      end
      if(_zz_3555_)begin
        int_reg_array_51_17_real <= _zz_3603_;
      end
      if(_zz_3556_)begin
        int_reg_array_51_18_real <= _zz_3603_;
      end
      if(_zz_3557_)begin
        int_reg_array_51_19_real <= _zz_3603_;
      end
      if(_zz_3558_)begin
        int_reg_array_51_20_real <= _zz_3603_;
      end
      if(_zz_3559_)begin
        int_reg_array_51_21_real <= _zz_3603_;
      end
      if(_zz_3560_)begin
        int_reg_array_51_22_real <= _zz_3603_;
      end
      if(_zz_3561_)begin
        int_reg_array_51_23_real <= _zz_3603_;
      end
      if(_zz_3562_)begin
        int_reg_array_51_24_real <= _zz_3603_;
      end
      if(_zz_3563_)begin
        int_reg_array_51_25_real <= _zz_3603_;
      end
      if(_zz_3564_)begin
        int_reg_array_51_26_real <= _zz_3603_;
      end
      if(_zz_3565_)begin
        int_reg_array_51_27_real <= _zz_3603_;
      end
      if(_zz_3566_)begin
        int_reg_array_51_28_real <= _zz_3603_;
      end
      if(_zz_3567_)begin
        int_reg_array_51_29_real <= _zz_3603_;
      end
      if(_zz_3568_)begin
        int_reg_array_51_30_real <= _zz_3603_;
      end
      if(_zz_3569_)begin
        int_reg_array_51_31_real <= _zz_3603_;
      end
      if(_zz_3570_)begin
        int_reg_array_51_32_real <= _zz_3603_;
      end
      if(_zz_3571_)begin
        int_reg_array_51_33_real <= _zz_3603_;
      end
      if(_zz_3572_)begin
        int_reg_array_51_34_real <= _zz_3603_;
      end
      if(_zz_3573_)begin
        int_reg_array_51_35_real <= _zz_3603_;
      end
      if(_zz_3574_)begin
        int_reg_array_51_36_real <= _zz_3603_;
      end
      if(_zz_3575_)begin
        int_reg_array_51_37_real <= _zz_3603_;
      end
      if(_zz_3576_)begin
        int_reg_array_51_38_real <= _zz_3603_;
      end
      if(_zz_3577_)begin
        int_reg_array_51_39_real <= _zz_3603_;
      end
      if(_zz_3578_)begin
        int_reg_array_51_40_real <= _zz_3603_;
      end
      if(_zz_3579_)begin
        int_reg_array_51_41_real <= _zz_3603_;
      end
      if(_zz_3580_)begin
        int_reg_array_51_42_real <= _zz_3603_;
      end
      if(_zz_3581_)begin
        int_reg_array_51_43_real <= _zz_3603_;
      end
      if(_zz_3582_)begin
        int_reg_array_51_44_real <= _zz_3603_;
      end
      if(_zz_3583_)begin
        int_reg_array_51_45_real <= _zz_3603_;
      end
      if(_zz_3584_)begin
        int_reg_array_51_46_real <= _zz_3603_;
      end
      if(_zz_3585_)begin
        int_reg_array_51_47_real <= _zz_3603_;
      end
      if(_zz_3586_)begin
        int_reg_array_51_48_real <= _zz_3603_;
      end
      if(_zz_3587_)begin
        int_reg_array_51_49_real <= _zz_3603_;
      end
      if(_zz_3588_)begin
        int_reg_array_51_50_real <= _zz_3603_;
      end
      if(_zz_3589_)begin
        int_reg_array_51_51_real <= _zz_3603_;
      end
      if(_zz_3590_)begin
        int_reg_array_51_52_real <= _zz_3603_;
      end
      if(_zz_3591_)begin
        int_reg_array_51_53_real <= _zz_3603_;
      end
      if(_zz_3592_)begin
        int_reg_array_51_54_real <= _zz_3603_;
      end
      if(_zz_3593_)begin
        int_reg_array_51_55_real <= _zz_3603_;
      end
      if(_zz_3594_)begin
        int_reg_array_51_56_real <= _zz_3603_;
      end
      if(_zz_3595_)begin
        int_reg_array_51_57_real <= _zz_3603_;
      end
      if(_zz_3596_)begin
        int_reg_array_51_58_real <= _zz_3603_;
      end
      if(_zz_3597_)begin
        int_reg_array_51_59_real <= _zz_3603_;
      end
      if(_zz_3598_)begin
        int_reg_array_51_60_real <= _zz_3603_;
      end
      if(_zz_3599_)begin
        int_reg_array_51_61_real <= _zz_3603_;
      end
      if(_zz_3600_)begin
        int_reg_array_51_62_real <= _zz_3603_;
      end
      if(_zz_3601_)begin
        int_reg_array_51_63_real <= _zz_3603_;
      end
      if(_zz_3538_)begin
        int_reg_array_51_0_imag <= _zz_3604_;
      end
      if(_zz_3539_)begin
        int_reg_array_51_1_imag <= _zz_3604_;
      end
      if(_zz_3540_)begin
        int_reg_array_51_2_imag <= _zz_3604_;
      end
      if(_zz_3541_)begin
        int_reg_array_51_3_imag <= _zz_3604_;
      end
      if(_zz_3542_)begin
        int_reg_array_51_4_imag <= _zz_3604_;
      end
      if(_zz_3543_)begin
        int_reg_array_51_5_imag <= _zz_3604_;
      end
      if(_zz_3544_)begin
        int_reg_array_51_6_imag <= _zz_3604_;
      end
      if(_zz_3545_)begin
        int_reg_array_51_7_imag <= _zz_3604_;
      end
      if(_zz_3546_)begin
        int_reg_array_51_8_imag <= _zz_3604_;
      end
      if(_zz_3547_)begin
        int_reg_array_51_9_imag <= _zz_3604_;
      end
      if(_zz_3548_)begin
        int_reg_array_51_10_imag <= _zz_3604_;
      end
      if(_zz_3549_)begin
        int_reg_array_51_11_imag <= _zz_3604_;
      end
      if(_zz_3550_)begin
        int_reg_array_51_12_imag <= _zz_3604_;
      end
      if(_zz_3551_)begin
        int_reg_array_51_13_imag <= _zz_3604_;
      end
      if(_zz_3552_)begin
        int_reg_array_51_14_imag <= _zz_3604_;
      end
      if(_zz_3553_)begin
        int_reg_array_51_15_imag <= _zz_3604_;
      end
      if(_zz_3554_)begin
        int_reg_array_51_16_imag <= _zz_3604_;
      end
      if(_zz_3555_)begin
        int_reg_array_51_17_imag <= _zz_3604_;
      end
      if(_zz_3556_)begin
        int_reg_array_51_18_imag <= _zz_3604_;
      end
      if(_zz_3557_)begin
        int_reg_array_51_19_imag <= _zz_3604_;
      end
      if(_zz_3558_)begin
        int_reg_array_51_20_imag <= _zz_3604_;
      end
      if(_zz_3559_)begin
        int_reg_array_51_21_imag <= _zz_3604_;
      end
      if(_zz_3560_)begin
        int_reg_array_51_22_imag <= _zz_3604_;
      end
      if(_zz_3561_)begin
        int_reg_array_51_23_imag <= _zz_3604_;
      end
      if(_zz_3562_)begin
        int_reg_array_51_24_imag <= _zz_3604_;
      end
      if(_zz_3563_)begin
        int_reg_array_51_25_imag <= _zz_3604_;
      end
      if(_zz_3564_)begin
        int_reg_array_51_26_imag <= _zz_3604_;
      end
      if(_zz_3565_)begin
        int_reg_array_51_27_imag <= _zz_3604_;
      end
      if(_zz_3566_)begin
        int_reg_array_51_28_imag <= _zz_3604_;
      end
      if(_zz_3567_)begin
        int_reg_array_51_29_imag <= _zz_3604_;
      end
      if(_zz_3568_)begin
        int_reg_array_51_30_imag <= _zz_3604_;
      end
      if(_zz_3569_)begin
        int_reg_array_51_31_imag <= _zz_3604_;
      end
      if(_zz_3570_)begin
        int_reg_array_51_32_imag <= _zz_3604_;
      end
      if(_zz_3571_)begin
        int_reg_array_51_33_imag <= _zz_3604_;
      end
      if(_zz_3572_)begin
        int_reg_array_51_34_imag <= _zz_3604_;
      end
      if(_zz_3573_)begin
        int_reg_array_51_35_imag <= _zz_3604_;
      end
      if(_zz_3574_)begin
        int_reg_array_51_36_imag <= _zz_3604_;
      end
      if(_zz_3575_)begin
        int_reg_array_51_37_imag <= _zz_3604_;
      end
      if(_zz_3576_)begin
        int_reg_array_51_38_imag <= _zz_3604_;
      end
      if(_zz_3577_)begin
        int_reg_array_51_39_imag <= _zz_3604_;
      end
      if(_zz_3578_)begin
        int_reg_array_51_40_imag <= _zz_3604_;
      end
      if(_zz_3579_)begin
        int_reg_array_51_41_imag <= _zz_3604_;
      end
      if(_zz_3580_)begin
        int_reg_array_51_42_imag <= _zz_3604_;
      end
      if(_zz_3581_)begin
        int_reg_array_51_43_imag <= _zz_3604_;
      end
      if(_zz_3582_)begin
        int_reg_array_51_44_imag <= _zz_3604_;
      end
      if(_zz_3583_)begin
        int_reg_array_51_45_imag <= _zz_3604_;
      end
      if(_zz_3584_)begin
        int_reg_array_51_46_imag <= _zz_3604_;
      end
      if(_zz_3585_)begin
        int_reg_array_51_47_imag <= _zz_3604_;
      end
      if(_zz_3586_)begin
        int_reg_array_51_48_imag <= _zz_3604_;
      end
      if(_zz_3587_)begin
        int_reg_array_51_49_imag <= _zz_3604_;
      end
      if(_zz_3588_)begin
        int_reg_array_51_50_imag <= _zz_3604_;
      end
      if(_zz_3589_)begin
        int_reg_array_51_51_imag <= _zz_3604_;
      end
      if(_zz_3590_)begin
        int_reg_array_51_52_imag <= _zz_3604_;
      end
      if(_zz_3591_)begin
        int_reg_array_51_53_imag <= _zz_3604_;
      end
      if(_zz_3592_)begin
        int_reg_array_51_54_imag <= _zz_3604_;
      end
      if(_zz_3593_)begin
        int_reg_array_51_55_imag <= _zz_3604_;
      end
      if(_zz_3594_)begin
        int_reg_array_51_56_imag <= _zz_3604_;
      end
      if(_zz_3595_)begin
        int_reg_array_51_57_imag <= _zz_3604_;
      end
      if(_zz_3596_)begin
        int_reg_array_51_58_imag <= _zz_3604_;
      end
      if(_zz_3597_)begin
        int_reg_array_51_59_imag <= _zz_3604_;
      end
      if(_zz_3598_)begin
        int_reg_array_51_60_imag <= _zz_3604_;
      end
      if(_zz_3599_)begin
        int_reg_array_51_61_imag <= _zz_3604_;
      end
      if(_zz_3600_)begin
        int_reg_array_51_62_imag <= _zz_3604_;
      end
      if(_zz_3601_)begin
        int_reg_array_51_63_imag <= _zz_3604_;
      end
      if(_zz_3607_)begin
        int_reg_array_52_0_real <= _zz_3672_;
      end
      if(_zz_3608_)begin
        int_reg_array_52_1_real <= _zz_3672_;
      end
      if(_zz_3609_)begin
        int_reg_array_52_2_real <= _zz_3672_;
      end
      if(_zz_3610_)begin
        int_reg_array_52_3_real <= _zz_3672_;
      end
      if(_zz_3611_)begin
        int_reg_array_52_4_real <= _zz_3672_;
      end
      if(_zz_3612_)begin
        int_reg_array_52_5_real <= _zz_3672_;
      end
      if(_zz_3613_)begin
        int_reg_array_52_6_real <= _zz_3672_;
      end
      if(_zz_3614_)begin
        int_reg_array_52_7_real <= _zz_3672_;
      end
      if(_zz_3615_)begin
        int_reg_array_52_8_real <= _zz_3672_;
      end
      if(_zz_3616_)begin
        int_reg_array_52_9_real <= _zz_3672_;
      end
      if(_zz_3617_)begin
        int_reg_array_52_10_real <= _zz_3672_;
      end
      if(_zz_3618_)begin
        int_reg_array_52_11_real <= _zz_3672_;
      end
      if(_zz_3619_)begin
        int_reg_array_52_12_real <= _zz_3672_;
      end
      if(_zz_3620_)begin
        int_reg_array_52_13_real <= _zz_3672_;
      end
      if(_zz_3621_)begin
        int_reg_array_52_14_real <= _zz_3672_;
      end
      if(_zz_3622_)begin
        int_reg_array_52_15_real <= _zz_3672_;
      end
      if(_zz_3623_)begin
        int_reg_array_52_16_real <= _zz_3672_;
      end
      if(_zz_3624_)begin
        int_reg_array_52_17_real <= _zz_3672_;
      end
      if(_zz_3625_)begin
        int_reg_array_52_18_real <= _zz_3672_;
      end
      if(_zz_3626_)begin
        int_reg_array_52_19_real <= _zz_3672_;
      end
      if(_zz_3627_)begin
        int_reg_array_52_20_real <= _zz_3672_;
      end
      if(_zz_3628_)begin
        int_reg_array_52_21_real <= _zz_3672_;
      end
      if(_zz_3629_)begin
        int_reg_array_52_22_real <= _zz_3672_;
      end
      if(_zz_3630_)begin
        int_reg_array_52_23_real <= _zz_3672_;
      end
      if(_zz_3631_)begin
        int_reg_array_52_24_real <= _zz_3672_;
      end
      if(_zz_3632_)begin
        int_reg_array_52_25_real <= _zz_3672_;
      end
      if(_zz_3633_)begin
        int_reg_array_52_26_real <= _zz_3672_;
      end
      if(_zz_3634_)begin
        int_reg_array_52_27_real <= _zz_3672_;
      end
      if(_zz_3635_)begin
        int_reg_array_52_28_real <= _zz_3672_;
      end
      if(_zz_3636_)begin
        int_reg_array_52_29_real <= _zz_3672_;
      end
      if(_zz_3637_)begin
        int_reg_array_52_30_real <= _zz_3672_;
      end
      if(_zz_3638_)begin
        int_reg_array_52_31_real <= _zz_3672_;
      end
      if(_zz_3639_)begin
        int_reg_array_52_32_real <= _zz_3672_;
      end
      if(_zz_3640_)begin
        int_reg_array_52_33_real <= _zz_3672_;
      end
      if(_zz_3641_)begin
        int_reg_array_52_34_real <= _zz_3672_;
      end
      if(_zz_3642_)begin
        int_reg_array_52_35_real <= _zz_3672_;
      end
      if(_zz_3643_)begin
        int_reg_array_52_36_real <= _zz_3672_;
      end
      if(_zz_3644_)begin
        int_reg_array_52_37_real <= _zz_3672_;
      end
      if(_zz_3645_)begin
        int_reg_array_52_38_real <= _zz_3672_;
      end
      if(_zz_3646_)begin
        int_reg_array_52_39_real <= _zz_3672_;
      end
      if(_zz_3647_)begin
        int_reg_array_52_40_real <= _zz_3672_;
      end
      if(_zz_3648_)begin
        int_reg_array_52_41_real <= _zz_3672_;
      end
      if(_zz_3649_)begin
        int_reg_array_52_42_real <= _zz_3672_;
      end
      if(_zz_3650_)begin
        int_reg_array_52_43_real <= _zz_3672_;
      end
      if(_zz_3651_)begin
        int_reg_array_52_44_real <= _zz_3672_;
      end
      if(_zz_3652_)begin
        int_reg_array_52_45_real <= _zz_3672_;
      end
      if(_zz_3653_)begin
        int_reg_array_52_46_real <= _zz_3672_;
      end
      if(_zz_3654_)begin
        int_reg_array_52_47_real <= _zz_3672_;
      end
      if(_zz_3655_)begin
        int_reg_array_52_48_real <= _zz_3672_;
      end
      if(_zz_3656_)begin
        int_reg_array_52_49_real <= _zz_3672_;
      end
      if(_zz_3657_)begin
        int_reg_array_52_50_real <= _zz_3672_;
      end
      if(_zz_3658_)begin
        int_reg_array_52_51_real <= _zz_3672_;
      end
      if(_zz_3659_)begin
        int_reg_array_52_52_real <= _zz_3672_;
      end
      if(_zz_3660_)begin
        int_reg_array_52_53_real <= _zz_3672_;
      end
      if(_zz_3661_)begin
        int_reg_array_52_54_real <= _zz_3672_;
      end
      if(_zz_3662_)begin
        int_reg_array_52_55_real <= _zz_3672_;
      end
      if(_zz_3663_)begin
        int_reg_array_52_56_real <= _zz_3672_;
      end
      if(_zz_3664_)begin
        int_reg_array_52_57_real <= _zz_3672_;
      end
      if(_zz_3665_)begin
        int_reg_array_52_58_real <= _zz_3672_;
      end
      if(_zz_3666_)begin
        int_reg_array_52_59_real <= _zz_3672_;
      end
      if(_zz_3667_)begin
        int_reg_array_52_60_real <= _zz_3672_;
      end
      if(_zz_3668_)begin
        int_reg_array_52_61_real <= _zz_3672_;
      end
      if(_zz_3669_)begin
        int_reg_array_52_62_real <= _zz_3672_;
      end
      if(_zz_3670_)begin
        int_reg_array_52_63_real <= _zz_3672_;
      end
      if(_zz_3607_)begin
        int_reg_array_52_0_imag <= _zz_3673_;
      end
      if(_zz_3608_)begin
        int_reg_array_52_1_imag <= _zz_3673_;
      end
      if(_zz_3609_)begin
        int_reg_array_52_2_imag <= _zz_3673_;
      end
      if(_zz_3610_)begin
        int_reg_array_52_3_imag <= _zz_3673_;
      end
      if(_zz_3611_)begin
        int_reg_array_52_4_imag <= _zz_3673_;
      end
      if(_zz_3612_)begin
        int_reg_array_52_5_imag <= _zz_3673_;
      end
      if(_zz_3613_)begin
        int_reg_array_52_6_imag <= _zz_3673_;
      end
      if(_zz_3614_)begin
        int_reg_array_52_7_imag <= _zz_3673_;
      end
      if(_zz_3615_)begin
        int_reg_array_52_8_imag <= _zz_3673_;
      end
      if(_zz_3616_)begin
        int_reg_array_52_9_imag <= _zz_3673_;
      end
      if(_zz_3617_)begin
        int_reg_array_52_10_imag <= _zz_3673_;
      end
      if(_zz_3618_)begin
        int_reg_array_52_11_imag <= _zz_3673_;
      end
      if(_zz_3619_)begin
        int_reg_array_52_12_imag <= _zz_3673_;
      end
      if(_zz_3620_)begin
        int_reg_array_52_13_imag <= _zz_3673_;
      end
      if(_zz_3621_)begin
        int_reg_array_52_14_imag <= _zz_3673_;
      end
      if(_zz_3622_)begin
        int_reg_array_52_15_imag <= _zz_3673_;
      end
      if(_zz_3623_)begin
        int_reg_array_52_16_imag <= _zz_3673_;
      end
      if(_zz_3624_)begin
        int_reg_array_52_17_imag <= _zz_3673_;
      end
      if(_zz_3625_)begin
        int_reg_array_52_18_imag <= _zz_3673_;
      end
      if(_zz_3626_)begin
        int_reg_array_52_19_imag <= _zz_3673_;
      end
      if(_zz_3627_)begin
        int_reg_array_52_20_imag <= _zz_3673_;
      end
      if(_zz_3628_)begin
        int_reg_array_52_21_imag <= _zz_3673_;
      end
      if(_zz_3629_)begin
        int_reg_array_52_22_imag <= _zz_3673_;
      end
      if(_zz_3630_)begin
        int_reg_array_52_23_imag <= _zz_3673_;
      end
      if(_zz_3631_)begin
        int_reg_array_52_24_imag <= _zz_3673_;
      end
      if(_zz_3632_)begin
        int_reg_array_52_25_imag <= _zz_3673_;
      end
      if(_zz_3633_)begin
        int_reg_array_52_26_imag <= _zz_3673_;
      end
      if(_zz_3634_)begin
        int_reg_array_52_27_imag <= _zz_3673_;
      end
      if(_zz_3635_)begin
        int_reg_array_52_28_imag <= _zz_3673_;
      end
      if(_zz_3636_)begin
        int_reg_array_52_29_imag <= _zz_3673_;
      end
      if(_zz_3637_)begin
        int_reg_array_52_30_imag <= _zz_3673_;
      end
      if(_zz_3638_)begin
        int_reg_array_52_31_imag <= _zz_3673_;
      end
      if(_zz_3639_)begin
        int_reg_array_52_32_imag <= _zz_3673_;
      end
      if(_zz_3640_)begin
        int_reg_array_52_33_imag <= _zz_3673_;
      end
      if(_zz_3641_)begin
        int_reg_array_52_34_imag <= _zz_3673_;
      end
      if(_zz_3642_)begin
        int_reg_array_52_35_imag <= _zz_3673_;
      end
      if(_zz_3643_)begin
        int_reg_array_52_36_imag <= _zz_3673_;
      end
      if(_zz_3644_)begin
        int_reg_array_52_37_imag <= _zz_3673_;
      end
      if(_zz_3645_)begin
        int_reg_array_52_38_imag <= _zz_3673_;
      end
      if(_zz_3646_)begin
        int_reg_array_52_39_imag <= _zz_3673_;
      end
      if(_zz_3647_)begin
        int_reg_array_52_40_imag <= _zz_3673_;
      end
      if(_zz_3648_)begin
        int_reg_array_52_41_imag <= _zz_3673_;
      end
      if(_zz_3649_)begin
        int_reg_array_52_42_imag <= _zz_3673_;
      end
      if(_zz_3650_)begin
        int_reg_array_52_43_imag <= _zz_3673_;
      end
      if(_zz_3651_)begin
        int_reg_array_52_44_imag <= _zz_3673_;
      end
      if(_zz_3652_)begin
        int_reg_array_52_45_imag <= _zz_3673_;
      end
      if(_zz_3653_)begin
        int_reg_array_52_46_imag <= _zz_3673_;
      end
      if(_zz_3654_)begin
        int_reg_array_52_47_imag <= _zz_3673_;
      end
      if(_zz_3655_)begin
        int_reg_array_52_48_imag <= _zz_3673_;
      end
      if(_zz_3656_)begin
        int_reg_array_52_49_imag <= _zz_3673_;
      end
      if(_zz_3657_)begin
        int_reg_array_52_50_imag <= _zz_3673_;
      end
      if(_zz_3658_)begin
        int_reg_array_52_51_imag <= _zz_3673_;
      end
      if(_zz_3659_)begin
        int_reg_array_52_52_imag <= _zz_3673_;
      end
      if(_zz_3660_)begin
        int_reg_array_52_53_imag <= _zz_3673_;
      end
      if(_zz_3661_)begin
        int_reg_array_52_54_imag <= _zz_3673_;
      end
      if(_zz_3662_)begin
        int_reg_array_52_55_imag <= _zz_3673_;
      end
      if(_zz_3663_)begin
        int_reg_array_52_56_imag <= _zz_3673_;
      end
      if(_zz_3664_)begin
        int_reg_array_52_57_imag <= _zz_3673_;
      end
      if(_zz_3665_)begin
        int_reg_array_52_58_imag <= _zz_3673_;
      end
      if(_zz_3666_)begin
        int_reg_array_52_59_imag <= _zz_3673_;
      end
      if(_zz_3667_)begin
        int_reg_array_52_60_imag <= _zz_3673_;
      end
      if(_zz_3668_)begin
        int_reg_array_52_61_imag <= _zz_3673_;
      end
      if(_zz_3669_)begin
        int_reg_array_52_62_imag <= _zz_3673_;
      end
      if(_zz_3670_)begin
        int_reg_array_52_63_imag <= _zz_3673_;
      end
      if(_zz_3676_)begin
        int_reg_array_53_0_real <= _zz_3741_;
      end
      if(_zz_3677_)begin
        int_reg_array_53_1_real <= _zz_3741_;
      end
      if(_zz_3678_)begin
        int_reg_array_53_2_real <= _zz_3741_;
      end
      if(_zz_3679_)begin
        int_reg_array_53_3_real <= _zz_3741_;
      end
      if(_zz_3680_)begin
        int_reg_array_53_4_real <= _zz_3741_;
      end
      if(_zz_3681_)begin
        int_reg_array_53_5_real <= _zz_3741_;
      end
      if(_zz_3682_)begin
        int_reg_array_53_6_real <= _zz_3741_;
      end
      if(_zz_3683_)begin
        int_reg_array_53_7_real <= _zz_3741_;
      end
      if(_zz_3684_)begin
        int_reg_array_53_8_real <= _zz_3741_;
      end
      if(_zz_3685_)begin
        int_reg_array_53_9_real <= _zz_3741_;
      end
      if(_zz_3686_)begin
        int_reg_array_53_10_real <= _zz_3741_;
      end
      if(_zz_3687_)begin
        int_reg_array_53_11_real <= _zz_3741_;
      end
      if(_zz_3688_)begin
        int_reg_array_53_12_real <= _zz_3741_;
      end
      if(_zz_3689_)begin
        int_reg_array_53_13_real <= _zz_3741_;
      end
      if(_zz_3690_)begin
        int_reg_array_53_14_real <= _zz_3741_;
      end
      if(_zz_3691_)begin
        int_reg_array_53_15_real <= _zz_3741_;
      end
      if(_zz_3692_)begin
        int_reg_array_53_16_real <= _zz_3741_;
      end
      if(_zz_3693_)begin
        int_reg_array_53_17_real <= _zz_3741_;
      end
      if(_zz_3694_)begin
        int_reg_array_53_18_real <= _zz_3741_;
      end
      if(_zz_3695_)begin
        int_reg_array_53_19_real <= _zz_3741_;
      end
      if(_zz_3696_)begin
        int_reg_array_53_20_real <= _zz_3741_;
      end
      if(_zz_3697_)begin
        int_reg_array_53_21_real <= _zz_3741_;
      end
      if(_zz_3698_)begin
        int_reg_array_53_22_real <= _zz_3741_;
      end
      if(_zz_3699_)begin
        int_reg_array_53_23_real <= _zz_3741_;
      end
      if(_zz_3700_)begin
        int_reg_array_53_24_real <= _zz_3741_;
      end
      if(_zz_3701_)begin
        int_reg_array_53_25_real <= _zz_3741_;
      end
      if(_zz_3702_)begin
        int_reg_array_53_26_real <= _zz_3741_;
      end
      if(_zz_3703_)begin
        int_reg_array_53_27_real <= _zz_3741_;
      end
      if(_zz_3704_)begin
        int_reg_array_53_28_real <= _zz_3741_;
      end
      if(_zz_3705_)begin
        int_reg_array_53_29_real <= _zz_3741_;
      end
      if(_zz_3706_)begin
        int_reg_array_53_30_real <= _zz_3741_;
      end
      if(_zz_3707_)begin
        int_reg_array_53_31_real <= _zz_3741_;
      end
      if(_zz_3708_)begin
        int_reg_array_53_32_real <= _zz_3741_;
      end
      if(_zz_3709_)begin
        int_reg_array_53_33_real <= _zz_3741_;
      end
      if(_zz_3710_)begin
        int_reg_array_53_34_real <= _zz_3741_;
      end
      if(_zz_3711_)begin
        int_reg_array_53_35_real <= _zz_3741_;
      end
      if(_zz_3712_)begin
        int_reg_array_53_36_real <= _zz_3741_;
      end
      if(_zz_3713_)begin
        int_reg_array_53_37_real <= _zz_3741_;
      end
      if(_zz_3714_)begin
        int_reg_array_53_38_real <= _zz_3741_;
      end
      if(_zz_3715_)begin
        int_reg_array_53_39_real <= _zz_3741_;
      end
      if(_zz_3716_)begin
        int_reg_array_53_40_real <= _zz_3741_;
      end
      if(_zz_3717_)begin
        int_reg_array_53_41_real <= _zz_3741_;
      end
      if(_zz_3718_)begin
        int_reg_array_53_42_real <= _zz_3741_;
      end
      if(_zz_3719_)begin
        int_reg_array_53_43_real <= _zz_3741_;
      end
      if(_zz_3720_)begin
        int_reg_array_53_44_real <= _zz_3741_;
      end
      if(_zz_3721_)begin
        int_reg_array_53_45_real <= _zz_3741_;
      end
      if(_zz_3722_)begin
        int_reg_array_53_46_real <= _zz_3741_;
      end
      if(_zz_3723_)begin
        int_reg_array_53_47_real <= _zz_3741_;
      end
      if(_zz_3724_)begin
        int_reg_array_53_48_real <= _zz_3741_;
      end
      if(_zz_3725_)begin
        int_reg_array_53_49_real <= _zz_3741_;
      end
      if(_zz_3726_)begin
        int_reg_array_53_50_real <= _zz_3741_;
      end
      if(_zz_3727_)begin
        int_reg_array_53_51_real <= _zz_3741_;
      end
      if(_zz_3728_)begin
        int_reg_array_53_52_real <= _zz_3741_;
      end
      if(_zz_3729_)begin
        int_reg_array_53_53_real <= _zz_3741_;
      end
      if(_zz_3730_)begin
        int_reg_array_53_54_real <= _zz_3741_;
      end
      if(_zz_3731_)begin
        int_reg_array_53_55_real <= _zz_3741_;
      end
      if(_zz_3732_)begin
        int_reg_array_53_56_real <= _zz_3741_;
      end
      if(_zz_3733_)begin
        int_reg_array_53_57_real <= _zz_3741_;
      end
      if(_zz_3734_)begin
        int_reg_array_53_58_real <= _zz_3741_;
      end
      if(_zz_3735_)begin
        int_reg_array_53_59_real <= _zz_3741_;
      end
      if(_zz_3736_)begin
        int_reg_array_53_60_real <= _zz_3741_;
      end
      if(_zz_3737_)begin
        int_reg_array_53_61_real <= _zz_3741_;
      end
      if(_zz_3738_)begin
        int_reg_array_53_62_real <= _zz_3741_;
      end
      if(_zz_3739_)begin
        int_reg_array_53_63_real <= _zz_3741_;
      end
      if(_zz_3676_)begin
        int_reg_array_53_0_imag <= _zz_3742_;
      end
      if(_zz_3677_)begin
        int_reg_array_53_1_imag <= _zz_3742_;
      end
      if(_zz_3678_)begin
        int_reg_array_53_2_imag <= _zz_3742_;
      end
      if(_zz_3679_)begin
        int_reg_array_53_3_imag <= _zz_3742_;
      end
      if(_zz_3680_)begin
        int_reg_array_53_4_imag <= _zz_3742_;
      end
      if(_zz_3681_)begin
        int_reg_array_53_5_imag <= _zz_3742_;
      end
      if(_zz_3682_)begin
        int_reg_array_53_6_imag <= _zz_3742_;
      end
      if(_zz_3683_)begin
        int_reg_array_53_7_imag <= _zz_3742_;
      end
      if(_zz_3684_)begin
        int_reg_array_53_8_imag <= _zz_3742_;
      end
      if(_zz_3685_)begin
        int_reg_array_53_9_imag <= _zz_3742_;
      end
      if(_zz_3686_)begin
        int_reg_array_53_10_imag <= _zz_3742_;
      end
      if(_zz_3687_)begin
        int_reg_array_53_11_imag <= _zz_3742_;
      end
      if(_zz_3688_)begin
        int_reg_array_53_12_imag <= _zz_3742_;
      end
      if(_zz_3689_)begin
        int_reg_array_53_13_imag <= _zz_3742_;
      end
      if(_zz_3690_)begin
        int_reg_array_53_14_imag <= _zz_3742_;
      end
      if(_zz_3691_)begin
        int_reg_array_53_15_imag <= _zz_3742_;
      end
      if(_zz_3692_)begin
        int_reg_array_53_16_imag <= _zz_3742_;
      end
      if(_zz_3693_)begin
        int_reg_array_53_17_imag <= _zz_3742_;
      end
      if(_zz_3694_)begin
        int_reg_array_53_18_imag <= _zz_3742_;
      end
      if(_zz_3695_)begin
        int_reg_array_53_19_imag <= _zz_3742_;
      end
      if(_zz_3696_)begin
        int_reg_array_53_20_imag <= _zz_3742_;
      end
      if(_zz_3697_)begin
        int_reg_array_53_21_imag <= _zz_3742_;
      end
      if(_zz_3698_)begin
        int_reg_array_53_22_imag <= _zz_3742_;
      end
      if(_zz_3699_)begin
        int_reg_array_53_23_imag <= _zz_3742_;
      end
      if(_zz_3700_)begin
        int_reg_array_53_24_imag <= _zz_3742_;
      end
      if(_zz_3701_)begin
        int_reg_array_53_25_imag <= _zz_3742_;
      end
      if(_zz_3702_)begin
        int_reg_array_53_26_imag <= _zz_3742_;
      end
      if(_zz_3703_)begin
        int_reg_array_53_27_imag <= _zz_3742_;
      end
      if(_zz_3704_)begin
        int_reg_array_53_28_imag <= _zz_3742_;
      end
      if(_zz_3705_)begin
        int_reg_array_53_29_imag <= _zz_3742_;
      end
      if(_zz_3706_)begin
        int_reg_array_53_30_imag <= _zz_3742_;
      end
      if(_zz_3707_)begin
        int_reg_array_53_31_imag <= _zz_3742_;
      end
      if(_zz_3708_)begin
        int_reg_array_53_32_imag <= _zz_3742_;
      end
      if(_zz_3709_)begin
        int_reg_array_53_33_imag <= _zz_3742_;
      end
      if(_zz_3710_)begin
        int_reg_array_53_34_imag <= _zz_3742_;
      end
      if(_zz_3711_)begin
        int_reg_array_53_35_imag <= _zz_3742_;
      end
      if(_zz_3712_)begin
        int_reg_array_53_36_imag <= _zz_3742_;
      end
      if(_zz_3713_)begin
        int_reg_array_53_37_imag <= _zz_3742_;
      end
      if(_zz_3714_)begin
        int_reg_array_53_38_imag <= _zz_3742_;
      end
      if(_zz_3715_)begin
        int_reg_array_53_39_imag <= _zz_3742_;
      end
      if(_zz_3716_)begin
        int_reg_array_53_40_imag <= _zz_3742_;
      end
      if(_zz_3717_)begin
        int_reg_array_53_41_imag <= _zz_3742_;
      end
      if(_zz_3718_)begin
        int_reg_array_53_42_imag <= _zz_3742_;
      end
      if(_zz_3719_)begin
        int_reg_array_53_43_imag <= _zz_3742_;
      end
      if(_zz_3720_)begin
        int_reg_array_53_44_imag <= _zz_3742_;
      end
      if(_zz_3721_)begin
        int_reg_array_53_45_imag <= _zz_3742_;
      end
      if(_zz_3722_)begin
        int_reg_array_53_46_imag <= _zz_3742_;
      end
      if(_zz_3723_)begin
        int_reg_array_53_47_imag <= _zz_3742_;
      end
      if(_zz_3724_)begin
        int_reg_array_53_48_imag <= _zz_3742_;
      end
      if(_zz_3725_)begin
        int_reg_array_53_49_imag <= _zz_3742_;
      end
      if(_zz_3726_)begin
        int_reg_array_53_50_imag <= _zz_3742_;
      end
      if(_zz_3727_)begin
        int_reg_array_53_51_imag <= _zz_3742_;
      end
      if(_zz_3728_)begin
        int_reg_array_53_52_imag <= _zz_3742_;
      end
      if(_zz_3729_)begin
        int_reg_array_53_53_imag <= _zz_3742_;
      end
      if(_zz_3730_)begin
        int_reg_array_53_54_imag <= _zz_3742_;
      end
      if(_zz_3731_)begin
        int_reg_array_53_55_imag <= _zz_3742_;
      end
      if(_zz_3732_)begin
        int_reg_array_53_56_imag <= _zz_3742_;
      end
      if(_zz_3733_)begin
        int_reg_array_53_57_imag <= _zz_3742_;
      end
      if(_zz_3734_)begin
        int_reg_array_53_58_imag <= _zz_3742_;
      end
      if(_zz_3735_)begin
        int_reg_array_53_59_imag <= _zz_3742_;
      end
      if(_zz_3736_)begin
        int_reg_array_53_60_imag <= _zz_3742_;
      end
      if(_zz_3737_)begin
        int_reg_array_53_61_imag <= _zz_3742_;
      end
      if(_zz_3738_)begin
        int_reg_array_53_62_imag <= _zz_3742_;
      end
      if(_zz_3739_)begin
        int_reg_array_53_63_imag <= _zz_3742_;
      end
      if(_zz_3745_)begin
        int_reg_array_54_0_real <= _zz_3810_;
      end
      if(_zz_3746_)begin
        int_reg_array_54_1_real <= _zz_3810_;
      end
      if(_zz_3747_)begin
        int_reg_array_54_2_real <= _zz_3810_;
      end
      if(_zz_3748_)begin
        int_reg_array_54_3_real <= _zz_3810_;
      end
      if(_zz_3749_)begin
        int_reg_array_54_4_real <= _zz_3810_;
      end
      if(_zz_3750_)begin
        int_reg_array_54_5_real <= _zz_3810_;
      end
      if(_zz_3751_)begin
        int_reg_array_54_6_real <= _zz_3810_;
      end
      if(_zz_3752_)begin
        int_reg_array_54_7_real <= _zz_3810_;
      end
      if(_zz_3753_)begin
        int_reg_array_54_8_real <= _zz_3810_;
      end
      if(_zz_3754_)begin
        int_reg_array_54_9_real <= _zz_3810_;
      end
      if(_zz_3755_)begin
        int_reg_array_54_10_real <= _zz_3810_;
      end
      if(_zz_3756_)begin
        int_reg_array_54_11_real <= _zz_3810_;
      end
      if(_zz_3757_)begin
        int_reg_array_54_12_real <= _zz_3810_;
      end
      if(_zz_3758_)begin
        int_reg_array_54_13_real <= _zz_3810_;
      end
      if(_zz_3759_)begin
        int_reg_array_54_14_real <= _zz_3810_;
      end
      if(_zz_3760_)begin
        int_reg_array_54_15_real <= _zz_3810_;
      end
      if(_zz_3761_)begin
        int_reg_array_54_16_real <= _zz_3810_;
      end
      if(_zz_3762_)begin
        int_reg_array_54_17_real <= _zz_3810_;
      end
      if(_zz_3763_)begin
        int_reg_array_54_18_real <= _zz_3810_;
      end
      if(_zz_3764_)begin
        int_reg_array_54_19_real <= _zz_3810_;
      end
      if(_zz_3765_)begin
        int_reg_array_54_20_real <= _zz_3810_;
      end
      if(_zz_3766_)begin
        int_reg_array_54_21_real <= _zz_3810_;
      end
      if(_zz_3767_)begin
        int_reg_array_54_22_real <= _zz_3810_;
      end
      if(_zz_3768_)begin
        int_reg_array_54_23_real <= _zz_3810_;
      end
      if(_zz_3769_)begin
        int_reg_array_54_24_real <= _zz_3810_;
      end
      if(_zz_3770_)begin
        int_reg_array_54_25_real <= _zz_3810_;
      end
      if(_zz_3771_)begin
        int_reg_array_54_26_real <= _zz_3810_;
      end
      if(_zz_3772_)begin
        int_reg_array_54_27_real <= _zz_3810_;
      end
      if(_zz_3773_)begin
        int_reg_array_54_28_real <= _zz_3810_;
      end
      if(_zz_3774_)begin
        int_reg_array_54_29_real <= _zz_3810_;
      end
      if(_zz_3775_)begin
        int_reg_array_54_30_real <= _zz_3810_;
      end
      if(_zz_3776_)begin
        int_reg_array_54_31_real <= _zz_3810_;
      end
      if(_zz_3777_)begin
        int_reg_array_54_32_real <= _zz_3810_;
      end
      if(_zz_3778_)begin
        int_reg_array_54_33_real <= _zz_3810_;
      end
      if(_zz_3779_)begin
        int_reg_array_54_34_real <= _zz_3810_;
      end
      if(_zz_3780_)begin
        int_reg_array_54_35_real <= _zz_3810_;
      end
      if(_zz_3781_)begin
        int_reg_array_54_36_real <= _zz_3810_;
      end
      if(_zz_3782_)begin
        int_reg_array_54_37_real <= _zz_3810_;
      end
      if(_zz_3783_)begin
        int_reg_array_54_38_real <= _zz_3810_;
      end
      if(_zz_3784_)begin
        int_reg_array_54_39_real <= _zz_3810_;
      end
      if(_zz_3785_)begin
        int_reg_array_54_40_real <= _zz_3810_;
      end
      if(_zz_3786_)begin
        int_reg_array_54_41_real <= _zz_3810_;
      end
      if(_zz_3787_)begin
        int_reg_array_54_42_real <= _zz_3810_;
      end
      if(_zz_3788_)begin
        int_reg_array_54_43_real <= _zz_3810_;
      end
      if(_zz_3789_)begin
        int_reg_array_54_44_real <= _zz_3810_;
      end
      if(_zz_3790_)begin
        int_reg_array_54_45_real <= _zz_3810_;
      end
      if(_zz_3791_)begin
        int_reg_array_54_46_real <= _zz_3810_;
      end
      if(_zz_3792_)begin
        int_reg_array_54_47_real <= _zz_3810_;
      end
      if(_zz_3793_)begin
        int_reg_array_54_48_real <= _zz_3810_;
      end
      if(_zz_3794_)begin
        int_reg_array_54_49_real <= _zz_3810_;
      end
      if(_zz_3795_)begin
        int_reg_array_54_50_real <= _zz_3810_;
      end
      if(_zz_3796_)begin
        int_reg_array_54_51_real <= _zz_3810_;
      end
      if(_zz_3797_)begin
        int_reg_array_54_52_real <= _zz_3810_;
      end
      if(_zz_3798_)begin
        int_reg_array_54_53_real <= _zz_3810_;
      end
      if(_zz_3799_)begin
        int_reg_array_54_54_real <= _zz_3810_;
      end
      if(_zz_3800_)begin
        int_reg_array_54_55_real <= _zz_3810_;
      end
      if(_zz_3801_)begin
        int_reg_array_54_56_real <= _zz_3810_;
      end
      if(_zz_3802_)begin
        int_reg_array_54_57_real <= _zz_3810_;
      end
      if(_zz_3803_)begin
        int_reg_array_54_58_real <= _zz_3810_;
      end
      if(_zz_3804_)begin
        int_reg_array_54_59_real <= _zz_3810_;
      end
      if(_zz_3805_)begin
        int_reg_array_54_60_real <= _zz_3810_;
      end
      if(_zz_3806_)begin
        int_reg_array_54_61_real <= _zz_3810_;
      end
      if(_zz_3807_)begin
        int_reg_array_54_62_real <= _zz_3810_;
      end
      if(_zz_3808_)begin
        int_reg_array_54_63_real <= _zz_3810_;
      end
      if(_zz_3745_)begin
        int_reg_array_54_0_imag <= _zz_3811_;
      end
      if(_zz_3746_)begin
        int_reg_array_54_1_imag <= _zz_3811_;
      end
      if(_zz_3747_)begin
        int_reg_array_54_2_imag <= _zz_3811_;
      end
      if(_zz_3748_)begin
        int_reg_array_54_3_imag <= _zz_3811_;
      end
      if(_zz_3749_)begin
        int_reg_array_54_4_imag <= _zz_3811_;
      end
      if(_zz_3750_)begin
        int_reg_array_54_5_imag <= _zz_3811_;
      end
      if(_zz_3751_)begin
        int_reg_array_54_6_imag <= _zz_3811_;
      end
      if(_zz_3752_)begin
        int_reg_array_54_7_imag <= _zz_3811_;
      end
      if(_zz_3753_)begin
        int_reg_array_54_8_imag <= _zz_3811_;
      end
      if(_zz_3754_)begin
        int_reg_array_54_9_imag <= _zz_3811_;
      end
      if(_zz_3755_)begin
        int_reg_array_54_10_imag <= _zz_3811_;
      end
      if(_zz_3756_)begin
        int_reg_array_54_11_imag <= _zz_3811_;
      end
      if(_zz_3757_)begin
        int_reg_array_54_12_imag <= _zz_3811_;
      end
      if(_zz_3758_)begin
        int_reg_array_54_13_imag <= _zz_3811_;
      end
      if(_zz_3759_)begin
        int_reg_array_54_14_imag <= _zz_3811_;
      end
      if(_zz_3760_)begin
        int_reg_array_54_15_imag <= _zz_3811_;
      end
      if(_zz_3761_)begin
        int_reg_array_54_16_imag <= _zz_3811_;
      end
      if(_zz_3762_)begin
        int_reg_array_54_17_imag <= _zz_3811_;
      end
      if(_zz_3763_)begin
        int_reg_array_54_18_imag <= _zz_3811_;
      end
      if(_zz_3764_)begin
        int_reg_array_54_19_imag <= _zz_3811_;
      end
      if(_zz_3765_)begin
        int_reg_array_54_20_imag <= _zz_3811_;
      end
      if(_zz_3766_)begin
        int_reg_array_54_21_imag <= _zz_3811_;
      end
      if(_zz_3767_)begin
        int_reg_array_54_22_imag <= _zz_3811_;
      end
      if(_zz_3768_)begin
        int_reg_array_54_23_imag <= _zz_3811_;
      end
      if(_zz_3769_)begin
        int_reg_array_54_24_imag <= _zz_3811_;
      end
      if(_zz_3770_)begin
        int_reg_array_54_25_imag <= _zz_3811_;
      end
      if(_zz_3771_)begin
        int_reg_array_54_26_imag <= _zz_3811_;
      end
      if(_zz_3772_)begin
        int_reg_array_54_27_imag <= _zz_3811_;
      end
      if(_zz_3773_)begin
        int_reg_array_54_28_imag <= _zz_3811_;
      end
      if(_zz_3774_)begin
        int_reg_array_54_29_imag <= _zz_3811_;
      end
      if(_zz_3775_)begin
        int_reg_array_54_30_imag <= _zz_3811_;
      end
      if(_zz_3776_)begin
        int_reg_array_54_31_imag <= _zz_3811_;
      end
      if(_zz_3777_)begin
        int_reg_array_54_32_imag <= _zz_3811_;
      end
      if(_zz_3778_)begin
        int_reg_array_54_33_imag <= _zz_3811_;
      end
      if(_zz_3779_)begin
        int_reg_array_54_34_imag <= _zz_3811_;
      end
      if(_zz_3780_)begin
        int_reg_array_54_35_imag <= _zz_3811_;
      end
      if(_zz_3781_)begin
        int_reg_array_54_36_imag <= _zz_3811_;
      end
      if(_zz_3782_)begin
        int_reg_array_54_37_imag <= _zz_3811_;
      end
      if(_zz_3783_)begin
        int_reg_array_54_38_imag <= _zz_3811_;
      end
      if(_zz_3784_)begin
        int_reg_array_54_39_imag <= _zz_3811_;
      end
      if(_zz_3785_)begin
        int_reg_array_54_40_imag <= _zz_3811_;
      end
      if(_zz_3786_)begin
        int_reg_array_54_41_imag <= _zz_3811_;
      end
      if(_zz_3787_)begin
        int_reg_array_54_42_imag <= _zz_3811_;
      end
      if(_zz_3788_)begin
        int_reg_array_54_43_imag <= _zz_3811_;
      end
      if(_zz_3789_)begin
        int_reg_array_54_44_imag <= _zz_3811_;
      end
      if(_zz_3790_)begin
        int_reg_array_54_45_imag <= _zz_3811_;
      end
      if(_zz_3791_)begin
        int_reg_array_54_46_imag <= _zz_3811_;
      end
      if(_zz_3792_)begin
        int_reg_array_54_47_imag <= _zz_3811_;
      end
      if(_zz_3793_)begin
        int_reg_array_54_48_imag <= _zz_3811_;
      end
      if(_zz_3794_)begin
        int_reg_array_54_49_imag <= _zz_3811_;
      end
      if(_zz_3795_)begin
        int_reg_array_54_50_imag <= _zz_3811_;
      end
      if(_zz_3796_)begin
        int_reg_array_54_51_imag <= _zz_3811_;
      end
      if(_zz_3797_)begin
        int_reg_array_54_52_imag <= _zz_3811_;
      end
      if(_zz_3798_)begin
        int_reg_array_54_53_imag <= _zz_3811_;
      end
      if(_zz_3799_)begin
        int_reg_array_54_54_imag <= _zz_3811_;
      end
      if(_zz_3800_)begin
        int_reg_array_54_55_imag <= _zz_3811_;
      end
      if(_zz_3801_)begin
        int_reg_array_54_56_imag <= _zz_3811_;
      end
      if(_zz_3802_)begin
        int_reg_array_54_57_imag <= _zz_3811_;
      end
      if(_zz_3803_)begin
        int_reg_array_54_58_imag <= _zz_3811_;
      end
      if(_zz_3804_)begin
        int_reg_array_54_59_imag <= _zz_3811_;
      end
      if(_zz_3805_)begin
        int_reg_array_54_60_imag <= _zz_3811_;
      end
      if(_zz_3806_)begin
        int_reg_array_54_61_imag <= _zz_3811_;
      end
      if(_zz_3807_)begin
        int_reg_array_54_62_imag <= _zz_3811_;
      end
      if(_zz_3808_)begin
        int_reg_array_54_63_imag <= _zz_3811_;
      end
      if(_zz_3814_)begin
        int_reg_array_55_0_real <= _zz_3879_;
      end
      if(_zz_3815_)begin
        int_reg_array_55_1_real <= _zz_3879_;
      end
      if(_zz_3816_)begin
        int_reg_array_55_2_real <= _zz_3879_;
      end
      if(_zz_3817_)begin
        int_reg_array_55_3_real <= _zz_3879_;
      end
      if(_zz_3818_)begin
        int_reg_array_55_4_real <= _zz_3879_;
      end
      if(_zz_3819_)begin
        int_reg_array_55_5_real <= _zz_3879_;
      end
      if(_zz_3820_)begin
        int_reg_array_55_6_real <= _zz_3879_;
      end
      if(_zz_3821_)begin
        int_reg_array_55_7_real <= _zz_3879_;
      end
      if(_zz_3822_)begin
        int_reg_array_55_8_real <= _zz_3879_;
      end
      if(_zz_3823_)begin
        int_reg_array_55_9_real <= _zz_3879_;
      end
      if(_zz_3824_)begin
        int_reg_array_55_10_real <= _zz_3879_;
      end
      if(_zz_3825_)begin
        int_reg_array_55_11_real <= _zz_3879_;
      end
      if(_zz_3826_)begin
        int_reg_array_55_12_real <= _zz_3879_;
      end
      if(_zz_3827_)begin
        int_reg_array_55_13_real <= _zz_3879_;
      end
      if(_zz_3828_)begin
        int_reg_array_55_14_real <= _zz_3879_;
      end
      if(_zz_3829_)begin
        int_reg_array_55_15_real <= _zz_3879_;
      end
      if(_zz_3830_)begin
        int_reg_array_55_16_real <= _zz_3879_;
      end
      if(_zz_3831_)begin
        int_reg_array_55_17_real <= _zz_3879_;
      end
      if(_zz_3832_)begin
        int_reg_array_55_18_real <= _zz_3879_;
      end
      if(_zz_3833_)begin
        int_reg_array_55_19_real <= _zz_3879_;
      end
      if(_zz_3834_)begin
        int_reg_array_55_20_real <= _zz_3879_;
      end
      if(_zz_3835_)begin
        int_reg_array_55_21_real <= _zz_3879_;
      end
      if(_zz_3836_)begin
        int_reg_array_55_22_real <= _zz_3879_;
      end
      if(_zz_3837_)begin
        int_reg_array_55_23_real <= _zz_3879_;
      end
      if(_zz_3838_)begin
        int_reg_array_55_24_real <= _zz_3879_;
      end
      if(_zz_3839_)begin
        int_reg_array_55_25_real <= _zz_3879_;
      end
      if(_zz_3840_)begin
        int_reg_array_55_26_real <= _zz_3879_;
      end
      if(_zz_3841_)begin
        int_reg_array_55_27_real <= _zz_3879_;
      end
      if(_zz_3842_)begin
        int_reg_array_55_28_real <= _zz_3879_;
      end
      if(_zz_3843_)begin
        int_reg_array_55_29_real <= _zz_3879_;
      end
      if(_zz_3844_)begin
        int_reg_array_55_30_real <= _zz_3879_;
      end
      if(_zz_3845_)begin
        int_reg_array_55_31_real <= _zz_3879_;
      end
      if(_zz_3846_)begin
        int_reg_array_55_32_real <= _zz_3879_;
      end
      if(_zz_3847_)begin
        int_reg_array_55_33_real <= _zz_3879_;
      end
      if(_zz_3848_)begin
        int_reg_array_55_34_real <= _zz_3879_;
      end
      if(_zz_3849_)begin
        int_reg_array_55_35_real <= _zz_3879_;
      end
      if(_zz_3850_)begin
        int_reg_array_55_36_real <= _zz_3879_;
      end
      if(_zz_3851_)begin
        int_reg_array_55_37_real <= _zz_3879_;
      end
      if(_zz_3852_)begin
        int_reg_array_55_38_real <= _zz_3879_;
      end
      if(_zz_3853_)begin
        int_reg_array_55_39_real <= _zz_3879_;
      end
      if(_zz_3854_)begin
        int_reg_array_55_40_real <= _zz_3879_;
      end
      if(_zz_3855_)begin
        int_reg_array_55_41_real <= _zz_3879_;
      end
      if(_zz_3856_)begin
        int_reg_array_55_42_real <= _zz_3879_;
      end
      if(_zz_3857_)begin
        int_reg_array_55_43_real <= _zz_3879_;
      end
      if(_zz_3858_)begin
        int_reg_array_55_44_real <= _zz_3879_;
      end
      if(_zz_3859_)begin
        int_reg_array_55_45_real <= _zz_3879_;
      end
      if(_zz_3860_)begin
        int_reg_array_55_46_real <= _zz_3879_;
      end
      if(_zz_3861_)begin
        int_reg_array_55_47_real <= _zz_3879_;
      end
      if(_zz_3862_)begin
        int_reg_array_55_48_real <= _zz_3879_;
      end
      if(_zz_3863_)begin
        int_reg_array_55_49_real <= _zz_3879_;
      end
      if(_zz_3864_)begin
        int_reg_array_55_50_real <= _zz_3879_;
      end
      if(_zz_3865_)begin
        int_reg_array_55_51_real <= _zz_3879_;
      end
      if(_zz_3866_)begin
        int_reg_array_55_52_real <= _zz_3879_;
      end
      if(_zz_3867_)begin
        int_reg_array_55_53_real <= _zz_3879_;
      end
      if(_zz_3868_)begin
        int_reg_array_55_54_real <= _zz_3879_;
      end
      if(_zz_3869_)begin
        int_reg_array_55_55_real <= _zz_3879_;
      end
      if(_zz_3870_)begin
        int_reg_array_55_56_real <= _zz_3879_;
      end
      if(_zz_3871_)begin
        int_reg_array_55_57_real <= _zz_3879_;
      end
      if(_zz_3872_)begin
        int_reg_array_55_58_real <= _zz_3879_;
      end
      if(_zz_3873_)begin
        int_reg_array_55_59_real <= _zz_3879_;
      end
      if(_zz_3874_)begin
        int_reg_array_55_60_real <= _zz_3879_;
      end
      if(_zz_3875_)begin
        int_reg_array_55_61_real <= _zz_3879_;
      end
      if(_zz_3876_)begin
        int_reg_array_55_62_real <= _zz_3879_;
      end
      if(_zz_3877_)begin
        int_reg_array_55_63_real <= _zz_3879_;
      end
      if(_zz_3814_)begin
        int_reg_array_55_0_imag <= _zz_3880_;
      end
      if(_zz_3815_)begin
        int_reg_array_55_1_imag <= _zz_3880_;
      end
      if(_zz_3816_)begin
        int_reg_array_55_2_imag <= _zz_3880_;
      end
      if(_zz_3817_)begin
        int_reg_array_55_3_imag <= _zz_3880_;
      end
      if(_zz_3818_)begin
        int_reg_array_55_4_imag <= _zz_3880_;
      end
      if(_zz_3819_)begin
        int_reg_array_55_5_imag <= _zz_3880_;
      end
      if(_zz_3820_)begin
        int_reg_array_55_6_imag <= _zz_3880_;
      end
      if(_zz_3821_)begin
        int_reg_array_55_7_imag <= _zz_3880_;
      end
      if(_zz_3822_)begin
        int_reg_array_55_8_imag <= _zz_3880_;
      end
      if(_zz_3823_)begin
        int_reg_array_55_9_imag <= _zz_3880_;
      end
      if(_zz_3824_)begin
        int_reg_array_55_10_imag <= _zz_3880_;
      end
      if(_zz_3825_)begin
        int_reg_array_55_11_imag <= _zz_3880_;
      end
      if(_zz_3826_)begin
        int_reg_array_55_12_imag <= _zz_3880_;
      end
      if(_zz_3827_)begin
        int_reg_array_55_13_imag <= _zz_3880_;
      end
      if(_zz_3828_)begin
        int_reg_array_55_14_imag <= _zz_3880_;
      end
      if(_zz_3829_)begin
        int_reg_array_55_15_imag <= _zz_3880_;
      end
      if(_zz_3830_)begin
        int_reg_array_55_16_imag <= _zz_3880_;
      end
      if(_zz_3831_)begin
        int_reg_array_55_17_imag <= _zz_3880_;
      end
      if(_zz_3832_)begin
        int_reg_array_55_18_imag <= _zz_3880_;
      end
      if(_zz_3833_)begin
        int_reg_array_55_19_imag <= _zz_3880_;
      end
      if(_zz_3834_)begin
        int_reg_array_55_20_imag <= _zz_3880_;
      end
      if(_zz_3835_)begin
        int_reg_array_55_21_imag <= _zz_3880_;
      end
      if(_zz_3836_)begin
        int_reg_array_55_22_imag <= _zz_3880_;
      end
      if(_zz_3837_)begin
        int_reg_array_55_23_imag <= _zz_3880_;
      end
      if(_zz_3838_)begin
        int_reg_array_55_24_imag <= _zz_3880_;
      end
      if(_zz_3839_)begin
        int_reg_array_55_25_imag <= _zz_3880_;
      end
      if(_zz_3840_)begin
        int_reg_array_55_26_imag <= _zz_3880_;
      end
      if(_zz_3841_)begin
        int_reg_array_55_27_imag <= _zz_3880_;
      end
      if(_zz_3842_)begin
        int_reg_array_55_28_imag <= _zz_3880_;
      end
      if(_zz_3843_)begin
        int_reg_array_55_29_imag <= _zz_3880_;
      end
      if(_zz_3844_)begin
        int_reg_array_55_30_imag <= _zz_3880_;
      end
      if(_zz_3845_)begin
        int_reg_array_55_31_imag <= _zz_3880_;
      end
      if(_zz_3846_)begin
        int_reg_array_55_32_imag <= _zz_3880_;
      end
      if(_zz_3847_)begin
        int_reg_array_55_33_imag <= _zz_3880_;
      end
      if(_zz_3848_)begin
        int_reg_array_55_34_imag <= _zz_3880_;
      end
      if(_zz_3849_)begin
        int_reg_array_55_35_imag <= _zz_3880_;
      end
      if(_zz_3850_)begin
        int_reg_array_55_36_imag <= _zz_3880_;
      end
      if(_zz_3851_)begin
        int_reg_array_55_37_imag <= _zz_3880_;
      end
      if(_zz_3852_)begin
        int_reg_array_55_38_imag <= _zz_3880_;
      end
      if(_zz_3853_)begin
        int_reg_array_55_39_imag <= _zz_3880_;
      end
      if(_zz_3854_)begin
        int_reg_array_55_40_imag <= _zz_3880_;
      end
      if(_zz_3855_)begin
        int_reg_array_55_41_imag <= _zz_3880_;
      end
      if(_zz_3856_)begin
        int_reg_array_55_42_imag <= _zz_3880_;
      end
      if(_zz_3857_)begin
        int_reg_array_55_43_imag <= _zz_3880_;
      end
      if(_zz_3858_)begin
        int_reg_array_55_44_imag <= _zz_3880_;
      end
      if(_zz_3859_)begin
        int_reg_array_55_45_imag <= _zz_3880_;
      end
      if(_zz_3860_)begin
        int_reg_array_55_46_imag <= _zz_3880_;
      end
      if(_zz_3861_)begin
        int_reg_array_55_47_imag <= _zz_3880_;
      end
      if(_zz_3862_)begin
        int_reg_array_55_48_imag <= _zz_3880_;
      end
      if(_zz_3863_)begin
        int_reg_array_55_49_imag <= _zz_3880_;
      end
      if(_zz_3864_)begin
        int_reg_array_55_50_imag <= _zz_3880_;
      end
      if(_zz_3865_)begin
        int_reg_array_55_51_imag <= _zz_3880_;
      end
      if(_zz_3866_)begin
        int_reg_array_55_52_imag <= _zz_3880_;
      end
      if(_zz_3867_)begin
        int_reg_array_55_53_imag <= _zz_3880_;
      end
      if(_zz_3868_)begin
        int_reg_array_55_54_imag <= _zz_3880_;
      end
      if(_zz_3869_)begin
        int_reg_array_55_55_imag <= _zz_3880_;
      end
      if(_zz_3870_)begin
        int_reg_array_55_56_imag <= _zz_3880_;
      end
      if(_zz_3871_)begin
        int_reg_array_55_57_imag <= _zz_3880_;
      end
      if(_zz_3872_)begin
        int_reg_array_55_58_imag <= _zz_3880_;
      end
      if(_zz_3873_)begin
        int_reg_array_55_59_imag <= _zz_3880_;
      end
      if(_zz_3874_)begin
        int_reg_array_55_60_imag <= _zz_3880_;
      end
      if(_zz_3875_)begin
        int_reg_array_55_61_imag <= _zz_3880_;
      end
      if(_zz_3876_)begin
        int_reg_array_55_62_imag <= _zz_3880_;
      end
      if(_zz_3877_)begin
        int_reg_array_55_63_imag <= _zz_3880_;
      end
      if(_zz_3883_)begin
        int_reg_array_56_0_real <= _zz_3948_;
      end
      if(_zz_3884_)begin
        int_reg_array_56_1_real <= _zz_3948_;
      end
      if(_zz_3885_)begin
        int_reg_array_56_2_real <= _zz_3948_;
      end
      if(_zz_3886_)begin
        int_reg_array_56_3_real <= _zz_3948_;
      end
      if(_zz_3887_)begin
        int_reg_array_56_4_real <= _zz_3948_;
      end
      if(_zz_3888_)begin
        int_reg_array_56_5_real <= _zz_3948_;
      end
      if(_zz_3889_)begin
        int_reg_array_56_6_real <= _zz_3948_;
      end
      if(_zz_3890_)begin
        int_reg_array_56_7_real <= _zz_3948_;
      end
      if(_zz_3891_)begin
        int_reg_array_56_8_real <= _zz_3948_;
      end
      if(_zz_3892_)begin
        int_reg_array_56_9_real <= _zz_3948_;
      end
      if(_zz_3893_)begin
        int_reg_array_56_10_real <= _zz_3948_;
      end
      if(_zz_3894_)begin
        int_reg_array_56_11_real <= _zz_3948_;
      end
      if(_zz_3895_)begin
        int_reg_array_56_12_real <= _zz_3948_;
      end
      if(_zz_3896_)begin
        int_reg_array_56_13_real <= _zz_3948_;
      end
      if(_zz_3897_)begin
        int_reg_array_56_14_real <= _zz_3948_;
      end
      if(_zz_3898_)begin
        int_reg_array_56_15_real <= _zz_3948_;
      end
      if(_zz_3899_)begin
        int_reg_array_56_16_real <= _zz_3948_;
      end
      if(_zz_3900_)begin
        int_reg_array_56_17_real <= _zz_3948_;
      end
      if(_zz_3901_)begin
        int_reg_array_56_18_real <= _zz_3948_;
      end
      if(_zz_3902_)begin
        int_reg_array_56_19_real <= _zz_3948_;
      end
      if(_zz_3903_)begin
        int_reg_array_56_20_real <= _zz_3948_;
      end
      if(_zz_3904_)begin
        int_reg_array_56_21_real <= _zz_3948_;
      end
      if(_zz_3905_)begin
        int_reg_array_56_22_real <= _zz_3948_;
      end
      if(_zz_3906_)begin
        int_reg_array_56_23_real <= _zz_3948_;
      end
      if(_zz_3907_)begin
        int_reg_array_56_24_real <= _zz_3948_;
      end
      if(_zz_3908_)begin
        int_reg_array_56_25_real <= _zz_3948_;
      end
      if(_zz_3909_)begin
        int_reg_array_56_26_real <= _zz_3948_;
      end
      if(_zz_3910_)begin
        int_reg_array_56_27_real <= _zz_3948_;
      end
      if(_zz_3911_)begin
        int_reg_array_56_28_real <= _zz_3948_;
      end
      if(_zz_3912_)begin
        int_reg_array_56_29_real <= _zz_3948_;
      end
      if(_zz_3913_)begin
        int_reg_array_56_30_real <= _zz_3948_;
      end
      if(_zz_3914_)begin
        int_reg_array_56_31_real <= _zz_3948_;
      end
      if(_zz_3915_)begin
        int_reg_array_56_32_real <= _zz_3948_;
      end
      if(_zz_3916_)begin
        int_reg_array_56_33_real <= _zz_3948_;
      end
      if(_zz_3917_)begin
        int_reg_array_56_34_real <= _zz_3948_;
      end
      if(_zz_3918_)begin
        int_reg_array_56_35_real <= _zz_3948_;
      end
      if(_zz_3919_)begin
        int_reg_array_56_36_real <= _zz_3948_;
      end
      if(_zz_3920_)begin
        int_reg_array_56_37_real <= _zz_3948_;
      end
      if(_zz_3921_)begin
        int_reg_array_56_38_real <= _zz_3948_;
      end
      if(_zz_3922_)begin
        int_reg_array_56_39_real <= _zz_3948_;
      end
      if(_zz_3923_)begin
        int_reg_array_56_40_real <= _zz_3948_;
      end
      if(_zz_3924_)begin
        int_reg_array_56_41_real <= _zz_3948_;
      end
      if(_zz_3925_)begin
        int_reg_array_56_42_real <= _zz_3948_;
      end
      if(_zz_3926_)begin
        int_reg_array_56_43_real <= _zz_3948_;
      end
      if(_zz_3927_)begin
        int_reg_array_56_44_real <= _zz_3948_;
      end
      if(_zz_3928_)begin
        int_reg_array_56_45_real <= _zz_3948_;
      end
      if(_zz_3929_)begin
        int_reg_array_56_46_real <= _zz_3948_;
      end
      if(_zz_3930_)begin
        int_reg_array_56_47_real <= _zz_3948_;
      end
      if(_zz_3931_)begin
        int_reg_array_56_48_real <= _zz_3948_;
      end
      if(_zz_3932_)begin
        int_reg_array_56_49_real <= _zz_3948_;
      end
      if(_zz_3933_)begin
        int_reg_array_56_50_real <= _zz_3948_;
      end
      if(_zz_3934_)begin
        int_reg_array_56_51_real <= _zz_3948_;
      end
      if(_zz_3935_)begin
        int_reg_array_56_52_real <= _zz_3948_;
      end
      if(_zz_3936_)begin
        int_reg_array_56_53_real <= _zz_3948_;
      end
      if(_zz_3937_)begin
        int_reg_array_56_54_real <= _zz_3948_;
      end
      if(_zz_3938_)begin
        int_reg_array_56_55_real <= _zz_3948_;
      end
      if(_zz_3939_)begin
        int_reg_array_56_56_real <= _zz_3948_;
      end
      if(_zz_3940_)begin
        int_reg_array_56_57_real <= _zz_3948_;
      end
      if(_zz_3941_)begin
        int_reg_array_56_58_real <= _zz_3948_;
      end
      if(_zz_3942_)begin
        int_reg_array_56_59_real <= _zz_3948_;
      end
      if(_zz_3943_)begin
        int_reg_array_56_60_real <= _zz_3948_;
      end
      if(_zz_3944_)begin
        int_reg_array_56_61_real <= _zz_3948_;
      end
      if(_zz_3945_)begin
        int_reg_array_56_62_real <= _zz_3948_;
      end
      if(_zz_3946_)begin
        int_reg_array_56_63_real <= _zz_3948_;
      end
      if(_zz_3883_)begin
        int_reg_array_56_0_imag <= _zz_3949_;
      end
      if(_zz_3884_)begin
        int_reg_array_56_1_imag <= _zz_3949_;
      end
      if(_zz_3885_)begin
        int_reg_array_56_2_imag <= _zz_3949_;
      end
      if(_zz_3886_)begin
        int_reg_array_56_3_imag <= _zz_3949_;
      end
      if(_zz_3887_)begin
        int_reg_array_56_4_imag <= _zz_3949_;
      end
      if(_zz_3888_)begin
        int_reg_array_56_5_imag <= _zz_3949_;
      end
      if(_zz_3889_)begin
        int_reg_array_56_6_imag <= _zz_3949_;
      end
      if(_zz_3890_)begin
        int_reg_array_56_7_imag <= _zz_3949_;
      end
      if(_zz_3891_)begin
        int_reg_array_56_8_imag <= _zz_3949_;
      end
      if(_zz_3892_)begin
        int_reg_array_56_9_imag <= _zz_3949_;
      end
      if(_zz_3893_)begin
        int_reg_array_56_10_imag <= _zz_3949_;
      end
      if(_zz_3894_)begin
        int_reg_array_56_11_imag <= _zz_3949_;
      end
      if(_zz_3895_)begin
        int_reg_array_56_12_imag <= _zz_3949_;
      end
      if(_zz_3896_)begin
        int_reg_array_56_13_imag <= _zz_3949_;
      end
      if(_zz_3897_)begin
        int_reg_array_56_14_imag <= _zz_3949_;
      end
      if(_zz_3898_)begin
        int_reg_array_56_15_imag <= _zz_3949_;
      end
      if(_zz_3899_)begin
        int_reg_array_56_16_imag <= _zz_3949_;
      end
      if(_zz_3900_)begin
        int_reg_array_56_17_imag <= _zz_3949_;
      end
      if(_zz_3901_)begin
        int_reg_array_56_18_imag <= _zz_3949_;
      end
      if(_zz_3902_)begin
        int_reg_array_56_19_imag <= _zz_3949_;
      end
      if(_zz_3903_)begin
        int_reg_array_56_20_imag <= _zz_3949_;
      end
      if(_zz_3904_)begin
        int_reg_array_56_21_imag <= _zz_3949_;
      end
      if(_zz_3905_)begin
        int_reg_array_56_22_imag <= _zz_3949_;
      end
      if(_zz_3906_)begin
        int_reg_array_56_23_imag <= _zz_3949_;
      end
      if(_zz_3907_)begin
        int_reg_array_56_24_imag <= _zz_3949_;
      end
      if(_zz_3908_)begin
        int_reg_array_56_25_imag <= _zz_3949_;
      end
      if(_zz_3909_)begin
        int_reg_array_56_26_imag <= _zz_3949_;
      end
      if(_zz_3910_)begin
        int_reg_array_56_27_imag <= _zz_3949_;
      end
      if(_zz_3911_)begin
        int_reg_array_56_28_imag <= _zz_3949_;
      end
      if(_zz_3912_)begin
        int_reg_array_56_29_imag <= _zz_3949_;
      end
      if(_zz_3913_)begin
        int_reg_array_56_30_imag <= _zz_3949_;
      end
      if(_zz_3914_)begin
        int_reg_array_56_31_imag <= _zz_3949_;
      end
      if(_zz_3915_)begin
        int_reg_array_56_32_imag <= _zz_3949_;
      end
      if(_zz_3916_)begin
        int_reg_array_56_33_imag <= _zz_3949_;
      end
      if(_zz_3917_)begin
        int_reg_array_56_34_imag <= _zz_3949_;
      end
      if(_zz_3918_)begin
        int_reg_array_56_35_imag <= _zz_3949_;
      end
      if(_zz_3919_)begin
        int_reg_array_56_36_imag <= _zz_3949_;
      end
      if(_zz_3920_)begin
        int_reg_array_56_37_imag <= _zz_3949_;
      end
      if(_zz_3921_)begin
        int_reg_array_56_38_imag <= _zz_3949_;
      end
      if(_zz_3922_)begin
        int_reg_array_56_39_imag <= _zz_3949_;
      end
      if(_zz_3923_)begin
        int_reg_array_56_40_imag <= _zz_3949_;
      end
      if(_zz_3924_)begin
        int_reg_array_56_41_imag <= _zz_3949_;
      end
      if(_zz_3925_)begin
        int_reg_array_56_42_imag <= _zz_3949_;
      end
      if(_zz_3926_)begin
        int_reg_array_56_43_imag <= _zz_3949_;
      end
      if(_zz_3927_)begin
        int_reg_array_56_44_imag <= _zz_3949_;
      end
      if(_zz_3928_)begin
        int_reg_array_56_45_imag <= _zz_3949_;
      end
      if(_zz_3929_)begin
        int_reg_array_56_46_imag <= _zz_3949_;
      end
      if(_zz_3930_)begin
        int_reg_array_56_47_imag <= _zz_3949_;
      end
      if(_zz_3931_)begin
        int_reg_array_56_48_imag <= _zz_3949_;
      end
      if(_zz_3932_)begin
        int_reg_array_56_49_imag <= _zz_3949_;
      end
      if(_zz_3933_)begin
        int_reg_array_56_50_imag <= _zz_3949_;
      end
      if(_zz_3934_)begin
        int_reg_array_56_51_imag <= _zz_3949_;
      end
      if(_zz_3935_)begin
        int_reg_array_56_52_imag <= _zz_3949_;
      end
      if(_zz_3936_)begin
        int_reg_array_56_53_imag <= _zz_3949_;
      end
      if(_zz_3937_)begin
        int_reg_array_56_54_imag <= _zz_3949_;
      end
      if(_zz_3938_)begin
        int_reg_array_56_55_imag <= _zz_3949_;
      end
      if(_zz_3939_)begin
        int_reg_array_56_56_imag <= _zz_3949_;
      end
      if(_zz_3940_)begin
        int_reg_array_56_57_imag <= _zz_3949_;
      end
      if(_zz_3941_)begin
        int_reg_array_56_58_imag <= _zz_3949_;
      end
      if(_zz_3942_)begin
        int_reg_array_56_59_imag <= _zz_3949_;
      end
      if(_zz_3943_)begin
        int_reg_array_56_60_imag <= _zz_3949_;
      end
      if(_zz_3944_)begin
        int_reg_array_56_61_imag <= _zz_3949_;
      end
      if(_zz_3945_)begin
        int_reg_array_56_62_imag <= _zz_3949_;
      end
      if(_zz_3946_)begin
        int_reg_array_56_63_imag <= _zz_3949_;
      end
      if(_zz_3952_)begin
        int_reg_array_57_0_real <= _zz_4017_;
      end
      if(_zz_3953_)begin
        int_reg_array_57_1_real <= _zz_4017_;
      end
      if(_zz_3954_)begin
        int_reg_array_57_2_real <= _zz_4017_;
      end
      if(_zz_3955_)begin
        int_reg_array_57_3_real <= _zz_4017_;
      end
      if(_zz_3956_)begin
        int_reg_array_57_4_real <= _zz_4017_;
      end
      if(_zz_3957_)begin
        int_reg_array_57_5_real <= _zz_4017_;
      end
      if(_zz_3958_)begin
        int_reg_array_57_6_real <= _zz_4017_;
      end
      if(_zz_3959_)begin
        int_reg_array_57_7_real <= _zz_4017_;
      end
      if(_zz_3960_)begin
        int_reg_array_57_8_real <= _zz_4017_;
      end
      if(_zz_3961_)begin
        int_reg_array_57_9_real <= _zz_4017_;
      end
      if(_zz_3962_)begin
        int_reg_array_57_10_real <= _zz_4017_;
      end
      if(_zz_3963_)begin
        int_reg_array_57_11_real <= _zz_4017_;
      end
      if(_zz_3964_)begin
        int_reg_array_57_12_real <= _zz_4017_;
      end
      if(_zz_3965_)begin
        int_reg_array_57_13_real <= _zz_4017_;
      end
      if(_zz_3966_)begin
        int_reg_array_57_14_real <= _zz_4017_;
      end
      if(_zz_3967_)begin
        int_reg_array_57_15_real <= _zz_4017_;
      end
      if(_zz_3968_)begin
        int_reg_array_57_16_real <= _zz_4017_;
      end
      if(_zz_3969_)begin
        int_reg_array_57_17_real <= _zz_4017_;
      end
      if(_zz_3970_)begin
        int_reg_array_57_18_real <= _zz_4017_;
      end
      if(_zz_3971_)begin
        int_reg_array_57_19_real <= _zz_4017_;
      end
      if(_zz_3972_)begin
        int_reg_array_57_20_real <= _zz_4017_;
      end
      if(_zz_3973_)begin
        int_reg_array_57_21_real <= _zz_4017_;
      end
      if(_zz_3974_)begin
        int_reg_array_57_22_real <= _zz_4017_;
      end
      if(_zz_3975_)begin
        int_reg_array_57_23_real <= _zz_4017_;
      end
      if(_zz_3976_)begin
        int_reg_array_57_24_real <= _zz_4017_;
      end
      if(_zz_3977_)begin
        int_reg_array_57_25_real <= _zz_4017_;
      end
      if(_zz_3978_)begin
        int_reg_array_57_26_real <= _zz_4017_;
      end
      if(_zz_3979_)begin
        int_reg_array_57_27_real <= _zz_4017_;
      end
      if(_zz_3980_)begin
        int_reg_array_57_28_real <= _zz_4017_;
      end
      if(_zz_3981_)begin
        int_reg_array_57_29_real <= _zz_4017_;
      end
      if(_zz_3982_)begin
        int_reg_array_57_30_real <= _zz_4017_;
      end
      if(_zz_3983_)begin
        int_reg_array_57_31_real <= _zz_4017_;
      end
      if(_zz_3984_)begin
        int_reg_array_57_32_real <= _zz_4017_;
      end
      if(_zz_3985_)begin
        int_reg_array_57_33_real <= _zz_4017_;
      end
      if(_zz_3986_)begin
        int_reg_array_57_34_real <= _zz_4017_;
      end
      if(_zz_3987_)begin
        int_reg_array_57_35_real <= _zz_4017_;
      end
      if(_zz_3988_)begin
        int_reg_array_57_36_real <= _zz_4017_;
      end
      if(_zz_3989_)begin
        int_reg_array_57_37_real <= _zz_4017_;
      end
      if(_zz_3990_)begin
        int_reg_array_57_38_real <= _zz_4017_;
      end
      if(_zz_3991_)begin
        int_reg_array_57_39_real <= _zz_4017_;
      end
      if(_zz_3992_)begin
        int_reg_array_57_40_real <= _zz_4017_;
      end
      if(_zz_3993_)begin
        int_reg_array_57_41_real <= _zz_4017_;
      end
      if(_zz_3994_)begin
        int_reg_array_57_42_real <= _zz_4017_;
      end
      if(_zz_3995_)begin
        int_reg_array_57_43_real <= _zz_4017_;
      end
      if(_zz_3996_)begin
        int_reg_array_57_44_real <= _zz_4017_;
      end
      if(_zz_3997_)begin
        int_reg_array_57_45_real <= _zz_4017_;
      end
      if(_zz_3998_)begin
        int_reg_array_57_46_real <= _zz_4017_;
      end
      if(_zz_3999_)begin
        int_reg_array_57_47_real <= _zz_4017_;
      end
      if(_zz_4000_)begin
        int_reg_array_57_48_real <= _zz_4017_;
      end
      if(_zz_4001_)begin
        int_reg_array_57_49_real <= _zz_4017_;
      end
      if(_zz_4002_)begin
        int_reg_array_57_50_real <= _zz_4017_;
      end
      if(_zz_4003_)begin
        int_reg_array_57_51_real <= _zz_4017_;
      end
      if(_zz_4004_)begin
        int_reg_array_57_52_real <= _zz_4017_;
      end
      if(_zz_4005_)begin
        int_reg_array_57_53_real <= _zz_4017_;
      end
      if(_zz_4006_)begin
        int_reg_array_57_54_real <= _zz_4017_;
      end
      if(_zz_4007_)begin
        int_reg_array_57_55_real <= _zz_4017_;
      end
      if(_zz_4008_)begin
        int_reg_array_57_56_real <= _zz_4017_;
      end
      if(_zz_4009_)begin
        int_reg_array_57_57_real <= _zz_4017_;
      end
      if(_zz_4010_)begin
        int_reg_array_57_58_real <= _zz_4017_;
      end
      if(_zz_4011_)begin
        int_reg_array_57_59_real <= _zz_4017_;
      end
      if(_zz_4012_)begin
        int_reg_array_57_60_real <= _zz_4017_;
      end
      if(_zz_4013_)begin
        int_reg_array_57_61_real <= _zz_4017_;
      end
      if(_zz_4014_)begin
        int_reg_array_57_62_real <= _zz_4017_;
      end
      if(_zz_4015_)begin
        int_reg_array_57_63_real <= _zz_4017_;
      end
      if(_zz_3952_)begin
        int_reg_array_57_0_imag <= _zz_4018_;
      end
      if(_zz_3953_)begin
        int_reg_array_57_1_imag <= _zz_4018_;
      end
      if(_zz_3954_)begin
        int_reg_array_57_2_imag <= _zz_4018_;
      end
      if(_zz_3955_)begin
        int_reg_array_57_3_imag <= _zz_4018_;
      end
      if(_zz_3956_)begin
        int_reg_array_57_4_imag <= _zz_4018_;
      end
      if(_zz_3957_)begin
        int_reg_array_57_5_imag <= _zz_4018_;
      end
      if(_zz_3958_)begin
        int_reg_array_57_6_imag <= _zz_4018_;
      end
      if(_zz_3959_)begin
        int_reg_array_57_7_imag <= _zz_4018_;
      end
      if(_zz_3960_)begin
        int_reg_array_57_8_imag <= _zz_4018_;
      end
      if(_zz_3961_)begin
        int_reg_array_57_9_imag <= _zz_4018_;
      end
      if(_zz_3962_)begin
        int_reg_array_57_10_imag <= _zz_4018_;
      end
      if(_zz_3963_)begin
        int_reg_array_57_11_imag <= _zz_4018_;
      end
      if(_zz_3964_)begin
        int_reg_array_57_12_imag <= _zz_4018_;
      end
      if(_zz_3965_)begin
        int_reg_array_57_13_imag <= _zz_4018_;
      end
      if(_zz_3966_)begin
        int_reg_array_57_14_imag <= _zz_4018_;
      end
      if(_zz_3967_)begin
        int_reg_array_57_15_imag <= _zz_4018_;
      end
      if(_zz_3968_)begin
        int_reg_array_57_16_imag <= _zz_4018_;
      end
      if(_zz_3969_)begin
        int_reg_array_57_17_imag <= _zz_4018_;
      end
      if(_zz_3970_)begin
        int_reg_array_57_18_imag <= _zz_4018_;
      end
      if(_zz_3971_)begin
        int_reg_array_57_19_imag <= _zz_4018_;
      end
      if(_zz_3972_)begin
        int_reg_array_57_20_imag <= _zz_4018_;
      end
      if(_zz_3973_)begin
        int_reg_array_57_21_imag <= _zz_4018_;
      end
      if(_zz_3974_)begin
        int_reg_array_57_22_imag <= _zz_4018_;
      end
      if(_zz_3975_)begin
        int_reg_array_57_23_imag <= _zz_4018_;
      end
      if(_zz_3976_)begin
        int_reg_array_57_24_imag <= _zz_4018_;
      end
      if(_zz_3977_)begin
        int_reg_array_57_25_imag <= _zz_4018_;
      end
      if(_zz_3978_)begin
        int_reg_array_57_26_imag <= _zz_4018_;
      end
      if(_zz_3979_)begin
        int_reg_array_57_27_imag <= _zz_4018_;
      end
      if(_zz_3980_)begin
        int_reg_array_57_28_imag <= _zz_4018_;
      end
      if(_zz_3981_)begin
        int_reg_array_57_29_imag <= _zz_4018_;
      end
      if(_zz_3982_)begin
        int_reg_array_57_30_imag <= _zz_4018_;
      end
      if(_zz_3983_)begin
        int_reg_array_57_31_imag <= _zz_4018_;
      end
      if(_zz_3984_)begin
        int_reg_array_57_32_imag <= _zz_4018_;
      end
      if(_zz_3985_)begin
        int_reg_array_57_33_imag <= _zz_4018_;
      end
      if(_zz_3986_)begin
        int_reg_array_57_34_imag <= _zz_4018_;
      end
      if(_zz_3987_)begin
        int_reg_array_57_35_imag <= _zz_4018_;
      end
      if(_zz_3988_)begin
        int_reg_array_57_36_imag <= _zz_4018_;
      end
      if(_zz_3989_)begin
        int_reg_array_57_37_imag <= _zz_4018_;
      end
      if(_zz_3990_)begin
        int_reg_array_57_38_imag <= _zz_4018_;
      end
      if(_zz_3991_)begin
        int_reg_array_57_39_imag <= _zz_4018_;
      end
      if(_zz_3992_)begin
        int_reg_array_57_40_imag <= _zz_4018_;
      end
      if(_zz_3993_)begin
        int_reg_array_57_41_imag <= _zz_4018_;
      end
      if(_zz_3994_)begin
        int_reg_array_57_42_imag <= _zz_4018_;
      end
      if(_zz_3995_)begin
        int_reg_array_57_43_imag <= _zz_4018_;
      end
      if(_zz_3996_)begin
        int_reg_array_57_44_imag <= _zz_4018_;
      end
      if(_zz_3997_)begin
        int_reg_array_57_45_imag <= _zz_4018_;
      end
      if(_zz_3998_)begin
        int_reg_array_57_46_imag <= _zz_4018_;
      end
      if(_zz_3999_)begin
        int_reg_array_57_47_imag <= _zz_4018_;
      end
      if(_zz_4000_)begin
        int_reg_array_57_48_imag <= _zz_4018_;
      end
      if(_zz_4001_)begin
        int_reg_array_57_49_imag <= _zz_4018_;
      end
      if(_zz_4002_)begin
        int_reg_array_57_50_imag <= _zz_4018_;
      end
      if(_zz_4003_)begin
        int_reg_array_57_51_imag <= _zz_4018_;
      end
      if(_zz_4004_)begin
        int_reg_array_57_52_imag <= _zz_4018_;
      end
      if(_zz_4005_)begin
        int_reg_array_57_53_imag <= _zz_4018_;
      end
      if(_zz_4006_)begin
        int_reg_array_57_54_imag <= _zz_4018_;
      end
      if(_zz_4007_)begin
        int_reg_array_57_55_imag <= _zz_4018_;
      end
      if(_zz_4008_)begin
        int_reg_array_57_56_imag <= _zz_4018_;
      end
      if(_zz_4009_)begin
        int_reg_array_57_57_imag <= _zz_4018_;
      end
      if(_zz_4010_)begin
        int_reg_array_57_58_imag <= _zz_4018_;
      end
      if(_zz_4011_)begin
        int_reg_array_57_59_imag <= _zz_4018_;
      end
      if(_zz_4012_)begin
        int_reg_array_57_60_imag <= _zz_4018_;
      end
      if(_zz_4013_)begin
        int_reg_array_57_61_imag <= _zz_4018_;
      end
      if(_zz_4014_)begin
        int_reg_array_57_62_imag <= _zz_4018_;
      end
      if(_zz_4015_)begin
        int_reg_array_57_63_imag <= _zz_4018_;
      end
      if(_zz_4021_)begin
        int_reg_array_58_0_real <= _zz_4086_;
      end
      if(_zz_4022_)begin
        int_reg_array_58_1_real <= _zz_4086_;
      end
      if(_zz_4023_)begin
        int_reg_array_58_2_real <= _zz_4086_;
      end
      if(_zz_4024_)begin
        int_reg_array_58_3_real <= _zz_4086_;
      end
      if(_zz_4025_)begin
        int_reg_array_58_4_real <= _zz_4086_;
      end
      if(_zz_4026_)begin
        int_reg_array_58_5_real <= _zz_4086_;
      end
      if(_zz_4027_)begin
        int_reg_array_58_6_real <= _zz_4086_;
      end
      if(_zz_4028_)begin
        int_reg_array_58_7_real <= _zz_4086_;
      end
      if(_zz_4029_)begin
        int_reg_array_58_8_real <= _zz_4086_;
      end
      if(_zz_4030_)begin
        int_reg_array_58_9_real <= _zz_4086_;
      end
      if(_zz_4031_)begin
        int_reg_array_58_10_real <= _zz_4086_;
      end
      if(_zz_4032_)begin
        int_reg_array_58_11_real <= _zz_4086_;
      end
      if(_zz_4033_)begin
        int_reg_array_58_12_real <= _zz_4086_;
      end
      if(_zz_4034_)begin
        int_reg_array_58_13_real <= _zz_4086_;
      end
      if(_zz_4035_)begin
        int_reg_array_58_14_real <= _zz_4086_;
      end
      if(_zz_4036_)begin
        int_reg_array_58_15_real <= _zz_4086_;
      end
      if(_zz_4037_)begin
        int_reg_array_58_16_real <= _zz_4086_;
      end
      if(_zz_4038_)begin
        int_reg_array_58_17_real <= _zz_4086_;
      end
      if(_zz_4039_)begin
        int_reg_array_58_18_real <= _zz_4086_;
      end
      if(_zz_4040_)begin
        int_reg_array_58_19_real <= _zz_4086_;
      end
      if(_zz_4041_)begin
        int_reg_array_58_20_real <= _zz_4086_;
      end
      if(_zz_4042_)begin
        int_reg_array_58_21_real <= _zz_4086_;
      end
      if(_zz_4043_)begin
        int_reg_array_58_22_real <= _zz_4086_;
      end
      if(_zz_4044_)begin
        int_reg_array_58_23_real <= _zz_4086_;
      end
      if(_zz_4045_)begin
        int_reg_array_58_24_real <= _zz_4086_;
      end
      if(_zz_4046_)begin
        int_reg_array_58_25_real <= _zz_4086_;
      end
      if(_zz_4047_)begin
        int_reg_array_58_26_real <= _zz_4086_;
      end
      if(_zz_4048_)begin
        int_reg_array_58_27_real <= _zz_4086_;
      end
      if(_zz_4049_)begin
        int_reg_array_58_28_real <= _zz_4086_;
      end
      if(_zz_4050_)begin
        int_reg_array_58_29_real <= _zz_4086_;
      end
      if(_zz_4051_)begin
        int_reg_array_58_30_real <= _zz_4086_;
      end
      if(_zz_4052_)begin
        int_reg_array_58_31_real <= _zz_4086_;
      end
      if(_zz_4053_)begin
        int_reg_array_58_32_real <= _zz_4086_;
      end
      if(_zz_4054_)begin
        int_reg_array_58_33_real <= _zz_4086_;
      end
      if(_zz_4055_)begin
        int_reg_array_58_34_real <= _zz_4086_;
      end
      if(_zz_4056_)begin
        int_reg_array_58_35_real <= _zz_4086_;
      end
      if(_zz_4057_)begin
        int_reg_array_58_36_real <= _zz_4086_;
      end
      if(_zz_4058_)begin
        int_reg_array_58_37_real <= _zz_4086_;
      end
      if(_zz_4059_)begin
        int_reg_array_58_38_real <= _zz_4086_;
      end
      if(_zz_4060_)begin
        int_reg_array_58_39_real <= _zz_4086_;
      end
      if(_zz_4061_)begin
        int_reg_array_58_40_real <= _zz_4086_;
      end
      if(_zz_4062_)begin
        int_reg_array_58_41_real <= _zz_4086_;
      end
      if(_zz_4063_)begin
        int_reg_array_58_42_real <= _zz_4086_;
      end
      if(_zz_4064_)begin
        int_reg_array_58_43_real <= _zz_4086_;
      end
      if(_zz_4065_)begin
        int_reg_array_58_44_real <= _zz_4086_;
      end
      if(_zz_4066_)begin
        int_reg_array_58_45_real <= _zz_4086_;
      end
      if(_zz_4067_)begin
        int_reg_array_58_46_real <= _zz_4086_;
      end
      if(_zz_4068_)begin
        int_reg_array_58_47_real <= _zz_4086_;
      end
      if(_zz_4069_)begin
        int_reg_array_58_48_real <= _zz_4086_;
      end
      if(_zz_4070_)begin
        int_reg_array_58_49_real <= _zz_4086_;
      end
      if(_zz_4071_)begin
        int_reg_array_58_50_real <= _zz_4086_;
      end
      if(_zz_4072_)begin
        int_reg_array_58_51_real <= _zz_4086_;
      end
      if(_zz_4073_)begin
        int_reg_array_58_52_real <= _zz_4086_;
      end
      if(_zz_4074_)begin
        int_reg_array_58_53_real <= _zz_4086_;
      end
      if(_zz_4075_)begin
        int_reg_array_58_54_real <= _zz_4086_;
      end
      if(_zz_4076_)begin
        int_reg_array_58_55_real <= _zz_4086_;
      end
      if(_zz_4077_)begin
        int_reg_array_58_56_real <= _zz_4086_;
      end
      if(_zz_4078_)begin
        int_reg_array_58_57_real <= _zz_4086_;
      end
      if(_zz_4079_)begin
        int_reg_array_58_58_real <= _zz_4086_;
      end
      if(_zz_4080_)begin
        int_reg_array_58_59_real <= _zz_4086_;
      end
      if(_zz_4081_)begin
        int_reg_array_58_60_real <= _zz_4086_;
      end
      if(_zz_4082_)begin
        int_reg_array_58_61_real <= _zz_4086_;
      end
      if(_zz_4083_)begin
        int_reg_array_58_62_real <= _zz_4086_;
      end
      if(_zz_4084_)begin
        int_reg_array_58_63_real <= _zz_4086_;
      end
      if(_zz_4021_)begin
        int_reg_array_58_0_imag <= _zz_4087_;
      end
      if(_zz_4022_)begin
        int_reg_array_58_1_imag <= _zz_4087_;
      end
      if(_zz_4023_)begin
        int_reg_array_58_2_imag <= _zz_4087_;
      end
      if(_zz_4024_)begin
        int_reg_array_58_3_imag <= _zz_4087_;
      end
      if(_zz_4025_)begin
        int_reg_array_58_4_imag <= _zz_4087_;
      end
      if(_zz_4026_)begin
        int_reg_array_58_5_imag <= _zz_4087_;
      end
      if(_zz_4027_)begin
        int_reg_array_58_6_imag <= _zz_4087_;
      end
      if(_zz_4028_)begin
        int_reg_array_58_7_imag <= _zz_4087_;
      end
      if(_zz_4029_)begin
        int_reg_array_58_8_imag <= _zz_4087_;
      end
      if(_zz_4030_)begin
        int_reg_array_58_9_imag <= _zz_4087_;
      end
      if(_zz_4031_)begin
        int_reg_array_58_10_imag <= _zz_4087_;
      end
      if(_zz_4032_)begin
        int_reg_array_58_11_imag <= _zz_4087_;
      end
      if(_zz_4033_)begin
        int_reg_array_58_12_imag <= _zz_4087_;
      end
      if(_zz_4034_)begin
        int_reg_array_58_13_imag <= _zz_4087_;
      end
      if(_zz_4035_)begin
        int_reg_array_58_14_imag <= _zz_4087_;
      end
      if(_zz_4036_)begin
        int_reg_array_58_15_imag <= _zz_4087_;
      end
      if(_zz_4037_)begin
        int_reg_array_58_16_imag <= _zz_4087_;
      end
      if(_zz_4038_)begin
        int_reg_array_58_17_imag <= _zz_4087_;
      end
      if(_zz_4039_)begin
        int_reg_array_58_18_imag <= _zz_4087_;
      end
      if(_zz_4040_)begin
        int_reg_array_58_19_imag <= _zz_4087_;
      end
      if(_zz_4041_)begin
        int_reg_array_58_20_imag <= _zz_4087_;
      end
      if(_zz_4042_)begin
        int_reg_array_58_21_imag <= _zz_4087_;
      end
      if(_zz_4043_)begin
        int_reg_array_58_22_imag <= _zz_4087_;
      end
      if(_zz_4044_)begin
        int_reg_array_58_23_imag <= _zz_4087_;
      end
      if(_zz_4045_)begin
        int_reg_array_58_24_imag <= _zz_4087_;
      end
      if(_zz_4046_)begin
        int_reg_array_58_25_imag <= _zz_4087_;
      end
      if(_zz_4047_)begin
        int_reg_array_58_26_imag <= _zz_4087_;
      end
      if(_zz_4048_)begin
        int_reg_array_58_27_imag <= _zz_4087_;
      end
      if(_zz_4049_)begin
        int_reg_array_58_28_imag <= _zz_4087_;
      end
      if(_zz_4050_)begin
        int_reg_array_58_29_imag <= _zz_4087_;
      end
      if(_zz_4051_)begin
        int_reg_array_58_30_imag <= _zz_4087_;
      end
      if(_zz_4052_)begin
        int_reg_array_58_31_imag <= _zz_4087_;
      end
      if(_zz_4053_)begin
        int_reg_array_58_32_imag <= _zz_4087_;
      end
      if(_zz_4054_)begin
        int_reg_array_58_33_imag <= _zz_4087_;
      end
      if(_zz_4055_)begin
        int_reg_array_58_34_imag <= _zz_4087_;
      end
      if(_zz_4056_)begin
        int_reg_array_58_35_imag <= _zz_4087_;
      end
      if(_zz_4057_)begin
        int_reg_array_58_36_imag <= _zz_4087_;
      end
      if(_zz_4058_)begin
        int_reg_array_58_37_imag <= _zz_4087_;
      end
      if(_zz_4059_)begin
        int_reg_array_58_38_imag <= _zz_4087_;
      end
      if(_zz_4060_)begin
        int_reg_array_58_39_imag <= _zz_4087_;
      end
      if(_zz_4061_)begin
        int_reg_array_58_40_imag <= _zz_4087_;
      end
      if(_zz_4062_)begin
        int_reg_array_58_41_imag <= _zz_4087_;
      end
      if(_zz_4063_)begin
        int_reg_array_58_42_imag <= _zz_4087_;
      end
      if(_zz_4064_)begin
        int_reg_array_58_43_imag <= _zz_4087_;
      end
      if(_zz_4065_)begin
        int_reg_array_58_44_imag <= _zz_4087_;
      end
      if(_zz_4066_)begin
        int_reg_array_58_45_imag <= _zz_4087_;
      end
      if(_zz_4067_)begin
        int_reg_array_58_46_imag <= _zz_4087_;
      end
      if(_zz_4068_)begin
        int_reg_array_58_47_imag <= _zz_4087_;
      end
      if(_zz_4069_)begin
        int_reg_array_58_48_imag <= _zz_4087_;
      end
      if(_zz_4070_)begin
        int_reg_array_58_49_imag <= _zz_4087_;
      end
      if(_zz_4071_)begin
        int_reg_array_58_50_imag <= _zz_4087_;
      end
      if(_zz_4072_)begin
        int_reg_array_58_51_imag <= _zz_4087_;
      end
      if(_zz_4073_)begin
        int_reg_array_58_52_imag <= _zz_4087_;
      end
      if(_zz_4074_)begin
        int_reg_array_58_53_imag <= _zz_4087_;
      end
      if(_zz_4075_)begin
        int_reg_array_58_54_imag <= _zz_4087_;
      end
      if(_zz_4076_)begin
        int_reg_array_58_55_imag <= _zz_4087_;
      end
      if(_zz_4077_)begin
        int_reg_array_58_56_imag <= _zz_4087_;
      end
      if(_zz_4078_)begin
        int_reg_array_58_57_imag <= _zz_4087_;
      end
      if(_zz_4079_)begin
        int_reg_array_58_58_imag <= _zz_4087_;
      end
      if(_zz_4080_)begin
        int_reg_array_58_59_imag <= _zz_4087_;
      end
      if(_zz_4081_)begin
        int_reg_array_58_60_imag <= _zz_4087_;
      end
      if(_zz_4082_)begin
        int_reg_array_58_61_imag <= _zz_4087_;
      end
      if(_zz_4083_)begin
        int_reg_array_58_62_imag <= _zz_4087_;
      end
      if(_zz_4084_)begin
        int_reg_array_58_63_imag <= _zz_4087_;
      end
      if(_zz_4090_)begin
        int_reg_array_59_0_real <= _zz_4155_;
      end
      if(_zz_4091_)begin
        int_reg_array_59_1_real <= _zz_4155_;
      end
      if(_zz_4092_)begin
        int_reg_array_59_2_real <= _zz_4155_;
      end
      if(_zz_4093_)begin
        int_reg_array_59_3_real <= _zz_4155_;
      end
      if(_zz_4094_)begin
        int_reg_array_59_4_real <= _zz_4155_;
      end
      if(_zz_4095_)begin
        int_reg_array_59_5_real <= _zz_4155_;
      end
      if(_zz_4096_)begin
        int_reg_array_59_6_real <= _zz_4155_;
      end
      if(_zz_4097_)begin
        int_reg_array_59_7_real <= _zz_4155_;
      end
      if(_zz_4098_)begin
        int_reg_array_59_8_real <= _zz_4155_;
      end
      if(_zz_4099_)begin
        int_reg_array_59_9_real <= _zz_4155_;
      end
      if(_zz_4100_)begin
        int_reg_array_59_10_real <= _zz_4155_;
      end
      if(_zz_4101_)begin
        int_reg_array_59_11_real <= _zz_4155_;
      end
      if(_zz_4102_)begin
        int_reg_array_59_12_real <= _zz_4155_;
      end
      if(_zz_4103_)begin
        int_reg_array_59_13_real <= _zz_4155_;
      end
      if(_zz_4104_)begin
        int_reg_array_59_14_real <= _zz_4155_;
      end
      if(_zz_4105_)begin
        int_reg_array_59_15_real <= _zz_4155_;
      end
      if(_zz_4106_)begin
        int_reg_array_59_16_real <= _zz_4155_;
      end
      if(_zz_4107_)begin
        int_reg_array_59_17_real <= _zz_4155_;
      end
      if(_zz_4108_)begin
        int_reg_array_59_18_real <= _zz_4155_;
      end
      if(_zz_4109_)begin
        int_reg_array_59_19_real <= _zz_4155_;
      end
      if(_zz_4110_)begin
        int_reg_array_59_20_real <= _zz_4155_;
      end
      if(_zz_4111_)begin
        int_reg_array_59_21_real <= _zz_4155_;
      end
      if(_zz_4112_)begin
        int_reg_array_59_22_real <= _zz_4155_;
      end
      if(_zz_4113_)begin
        int_reg_array_59_23_real <= _zz_4155_;
      end
      if(_zz_4114_)begin
        int_reg_array_59_24_real <= _zz_4155_;
      end
      if(_zz_4115_)begin
        int_reg_array_59_25_real <= _zz_4155_;
      end
      if(_zz_4116_)begin
        int_reg_array_59_26_real <= _zz_4155_;
      end
      if(_zz_4117_)begin
        int_reg_array_59_27_real <= _zz_4155_;
      end
      if(_zz_4118_)begin
        int_reg_array_59_28_real <= _zz_4155_;
      end
      if(_zz_4119_)begin
        int_reg_array_59_29_real <= _zz_4155_;
      end
      if(_zz_4120_)begin
        int_reg_array_59_30_real <= _zz_4155_;
      end
      if(_zz_4121_)begin
        int_reg_array_59_31_real <= _zz_4155_;
      end
      if(_zz_4122_)begin
        int_reg_array_59_32_real <= _zz_4155_;
      end
      if(_zz_4123_)begin
        int_reg_array_59_33_real <= _zz_4155_;
      end
      if(_zz_4124_)begin
        int_reg_array_59_34_real <= _zz_4155_;
      end
      if(_zz_4125_)begin
        int_reg_array_59_35_real <= _zz_4155_;
      end
      if(_zz_4126_)begin
        int_reg_array_59_36_real <= _zz_4155_;
      end
      if(_zz_4127_)begin
        int_reg_array_59_37_real <= _zz_4155_;
      end
      if(_zz_4128_)begin
        int_reg_array_59_38_real <= _zz_4155_;
      end
      if(_zz_4129_)begin
        int_reg_array_59_39_real <= _zz_4155_;
      end
      if(_zz_4130_)begin
        int_reg_array_59_40_real <= _zz_4155_;
      end
      if(_zz_4131_)begin
        int_reg_array_59_41_real <= _zz_4155_;
      end
      if(_zz_4132_)begin
        int_reg_array_59_42_real <= _zz_4155_;
      end
      if(_zz_4133_)begin
        int_reg_array_59_43_real <= _zz_4155_;
      end
      if(_zz_4134_)begin
        int_reg_array_59_44_real <= _zz_4155_;
      end
      if(_zz_4135_)begin
        int_reg_array_59_45_real <= _zz_4155_;
      end
      if(_zz_4136_)begin
        int_reg_array_59_46_real <= _zz_4155_;
      end
      if(_zz_4137_)begin
        int_reg_array_59_47_real <= _zz_4155_;
      end
      if(_zz_4138_)begin
        int_reg_array_59_48_real <= _zz_4155_;
      end
      if(_zz_4139_)begin
        int_reg_array_59_49_real <= _zz_4155_;
      end
      if(_zz_4140_)begin
        int_reg_array_59_50_real <= _zz_4155_;
      end
      if(_zz_4141_)begin
        int_reg_array_59_51_real <= _zz_4155_;
      end
      if(_zz_4142_)begin
        int_reg_array_59_52_real <= _zz_4155_;
      end
      if(_zz_4143_)begin
        int_reg_array_59_53_real <= _zz_4155_;
      end
      if(_zz_4144_)begin
        int_reg_array_59_54_real <= _zz_4155_;
      end
      if(_zz_4145_)begin
        int_reg_array_59_55_real <= _zz_4155_;
      end
      if(_zz_4146_)begin
        int_reg_array_59_56_real <= _zz_4155_;
      end
      if(_zz_4147_)begin
        int_reg_array_59_57_real <= _zz_4155_;
      end
      if(_zz_4148_)begin
        int_reg_array_59_58_real <= _zz_4155_;
      end
      if(_zz_4149_)begin
        int_reg_array_59_59_real <= _zz_4155_;
      end
      if(_zz_4150_)begin
        int_reg_array_59_60_real <= _zz_4155_;
      end
      if(_zz_4151_)begin
        int_reg_array_59_61_real <= _zz_4155_;
      end
      if(_zz_4152_)begin
        int_reg_array_59_62_real <= _zz_4155_;
      end
      if(_zz_4153_)begin
        int_reg_array_59_63_real <= _zz_4155_;
      end
      if(_zz_4090_)begin
        int_reg_array_59_0_imag <= _zz_4156_;
      end
      if(_zz_4091_)begin
        int_reg_array_59_1_imag <= _zz_4156_;
      end
      if(_zz_4092_)begin
        int_reg_array_59_2_imag <= _zz_4156_;
      end
      if(_zz_4093_)begin
        int_reg_array_59_3_imag <= _zz_4156_;
      end
      if(_zz_4094_)begin
        int_reg_array_59_4_imag <= _zz_4156_;
      end
      if(_zz_4095_)begin
        int_reg_array_59_5_imag <= _zz_4156_;
      end
      if(_zz_4096_)begin
        int_reg_array_59_6_imag <= _zz_4156_;
      end
      if(_zz_4097_)begin
        int_reg_array_59_7_imag <= _zz_4156_;
      end
      if(_zz_4098_)begin
        int_reg_array_59_8_imag <= _zz_4156_;
      end
      if(_zz_4099_)begin
        int_reg_array_59_9_imag <= _zz_4156_;
      end
      if(_zz_4100_)begin
        int_reg_array_59_10_imag <= _zz_4156_;
      end
      if(_zz_4101_)begin
        int_reg_array_59_11_imag <= _zz_4156_;
      end
      if(_zz_4102_)begin
        int_reg_array_59_12_imag <= _zz_4156_;
      end
      if(_zz_4103_)begin
        int_reg_array_59_13_imag <= _zz_4156_;
      end
      if(_zz_4104_)begin
        int_reg_array_59_14_imag <= _zz_4156_;
      end
      if(_zz_4105_)begin
        int_reg_array_59_15_imag <= _zz_4156_;
      end
      if(_zz_4106_)begin
        int_reg_array_59_16_imag <= _zz_4156_;
      end
      if(_zz_4107_)begin
        int_reg_array_59_17_imag <= _zz_4156_;
      end
      if(_zz_4108_)begin
        int_reg_array_59_18_imag <= _zz_4156_;
      end
      if(_zz_4109_)begin
        int_reg_array_59_19_imag <= _zz_4156_;
      end
      if(_zz_4110_)begin
        int_reg_array_59_20_imag <= _zz_4156_;
      end
      if(_zz_4111_)begin
        int_reg_array_59_21_imag <= _zz_4156_;
      end
      if(_zz_4112_)begin
        int_reg_array_59_22_imag <= _zz_4156_;
      end
      if(_zz_4113_)begin
        int_reg_array_59_23_imag <= _zz_4156_;
      end
      if(_zz_4114_)begin
        int_reg_array_59_24_imag <= _zz_4156_;
      end
      if(_zz_4115_)begin
        int_reg_array_59_25_imag <= _zz_4156_;
      end
      if(_zz_4116_)begin
        int_reg_array_59_26_imag <= _zz_4156_;
      end
      if(_zz_4117_)begin
        int_reg_array_59_27_imag <= _zz_4156_;
      end
      if(_zz_4118_)begin
        int_reg_array_59_28_imag <= _zz_4156_;
      end
      if(_zz_4119_)begin
        int_reg_array_59_29_imag <= _zz_4156_;
      end
      if(_zz_4120_)begin
        int_reg_array_59_30_imag <= _zz_4156_;
      end
      if(_zz_4121_)begin
        int_reg_array_59_31_imag <= _zz_4156_;
      end
      if(_zz_4122_)begin
        int_reg_array_59_32_imag <= _zz_4156_;
      end
      if(_zz_4123_)begin
        int_reg_array_59_33_imag <= _zz_4156_;
      end
      if(_zz_4124_)begin
        int_reg_array_59_34_imag <= _zz_4156_;
      end
      if(_zz_4125_)begin
        int_reg_array_59_35_imag <= _zz_4156_;
      end
      if(_zz_4126_)begin
        int_reg_array_59_36_imag <= _zz_4156_;
      end
      if(_zz_4127_)begin
        int_reg_array_59_37_imag <= _zz_4156_;
      end
      if(_zz_4128_)begin
        int_reg_array_59_38_imag <= _zz_4156_;
      end
      if(_zz_4129_)begin
        int_reg_array_59_39_imag <= _zz_4156_;
      end
      if(_zz_4130_)begin
        int_reg_array_59_40_imag <= _zz_4156_;
      end
      if(_zz_4131_)begin
        int_reg_array_59_41_imag <= _zz_4156_;
      end
      if(_zz_4132_)begin
        int_reg_array_59_42_imag <= _zz_4156_;
      end
      if(_zz_4133_)begin
        int_reg_array_59_43_imag <= _zz_4156_;
      end
      if(_zz_4134_)begin
        int_reg_array_59_44_imag <= _zz_4156_;
      end
      if(_zz_4135_)begin
        int_reg_array_59_45_imag <= _zz_4156_;
      end
      if(_zz_4136_)begin
        int_reg_array_59_46_imag <= _zz_4156_;
      end
      if(_zz_4137_)begin
        int_reg_array_59_47_imag <= _zz_4156_;
      end
      if(_zz_4138_)begin
        int_reg_array_59_48_imag <= _zz_4156_;
      end
      if(_zz_4139_)begin
        int_reg_array_59_49_imag <= _zz_4156_;
      end
      if(_zz_4140_)begin
        int_reg_array_59_50_imag <= _zz_4156_;
      end
      if(_zz_4141_)begin
        int_reg_array_59_51_imag <= _zz_4156_;
      end
      if(_zz_4142_)begin
        int_reg_array_59_52_imag <= _zz_4156_;
      end
      if(_zz_4143_)begin
        int_reg_array_59_53_imag <= _zz_4156_;
      end
      if(_zz_4144_)begin
        int_reg_array_59_54_imag <= _zz_4156_;
      end
      if(_zz_4145_)begin
        int_reg_array_59_55_imag <= _zz_4156_;
      end
      if(_zz_4146_)begin
        int_reg_array_59_56_imag <= _zz_4156_;
      end
      if(_zz_4147_)begin
        int_reg_array_59_57_imag <= _zz_4156_;
      end
      if(_zz_4148_)begin
        int_reg_array_59_58_imag <= _zz_4156_;
      end
      if(_zz_4149_)begin
        int_reg_array_59_59_imag <= _zz_4156_;
      end
      if(_zz_4150_)begin
        int_reg_array_59_60_imag <= _zz_4156_;
      end
      if(_zz_4151_)begin
        int_reg_array_59_61_imag <= _zz_4156_;
      end
      if(_zz_4152_)begin
        int_reg_array_59_62_imag <= _zz_4156_;
      end
      if(_zz_4153_)begin
        int_reg_array_59_63_imag <= _zz_4156_;
      end
      if(_zz_4159_)begin
        int_reg_array_60_0_real <= _zz_4224_;
      end
      if(_zz_4160_)begin
        int_reg_array_60_1_real <= _zz_4224_;
      end
      if(_zz_4161_)begin
        int_reg_array_60_2_real <= _zz_4224_;
      end
      if(_zz_4162_)begin
        int_reg_array_60_3_real <= _zz_4224_;
      end
      if(_zz_4163_)begin
        int_reg_array_60_4_real <= _zz_4224_;
      end
      if(_zz_4164_)begin
        int_reg_array_60_5_real <= _zz_4224_;
      end
      if(_zz_4165_)begin
        int_reg_array_60_6_real <= _zz_4224_;
      end
      if(_zz_4166_)begin
        int_reg_array_60_7_real <= _zz_4224_;
      end
      if(_zz_4167_)begin
        int_reg_array_60_8_real <= _zz_4224_;
      end
      if(_zz_4168_)begin
        int_reg_array_60_9_real <= _zz_4224_;
      end
      if(_zz_4169_)begin
        int_reg_array_60_10_real <= _zz_4224_;
      end
      if(_zz_4170_)begin
        int_reg_array_60_11_real <= _zz_4224_;
      end
      if(_zz_4171_)begin
        int_reg_array_60_12_real <= _zz_4224_;
      end
      if(_zz_4172_)begin
        int_reg_array_60_13_real <= _zz_4224_;
      end
      if(_zz_4173_)begin
        int_reg_array_60_14_real <= _zz_4224_;
      end
      if(_zz_4174_)begin
        int_reg_array_60_15_real <= _zz_4224_;
      end
      if(_zz_4175_)begin
        int_reg_array_60_16_real <= _zz_4224_;
      end
      if(_zz_4176_)begin
        int_reg_array_60_17_real <= _zz_4224_;
      end
      if(_zz_4177_)begin
        int_reg_array_60_18_real <= _zz_4224_;
      end
      if(_zz_4178_)begin
        int_reg_array_60_19_real <= _zz_4224_;
      end
      if(_zz_4179_)begin
        int_reg_array_60_20_real <= _zz_4224_;
      end
      if(_zz_4180_)begin
        int_reg_array_60_21_real <= _zz_4224_;
      end
      if(_zz_4181_)begin
        int_reg_array_60_22_real <= _zz_4224_;
      end
      if(_zz_4182_)begin
        int_reg_array_60_23_real <= _zz_4224_;
      end
      if(_zz_4183_)begin
        int_reg_array_60_24_real <= _zz_4224_;
      end
      if(_zz_4184_)begin
        int_reg_array_60_25_real <= _zz_4224_;
      end
      if(_zz_4185_)begin
        int_reg_array_60_26_real <= _zz_4224_;
      end
      if(_zz_4186_)begin
        int_reg_array_60_27_real <= _zz_4224_;
      end
      if(_zz_4187_)begin
        int_reg_array_60_28_real <= _zz_4224_;
      end
      if(_zz_4188_)begin
        int_reg_array_60_29_real <= _zz_4224_;
      end
      if(_zz_4189_)begin
        int_reg_array_60_30_real <= _zz_4224_;
      end
      if(_zz_4190_)begin
        int_reg_array_60_31_real <= _zz_4224_;
      end
      if(_zz_4191_)begin
        int_reg_array_60_32_real <= _zz_4224_;
      end
      if(_zz_4192_)begin
        int_reg_array_60_33_real <= _zz_4224_;
      end
      if(_zz_4193_)begin
        int_reg_array_60_34_real <= _zz_4224_;
      end
      if(_zz_4194_)begin
        int_reg_array_60_35_real <= _zz_4224_;
      end
      if(_zz_4195_)begin
        int_reg_array_60_36_real <= _zz_4224_;
      end
      if(_zz_4196_)begin
        int_reg_array_60_37_real <= _zz_4224_;
      end
      if(_zz_4197_)begin
        int_reg_array_60_38_real <= _zz_4224_;
      end
      if(_zz_4198_)begin
        int_reg_array_60_39_real <= _zz_4224_;
      end
      if(_zz_4199_)begin
        int_reg_array_60_40_real <= _zz_4224_;
      end
      if(_zz_4200_)begin
        int_reg_array_60_41_real <= _zz_4224_;
      end
      if(_zz_4201_)begin
        int_reg_array_60_42_real <= _zz_4224_;
      end
      if(_zz_4202_)begin
        int_reg_array_60_43_real <= _zz_4224_;
      end
      if(_zz_4203_)begin
        int_reg_array_60_44_real <= _zz_4224_;
      end
      if(_zz_4204_)begin
        int_reg_array_60_45_real <= _zz_4224_;
      end
      if(_zz_4205_)begin
        int_reg_array_60_46_real <= _zz_4224_;
      end
      if(_zz_4206_)begin
        int_reg_array_60_47_real <= _zz_4224_;
      end
      if(_zz_4207_)begin
        int_reg_array_60_48_real <= _zz_4224_;
      end
      if(_zz_4208_)begin
        int_reg_array_60_49_real <= _zz_4224_;
      end
      if(_zz_4209_)begin
        int_reg_array_60_50_real <= _zz_4224_;
      end
      if(_zz_4210_)begin
        int_reg_array_60_51_real <= _zz_4224_;
      end
      if(_zz_4211_)begin
        int_reg_array_60_52_real <= _zz_4224_;
      end
      if(_zz_4212_)begin
        int_reg_array_60_53_real <= _zz_4224_;
      end
      if(_zz_4213_)begin
        int_reg_array_60_54_real <= _zz_4224_;
      end
      if(_zz_4214_)begin
        int_reg_array_60_55_real <= _zz_4224_;
      end
      if(_zz_4215_)begin
        int_reg_array_60_56_real <= _zz_4224_;
      end
      if(_zz_4216_)begin
        int_reg_array_60_57_real <= _zz_4224_;
      end
      if(_zz_4217_)begin
        int_reg_array_60_58_real <= _zz_4224_;
      end
      if(_zz_4218_)begin
        int_reg_array_60_59_real <= _zz_4224_;
      end
      if(_zz_4219_)begin
        int_reg_array_60_60_real <= _zz_4224_;
      end
      if(_zz_4220_)begin
        int_reg_array_60_61_real <= _zz_4224_;
      end
      if(_zz_4221_)begin
        int_reg_array_60_62_real <= _zz_4224_;
      end
      if(_zz_4222_)begin
        int_reg_array_60_63_real <= _zz_4224_;
      end
      if(_zz_4159_)begin
        int_reg_array_60_0_imag <= _zz_4225_;
      end
      if(_zz_4160_)begin
        int_reg_array_60_1_imag <= _zz_4225_;
      end
      if(_zz_4161_)begin
        int_reg_array_60_2_imag <= _zz_4225_;
      end
      if(_zz_4162_)begin
        int_reg_array_60_3_imag <= _zz_4225_;
      end
      if(_zz_4163_)begin
        int_reg_array_60_4_imag <= _zz_4225_;
      end
      if(_zz_4164_)begin
        int_reg_array_60_5_imag <= _zz_4225_;
      end
      if(_zz_4165_)begin
        int_reg_array_60_6_imag <= _zz_4225_;
      end
      if(_zz_4166_)begin
        int_reg_array_60_7_imag <= _zz_4225_;
      end
      if(_zz_4167_)begin
        int_reg_array_60_8_imag <= _zz_4225_;
      end
      if(_zz_4168_)begin
        int_reg_array_60_9_imag <= _zz_4225_;
      end
      if(_zz_4169_)begin
        int_reg_array_60_10_imag <= _zz_4225_;
      end
      if(_zz_4170_)begin
        int_reg_array_60_11_imag <= _zz_4225_;
      end
      if(_zz_4171_)begin
        int_reg_array_60_12_imag <= _zz_4225_;
      end
      if(_zz_4172_)begin
        int_reg_array_60_13_imag <= _zz_4225_;
      end
      if(_zz_4173_)begin
        int_reg_array_60_14_imag <= _zz_4225_;
      end
      if(_zz_4174_)begin
        int_reg_array_60_15_imag <= _zz_4225_;
      end
      if(_zz_4175_)begin
        int_reg_array_60_16_imag <= _zz_4225_;
      end
      if(_zz_4176_)begin
        int_reg_array_60_17_imag <= _zz_4225_;
      end
      if(_zz_4177_)begin
        int_reg_array_60_18_imag <= _zz_4225_;
      end
      if(_zz_4178_)begin
        int_reg_array_60_19_imag <= _zz_4225_;
      end
      if(_zz_4179_)begin
        int_reg_array_60_20_imag <= _zz_4225_;
      end
      if(_zz_4180_)begin
        int_reg_array_60_21_imag <= _zz_4225_;
      end
      if(_zz_4181_)begin
        int_reg_array_60_22_imag <= _zz_4225_;
      end
      if(_zz_4182_)begin
        int_reg_array_60_23_imag <= _zz_4225_;
      end
      if(_zz_4183_)begin
        int_reg_array_60_24_imag <= _zz_4225_;
      end
      if(_zz_4184_)begin
        int_reg_array_60_25_imag <= _zz_4225_;
      end
      if(_zz_4185_)begin
        int_reg_array_60_26_imag <= _zz_4225_;
      end
      if(_zz_4186_)begin
        int_reg_array_60_27_imag <= _zz_4225_;
      end
      if(_zz_4187_)begin
        int_reg_array_60_28_imag <= _zz_4225_;
      end
      if(_zz_4188_)begin
        int_reg_array_60_29_imag <= _zz_4225_;
      end
      if(_zz_4189_)begin
        int_reg_array_60_30_imag <= _zz_4225_;
      end
      if(_zz_4190_)begin
        int_reg_array_60_31_imag <= _zz_4225_;
      end
      if(_zz_4191_)begin
        int_reg_array_60_32_imag <= _zz_4225_;
      end
      if(_zz_4192_)begin
        int_reg_array_60_33_imag <= _zz_4225_;
      end
      if(_zz_4193_)begin
        int_reg_array_60_34_imag <= _zz_4225_;
      end
      if(_zz_4194_)begin
        int_reg_array_60_35_imag <= _zz_4225_;
      end
      if(_zz_4195_)begin
        int_reg_array_60_36_imag <= _zz_4225_;
      end
      if(_zz_4196_)begin
        int_reg_array_60_37_imag <= _zz_4225_;
      end
      if(_zz_4197_)begin
        int_reg_array_60_38_imag <= _zz_4225_;
      end
      if(_zz_4198_)begin
        int_reg_array_60_39_imag <= _zz_4225_;
      end
      if(_zz_4199_)begin
        int_reg_array_60_40_imag <= _zz_4225_;
      end
      if(_zz_4200_)begin
        int_reg_array_60_41_imag <= _zz_4225_;
      end
      if(_zz_4201_)begin
        int_reg_array_60_42_imag <= _zz_4225_;
      end
      if(_zz_4202_)begin
        int_reg_array_60_43_imag <= _zz_4225_;
      end
      if(_zz_4203_)begin
        int_reg_array_60_44_imag <= _zz_4225_;
      end
      if(_zz_4204_)begin
        int_reg_array_60_45_imag <= _zz_4225_;
      end
      if(_zz_4205_)begin
        int_reg_array_60_46_imag <= _zz_4225_;
      end
      if(_zz_4206_)begin
        int_reg_array_60_47_imag <= _zz_4225_;
      end
      if(_zz_4207_)begin
        int_reg_array_60_48_imag <= _zz_4225_;
      end
      if(_zz_4208_)begin
        int_reg_array_60_49_imag <= _zz_4225_;
      end
      if(_zz_4209_)begin
        int_reg_array_60_50_imag <= _zz_4225_;
      end
      if(_zz_4210_)begin
        int_reg_array_60_51_imag <= _zz_4225_;
      end
      if(_zz_4211_)begin
        int_reg_array_60_52_imag <= _zz_4225_;
      end
      if(_zz_4212_)begin
        int_reg_array_60_53_imag <= _zz_4225_;
      end
      if(_zz_4213_)begin
        int_reg_array_60_54_imag <= _zz_4225_;
      end
      if(_zz_4214_)begin
        int_reg_array_60_55_imag <= _zz_4225_;
      end
      if(_zz_4215_)begin
        int_reg_array_60_56_imag <= _zz_4225_;
      end
      if(_zz_4216_)begin
        int_reg_array_60_57_imag <= _zz_4225_;
      end
      if(_zz_4217_)begin
        int_reg_array_60_58_imag <= _zz_4225_;
      end
      if(_zz_4218_)begin
        int_reg_array_60_59_imag <= _zz_4225_;
      end
      if(_zz_4219_)begin
        int_reg_array_60_60_imag <= _zz_4225_;
      end
      if(_zz_4220_)begin
        int_reg_array_60_61_imag <= _zz_4225_;
      end
      if(_zz_4221_)begin
        int_reg_array_60_62_imag <= _zz_4225_;
      end
      if(_zz_4222_)begin
        int_reg_array_60_63_imag <= _zz_4225_;
      end
      if(_zz_4228_)begin
        int_reg_array_61_0_real <= _zz_4293_;
      end
      if(_zz_4229_)begin
        int_reg_array_61_1_real <= _zz_4293_;
      end
      if(_zz_4230_)begin
        int_reg_array_61_2_real <= _zz_4293_;
      end
      if(_zz_4231_)begin
        int_reg_array_61_3_real <= _zz_4293_;
      end
      if(_zz_4232_)begin
        int_reg_array_61_4_real <= _zz_4293_;
      end
      if(_zz_4233_)begin
        int_reg_array_61_5_real <= _zz_4293_;
      end
      if(_zz_4234_)begin
        int_reg_array_61_6_real <= _zz_4293_;
      end
      if(_zz_4235_)begin
        int_reg_array_61_7_real <= _zz_4293_;
      end
      if(_zz_4236_)begin
        int_reg_array_61_8_real <= _zz_4293_;
      end
      if(_zz_4237_)begin
        int_reg_array_61_9_real <= _zz_4293_;
      end
      if(_zz_4238_)begin
        int_reg_array_61_10_real <= _zz_4293_;
      end
      if(_zz_4239_)begin
        int_reg_array_61_11_real <= _zz_4293_;
      end
      if(_zz_4240_)begin
        int_reg_array_61_12_real <= _zz_4293_;
      end
      if(_zz_4241_)begin
        int_reg_array_61_13_real <= _zz_4293_;
      end
      if(_zz_4242_)begin
        int_reg_array_61_14_real <= _zz_4293_;
      end
      if(_zz_4243_)begin
        int_reg_array_61_15_real <= _zz_4293_;
      end
      if(_zz_4244_)begin
        int_reg_array_61_16_real <= _zz_4293_;
      end
      if(_zz_4245_)begin
        int_reg_array_61_17_real <= _zz_4293_;
      end
      if(_zz_4246_)begin
        int_reg_array_61_18_real <= _zz_4293_;
      end
      if(_zz_4247_)begin
        int_reg_array_61_19_real <= _zz_4293_;
      end
      if(_zz_4248_)begin
        int_reg_array_61_20_real <= _zz_4293_;
      end
      if(_zz_4249_)begin
        int_reg_array_61_21_real <= _zz_4293_;
      end
      if(_zz_4250_)begin
        int_reg_array_61_22_real <= _zz_4293_;
      end
      if(_zz_4251_)begin
        int_reg_array_61_23_real <= _zz_4293_;
      end
      if(_zz_4252_)begin
        int_reg_array_61_24_real <= _zz_4293_;
      end
      if(_zz_4253_)begin
        int_reg_array_61_25_real <= _zz_4293_;
      end
      if(_zz_4254_)begin
        int_reg_array_61_26_real <= _zz_4293_;
      end
      if(_zz_4255_)begin
        int_reg_array_61_27_real <= _zz_4293_;
      end
      if(_zz_4256_)begin
        int_reg_array_61_28_real <= _zz_4293_;
      end
      if(_zz_4257_)begin
        int_reg_array_61_29_real <= _zz_4293_;
      end
      if(_zz_4258_)begin
        int_reg_array_61_30_real <= _zz_4293_;
      end
      if(_zz_4259_)begin
        int_reg_array_61_31_real <= _zz_4293_;
      end
      if(_zz_4260_)begin
        int_reg_array_61_32_real <= _zz_4293_;
      end
      if(_zz_4261_)begin
        int_reg_array_61_33_real <= _zz_4293_;
      end
      if(_zz_4262_)begin
        int_reg_array_61_34_real <= _zz_4293_;
      end
      if(_zz_4263_)begin
        int_reg_array_61_35_real <= _zz_4293_;
      end
      if(_zz_4264_)begin
        int_reg_array_61_36_real <= _zz_4293_;
      end
      if(_zz_4265_)begin
        int_reg_array_61_37_real <= _zz_4293_;
      end
      if(_zz_4266_)begin
        int_reg_array_61_38_real <= _zz_4293_;
      end
      if(_zz_4267_)begin
        int_reg_array_61_39_real <= _zz_4293_;
      end
      if(_zz_4268_)begin
        int_reg_array_61_40_real <= _zz_4293_;
      end
      if(_zz_4269_)begin
        int_reg_array_61_41_real <= _zz_4293_;
      end
      if(_zz_4270_)begin
        int_reg_array_61_42_real <= _zz_4293_;
      end
      if(_zz_4271_)begin
        int_reg_array_61_43_real <= _zz_4293_;
      end
      if(_zz_4272_)begin
        int_reg_array_61_44_real <= _zz_4293_;
      end
      if(_zz_4273_)begin
        int_reg_array_61_45_real <= _zz_4293_;
      end
      if(_zz_4274_)begin
        int_reg_array_61_46_real <= _zz_4293_;
      end
      if(_zz_4275_)begin
        int_reg_array_61_47_real <= _zz_4293_;
      end
      if(_zz_4276_)begin
        int_reg_array_61_48_real <= _zz_4293_;
      end
      if(_zz_4277_)begin
        int_reg_array_61_49_real <= _zz_4293_;
      end
      if(_zz_4278_)begin
        int_reg_array_61_50_real <= _zz_4293_;
      end
      if(_zz_4279_)begin
        int_reg_array_61_51_real <= _zz_4293_;
      end
      if(_zz_4280_)begin
        int_reg_array_61_52_real <= _zz_4293_;
      end
      if(_zz_4281_)begin
        int_reg_array_61_53_real <= _zz_4293_;
      end
      if(_zz_4282_)begin
        int_reg_array_61_54_real <= _zz_4293_;
      end
      if(_zz_4283_)begin
        int_reg_array_61_55_real <= _zz_4293_;
      end
      if(_zz_4284_)begin
        int_reg_array_61_56_real <= _zz_4293_;
      end
      if(_zz_4285_)begin
        int_reg_array_61_57_real <= _zz_4293_;
      end
      if(_zz_4286_)begin
        int_reg_array_61_58_real <= _zz_4293_;
      end
      if(_zz_4287_)begin
        int_reg_array_61_59_real <= _zz_4293_;
      end
      if(_zz_4288_)begin
        int_reg_array_61_60_real <= _zz_4293_;
      end
      if(_zz_4289_)begin
        int_reg_array_61_61_real <= _zz_4293_;
      end
      if(_zz_4290_)begin
        int_reg_array_61_62_real <= _zz_4293_;
      end
      if(_zz_4291_)begin
        int_reg_array_61_63_real <= _zz_4293_;
      end
      if(_zz_4228_)begin
        int_reg_array_61_0_imag <= _zz_4294_;
      end
      if(_zz_4229_)begin
        int_reg_array_61_1_imag <= _zz_4294_;
      end
      if(_zz_4230_)begin
        int_reg_array_61_2_imag <= _zz_4294_;
      end
      if(_zz_4231_)begin
        int_reg_array_61_3_imag <= _zz_4294_;
      end
      if(_zz_4232_)begin
        int_reg_array_61_4_imag <= _zz_4294_;
      end
      if(_zz_4233_)begin
        int_reg_array_61_5_imag <= _zz_4294_;
      end
      if(_zz_4234_)begin
        int_reg_array_61_6_imag <= _zz_4294_;
      end
      if(_zz_4235_)begin
        int_reg_array_61_7_imag <= _zz_4294_;
      end
      if(_zz_4236_)begin
        int_reg_array_61_8_imag <= _zz_4294_;
      end
      if(_zz_4237_)begin
        int_reg_array_61_9_imag <= _zz_4294_;
      end
      if(_zz_4238_)begin
        int_reg_array_61_10_imag <= _zz_4294_;
      end
      if(_zz_4239_)begin
        int_reg_array_61_11_imag <= _zz_4294_;
      end
      if(_zz_4240_)begin
        int_reg_array_61_12_imag <= _zz_4294_;
      end
      if(_zz_4241_)begin
        int_reg_array_61_13_imag <= _zz_4294_;
      end
      if(_zz_4242_)begin
        int_reg_array_61_14_imag <= _zz_4294_;
      end
      if(_zz_4243_)begin
        int_reg_array_61_15_imag <= _zz_4294_;
      end
      if(_zz_4244_)begin
        int_reg_array_61_16_imag <= _zz_4294_;
      end
      if(_zz_4245_)begin
        int_reg_array_61_17_imag <= _zz_4294_;
      end
      if(_zz_4246_)begin
        int_reg_array_61_18_imag <= _zz_4294_;
      end
      if(_zz_4247_)begin
        int_reg_array_61_19_imag <= _zz_4294_;
      end
      if(_zz_4248_)begin
        int_reg_array_61_20_imag <= _zz_4294_;
      end
      if(_zz_4249_)begin
        int_reg_array_61_21_imag <= _zz_4294_;
      end
      if(_zz_4250_)begin
        int_reg_array_61_22_imag <= _zz_4294_;
      end
      if(_zz_4251_)begin
        int_reg_array_61_23_imag <= _zz_4294_;
      end
      if(_zz_4252_)begin
        int_reg_array_61_24_imag <= _zz_4294_;
      end
      if(_zz_4253_)begin
        int_reg_array_61_25_imag <= _zz_4294_;
      end
      if(_zz_4254_)begin
        int_reg_array_61_26_imag <= _zz_4294_;
      end
      if(_zz_4255_)begin
        int_reg_array_61_27_imag <= _zz_4294_;
      end
      if(_zz_4256_)begin
        int_reg_array_61_28_imag <= _zz_4294_;
      end
      if(_zz_4257_)begin
        int_reg_array_61_29_imag <= _zz_4294_;
      end
      if(_zz_4258_)begin
        int_reg_array_61_30_imag <= _zz_4294_;
      end
      if(_zz_4259_)begin
        int_reg_array_61_31_imag <= _zz_4294_;
      end
      if(_zz_4260_)begin
        int_reg_array_61_32_imag <= _zz_4294_;
      end
      if(_zz_4261_)begin
        int_reg_array_61_33_imag <= _zz_4294_;
      end
      if(_zz_4262_)begin
        int_reg_array_61_34_imag <= _zz_4294_;
      end
      if(_zz_4263_)begin
        int_reg_array_61_35_imag <= _zz_4294_;
      end
      if(_zz_4264_)begin
        int_reg_array_61_36_imag <= _zz_4294_;
      end
      if(_zz_4265_)begin
        int_reg_array_61_37_imag <= _zz_4294_;
      end
      if(_zz_4266_)begin
        int_reg_array_61_38_imag <= _zz_4294_;
      end
      if(_zz_4267_)begin
        int_reg_array_61_39_imag <= _zz_4294_;
      end
      if(_zz_4268_)begin
        int_reg_array_61_40_imag <= _zz_4294_;
      end
      if(_zz_4269_)begin
        int_reg_array_61_41_imag <= _zz_4294_;
      end
      if(_zz_4270_)begin
        int_reg_array_61_42_imag <= _zz_4294_;
      end
      if(_zz_4271_)begin
        int_reg_array_61_43_imag <= _zz_4294_;
      end
      if(_zz_4272_)begin
        int_reg_array_61_44_imag <= _zz_4294_;
      end
      if(_zz_4273_)begin
        int_reg_array_61_45_imag <= _zz_4294_;
      end
      if(_zz_4274_)begin
        int_reg_array_61_46_imag <= _zz_4294_;
      end
      if(_zz_4275_)begin
        int_reg_array_61_47_imag <= _zz_4294_;
      end
      if(_zz_4276_)begin
        int_reg_array_61_48_imag <= _zz_4294_;
      end
      if(_zz_4277_)begin
        int_reg_array_61_49_imag <= _zz_4294_;
      end
      if(_zz_4278_)begin
        int_reg_array_61_50_imag <= _zz_4294_;
      end
      if(_zz_4279_)begin
        int_reg_array_61_51_imag <= _zz_4294_;
      end
      if(_zz_4280_)begin
        int_reg_array_61_52_imag <= _zz_4294_;
      end
      if(_zz_4281_)begin
        int_reg_array_61_53_imag <= _zz_4294_;
      end
      if(_zz_4282_)begin
        int_reg_array_61_54_imag <= _zz_4294_;
      end
      if(_zz_4283_)begin
        int_reg_array_61_55_imag <= _zz_4294_;
      end
      if(_zz_4284_)begin
        int_reg_array_61_56_imag <= _zz_4294_;
      end
      if(_zz_4285_)begin
        int_reg_array_61_57_imag <= _zz_4294_;
      end
      if(_zz_4286_)begin
        int_reg_array_61_58_imag <= _zz_4294_;
      end
      if(_zz_4287_)begin
        int_reg_array_61_59_imag <= _zz_4294_;
      end
      if(_zz_4288_)begin
        int_reg_array_61_60_imag <= _zz_4294_;
      end
      if(_zz_4289_)begin
        int_reg_array_61_61_imag <= _zz_4294_;
      end
      if(_zz_4290_)begin
        int_reg_array_61_62_imag <= _zz_4294_;
      end
      if(_zz_4291_)begin
        int_reg_array_61_63_imag <= _zz_4294_;
      end
      if(_zz_4297_)begin
        int_reg_array_62_0_real <= _zz_4362_;
      end
      if(_zz_4298_)begin
        int_reg_array_62_1_real <= _zz_4362_;
      end
      if(_zz_4299_)begin
        int_reg_array_62_2_real <= _zz_4362_;
      end
      if(_zz_4300_)begin
        int_reg_array_62_3_real <= _zz_4362_;
      end
      if(_zz_4301_)begin
        int_reg_array_62_4_real <= _zz_4362_;
      end
      if(_zz_4302_)begin
        int_reg_array_62_5_real <= _zz_4362_;
      end
      if(_zz_4303_)begin
        int_reg_array_62_6_real <= _zz_4362_;
      end
      if(_zz_4304_)begin
        int_reg_array_62_7_real <= _zz_4362_;
      end
      if(_zz_4305_)begin
        int_reg_array_62_8_real <= _zz_4362_;
      end
      if(_zz_4306_)begin
        int_reg_array_62_9_real <= _zz_4362_;
      end
      if(_zz_4307_)begin
        int_reg_array_62_10_real <= _zz_4362_;
      end
      if(_zz_4308_)begin
        int_reg_array_62_11_real <= _zz_4362_;
      end
      if(_zz_4309_)begin
        int_reg_array_62_12_real <= _zz_4362_;
      end
      if(_zz_4310_)begin
        int_reg_array_62_13_real <= _zz_4362_;
      end
      if(_zz_4311_)begin
        int_reg_array_62_14_real <= _zz_4362_;
      end
      if(_zz_4312_)begin
        int_reg_array_62_15_real <= _zz_4362_;
      end
      if(_zz_4313_)begin
        int_reg_array_62_16_real <= _zz_4362_;
      end
      if(_zz_4314_)begin
        int_reg_array_62_17_real <= _zz_4362_;
      end
      if(_zz_4315_)begin
        int_reg_array_62_18_real <= _zz_4362_;
      end
      if(_zz_4316_)begin
        int_reg_array_62_19_real <= _zz_4362_;
      end
      if(_zz_4317_)begin
        int_reg_array_62_20_real <= _zz_4362_;
      end
      if(_zz_4318_)begin
        int_reg_array_62_21_real <= _zz_4362_;
      end
      if(_zz_4319_)begin
        int_reg_array_62_22_real <= _zz_4362_;
      end
      if(_zz_4320_)begin
        int_reg_array_62_23_real <= _zz_4362_;
      end
      if(_zz_4321_)begin
        int_reg_array_62_24_real <= _zz_4362_;
      end
      if(_zz_4322_)begin
        int_reg_array_62_25_real <= _zz_4362_;
      end
      if(_zz_4323_)begin
        int_reg_array_62_26_real <= _zz_4362_;
      end
      if(_zz_4324_)begin
        int_reg_array_62_27_real <= _zz_4362_;
      end
      if(_zz_4325_)begin
        int_reg_array_62_28_real <= _zz_4362_;
      end
      if(_zz_4326_)begin
        int_reg_array_62_29_real <= _zz_4362_;
      end
      if(_zz_4327_)begin
        int_reg_array_62_30_real <= _zz_4362_;
      end
      if(_zz_4328_)begin
        int_reg_array_62_31_real <= _zz_4362_;
      end
      if(_zz_4329_)begin
        int_reg_array_62_32_real <= _zz_4362_;
      end
      if(_zz_4330_)begin
        int_reg_array_62_33_real <= _zz_4362_;
      end
      if(_zz_4331_)begin
        int_reg_array_62_34_real <= _zz_4362_;
      end
      if(_zz_4332_)begin
        int_reg_array_62_35_real <= _zz_4362_;
      end
      if(_zz_4333_)begin
        int_reg_array_62_36_real <= _zz_4362_;
      end
      if(_zz_4334_)begin
        int_reg_array_62_37_real <= _zz_4362_;
      end
      if(_zz_4335_)begin
        int_reg_array_62_38_real <= _zz_4362_;
      end
      if(_zz_4336_)begin
        int_reg_array_62_39_real <= _zz_4362_;
      end
      if(_zz_4337_)begin
        int_reg_array_62_40_real <= _zz_4362_;
      end
      if(_zz_4338_)begin
        int_reg_array_62_41_real <= _zz_4362_;
      end
      if(_zz_4339_)begin
        int_reg_array_62_42_real <= _zz_4362_;
      end
      if(_zz_4340_)begin
        int_reg_array_62_43_real <= _zz_4362_;
      end
      if(_zz_4341_)begin
        int_reg_array_62_44_real <= _zz_4362_;
      end
      if(_zz_4342_)begin
        int_reg_array_62_45_real <= _zz_4362_;
      end
      if(_zz_4343_)begin
        int_reg_array_62_46_real <= _zz_4362_;
      end
      if(_zz_4344_)begin
        int_reg_array_62_47_real <= _zz_4362_;
      end
      if(_zz_4345_)begin
        int_reg_array_62_48_real <= _zz_4362_;
      end
      if(_zz_4346_)begin
        int_reg_array_62_49_real <= _zz_4362_;
      end
      if(_zz_4347_)begin
        int_reg_array_62_50_real <= _zz_4362_;
      end
      if(_zz_4348_)begin
        int_reg_array_62_51_real <= _zz_4362_;
      end
      if(_zz_4349_)begin
        int_reg_array_62_52_real <= _zz_4362_;
      end
      if(_zz_4350_)begin
        int_reg_array_62_53_real <= _zz_4362_;
      end
      if(_zz_4351_)begin
        int_reg_array_62_54_real <= _zz_4362_;
      end
      if(_zz_4352_)begin
        int_reg_array_62_55_real <= _zz_4362_;
      end
      if(_zz_4353_)begin
        int_reg_array_62_56_real <= _zz_4362_;
      end
      if(_zz_4354_)begin
        int_reg_array_62_57_real <= _zz_4362_;
      end
      if(_zz_4355_)begin
        int_reg_array_62_58_real <= _zz_4362_;
      end
      if(_zz_4356_)begin
        int_reg_array_62_59_real <= _zz_4362_;
      end
      if(_zz_4357_)begin
        int_reg_array_62_60_real <= _zz_4362_;
      end
      if(_zz_4358_)begin
        int_reg_array_62_61_real <= _zz_4362_;
      end
      if(_zz_4359_)begin
        int_reg_array_62_62_real <= _zz_4362_;
      end
      if(_zz_4360_)begin
        int_reg_array_62_63_real <= _zz_4362_;
      end
      if(_zz_4297_)begin
        int_reg_array_62_0_imag <= _zz_4363_;
      end
      if(_zz_4298_)begin
        int_reg_array_62_1_imag <= _zz_4363_;
      end
      if(_zz_4299_)begin
        int_reg_array_62_2_imag <= _zz_4363_;
      end
      if(_zz_4300_)begin
        int_reg_array_62_3_imag <= _zz_4363_;
      end
      if(_zz_4301_)begin
        int_reg_array_62_4_imag <= _zz_4363_;
      end
      if(_zz_4302_)begin
        int_reg_array_62_5_imag <= _zz_4363_;
      end
      if(_zz_4303_)begin
        int_reg_array_62_6_imag <= _zz_4363_;
      end
      if(_zz_4304_)begin
        int_reg_array_62_7_imag <= _zz_4363_;
      end
      if(_zz_4305_)begin
        int_reg_array_62_8_imag <= _zz_4363_;
      end
      if(_zz_4306_)begin
        int_reg_array_62_9_imag <= _zz_4363_;
      end
      if(_zz_4307_)begin
        int_reg_array_62_10_imag <= _zz_4363_;
      end
      if(_zz_4308_)begin
        int_reg_array_62_11_imag <= _zz_4363_;
      end
      if(_zz_4309_)begin
        int_reg_array_62_12_imag <= _zz_4363_;
      end
      if(_zz_4310_)begin
        int_reg_array_62_13_imag <= _zz_4363_;
      end
      if(_zz_4311_)begin
        int_reg_array_62_14_imag <= _zz_4363_;
      end
      if(_zz_4312_)begin
        int_reg_array_62_15_imag <= _zz_4363_;
      end
      if(_zz_4313_)begin
        int_reg_array_62_16_imag <= _zz_4363_;
      end
      if(_zz_4314_)begin
        int_reg_array_62_17_imag <= _zz_4363_;
      end
      if(_zz_4315_)begin
        int_reg_array_62_18_imag <= _zz_4363_;
      end
      if(_zz_4316_)begin
        int_reg_array_62_19_imag <= _zz_4363_;
      end
      if(_zz_4317_)begin
        int_reg_array_62_20_imag <= _zz_4363_;
      end
      if(_zz_4318_)begin
        int_reg_array_62_21_imag <= _zz_4363_;
      end
      if(_zz_4319_)begin
        int_reg_array_62_22_imag <= _zz_4363_;
      end
      if(_zz_4320_)begin
        int_reg_array_62_23_imag <= _zz_4363_;
      end
      if(_zz_4321_)begin
        int_reg_array_62_24_imag <= _zz_4363_;
      end
      if(_zz_4322_)begin
        int_reg_array_62_25_imag <= _zz_4363_;
      end
      if(_zz_4323_)begin
        int_reg_array_62_26_imag <= _zz_4363_;
      end
      if(_zz_4324_)begin
        int_reg_array_62_27_imag <= _zz_4363_;
      end
      if(_zz_4325_)begin
        int_reg_array_62_28_imag <= _zz_4363_;
      end
      if(_zz_4326_)begin
        int_reg_array_62_29_imag <= _zz_4363_;
      end
      if(_zz_4327_)begin
        int_reg_array_62_30_imag <= _zz_4363_;
      end
      if(_zz_4328_)begin
        int_reg_array_62_31_imag <= _zz_4363_;
      end
      if(_zz_4329_)begin
        int_reg_array_62_32_imag <= _zz_4363_;
      end
      if(_zz_4330_)begin
        int_reg_array_62_33_imag <= _zz_4363_;
      end
      if(_zz_4331_)begin
        int_reg_array_62_34_imag <= _zz_4363_;
      end
      if(_zz_4332_)begin
        int_reg_array_62_35_imag <= _zz_4363_;
      end
      if(_zz_4333_)begin
        int_reg_array_62_36_imag <= _zz_4363_;
      end
      if(_zz_4334_)begin
        int_reg_array_62_37_imag <= _zz_4363_;
      end
      if(_zz_4335_)begin
        int_reg_array_62_38_imag <= _zz_4363_;
      end
      if(_zz_4336_)begin
        int_reg_array_62_39_imag <= _zz_4363_;
      end
      if(_zz_4337_)begin
        int_reg_array_62_40_imag <= _zz_4363_;
      end
      if(_zz_4338_)begin
        int_reg_array_62_41_imag <= _zz_4363_;
      end
      if(_zz_4339_)begin
        int_reg_array_62_42_imag <= _zz_4363_;
      end
      if(_zz_4340_)begin
        int_reg_array_62_43_imag <= _zz_4363_;
      end
      if(_zz_4341_)begin
        int_reg_array_62_44_imag <= _zz_4363_;
      end
      if(_zz_4342_)begin
        int_reg_array_62_45_imag <= _zz_4363_;
      end
      if(_zz_4343_)begin
        int_reg_array_62_46_imag <= _zz_4363_;
      end
      if(_zz_4344_)begin
        int_reg_array_62_47_imag <= _zz_4363_;
      end
      if(_zz_4345_)begin
        int_reg_array_62_48_imag <= _zz_4363_;
      end
      if(_zz_4346_)begin
        int_reg_array_62_49_imag <= _zz_4363_;
      end
      if(_zz_4347_)begin
        int_reg_array_62_50_imag <= _zz_4363_;
      end
      if(_zz_4348_)begin
        int_reg_array_62_51_imag <= _zz_4363_;
      end
      if(_zz_4349_)begin
        int_reg_array_62_52_imag <= _zz_4363_;
      end
      if(_zz_4350_)begin
        int_reg_array_62_53_imag <= _zz_4363_;
      end
      if(_zz_4351_)begin
        int_reg_array_62_54_imag <= _zz_4363_;
      end
      if(_zz_4352_)begin
        int_reg_array_62_55_imag <= _zz_4363_;
      end
      if(_zz_4353_)begin
        int_reg_array_62_56_imag <= _zz_4363_;
      end
      if(_zz_4354_)begin
        int_reg_array_62_57_imag <= _zz_4363_;
      end
      if(_zz_4355_)begin
        int_reg_array_62_58_imag <= _zz_4363_;
      end
      if(_zz_4356_)begin
        int_reg_array_62_59_imag <= _zz_4363_;
      end
      if(_zz_4357_)begin
        int_reg_array_62_60_imag <= _zz_4363_;
      end
      if(_zz_4358_)begin
        int_reg_array_62_61_imag <= _zz_4363_;
      end
      if(_zz_4359_)begin
        int_reg_array_62_62_imag <= _zz_4363_;
      end
      if(_zz_4360_)begin
        int_reg_array_62_63_imag <= _zz_4363_;
      end
      if(_zz_4366_)begin
        int_reg_array_63_0_real <= _zz_4431_;
      end
      if(_zz_4367_)begin
        int_reg_array_63_1_real <= _zz_4431_;
      end
      if(_zz_4368_)begin
        int_reg_array_63_2_real <= _zz_4431_;
      end
      if(_zz_4369_)begin
        int_reg_array_63_3_real <= _zz_4431_;
      end
      if(_zz_4370_)begin
        int_reg_array_63_4_real <= _zz_4431_;
      end
      if(_zz_4371_)begin
        int_reg_array_63_5_real <= _zz_4431_;
      end
      if(_zz_4372_)begin
        int_reg_array_63_6_real <= _zz_4431_;
      end
      if(_zz_4373_)begin
        int_reg_array_63_7_real <= _zz_4431_;
      end
      if(_zz_4374_)begin
        int_reg_array_63_8_real <= _zz_4431_;
      end
      if(_zz_4375_)begin
        int_reg_array_63_9_real <= _zz_4431_;
      end
      if(_zz_4376_)begin
        int_reg_array_63_10_real <= _zz_4431_;
      end
      if(_zz_4377_)begin
        int_reg_array_63_11_real <= _zz_4431_;
      end
      if(_zz_4378_)begin
        int_reg_array_63_12_real <= _zz_4431_;
      end
      if(_zz_4379_)begin
        int_reg_array_63_13_real <= _zz_4431_;
      end
      if(_zz_4380_)begin
        int_reg_array_63_14_real <= _zz_4431_;
      end
      if(_zz_4381_)begin
        int_reg_array_63_15_real <= _zz_4431_;
      end
      if(_zz_4382_)begin
        int_reg_array_63_16_real <= _zz_4431_;
      end
      if(_zz_4383_)begin
        int_reg_array_63_17_real <= _zz_4431_;
      end
      if(_zz_4384_)begin
        int_reg_array_63_18_real <= _zz_4431_;
      end
      if(_zz_4385_)begin
        int_reg_array_63_19_real <= _zz_4431_;
      end
      if(_zz_4386_)begin
        int_reg_array_63_20_real <= _zz_4431_;
      end
      if(_zz_4387_)begin
        int_reg_array_63_21_real <= _zz_4431_;
      end
      if(_zz_4388_)begin
        int_reg_array_63_22_real <= _zz_4431_;
      end
      if(_zz_4389_)begin
        int_reg_array_63_23_real <= _zz_4431_;
      end
      if(_zz_4390_)begin
        int_reg_array_63_24_real <= _zz_4431_;
      end
      if(_zz_4391_)begin
        int_reg_array_63_25_real <= _zz_4431_;
      end
      if(_zz_4392_)begin
        int_reg_array_63_26_real <= _zz_4431_;
      end
      if(_zz_4393_)begin
        int_reg_array_63_27_real <= _zz_4431_;
      end
      if(_zz_4394_)begin
        int_reg_array_63_28_real <= _zz_4431_;
      end
      if(_zz_4395_)begin
        int_reg_array_63_29_real <= _zz_4431_;
      end
      if(_zz_4396_)begin
        int_reg_array_63_30_real <= _zz_4431_;
      end
      if(_zz_4397_)begin
        int_reg_array_63_31_real <= _zz_4431_;
      end
      if(_zz_4398_)begin
        int_reg_array_63_32_real <= _zz_4431_;
      end
      if(_zz_4399_)begin
        int_reg_array_63_33_real <= _zz_4431_;
      end
      if(_zz_4400_)begin
        int_reg_array_63_34_real <= _zz_4431_;
      end
      if(_zz_4401_)begin
        int_reg_array_63_35_real <= _zz_4431_;
      end
      if(_zz_4402_)begin
        int_reg_array_63_36_real <= _zz_4431_;
      end
      if(_zz_4403_)begin
        int_reg_array_63_37_real <= _zz_4431_;
      end
      if(_zz_4404_)begin
        int_reg_array_63_38_real <= _zz_4431_;
      end
      if(_zz_4405_)begin
        int_reg_array_63_39_real <= _zz_4431_;
      end
      if(_zz_4406_)begin
        int_reg_array_63_40_real <= _zz_4431_;
      end
      if(_zz_4407_)begin
        int_reg_array_63_41_real <= _zz_4431_;
      end
      if(_zz_4408_)begin
        int_reg_array_63_42_real <= _zz_4431_;
      end
      if(_zz_4409_)begin
        int_reg_array_63_43_real <= _zz_4431_;
      end
      if(_zz_4410_)begin
        int_reg_array_63_44_real <= _zz_4431_;
      end
      if(_zz_4411_)begin
        int_reg_array_63_45_real <= _zz_4431_;
      end
      if(_zz_4412_)begin
        int_reg_array_63_46_real <= _zz_4431_;
      end
      if(_zz_4413_)begin
        int_reg_array_63_47_real <= _zz_4431_;
      end
      if(_zz_4414_)begin
        int_reg_array_63_48_real <= _zz_4431_;
      end
      if(_zz_4415_)begin
        int_reg_array_63_49_real <= _zz_4431_;
      end
      if(_zz_4416_)begin
        int_reg_array_63_50_real <= _zz_4431_;
      end
      if(_zz_4417_)begin
        int_reg_array_63_51_real <= _zz_4431_;
      end
      if(_zz_4418_)begin
        int_reg_array_63_52_real <= _zz_4431_;
      end
      if(_zz_4419_)begin
        int_reg_array_63_53_real <= _zz_4431_;
      end
      if(_zz_4420_)begin
        int_reg_array_63_54_real <= _zz_4431_;
      end
      if(_zz_4421_)begin
        int_reg_array_63_55_real <= _zz_4431_;
      end
      if(_zz_4422_)begin
        int_reg_array_63_56_real <= _zz_4431_;
      end
      if(_zz_4423_)begin
        int_reg_array_63_57_real <= _zz_4431_;
      end
      if(_zz_4424_)begin
        int_reg_array_63_58_real <= _zz_4431_;
      end
      if(_zz_4425_)begin
        int_reg_array_63_59_real <= _zz_4431_;
      end
      if(_zz_4426_)begin
        int_reg_array_63_60_real <= _zz_4431_;
      end
      if(_zz_4427_)begin
        int_reg_array_63_61_real <= _zz_4431_;
      end
      if(_zz_4428_)begin
        int_reg_array_63_62_real <= _zz_4431_;
      end
      if(_zz_4429_)begin
        int_reg_array_63_63_real <= _zz_4431_;
      end
      if(_zz_4366_)begin
        int_reg_array_63_0_imag <= _zz_4432_;
      end
      if(_zz_4367_)begin
        int_reg_array_63_1_imag <= _zz_4432_;
      end
      if(_zz_4368_)begin
        int_reg_array_63_2_imag <= _zz_4432_;
      end
      if(_zz_4369_)begin
        int_reg_array_63_3_imag <= _zz_4432_;
      end
      if(_zz_4370_)begin
        int_reg_array_63_4_imag <= _zz_4432_;
      end
      if(_zz_4371_)begin
        int_reg_array_63_5_imag <= _zz_4432_;
      end
      if(_zz_4372_)begin
        int_reg_array_63_6_imag <= _zz_4432_;
      end
      if(_zz_4373_)begin
        int_reg_array_63_7_imag <= _zz_4432_;
      end
      if(_zz_4374_)begin
        int_reg_array_63_8_imag <= _zz_4432_;
      end
      if(_zz_4375_)begin
        int_reg_array_63_9_imag <= _zz_4432_;
      end
      if(_zz_4376_)begin
        int_reg_array_63_10_imag <= _zz_4432_;
      end
      if(_zz_4377_)begin
        int_reg_array_63_11_imag <= _zz_4432_;
      end
      if(_zz_4378_)begin
        int_reg_array_63_12_imag <= _zz_4432_;
      end
      if(_zz_4379_)begin
        int_reg_array_63_13_imag <= _zz_4432_;
      end
      if(_zz_4380_)begin
        int_reg_array_63_14_imag <= _zz_4432_;
      end
      if(_zz_4381_)begin
        int_reg_array_63_15_imag <= _zz_4432_;
      end
      if(_zz_4382_)begin
        int_reg_array_63_16_imag <= _zz_4432_;
      end
      if(_zz_4383_)begin
        int_reg_array_63_17_imag <= _zz_4432_;
      end
      if(_zz_4384_)begin
        int_reg_array_63_18_imag <= _zz_4432_;
      end
      if(_zz_4385_)begin
        int_reg_array_63_19_imag <= _zz_4432_;
      end
      if(_zz_4386_)begin
        int_reg_array_63_20_imag <= _zz_4432_;
      end
      if(_zz_4387_)begin
        int_reg_array_63_21_imag <= _zz_4432_;
      end
      if(_zz_4388_)begin
        int_reg_array_63_22_imag <= _zz_4432_;
      end
      if(_zz_4389_)begin
        int_reg_array_63_23_imag <= _zz_4432_;
      end
      if(_zz_4390_)begin
        int_reg_array_63_24_imag <= _zz_4432_;
      end
      if(_zz_4391_)begin
        int_reg_array_63_25_imag <= _zz_4432_;
      end
      if(_zz_4392_)begin
        int_reg_array_63_26_imag <= _zz_4432_;
      end
      if(_zz_4393_)begin
        int_reg_array_63_27_imag <= _zz_4432_;
      end
      if(_zz_4394_)begin
        int_reg_array_63_28_imag <= _zz_4432_;
      end
      if(_zz_4395_)begin
        int_reg_array_63_29_imag <= _zz_4432_;
      end
      if(_zz_4396_)begin
        int_reg_array_63_30_imag <= _zz_4432_;
      end
      if(_zz_4397_)begin
        int_reg_array_63_31_imag <= _zz_4432_;
      end
      if(_zz_4398_)begin
        int_reg_array_63_32_imag <= _zz_4432_;
      end
      if(_zz_4399_)begin
        int_reg_array_63_33_imag <= _zz_4432_;
      end
      if(_zz_4400_)begin
        int_reg_array_63_34_imag <= _zz_4432_;
      end
      if(_zz_4401_)begin
        int_reg_array_63_35_imag <= _zz_4432_;
      end
      if(_zz_4402_)begin
        int_reg_array_63_36_imag <= _zz_4432_;
      end
      if(_zz_4403_)begin
        int_reg_array_63_37_imag <= _zz_4432_;
      end
      if(_zz_4404_)begin
        int_reg_array_63_38_imag <= _zz_4432_;
      end
      if(_zz_4405_)begin
        int_reg_array_63_39_imag <= _zz_4432_;
      end
      if(_zz_4406_)begin
        int_reg_array_63_40_imag <= _zz_4432_;
      end
      if(_zz_4407_)begin
        int_reg_array_63_41_imag <= _zz_4432_;
      end
      if(_zz_4408_)begin
        int_reg_array_63_42_imag <= _zz_4432_;
      end
      if(_zz_4409_)begin
        int_reg_array_63_43_imag <= _zz_4432_;
      end
      if(_zz_4410_)begin
        int_reg_array_63_44_imag <= _zz_4432_;
      end
      if(_zz_4411_)begin
        int_reg_array_63_45_imag <= _zz_4432_;
      end
      if(_zz_4412_)begin
        int_reg_array_63_46_imag <= _zz_4432_;
      end
      if(_zz_4413_)begin
        int_reg_array_63_47_imag <= _zz_4432_;
      end
      if(_zz_4414_)begin
        int_reg_array_63_48_imag <= _zz_4432_;
      end
      if(_zz_4415_)begin
        int_reg_array_63_49_imag <= _zz_4432_;
      end
      if(_zz_4416_)begin
        int_reg_array_63_50_imag <= _zz_4432_;
      end
      if(_zz_4417_)begin
        int_reg_array_63_51_imag <= _zz_4432_;
      end
      if(_zz_4418_)begin
        int_reg_array_63_52_imag <= _zz_4432_;
      end
      if(_zz_4419_)begin
        int_reg_array_63_53_imag <= _zz_4432_;
      end
      if(_zz_4420_)begin
        int_reg_array_63_54_imag <= _zz_4432_;
      end
      if(_zz_4421_)begin
        int_reg_array_63_55_imag <= _zz_4432_;
      end
      if(_zz_4422_)begin
        int_reg_array_63_56_imag <= _zz_4432_;
      end
      if(_zz_4423_)begin
        int_reg_array_63_57_imag <= _zz_4432_;
      end
      if(_zz_4424_)begin
        int_reg_array_63_58_imag <= _zz_4432_;
      end
      if(_zz_4425_)begin
        int_reg_array_63_59_imag <= _zz_4432_;
      end
      if(_zz_4426_)begin
        int_reg_array_63_60_imag <= _zz_4432_;
      end
      if(_zz_4427_)begin
        int_reg_array_63_61_imag <= _zz_4432_;
      end
      if(_zz_4428_)begin
        int_reg_array_63_62_imag <= _zz_4432_;
      end
      if(_zz_4429_)begin
        int_reg_array_63_63_imag <= _zz_4432_;
      end
    end
  end

  always @ (posedge clk or posedge reset) begin
    if (reset) begin
      load_data_area_current_addr <= 32'h0;
    end else begin
      if(_zz_7_)begin
        load_data_area_current_addr <= Axi4Incr_result;
      end
    end
  end

  always @ (posedge clk) begin
    _zz_9__regNext <= _zz_9_;
  end


endmodule
