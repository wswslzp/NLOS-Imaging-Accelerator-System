// Generator : SpinalHDL v1.4.1    git head : d1b4746673438bc5f242515335278fa39a666c38
// Component : SFFT
// Git hash  : 5b9162698fb44411d3965102ba2614672aab0931



module SFFT (
  input               data_in_valid,
  input      [15:0]   data_in_payload_real,
  input      [15:0]   data_in_payload_imag,
  output              data_out_valid,
  output     [15:0]   data_out_payload_real,
  output     [15:0]   data_out_payload_imag,
  input               clk,
  input               reset
);
  reg        [15:0]   _zz_257;
  reg        [15:0]   _zz_258;
  wire                myFFT_1_sdata_out_valid;
  wire       [15:0]   myFFT_1_sdata_out_payload_0_real;
  wire       [15:0]   myFFT_1_sdata_out_payload_0_imag;
  wire       [15:0]   myFFT_1_sdata_out_payload_1_real;
  wire       [15:0]   myFFT_1_sdata_out_payload_1_imag;
  wire       [15:0]   myFFT_1_sdata_out_payload_2_real;
  wire       [15:0]   myFFT_1_sdata_out_payload_2_imag;
  wire       [15:0]   myFFT_1_sdata_out_payload_3_real;
  wire       [15:0]   myFFT_1_sdata_out_payload_3_imag;
  wire       [15:0]   myFFT_1_sdata_out_payload_4_real;
  wire       [15:0]   myFFT_1_sdata_out_payload_4_imag;
  wire       [15:0]   myFFT_1_sdata_out_payload_5_real;
  wire       [15:0]   myFFT_1_sdata_out_payload_5_imag;
  wire       [15:0]   myFFT_1_sdata_out_payload_6_real;
  wire       [15:0]   myFFT_1_sdata_out_payload_6_imag;
  wire       [15:0]   myFFT_1_sdata_out_payload_7_real;
  wire       [15:0]   myFFT_1_sdata_out_payload_7_imag;
  wire       [15:0]   myFFT_1_sdata_out_payload_8_real;
  wire       [15:0]   myFFT_1_sdata_out_payload_8_imag;
  wire       [15:0]   myFFT_1_sdata_out_payload_9_real;
  wire       [15:0]   myFFT_1_sdata_out_payload_9_imag;
  wire       [15:0]   myFFT_1_sdata_out_payload_10_real;
  wire       [15:0]   myFFT_1_sdata_out_payload_10_imag;
  wire       [15:0]   myFFT_1_sdata_out_payload_11_real;
  wire       [15:0]   myFFT_1_sdata_out_payload_11_imag;
  wire       [15:0]   myFFT_1_sdata_out_payload_12_real;
  wire       [15:0]   myFFT_1_sdata_out_payload_12_imag;
  wire       [15:0]   myFFT_1_sdata_out_payload_13_real;
  wire       [15:0]   myFFT_1_sdata_out_payload_13_imag;
  wire       [15:0]   myFFT_1_sdata_out_payload_14_real;
  wire       [15:0]   myFFT_1_sdata_out_payload_14_imag;
  wire       [15:0]   myFFT_1_sdata_out_payload_15_real;
  wire       [15:0]   myFFT_1_sdata_out_payload_15_imag;
  wire       [15:0]   myFFT_1_sdata_out_payload_16_real;
  wire       [15:0]   myFFT_1_sdata_out_payload_16_imag;
  wire       [15:0]   myFFT_1_sdata_out_payload_17_real;
  wire       [15:0]   myFFT_1_sdata_out_payload_17_imag;
  wire       [15:0]   myFFT_1_sdata_out_payload_18_real;
  wire       [15:0]   myFFT_1_sdata_out_payload_18_imag;
  wire       [15:0]   myFFT_1_sdata_out_payload_19_real;
  wire       [15:0]   myFFT_1_sdata_out_payload_19_imag;
  wire       [15:0]   myFFT_1_sdata_out_payload_20_real;
  wire       [15:0]   myFFT_1_sdata_out_payload_20_imag;
  wire       [15:0]   myFFT_1_sdata_out_payload_21_real;
  wire       [15:0]   myFFT_1_sdata_out_payload_21_imag;
  wire       [15:0]   myFFT_1_sdata_out_payload_22_real;
  wire       [15:0]   myFFT_1_sdata_out_payload_22_imag;
  wire       [15:0]   myFFT_1_sdata_out_payload_23_real;
  wire       [15:0]   myFFT_1_sdata_out_payload_23_imag;
  wire       [15:0]   myFFT_1_sdata_out_payload_24_real;
  wire       [15:0]   myFFT_1_sdata_out_payload_24_imag;
  wire       [15:0]   myFFT_1_sdata_out_payload_25_real;
  wire       [15:0]   myFFT_1_sdata_out_payload_25_imag;
  wire       [15:0]   myFFT_1_sdata_out_payload_26_real;
  wire       [15:0]   myFFT_1_sdata_out_payload_26_imag;
  wire       [15:0]   myFFT_1_sdata_out_payload_27_real;
  wire       [15:0]   myFFT_1_sdata_out_payload_27_imag;
  wire       [15:0]   myFFT_1_sdata_out_payload_28_real;
  wire       [15:0]   myFFT_1_sdata_out_payload_28_imag;
  wire       [15:0]   myFFT_1_sdata_out_payload_29_real;
  wire       [15:0]   myFFT_1_sdata_out_payload_29_imag;
  wire       [15:0]   myFFT_1_sdata_out_payload_30_real;
  wire       [15:0]   myFFT_1_sdata_out_payload_30_imag;
  wire       [15:0]   myFFT_1_sdata_out_payload_31_real;
  wire       [15:0]   myFFT_1_sdata_out_payload_31_imag;
  wire       [15:0]   myFFT_1_sdata_out_payload_32_real;
  wire       [15:0]   myFFT_1_sdata_out_payload_32_imag;
  wire       [15:0]   myFFT_1_sdata_out_payload_33_real;
  wire       [15:0]   myFFT_1_sdata_out_payload_33_imag;
  wire       [15:0]   myFFT_1_sdata_out_payload_34_real;
  wire       [15:0]   myFFT_1_sdata_out_payload_34_imag;
  wire       [15:0]   myFFT_1_sdata_out_payload_35_real;
  wire       [15:0]   myFFT_1_sdata_out_payload_35_imag;
  wire       [15:0]   myFFT_1_sdata_out_payload_36_real;
  wire       [15:0]   myFFT_1_sdata_out_payload_36_imag;
  wire       [15:0]   myFFT_1_sdata_out_payload_37_real;
  wire       [15:0]   myFFT_1_sdata_out_payload_37_imag;
  wire       [15:0]   myFFT_1_sdata_out_payload_38_real;
  wire       [15:0]   myFFT_1_sdata_out_payload_38_imag;
  wire       [15:0]   myFFT_1_sdata_out_payload_39_real;
  wire       [15:0]   myFFT_1_sdata_out_payload_39_imag;
  wire       [15:0]   myFFT_1_sdata_out_payload_40_real;
  wire       [15:0]   myFFT_1_sdata_out_payload_40_imag;
  wire       [15:0]   myFFT_1_sdata_out_payload_41_real;
  wire       [15:0]   myFFT_1_sdata_out_payload_41_imag;
  wire       [15:0]   myFFT_1_sdata_out_payload_42_real;
  wire       [15:0]   myFFT_1_sdata_out_payload_42_imag;
  wire       [15:0]   myFFT_1_sdata_out_payload_43_real;
  wire       [15:0]   myFFT_1_sdata_out_payload_43_imag;
  wire       [15:0]   myFFT_1_sdata_out_payload_44_real;
  wire       [15:0]   myFFT_1_sdata_out_payload_44_imag;
  wire       [15:0]   myFFT_1_sdata_out_payload_45_real;
  wire       [15:0]   myFFT_1_sdata_out_payload_45_imag;
  wire       [15:0]   myFFT_1_sdata_out_payload_46_real;
  wire       [15:0]   myFFT_1_sdata_out_payload_46_imag;
  wire       [15:0]   myFFT_1_sdata_out_payload_47_real;
  wire       [15:0]   myFFT_1_sdata_out_payload_47_imag;
  wire       [15:0]   myFFT_1_sdata_out_payload_48_real;
  wire       [15:0]   myFFT_1_sdata_out_payload_48_imag;
  wire       [15:0]   myFFT_1_sdata_out_payload_49_real;
  wire       [15:0]   myFFT_1_sdata_out_payload_49_imag;
  wire       [15:0]   myFFT_1_sdata_out_payload_50_real;
  wire       [15:0]   myFFT_1_sdata_out_payload_50_imag;
  wire       [15:0]   myFFT_1_sdata_out_payload_51_real;
  wire       [15:0]   myFFT_1_sdata_out_payload_51_imag;
  wire       [15:0]   myFFT_1_sdata_out_payload_52_real;
  wire       [15:0]   myFFT_1_sdata_out_payload_52_imag;
  wire       [15:0]   myFFT_1_sdata_out_payload_53_real;
  wire       [15:0]   myFFT_1_sdata_out_payload_53_imag;
  wire       [15:0]   myFFT_1_sdata_out_payload_54_real;
  wire       [15:0]   myFFT_1_sdata_out_payload_54_imag;
  wire       [15:0]   myFFT_1_sdata_out_payload_55_real;
  wire       [15:0]   myFFT_1_sdata_out_payload_55_imag;
  wire       [15:0]   myFFT_1_sdata_out_payload_56_real;
  wire       [15:0]   myFFT_1_sdata_out_payload_56_imag;
  wire       [15:0]   myFFT_1_sdata_out_payload_57_real;
  wire       [15:0]   myFFT_1_sdata_out_payload_57_imag;
  wire       [15:0]   myFFT_1_sdata_out_payload_58_real;
  wire       [15:0]   myFFT_1_sdata_out_payload_58_imag;
  wire       [15:0]   myFFT_1_sdata_out_payload_59_real;
  wire       [15:0]   myFFT_1_sdata_out_payload_59_imag;
  wire       [15:0]   myFFT_1_sdata_out_payload_60_real;
  wire       [15:0]   myFFT_1_sdata_out_payload_60_imag;
  wire       [15:0]   myFFT_1_sdata_out_payload_61_real;
  wire       [15:0]   myFFT_1_sdata_out_payload_61_imag;
  wire       [15:0]   myFFT_1_sdata_out_payload_62_real;
  wire       [15:0]   myFFT_1_sdata_out_payload_62_imag;
  wire       [15:0]   myFFT_1_sdata_out_payload_63_real;
  wire       [15:0]   myFFT_1_sdata_out_payload_63_imag;
  wire       [15:0]   myFFT_1_sdata_out_payload_64_real;
  wire       [15:0]   myFFT_1_sdata_out_payload_64_imag;
  wire       [15:0]   myFFT_1_sdata_out_payload_65_real;
  wire       [15:0]   myFFT_1_sdata_out_payload_65_imag;
  wire       [15:0]   myFFT_1_sdata_out_payload_66_real;
  wire       [15:0]   myFFT_1_sdata_out_payload_66_imag;
  wire       [15:0]   myFFT_1_sdata_out_payload_67_real;
  wire       [15:0]   myFFT_1_sdata_out_payload_67_imag;
  wire       [15:0]   myFFT_1_sdata_out_payload_68_real;
  wire       [15:0]   myFFT_1_sdata_out_payload_68_imag;
  wire       [15:0]   myFFT_1_sdata_out_payload_69_real;
  wire       [15:0]   myFFT_1_sdata_out_payload_69_imag;
  wire       [15:0]   myFFT_1_sdata_out_payload_70_real;
  wire       [15:0]   myFFT_1_sdata_out_payload_70_imag;
  wire       [15:0]   myFFT_1_sdata_out_payload_71_real;
  wire       [15:0]   myFFT_1_sdata_out_payload_71_imag;
  wire       [15:0]   myFFT_1_sdata_out_payload_72_real;
  wire       [15:0]   myFFT_1_sdata_out_payload_72_imag;
  wire       [15:0]   myFFT_1_sdata_out_payload_73_real;
  wire       [15:0]   myFFT_1_sdata_out_payload_73_imag;
  wire       [15:0]   myFFT_1_sdata_out_payload_74_real;
  wire       [15:0]   myFFT_1_sdata_out_payload_74_imag;
  wire       [15:0]   myFFT_1_sdata_out_payload_75_real;
  wire       [15:0]   myFFT_1_sdata_out_payload_75_imag;
  wire       [15:0]   myFFT_1_sdata_out_payload_76_real;
  wire       [15:0]   myFFT_1_sdata_out_payload_76_imag;
  wire       [15:0]   myFFT_1_sdata_out_payload_77_real;
  wire       [15:0]   myFFT_1_sdata_out_payload_77_imag;
  wire       [15:0]   myFFT_1_sdata_out_payload_78_real;
  wire       [15:0]   myFFT_1_sdata_out_payload_78_imag;
  wire       [15:0]   myFFT_1_sdata_out_payload_79_real;
  wire       [15:0]   myFFT_1_sdata_out_payload_79_imag;
  wire       [15:0]   myFFT_1_sdata_out_payload_80_real;
  wire       [15:0]   myFFT_1_sdata_out_payload_80_imag;
  wire       [15:0]   myFFT_1_sdata_out_payload_81_real;
  wire       [15:0]   myFFT_1_sdata_out_payload_81_imag;
  wire       [15:0]   myFFT_1_sdata_out_payload_82_real;
  wire       [15:0]   myFFT_1_sdata_out_payload_82_imag;
  wire       [15:0]   myFFT_1_sdata_out_payload_83_real;
  wire       [15:0]   myFFT_1_sdata_out_payload_83_imag;
  wire       [15:0]   myFFT_1_sdata_out_payload_84_real;
  wire       [15:0]   myFFT_1_sdata_out_payload_84_imag;
  wire       [15:0]   myFFT_1_sdata_out_payload_85_real;
  wire       [15:0]   myFFT_1_sdata_out_payload_85_imag;
  wire       [15:0]   myFFT_1_sdata_out_payload_86_real;
  wire       [15:0]   myFFT_1_sdata_out_payload_86_imag;
  wire       [15:0]   myFFT_1_sdata_out_payload_87_real;
  wire       [15:0]   myFFT_1_sdata_out_payload_87_imag;
  wire       [15:0]   myFFT_1_sdata_out_payload_88_real;
  wire       [15:0]   myFFT_1_sdata_out_payload_88_imag;
  wire       [15:0]   myFFT_1_sdata_out_payload_89_real;
  wire       [15:0]   myFFT_1_sdata_out_payload_89_imag;
  wire       [15:0]   myFFT_1_sdata_out_payload_90_real;
  wire       [15:0]   myFFT_1_sdata_out_payload_90_imag;
  wire       [15:0]   myFFT_1_sdata_out_payload_91_real;
  wire       [15:0]   myFFT_1_sdata_out_payload_91_imag;
  wire       [15:0]   myFFT_1_sdata_out_payload_92_real;
  wire       [15:0]   myFFT_1_sdata_out_payload_92_imag;
  wire       [15:0]   myFFT_1_sdata_out_payload_93_real;
  wire       [15:0]   myFFT_1_sdata_out_payload_93_imag;
  wire       [15:0]   myFFT_1_sdata_out_payload_94_real;
  wire       [15:0]   myFFT_1_sdata_out_payload_94_imag;
  wire       [15:0]   myFFT_1_sdata_out_payload_95_real;
  wire       [15:0]   myFFT_1_sdata_out_payload_95_imag;
  wire       [15:0]   myFFT_1_sdata_out_payload_96_real;
  wire       [15:0]   myFFT_1_sdata_out_payload_96_imag;
  wire       [15:0]   myFFT_1_sdata_out_payload_97_real;
  wire       [15:0]   myFFT_1_sdata_out_payload_97_imag;
  wire       [15:0]   myFFT_1_sdata_out_payload_98_real;
  wire       [15:0]   myFFT_1_sdata_out_payload_98_imag;
  wire       [15:0]   myFFT_1_sdata_out_payload_99_real;
  wire       [15:0]   myFFT_1_sdata_out_payload_99_imag;
  wire       [15:0]   myFFT_1_sdata_out_payload_100_real;
  wire       [15:0]   myFFT_1_sdata_out_payload_100_imag;
  wire       [15:0]   myFFT_1_sdata_out_payload_101_real;
  wire       [15:0]   myFFT_1_sdata_out_payload_101_imag;
  wire       [15:0]   myFFT_1_sdata_out_payload_102_real;
  wire       [15:0]   myFFT_1_sdata_out_payload_102_imag;
  wire       [15:0]   myFFT_1_sdata_out_payload_103_real;
  wire       [15:0]   myFFT_1_sdata_out_payload_103_imag;
  wire       [15:0]   myFFT_1_sdata_out_payload_104_real;
  wire       [15:0]   myFFT_1_sdata_out_payload_104_imag;
  wire       [15:0]   myFFT_1_sdata_out_payload_105_real;
  wire       [15:0]   myFFT_1_sdata_out_payload_105_imag;
  wire       [15:0]   myFFT_1_sdata_out_payload_106_real;
  wire       [15:0]   myFFT_1_sdata_out_payload_106_imag;
  wire       [15:0]   myFFT_1_sdata_out_payload_107_real;
  wire       [15:0]   myFFT_1_sdata_out_payload_107_imag;
  wire       [15:0]   myFFT_1_sdata_out_payload_108_real;
  wire       [15:0]   myFFT_1_sdata_out_payload_108_imag;
  wire       [15:0]   myFFT_1_sdata_out_payload_109_real;
  wire       [15:0]   myFFT_1_sdata_out_payload_109_imag;
  wire       [15:0]   myFFT_1_sdata_out_payload_110_real;
  wire       [15:0]   myFFT_1_sdata_out_payload_110_imag;
  wire       [15:0]   myFFT_1_sdata_out_payload_111_real;
  wire       [15:0]   myFFT_1_sdata_out_payload_111_imag;
  wire       [15:0]   myFFT_1_sdata_out_payload_112_real;
  wire       [15:0]   myFFT_1_sdata_out_payload_112_imag;
  wire       [15:0]   myFFT_1_sdata_out_payload_113_real;
  wire       [15:0]   myFFT_1_sdata_out_payload_113_imag;
  wire       [15:0]   myFFT_1_sdata_out_payload_114_real;
  wire       [15:0]   myFFT_1_sdata_out_payload_114_imag;
  wire       [15:0]   myFFT_1_sdata_out_payload_115_real;
  wire       [15:0]   myFFT_1_sdata_out_payload_115_imag;
  wire       [15:0]   myFFT_1_sdata_out_payload_116_real;
  wire       [15:0]   myFFT_1_sdata_out_payload_116_imag;
  wire       [15:0]   myFFT_1_sdata_out_payload_117_real;
  wire       [15:0]   myFFT_1_sdata_out_payload_117_imag;
  wire       [15:0]   myFFT_1_sdata_out_payload_118_real;
  wire       [15:0]   myFFT_1_sdata_out_payload_118_imag;
  wire       [15:0]   myFFT_1_sdata_out_payload_119_real;
  wire       [15:0]   myFFT_1_sdata_out_payload_119_imag;
  wire       [15:0]   myFFT_1_sdata_out_payload_120_real;
  wire       [15:0]   myFFT_1_sdata_out_payload_120_imag;
  wire       [15:0]   myFFT_1_sdata_out_payload_121_real;
  wire       [15:0]   myFFT_1_sdata_out_payload_121_imag;
  wire       [15:0]   myFFT_1_sdata_out_payload_122_real;
  wire       [15:0]   myFFT_1_sdata_out_payload_122_imag;
  wire       [15:0]   myFFT_1_sdata_out_payload_123_real;
  wire       [15:0]   myFFT_1_sdata_out_payload_123_imag;
  wire       [15:0]   myFFT_1_sdata_out_payload_124_real;
  wire       [15:0]   myFFT_1_sdata_out_payload_124_imag;
  wire       [15:0]   myFFT_1_sdata_out_payload_125_real;
  wire       [15:0]   myFFT_1_sdata_out_payload_125_imag;
  wire       [15:0]   myFFT_1_sdata_out_payload_126_real;
  wire       [15:0]   myFFT_1_sdata_out_payload_126_imag;
  wire       [15:0]   myFFT_1_sdata_out_payload_127_real;
  wire       [15:0]   myFFT_1_sdata_out_payload_127_imag;
  wire       [0:0]    _zz_259;
  wire       [6:0]    _zz_260;
  wire       [0:0]    _zz_261;
  wire       [6:0]    _zz_262;
  wire       [15:0]   _zz_1;
  wire       [15:0]   _zz_2;
  reg        [15:0]   _zz_3;
  reg        [15:0]   _zz_4;
  reg        [15:0]   _zz_5;
  reg        [15:0]   _zz_6;
  reg        [15:0]   _zz_7;
  reg        [15:0]   _zz_8;
  reg        [15:0]   _zz_9;
  reg        [15:0]   _zz_10;
  reg        [15:0]   _zz_11;
  reg        [15:0]   _zz_12;
  reg        [15:0]   _zz_13;
  reg        [15:0]   _zz_14;
  reg        [15:0]   _zz_15;
  reg        [15:0]   _zz_16;
  reg        [15:0]   _zz_17;
  reg        [15:0]   _zz_18;
  reg        [15:0]   _zz_19;
  reg        [15:0]   _zz_20;
  reg        [15:0]   _zz_21;
  reg        [15:0]   _zz_22;
  reg        [15:0]   _zz_23;
  reg        [15:0]   _zz_24;
  reg        [15:0]   _zz_25;
  reg        [15:0]   _zz_26;
  reg        [15:0]   _zz_27;
  reg        [15:0]   _zz_28;
  reg        [15:0]   _zz_29;
  reg        [15:0]   _zz_30;
  reg        [15:0]   _zz_31;
  reg        [15:0]   _zz_32;
  reg        [15:0]   _zz_33;
  reg        [15:0]   _zz_34;
  reg        [15:0]   _zz_35;
  reg        [15:0]   _zz_36;
  reg        [15:0]   _zz_37;
  reg        [15:0]   _zz_38;
  reg        [15:0]   _zz_39;
  reg        [15:0]   _zz_40;
  reg        [15:0]   _zz_41;
  reg        [15:0]   _zz_42;
  reg        [15:0]   _zz_43;
  reg        [15:0]   _zz_44;
  reg        [15:0]   _zz_45;
  reg        [15:0]   _zz_46;
  reg        [15:0]   _zz_47;
  reg        [15:0]   _zz_48;
  reg        [15:0]   _zz_49;
  reg        [15:0]   _zz_50;
  reg        [15:0]   _zz_51;
  reg        [15:0]   _zz_52;
  reg        [15:0]   _zz_53;
  reg        [15:0]   _zz_54;
  reg        [15:0]   _zz_55;
  reg        [15:0]   _zz_56;
  reg        [15:0]   _zz_57;
  reg        [15:0]   _zz_58;
  reg        [15:0]   _zz_59;
  reg        [15:0]   _zz_60;
  reg        [15:0]   _zz_61;
  reg        [15:0]   _zz_62;
  reg        [15:0]   _zz_63;
  reg        [15:0]   _zz_64;
  reg        [15:0]   _zz_65;
  reg        [15:0]   _zz_66;
  reg        [15:0]   _zz_67;
  reg        [15:0]   _zz_68;
  reg        [15:0]   _zz_69;
  reg        [15:0]   _zz_70;
  reg        [15:0]   _zz_71;
  reg        [15:0]   _zz_72;
  reg        [15:0]   _zz_73;
  reg        [15:0]   _zz_74;
  reg        [15:0]   _zz_75;
  reg        [15:0]   _zz_76;
  reg        [15:0]   _zz_77;
  reg        [15:0]   _zz_78;
  reg        [15:0]   _zz_79;
  reg        [15:0]   _zz_80;
  reg        [15:0]   _zz_81;
  reg        [15:0]   _zz_82;
  reg        [15:0]   _zz_83;
  reg        [15:0]   _zz_84;
  reg        [15:0]   _zz_85;
  reg        [15:0]   _zz_86;
  reg        [15:0]   _zz_87;
  reg        [15:0]   _zz_88;
  reg        [15:0]   _zz_89;
  reg        [15:0]   _zz_90;
  reg        [15:0]   _zz_91;
  reg        [15:0]   _zz_92;
  reg        [15:0]   _zz_93;
  reg        [15:0]   _zz_94;
  reg        [15:0]   _zz_95;
  reg        [15:0]   _zz_96;
  reg        [15:0]   _zz_97;
  reg        [15:0]   _zz_98;
  reg        [15:0]   _zz_99;
  reg        [15:0]   _zz_100;
  reg        [15:0]   _zz_101;
  reg        [15:0]   _zz_102;
  reg        [15:0]   _zz_103;
  reg        [15:0]   _zz_104;
  reg        [15:0]   _zz_105;
  reg        [15:0]   _zz_106;
  reg        [15:0]   _zz_107;
  reg        [15:0]   _zz_108;
  reg        [15:0]   _zz_109;
  reg        [15:0]   _zz_110;
  reg        [15:0]   _zz_111;
  reg        [15:0]   _zz_112;
  reg        [15:0]   _zz_113;
  reg        [15:0]   _zz_114;
  reg        [15:0]   _zz_115;
  reg        [15:0]   _zz_116;
  reg        [15:0]   _zz_117;
  reg        [15:0]   _zz_118;
  reg        [15:0]   _zz_119;
  reg        [15:0]   _zz_120;
  reg        [15:0]   _zz_121;
  reg        [15:0]   _zz_122;
  reg        [15:0]   _zz_123;
  reg        [15:0]   _zz_124;
  reg        [15:0]   _zz_125;
  reg        [15:0]   _zz_126;
  reg        [15:0]   _zz_127;
  reg        [15:0]   _zz_128;
  reg        [15:0]   _zz_129;
  reg        [15:0]   _zz_130;
  reg        [15:0]   _zz_131;
  reg        [15:0]   _zz_132;
  reg        [15:0]   _zz_133;
  reg        [15:0]   _zz_134;
  reg        [15:0]   _zz_135;
  reg        [15:0]   _zz_136;
  reg        [15:0]   _zz_137;
  reg        [15:0]   _zz_138;
  reg        [15:0]   _zz_139;
  reg        [15:0]   _zz_140;
  reg        [15:0]   _zz_141;
  reg        [15:0]   _zz_142;
  reg        [15:0]   _zz_143;
  reg        [15:0]   _zz_144;
  reg        [15:0]   _zz_145;
  reg        [15:0]   _zz_146;
  reg        [15:0]   _zz_147;
  reg        [15:0]   _zz_148;
  reg        [15:0]   _zz_149;
  reg        [15:0]   _zz_150;
  reg        [15:0]   _zz_151;
  reg        [15:0]   _zz_152;
  reg        [15:0]   _zz_153;
  reg        [15:0]   _zz_154;
  reg        [15:0]   _zz_155;
  reg        [15:0]   _zz_156;
  reg        [15:0]   _zz_157;
  reg        [15:0]   _zz_158;
  reg        [15:0]   _zz_159;
  reg        [15:0]   _zz_160;
  reg        [15:0]   _zz_161;
  reg        [15:0]   _zz_162;
  reg        [15:0]   _zz_163;
  reg        [15:0]   _zz_164;
  reg        [15:0]   _zz_165;
  reg        [15:0]   _zz_166;
  reg        [15:0]   _zz_167;
  reg        [15:0]   _zz_168;
  reg        [15:0]   _zz_169;
  reg        [15:0]   _zz_170;
  reg        [15:0]   _zz_171;
  reg        [15:0]   _zz_172;
  reg        [15:0]   _zz_173;
  reg        [15:0]   _zz_174;
  reg        [15:0]   _zz_175;
  reg        [15:0]   _zz_176;
  reg        [15:0]   _zz_177;
  reg        [15:0]   _zz_178;
  reg        [15:0]   _zz_179;
  reg        [15:0]   _zz_180;
  reg        [15:0]   _zz_181;
  reg        [15:0]   _zz_182;
  reg        [15:0]   _zz_183;
  reg        [15:0]   _zz_184;
  reg        [15:0]   _zz_185;
  reg        [15:0]   _zz_186;
  reg        [15:0]   _zz_187;
  reg        [15:0]   _zz_188;
  reg        [15:0]   _zz_189;
  reg        [15:0]   _zz_190;
  reg        [15:0]   _zz_191;
  reg        [15:0]   _zz_192;
  reg        [15:0]   _zz_193;
  reg        [15:0]   _zz_194;
  reg        [15:0]   _zz_195;
  reg        [15:0]   _zz_196;
  reg        [15:0]   _zz_197;
  reg        [15:0]   _zz_198;
  reg        [15:0]   _zz_199;
  reg        [15:0]   _zz_200;
  reg        [15:0]   _zz_201;
  reg        [15:0]   _zz_202;
  reg        [15:0]   _zz_203;
  reg        [15:0]   _zz_204;
  reg        [15:0]   _zz_205;
  reg        [15:0]   _zz_206;
  reg        [15:0]   _zz_207;
  reg        [15:0]   _zz_208;
  reg        [15:0]   _zz_209;
  reg        [15:0]   _zz_210;
  reg        [15:0]   _zz_211;
  reg        [15:0]   _zz_212;
  reg        [15:0]   _zz_213;
  reg        [15:0]   _zz_214;
  reg        [15:0]   _zz_215;
  reg        [15:0]   _zz_216;
  reg        [15:0]   _zz_217;
  reg        [15:0]   _zz_218;
  reg        [15:0]   _zz_219;
  reg        [15:0]   _zz_220;
  reg        [15:0]   _zz_221;
  reg        [15:0]   _zz_222;
  reg        [15:0]   _zz_223;
  reg        [15:0]   _zz_224;
  reg        [15:0]   _zz_225;
  reg        [15:0]   _zz_226;
  reg        [15:0]   _zz_227;
  reg        [15:0]   _zz_228;
  reg        [15:0]   _zz_229;
  reg        [15:0]   _zz_230;
  reg        [15:0]   _zz_231;
  reg        [15:0]   _zz_232;
  reg        [15:0]   _zz_233;
  reg        [15:0]   _zz_234;
  reg        [15:0]   _zz_235;
  reg        [15:0]   _zz_236;
  reg        [15:0]   _zz_237;
  reg        [15:0]   _zz_238;
  reg        [15:0]   _zz_239;
  reg        [15:0]   _zz_240;
  reg        [15:0]   _zz_241;
  reg        [15:0]   _zz_242;
  reg        [15:0]   _zz_243;
  reg        [15:0]   _zz_244;
  reg        [15:0]   _zz_245;
  reg        [15:0]   _zz_246;
  reg        [15:0]   _zz_247;
  reg        [15:0]   _zz_248;
  reg        [15:0]   _zz_249;
  reg        [15:0]   _zz_250;
  reg        [15:0]   _zz_251;
  reg        [15:0]   _zz_252;
  reg        [15:0]   _zz_253;
  reg        [15:0]   _zz_254;
  reg        [15:0]   _zz_255;
  reg        [15:0]   _zz_256;
  wire                fft_input_flow_valid;
  wire       [15:0]   fft_input_flow_payload_0_real;
  wire       [15:0]   fft_input_flow_payload_0_imag;
  wire       [15:0]   fft_input_flow_payload_1_real;
  wire       [15:0]   fft_input_flow_payload_1_imag;
  wire       [15:0]   fft_input_flow_payload_2_real;
  wire       [15:0]   fft_input_flow_payload_2_imag;
  wire       [15:0]   fft_input_flow_payload_3_real;
  wire       [15:0]   fft_input_flow_payload_3_imag;
  wire       [15:0]   fft_input_flow_payload_4_real;
  wire       [15:0]   fft_input_flow_payload_4_imag;
  wire       [15:0]   fft_input_flow_payload_5_real;
  wire       [15:0]   fft_input_flow_payload_5_imag;
  wire       [15:0]   fft_input_flow_payload_6_real;
  wire       [15:0]   fft_input_flow_payload_6_imag;
  wire       [15:0]   fft_input_flow_payload_7_real;
  wire       [15:0]   fft_input_flow_payload_7_imag;
  wire       [15:0]   fft_input_flow_payload_8_real;
  wire       [15:0]   fft_input_flow_payload_8_imag;
  wire       [15:0]   fft_input_flow_payload_9_real;
  wire       [15:0]   fft_input_flow_payload_9_imag;
  wire       [15:0]   fft_input_flow_payload_10_real;
  wire       [15:0]   fft_input_flow_payload_10_imag;
  wire       [15:0]   fft_input_flow_payload_11_real;
  wire       [15:0]   fft_input_flow_payload_11_imag;
  wire       [15:0]   fft_input_flow_payload_12_real;
  wire       [15:0]   fft_input_flow_payload_12_imag;
  wire       [15:0]   fft_input_flow_payload_13_real;
  wire       [15:0]   fft_input_flow_payload_13_imag;
  wire       [15:0]   fft_input_flow_payload_14_real;
  wire       [15:0]   fft_input_flow_payload_14_imag;
  wire       [15:0]   fft_input_flow_payload_15_real;
  wire       [15:0]   fft_input_flow_payload_15_imag;
  wire       [15:0]   fft_input_flow_payload_16_real;
  wire       [15:0]   fft_input_flow_payload_16_imag;
  wire       [15:0]   fft_input_flow_payload_17_real;
  wire       [15:0]   fft_input_flow_payload_17_imag;
  wire       [15:0]   fft_input_flow_payload_18_real;
  wire       [15:0]   fft_input_flow_payload_18_imag;
  wire       [15:0]   fft_input_flow_payload_19_real;
  wire       [15:0]   fft_input_flow_payload_19_imag;
  wire       [15:0]   fft_input_flow_payload_20_real;
  wire       [15:0]   fft_input_flow_payload_20_imag;
  wire       [15:0]   fft_input_flow_payload_21_real;
  wire       [15:0]   fft_input_flow_payload_21_imag;
  wire       [15:0]   fft_input_flow_payload_22_real;
  wire       [15:0]   fft_input_flow_payload_22_imag;
  wire       [15:0]   fft_input_flow_payload_23_real;
  wire       [15:0]   fft_input_flow_payload_23_imag;
  wire       [15:0]   fft_input_flow_payload_24_real;
  wire       [15:0]   fft_input_flow_payload_24_imag;
  wire       [15:0]   fft_input_flow_payload_25_real;
  wire       [15:0]   fft_input_flow_payload_25_imag;
  wire       [15:0]   fft_input_flow_payload_26_real;
  wire       [15:0]   fft_input_flow_payload_26_imag;
  wire       [15:0]   fft_input_flow_payload_27_real;
  wire       [15:0]   fft_input_flow_payload_27_imag;
  wire       [15:0]   fft_input_flow_payload_28_real;
  wire       [15:0]   fft_input_flow_payload_28_imag;
  wire       [15:0]   fft_input_flow_payload_29_real;
  wire       [15:0]   fft_input_flow_payload_29_imag;
  wire       [15:0]   fft_input_flow_payload_30_real;
  wire       [15:0]   fft_input_flow_payload_30_imag;
  wire       [15:0]   fft_input_flow_payload_31_real;
  wire       [15:0]   fft_input_flow_payload_31_imag;
  wire       [15:0]   fft_input_flow_payload_32_real;
  wire       [15:0]   fft_input_flow_payload_32_imag;
  wire       [15:0]   fft_input_flow_payload_33_real;
  wire       [15:0]   fft_input_flow_payload_33_imag;
  wire       [15:0]   fft_input_flow_payload_34_real;
  wire       [15:0]   fft_input_flow_payload_34_imag;
  wire       [15:0]   fft_input_flow_payload_35_real;
  wire       [15:0]   fft_input_flow_payload_35_imag;
  wire       [15:0]   fft_input_flow_payload_36_real;
  wire       [15:0]   fft_input_flow_payload_36_imag;
  wire       [15:0]   fft_input_flow_payload_37_real;
  wire       [15:0]   fft_input_flow_payload_37_imag;
  wire       [15:0]   fft_input_flow_payload_38_real;
  wire       [15:0]   fft_input_flow_payload_38_imag;
  wire       [15:0]   fft_input_flow_payload_39_real;
  wire       [15:0]   fft_input_flow_payload_39_imag;
  wire       [15:0]   fft_input_flow_payload_40_real;
  wire       [15:0]   fft_input_flow_payload_40_imag;
  wire       [15:0]   fft_input_flow_payload_41_real;
  wire       [15:0]   fft_input_flow_payload_41_imag;
  wire       [15:0]   fft_input_flow_payload_42_real;
  wire       [15:0]   fft_input_flow_payload_42_imag;
  wire       [15:0]   fft_input_flow_payload_43_real;
  wire       [15:0]   fft_input_flow_payload_43_imag;
  wire       [15:0]   fft_input_flow_payload_44_real;
  wire       [15:0]   fft_input_flow_payload_44_imag;
  wire       [15:0]   fft_input_flow_payload_45_real;
  wire       [15:0]   fft_input_flow_payload_45_imag;
  wire       [15:0]   fft_input_flow_payload_46_real;
  wire       [15:0]   fft_input_flow_payload_46_imag;
  wire       [15:0]   fft_input_flow_payload_47_real;
  wire       [15:0]   fft_input_flow_payload_47_imag;
  wire       [15:0]   fft_input_flow_payload_48_real;
  wire       [15:0]   fft_input_flow_payload_48_imag;
  wire       [15:0]   fft_input_flow_payload_49_real;
  wire       [15:0]   fft_input_flow_payload_49_imag;
  wire       [15:0]   fft_input_flow_payload_50_real;
  wire       [15:0]   fft_input_flow_payload_50_imag;
  wire       [15:0]   fft_input_flow_payload_51_real;
  wire       [15:0]   fft_input_flow_payload_51_imag;
  wire       [15:0]   fft_input_flow_payload_52_real;
  wire       [15:0]   fft_input_flow_payload_52_imag;
  wire       [15:0]   fft_input_flow_payload_53_real;
  wire       [15:0]   fft_input_flow_payload_53_imag;
  wire       [15:0]   fft_input_flow_payload_54_real;
  wire       [15:0]   fft_input_flow_payload_54_imag;
  wire       [15:0]   fft_input_flow_payload_55_real;
  wire       [15:0]   fft_input_flow_payload_55_imag;
  wire       [15:0]   fft_input_flow_payload_56_real;
  wire       [15:0]   fft_input_flow_payload_56_imag;
  wire       [15:0]   fft_input_flow_payload_57_real;
  wire       [15:0]   fft_input_flow_payload_57_imag;
  wire       [15:0]   fft_input_flow_payload_58_real;
  wire       [15:0]   fft_input_flow_payload_58_imag;
  wire       [15:0]   fft_input_flow_payload_59_real;
  wire       [15:0]   fft_input_flow_payload_59_imag;
  wire       [15:0]   fft_input_flow_payload_60_real;
  wire       [15:0]   fft_input_flow_payload_60_imag;
  wire       [15:0]   fft_input_flow_payload_61_real;
  wire       [15:0]   fft_input_flow_payload_61_imag;
  wire       [15:0]   fft_input_flow_payload_62_real;
  wire       [15:0]   fft_input_flow_payload_62_imag;
  wire       [15:0]   fft_input_flow_payload_63_real;
  wire       [15:0]   fft_input_flow_payload_63_imag;
  wire       [15:0]   fft_input_flow_payload_64_real;
  wire       [15:0]   fft_input_flow_payload_64_imag;
  wire       [15:0]   fft_input_flow_payload_65_real;
  wire       [15:0]   fft_input_flow_payload_65_imag;
  wire       [15:0]   fft_input_flow_payload_66_real;
  wire       [15:0]   fft_input_flow_payload_66_imag;
  wire       [15:0]   fft_input_flow_payload_67_real;
  wire       [15:0]   fft_input_flow_payload_67_imag;
  wire       [15:0]   fft_input_flow_payload_68_real;
  wire       [15:0]   fft_input_flow_payload_68_imag;
  wire       [15:0]   fft_input_flow_payload_69_real;
  wire       [15:0]   fft_input_flow_payload_69_imag;
  wire       [15:0]   fft_input_flow_payload_70_real;
  wire       [15:0]   fft_input_flow_payload_70_imag;
  wire       [15:0]   fft_input_flow_payload_71_real;
  wire       [15:0]   fft_input_flow_payload_71_imag;
  wire       [15:0]   fft_input_flow_payload_72_real;
  wire       [15:0]   fft_input_flow_payload_72_imag;
  wire       [15:0]   fft_input_flow_payload_73_real;
  wire       [15:0]   fft_input_flow_payload_73_imag;
  wire       [15:0]   fft_input_flow_payload_74_real;
  wire       [15:0]   fft_input_flow_payload_74_imag;
  wire       [15:0]   fft_input_flow_payload_75_real;
  wire       [15:0]   fft_input_flow_payload_75_imag;
  wire       [15:0]   fft_input_flow_payload_76_real;
  wire       [15:0]   fft_input_flow_payload_76_imag;
  wire       [15:0]   fft_input_flow_payload_77_real;
  wire       [15:0]   fft_input_flow_payload_77_imag;
  wire       [15:0]   fft_input_flow_payload_78_real;
  wire       [15:0]   fft_input_flow_payload_78_imag;
  wire       [15:0]   fft_input_flow_payload_79_real;
  wire       [15:0]   fft_input_flow_payload_79_imag;
  wire       [15:0]   fft_input_flow_payload_80_real;
  wire       [15:0]   fft_input_flow_payload_80_imag;
  wire       [15:0]   fft_input_flow_payload_81_real;
  wire       [15:0]   fft_input_flow_payload_81_imag;
  wire       [15:0]   fft_input_flow_payload_82_real;
  wire       [15:0]   fft_input_flow_payload_82_imag;
  wire       [15:0]   fft_input_flow_payload_83_real;
  wire       [15:0]   fft_input_flow_payload_83_imag;
  wire       [15:0]   fft_input_flow_payload_84_real;
  wire       [15:0]   fft_input_flow_payload_84_imag;
  wire       [15:0]   fft_input_flow_payload_85_real;
  wire       [15:0]   fft_input_flow_payload_85_imag;
  wire       [15:0]   fft_input_flow_payload_86_real;
  wire       [15:0]   fft_input_flow_payload_86_imag;
  wire       [15:0]   fft_input_flow_payload_87_real;
  wire       [15:0]   fft_input_flow_payload_87_imag;
  wire       [15:0]   fft_input_flow_payload_88_real;
  wire       [15:0]   fft_input_flow_payload_88_imag;
  wire       [15:0]   fft_input_flow_payload_89_real;
  wire       [15:0]   fft_input_flow_payload_89_imag;
  wire       [15:0]   fft_input_flow_payload_90_real;
  wire       [15:0]   fft_input_flow_payload_90_imag;
  wire       [15:0]   fft_input_flow_payload_91_real;
  wire       [15:0]   fft_input_flow_payload_91_imag;
  wire       [15:0]   fft_input_flow_payload_92_real;
  wire       [15:0]   fft_input_flow_payload_92_imag;
  wire       [15:0]   fft_input_flow_payload_93_real;
  wire       [15:0]   fft_input_flow_payload_93_imag;
  wire       [15:0]   fft_input_flow_payload_94_real;
  wire       [15:0]   fft_input_flow_payload_94_imag;
  wire       [15:0]   fft_input_flow_payload_95_real;
  wire       [15:0]   fft_input_flow_payload_95_imag;
  wire       [15:0]   fft_input_flow_payload_96_real;
  wire       [15:0]   fft_input_flow_payload_96_imag;
  wire       [15:0]   fft_input_flow_payload_97_real;
  wire       [15:0]   fft_input_flow_payload_97_imag;
  wire       [15:0]   fft_input_flow_payload_98_real;
  wire       [15:0]   fft_input_flow_payload_98_imag;
  wire       [15:0]   fft_input_flow_payload_99_real;
  wire       [15:0]   fft_input_flow_payload_99_imag;
  wire       [15:0]   fft_input_flow_payload_100_real;
  wire       [15:0]   fft_input_flow_payload_100_imag;
  wire       [15:0]   fft_input_flow_payload_101_real;
  wire       [15:0]   fft_input_flow_payload_101_imag;
  wire       [15:0]   fft_input_flow_payload_102_real;
  wire       [15:0]   fft_input_flow_payload_102_imag;
  wire       [15:0]   fft_input_flow_payload_103_real;
  wire       [15:0]   fft_input_flow_payload_103_imag;
  wire       [15:0]   fft_input_flow_payload_104_real;
  wire       [15:0]   fft_input_flow_payload_104_imag;
  wire       [15:0]   fft_input_flow_payload_105_real;
  wire       [15:0]   fft_input_flow_payload_105_imag;
  wire       [15:0]   fft_input_flow_payload_106_real;
  wire       [15:0]   fft_input_flow_payload_106_imag;
  wire       [15:0]   fft_input_flow_payload_107_real;
  wire       [15:0]   fft_input_flow_payload_107_imag;
  wire       [15:0]   fft_input_flow_payload_108_real;
  wire       [15:0]   fft_input_flow_payload_108_imag;
  wire       [15:0]   fft_input_flow_payload_109_real;
  wire       [15:0]   fft_input_flow_payload_109_imag;
  wire       [15:0]   fft_input_flow_payload_110_real;
  wire       [15:0]   fft_input_flow_payload_110_imag;
  wire       [15:0]   fft_input_flow_payload_111_real;
  wire       [15:0]   fft_input_flow_payload_111_imag;
  wire       [15:0]   fft_input_flow_payload_112_real;
  wire       [15:0]   fft_input_flow_payload_112_imag;
  wire       [15:0]   fft_input_flow_payload_113_real;
  wire       [15:0]   fft_input_flow_payload_113_imag;
  wire       [15:0]   fft_input_flow_payload_114_real;
  wire       [15:0]   fft_input_flow_payload_114_imag;
  wire       [15:0]   fft_input_flow_payload_115_real;
  wire       [15:0]   fft_input_flow_payload_115_imag;
  wire       [15:0]   fft_input_flow_payload_116_real;
  wire       [15:0]   fft_input_flow_payload_116_imag;
  wire       [15:0]   fft_input_flow_payload_117_real;
  wire       [15:0]   fft_input_flow_payload_117_imag;
  wire       [15:0]   fft_input_flow_payload_118_real;
  wire       [15:0]   fft_input_flow_payload_118_imag;
  wire       [15:0]   fft_input_flow_payload_119_real;
  wire       [15:0]   fft_input_flow_payload_119_imag;
  wire       [15:0]   fft_input_flow_payload_120_real;
  wire       [15:0]   fft_input_flow_payload_120_imag;
  wire       [15:0]   fft_input_flow_payload_121_real;
  wire       [15:0]   fft_input_flow_payload_121_imag;
  wire       [15:0]   fft_input_flow_payload_122_real;
  wire       [15:0]   fft_input_flow_payload_122_imag;
  wire       [15:0]   fft_input_flow_payload_123_real;
  wire       [15:0]   fft_input_flow_payload_123_imag;
  wire       [15:0]   fft_input_flow_payload_124_real;
  wire       [15:0]   fft_input_flow_payload_124_imag;
  wire       [15:0]   fft_input_flow_payload_125_real;
  wire       [15:0]   fft_input_flow_payload_125_imag;
  wire       [15:0]   fft_input_flow_payload_126_real;
  wire       [15:0]   fft_input_flow_payload_126_imag;
  wire       [15:0]   fft_input_flow_payload_127_real;
  wire       [15:0]   fft_input_flow_payload_127_imag;
  reg                 count_up_inside_cnt_willIncrement;
  wire                count_up_inside_cnt_willClear;
  reg        [6:0]    count_up_inside_cnt_valueNext;
  reg        [6:0]    count_up_inside_cnt_value;
  wire                count_up_inside_cnt_willOverflowIfInc;
  wire                count_up_inside_cnt_willOverflow;
  reg                 myFFT_1_sdata_out_valid_regNext;
  reg                 null_cnt_willIncrement;
  wire                null_cnt_willClear;
  reg        [6:0]    null_cnt_valueNext;
  reg        [6:0]    null_cnt_value;
  wire                null_cnt_willOverflowIfInc;
  wire                null_cnt_willOverflow;
  reg                 null_cond_period_minus_1;
  wire                null_cond_period;
  reg        [15:0]   sdata_out_regs_0_real;
  reg        [15:0]   sdata_out_regs_0_imag;
  reg        [15:0]   sdata_out_regs_1_real;
  reg        [15:0]   sdata_out_regs_1_imag;
  reg        [15:0]   sdata_out_regs_2_real;
  reg        [15:0]   sdata_out_regs_2_imag;
  reg        [15:0]   sdata_out_regs_3_real;
  reg        [15:0]   sdata_out_regs_3_imag;
  reg        [15:0]   sdata_out_regs_4_real;
  reg        [15:0]   sdata_out_regs_4_imag;
  reg        [15:0]   sdata_out_regs_5_real;
  reg        [15:0]   sdata_out_regs_5_imag;
  reg        [15:0]   sdata_out_regs_6_real;
  reg        [15:0]   sdata_out_regs_6_imag;
  reg        [15:0]   sdata_out_regs_7_real;
  reg        [15:0]   sdata_out_regs_7_imag;
  reg        [15:0]   sdata_out_regs_8_real;
  reg        [15:0]   sdata_out_regs_8_imag;
  reg        [15:0]   sdata_out_regs_9_real;
  reg        [15:0]   sdata_out_regs_9_imag;
  reg        [15:0]   sdata_out_regs_10_real;
  reg        [15:0]   sdata_out_regs_10_imag;
  reg        [15:0]   sdata_out_regs_11_real;
  reg        [15:0]   sdata_out_regs_11_imag;
  reg        [15:0]   sdata_out_regs_12_real;
  reg        [15:0]   sdata_out_regs_12_imag;
  reg        [15:0]   sdata_out_regs_13_real;
  reg        [15:0]   sdata_out_regs_13_imag;
  reg        [15:0]   sdata_out_regs_14_real;
  reg        [15:0]   sdata_out_regs_14_imag;
  reg        [15:0]   sdata_out_regs_15_real;
  reg        [15:0]   sdata_out_regs_15_imag;
  reg        [15:0]   sdata_out_regs_16_real;
  reg        [15:0]   sdata_out_regs_16_imag;
  reg        [15:0]   sdata_out_regs_17_real;
  reg        [15:0]   sdata_out_regs_17_imag;
  reg        [15:0]   sdata_out_regs_18_real;
  reg        [15:0]   sdata_out_regs_18_imag;
  reg        [15:0]   sdata_out_regs_19_real;
  reg        [15:0]   sdata_out_regs_19_imag;
  reg        [15:0]   sdata_out_regs_20_real;
  reg        [15:0]   sdata_out_regs_20_imag;
  reg        [15:0]   sdata_out_regs_21_real;
  reg        [15:0]   sdata_out_regs_21_imag;
  reg        [15:0]   sdata_out_regs_22_real;
  reg        [15:0]   sdata_out_regs_22_imag;
  reg        [15:0]   sdata_out_regs_23_real;
  reg        [15:0]   sdata_out_regs_23_imag;
  reg        [15:0]   sdata_out_regs_24_real;
  reg        [15:0]   sdata_out_regs_24_imag;
  reg        [15:0]   sdata_out_regs_25_real;
  reg        [15:0]   sdata_out_regs_25_imag;
  reg        [15:0]   sdata_out_regs_26_real;
  reg        [15:0]   sdata_out_regs_26_imag;
  reg        [15:0]   sdata_out_regs_27_real;
  reg        [15:0]   sdata_out_regs_27_imag;
  reg        [15:0]   sdata_out_regs_28_real;
  reg        [15:0]   sdata_out_regs_28_imag;
  reg        [15:0]   sdata_out_regs_29_real;
  reg        [15:0]   sdata_out_regs_29_imag;
  reg        [15:0]   sdata_out_regs_30_real;
  reg        [15:0]   sdata_out_regs_30_imag;
  reg        [15:0]   sdata_out_regs_31_real;
  reg        [15:0]   sdata_out_regs_31_imag;
  reg        [15:0]   sdata_out_regs_32_real;
  reg        [15:0]   sdata_out_regs_32_imag;
  reg        [15:0]   sdata_out_regs_33_real;
  reg        [15:0]   sdata_out_regs_33_imag;
  reg        [15:0]   sdata_out_regs_34_real;
  reg        [15:0]   sdata_out_regs_34_imag;
  reg        [15:0]   sdata_out_regs_35_real;
  reg        [15:0]   sdata_out_regs_35_imag;
  reg        [15:0]   sdata_out_regs_36_real;
  reg        [15:0]   sdata_out_regs_36_imag;
  reg        [15:0]   sdata_out_regs_37_real;
  reg        [15:0]   sdata_out_regs_37_imag;
  reg        [15:0]   sdata_out_regs_38_real;
  reg        [15:0]   sdata_out_regs_38_imag;
  reg        [15:0]   sdata_out_regs_39_real;
  reg        [15:0]   sdata_out_regs_39_imag;
  reg        [15:0]   sdata_out_regs_40_real;
  reg        [15:0]   sdata_out_regs_40_imag;
  reg        [15:0]   sdata_out_regs_41_real;
  reg        [15:0]   sdata_out_regs_41_imag;
  reg        [15:0]   sdata_out_regs_42_real;
  reg        [15:0]   sdata_out_regs_42_imag;
  reg        [15:0]   sdata_out_regs_43_real;
  reg        [15:0]   sdata_out_regs_43_imag;
  reg        [15:0]   sdata_out_regs_44_real;
  reg        [15:0]   sdata_out_regs_44_imag;
  reg        [15:0]   sdata_out_regs_45_real;
  reg        [15:0]   sdata_out_regs_45_imag;
  reg        [15:0]   sdata_out_regs_46_real;
  reg        [15:0]   sdata_out_regs_46_imag;
  reg        [15:0]   sdata_out_regs_47_real;
  reg        [15:0]   sdata_out_regs_47_imag;
  reg        [15:0]   sdata_out_regs_48_real;
  reg        [15:0]   sdata_out_regs_48_imag;
  reg        [15:0]   sdata_out_regs_49_real;
  reg        [15:0]   sdata_out_regs_49_imag;
  reg        [15:0]   sdata_out_regs_50_real;
  reg        [15:0]   sdata_out_regs_50_imag;
  reg        [15:0]   sdata_out_regs_51_real;
  reg        [15:0]   sdata_out_regs_51_imag;
  reg        [15:0]   sdata_out_regs_52_real;
  reg        [15:0]   sdata_out_regs_52_imag;
  reg        [15:0]   sdata_out_regs_53_real;
  reg        [15:0]   sdata_out_regs_53_imag;
  reg        [15:0]   sdata_out_regs_54_real;
  reg        [15:0]   sdata_out_regs_54_imag;
  reg        [15:0]   sdata_out_regs_55_real;
  reg        [15:0]   sdata_out_regs_55_imag;
  reg        [15:0]   sdata_out_regs_56_real;
  reg        [15:0]   sdata_out_regs_56_imag;
  reg        [15:0]   sdata_out_regs_57_real;
  reg        [15:0]   sdata_out_regs_57_imag;
  reg        [15:0]   sdata_out_regs_58_real;
  reg        [15:0]   sdata_out_regs_58_imag;
  reg        [15:0]   sdata_out_regs_59_real;
  reg        [15:0]   sdata_out_regs_59_imag;
  reg        [15:0]   sdata_out_regs_60_real;
  reg        [15:0]   sdata_out_regs_60_imag;
  reg        [15:0]   sdata_out_regs_61_real;
  reg        [15:0]   sdata_out_regs_61_imag;
  reg        [15:0]   sdata_out_regs_62_real;
  reg        [15:0]   sdata_out_regs_62_imag;
  reg        [15:0]   sdata_out_regs_63_real;
  reg        [15:0]   sdata_out_regs_63_imag;
  reg        [15:0]   sdata_out_regs_64_real;
  reg        [15:0]   sdata_out_regs_64_imag;
  reg        [15:0]   sdata_out_regs_65_real;
  reg        [15:0]   sdata_out_regs_65_imag;
  reg        [15:0]   sdata_out_regs_66_real;
  reg        [15:0]   sdata_out_regs_66_imag;
  reg        [15:0]   sdata_out_regs_67_real;
  reg        [15:0]   sdata_out_regs_67_imag;
  reg        [15:0]   sdata_out_regs_68_real;
  reg        [15:0]   sdata_out_regs_68_imag;
  reg        [15:0]   sdata_out_regs_69_real;
  reg        [15:0]   sdata_out_regs_69_imag;
  reg        [15:0]   sdata_out_regs_70_real;
  reg        [15:0]   sdata_out_regs_70_imag;
  reg        [15:0]   sdata_out_regs_71_real;
  reg        [15:0]   sdata_out_regs_71_imag;
  reg        [15:0]   sdata_out_regs_72_real;
  reg        [15:0]   sdata_out_regs_72_imag;
  reg        [15:0]   sdata_out_regs_73_real;
  reg        [15:0]   sdata_out_regs_73_imag;
  reg        [15:0]   sdata_out_regs_74_real;
  reg        [15:0]   sdata_out_regs_74_imag;
  reg        [15:0]   sdata_out_regs_75_real;
  reg        [15:0]   sdata_out_regs_75_imag;
  reg        [15:0]   sdata_out_regs_76_real;
  reg        [15:0]   sdata_out_regs_76_imag;
  reg        [15:0]   sdata_out_regs_77_real;
  reg        [15:0]   sdata_out_regs_77_imag;
  reg        [15:0]   sdata_out_regs_78_real;
  reg        [15:0]   sdata_out_regs_78_imag;
  reg        [15:0]   sdata_out_regs_79_real;
  reg        [15:0]   sdata_out_regs_79_imag;
  reg        [15:0]   sdata_out_regs_80_real;
  reg        [15:0]   sdata_out_regs_80_imag;
  reg        [15:0]   sdata_out_regs_81_real;
  reg        [15:0]   sdata_out_regs_81_imag;
  reg        [15:0]   sdata_out_regs_82_real;
  reg        [15:0]   sdata_out_regs_82_imag;
  reg        [15:0]   sdata_out_regs_83_real;
  reg        [15:0]   sdata_out_regs_83_imag;
  reg        [15:0]   sdata_out_regs_84_real;
  reg        [15:0]   sdata_out_regs_84_imag;
  reg        [15:0]   sdata_out_regs_85_real;
  reg        [15:0]   sdata_out_regs_85_imag;
  reg        [15:0]   sdata_out_regs_86_real;
  reg        [15:0]   sdata_out_regs_86_imag;
  reg        [15:0]   sdata_out_regs_87_real;
  reg        [15:0]   sdata_out_regs_87_imag;
  reg        [15:0]   sdata_out_regs_88_real;
  reg        [15:0]   sdata_out_regs_88_imag;
  reg        [15:0]   sdata_out_regs_89_real;
  reg        [15:0]   sdata_out_regs_89_imag;
  reg        [15:0]   sdata_out_regs_90_real;
  reg        [15:0]   sdata_out_regs_90_imag;
  reg        [15:0]   sdata_out_regs_91_real;
  reg        [15:0]   sdata_out_regs_91_imag;
  reg        [15:0]   sdata_out_regs_92_real;
  reg        [15:0]   sdata_out_regs_92_imag;
  reg        [15:0]   sdata_out_regs_93_real;
  reg        [15:0]   sdata_out_regs_93_imag;
  reg        [15:0]   sdata_out_regs_94_real;
  reg        [15:0]   sdata_out_regs_94_imag;
  reg        [15:0]   sdata_out_regs_95_real;
  reg        [15:0]   sdata_out_regs_95_imag;
  reg        [15:0]   sdata_out_regs_96_real;
  reg        [15:0]   sdata_out_regs_96_imag;
  reg        [15:0]   sdata_out_regs_97_real;
  reg        [15:0]   sdata_out_regs_97_imag;
  reg        [15:0]   sdata_out_regs_98_real;
  reg        [15:0]   sdata_out_regs_98_imag;
  reg        [15:0]   sdata_out_regs_99_real;
  reg        [15:0]   sdata_out_regs_99_imag;
  reg        [15:0]   sdata_out_regs_100_real;
  reg        [15:0]   sdata_out_regs_100_imag;
  reg        [15:0]   sdata_out_regs_101_real;
  reg        [15:0]   sdata_out_regs_101_imag;
  reg        [15:0]   sdata_out_regs_102_real;
  reg        [15:0]   sdata_out_regs_102_imag;
  reg        [15:0]   sdata_out_regs_103_real;
  reg        [15:0]   sdata_out_regs_103_imag;
  reg        [15:0]   sdata_out_regs_104_real;
  reg        [15:0]   sdata_out_regs_104_imag;
  reg        [15:0]   sdata_out_regs_105_real;
  reg        [15:0]   sdata_out_regs_105_imag;
  reg        [15:0]   sdata_out_regs_106_real;
  reg        [15:0]   sdata_out_regs_106_imag;
  reg        [15:0]   sdata_out_regs_107_real;
  reg        [15:0]   sdata_out_regs_107_imag;
  reg        [15:0]   sdata_out_regs_108_real;
  reg        [15:0]   sdata_out_regs_108_imag;
  reg        [15:0]   sdata_out_regs_109_real;
  reg        [15:0]   sdata_out_regs_109_imag;
  reg        [15:0]   sdata_out_regs_110_real;
  reg        [15:0]   sdata_out_regs_110_imag;
  reg        [15:0]   sdata_out_regs_111_real;
  reg        [15:0]   sdata_out_regs_111_imag;
  reg        [15:0]   sdata_out_regs_112_real;
  reg        [15:0]   sdata_out_regs_112_imag;
  reg        [15:0]   sdata_out_regs_113_real;
  reg        [15:0]   sdata_out_regs_113_imag;
  reg        [15:0]   sdata_out_regs_114_real;
  reg        [15:0]   sdata_out_regs_114_imag;
  reg        [15:0]   sdata_out_regs_115_real;
  reg        [15:0]   sdata_out_regs_115_imag;
  reg        [15:0]   sdata_out_regs_116_real;
  reg        [15:0]   sdata_out_regs_116_imag;
  reg        [15:0]   sdata_out_regs_117_real;
  reg        [15:0]   sdata_out_regs_117_imag;
  reg        [15:0]   sdata_out_regs_118_real;
  reg        [15:0]   sdata_out_regs_118_imag;
  reg        [15:0]   sdata_out_regs_119_real;
  reg        [15:0]   sdata_out_regs_119_imag;
  reg        [15:0]   sdata_out_regs_120_real;
  reg        [15:0]   sdata_out_regs_120_imag;
  reg        [15:0]   sdata_out_regs_121_real;
  reg        [15:0]   sdata_out_regs_121_imag;
  reg        [15:0]   sdata_out_regs_122_real;
  reg        [15:0]   sdata_out_regs_122_imag;
  reg        [15:0]   sdata_out_regs_123_real;
  reg        [15:0]   sdata_out_regs_123_imag;
  reg        [15:0]   sdata_out_regs_124_real;
  reg        [15:0]   sdata_out_regs_124_imag;
  reg        [15:0]   sdata_out_regs_125_real;
  reg        [15:0]   sdata_out_regs_125_imag;
  reg        [15:0]   sdata_out_regs_126_real;
  reg        [15:0]   sdata_out_regs_126_imag;
  reg        [15:0]   sdata_out_regs_127_real;
  reg        [15:0]   sdata_out_regs_127_imag;
  wire                output_valid;
  wire       [15:0]   output_payload_real;
  wire       [15:0]   output_payload_imag;

  assign _zz_259 = count_up_inside_cnt_willIncrement;
  assign _zz_260 = {6'd0, _zz_259};
  assign _zz_261 = null_cnt_willIncrement;
  assign _zz_262 = {6'd0, _zz_261};
  MyFFT myFFT_1 (
    .io_data_in_valid               (fft_input_flow_valid                      ), //i
    .io_data_in_payload_0_real      (fft_input_flow_payload_0_real[15:0]       ), //i
    .io_data_in_payload_0_imag      (fft_input_flow_payload_0_imag[15:0]       ), //i
    .io_data_in_payload_1_real      (fft_input_flow_payload_1_real[15:0]       ), //i
    .io_data_in_payload_1_imag      (fft_input_flow_payload_1_imag[15:0]       ), //i
    .io_data_in_payload_2_real      (fft_input_flow_payload_2_real[15:0]       ), //i
    .io_data_in_payload_2_imag      (fft_input_flow_payload_2_imag[15:0]       ), //i
    .io_data_in_payload_3_real      (fft_input_flow_payload_3_real[15:0]       ), //i
    .io_data_in_payload_3_imag      (fft_input_flow_payload_3_imag[15:0]       ), //i
    .io_data_in_payload_4_real      (fft_input_flow_payload_4_real[15:0]       ), //i
    .io_data_in_payload_4_imag      (fft_input_flow_payload_4_imag[15:0]       ), //i
    .io_data_in_payload_5_real      (fft_input_flow_payload_5_real[15:0]       ), //i
    .io_data_in_payload_5_imag      (fft_input_flow_payload_5_imag[15:0]       ), //i
    .io_data_in_payload_6_real      (fft_input_flow_payload_6_real[15:0]       ), //i
    .io_data_in_payload_6_imag      (fft_input_flow_payload_6_imag[15:0]       ), //i
    .io_data_in_payload_7_real      (fft_input_flow_payload_7_real[15:0]       ), //i
    .io_data_in_payload_7_imag      (fft_input_flow_payload_7_imag[15:0]       ), //i
    .io_data_in_payload_8_real      (fft_input_flow_payload_8_real[15:0]       ), //i
    .io_data_in_payload_8_imag      (fft_input_flow_payload_8_imag[15:0]       ), //i
    .io_data_in_payload_9_real      (fft_input_flow_payload_9_real[15:0]       ), //i
    .io_data_in_payload_9_imag      (fft_input_flow_payload_9_imag[15:0]       ), //i
    .io_data_in_payload_10_real     (fft_input_flow_payload_10_real[15:0]      ), //i
    .io_data_in_payload_10_imag     (fft_input_flow_payload_10_imag[15:0]      ), //i
    .io_data_in_payload_11_real     (fft_input_flow_payload_11_real[15:0]      ), //i
    .io_data_in_payload_11_imag     (fft_input_flow_payload_11_imag[15:0]      ), //i
    .io_data_in_payload_12_real     (fft_input_flow_payload_12_real[15:0]      ), //i
    .io_data_in_payload_12_imag     (fft_input_flow_payload_12_imag[15:0]      ), //i
    .io_data_in_payload_13_real     (fft_input_flow_payload_13_real[15:0]      ), //i
    .io_data_in_payload_13_imag     (fft_input_flow_payload_13_imag[15:0]      ), //i
    .io_data_in_payload_14_real     (fft_input_flow_payload_14_real[15:0]      ), //i
    .io_data_in_payload_14_imag     (fft_input_flow_payload_14_imag[15:0]      ), //i
    .io_data_in_payload_15_real     (fft_input_flow_payload_15_real[15:0]      ), //i
    .io_data_in_payload_15_imag     (fft_input_flow_payload_15_imag[15:0]      ), //i
    .io_data_in_payload_16_real     (fft_input_flow_payload_16_real[15:0]      ), //i
    .io_data_in_payload_16_imag     (fft_input_flow_payload_16_imag[15:0]      ), //i
    .io_data_in_payload_17_real     (fft_input_flow_payload_17_real[15:0]      ), //i
    .io_data_in_payload_17_imag     (fft_input_flow_payload_17_imag[15:0]      ), //i
    .io_data_in_payload_18_real     (fft_input_flow_payload_18_real[15:0]      ), //i
    .io_data_in_payload_18_imag     (fft_input_flow_payload_18_imag[15:0]      ), //i
    .io_data_in_payload_19_real     (fft_input_flow_payload_19_real[15:0]      ), //i
    .io_data_in_payload_19_imag     (fft_input_flow_payload_19_imag[15:0]      ), //i
    .io_data_in_payload_20_real     (fft_input_flow_payload_20_real[15:0]      ), //i
    .io_data_in_payload_20_imag     (fft_input_flow_payload_20_imag[15:0]      ), //i
    .io_data_in_payload_21_real     (fft_input_flow_payload_21_real[15:0]      ), //i
    .io_data_in_payload_21_imag     (fft_input_flow_payload_21_imag[15:0]      ), //i
    .io_data_in_payload_22_real     (fft_input_flow_payload_22_real[15:0]      ), //i
    .io_data_in_payload_22_imag     (fft_input_flow_payload_22_imag[15:0]      ), //i
    .io_data_in_payload_23_real     (fft_input_flow_payload_23_real[15:0]      ), //i
    .io_data_in_payload_23_imag     (fft_input_flow_payload_23_imag[15:0]      ), //i
    .io_data_in_payload_24_real     (fft_input_flow_payload_24_real[15:0]      ), //i
    .io_data_in_payload_24_imag     (fft_input_flow_payload_24_imag[15:0]      ), //i
    .io_data_in_payload_25_real     (fft_input_flow_payload_25_real[15:0]      ), //i
    .io_data_in_payload_25_imag     (fft_input_flow_payload_25_imag[15:0]      ), //i
    .io_data_in_payload_26_real     (fft_input_flow_payload_26_real[15:0]      ), //i
    .io_data_in_payload_26_imag     (fft_input_flow_payload_26_imag[15:0]      ), //i
    .io_data_in_payload_27_real     (fft_input_flow_payload_27_real[15:0]      ), //i
    .io_data_in_payload_27_imag     (fft_input_flow_payload_27_imag[15:0]      ), //i
    .io_data_in_payload_28_real     (fft_input_flow_payload_28_real[15:0]      ), //i
    .io_data_in_payload_28_imag     (fft_input_flow_payload_28_imag[15:0]      ), //i
    .io_data_in_payload_29_real     (fft_input_flow_payload_29_real[15:0]      ), //i
    .io_data_in_payload_29_imag     (fft_input_flow_payload_29_imag[15:0]      ), //i
    .io_data_in_payload_30_real     (fft_input_flow_payload_30_real[15:0]      ), //i
    .io_data_in_payload_30_imag     (fft_input_flow_payload_30_imag[15:0]      ), //i
    .io_data_in_payload_31_real     (fft_input_flow_payload_31_real[15:0]      ), //i
    .io_data_in_payload_31_imag     (fft_input_flow_payload_31_imag[15:0]      ), //i
    .io_data_in_payload_32_real     (fft_input_flow_payload_32_real[15:0]      ), //i
    .io_data_in_payload_32_imag     (fft_input_flow_payload_32_imag[15:0]      ), //i
    .io_data_in_payload_33_real     (fft_input_flow_payload_33_real[15:0]      ), //i
    .io_data_in_payload_33_imag     (fft_input_flow_payload_33_imag[15:0]      ), //i
    .io_data_in_payload_34_real     (fft_input_flow_payload_34_real[15:0]      ), //i
    .io_data_in_payload_34_imag     (fft_input_flow_payload_34_imag[15:0]      ), //i
    .io_data_in_payload_35_real     (fft_input_flow_payload_35_real[15:0]      ), //i
    .io_data_in_payload_35_imag     (fft_input_flow_payload_35_imag[15:0]      ), //i
    .io_data_in_payload_36_real     (fft_input_flow_payload_36_real[15:0]      ), //i
    .io_data_in_payload_36_imag     (fft_input_flow_payload_36_imag[15:0]      ), //i
    .io_data_in_payload_37_real     (fft_input_flow_payload_37_real[15:0]      ), //i
    .io_data_in_payload_37_imag     (fft_input_flow_payload_37_imag[15:0]      ), //i
    .io_data_in_payload_38_real     (fft_input_flow_payload_38_real[15:0]      ), //i
    .io_data_in_payload_38_imag     (fft_input_flow_payload_38_imag[15:0]      ), //i
    .io_data_in_payload_39_real     (fft_input_flow_payload_39_real[15:0]      ), //i
    .io_data_in_payload_39_imag     (fft_input_flow_payload_39_imag[15:0]      ), //i
    .io_data_in_payload_40_real     (fft_input_flow_payload_40_real[15:0]      ), //i
    .io_data_in_payload_40_imag     (fft_input_flow_payload_40_imag[15:0]      ), //i
    .io_data_in_payload_41_real     (fft_input_flow_payload_41_real[15:0]      ), //i
    .io_data_in_payload_41_imag     (fft_input_flow_payload_41_imag[15:0]      ), //i
    .io_data_in_payload_42_real     (fft_input_flow_payload_42_real[15:0]      ), //i
    .io_data_in_payload_42_imag     (fft_input_flow_payload_42_imag[15:0]      ), //i
    .io_data_in_payload_43_real     (fft_input_flow_payload_43_real[15:0]      ), //i
    .io_data_in_payload_43_imag     (fft_input_flow_payload_43_imag[15:0]      ), //i
    .io_data_in_payload_44_real     (fft_input_flow_payload_44_real[15:0]      ), //i
    .io_data_in_payload_44_imag     (fft_input_flow_payload_44_imag[15:0]      ), //i
    .io_data_in_payload_45_real     (fft_input_flow_payload_45_real[15:0]      ), //i
    .io_data_in_payload_45_imag     (fft_input_flow_payload_45_imag[15:0]      ), //i
    .io_data_in_payload_46_real     (fft_input_flow_payload_46_real[15:0]      ), //i
    .io_data_in_payload_46_imag     (fft_input_flow_payload_46_imag[15:0]      ), //i
    .io_data_in_payload_47_real     (fft_input_flow_payload_47_real[15:0]      ), //i
    .io_data_in_payload_47_imag     (fft_input_flow_payload_47_imag[15:0]      ), //i
    .io_data_in_payload_48_real     (fft_input_flow_payload_48_real[15:0]      ), //i
    .io_data_in_payload_48_imag     (fft_input_flow_payload_48_imag[15:0]      ), //i
    .io_data_in_payload_49_real     (fft_input_flow_payload_49_real[15:0]      ), //i
    .io_data_in_payload_49_imag     (fft_input_flow_payload_49_imag[15:0]      ), //i
    .io_data_in_payload_50_real     (fft_input_flow_payload_50_real[15:0]      ), //i
    .io_data_in_payload_50_imag     (fft_input_flow_payload_50_imag[15:0]      ), //i
    .io_data_in_payload_51_real     (fft_input_flow_payload_51_real[15:0]      ), //i
    .io_data_in_payload_51_imag     (fft_input_flow_payload_51_imag[15:0]      ), //i
    .io_data_in_payload_52_real     (fft_input_flow_payload_52_real[15:0]      ), //i
    .io_data_in_payload_52_imag     (fft_input_flow_payload_52_imag[15:0]      ), //i
    .io_data_in_payload_53_real     (fft_input_flow_payload_53_real[15:0]      ), //i
    .io_data_in_payload_53_imag     (fft_input_flow_payload_53_imag[15:0]      ), //i
    .io_data_in_payload_54_real     (fft_input_flow_payload_54_real[15:0]      ), //i
    .io_data_in_payload_54_imag     (fft_input_flow_payload_54_imag[15:0]      ), //i
    .io_data_in_payload_55_real     (fft_input_flow_payload_55_real[15:0]      ), //i
    .io_data_in_payload_55_imag     (fft_input_flow_payload_55_imag[15:0]      ), //i
    .io_data_in_payload_56_real     (fft_input_flow_payload_56_real[15:0]      ), //i
    .io_data_in_payload_56_imag     (fft_input_flow_payload_56_imag[15:0]      ), //i
    .io_data_in_payload_57_real     (fft_input_flow_payload_57_real[15:0]      ), //i
    .io_data_in_payload_57_imag     (fft_input_flow_payload_57_imag[15:0]      ), //i
    .io_data_in_payload_58_real     (fft_input_flow_payload_58_real[15:0]      ), //i
    .io_data_in_payload_58_imag     (fft_input_flow_payload_58_imag[15:0]      ), //i
    .io_data_in_payload_59_real     (fft_input_flow_payload_59_real[15:0]      ), //i
    .io_data_in_payload_59_imag     (fft_input_flow_payload_59_imag[15:0]      ), //i
    .io_data_in_payload_60_real     (fft_input_flow_payload_60_real[15:0]      ), //i
    .io_data_in_payload_60_imag     (fft_input_flow_payload_60_imag[15:0]      ), //i
    .io_data_in_payload_61_real     (fft_input_flow_payload_61_real[15:0]      ), //i
    .io_data_in_payload_61_imag     (fft_input_flow_payload_61_imag[15:0]      ), //i
    .io_data_in_payload_62_real     (fft_input_flow_payload_62_real[15:0]      ), //i
    .io_data_in_payload_62_imag     (fft_input_flow_payload_62_imag[15:0]      ), //i
    .io_data_in_payload_63_real     (fft_input_flow_payload_63_real[15:0]      ), //i
    .io_data_in_payload_63_imag     (fft_input_flow_payload_63_imag[15:0]      ), //i
    .io_data_in_payload_64_real     (fft_input_flow_payload_64_real[15:0]      ), //i
    .io_data_in_payload_64_imag     (fft_input_flow_payload_64_imag[15:0]      ), //i
    .io_data_in_payload_65_real     (fft_input_flow_payload_65_real[15:0]      ), //i
    .io_data_in_payload_65_imag     (fft_input_flow_payload_65_imag[15:0]      ), //i
    .io_data_in_payload_66_real     (fft_input_flow_payload_66_real[15:0]      ), //i
    .io_data_in_payload_66_imag     (fft_input_flow_payload_66_imag[15:0]      ), //i
    .io_data_in_payload_67_real     (fft_input_flow_payload_67_real[15:0]      ), //i
    .io_data_in_payload_67_imag     (fft_input_flow_payload_67_imag[15:0]      ), //i
    .io_data_in_payload_68_real     (fft_input_flow_payload_68_real[15:0]      ), //i
    .io_data_in_payload_68_imag     (fft_input_flow_payload_68_imag[15:0]      ), //i
    .io_data_in_payload_69_real     (fft_input_flow_payload_69_real[15:0]      ), //i
    .io_data_in_payload_69_imag     (fft_input_flow_payload_69_imag[15:0]      ), //i
    .io_data_in_payload_70_real     (fft_input_flow_payload_70_real[15:0]      ), //i
    .io_data_in_payload_70_imag     (fft_input_flow_payload_70_imag[15:0]      ), //i
    .io_data_in_payload_71_real     (fft_input_flow_payload_71_real[15:0]      ), //i
    .io_data_in_payload_71_imag     (fft_input_flow_payload_71_imag[15:0]      ), //i
    .io_data_in_payload_72_real     (fft_input_flow_payload_72_real[15:0]      ), //i
    .io_data_in_payload_72_imag     (fft_input_flow_payload_72_imag[15:0]      ), //i
    .io_data_in_payload_73_real     (fft_input_flow_payload_73_real[15:0]      ), //i
    .io_data_in_payload_73_imag     (fft_input_flow_payload_73_imag[15:0]      ), //i
    .io_data_in_payload_74_real     (fft_input_flow_payload_74_real[15:0]      ), //i
    .io_data_in_payload_74_imag     (fft_input_flow_payload_74_imag[15:0]      ), //i
    .io_data_in_payload_75_real     (fft_input_flow_payload_75_real[15:0]      ), //i
    .io_data_in_payload_75_imag     (fft_input_flow_payload_75_imag[15:0]      ), //i
    .io_data_in_payload_76_real     (fft_input_flow_payload_76_real[15:0]      ), //i
    .io_data_in_payload_76_imag     (fft_input_flow_payload_76_imag[15:0]      ), //i
    .io_data_in_payload_77_real     (fft_input_flow_payload_77_real[15:0]      ), //i
    .io_data_in_payload_77_imag     (fft_input_flow_payload_77_imag[15:0]      ), //i
    .io_data_in_payload_78_real     (fft_input_flow_payload_78_real[15:0]      ), //i
    .io_data_in_payload_78_imag     (fft_input_flow_payload_78_imag[15:0]      ), //i
    .io_data_in_payload_79_real     (fft_input_flow_payload_79_real[15:0]      ), //i
    .io_data_in_payload_79_imag     (fft_input_flow_payload_79_imag[15:0]      ), //i
    .io_data_in_payload_80_real     (fft_input_flow_payload_80_real[15:0]      ), //i
    .io_data_in_payload_80_imag     (fft_input_flow_payload_80_imag[15:0]      ), //i
    .io_data_in_payload_81_real     (fft_input_flow_payload_81_real[15:0]      ), //i
    .io_data_in_payload_81_imag     (fft_input_flow_payload_81_imag[15:0]      ), //i
    .io_data_in_payload_82_real     (fft_input_flow_payload_82_real[15:0]      ), //i
    .io_data_in_payload_82_imag     (fft_input_flow_payload_82_imag[15:0]      ), //i
    .io_data_in_payload_83_real     (fft_input_flow_payload_83_real[15:0]      ), //i
    .io_data_in_payload_83_imag     (fft_input_flow_payload_83_imag[15:0]      ), //i
    .io_data_in_payload_84_real     (fft_input_flow_payload_84_real[15:0]      ), //i
    .io_data_in_payload_84_imag     (fft_input_flow_payload_84_imag[15:0]      ), //i
    .io_data_in_payload_85_real     (fft_input_flow_payload_85_real[15:0]      ), //i
    .io_data_in_payload_85_imag     (fft_input_flow_payload_85_imag[15:0]      ), //i
    .io_data_in_payload_86_real     (fft_input_flow_payload_86_real[15:0]      ), //i
    .io_data_in_payload_86_imag     (fft_input_flow_payload_86_imag[15:0]      ), //i
    .io_data_in_payload_87_real     (fft_input_flow_payload_87_real[15:0]      ), //i
    .io_data_in_payload_87_imag     (fft_input_flow_payload_87_imag[15:0]      ), //i
    .io_data_in_payload_88_real     (fft_input_flow_payload_88_real[15:0]      ), //i
    .io_data_in_payload_88_imag     (fft_input_flow_payload_88_imag[15:0]      ), //i
    .io_data_in_payload_89_real     (fft_input_flow_payload_89_real[15:0]      ), //i
    .io_data_in_payload_89_imag     (fft_input_flow_payload_89_imag[15:0]      ), //i
    .io_data_in_payload_90_real     (fft_input_flow_payload_90_real[15:0]      ), //i
    .io_data_in_payload_90_imag     (fft_input_flow_payload_90_imag[15:0]      ), //i
    .io_data_in_payload_91_real     (fft_input_flow_payload_91_real[15:0]      ), //i
    .io_data_in_payload_91_imag     (fft_input_flow_payload_91_imag[15:0]      ), //i
    .io_data_in_payload_92_real     (fft_input_flow_payload_92_real[15:0]      ), //i
    .io_data_in_payload_92_imag     (fft_input_flow_payload_92_imag[15:0]      ), //i
    .io_data_in_payload_93_real     (fft_input_flow_payload_93_real[15:0]      ), //i
    .io_data_in_payload_93_imag     (fft_input_flow_payload_93_imag[15:0]      ), //i
    .io_data_in_payload_94_real     (fft_input_flow_payload_94_real[15:0]      ), //i
    .io_data_in_payload_94_imag     (fft_input_flow_payload_94_imag[15:0]      ), //i
    .io_data_in_payload_95_real     (fft_input_flow_payload_95_real[15:0]      ), //i
    .io_data_in_payload_95_imag     (fft_input_flow_payload_95_imag[15:0]      ), //i
    .io_data_in_payload_96_real     (fft_input_flow_payload_96_real[15:0]      ), //i
    .io_data_in_payload_96_imag     (fft_input_flow_payload_96_imag[15:0]      ), //i
    .io_data_in_payload_97_real     (fft_input_flow_payload_97_real[15:0]      ), //i
    .io_data_in_payload_97_imag     (fft_input_flow_payload_97_imag[15:0]      ), //i
    .io_data_in_payload_98_real     (fft_input_flow_payload_98_real[15:0]      ), //i
    .io_data_in_payload_98_imag     (fft_input_flow_payload_98_imag[15:0]      ), //i
    .io_data_in_payload_99_real     (fft_input_flow_payload_99_real[15:0]      ), //i
    .io_data_in_payload_99_imag     (fft_input_flow_payload_99_imag[15:0]      ), //i
    .io_data_in_payload_100_real    (fft_input_flow_payload_100_real[15:0]     ), //i
    .io_data_in_payload_100_imag    (fft_input_flow_payload_100_imag[15:0]     ), //i
    .io_data_in_payload_101_real    (fft_input_flow_payload_101_real[15:0]     ), //i
    .io_data_in_payload_101_imag    (fft_input_flow_payload_101_imag[15:0]     ), //i
    .io_data_in_payload_102_real    (fft_input_flow_payload_102_real[15:0]     ), //i
    .io_data_in_payload_102_imag    (fft_input_flow_payload_102_imag[15:0]     ), //i
    .io_data_in_payload_103_real    (fft_input_flow_payload_103_real[15:0]     ), //i
    .io_data_in_payload_103_imag    (fft_input_flow_payload_103_imag[15:0]     ), //i
    .io_data_in_payload_104_real    (fft_input_flow_payload_104_real[15:0]     ), //i
    .io_data_in_payload_104_imag    (fft_input_flow_payload_104_imag[15:0]     ), //i
    .io_data_in_payload_105_real    (fft_input_flow_payload_105_real[15:0]     ), //i
    .io_data_in_payload_105_imag    (fft_input_flow_payload_105_imag[15:0]     ), //i
    .io_data_in_payload_106_real    (fft_input_flow_payload_106_real[15:0]     ), //i
    .io_data_in_payload_106_imag    (fft_input_flow_payload_106_imag[15:0]     ), //i
    .io_data_in_payload_107_real    (fft_input_flow_payload_107_real[15:0]     ), //i
    .io_data_in_payload_107_imag    (fft_input_flow_payload_107_imag[15:0]     ), //i
    .io_data_in_payload_108_real    (fft_input_flow_payload_108_real[15:0]     ), //i
    .io_data_in_payload_108_imag    (fft_input_flow_payload_108_imag[15:0]     ), //i
    .io_data_in_payload_109_real    (fft_input_flow_payload_109_real[15:0]     ), //i
    .io_data_in_payload_109_imag    (fft_input_flow_payload_109_imag[15:0]     ), //i
    .io_data_in_payload_110_real    (fft_input_flow_payload_110_real[15:0]     ), //i
    .io_data_in_payload_110_imag    (fft_input_flow_payload_110_imag[15:0]     ), //i
    .io_data_in_payload_111_real    (fft_input_flow_payload_111_real[15:0]     ), //i
    .io_data_in_payload_111_imag    (fft_input_flow_payload_111_imag[15:0]     ), //i
    .io_data_in_payload_112_real    (fft_input_flow_payload_112_real[15:0]     ), //i
    .io_data_in_payload_112_imag    (fft_input_flow_payload_112_imag[15:0]     ), //i
    .io_data_in_payload_113_real    (fft_input_flow_payload_113_real[15:0]     ), //i
    .io_data_in_payload_113_imag    (fft_input_flow_payload_113_imag[15:0]     ), //i
    .io_data_in_payload_114_real    (fft_input_flow_payload_114_real[15:0]     ), //i
    .io_data_in_payload_114_imag    (fft_input_flow_payload_114_imag[15:0]     ), //i
    .io_data_in_payload_115_real    (fft_input_flow_payload_115_real[15:0]     ), //i
    .io_data_in_payload_115_imag    (fft_input_flow_payload_115_imag[15:0]     ), //i
    .io_data_in_payload_116_real    (fft_input_flow_payload_116_real[15:0]     ), //i
    .io_data_in_payload_116_imag    (fft_input_flow_payload_116_imag[15:0]     ), //i
    .io_data_in_payload_117_real    (fft_input_flow_payload_117_real[15:0]     ), //i
    .io_data_in_payload_117_imag    (fft_input_flow_payload_117_imag[15:0]     ), //i
    .io_data_in_payload_118_real    (fft_input_flow_payload_118_real[15:0]     ), //i
    .io_data_in_payload_118_imag    (fft_input_flow_payload_118_imag[15:0]     ), //i
    .io_data_in_payload_119_real    (fft_input_flow_payload_119_real[15:0]     ), //i
    .io_data_in_payload_119_imag    (fft_input_flow_payload_119_imag[15:0]     ), //i
    .io_data_in_payload_120_real    (fft_input_flow_payload_120_real[15:0]     ), //i
    .io_data_in_payload_120_imag    (fft_input_flow_payload_120_imag[15:0]     ), //i
    .io_data_in_payload_121_real    (fft_input_flow_payload_121_real[15:0]     ), //i
    .io_data_in_payload_121_imag    (fft_input_flow_payload_121_imag[15:0]     ), //i
    .io_data_in_payload_122_real    (fft_input_flow_payload_122_real[15:0]     ), //i
    .io_data_in_payload_122_imag    (fft_input_flow_payload_122_imag[15:0]     ), //i
    .io_data_in_payload_123_real    (fft_input_flow_payload_123_real[15:0]     ), //i
    .io_data_in_payload_123_imag    (fft_input_flow_payload_123_imag[15:0]     ), //i
    .io_data_in_payload_124_real    (fft_input_flow_payload_124_real[15:0]     ), //i
    .io_data_in_payload_124_imag    (fft_input_flow_payload_124_imag[15:0]     ), //i
    .io_data_in_payload_125_real    (fft_input_flow_payload_125_real[15:0]     ), //i
    .io_data_in_payload_125_imag    (fft_input_flow_payload_125_imag[15:0]     ), //i
    .io_data_in_payload_126_real    (fft_input_flow_payload_126_real[15:0]     ), //i
    .io_data_in_payload_126_imag    (fft_input_flow_payload_126_imag[15:0]     ), //i
    .io_data_in_payload_127_real    (fft_input_flow_payload_127_real[15:0]     ), //i
    .io_data_in_payload_127_imag    (fft_input_flow_payload_127_imag[15:0]     ), //i
    .sdata_out_valid                (myFFT_1_sdata_out_valid                   ), //o
    .sdata_out_payload_0_real       (myFFT_1_sdata_out_payload_0_real[15:0]    ), //o
    .sdata_out_payload_0_imag       (myFFT_1_sdata_out_payload_0_imag[15:0]    ), //o
    .sdata_out_payload_1_real       (myFFT_1_sdata_out_payload_1_real[15:0]    ), //o
    .sdata_out_payload_1_imag       (myFFT_1_sdata_out_payload_1_imag[15:0]    ), //o
    .sdata_out_payload_2_real       (myFFT_1_sdata_out_payload_2_real[15:0]    ), //o
    .sdata_out_payload_2_imag       (myFFT_1_sdata_out_payload_2_imag[15:0]    ), //o
    .sdata_out_payload_3_real       (myFFT_1_sdata_out_payload_3_real[15:0]    ), //o
    .sdata_out_payload_3_imag       (myFFT_1_sdata_out_payload_3_imag[15:0]    ), //o
    .sdata_out_payload_4_real       (myFFT_1_sdata_out_payload_4_real[15:0]    ), //o
    .sdata_out_payload_4_imag       (myFFT_1_sdata_out_payload_4_imag[15:0]    ), //o
    .sdata_out_payload_5_real       (myFFT_1_sdata_out_payload_5_real[15:0]    ), //o
    .sdata_out_payload_5_imag       (myFFT_1_sdata_out_payload_5_imag[15:0]    ), //o
    .sdata_out_payload_6_real       (myFFT_1_sdata_out_payload_6_real[15:0]    ), //o
    .sdata_out_payload_6_imag       (myFFT_1_sdata_out_payload_6_imag[15:0]    ), //o
    .sdata_out_payload_7_real       (myFFT_1_sdata_out_payload_7_real[15:0]    ), //o
    .sdata_out_payload_7_imag       (myFFT_1_sdata_out_payload_7_imag[15:0]    ), //o
    .sdata_out_payload_8_real       (myFFT_1_sdata_out_payload_8_real[15:0]    ), //o
    .sdata_out_payload_8_imag       (myFFT_1_sdata_out_payload_8_imag[15:0]    ), //o
    .sdata_out_payload_9_real       (myFFT_1_sdata_out_payload_9_real[15:0]    ), //o
    .sdata_out_payload_9_imag       (myFFT_1_sdata_out_payload_9_imag[15:0]    ), //o
    .sdata_out_payload_10_real      (myFFT_1_sdata_out_payload_10_real[15:0]   ), //o
    .sdata_out_payload_10_imag      (myFFT_1_sdata_out_payload_10_imag[15:0]   ), //o
    .sdata_out_payload_11_real      (myFFT_1_sdata_out_payload_11_real[15:0]   ), //o
    .sdata_out_payload_11_imag      (myFFT_1_sdata_out_payload_11_imag[15:0]   ), //o
    .sdata_out_payload_12_real      (myFFT_1_sdata_out_payload_12_real[15:0]   ), //o
    .sdata_out_payload_12_imag      (myFFT_1_sdata_out_payload_12_imag[15:0]   ), //o
    .sdata_out_payload_13_real      (myFFT_1_sdata_out_payload_13_real[15:0]   ), //o
    .sdata_out_payload_13_imag      (myFFT_1_sdata_out_payload_13_imag[15:0]   ), //o
    .sdata_out_payload_14_real      (myFFT_1_sdata_out_payload_14_real[15:0]   ), //o
    .sdata_out_payload_14_imag      (myFFT_1_sdata_out_payload_14_imag[15:0]   ), //o
    .sdata_out_payload_15_real      (myFFT_1_sdata_out_payload_15_real[15:0]   ), //o
    .sdata_out_payload_15_imag      (myFFT_1_sdata_out_payload_15_imag[15:0]   ), //o
    .sdata_out_payload_16_real      (myFFT_1_sdata_out_payload_16_real[15:0]   ), //o
    .sdata_out_payload_16_imag      (myFFT_1_sdata_out_payload_16_imag[15:0]   ), //o
    .sdata_out_payload_17_real      (myFFT_1_sdata_out_payload_17_real[15:0]   ), //o
    .sdata_out_payload_17_imag      (myFFT_1_sdata_out_payload_17_imag[15:0]   ), //o
    .sdata_out_payload_18_real      (myFFT_1_sdata_out_payload_18_real[15:0]   ), //o
    .sdata_out_payload_18_imag      (myFFT_1_sdata_out_payload_18_imag[15:0]   ), //o
    .sdata_out_payload_19_real      (myFFT_1_sdata_out_payload_19_real[15:0]   ), //o
    .sdata_out_payload_19_imag      (myFFT_1_sdata_out_payload_19_imag[15:0]   ), //o
    .sdata_out_payload_20_real      (myFFT_1_sdata_out_payload_20_real[15:0]   ), //o
    .sdata_out_payload_20_imag      (myFFT_1_sdata_out_payload_20_imag[15:0]   ), //o
    .sdata_out_payload_21_real      (myFFT_1_sdata_out_payload_21_real[15:0]   ), //o
    .sdata_out_payload_21_imag      (myFFT_1_sdata_out_payload_21_imag[15:0]   ), //o
    .sdata_out_payload_22_real      (myFFT_1_sdata_out_payload_22_real[15:0]   ), //o
    .sdata_out_payload_22_imag      (myFFT_1_sdata_out_payload_22_imag[15:0]   ), //o
    .sdata_out_payload_23_real      (myFFT_1_sdata_out_payload_23_real[15:0]   ), //o
    .sdata_out_payload_23_imag      (myFFT_1_sdata_out_payload_23_imag[15:0]   ), //o
    .sdata_out_payload_24_real      (myFFT_1_sdata_out_payload_24_real[15:0]   ), //o
    .sdata_out_payload_24_imag      (myFFT_1_sdata_out_payload_24_imag[15:0]   ), //o
    .sdata_out_payload_25_real      (myFFT_1_sdata_out_payload_25_real[15:0]   ), //o
    .sdata_out_payload_25_imag      (myFFT_1_sdata_out_payload_25_imag[15:0]   ), //o
    .sdata_out_payload_26_real      (myFFT_1_sdata_out_payload_26_real[15:0]   ), //o
    .sdata_out_payload_26_imag      (myFFT_1_sdata_out_payload_26_imag[15:0]   ), //o
    .sdata_out_payload_27_real      (myFFT_1_sdata_out_payload_27_real[15:0]   ), //o
    .sdata_out_payload_27_imag      (myFFT_1_sdata_out_payload_27_imag[15:0]   ), //o
    .sdata_out_payload_28_real      (myFFT_1_sdata_out_payload_28_real[15:0]   ), //o
    .sdata_out_payload_28_imag      (myFFT_1_sdata_out_payload_28_imag[15:0]   ), //o
    .sdata_out_payload_29_real      (myFFT_1_sdata_out_payload_29_real[15:0]   ), //o
    .sdata_out_payload_29_imag      (myFFT_1_sdata_out_payload_29_imag[15:0]   ), //o
    .sdata_out_payload_30_real      (myFFT_1_sdata_out_payload_30_real[15:0]   ), //o
    .sdata_out_payload_30_imag      (myFFT_1_sdata_out_payload_30_imag[15:0]   ), //o
    .sdata_out_payload_31_real      (myFFT_1_sdata_out_payload_31_real[15:0]   ), //o
    .sdata_out_payload_31_imag      (myFFT_1_sdata_out_payload_31_imag[15:0]   ), //o
    .sdata_out_payload_32_real      (myFFT_1_sdata_out_payload_32_real[15:0]   ), //o
    .sdata_out_payload_32_imag      (myFFT_1_sdata_out_payload_32_imag[15:0]   ), //o
    .sdata_out_payload_33_real      (myFFT_1_sdata_out_payload_33_real[15:0]   ), //o
    .sdata_out_payload_33_imag      (myFFT_1_sdata_out_payload_33_imag[15:0]   ), //o
    .sdata_out_payload_34_real      (myFFT_1_sdata_out_payload_34_real[15:0]   ), //o
    .sdata_out_payload_34_imag      (myFFT_1_sdata_out_payload_34_imag[15:0]   ), //o
    .sdata_out_payload_35_real      (myFFT_1_sdata_out_payload_35_real[15:0]   ), //o
    .sdata_out_payload_35_imag      (myFFT_1_sdata_out_payload_35_imag[15:0]   ), //o
    .sdata_out_payload_36_real      (myFFT_1_sdata_out_payload_36_real[15:0]   ), //o
    .sdata_out_payload_36_imag      (myFFT_1_sdata_out_payload_36_imag[15:0]   ), //o
    .sdata_out_payload_37_real      (myFFT_1_sdata_out_payload_37_real[15:0]   ), //o
    .sdata_out_payload_37_imag      (myFFT_1_sdata_out_payload_37_imag[15:0]   ), //o
    .sdata_out_payload_38_real      (myFFT_1_sdata_out_payload_38_real[15:0]   ), //o
    .sdata_out_payload_38_imag      (myFFT_1_sdata_out_payload_38_imag[15:0]   ), //o
    .sdata_out_payload_39_real      (myFFT_1_sdata_out_payload_39_real[15:0]   ), //o
    .sdata_out_payload_39_imag      (myFFT_1_sdata_out_payload_39_imag[15:0]   ), //o
    .sdata_out_payload_40_real      (myFFT_1_sdata_out_payload_40_real[15:0]   ), //o
    .sdata_out_payload_40_imag      (myFFT_1_sdata_out_payload_40_imag[15:0]   ), //o
    .sdata_out_payload_41_real      (myFFT_1_sdata_out_payload_41_real[15:0]   ), //o
    .sdata_out_payload_41_imag      (myFFT_1_sdata_out_payload_41_imag[15:0]   ), //o
    .sdata_out_payload_42_real      (myFFT_1_sdata_out_payload_42_real[15:0]   ), //o
    .sdata_out_payload_42_imag      (myFFT_1_sdata_out_payload_42_imag[15:0]   ), //o
    .sdata_out_payload_43_real      (myFFT_1_sdata_out_payload_43_real[15:0]   ), //o
    .sdata_out_payload_43_imag      (myFFT_1_sdata_out_payload_43_imag[15:0]   ), //o
    .sdata_out_payload_44_real      (myFFT_1_sdata_out_payload_44_real[15:0]   ), //o
    .sdata_out_payload_44_imag      (myFFT_1_sdata_out_payload_44_imag[15:0]   ), //o
    .sdata_out_payload_45_real      (myFFT_1_sdata_out_payload_45_real[15:0]   ), //o
    .sdata_out_payload_45_imag      (myFFT_1_sdata_out_payload_45_imag[15:0]   ), //o
    .sdata_out_payload_46_real      (myFFT_1_sdata_out_payload_46_real[15:0]   ), //o
    .sdata_out_payload_46_imag      (myFFT_1_sdata_out_payload_46_imag[15:0]   ), //o
    .sdata_out_payload_47_real      (myFFT_1_sdata_out_payload_47_real[15:0]   ), //o
    .sdata_out_payload_47_imag      (myFFT_1_sdata_out_payload_47_imag[15:0]   ), //o
    .sdata_out_payload_48_real      (myFFT_1_sdata_out_payload_48_real[15:0]   ), //o
    .sdata_out_payload_48_imag      (myFFT_1_sdata_out_payload_48_imag[15:0]   ), //o
    .sdata_out_payload_49_real      (myFFT_1_sdata_out_payload_49_real[15:0]   ), //o
    .sdata_out_payload_49_imag      (myFFT_1_sdata_out_payload_49_imag[15:0]   ), //o
    .sdata_out_payload_50_real      (myFFT_1_sdata_out_payload_50_real[15:0]   ), //o
    .sdata_out_payload_50_imag      (myFFT_1_sdata_out_payload_50_imag[15:0]   ), //o
    .sdata_out_payload_51_real      (myFFT_1_sdata_out_payload_51_real[15:0]   ), //o
    .sdata_out_payload_51_imag      (myFFT_1_sdata_out_payload_51_imag[15:0]   ), //o
    .sdata_out_payload_52_real      (myFFT_1_sdata_out_payload_52_real[15:0]   ), //o
    .sdata_out_payload_52_imag      (myFFT_1_sdata_out_payload_52_imag[15:0]   ), //o
    .sdata_out_payload_53_real      (myFFT_1_sdata_out_payload_53_real[15:0]   ), //o
    .sdata_out_payload_53_imag      (myFFT_1_sdata_out_payload_53_imag[15:0]   ), //o
    .sdata_out_payload_54_real      (myFFT_1_sdata_out_payload_54_real[15:0]   ), //o
    .sdata_out_payload_54_imag      (myFFT_1_sdata_out_payload_54_imag[15:0]   ), //o
    .sdata_out_payload_55_real      (myFFT_1_sdata_out_payload_55_real[15:0]   ), //o
    .sdata_out_payload_55_imag      (myFFT_1_sdata_out_payload_55_imag[15:0]   ), //o
    .sdata_out_payload_56_real      (myFFT_1_sdata_out_payload_56_real[15:0]   ), //o
    .sdata_out_payload_56_imag      (myFFT_1_sdata_out_payload_56_imag[15:0]   ), //o
    .sdata_out_payload_57_real      (myFFT_1_sdata_out_payload_57_real[15:0]   ), //o
    .sdata_out_payload_57_imag      (myFFT_1_sdata_out_payload_57_imag[15:0]   ), //o
    .sdata_out_payload_58_real      (myFFT_1_sdata_out_payload_58_real[15:0]   ), //o
    .sdata_out_payload_58_imag      (myFFT_1_sdata_out_payload_58_imag[15:0]   ), //o
    .sdata_out_payload_59_real      (myFFT_1_sdata_out_payload_59_real[15:0]   ), //o
    .sdata_out_payload_59_imag      (myFFT_1_sdata_out_payload_59_imag[15:0]   ), //o
    .sdata_out_payload_60_real      (myFFT_1_sdata_out_payload_60_real[15:0]   ), //o
    .sdata_out_payload_60_imag      (myFFT_1_sdata_out_payload_60_imag[15:0]   ), //o
    .sdata_out_payload_61_real      (myFFT_1_sdata_out_payload_61_real[15:0]   ), //o
    .sdata_out_payload_61_imag      (myFFT_1_sdata_out_payload_61_imag[15:0]   ), //o
    .sdata_out_payload_62_real      (myFFT_1_sdata_out_payload_62_real[15:0]   ), //o
    .sdata_out_payload_62_imag      (myFFT_1_sdata_out_payload_62_imag[15:0]   ), //o
    .sdata_out_payload_63_real      (myFFT_1_sdata_out_payload_63_real[15:0]   ), //o
    .sdata_out_payload_63_imag      (myFFT_1_sdata_out_payload_63_imag[15:0]   ), //o
    .sdata_out_payload_64_real      (myFFT_1_sdata_out_payload_64_real[15:0]   ), //o
    .sdata_out_payload_64_imag      (myFFT_1_sdata_out_payload_64_imag[15:0]   ), //o
    .sdata_out_payload_65_real      (myFFT_1_sdata_out_payload_65_real[15:0]   ), //o
    .sdata_out_payload_65_imag      (myFFT_1_sdata_out_payload_65_imag[15:0]   ), //o
    .sdata_out_payload_66_real      (myFFT_1_sdata_out_payload_66_real[15:0]   ), //o
    .sdata_out_payload_66_imag      (myFFT_1_sdata_out_payload_66_imag[15:0]   ), //o
    .sdata_out_payload_67_real      (myFFT_1_sdata_out_payload_67_real[15:0]   ), //o
    .sdata_out_payload_67_imag      (myFFT_1_sdata_out_payload_67_imag[15:0]   ), //o
    .sdata_out_payload_68_real      (myFFT_1_sdata_out_payload_68_real[15:0]   ), //o
    .sdata_out_payload_68_imag      (myFFT_1_sdata_out_payload_68_imag[15:0]   ), //o
    .sdata_out_payload_69_real      (myFFT_1_sdata_out_payload_69_real[15:0]   ), //o
    .sdata_out_payload_69_imag      (myFFT_1_sdata_out_payload_69_imag[15:0]   ), //o
    .sdata_out_payload_70_real      (myFFT_1_sdata_out_payload_70_real[15:0]   ), //o
    .sdata_out_payload_70_imag      (myFFT_1_sdata_out_payload_70_imag[15:0]   ), //o
    .sdata_out_payload_71_real      (myFFT_1_sdata_out_payload_71_real[15:0]   ), //o
    .sdata_out_payload_71_imag      (myFFT_1_sdata_out_payload_71_imag[15:0]   ), //o
    .sdata_out_payload_72_real      (myFFT_1_sdata_out_payload_72_real[15:0]   ), //o
    .sdata_out_payload_72_imag      (myFFT_1_sdata_out_payload_72_imag[15:0]   ), //o
    .sdata_out_payload_73_real      (myFFT_1_sdata_out_payload_73_real[15:0]   ), //o
    .sdata_out_payload_73_imag      (myFFT_1_sdata_out_payload_73_imag[15:0]   ), //o
    .sdata_out_payload_74_real      (myFFT_1_sdata_out_payload_74_real[15:0]   ), //o
    .sdata_out_payload_74_imag      (myFFT_1_sdata_out_payload_74_imag[15:0]   ), //o
    .sdata_out_payload_75_real      (myFFT_1_sdata_out_payload_75_real[15:0]   ), //o
    .sdata_out_payload_75_imag      (myFFT_1_sdata_out_payload_75_imag[15:0]   ), //o
    .sdata_out_payload_76_real      (myFFT_1_sdata_out_payload_76_real[15:0]   ), //o
    .sdata_out_payload_76_imag      (myFFT_1_sdata_out_payload_76_imag[15:0]   ), //o
    .sdata_out_payload_77_real      (myFFT_1_sdata_out_payload_77_real[15:0]   ), //o
    .sdata_out_payload_77_imag      (myFFT_1_sdata_out_payload_77_imag[15:0]   ), //o
    .sdata_out_payload_78_real      (myFFT_1_sdata_out_payload_78_real[15:0]   ), //o
    .sdata_out_payload_78_imag      (myFFT_1_sdata_out_payload_78_imag[15:0]   ), //o
    .sdata_out_payload_79_real      (myFFT_1_sdata_out_payload_79_real[15:0]   ), //o
    .sdata_out_payload_79_imag      (myFFT_1_sdata_out_payload_79_imag[15:0]   ), //o
    .sdata_out_payload_80_real      (myFFT_1_sdata_out_payload_80_real[15:0]   ), //o
    .sdata_out_payload_80_imag      (myFFT_1_sdata_out_payload_80_imag[15:0]   ), //o
    .sdata_out_payload_81_real      (myFFT_1_sdata_out_payload_81_real[15:0]   ), //o
    .sdata_out_payload_81_imag      (myFFT_1_sdata_out_payload_81_imag[15:0]   ), //o
    .sdata_out_payload_82_real      (myFFT_1_sdata_out_payload_82_real[15:0]   ), //o
    .sdata_out_payload_82_imag      (myFFT_1_sdata_out_payload_82_imag[15:0]   ), //o
    .sdata_out_payload_83_real      (myFFT_1_sdata_out_payload_83_real[15:0]   ), //o
    .sdata_out_payload_83_imag      (myFFT_1_sdata_out_payload_83_imag[15:0]   ), //o
    .sdata_out_payload_84_real      (myFFT_1_sdata_out_payload_84_real[15:0]   ), //o
    .sdata_out_payload_84_imag      (myFFT_1_sdata_out_payload_84_imag[15:0]   ), //o
    .sdata_out_payload_85_real      (myFFT_1_sdata_out_payload_85_real[15:0]   ), //o
    .sdata_out_payload_85_imag      (myFFT_1_sdata_out_payload_85_imag[15:0]   ), //o
    .sdata_out_payload_86_real      (myFFT_1_sdata_out_payload_86_real[15:0]   ), //o
    .sdata_out_payload_86_imag      (myFFT_1_sdata_out_payload_86_imag[15:0]   ), //o
    .sdata_out_payload_87_real      (myFFT_1_sdata_out_payload_87_real[15:0]   ), //o
    .sdata_out_payload_87_imag      (myFFT_1_sdata_out_payload_87_imag[15:0]   ), //o
    .sdata_out_payload_88_real      (myFFT_1_sdata_out_payload_88_real[15:0]   ), //o
    .sdata_out_payload_88_imag      (myFFT_1_sdata_out_payload_88_imag[15:0]   ), //o
    .sdata_out_payload_89_real      (myFFT_1_sdata_out_payload_89_real[15:0]   ), //o
    .sdata_out_payload_89_imag      (myFFT_1_sdata_out_payload_89_imag[15:0]   ), //o
    .sdata_out_payload_90_real      (myFFT_1_sdata_out_payload_90_real[15:0]   ), //o
    .sdata_out_payload_90_imag      (myFFT_1_sdata_out_payload_90_imag[15:0]   ), //o
    .sdata_out_payload_91_real      (myFFT_1_sdata_out_payload_91_real[15:0]   ), //o
    .sdata_out_payload_91_imag      (myFFT_1_sdata_out_payload_91_imag[15:0]   ), //o
    .sdata_out_payload_92_real      (myFFT_1_sdata_out_payload_92_real[15:0]   ), //o
    .sdata_out_payload_92_imag      (myFFT_1_sdata_out_payload_92_imag[15:0]   ), //o
    .sdata_out_payload_93_real      (myFFT_1_sdata_out_payload_93_real[15:0]   ), //o
    .sdata_out_payload_93_imag      (myFFT_1_sdata_out_payload_93_imag[15:0]   ), //o
    .sdata_out_payload_94_real      (myFFT_1_sdata_out_payload_94_real[15:0]   ), //o
    .sdata_out_payload_94_imag      (myFFT_1_sdata_out_payload_94_imag[15:0]   ), //o
    .sdata_out_payload_95_real      (myFFT_1_sdata_out_payload_95_real[15:0]   ), //o
    .sdata_out_payload_95_imag      (myFFT_1_sdata_out_payload_95_imag[15:0]   ), //o
    .sdata_out_payload_96_real      (myFFT_1_sdata_out_payload_96_real[15:0]   ), //o
    .sdata_out_payload_96_imag      (myFFT_1_sdata_out_payload_96_imag[15:0]   ), //o
    .sdata_out_payload_97_real      (myFFT_1_sdata_out_payload_97_real[15:0]   ), //o
    .sdata_out_payload_97_imag      (myFFT_1_sdata_out_payload_97_imag[15:0]   ), //o
    .sdata_out_payload_98_real      (myFFT_1_sdata_out_payload_98_real[15:0]   ), //o
    .sdata_out_payload_98_imag      (myFFT_1_sdata_out_payload_98_imag[15:0]   ), //o
    .sdata_out_payload_99_real      (myFFT_1_sdata_out_payload_99_real[15:0]   ), //o
    .sdata_out_payload_99_imag      (myFFT_1_sdata_out_payload_99_imag[15:0]   ), //o
    .sdata_out_payload_100_real     (myFFT_1_sdata_out_payload_100_real[15:0]  ), //o
    .sdata_out_payload_100_imag     (myFFT_1_sdata_out_payload_100_imag[15:0]  ), //o
    .sdata_out_payload_101_real     (myFFT_1_sdata_out_payload_101_real[15:0]  ), //o
    .sdata_out_payload_101_imag     (myFFT_1_sdata_out_payload_101_imag[15:0]  ), //o
    .sdata_out_payload_102_real     (myFFT_1_sdata_out_payload_102_real[15:0]  ), //o
    .sdata_out_payload_102_imag     (myFFT_1_sdata_out_payload_102_imag[15:0]  ), //o
    .sdata_out_payload_103_real     (myFFT_1_sdata_out_payload_103_real[15:0]  ), //o
    .sdata_out_payload_103_imag     (myFFT_1_sdata_out_payload_103_imag[15:0]  ), //o
    .sdata_out_payload_104_real     (myFFT_1_sdata_out_payload_104_real[15:0]  ), //o
    .sdata_out_payload_104_imag     (myFFT_1_sdata_out_payload_104_imag[15:0]  ), //o
    .sdata_out_payload_105_real     (myFFT_1_sdata_out_payload_105_real[15:0]  ), //o
    .sdata_out_payload_105_imag     (myFFT_1_sdata_out_payload_105_imag[15:0]  ), //o
    .sdata_out_payload_106_real     (myFFT_1_sdata_out_payload_106_real[15:0]  ), //o
    .sdata_out_payload_106_imag     (myFFT_1_sdata_out_payload_106_imag[15:0]  ), //o
    .sdata_out_payload_107_real     (myFFT_1_sdata_out_payload_107_real[15:0]  ), //o
    .sdata_out_payload_107_imag     (myFFT_1_sdata_out_payload_107_imag[15:0]  ), //o
    .sdata_out_payload_108_real     (myFFT_1_sdata_out_payload_108_real[15:0]  ), //o
    .sdata_out_payload_108_imag     (myFFT_1_sdata_out_payload_108_imag[15:0]  ), //o
    .sdata_out_payload_109_real     (myFFT_1_sdata_out_payload_109_real[15:0]  ), //o
    .sdata_out_payload_109_imag     (myFFT_1_sdata_out_payload_109_imag[15:0]  ), //o
    .sdata_out_payload_110_real     (myFFT_1_sdata_out_payload_110_real[15:0]  ), //o
    .sdata_out_payload_110_imag     (myFFT_1_sdata_out_payload_110_imag[15:0]  ), //o
    .sdata_out_payload_111_real     (myFFT_1_sdata_out_payload_111_real[15:0]  ), //o
    .sdata_out_payload_111_imag     (myFFT_1_sdata_out_payload_111_imag[15:0]  ), //o
    .sdata_out_payload_112_real     (myFFT_1_sdata_out_payload_112_real[15:0]  ), //o
    .sdata_out_payload_112_imag     (myFFT_1_sdata_out_payload_112_imag[15:0]  ), //o
    .sdata_out_payload_113_real     (myFFT_1_sdata_out_payload_113_real[15:0]  ), //o
    .sdata_out_payload_113_imag     (myFFT_1_sdata_out_payload_113_imag[15:0]  ), //o
    .sdata_out_payload_114_real     (myFFT_1_sdata_out_payload_114_real[15:0]  ), //o
    .sdata_out_payload_114_imag     (myFFT_1_sdata_out_payload_114_imag[15:0]  ), //o
    .sdata_out_payload_115_real     (myFFT_1_sdata_out_payload_115_real[15:0]  ), //o
    .sdata_out_payload_115_imag     (myFFT_1_sdata_out_payload_115_imag[15:0]  ), //o
    .sdata_out_payload_116_real     (myFFT_1_sdata_out_payload_116_real[15:0]  ), //o
    .sdata_out_payload_116_imag     (myFFT_1_sdata_out_payload_116_imag[15:0]  ), //o
    .sdata_out_payload_117_real     (myFFT_1_sdata_out_payload_117_real[15:0]  ), //o
    .sdata_out_payload_117_imag     (myFFT_1_sdata_out_payload_117_imag[15:0]  ), //o
    .sdata_out_payload_118_real     (myFFT_1_sdata_out_payload_118_real[15:0]  ), //o
    .sdata_out_payload_118_imag     (myFFT_1_sdata_out_payload_118_imag[15:0]  ), //o
    .sdata_out_payload_119_real     (myFFT_1_sdata_out_payload_119_real[15:0]  ), //o
    .sdata_out_payload_119_imag     (myFFT_1_sdata_out_payload_119_imag[15:0]  ), //o
    .sdata_out_payload_120_real     (myFFT_1_sdata_out_payload_120_real[15:0]  ), //o
    .sdata_out_payload_120_imag     (myFFT_1_sdata_out_payload_120_imag[15:0]  ), //o
    .sdata_out_payload_121_real     (myFFT_1_sdata_out_payload_121_real[15:0]  ), //o
    .sdata_out_payload_121_imag     (myFFT_1_sdata_out_payload_121_imag[15:0]  ), //o
    .sdata_out_payload_122_real     (myFFT_1_sdata_out_payload_122_real[15:0]  ), //o
    .sdata_out_payload_122_imag     (myFFT_1_sdata_out_payload_122_imag[15:0]  ), //o
    .sdata_out_payload_123_real     (myFFT_1_sdata_out_payload_123_real[15:0]  ), //o
    .sdata_out_payload_123_imag     (myFFT_1_sdata_out_payload_123_imag[15:0]  ), //o
    .sdata_out_payload_124_real     (myFFT_1_sdata_out_payload_124_real[15:0]  ), //o
    .sdata_out_payload_124_imag     (myFFT_1_sdata_out_payload_124_imag[15:0]  ), //o
    .sdata_out_payload_125_real     (myFFT_1_sdata_out_payload_125_real[15:0]  ), //o
    .sdata_out_payload_125_imag     (myFFT_1_sdata_out_payload_125_imag[15:0]  ), //o
    .sdata_out_payload_126_real     (myFFT_1_sdata_out_payload_126_real[15:0]  ), //o
    .sdata_out_payload_126_imag     (myFFT_1_sdata_out_payload_126_imag[15:0]  ), //o
    .sdata_out_payload_127_real     (myFFT_1_sdata_out_payload_127_real[15:0]  ), //o
    .sdata_out_payload_127_imag     (myFFT_1_sdata_out_payload_127_imag[15:0]  ), //o
    .clk                            (clk                                       ), //i
    .reset                          (reset                                     )  //i
  );
  always @(*) begin
    case(null_cnt_value)
      7'b0000000 : begin
        _zz_257 = sdata_out_regs_0_real;
        _zz_258 = sdata_out_regs_0_imag;
      end
      7'b0000001 : begin
        _zz_257 = sdata_out_regs_1_real;
        _zz_258 = sdata_out_regs_1_imag;
      end
      7'b0000010 : begin
        _zz_257 = sdata_out_regs_2_real;
        _zz_258 = sdata_out_regs_2_imag;
      end
      7'b0000011 : begin
        _zz_257 = sdata_out_regs_3_real;
        _zz_258 = sdata_out_regs_3_imag;
      end
      7'b0000100 : begin
        _zz_257 = sdata_out_regs_4_real;
        _zz_258 = sdata_out_regs_4_imag;
      end
      7'b0000101 : begin
        _zz_257 = sdata_out_regs_5_real;
        _zz_258 = sdata_out_regs_5_imag;
      end
      7'b0000110 : begin
        _zz_257 = sdata_out_regs_6_real;
        _zz_258 = sdata_out_regs_6_imag;
      end
      7'b0000111 : begin
        _zz_257 = sdata_out_regs_7_real;
        _zz_258 = sdata_out_regs_7_imag;
      end
      7'b0001000 : begin
        _zz_257 = sdata_out_regs_8_real;
        _zz_258 = sdata_out_regs_8_imag;
      end
      7'b0001001 : begin
        _zz_257 = sdata_out_regs_9_real;
        _zz_258 = sdata_out_regs_9_imag;
      end
      7'b0001010 : begin
        _zz_257 = sdata_out_regs_10_real;
        _zz_258 = sdata_out_regs_10_imag;
      end
      7'b0001011 : begin
        _zz_257 = sdata_out_regs_11_real;
        _zz_258 = sdata_out_regs_11_imag;
      end
      7'b0001100 : begin
        _zz_257 = sdata_out_regs_12_real;
        _zz_258 = sdata_out_regs_12_imag;
      end
      7'b0001101 : begin
        _zz_257 = sdata_out_regs_13_real;
        _zz_258 = sdata_out_regs_13_imag;
      end
      7'b0001110 : begin
        _zz_257 = sdata_out_regs_14_real;
        _zz_258 = sdata_out_regs_14_imag;
      end
      7'b0001111 : begin
        _zz_257 = sdata_out_regs_15_real;
        _zz_258 = sdata_out_regs_15_imag;
      end
      7'b0010000 : begin
        _zz_257 = sdata_out_regs_16_real;
        _zz_258 = sdata_out_regs_16_imag;
      end
      7'b0010001 : begin
        _zz_257 = sdata_out_regs_17_real;
        _zz_258 = sdata_out_regs_17_imag;
      end
      7'b0010010 : begin
        _zz_257 = sdata_out_regs_18_real;
        _zz_258 = sdata_out_regs_18_imag;
      end
      7'b0010011 : begin
        _zz_257 = sdata_out_regs_19_real;
        _zz_258 = sdata_out_regs_19_imag;
      end
      7'b0010100 : begin
        _zz_257 = sdata_out_regs_20_real;
        _zz_258 = sdata_out_regs_20_imag;
      end
      7'b0010101 : begin
        _zz_257 = sdata_out_regs_21_real;
        _zz_258 = sdata_out_regs_21_imag;
      end
      7'b0010110 : begin
        _zz_257 = sdata_out_regs_22_real;
        _zz_258 = sdata_out_regs_22_imag;
      end
      7'b0010111 : begin
        _zz_257 = sdata_out_regs_23_real;
        _zz_258 = sdata_out_regs_23_imag;
      end
      7'b0011000 : begin
        _zz_257 = sdata_out_regs_24_real;
        _zz_258 = sdata_out_regs_24_imag;
      end
      7'b0011001 : begin
        _zz_257 = sdata_out_regs_25_real;
        _zz_258 = sdata_out_regs_25_imag;
      end
      7'b0011010 : begin
        _zz_257 = sdata_out_regs_26_real;
        _zz_258 = sdata_out_regs_26_imag;
      end
      7'b0011011 : begin
        _zz_257 = sdata_out_regs_27_real;
        _zz_258 = sdata_out_regs_27_imag;
      end
      7'b0011100 : begin
        _zz_257 = sdata_out_regs_28_real;
        _zz_258 = sdata_out_regs_28_imag;
      end
      7'b0011101 : begin
        _zz_257 = sdata_out_regs_29_real;
        _zz_258 = sdata_out_regs_29_imag;
      end
      7'b0011110 : begin
        _zz_257 = sdata_out_regs_30_real;
        _zz_258 = sdata_out_regs_30_imag;
      end
      7'b0011111 : begin
        _zz_257 = sdata_out_regs_31_real;
        _zz_258 = sdata_out_regs_31_imag;
      end
      7'b0100000 : begin
        _zz_257 = sdata_out_regs_32_real;
        _zz_258 = sdata_out_regs_32_imag;
      end
      7'b0100001 : begin
        _zz_257 = sdata_out_regs_33_real;
        _zz_258 = sdata_out_regs_33_imag;
      end
      7'b0100010 : begin
        _zz_257 = sdata_out_regs_34_real;
        _zz_258 = sdata_out_regs_34_imag;
      end
      7'b0100011 : begin
        _zz_257 = sdata_out_regs_35_real;
        _zz_258 = sdata_out_regs_35_imag;
      end
      7'b0100100 : begin
        _zz_257 = sdata_out_regs_36_real;
        _zz_258 = sdata_out_regs_36_imag;
      end
      7'b0100101 : begin
        _zz_257 = sdata_out_regs_37_real;
        _zz_258 = sdata_out_regs_37_imag;
      end
      7'b0100110 : begin
        _zz_257 = sdata_out_regs_38_real;
        _zz_258 = sdata_out_regs_38_imag;
      end
      7'b0100111 : begin
        _zz_257 = sdata_out_regs_39_real;
        _zz_258 = sdata_out_regs_39_imag;
      end
      7'b0101000 : begin
        _zz_257 = sdata_out_regs_40_real;
        _zz_258 = sdata_out_regs_40_imag;
      end
      7'b0101001 : begin
        _zz_257 = sdata_out_regs_41_real;
        _zz_258 = sdata_out_regs_41_imag;
      end
      7'b0101010 : begin
        _zz_257 = sdata_out_regs_42_real;
        _zz_258 = sdata_out_regs_42_imag;
      end
      7'b0101011 : begin
        _zz_257 = sdata_out_regs_43_real;
        _zz_258 = sdata_out_regs_43_imag;
      end
      7'b0101100 : begin
        _zz_257 = sdata_out_regs_44_real;
        _zz_258 = sdata_out_regs_44_imag;
      end
      7'b0101101 : begin
        _zz_257 = sdata_out_regs_45_real;
        _zz_258 = sdata_out_regs_45_imag;
      end
      7'b0101110 : begin
        _zz_257 = sdata_out_regs_46_real;
        _zz_258 = sdata_out_regs_46_imag;
      end
      7'b0101111 : begin
        _zz_257 = sdata_out_regs_47_real;
        _zz_258 = sdata_out_regs_47_imag;
      end
      7'b0110000 : begin
        _zz_257 = sdata_out_regs_48_real;
        _zz_258 = sdata_out_regs_48_imag;
      end
      7'b0110001 : begin
        _zz_257 = sdata_out_regs_49_real;
        _zz_258 = sdata_out_regs_49_imag;
      end
      7'b0110010 : begin
        _zz_257 = sdata_out_regs_50_real;
        _zz_258 = sdata_out_regs_50_imag;
      end
      7'b0110011 : begin
        _zz_257 = sdata_out_regs_51_real;
        _zz_258 = sdata_out_regs_51_imag;
      end
      7'b0110100 : begin
        _zz_257 = sdata_out_regs_52_real;
        _zz_258 = sdata_out_regs_52_imag;
      end
      7'b0110101 : begin
        _zz_257 = sdata_out_regs_53_real;
        _zz_258 = sdata_out_regs_53_imag;
      end
      7'b0110110 : begin
        _zz_257 = sdata_out_regs_54_real;
        _zz_258 = sdata_out_regs_54_imag;
      end
      7'b0110111 : begin
        _zz_257 = sdata_out_regs_55_real;
        _zz_258 = sdata_out_regs_55_imag;
      end
      7'b0111000 : begin
        _zz_257 = sdata_out_regs_56_real;
        _zz_258 = sdata_out_regs_56_imag;
      end
      7'b0111001 : begin
        _zz_257 = sdata_out_regs_57_real;
        _zz_258 = sdata_out_regs_57_imag;
      end
      7'b0111010 : begin
        _zz_257 = sdata_out_regs_58_real;
        _zz_258 = sdata_out_regs_58_imag;
      end
      7'b0111011 : begin
        _zz_257 = sdata_out_regs_59_real;
        _zz_258 = sdata_out_regs_59_imag;
      end
      7'b0111100 : begin
        _zz_257 = sdata_out_regs_60_real;
        _zz_258 = sdata_out_regs_60_imag;
      end
      7'b0111101 : begin
        _zz_257 = sdata_out_regs_61_real;
        _zz_258 = sdata_out_regs_61_imag;
      end
      7'b0111110 : begin
        _zz_257 = sdata_out_regs_62_real;
        _zz_258 = sdata_out_regs_62_imag;
      end
      7'b0111111 : begin
        _zz_257 = sdata_out_regs_63_real;
        _zz_258 = sdata_out_regs_63_imag;
      end
      7'b1000000 : begin
        _zz_257 = sdata_out_regs_64_real;
        _zz_258 = sdata_out_regs_64_imag;
      end
      7'b1000001 : begin
        _zz_257 = sdata_out_regs_65_real;
        _zz_258 = sdata_out_regs_65_imag;
      end
      7'b1000010 : begin
        _zz_257 = sdata_out_regs_66_real;
        _zz_258 = sdata_out_regs_66_imag;
      end
      7'b1000011 : begin
        _zz_257 = sdata_out_regs_67_real;
        _zz_258 = sdata_out_regs_67_imag;
      end
      7'b1000100 : begin
        _zz_257 = sdata_out_regs_68_real;
        _zz_258 = sdata_out_regs_68_imag;
      end
      7'b1000101 : begin
        _zz_257 = sdata_out_regs_69_real;
        _zz_258 = sdata_out_regs_69_imag;
      end
      7'b1000110 : begin
        _zz_257 = sdata_out_regs_70_real;
        _zz_258 = sdata_out_regs_70_imag;
      end
      7'b1000111 : begin
        _zz_257 = sdata_out_regs_71_real;
        _zz_258 = sdata_out_regs_71_imag;
      end
      7'b1001000 : begin
        _zz_257 = sdata_out_regs_72_real;
        _zz_258 = sdata_out_regs_72_imag;
      end
      7'b1001001 : begin
        _zz_257 = sdata_out_regs_73_real;
        _zz_258 = sdata_out_regs_73_imag;
      end
      7'b1001010 : begin
        _zz_257 = sdata_out_regs_74_real;
        _zz_258 = sdata_out_regs_74_imag;
      end
      7'b1001011 : begin
        _zz_257 = sdata_out_regs_75_real;
        _zz_258 = sdata_out_regs_75_imag;
      end
      7'b1001100 : begin
        _zz_257 = sdata_out_regs_76_real;
        _zz_258 = sdata_out_regs_76_imag;
      end
      7'b1001101 : begin
        _zz_257 = sdata_out_regs_77_real;
        _zz_258 = sdata_out_regs_77_imag;
      end
      7'b1001110 : begin
        _zz_257 = sdata_out_regs_78_real;
        _zz_258 = sdata_out_regs_78_imag;
      end
      7'b1001111 : begin
        _zz_257 = sdata_out_regs_79_real;
        _zz_258 = sdata_out_regs_79_imag;
      end
      7'b1010000 : begin
        _zz_257 = sdata_out_regs_80_real;
        _zz_258 = sdata_out_regs_80_imag;
      end
      7'b1010001 : begin
        _zz_257 = sdata_out_regs_81_real;
        _zz_258 = sdata_out_regs_81_imag;
      end
      7'b1010010 : begin
        _zz_257 = sdata_out_regs_82_real;
        _zz_258 = sdata_out_regs_82_imag;
      end
      7'b1010011 : begin
        _zz_257 = sdata_out_regs_83_real;
        _zz_258 = sdata_out_regs_83_imag;
      end
      7'b1010100 : begin
        _zz_257 = sdata_out_regs_84_real;
        _zz_258 = sdata_out_regs_84_imag;
      end
      7'b1010101 : begin
        _zz_257 = sdata_out_regs_85_real;
        _zz_258 = sdata_out_regs_85_imag;
      end
      7'b1010110 : begin
        _zz_257 = sdata_out_regs_86_real;
        _zz_258 = sdata_out_regs_86_imag;
      end
      7'b1010111 : begin
        _zz_257 = sdata_out_regs_87_real;
        _zz_258 = sdata_out_regs_87_imag;
      end
      7'b1011000 : begin
        _zz_257 = sdata_out_regs_88_real;
        _zz_258 = sdata_out_regs_88_imag;
      end
      7'b1011001 : begin
        _zz_257 = sdata_out_regs_89_real;
        _zz_258 = sdata_out_regs_89_imag;
      end
      7'b1011010 : begin
        _zz_257 = sdata_out_regs_90_real;
        _zz_258 = sdata_out_regs_90_imag;
      end
      7'b1011011 : begin
        _zz_257 = sdata_out_regs_91_real;
        _zz_258 = sdata_out_regs_91_imag;
      end
      7'b1011100 : begin
        _zz_257 = sdata_out_regs_92_real;
        _zz_258 = sdata_out_regs_92_imag;
      end
      7'b1011101 : begin
        _zz_257 = sdata_out_regs_93_real;
        _zz_258 = sdata_out_regs_93_imag;
      end
      7'b1011110 : begin
        _zz_257 = sdata_out_regs_94_real;
        _zz_258 = sdata_out_regs_94_imag;
      end
      7'b1011111 : begin
        _zz_257 = sdata_out_regs_95_real;
        _zz_258 = sdata_out_regs_95_imag;
      end
      7'b1100000 : begin
        _zz_257 = sdata_out_regs_96_real;
        _zz_258 = sdata_out_regs_96_imag;
      end
      7'b1100001 : begin
        _zz_257 = sdata_out_regs_97_real;
        _zz_258 = sdata_out_regs_97_imag;
      end
      7'b1100010 : begin
        _zz_257 = sdata_out_regs_98_real;
        _zz_258 = sdata_out_regs_98_imag;
      end
      7'b1100011 : begin
        _zz_257 = sdata_out_regs_99_real;
        _zz_258 = sdata_out_regs_99_imag;
      end
      7'b1100100 : begin
        _zz_257 = sdata_out_regs_100_real;
        _zz_258 = sdata_out_regs_100_imag;
      end
      7'b1100101 : begin
        _zz_257 = sdata_out_regs_101_real;
        _zz_258 = sdata_out_regs_101_imag;
      end
      7'b1100110 : begin
        _zz_257 = sdata_out_regs_102_real;
        _zz_258 = sdata_out_regs_102_imag;
      end
      7'b1100111 : begin
        _zz_257 = sdata_out_regs_103_real;
        _zz_258 = sdata_out_regs_103_imag;
      end
      7'b1101000 : begin
        _zz_257 = sdata_out_regs_104_real;
        _zz_258 = sdata_out_regs_104_imag;
      end
      7'b1101001 : begin
        _zz_257 = sdata_out_regs_105_real;
        _zz_258 = sdata_out_regs_105_imag;
      end
      7'b1101010 : begin
        _zz_257 = sdata_out_regs_106_real;
        _zz_258 = sdata_out_regs_106_imag;
      end
      7'b1101011 : begin
        _zz_257 = sdata_out_regs_107_real;
        _zz_258 = sdata_out_regs_107_imag;
      end
      7'b1101100 : begin
        _zz_257 = sdata_out_regs_108_real;
        _zz_258 = sdata_out_regs_108_imag;
      end
      7'b1101101 : begin
        _zz_257 = sdata_out_regs_109_real;
        _zz_258 = sdata_out_regs_109_imag;
      end
      7'b1101110 : begin
        _zz_257 = sdata_out_regs_110_real;
        _zz_258 = sdata_out_regs_110_imag;
      end
      7'b1101111 : begin
        _zz_257 = sdata_out_regs_111_real;
        _zz_258 = sdata_out_regs_111_imag;
      end
      7'b1110000 : begin
        _zz_257 = sdata_out_regs_112_real;
        _zz_258 = sdata_out_regs_112_imag;
      end
      7'b1110001 : begin
        _zz_257 = sdata_out_regs_113_real;
        _zz_258 = sdata_out_regs_113_imag;
      end
      7'b1110010 : begin
        _zz_257 = sdata_out_regs_114_real;
        _zz_258 = sdata_out_regs_114_imag;
      end
      7'b1110011 : begin
        _zz_257 = sdata_out_regs_115_real;
        _zz_258 = sdata_out_regs_115_imag;
      end
      7'b1110100 : begin
        _zz_257 = sdata_out_regs_116_real;
        _zz_258 = sdata_out_regs_116_imag;
      end
      7'b1110101 : begin
        _zz_257 = sdata_out_regs_117_real;
        _zz_258 = sdata_out_regs_117_imag;
      end
      7'b1110110 : begin
        _zz_257 = sdata_out_regs_118_real;
        _zz_258 = sdata_out_regs_118_imag;
      end
      7'b1110111 : begin
        _zz_257 = sdata_out_regs_119_real;
        _zz_258 = sdata_out_regs_119_imag;
      end
      7'b1111000 : begin
        _zz_257 = sdata_out_regs_120_real;
        _zz_258 = sdata_out_regs_120_imag;
      end
      7'b1111001 : begin
        _zz_257 = sdata_out_regs_121_real;
        _zz_258 = sdata_out_regs_121_imag;
      end
      7'b1111010 : begin
        _zz_257 = sdata_out_regs_122_real;
        _zz_258 = sdata_out_regs_122_imag;
      end
      7'b1111011 : begin
        _zz_257 = sdata_out_regs_123_real;
        _zz_258 = sdata_out_regs_123_imag;
      end
      7'b1111100 : begin
        _zz_257 = sdata_out_regs_124_real;
        _zz_258 = sdata_out_regs_124_imag;
      end
      7'b1111101 : begin
        _zz_257 = sdata_out_regs_125_real;
        _zz_258 = sdata_out_regs_125_imag;
      end
      7'b1111110 : begin
        _zz_257 = sdata_out_regs_126_real;
        _zz_258 = sdata_out_regs_126_imag;
      end
      default : begin
        _zz_257 = sdata_out_regs_127_real;
        _zz_258 = sdata_out_regs_127_imag;
      end
    endcase
  end

  assign _zz_1 = data_in_payload_real;
  assign _zz_2 = data_in_payload_imag;
  assign fft_input_flow_payload_0_real = _zz_255;
  assign fft_input_flow_payload_0_imag = _zz_256;
  assign fft_input_flow_payload_1_real = _zz_253;
  assign fft_input_flow_payload_1_imag = _zz_254;
  assign fft_input_flow_payload_2_real = _zz_251;
  assign fft_input_flow_payload_2_imag = _zz_252;
  assign fft_input_flow_payload_3_real = _zz_249;
  assign fft_input_flow_payload_3_imag = _zz_250;
  assign fft_input_flow_payload_4_real = _zz_247;
  assign fft_input_flow_payload_4_imag = _zz_248;
  assign fft_input_flow_payload_5_real = _zz_245;
  assign fft_input_flow_payload_5_imag = _zz_246;
  assign fft_input_flow_payload_6_real = _zz_243;
  assign fft_input_flow_payload_6_imag = _zz_244;
  assign fft_input_flow_payload_7_real = _zz_241;
  assign fft_input_flow_payload_7_imag = _zz_242;
  assign fft_input_flow_payload_8_real = _zz_239;
  assign fft_input_flow_payload_8_imag = _zz_240;
  assign fft_input_flow_payload_9_real = _zz_237;
  assign fft_input_flow_payload_9_imag = _zz_238;
  assign fft_input_flow_payload_10_real = _zz_235;
  assign fft_input_flow_payload_10_imag = _zz_236;
  assign fft_input_flow_payload_11_real = _zz_233;
  assign fft_input_flow_payload_11_imag = _zz_234;
  assign fft_input_flow_payload_12_real = _zz_231;
  assign fft_input_flow_payload_12_imag = _zz_232;
  assign fft_input_flow_payload_13_real = _zz_229;
  assign fft_input_flow_payload_13_imag = _zz_230;
  assign fft_input_flow_payload_14_real = _zz_227;
  assign fft_input_flow_payload_14_imag = _zz_228;
  assign fft_input_flow_payload_15_real = _zz_225;
  assign fft_input_flow_payload_15_imag = _zz_226;
  assign fft_input_flow_payload_16_real = _zz_223;
  assign fft_input_flow_payload_16_imag = _zz_224;
  assign fft_input_flow_payload_17_real = _zz_221;
  assign fft_input_flow_payload_17_imag = _zz_222;
  assign fft_input_flow_payload_18_real = _zz_219;
  assign fft_input_flow_payload_18_imag = _zz_220;
  assign fft_input_flow_payload_19_real = _zz_217;
  assign fft_input_flow_payload_19_imag = _zz_218;
  assign fft_input_flow_payload_20_real = _zz_215;
  assign fft_input_flow_payload_20_imag = _zz_216;
  assign fft_input_flow_payload_21_real = _zz_213;
  assign fft_input_flow_payload_21_imag = _zz_214;
  assign fft_input_flow_payload_22_real = _zz_211;
  assign fft_input_flow_payload_22_imag = _zz_212;
  assign fft_input_flow_payload_23_real = _zz_209;
  assign fft_input_flow_payload_23_imag = _zz_210;
  assign fft_input_flow_payload_24_real = _zz_207;
  assign fft_input_flow_payload_24_imag = _zz_208;
  assign fft_input_flow_payload_25_real = _zz_205;
  assign fft_input_flow_payload_25_imag = _zz_206;
  assign fft_input_flow_payload_26_real = _zz_203;
  assign fft_input_flow_payload_26_imag = _zz_204;
  assign fft_input_flow_payload_27_real = _zz_201;
  assign fft_input_flow_payload_27_imag = _zz_202;
  assign fft_input_flow_payload_28_real = _zz_199;
  assign fft_input_flow_payload_28_imag = _zz_200;
  assign fft_input_flow_payload_29_real = _zz_197;
  assign fft_input_flow_payload_29_imag = _zz_198;
  assign fft_input_flow_payload_30_real = _zz_195;
  assign fft_input_flow_payload_30_imag = _zz_196;
  assign fft_input_flow_payload_31_real = _zz_193;
  assign fft_input_flow_payload_31_imag = _zz_194;
  assign fft_input_flow_payload_32_real = _zz_191;
  assign fft_input_flow_payload_32_imag = _zz_192;
  assign fft_input_flow_payload_33_real = _zz_189;
  assign fft_input_flow_payload_33_imag = _zz_190;
  assign fft_input_flow_payload_34_real = _zz_187;
  assign fft_input_flow_payload_34_imag = _zz_188;
  assign fft_input_flow_payload_35_real = _zz_185;
  assign fft_input_flow_payload_35_imag = _zz_186;
  assign fft_input_flow_payload_36_real = _zz_183;
  assign fft_input_flow_payload_36_imag = _zz_184;
  assign fft_input_flow_payload_37_real = _zz_181;
  assign fft_input_flow_payload_37_imag = _zz_182;
  assign fft_input_flow_payload_38_real = _zz_179;
  assign fft_input_flow_payload_38_imag = _zz_180;
  assign fft_input_flow_payload_39_real = _zz_177;
  assign fft_input_flow_payload_39_imag = _zz_178;
  assign fft_input_flow_payload_40_real = _zz_175;
  assign fft_input_flow_payload_40_imag = _zz_176;
  assign fft_input_flow_payload_41_real = _zz_173;
  assign fft_input_flow_payload_41_imag = _zz_174;
  assign fft_input_flow_payload_42_real = _zz_171;
  assign fft_input_flow_payload_42_imag = _zz_172;
  assign fft_input_flow_payload_43_real = _zz_169;
  assign fft_input_flow_payload_43_imag = _zz_170;
  assign fft_input_flow_payload_44_real = _zz_167;
  assign fft_input_flow_payload_44_imag = _zz_168;
  assign fft_input_flow_payload_45_real = _zz_165;
  assign fft_input_flow_payload_45_imag = _zz_166;
  assign fft_input_flow_payload_46_real = _zz_163;
  assign fft_input_flow_payload_46_imag = _zz_164;
  assign fft_input_flow_payload_47_real = _zz_161;
  assign fft_input_flow_payload_47_imag = _zz_162;
  assign fft_input_flow_payload_48_real = _zz_159;
  assign fft_input_flow_payload_48_imag = _zz_160;
  assign fft_input_flow_payload_49_real = _zz_157;
  assign fft_input_flow_payload_49_imag = _zz_158;
  assign fft_input_flow_payload_50_real = _zz_155;
  assign fft_input_flow_payload_50_imag = _zz_156;
  assign fft_input_flow_payload_51_real = _zz_153;
  assign fft_input_flow_payload_51_imag = _zz_154;
  assign fft_input_flow_payload_52_real = _zz_151;
  assign fft_input_flow_payload_52_imag = _zz_152;
  assign fft_input_flow_payload_53_real = _zz_149;
  assign fft_input_flow_payload_53_imag = _zz_150;
  assign fft_input_flow_payload_54_real = _zz_147;
  assign fft_input_flow_payload_54_imag = _zz_148;
  assign fft_input_flow_payload_55_real = _zz_145;
  assign fft_input_flow_payload_55_imag = _zz_146;
  assign fft_input_flow_payload_56_real = _zz_143;
  assign fft_input_flow_payload_56_imag = _zz_144;
  assign fft_input_flow_payload_57_real = _zz_141;
  assign fft_input_flow_payload_57_imag = _zz_142;
  assign fft_input_flow_payload_58_real = _zz_139;
  assign fft_input_flow_payload_58_imag = _zz_140;
  assign fft_input_flow_payload_59_real = _zz_137;
  assign fft_input_flow_payload_59_imag = _zz_138;
  assign fft_input_flow_payload_60_real = _zz_135;
  assign fft_input_flow_payload_60_imag = _zz_136;
  assign fft_input_flow_payload_61_real = _zz_133;
  assign fft_input_flow_payload_61_imag = _zz_134;
  assign fft_input_flow_payload_62_real = _zz_131;
  assign fft_input_flow_payload_62_imag = _zz_132;
  assign fft_input_flow_payload_63_real = _zz_129;
  assign fft_input_flow_payload_63_imag = _zz_130;
  assign fft_input_flow_payload_64_real = _zz_127;
  assign fft_input_flow_payload_64_imag = _zz_128;
  assign fft_input_flow_payload_65_real = _zz_125;
  assign fft_input_flow_payload_65_imag = _zz_126;
  assign fft_input_flow_payload_66_real = _zz_123;
  assign fft_input_flow_payload_66_imag = _zz_124;
  assign fft_input_flow_payload_67_real = _zz_121;
  assign fft_input_flow_payload_67_imag = _zz_122;
  assign fft_input_flow_payload_68_real = _zz_119;
  assign fft_input_flow_payload_68_imag = _zz_120;
  assign fft_input_flow_payload_69_real = _zz_117;
  assign fft_input_flow_payload_69_imag = _zz_118;
  assign fft_input_flow_payload_70_real = _zz_115;
  assign fft_input_flow_payload_70_imag = _zz_116;
  assign fft_input_flow_payload_71_real = _zz_113;
  assign fft_input_flow_payload_71_imag = _zz_114;
  assign fft_input_flow_payload_72_real = _zz_111;
  assign fft_input_flow_payload_72_imag = _zz_112;
  assign fft_input_flow_payload_73_real = _zz_109;
  assign fft_input_flow_payload_73_imag = _zz_110;
  assign fft_input_flow_payload_74_real = _zz_107;
  assign fft_input_flow_payload_74_imag = _zz_108;
  assign fft_input_flow_payload_75_real = _zz_105;
  assign fft_input_flow_payload_75_imag = _zz_106;
  assign fft_input_flow_payload_76_real = _zz_103;
  assign fft_input_flow_payload_76_imag = _zz_104;
  assign fft_input_flow_payload_77_real = _zz_101;
  assign fft_input_flow_payload_77_imag = _zz_102;
  assign fft_input_flow_payload_78_real = _zz_99;
  assign fft_input_flow_payload_78_imag = _zz_100;
  assign fft_input_flow_payload_79_real = _zz_97;
  assign fft_input_flow_payload_79_imag = _zz_98;
  assign fft_input_flow_payload_80_real = _zz_95;
  assign fft_input_flow_payload_80_imag = _zz_96;
  assign fft_input_flow_payload_81_real = _zz_93;
  assign fft_input_flow_payload_81_imag = _zz_94;
  assign fft_input_flow_payload_82_real = _zz_91;
  assign fft_input_flow_payload_82_imag = _zz_92;
  assign fft_input_flow_payload_83_real = _zz_89;
  assign fft_input_flow_payload_83_imag = _zz_90;
  assign fft_input_flow_payload_84_real = _zz_87;
  assign fft_input_flow_payload_84_imag = _zz_88;
  assign fft_input_flow_payload_85_real = _zz_85;
  assign fft_input_flow_payload_85_imag = _zz_86;
  assign fft_input_flow_payload_86_real = _zz_83;
  assign fft_input_flow_payload_86_imag = _zz_84;
  assign fft_input_flow_payload_87_real = _zz_81;
  assign fft_input_flow_payload_87_imag = _zz_82;
  assign fft_input_flow_payload_88_real = _zz_79;
  assign fft_input_flow_payload_88_imag = _zz_80;
  assign fft_input_flow_payload_89_real = _zz_77;
  assign fft_input_flow_payload_89_imag = _zz_78;
  assign fft_input_flow_payload_90_real = _zz_75;
  assign fft_input_flow_payload_90_imag = _zz_76;
  assign fft_input_flow_payload_91_real = _zz_73;
  assign fft_input_flow_payload_91_imag = _zz_74;
  assign fft_input_flow_payload_92_real = _zz_71;
  assign fft_input_flow_payload_92_imag = _zz_72;
  assign fft_input_flow_payload_93_real = _zz_69;
  assign fft_input_flow_payload_93_imag = _zz_70;
  assign fft_input_flow_payload_94_real = _zz_67;
  assign fft_input_flow_payload_94_imag = _zz_68;
  assign fft_input_flow_payload_95_real = _zz_65;
  assign fft_input_flow_payload_95_imag = _zz_66;
  assign fft_input_flow_payload_96_real = _zz_63;
  assign fft_input_flow_payload_96_imag = _zz_64;
  assign fft_input_flow_payload_97_real = _zz_61;
  assign fft_input_flow_payload_97_imag = _zz_62;
  assign fft_input_flow_payload_98_real = _zz_59;
  assign fft_input_flow_payload_98_imag = _zz_60;
  assign fft_input_flow_payload_99_real = _zz_57;
  assign fft_input_flow_payload_99_imag = _zz_58;
  assign fft_input_flow_payload_100_real = _zz_55;
  assign fft_input_flow_payload_100_imag = _zz_56;
  assign fft_input_flow_payload_101_real = _zz_53;
  assign fft_input_flow_payload_101_imag = _zz_54;
  assign fft_input_flow_payload_102_real = _zz_51;
  assign fft_input_flow_payload_102_imag = _zz_52;
  assign fft_input_flow_payload_103_real = _zz_49;
  assign fft_input_flow_payload_103_imag = _zz_50;
  assign fft_input_flow_payload_104_real = _zz_47;
  assign fft_input_flow_payload_104_imag = _zz_48;
  assign fft_input_flow_payload_105_real = _zz_45;
  assign fft_input_flow_payload_105_imag = _zz_46;
  assign fft_input_flow_payload_106_real = _zz_43;
  assign fft_input_flow_payload_106_imag = _zz_44;
  assign fft_input_flow_payload_107_real = _zz_41;
  assign fft_input_flow_payload_107_imag = _zz_42;
  assign fft_input_flow_payload_108_real = _zz_39;
  assign fft_input_flow_payload_108_imag = _zz_40;
  assign fft_input_flow_payload_109_real = _zz_37;
  assign fft_input_flow_payload_109_imag = _zz_38;
  assign fft_input_flow_payload_110_real = _zz_35;
  assign fft_input_flow_payload_110_imag = _zz_36;
  assign fft_input_flow_payload_111_real = _zz_33;
  assign fft_input_flow_payload_111_imag = _zz_34;
  assign fft_input_flow_payload_112_real = _zz_31;
  assign fft_input_flow_payload_112_imag = _zz_32;
  assign fft_input_flow_payload_113_real = _zz_29;
  assign fft_input_flow_payload_113_imag = _zz_30;
  assign fft_input_flow_payload_114_real = _zz_27;
  assign fft_input_flow_payload_114_imag = _zz_28;
  assign fft_input_flow_payload_115_real = _zz_25;
  assign fft_input_flow_payload_115_imag = _zz_26;
  assign fft_input_flow_payload_116_real = _zz_23;
  assign fft_input_flow_payload_116_imag = _zz_24;
  assign fft_input_flow_payload_117_real = _zz_21;
  assign fft_input_flow_payload_117_imag = _zz_22;
  assign fft_input_flow_payload_118_real = _zz_19;
  assign fft_input_flow_payload_118_imag = _zz_20;
  assign fft_input_flow_payload_119_real = _zz_17;
  assign fft_input_flow_payload_119_imag = _zz_18;
  assign fft_input_flow_payload_120_real = _zz_15;
  assign fft_input_flow_payload_120_imag = _zz_16;
  assign fft_input_flow_payload_121_real = _zz_13;
  assign fft_input_flow_payload_121_imag = _zz_14;
  assign fft_input_flow_payload_122_real = _zz_11;
  assign fft_input_flow_payload_122_imag = _zz_12;
  assign fft_input_flow_payload_123_real = _zz_9;
  assign fft_input_flow_payload_123_imag = _zz_10;
  assign fft_input_flow_payload_124_real = _zz_7;
  assign fft_input_flow_payload_124_imag = _zz_8;
  assign fft_input_flow_payload_125_real = _zz_5;
  assign fft_input_flow_payload_125_imag = _zz_6;
  assign fft_input_flow_payload_126_real = _zz_3;
  assign fft_input_flow_payload_126_imag = _zz_4;
  assign fft_input_flow_payload_127_real = _zz_1;
  assign fft_input_flow_payload_127_imag = _zz_2;
  always @ (*) begin
    count_up_inside_cnt_willIncrement = 1'b0;
    if(data_in_valid)begin
      count_up_inside_cnt_willIncrement = 1'b1;
    end
  end

  assign count_up_inside_cnt_willClear = 1'b0;
  assign count_up_inside_cnt_willOverflowIfInc = (count_up_inside_cnt_value == 7'h7f);
  assign count_up_inside_cnt_willOverflow = (count_up_inside_cnt_willOverflowIfInc && count_up_inside_cnt_willIncrement);
  always @ (*) begin
    count_up_inside_cnt_valueNext = (count_up_inside_cnt_value + _zz_260);
    if(count_up_inside_cnt_willClear)begin
      count_up_inside_cnt_valueNext = 7'h0;
    end
  end

  assign fft_input_flow_valid = count_up_inside_cnt_willOverflow;
  always @ (*) begin
    null_cnt_willIncrement = 1'b0;
    if(null_cond_period)begin
      null_cnt_willIncrement = 1'b1;
    end
  end

  assign null_cnt_willClear = 1'b0;
  assign null_cnt_willOverflowIfInc = (null_cnt_value == 7'h7f);
  assign null_cnt_willOverflow = (null_cnt_willOverflowIfInc && null_cnt_willIncrement);
  always @ (*) begin
    null_cnt_valueNext = (null_cnt_value + _zz_262);
    if(null_cnt_willClear)begin
      null_cnt_valueNext = 7'h0;
    end
  end

  assign null_cond_period = (myFFT_1_sdata_out_valid_regNext || null_cond_period_minus_1);
  assign output_payload_real = _zz_257;
  assign output_payload_imag = _zz_258;
  assign output_valid = null_cond_period;
  assign data_out_valid = output_valid;
  assign data_out_payload_real = output_payload_real;
  assign data_out_payload_imag = output_payload_imag;
  always @ (posedge clk) begin
    if(data_in_valid)begin
      _zz_3 <= _zz_1;
      _zz_4 <= _zz_2;
    end
    if(data_in_valid)begin
      _zz_5 <= _zz_3;
      _zz_6 <= _zz_4;
    end
    if(data_in_valid)begin
      _zz_7 <= _zz_5;
      _zz_8 <= _zz_6;
    end
    if(data_in_valid)begin
      _zz_9 <= _zz_7;
      _zz_10 <= _zz_8;
    end
    if(data_in_valid)begin
      _zz_11 <= _zz_9;
      _zz_12 <= _zz_10;
    end
    if(data_in_valid)begin
      _zz_13 <= _zz_11;
      _zz_14 <= _zz_12;
    end
    if(data_in_valid)begin
      _zz_15 <= _zz_13;
      _zz_16 <= _zz_14;
    end
    if(data_in_valid)begin
      _zz_17 <= _zz_15;
      _zz_18 <= _zz_16;
    end
    if(data_in_valid)begin
      _zz_19 <= _zz_17;
      _zz_20 <= _zz_18;
    end
    if(data_in_valid)begin
      _zz_21 <= _zz_19;
      _zz_22 <= _zz_20;
    end
    if(data_in_valid)begin
      _zz_23 <= _zz_21;
      _zz_24 <= _zz_22;
    end
    if(data_in_valid)begin
      _zz_25 <= _zz_23;
      _zz_26 <= _zz_24;
    end
    if(data_in_valid)begin
      _zz_27 <= _zz_25;
      _zz_28 <= _zz_26;
    end
    if(data_in_valid)begin
      _zz_29 <= _zz_27;
      _zz_30 <= _zz_28;
    end
    if(data_in_valid)begin
      _zz_31 <= _zz_29;
      _zz_32 <= _zz_30;
    end
    if(data_in_valid)begin
      _zz_33 <= _zz_31;
      _zz_34 <= _zz_32;
    end
    if(data_in_valid)begin
      _zz_35 <= _zz_33;
      _zz_36 <= _zz_34;
    end
    if(data_in_valid)begin
      _zz_37 <= _zz_35;
      _zz_38 <= _zz_36;
    end
    if(data_in_valid)begin
      _zz_39 <= _zz_37;
      _zz_40 <= _zz_38;
    end
    if(data_in_valid)begin
      _zz_41 <= _zz_39;
      _zz_42 <= _zz_40;
    end
    if(data_in_valid)begin
      _zz_43 <= _zz_41;
      _zz_44 <= _zz_42;
    end
    if(data_in_valid)begin
      _zz_45 <= _zz_43;
      _zz_46 <= _zz_44;
    end
    if(data_in_valid)begin
      _zz_47 <= _zz_45;
      _zz_48 <= _zz_46;
    end
    if(data_in_valid)begin
      _zz_49 <= _zz_47;
      _zz_50 <= _zz_48;
    end
    if(data_in_valid)begin
      _zz_51 <= _zz_49;
      _zz_52 <= _zz_50;
    end
    if(data_in_valid)begin
      _zz_53 <= _zz_51;
      _zz_54 <= _zz_52;
    end
    if(data_in_valid)begin
      _zz_55 <= _zz_53;
      _zz_56 <= _zz_54;
    end
    if(data_in_valid)begin
      _zz_57 <= _zz_55;
      _zz_58 <= _zz_56;
    end
    if(data_in_valid)begin
      _zz_59 <= _zz_57;
      _zz_60 <= _zz_58;
    end
    if(data_in_valid)begin
      _zz_61 <= _zz_59;
      _zz_62 <= _zz_60;
    end
    if(data_in_valid)begin
      _zz_63 <= _zz_61;
      _zz_64 <= _zz_62;
    end
    if(data_in_valid)begin
      _zz_65 <= _zz_63;
      _zz_66 <= _zz_64;
    end
    if(data_in_valid)begin
      _zz_67 <= _zz_65;
      _zz_68 <= _zz_66;
    end
    if(data_in_valid)begin
      _zz_69 <= _zz_67;
      _zz_70 <= _zz_68;
    end
    if(data_in_valid)begin
      _zz_71 <= _zz_69;
      _zz_72 <= _zz_70;
    end
    if(data_in_valid)begin
      _zz_73 <= _zz_71;
      _zz_74 <= _zz_72;
    end
    if(data_in_valid)begin
      _zz_75 <= _zz_73;
      _zz_76 <= _zz_74;
    end
    if(data_in_valid)begin
      _zz_77 <= _zz_75;
      _zz_78 <= _zz_76;
    end
    if(data_in_valid)begin
      _zz_79 <= _zz_77;
      _zz_80 <= _zz_78;
    end
    if(data_in_valid)begin
      _zz_81 <= _zz_79;
      _zz_82 <= _zz_80;
    end
    if(data_in_valid)begin
      _zz_83 <= _zz_81;
      _zz_84 <= _zz_82;
    end
    if(data_in_valid)begin
      _zz_85 <= _zz_83;
      _zz_86 <= _zz_84;
    end
    if(data_in_valid)begin
      _zz_87 <= _zz_85;
      _zz_88 <= _zz_86;
    end
    if(data_in_valid)begin
      _zz_89 <= _zz_87;
      _zz_90 <= _zz_88;
    end
    if(data_in_valid)begin
      _zz_91 <= _zz_89;
      _zz_92 <= _zz_90;
    end
    if(data_in_valid)begin
      _zz_93 <= _zz_91;
      _zz_94 <= _zz_92;
    end
    if(data_in_valid)begin
      _zz_95 <= _zz_93;
      _zz_96 <= _zz_94;
    end
    if(data_in_valid)begin
      _zz_97 <= _zz_95;
      _zz_98 <= _zz_96;
    end
    if(data_in_valid)begin
      _zz_99 <= _zz_97;
      _zz_100 <= _zz_98;
    end
    if(data_in_valid)begin
      _zz_101 <= _zz_99;
      _zz_102 <= _zz_100;
    end
    if(data_in_valid)begin
      _zz_103 <= _zz_101;
      _zz_104 <= _zz_102;
    end
    if(data_in_valid)begin
      _zz_105 <= _zz_103;
      _zz_106 <= _zz_104;
    end
    if(data_in_valid)begin
      _zz_107 <= _zz_105;
      _zz_108 <= _zz_106;
    end
    if(data_in_valid)begin
      _zz_109 <= _zz_107;
      _zz_110 <= _zz_108;
    end
    if(data_in_valid)begin
      _zz_111 <= _zz_109;
      _zz_112 <= _zz_110;
    end
    if(data_in_valid)begin
      _zz_113 <= _zz_111;
      _zz_114 <= _zz_112;
    end
    if(data_in_valid)begin
      _zz_115 <= _zz_113;
      _zz_116 <= _zz_114;
    end
    if(data_in_valid)begin
      _zz_117 <= _zz_115;
      _zz_118 <= _zz_116;
    end
    if(data_in_valid)begin
      _zz_119 <= _zz_117;
      _zz_120 <= _zz_118;
    end
    if(data_in_valid)begin
      _zz_121 <= _zz_119;
      _zz_122 <= _zz_120;
    end
    if(data_in_valid)begin
      _zz_123 <= _zz_121;
      _zz_124 <= _zz_122;
    end
    if(data_in_valid)begin
      _zz_125 <= _zz_123;
      _zz_126 <= _zz_124;
    end
    if(data_in_valid)begin
      _zz_127 <= _zz_125;
      _zz_128 <= _zz_126;
    end
    if(data_in_valid)begin
      _zz_129 <= _zz_127;
      _zz_130 <= _zz_128;
    end
    if(data_in_valid)begin
      _zz_131 <= _zz_129;
      _zz_132 <= _zz_130;
    end
    if(data_in_valid)begin
      _zz_133 <= _zz_131;
      _zz_134 <= _zz_132;
    end
    if(data_in_valid)begin
      _zz_135 <= _zz_133;
      _zz_136 <= _zz_134;
    end
    if(data_in_valid)begin
      _zz_137 <= _zz_135;
      _zz_138 <= _zz_136;
    end
    if(data_in_valid)begin
      _zz_139 <= _zz_137;
      _zz_140 <= _zz_138;
    end
    if(data_in_valid)begin
      _zz_141 <= _zz_139;
      _zz_142 <= _zz_140;
    end
    if(data_in_valid)begin
      _zz_143 <= _zz_141;
      _zz_144 <= _zz_142;
    end
    if(data_in_valid)begin
      _zz_145 <= _zz_143;
      _zz_146 <= _zz_144;
    end
    if(data_in_valid)begin
      _zz_147 <= _zz_145;
      _zz_148 <= _zz_146;
    end
    if(data_in_valid)begin
      _zz_149 <= _zz_147;
      _zz_150 <= _zz_148;
    end
    if(data_in_valid)begin
      _zz_151 <= _zz_149;
      _zz_152 <= _zz_150;
    end
    if(data_in_valid)begin
      _zz_153 <= _zz_151;
      _zz_154 <= _zz_152;
    end
    if(data_in_valid)begin
      _zz_155 <= _zz_153;
      _zz_156 <= _zz_154;
    end
    if(data_in_valid)begin
      _zz_157 <= _zz_155;
      _zz_158 <= _zz_156;
    end
    if(data_in_valid)begin
      _zz_159 <= _zz_157;
      _zz_160 <= _zz_158;
    end
    if(data_in_valid)begin
      _zz_161 <= _zz_159;
      _zz_162 <= _zz_160;
    end
    if(data_in_valid)begin
      _zz_163 <= _zz_161;
      _zz_164 <= _zz_162;
    end
    if(data_in_valid)begin
      _zz_165 <= _zz_163;
      _zz_166 <= _zz_164;
    end
    if(data_in_valid)begin
      _zz_167 <= _zz_165;
      _zz_168 <= _zz_166;
    end
    if(data_in_valid)begin
      _zz_169 <= _zz_167;
      _zz_170 <= _zz_168;
    end
    if(data_in_valid)begin
      _zz_171 <= _zz_169;
      _zz_172 <= _zz_170;
    end
    if(data_in_valid)begin
      _zz_173 <= _zz_171;
      _zz_174 <= _zz_172;
    end
    if(data_in_valid)begin
      _zz_175 <= _zz_173;
      _zz_176 <= _zz_174;
    end
    if(data_in_valid)begin
      _zz_177 <= _zz_175;
      _zz_178 <= _zz_176;
    end
    if(data_in_valid)begin
      _zz_179 <= _zz_177;
      _zz_180 <= _zz_178;
    end
    if(data_in_valid)begin
      _zz_181 <= _zz_179;
      _zz_182 <= _zz_180;
    end
    if(data_in_valid)begin
      _zz_183 <= _zz_181;
      _zz_184 <= _zz_182;
    end
    if(data_in_valid)begin
      _zz_185 <= _zz_183;
      _zz_186 <= _zz_184;
    end
    if(data_in_valid)begin
      _zz_187 <= _zz_185;
      _zz_188 <= _zz_186;
    end
    if(data_in_valid)begin
      _zz_189 <= _zz_187;
      _zz_190 <= _zz_188;
    end
    if(data_in_valid)begin
      _zz_191 <= _zz_189;
      _zz_192 <= _zz_190;
    end
    if(data_in_valid)begin
      _zz_193 <= _zz_191;
      _zz_194 <= _zz_192;
    end
    if(data_in_valid)begin
      _zz_195 <= _zz_193;
      _zz_196 <= _zz_194;
    end
    if(data_in_valid)begin
      _zz_197 <= _zz_195;
      _zz_198 <= _zz_196;
    end
    if(data_in_valid)begin
      _zz_199 <= _zz_197;
      _zz_200 <= _zz_198;
    end
    if(data_in_valid)begin
      _zz_201 <= _zz_199;
      _zz_202 <= _zz_200;
    end
    if(data_in_valid)begin
      _zz_203 <= _zz_201;
      _zz_204 <= _zz_202;
    end
    if(data_in_valid)begin
      _zz_205 <= _zz_203;
      _zz_206 <= _zz_204;
    end
    if(data_in_valid)begin
      _zz_207 <= _zz_205;
      _zz_208 <= _zz_206;
    end
    if(data_in_valid)begin
      _zz_209 <= _zz_207;
      _zz_210 <= _zz_208;
    end
    if(data_in_valid)begin
      _zz_211 <= _zz_209;
      _zz_212 <= _zz_210;
    end
    if(data_in_valid)begin
      _zz_213 <= _zz_211;
      _zz_214 <= _zz_212;
    end
    if(data_in_valid)begin
      _zz_215 <= _zz_213;
      _zz_216 <= _zz_214;
    end
    if(data_in_valid)begin
      _zz_217 <= _zz_215;
      _zz_218 <= _zz_216;
    end
    if(data_in_valid)begin
      _zz_219 <= _zz_217;
      _zz_220 <= _zz_218;
    end
    if(data_in_valid)begin
      _zz_221 <= _zz_219;
      _zz_222 <= _zz_220;
    end
    if(data_in_valid)begin
      _zz_223 <= _zz_221;
      _zz_224 <= _zz_222;
    end
    if(data_in_valid)begin
      _zz_225 <= _zz_223;
      _zz_226 <= _zz_224;
    end
    if(data_in_valid)begin
      _zz_227 <= _zz_225;
      _zz_228 <= _zz_226;
    end
    if(data_in_valid)begin
      _zz_229 <= _zz_227;
      _zz_230 <= _zz_228;
    end
    if(data_in_valid)begin
      _zz_231 <= _zz_229;
      _zz_232 <= _zz_230;
    end
    if(data_in_valid)begin
      _zz_233 <= _zz_231;
      _zz_234 <= _zz_232;
    end
    if(data_in_valid)begin
      _zz_235 <= _zz_233;
      _zz_236 <= _zz_234;
    end
    if(data_in_valid)begin
      _zz_237 <= _zz_235;
      _zz_238 <= _zz_236;
    end
    if(data_in_valid)begin
      _zz_239 <= _zz_237;
      _zz_240 <= _zz_238;
    end
    if(data_in_valid)begin
      _zz_241 <= _zz_239;
      _zz_242 <= _zz_240;
    end
    if(data_in_valid)begin
      _zz_243 <= _zz_241;
      _zz_244 <= _zz_242;
    end
    if(data_in_valid)begin
      _zz_245 <= _zz_243;
      _zz_246 <= _zz_244;
    end
    if(data_in_valid)begin
      _zz_247 <= _zz_245;
      _zz_248 <= _zz_246;
    end
    if(data_in_valid)begin
      _zz_249 <= _zz_247;
      _zz_250 <= _zz_248;
    end
    if(data_in_valid)begin
      _zz_251 <= _zz_249;
      _zz_252 <= _zz_250;
    end
    if(data_in_valid)begin
      _zz_253 <= _zz_251;
      _zz_254 <= _zz_252;
    end
    if(data_in_valid)begin
      _zz_255 <= _zz_253;
      _zz_256 <= _zz_254;
    end
    if(myFFT_1_sdata_out_valid)begin
      sdata_out_regs_0_real <= myFFT_1_sdata_out_payload_0_real;
      sdata_out_regs_0_imag <= myFFT_1_sdata_out_payload_0_imag;
      sdata_out_regs_1_real <= myFFT_1_sdata_out_payload_1_real;
      sdata_out_regs_1_imag <= myFFT_1_sdata_out_payload_1_imag;
      sdata_out_regs_2_real <= myFFT_1_sdata_out_payload_2_real;
      sdata_out_regs_2_imag <= myFFT_1_sdata_out_payload_2_imag;
      sdata_out_regs_3_real <= myFFT_1_sdata_out_payload_3_real;
      sdata_out_regs_3_imag <= myFFT_1_sdata_out_payload_3_imag;
      sdata_out_regs_4_real <= myFFT_1_sdata_out_payload_4_real;
      sdata_out_regs_4_imag <= myFFT_1_sdata_out_payload_4_imag;
      sdata_out_regs_5_real <= myFFT_1_sdata_out_payload_5_real;
      sdata_out_regs_5_imag <= myFFT_1_sdata_out_payload_5_imag;
      sdata_out_regs_6_real <= myFFT_1_sdata_out_payload_6_real;
      sdata_out_regs_6_imag <= myFFT_1_sdata_out_payload_6_imag;
      sdata_out_regs_7_real <= myFFT_1_sdata_out_payload_7_real;
      sdata_out_regs_7_imag <= myFFT_1_sdata_out_payload_7_imag;
      sdata_out_regs_8_real <= myFFT_1_sdata_out_payload_8_real;
      sdata_out_regs_8_imag <= myFFT_1_sdata_out_payload_8_imag;
      sdata_out_regs_9_real <= myFFT_1_sdata_out_payload_9_real;
      sdata_out_regs_9_imag <= myFFT_1_sdata_out_payload_9_imag;
      sdata_out_regs_10_real <= myFFT_1_sdata_out_payload_10_real;
      sdata_out_regs_10_imag <= myFFT_1_sdata_out_payload_10_imag;
      sdata_out_regs_11_real <= myFFT_1_sdata_out_payload_11_real;
      sdata_out_regs_11_imag <= myFFT_1_sdata_out_payload_11_imag;
      sdata_out_regs_12_real <= myFFT_1_sdata_out_payload_12_real;
      sdata_out_regs_12_imag <= myFFT_1_sdata_out_payload_12_imag;
      sdata_out_regs_13_real <= myFFT_1_sdata_out_payload_13_real;
      sdata_out_regs_13_imag <= myFFT_1_sdata_out_payload_13_imag;
      sdata_out_regs_14_real <= myFFT_1_sdata_out_payload_14_real;
      sdata_out_regs_14_imag <= myFFT_1_sdata_out_payload_14_imag;
      sdata_out_regs_15_real <= myFFT_1_sdata_out_payload_15_real;
      sdata_out_regs_15_imag <= myFFT_1_sdata_out_payload_15_imag;
      sdata_out_regs_16_real <= myFFT_1_sdata_out_payload_16_real;
      sdata_out_regs_16_imag <= myFFT_1_sdata_out_payload_16_imag;
      sdata_out_regs_17_real <= myFFT_1_sdata_out_payload_17_real;
      sdata_out_regs_17_imag <= myFFT_1_sdata_out_payload_17_imag;
      sdata_out_regs_18_real <= myFFT_1_sdata_out_payload_18_real;
      sdata_out_regs_18_imag <= myFFT_1_sdata_out_payload_18_imag;
      sdata_out_regs_19_real <= myFFT_1_sdata_out_payload_19_real;
      sdata_out_regs_19_imag <= myFFT_1_sdata_out_payload_19_imag;
      sdata_out_regs_20_real <= myFFT_1_sdata_out_payload_20_real;
      sdata_out_regs_20_imag <= myFFT_1_sdata_out_payload_20_imag;
      sdata_out_regs_21_real <= myFFT_1_sdata_out_payload_21_real;
      sdata_out_regs_21_imag <= myFFT_1_sdata_out_payload_21_imag;
      sdata_out_regs_22_real <= myFFT_1_sdata_out_payload_22_real;
      sdata_out_regs_22_imag <= myFFT_1_sdata_out_payload_22_imag;
      sdata_out_regs_23_real <= myFFT_1_sdata_out_payload_23_real;
      sdata_out_regs_23_imag <= myFFT_1_sdata_out_payload_23_imag;
      sdata_out_regs_24_real <= myFFT_1_sdata_out_payload_24_real;
      sdata_out_regs_24_imag <= myFFT_1_sdata_out_payload_24_imag;
      sdata_out_regs_25_real <= myFFT_1_sdata_out_payload_25_real;
      sdata_out_regs_25_imag <= myFFT_1_sdata_out_payload_25_imag;
      sdata_out_regs_26_real <= myFFT_1_sdata_out_payload_26_real;
      sdata_out_regs_26_imag <= myFFT_1_sdata_out_payload_26_imag;
      sdata_out_regs_27_real <= myFFT_1_sdata_out_payload_27_real;
      sdata_out_regs_27_imag <= myFFT_1_sdata_out_payload_27_imag;
      sdata_out_regs_28_real <= myFFT_1_sdata_out_payload_28_real;
      sdata_out_regs_28_imag <= myFFT_1_sdata_out_payload_28_imag;
      sdata_out_regs_29_real <= myFFT_1_sdata_out_payload_29_real;
      sdata_out_regs_29_imag <= myFFT_1_sdata_out_payload_29_imag;
      sdata_out_regs_30_real <= myFFT_1_sdata_out_payload_30_real;
      sdata_out_regs_30_imag <= myFFT_1_sdata_out_payload_30_imag;
      sdata_out_regs_31_real <= myFFT_1_sdata_out_payload_31_real;
      sdata_out_regs_31_imag <= myFFT_1_sdata_out_payload_31_imag;
      sdata_out_regs_32_real <= myFFT_1_sdata_out_payload_32_real;
      sdata_out_regs_32_imag <= myFFT_1_sdata_out_payload_32_imag;
      sdata_out_regs_33_real <= myFFT_1_sdata_out_payload_33_real;
      sdata_out_regs_33_imag <= myFFT_1_sdata_out_payload_33_imag;
      sdata_out_regs_34_real <= myFFT_1_sdata_out_payload_34_real;
      sdata_out_regs_34_imag <= myFFT_1_sdata_out_payload_34_imag;
      sdata_out_regs_35_real <= myFFT_1_sdata_out_payload_35_real;
      sdata_out_regs_35_imag <= myFFT_1_sdata_out_payload_35_imag;
      sdata_out_regs_36_real <= myFFT_1_sdata_out_payload_36_real;
      sdata_out_regs_36_imag <= myFFT_1_sdata_out_payload_36_imag;
      sdata_out_regs_37_real <= myFFT_1_sdata_out_payload_37_real;
      sdata_out_regs_37_imag <= myFFT_1_sdata_out_payload_37_imag;
      sdata_out_regs_38_real <= myFFT_1_sdata_out_payload_38_real;
      sdata_out_regs_38_imag <= myFFT_1_sdata_out_payload_38_imag;
      sdata_out_regs_39_real <= myFFT_1_sdata_out_payload_39_real;
      sdata_out_regs_39_imag <= myFFT_1_sdata_out_payload_39_imag;
      sdata_out_regs_40_real <= myFFT_1_sdata_out_payload_40_real;
      sdata_out_regs_40_imag <= myFFT_1_sdata_out_payload_40_imag;
      sdata_out_regs_41_real <= myFFT_1_sdata_out_payload_41_real;
      sdata_out_regs_41_imag <= myFFT_1_sdata_out_payload_41_imag;
      sdata_out_regs_42_real <= myFFT_1_sdata_out_payload_42_real;
      sdata_out_regs_42_imag <= myFFT_1_sdata_out_payload_42_imag;
      sdata_out_regs_43_real <= myFFT_1_sdata_out_payload_43_real;
      sdata_out_regs_43_imag <= myFFT_1_sdata_out_payload_43_imag;
      sdata_out_regs_44_real <= myFFT_1_sdata_out_payload_44_real;
      sdata_out_regs_44_imag <= myFFT_1_sdata_out_payload_44_imag;
      sdata_out_regs_45_real <= myFFT_1_sdata_out_payload_45_real;
      sdata_out_regs_45_imag <= myFFT_1_sdata_out_payload_45_imag;
      sdata_out_regs_46_real <= myFFT_1_sdata_out_payload_46_real;
      sdata_out_regs_46_imag <= myFFT_1_sdata_out_payload_46_imag;
      sdata_out_regs_47_real <= myFFT_1_sdata_out_payload_47_real;
      sdata_out_regs_47_imag <= myFFT_1_sdata_out_payload_47_imag;
      sdata_out_regs_48_real <= myFFT_1_sdata_out_payload_48_real;
      sdata_out_regs_48_imag <= myFFT_1_sdata_out_payload_48_imag;
      sdata_out_regs_49_real <= myFFT_1_sdata_out_payload_49_real;
      sdata_out_regs_49_imag <= myFFT_1_sdata_out_payload_49_imag;
      sdata_out_regs_50_real <= myFFT_1_sdata_out_payload_50_real;
      sdata_out_regs_50_imag <= myFFT_1_sdata_out_payload_50_imag;
      sdata_out_regs_51_real <= myFFT_1_sdata_out_payload_51_real;
      sdata_out_regs_51_imag <= myFFT_1_sdata_out_payload_51_imag;
      sdata_out_regs_52_real <= myFFT_1_sdata_out_payload_52_real;
      sdata_out_regs_52_imag <= myFFT_1_sdata_out_payload_52_imag;
      sdata_out_regs_53_real <= myFFT_1_sdata_out_payload_53_real;
      sdata_out_regs_53_imag <= myFFT_1_sdata_out_payload_53_imag;
      sdata_out_regs_54_real <= myFFT_1_sdata_out_payload_54_real;
      sdata_out_regs_54_imag <= myFFT_1_sdata_out_payload_54_imag;
      sdata_out_regs_55_real <= myFFT_1_sdata_out_payload_55_real;
      sdata_out_regs_55_imag <= myFFT_1_sdata_out_payload_55_imag;
      sdata_out_regs_56_real <= myFFT_1_sdata_out_payload_56_real;
      sdata_out_regs_56_imag <= myFFT_1_sdata_out_payload_56_imag;
      sdata_out_regs_57_real <= myFFT_1_sdata_out_payload_57_real;
      sdata_out_regs_57_imag <= myFFT_1_sdata_out_payload_57_imag;
      sdata_out_regs_58_real <= myFFT_1_sdata_out_payload_58_real;
      sdata_out_regs_58_imag <= myFFT_1_sdata_out_payload_58_imag;
      sdata_out_regs_59_real <= myFFT_1_sdata_out_payload_59_real;
      sdata_out_regs_59_imag <= myFFT_1_sdata_out_payload_59_imag;
      sdata_out_regs_60_real <= myFFT_1_sdata_out_payload_60_real;
      sdata_out_regs_60_imag <= myFFT_1_sdata_out_payload_60_imag;
      sdata_out_regs_61_real <= myFFT_1_sdata_out_payload_61_real;
      sdata_out_regs_61_imag <= myFFT_1_sdata_out_payload_61_imag;
      sdata_out_regs_62_real <= myFFT_1_sdata_out_payload_62_real;
      sdata_out_regs_62_imag <= myFFT_1_sdata_out_payload_62_imag;
      sdata_out_regs_63_real <= myFFT_1_sdata_out_payload_63_real;
      sdata_out_regs_63_imag <= myFFT_1_sdata_out_payload_63_imag;
      sdata_out_regs_64_real <= myFFT_1_sdata_out_payload_64_real;
      sdata_out_regs_64_imag <= myFFT_1_sdata_out_payload_64_imag;
      sdata_out_regs_65_real <= myFFT_1_sdata_out_payload_65_real;
      sdata_out_regs_65_imag <= myFFT_1_sdata_out_payload_65_imag;
      sdata_out_regs_66_real <= myFFT_1_sdata_out_payload_66_real;
      sdata_out_regs_66_imag <= myFFT_1_sdata_out_payload_66_imag;
      sdata_out_regs_67_real <= myFFT_1_sdata_out_payload_67_real;
      sdata_out_regs_67_imag <= myFFT_1_sdata_out_payload_67_imag;
      sdata_out_regs_68_real <= myFFT_1_sdata_out_payload_68_real;
      sdata_out_regs_68_imag <= myFFT_1_sdata_out_payload_68_imag;
      sdata_out_regs_69_real <= myFFT_1_sdata_out_payload_69_real;
      sdata_out_regs_69_imag <= myFFT_1_sdata_out_payload_69_imag;
      sdata_out_regs_70_real <= myFFT_1_sdata_out_payload_70_real;
      sdata_out_regs_70_imag <= myFFT_1_sdata_out_payload_70_imag;
      sdata_out_regs_71_real <= myFFT_1_sdata_out_payload_71_real;
      sdata_out_regs_71_imag <= myFFT_1_sdata_out_payload_71_imag;
      sdata_out_regs_72_real <= myFFT_1_sdata_out_payload_72_real;
      sdata_out_regs_72_imag <= myFFT_1_sdata_out_payload_72_imag;
      sdata_out_regs_73_real <= myFFT_1_sdata_out_payload_73_real;
      sdata_out_regs_73_imag <= myFFT_1_sdata_out_payload_73_imag;
      sdata_out_regs_74_real <= myFFT_1_sdata_out_payload_74_real;
      sdata_out_regs_74_imag <= myFFT_1_sdata_out_payload_74_imag;
      sdata_out_regs_75_real <= myFFT_1_sdata_out_payload_75_real;
      sdata_out_regs_75_imag <= myFFT_1_sdata_out_payload_75_imag;
      sdata_out_regs_76_real <= myFFT_1_sdata_out_payload_76_real;
      sdata_out_regs_76_imag <= myFFT_1_sdata_out_payload_76_imag;
      sdata_out_regs_77_real <= myFFT_1_sdata_out_payload_77_real;
      sdata_out_regs_77_imag <= myFFT_1_sdata_out_payload_77_imag;
      sdata_out_regs_78_real <= myFFT_1_sdata_out_payload_78_real;
      sdata_out_regs_78_imag <= myFFT_1_sdata_out_payload_78_imag;
      sdata_out_regs_79_real <= myFFT_1_sdata_out_payload_79_real;
      sdata_out_regs_79_imag <= myFFT_1_sdata_out_payload_79_imag;
      sdata_out_regs_80_real <= myFFT_1_sdata_out_payload_80_real;
      sdata_out_regs_80_imag <= myFFT_1_sdata_out_payload_80_imag;
      sdata_out_regs_81_real <= myFFT_1_sdata_out_payload_81_real;
      sdata_out_regs_81_imag <= myFFT_1_sdata_out_payload_81_imag;
      sdata_out_regs_82_real <= myFFT_1_sdata_out_payload_82_real;
      sdata_out_regs_82_imag <= myFFT_1_sdata_out_payload_82_imag;
      sdata_out_regs_83_real <= myFFT_1_sdata_out_payload_83_real;
      sdata_out_regs_83_imag <= myFFT_1_sdata_out_payload_83_imag;
      sdata_out_regs_84_real <= myFFT_1_sdata_out_payload_84_real;
      sdata_out_regs_84_imag <= myFFT_1_sdata_out_payload_84_imag;
      sdata_out_regs_85_real <= myFFT_1_sdata_out_payload_85_real;
      sdata_out_regs_85_imag <= myFFT_1_sdata_out_payload_85_imag;
      sdata_out_regs_86_real <= myFFT_1_sdata_out_payload_86_real;
      sdata_out_regs_86_imag <= myFFT_1_sdata_out_payload_86_imag;
      sdata_out_regs_87_real <= myFFT_1_sdata_out_payload_87_real;
      sdata_out_regs_87_imag <= myFFT_1_sdata_out_payload_87_imag;
      sdata_out_regs_88_real <= myFFT_1_sdata_out_payload_88_real;
      sdata_out_regs_88_imag <= myFFT_1_sdata_out_payload_88_imag;
      sdata_out_regs_89_real <= myFFT_1_sdata_out_payload_89_real;
      sdata_out_regs_89_imag <= myFFT_1_sdata_out_payload_89_imag;
      sdata_out_regs_90_real <= myFFT_1_sdata_out_payload_90_real;
      sdata_out_regs_90_imag <= myFFT_1_sdata_out_payload_90_imag;
      sdata_out_regs_91_real <= myFFT_1_sdata_out_payload_91_real;
      sdata_out_regs_91_imag <= myFFT_1_sdata_out_payload_91_imag;
      sdata_out_regs_92_real <= myFFT_1_sdata_out_payload_92_real;
      sdata_out_regs_92_imag <= myFFT_1_sdata_out_payload_92_imag;
      sdata_out_regs_93_real <= myFFT_1_sdata_out_payload_93_real;
      sdata_out_regs_93_imag <= myFFT_1_sdata_out_payload_93_imag;
      sdata_out_regs_94_real <= myFFT_1_sdata_out_payload_94_real;
      sdata_out_regs_94_imag <= myFFT_1_sdata_out_payload_94_imag;
      sdata_out_regs_95_real <= myFFT_1_sdata_out_payload_95_real;
      sdata_out_regs_95_imag <= myFFT_1_sdata_out_payload_95_imag;
      sdata_out_regs_96_real <= myFFT_1_sdata_out_payload_96_real;
      sdata_out_regs_96_imag <= myFFT_1_sdata_out_payload_96_imag;
      sdata_out_regs_97_real <= myFFT_1_sdata_out_payload_97_real;
      sdata_out_regs_97_imag <= myFFT_1_sdata_out_payload_97_imag;
      sdata_out_regs_98_real <= myFFT_1_sdata_out_payload_98_real;
      sdata_out_regs_98_imag <= myFFT_1_sdata_out_payload_98_imag;
      sdata_out_regs_99_real <= myFFT_1_sdata_out_payload_99_real;
      sdata_out_regs_99_imag <= myFFT_1_sdata_out_payload_99_imag;
      sdata_out_regs_100_real <= myFFT_1_sdata_out_payload_100_real;
      sdata_out_regs_100_imag <= myFFT_1_sdata_out_payload_100_imag;
      sdata_out_regs_101_real <= myFFT_1_sdata_out_payload_101_real;
      sdata_out_regs_101_imag <= myFFT_1_sdata_out_payload_101_imag;
      sdata_out_regs_102_real <= myFFT_1_sdata_out_payload_102_real;
      sdata_out_regs_102_imag <= myFFT_1_sdata_out_payload_102_imag;
      sdata_out_regs_103_real <= myFFT_1_sdata_out_payload_103_real;
      sdata_out_regs_103_imag <= myFFT_1_sdata_out_payload_103_imag;
      sdata_out_regs_104_real <= myFFT_1_sdata_out_payload_104_real;
      sdata_out_regs_104_imag <= myFFT_1_sdata_out_payload_104_imag;
      sdata_out_regs_105_real <= myFFT_1_sdata_out_payload_105_real;
      sdata_out_regs_105_imag <= myFFT_1_sdata_out_payload_105_imag;
      sdata_out_regs_106_real <= myFFT_1_sdata_out_payload_106_real;
      sdata_out_regs_106_imag <= myFFT_1_sdata_out_payload_106_imag;
      sdata_out_regs_107_real <= myFFT_1_sdata_out_payload_107_real;
      sdata_out_regs_107_imag <= myFFT_1_sdata_out_payload_107_imag;
      sdata_out_regs_108_real <= myFFT_1_sdata_out_payload_108_real;
      sdata_out_regs_108_imag <= myFFT_1_sdata_out_payload_108_imag;
      sdata_out_regs_109_real <= myFFT_1_sdata_out_payload_109_real;
      sdata_out_regs_109_imag <= myFFT_1_sdata_out_payload_109_imag;
      sdata_out_regs_110_real <= myFFT_1_sdata_out_payload_110_real;
      sdata_out_regs_110_imag <= myFFT_1_sdata_out_payload_110_imag;
      sdata_out_regs_111_real <= myFFT_1_sdata_out_payload_111_real;
      sdata_out_regs_111_imag <= myFFT_1_sdata_out_payload_111_imag;
      sdata_out_regs_112_real <= myFFT_1_sdata_out_payload_112_real;
      sdata_out_regs_112_imag <= myFFT_1_sdata_out_payload_112_imag;
      sdata_out_regs_113_real <= myFFT_1_sdata_out_payload_113_real;
      sdata_out_regs_113_imag <= myFFT_1_sdata_out_payload_113_imag;
      sdata_out_regs_114_real <= myFFT_1_sdata_out_payload_114_real;
      sdata_out_regs_114_imag <= myFFT_1_sdata_out_payload_114_imag;
      sdata_out_regs_115_real <= myFFT_1_sdata_out_payload_115_real;
      sdata_out_regs_115_imag <= myFFT_1_sdata_out_payload_115_imag;
      sdata_out_regs_116_real <= myFFT_1_sdata_out_payload_116_real;
      sdata_out_regs_116_imag <= myFFT_1_sdata_out_payload_116_imag;
      sdata_out_regs_117_real <= myFFT_1_sdata_out_payload_117_real;
      sdata_out_regs_117_imag <= myFFT_1_sdata_out_payload_117_imag;
      sdata_out_regs_118_real <= myFFT_1_sdata_out_payload_118_real;
      sdata_out_regs_118_imag <= myFFT_1_sdata_out_payload_118_imag;
      sdata_out_regs_119_real <= myFFT_1_sdata_out_payload_119_real;
      sdata_out_regs_119_imag <= myFFT_1_sdata_out_payload_119_imag;
      sdata_out_regs_120_real <= myFFT_1_sdata_out_payload_120_real;
      sdata_out_regs_120_imag <= myFFT_1_sdata_out_payload_120_imag;
      sdata_out_regs_121_real <= myFFT_1_sdata_out_payload_121_real;
      sdata_out_regs_121_imag <= myFFT_1_sdata_out_payload_121_imag;
      sdata_out_regs_122_real <= myFFT_1_sdata_out_payload_122_real;
      sdata_out_regs_122_imag <= myFFT_1_sdata_out_payload_122_imag;
      sdata_out_regs_123_real <= myFFT_1_sdata_out_payload_123_real;
      sdata_out_regs_123_imag <= myFFT_1_sdata_out_payload_123_imag;
      sdata_out_regs_124_real <= myFFT_1_sdata_out_payload_124_real;
      sdata_out_regs_124_imag <= myFFT_1_sdata_out_payload_124_imag;
      sdata_out_regs_125_real <= myFFT_1_sdata_out_payload_125_real;
      sdata_out_regs_125_imag <= myFFT_1_sdata_out_payload_125_imag;
      sdata_out_regs_126_real <= myFFT_1_sdata_out_payload_126_real;
      sdata_out_regs_126_imag <= myFFT_1_sdata_out_payload_126_imag;
      sdata_out_regs_127_real <= myFFT_1_sdata_out_payload_127_real;
      sdata_out_regs_127_imag <= myFFT_1_sdata_out_payload_127_imag;
    end
  end

  always @ (posedge clk or posedge reset) begin
    if (reset) begin
      count_up_inside_cnt_value <= 7'h0;
      myFFT_1_sdata_out_valid_regNext <= 1'b0;
      null_cnt_value <= 7'h0;
      null_cond_period_minus_1 <= 1'b0;
    end else begin
      count_up_inside_cnt_value <= count_up_inside_cnt_valueNext;
      myFFT_1_sdata_out_valid_regNext <= myFFT_1_sdata_out_valid;
      null_cnt_value <= null_cnt_valueNext;
      if(myFFT_1_sdata_out_valid_regNext)begin
        null_cond_period_minus_1 <= 1'b1;
      end else begin
        if(null_cnt_willOverflow)begin
          null_cond_period_minus_1 <= 1'b0;
        end
      end
    end
  end


endmodule

module MyFFT (
  input               io_data_in_valid,
  input      [15:0]   io_data_in_payload_0_real,
  input      [15:0]   io_data_in_payload_0_imag,
  input      [15:0]   io_data_in_payload_1_real,
  input      [15:0]   io_data_in_payload_1_imag,
  input      [15:0]   io_data_in_payload_2_real,
  input      [15:0]   io_data_in_payload_2_imag,
  input      [15:0]   io_data_in_payload_3_real,
  input      [15:0]   io_data_in_payload_3_imag,
  input      [15:0]   io_data_in_payload_4_real,
  input      [15:0]   io_data_in_payload_4_imag,
  input      [15:0]   io_data_in_payload_5_real,
  input      [15:0]   io_data_in_payload_5_imag,
  input      [15:0]   io_data_in_payload_6_real,
  input      [15:0]   io_data_in_payload_6_imag,
  input      [15:0]   io_data_in_payload_7_real,
  input      [15:0]   io_data_in_payload_7_imag,
  input      [15:0]   io_data_in_payload_8_real,
  input      [15:0]   io_data_in_payload_8_imag,
  input      [15:0]   io_data_in_payload_9_real,
  input      [15:0]   io_data_in_payload_9_imag,
  input      [15:0]   io_data_in_payload_10_real,
  input      [15:0]   io_data_in_payload_10_imag,
  input      [15:0]   io_data_in_payload_11_real,
  input      [15:0]   io_data_in_payload_11_imag,
  input      [15:0]   io_data_in_payload_12_real,
  input      [15:0]   io_data_in_payload_12_imag,
  input      [15:0]   io_data_in_payload_13_real,
  input      [15:0]   io_data_in_payload_13_imag,
  input      [15:0]   io_data_in_payload_14_real,
  input      [15:0]   io_data_in_payload_14_imag,
  input      [15:0]   io_data_in_payload_15_real,
  input      [15:0]   io_data_in_payload_15_imag,
  input      [15:0]   io_data_in_payload_16_real,
  input      [15:0]   io_data_in_payload_16_imag,
  input      [15:0]   io_data_in_payload_17_real,
  input      [15:0]   io_data_in_payload_17_imag,
  input      [15:0]   io_data_in_payload_18_real,
  input      [15:0]   io_data_in_payload_18_imag,
  input      [15:0]   io_data_in_payload_19_real,
  input      [15:0]   io_data_in_payload_19_imag,
  input      [15:0]   io_data_in_payload_20_real,
  input      [15:0]   io_data_in_payload_20_imag,
  input      [15:0]   io_data_in_payload_21_real,
  input      [15:0]   io_data_in_payload_21_imag,
  input      [15:0]   io_data_in_payload_22_real,
  input      [15:0]   io_data_in_payload_22_imag,
  input      [15:0]   io_data_in_payload_23_real,
  input      [15:0]   io_data_in_payload_23_imag,
  input      [15:0]   io_data_in_payload_24_real,
  input      [15:0]   io_data_in_payload_24_imag,
  input      [15:0]   io_data_in_payload_25_real,
  input      [15:0]   io_data_in_payload_25_imag,
  input      [15:0]   io_data_in_payload_26_real,
  input      [15:0]   io_data_in_payload_26_imag,
  input      [15:0]   io_data_in_payload_27_real,
  input      [15:0]   io_data_in_payload_27_imag,
  input      [15:0]   io_data_in_payload_28_real,
  input      [15:0]   io_data_in_payload_28_imag,
  input      [15:0]   io_data_in_payload_29_real,
  input      [15:0]   io_data_in_payload_29_imag,
  input      [15:0]   io_data_in_payload_30_real,
  input      [15:0]   io_data_in_payload_30_imag,
  input      [15:0]   io_data_in_payload_31_real,
  input      [15:0]   io_data_in_payload_31_imag,
  input      [15:0]   io_data_in_payload_32_real,
  input      [15:0]   io_data_in_payload_32_imag,
  input      [15:0]   io_data_in_payload_33_real,
  input      [15:0]   io_data_in_payload_33_imag,
  input      [15:0]   io_data_in_payload_34_real,
  input      [15:0]   io_data_in_payload_34_imag,
  input      [15:0]   io_data_in_payload_35_real,
  input      [15:0]   io_data_in_payload_35_imag,
  input      [15:0]   io_data_in_payload_36_real,
  input      [15:0]   io_data_in_payload_36_imag,
  input      [15:0]   io_data_in_payload_37_real,
  input      [15:0]   io_data_in_payload_37_imag,
  input      [15:0]   io_data_in_payload_38_real,
  input      [15:0]   io_data_in_payload_38_imag,
  input      [15:0]   io_data_in_payload_39_real,
  input      [15:0]   io_data_in_payload_39_imag,
  input      [15:0]   io_data_in_payload_40_real,
  input      [15:0]   io_data_in_payload_40_imag,
  input      [15:0]   io_data_in_payload_41_real,
  input      [15:0]   io_data_in_payload_41_imag,
  input      [15:0]   io_data_in_payload_42_real,
  input      [15:0]   io_data_in_payload_42_imag,
  input      [15:0]   io_data_in_payload_43_real,
  input      [15:0]   io_data_in_payload_43_imag,
  input      [15:0]   io_data_in_payload_44_real,
  input      [15:0]   io_data_in_payload_44_imag,
  input      [15:0]   io_data_in_payload_45_real,
  input      [15:0]   io_data_in_payload_45_imag,
  input      [15:0]   io_data_in_payload_46_real,
  input      [15:0]   io_data_in_payload_46_imag,
  input      [15:0]   io_data_in_payload_47_real,
  input      [15:0]   io_data_in_payload_47_imag,
  input      [15:0]   io_data_in_payload_48_real,
  input      [15:0]   io_data_in_payload_48_imag,
  input      [15:0]   io_data_in_payload_49_real,
  input      [15:0]   io_data_in_payload_49_imag,
  input      [15:0]   io_data_in_payload_50_real,
  input      [15:0]   io_data_in_payload_50_imag,
  input      [15:0]   io_data_in_payload_51_real,
  input      [15:0]   io_data_in_payload_51_imag,
  input      [15:0]   io_data_in_payload_52_real,
  input      [15:0]   io_data_in_payload_52_imag,
  input      [15:0]   io_data_in_payload_53_real,
  input      [15:0]   io_data_in_payload_53_imag,
  input      [15:0]   io_data_in_payload_54_real,
  input      [15:0]   io_data_in_payload_54_imag,
  input      [15:0]   io_data_in_payload_55_real,
  input      [15:0]   io_data_in_payload_55_imag,
  input      [15:0]   io_data_in_payload_56_real,
  input      [15:0]   io_data_in_payload_56_imag,
  input      [15:0]   io_data_in_payload_57_real,
  input      [15:0]   io_data_in_payload_57_imag,
  input      [15:0]   io_data_in_payload_58_real,
  input      [15:0]   io_data_in_payload_58_imag,
  input      [15:0]   io_data_in_payload_59_real,
  input      [15:0]   io_data_in_payload_59_imag,
  input      [15:0]   io_data_in_payload_60_real,
  input      [15:0]   io_data_in_payload_60_imag,
  input      [15:0]   io_data_in_payload_61_real,
  input      [15:0]   io_data_in_payload_61_imag,
  input      [15:0]   io_data_in_payload_62_real,
  input      [15:0]   io_data_in_payload_62_imag,
  input      [15:0]   io_data_in_payload_63_real,
  input      [15:0]   io_data_in_payload_63_imag,
  input      [15:0]   io_data_in_payload_64_real,
  input      [15:0]   io_data_in_payload_64_imag,
  input      [15:0]   io_data_in_payload_65_real,
  input      [15:0]   io_data_in_payload_65_imag,
  input      [15:0]   io_data_in_payload_66_real,
  input      [15:0]   io_data_in_payload_66_imag,
  input      [15:0]   io_data_in_payload_67_real,
  input      [15:0]   io_data_in_payload_67_imag,
  input      [15:0]   io_data_in_payload_68_real,
  input      [15:0]   io_data_in_payload_68_imag,
  input      [15:0]   io_data_in_payload_69_real,
  input      [15:0]   io_data_in_payload_69_imag,
  input      [15:0]   io_data_in_payload_70_real,
  input      [15:0]   io_data_in_payload_70_imag,
  input      [15:0]   io_data_in_payload_71_real,
  input      [15:0]   io_data_in_payload_71_imag,
  input      [15:0]   io_data_in_payload_72_real,
  input      [15:0]   io_data_in_payload_72_imag,
  input      [15:0]   io_data_in_payload_73_real,
  input      [15:0]   io_data_in_payload_73_imag,
  input      [15:0]   io_data_in_payload_74_real,
  input      [15:0]   io_data_in_payload_74_imag,
  input      [15:0]   io_data_in_payload_75_real,
  input      [15:0]   io_data_in_payload_75_imag,
  input      [15:0]   io_data_in_payload_76_real,
  input      [15:0]   io_data_in_payload_76_imag,
  input      [15:0]   io_data_in_payload_77_real,
  input      [15:0]   io_data_in_payload_77_imag,
  input      [15:0]   io_data_in_payload_78_real,
  input      [15:0]   io_data_in_payload_78_imag,
  input      [15:0]   io_data_in_payload_79_real,
  input      [15:0]   io_data_in_payload_79_imag,
  input      [15:0]   io_data_in_payload_80_real,
  input      [15:0]   io_data_in_payload_80_imag,
  input      [15:0]   io_data_in_payload_81_real,
  input      [15:0]   io_data_in_payload_81_imag,
  input      [15:0]   io_data_in_payload_82_real,
  input      [15:0]   io_data_in_payload_82_imag,
  input      [15:0]   io_data_in_payload_83_real,
  input      [15:0]   io_data_in_payload_83_imag,
  input      [15:0]   io_data_in_payload_84_real,
  input      [15:0]   io_data_in_payload_84_imag,
  input      [15:0]   io_data_in_payload_85_real,
  input      [15:0]   io_data_in_payload_85_imag,
  input      [15:0]   io_data_in_payload_86_real,
  input      [15:0]   io_data_in_payload_86_imag,
  input      [15:0]   io_data_in_payload_87_real,
  input      [15:0]   io_data_in_payload_87_imag,
  input      [15:0]   io_data_in_payload_88_real,
  input      [15:0]   io_data_in_payload_88_imag,
  input      [15:0]   io_data_in_payload_89_real,
  input      [15:0]   io_data_in_payload_89_imag,
  input      [15:0]   io_data_in_payload_90_real,
  input      [15:0]   io_data_in_payload_90_imag,
  input      [15:0]   io_data_in_payload_91_real,
  input      [15:0]   io_data_in_payload_91_imag,
  input      [15:0]   io_data_in_payload_92_real,
  input      [15:0]   io_data_in_payload_92_imag,
  input      [15:0]   io_data_in_payload_93_real,
  input      [15:0]   io_data_in_payload_93_imag,
  input      [15:0]   io_data_in_payload_94_real,
  input      [15:0]   io_data_in_payload_94_imag,
  input      [15:0]   io_data_in_payload_95_real,
  input      [15:0]   io_data_in_payload_95_imag,
  input      [15:0]   io_data_in_payload_96_real,
  input      [15:0]   io_data_in_payload_96_imag,
  input      [15:0]   io_data_in_payload_97_real,
  input      [15:0]   io_data_in_payload_97_imag,
  input      [15:0]   io_data_in_payload_98_real,
  input      [15:0]   io_data_in_payload_98_imag,
  input      [15:0]   io_data_in_payload_99_real,
  input      [15:0]   io_data_in_payload_99_imag,
  input      [15:0]   io_data_in_payload_100_real,
  input      [15:0]   io_data_in_payload_100_imag,
  input      [15:0]   io_data_in_payload_101_real,
  input      [15:0]   io_data_in_payload_101_imag,
  input      [15:0]   io_data_in_payload_102_real,
  input      [15:0]   io_data_in_payload_102_imag,
  input      [15:0]   io_data_in_payload_103_real,
  input      [15:0]   io_data_in_payload_103_imag,
  input      [15:0]   io_data_in_payload_104_real,
  input      [15:0]   io_data_in_payload_104_imag,
  input      [15:0]   io_data_in_payload_105_real,
  input      [15:0]   io_data_in_payload_105_imag,
  input      [15:0]   io_data_in_payload_106_real,
  input      [15:0]   io_data_in_payload_106_imag,
  input      [15:0]   io_data_in_payload_107_real,
  input      [15:0]   io_data_in_payload_107_imag,
  input      [15:0]   io_data_in_payload_108_real,
  input      [15:0]   io_data_in_payload_108_imag,
  input      [15:0]   io_data_in_payload_109_real,
  input      [15:0]   io_data_in_payload_109_imag,
  input      [15:0]   io_data_in_payload_110_real,
  input      [15:0]   io_data_in_payload_110_imag,
  input      [15:0]   io_data_in_payload_111_real,
  input      [15:0]   io_data_in_payload_111_imag,
  input      [15:0]   io_data_in_payload_112_real,
  input      [15:0]   io_data_in_payload_112_imag,
  input      [15:0]   io_data_in_payload_113_real,
  input      [15:0]   io_data_in_payload_113_imag,
  input      [15:0]   io_data_in_payload_114_real,
  input      [15:0]   io_data_in_payload_114_imag,
  input      [15:0]   io_data_in_payload_115_real,
  input      [15:0]   io_data_in_payload_115_imag,
  input      [15:0]   io_data_in_payload_116_real,
  input      [15:0]   io_data_in_payload_116_imag,
  input      [15:0]   io_data_in_payload_117_real,
  input      [15:0]   io_data_in_payload_117_imag,
  input      [15:0]   io_data_in_payload_118_real,
  input      [15:0]   io_data_in_payload_118_imag,
  input      [15:0]   io_data_in_payload_119_real,
  input      [15:0]   io_data_in_payload_119_imag,
  input      [15:0]   io_data_in_payload_120_real,
  input      [15:0]   io_data_in_payload_120_imag,
  input      [15:0]   io_data_in_payload_121_real,
  input      [15:0]   io_data_in_payload_121_imag,
  input      [15:0]   io_data_in_payload_122_real,
  input      [15:0]   io_data_in_payload_122_imag,
  input      [15:0]   io_data_in_payload_123_real,
  input      [15:0]   io_data_in_payload_123_imag,
  input      [15:0]   io_data_in_payload_124_real,
  input      [15:0]   io_data_in_payload_124_imag,
  input      [15:0]   io_data_in_payload_125_real,
  input      [15:0]   io_data_in_payload_125_imag,
  input      [15:0]   io_data_in_payload_126_real,
  input      [15:0]   io_data_in_payload_126_imag,
  input      [15:0]   io_data_in_payload_127_real,
  input      [15:0]   io_data_in_payload_127_imag,
  output              sdata_out_valid,
  output     [15:0]   sdata_out_payload_0_real,
  output     [15:0]   sdata_out_payload_0_imag,
  output     [15:0]   sdata_out_payload_1_real,
  output     [15:0]   sdata_out_payload_1_imag,
  output     [15:0]   sdata_out_payload_2_real,
  output     [15:0]   sdata_out_payload_2_imag,
  output     [15:0]   sdata_out_payload_3_real,
  output     [15:0]   sdata_out_payload_3_imag,
  output     [15:0]   sdata_out_payload_4_real,
  output     [15:0]   sdata_out_payload_4_imag,
  output     [15:0]   sdata_out_payload_5_real,
  output     [15:0]   sdata_out_payload_5_imag,
  output     [15:0]   sdata_out_payload_6_real,
  output     [15:0]   sdata_out_payload_6_imag,
  output     [15:0]   sdata_out_payload_7_real,
  output     [15:0]   sdata_out_payload_7_imag,
  output     [15:0]   sdata_out_payload_8_real,
  output     [15:0]   sdata_out_payload_8_imag,
  output     [15:0]   sdata_out_payload_9_real,
  output     [15:0]   sdata_out_payload_9_imag,
  output     [15:0]   sdata_out_payload_10_real,
  output     [15:0]   sdata_out_payload_10_imag,
  output     [15:0]   sdata_out_payload_11_real,
  output     [15:0]   sdata_out_payload_11_imag,
  output     [15:0]   sdata_out_payload_12_real,
  output     [15:0]   sdata_out_payload_12_imag,
  output     [15:0]   sdata_out_payload_13_real,
  output     [15:0]   sdata_out_payload_13_imag,
  output     [15:0]   sdata_out_payload_14_real,
  output     [15:0]   sdata_out_payload_14_imag,
  output     [15:0]   sdata_out_payload_15_real,
  output     [15:0]   sdata_out_payload_15_imag,
  output     [15:0]   sdata_out_payload_16_real,
  output     [15:0]   sdata_out_payload_16_imag,
  output     [15:0]   sdata_out_payload_17_real,
  output     [15:0]   sdata_out_payload_17_imag,
  output     [15:0]   sdata_out_payload_18_real,
  output     [15:0]   sdata_out_payload_18_imag,
  output     [15:0]   sdata_out_payload_19_real,
  output     [15:0]   sdata_out_payload_19_imag,
  output     [15:0]   sdata_out_payload_20_real,
  output     [15:0]   sdata_out_payload_20_imag,
  output     [15:0]   sdata_out_payload_21_real,
  output     [15:0]   sdata_out_payload_21_imag,
  output     [15:0]   sdata_out_payload_22_real,
  output     [15:0]   sdata_out_payload_22_imag,
  output     [15:0]   sdata_out_payload_23_real,
  output     [15:0]   sdata_out_payload_23_imag,
  output     [15:0]   sdata_out_payload_24_real,
  output     [15:0]   sdata_out_payload_24_imag,
  output     [15:0]   sdata_out_payload_25_real,
  output     [15:0]   sdata_out_payload_25_imag,
  output     [15:0]   sdata_out_payload_26_real,
  output     [15:0]   sdata_out_payload_26_imag,
  output     [15:0]   sdata_out_payload_27_real,
  output     [15:0]   sdata_out_payload_27_imag,
  output     [15:0]   sdata_out_payload_28_real,
  output     [15:0]   sdata_out_payload_28_imag,
  output     [15:0]   sdata_out_payload_29_real,
  output     [15:0]   sdata_out_payload_29_imag,
  output     [15:0]   sdata_out_payload_30_real,
  output     [15:0]   sdata_out_payload_30_imag,
  output     [15:0]   sdata_out_payload_31_real,
  output     [15:0]   sdata_out_payload_31_imag,
  output     [15:0]   sdata_out_payload_32_real,
  output     [15:0]   sdata_out_payload_32_imag,
  output     [15:0]   sdata_out_payload_33_real,
  output     [15:0]   sdata_out_payload_33_imag,
  output     [15:0]   sdata_out_payload_34_real,
  output     [15:0]   sdata_out_payload_34_imag,
  output     [15:0]   sdata_out_payload_35_real,
  output     [15:0]   sdata_out_payload_35_imag,
  output     [15:0]   sdata_out_payload_36_real,
  output     [15:0]   sdata_out_payload_36_imag,
  output     [15:0]   sdata_out_payload_37_real,
  output     [15:0]   sdata_out_payload_37_imag,
  output     [15:0]   sdata_out_payload_38_real,
  output     [15:0]   sdata_out_payload_38_imag,
  output     [15:0]   sdata_out_payload_39_real,
  output     [15:0]   sdata_out_payload_39_imag,
  output     [15:0]   sdata_out_payload_40_real,
  output     [15:0]   sdata_out_payload_40_imag,
  output     [15:0]   sdata_out_payload_41_real,
  output     [15:0]   sdata_out_payload_41_imag,
  output     [15:0]   sdata_out_payload_42_real,
  output     [15:0]   sdata_out_payload_42_imag,
  output     [15:0]   sdata_out_payload_43_real,
  output     [15:0]   sdata_out_payload_43_imag,
  output     [15:0]   sdata_out_payload_44_real,
  output     [15:0]   sdata_out_payload_44_imag,
  output     [15:0]   sdata_out_payload_45_real,
  output     [15:0]   sdata_out_payload_45_imag,
  output     [15:0]   sdata_out_payload_46_real,
  output     [15:0]   sdata_out_payload_46_imag,
  output     [15:0]   sdata_out_payload_47_real,
  output     [15:0]   sdata_out_payload_47_imag,
  output     [15:0]   sdata_out_payload_48_real,
  output     [15:0]   sdata_out_payload_48_imag,
  output     [15:0]   sdata_out_payload_49_real,
  output     [15:0]   sdata_out_payload_49_imag,
  output     [15:0]   sdata_out_payload_50_real,
  output     [15:0]   sdata_out_payload_50_imag,
  output     [15:0]   sdata_out_payload_51_real,
  output     [15:0]   sdata_out_payload_51_imag,
  output     [15:0]   sdata_out_payload_52_real,
  output     [15:0]   sdata_out_payload_52_imag,
  output     [15:0]   sdata_out_payload_53_real,
  output     [15:0]   sdata_out_payload_53_imag,
  output     [15:0]   sdata_out_payload_54_real,
  output     [15:0]   sdata_out_payload_54_imag,
  output     [15:0]   sdata_out_payload_55_real,
  output     [15:0]   sdata_out_payload_55_imag,
  output     [15:0]   sdata_out_payload_56_real,
  output     [15:0]   sdata_out_payload_56_imag,
  output     [15:0]   sdata_out_payload_57_real,
  output     [15:0]   sdata_out_payload_57_imag,
  output     [15:0]   sdata_out_payload_58_real,
  output     [15:0]   sdata_out_payload_58_imag,
  output     [15:0]   sdata_out_payload_59_real,
  output     [15:0]   sdata_out_payload_59_imag,
  output     [15:0]   sdata_out_payload_60_real,
  output     [15:0]   sdata_out_payload_60_imag,
  output     [15:0]   sdata_out_payload_61_real,
  output     [15:0]   sdata_out_payload_61_imag,
  output     [15:0]   sdata_out_payload_62_real,
  output     [15:0]   sdata_out_payload_62_imag,
  output     [15:0]   sdata_out_payload_63_real,
  output     [15:0]   sdata_out_payload_63_imag,
  output     [15:0]   sdata_out_payload_64_real,
  output     [15:0]   sdata_out_payload_64_imag,
  output     [15:0]   sdata_out_payload_65_real,
  output     [15:0]   sdata_out_payload_65_imag,
  output     [15:0]   sdata_out_payload_66_real,
  output     [15:0]   sdata_out_payload_66_imag,
  output     [15:0]   sdata_out_payload_67_real,
  output     [15:0]   sdata_out_payload_67_imag,
  output     [15:0]   sdata_out_payload_68_real,
  output     [15:0]   sdata_out_payload_68_imag,
  output     [15:0]   sdata_out_payload_69_real,
  output     [15:0]   sdata_out_payload_69_imag,
  output     [15:0]   sdata_out_payload_70_real,
  output     [15:0]   sdata_out_payload_70_imag,
  output     [15:0]   sdata_out_payload_71_real,
  output     [15:0]   sdata_out_payload_71_imag,
  output     [15:0]   sdata_out_payload_72_real,
  output     [15:0]   sdata_out_payload_72_imag,
  output     [15:0]   sdata_out_payload_73_real,
  output     [15:0]   sdata_out_payload_73_imag,
  output     [15:0]   sdata_out_payload_74_real,
  output     [15:0]   sdata_out_payload_74_imag,
  output     [15:0]   sdata_out_payload_75_real,
  output     [15:0]   sdata_out_payload_75_imag,
  output     [15:0]   sdata_out_payload_76_real,
  output     [15:0]   sdata_out_payload_76_imag,
  output     [15:0]   sdata_out_payload_77_real,
  output     [15:0]   sdata_out_payload_77_imag,
  output     [15:0]   sdata_out_payload_78_real,
  output     [15:0]   sdata_out_payload_78_imag,
  output     [15:0]   sdata_out_payload_79_real,
  output     [15:0]   sdata_out_payload_79_imag,
  output     [15:0]   sdata_out_payload_80_real,
  output     [15:0]   sdata_out_payload_80_imag,
  output     [15:0]   sdata_out_payload_81_real,
  output     [15:0]   sdata_out_payload_81_imag,
  output     [15:0]   sdata_out_payload_82_real,
  output     [15:0]   sdata_out_payload_82_imag,
  output     [15:0]   sdata_out_payload_83_real,
  output     [15:0]   sdata_out_payload_83_imag,
  output     [15:0]   sdata_out_payload_84_real,
  output     [15:0]   sdata_out_payload_84_imag,
  output     [15:0]   sdata_out_payload_85_real,
  output     [15:0]   sdata_out_payload_85_imag,
  output     [15:0]   sdata_out_payload_86_real,
  output     [15:0]   sdata_out_payload_86_imag,
  output     [15:0]   sdata_out_payload_87_real,
  output     [15:0]   sdata_out_payload_87_imag,
  output     [15:0]   sdata_out_payload_88_real,
  output     [15:0]   sdata_out_payload_88_imag,
  output     [15:0]   sdata_out_payload_89_real,
  output     [15:0]   sdata_out_payload_89_imag,
  output     [15:0]   sdata_out_payload_90_real,
  output     [15:0]   sdata_out_payload_90_imag,
  output     [15:0]   sdata_out_payload_91_real,
  output     [15:0]   sdata_out_payload_91_imag,
  output     [15:0]   sdata_out_payload_92_real,
  output     [15:0]   sdata_out_payload_92_imag,
  output     [15:0]   sdata_out_payload_93_real,
  output     [15:0]   sdata_out_payload_93_imag,
  output     [15:0]   sdata_out_payload_94_real,
  output     [15:0]   sdata_out_payload_94_imag,
  output     [15:0]   sdata_out_payload_95_real,
  output     [15:0]   sdata_out_payload_95_imag,
  output     [15:0]   sdata_out_payload_96_real,
  output     [15:0]   sdata_out_payload_96_imag,
  output     [15:0]   sdata_out_payload_97_real,
  output     [15:0]   sdata_out_payload_97_imag,
  output     [15:0]   sdata_out_payload_98_real,
  output     [15:0]   sdata_out_payload_98_imag,
  output     [15:0]   sdata_out_payload_99_real,
  output     [15:0]   sdata_out_payload_99_imag,
  output     [15:0]   sdata_out_payload_100_real,
  output     [15:0]   sdata_out_payload_100_imag,
  output     [15:0]   sdata_out_payload_101_real,
  output     [15:0]   sdata_out_payload_101_imag,
  output     [15:0]   sdata_out_payload_102_real,
  output     [15:0]   sdata_out_payload_102_imag,
  output     [15:0]   sdata_out_payload_103_real,
  output     [15:0]   sdata_out_payload_103_imag,
  output     [15:0]   sdata_out_payload_104_real,
  output     [15:0]   sdata_out_payload_104_imag,
  output     [15:0]   sdata_out_payload_105_real,
  output     [15:0]   sdata_out_payload_105_imag,
  output     [15:0]   sdata_out_payload_106_real,
  output     [15:0]   sdata_out_payload_106_imag,
  output     [15:0]   sdata_out_payload_107_real,
  output     [15:0]   sdata_out_payload_107_imag,
  output     [15:0]   sdata_out_payload_108_real,
  output     [15:0]   sdata_out_payload_108_imag,
  output     [15:0]   sdata_out_payload_109_real,
  output     [15:0]   sdata_out_payload_109_imag,
  output     [15:0]   sdata_out_payload_110_real,
  output     [15:0]   sdata_out_payload_110_imag,
  output     [15:0]   sdata_out_payload_111_real,
  output     [15:0]   sdata_out_payload_111_imag,
  output     [15:0]   sdata_out_payload_112_real,
  output     [15:0]   sdata_out_payload_112_imag,
  output     [15:0]   sdata_out_payload_113_real,
  output     [15:0]   sdata_out_payload_113_imag,
  output     [15:0]   sdata_out_payload_114_real,
  output     [15:0]   sdata_out_payload_114_imag,
  output     [15:0]   sdata_out_payload_115_real,
  output     [15:0]   sdata_out_payload_115_imag,
  output     [15:0]   sdata_out_payload_116_real,
  output     [15:0]   sdata_out_payload_116_imag,
  output     [15:0]   sdata_out_payload_117_real,
  output     [15:0]   sdata_out_payload_117_imag,
  output     [15:0]   sdata_out_payload_118_real,
  output     [15:0]   sdata_out_payload_118_imag,
  output     [15:0]   sdata_out_payload_119_real,
  output     [15:0]   sdata_out_payload_119_imag,
  output     [15:0]   sdata_out_payload_120_real,
  output     [15:0]   sdata_out_payload_120_imag,
  output     [15:0]   sdata_out_payload_121_real,
  output     [15:0]   sdata_out_payload_121_imag,
  output     [15:0]   sdata_out_payload_122_real,
  output     [15:0]   sdata_out_payload_122_imag,
  output     [15:0]   sdata_out_payload_123_real,
  output     [15:0]   sdata_out_payload_123_imag,
  output     [15:0]   sdata_out_payload_124_real,
  output     [15:0]   sdata_out_payload_124_imag,
  output     [15:0]   sdata_out_payload_125_real,
  output     [15:0]   sdata_out_payload_125_imag,
  output     [15:0]   sdata_out_payload_126_real,
  output     [15:0]   sdata_out_payload_126_imag,
  output     [15:0]   sdata_out_payload_127_real,
  output     [15:0]   sdata_out_payload_127_imag,
  input               clk,
  input               reset
);
  wire       [31:0]   _zz_2241;
  wire       [31:0]   _zz_2242;
  wire       [31:0]   _zz_2243;
  wire       [31:0]   _zz_2244;
  wire       [31:0]   _zz_2245;
  wire       [31:0]   _zz_2246;
  wire       [31:0]   _zz_2247;
  wire       [31:0]   _zz_2248;
  wire       [31:0]   _zz_2249;
  wire       [31:0]   _zz_2250;
  wire       [31:0]   _zz_2251;
  wire       [31:0]   _zz_2252;
  wire       [31:0]   _zz_2253;
  wire       [31:0]   _zz_2254;
  wire       [31:0]   _zz_2255;
  wire       [31:0]   _zz_2256;
  wire       [31:0]   _zz_2257;
  wire       [31:0]   _zz_2258;
  wire       [31:0]   _zz_2259;
  wire       [31:0]   _zz_2260;
  wire       [31:0]   _zz_2261;
  wire       [31:0]   _zz_2262;
  wire       [31:0]   _zz_2263;
  wire       [31:0]   _zz_2264;
  wire       [31:0]   _zz_2265;
  wire       [31:0]   _zz_2266;
  wire       [31:0]   _zz_2267;
  wire       [31:0]   _zz_2268;
  wire       [31:0]   _zz_2269;
  wire       [31:0]   _zz_2270;
  wire       [31:0]   _zz_2271;
  wire       [31:0]   _zz_2272;
  wire       [31:0]   _zz_2273;
  wire       [31:0]   _zz_2274;
  wire       [31:0]   _zz_2275;
  wire       [31:0]   _zz_2276;
  wire       [31:0]   _zz_2277;
  wire       [31:0]   _zz_2278;
  wire       [31:0]   _zz_2279;
  wire       [31:0]   _zz_2280;
  wire       [31:0]   _zz_2281;
  wire       [31:0]   _zz_2282;
  wire       [31:0]   _zz_2283;
  wire       [31:0]   _zz_2284;
  wire       [31:0]   _zz_2285;
  wire       [31:0]   _zz_2286;
  wire       [31:0]   _zz_2287;
  wire       [31:0]   _zz_2288;
  wire       [31:0]   _zz_2289;
  wire       [31:0]   _zz_2290;
  wire       [31:0]   _zz_2291;
  wire       [31:0]   _zz_2292;
  wire       [31:0]   _zz_2293;
  wire       [31:0]   _zz_2294;
  wire       [31:0]   _zz_2295;
  wire       [31:0]   _zz_2296;
  wire       [31:0]   _zz_2297;
  wire       [31:0]   _zz_2298;
  wire       [31:0]   _zz_2299;
  wire       [31:0]   _zz_2300;
  wire       [31:0]   _zz_2301;
  wire       [31:0]   _zz_2302;
  wire       [31:0]   _zz_2303;
  wire       [31:0]   _zz_2304;
  wire       [31:0]   _zz_2305;
  wire       [31:0]   _zz_2306;
  wire       [31:0]   _zz_2307;
  wire       [31:0]   _zz_2308;
  wire       [31:0]   _zz_2309;
  wire       [31:0]   _zz_2310;
  wire       [31:0]   _zz_2311;
  wire       [31:0]   _zz_2312;
  wire       [31:0]   _zz_2313;
  wire       [31:0]   _zz_2314;
  wire       [31:0]   _zz_2315;
  wire       [31:0]   _zz_2316;
  wire       [31:0]   _zz_2317;
  wire       [31:0]   _zz_2318;
  wire       [31:0]   _zz_2319;
  wire       [31:0]   _zz_2320;
  wire       [31:0]   _zz_2321;
  wire       [31:0]   _zz_2322;
  wire       [31:0]   _zz_2323;
  wire       [31:0]   _zz_2324;
  wire       [31:0]   _zz_2325;
  wire       [31:0]   _zz_2326;
  wire       [31:0]   _zz_2327;
  wire       [31:0]   _zz_2328;
  wire       [31:0]   _zz_2329;
  wire       [31:0]   _zz_2330;
  wire       [31:0]   _zz_2331;
  wire       [31:0]   _zz_2332;
  wire       [31:0]   _zz_2333;
  wire       [31:0]   _zz_2334;
  wire       [31:0]   _zz_2335;
  wire       [31:0]   _zz_2336;
  wire       [31:0]   _zz_2337;
  wire       [31:0]   _zz_2338;
  wire       [31:0]   _zz_2339;
  wire       [31:0]   _zz_2340;
  wire       [31:0]   _zz_2341;
  wire       [31:0]   _zz_2342;
  wire       [31:0]   _zz_2343;
  wire       [31:0]   _zz_2344;
  wire       [31:0]   _zz_2345;
  wire       [31:0]   _zz_2346;
  wire       [31:0]   _zz_2347;
  wire       [31:0]   _zz_2348;
  wire       [31:0]   _zz_2349;
  wire       [31:0]   _zz_2350;
  wire       [31:0]   _zz_2351;
  wire       [31:0]   _zz_2352;
  wire       [31:0]   _zz_2353;
  wire       [31:0]   _zz_2354;
  wire       [31:0]   _zz_2355;
  wire       [31:0]   _zz_2356;
  wire       [31:0]   _zz_2357;
  wire       [31:0]   _zz_2358;
  wire       [31:0]   _zz_2359;
  wire       [31:0]   _zz_2360;
  wire       [31:0]   _zz_2361;
  wire       [31:0]   _zz_2362;
  wire       [31:0]   _zz_2363;
  wire       [31:0]   _zz_2364;
  wire       [31:0]   _zz_2365;
  wire       [31:0]   _zz_2366;
  wire       [31:0]   _zz_2367;
  wire       [31:0]   _zz_2368;
  wire       [31:0]   _zz_2369;
  wire       [31:0]   _zz_2370;
  wire       [31:0]   _zz_2371;
  wire       [31:0]   _zz_2372;
  wire       [31:0]   _zz_2373;
  wire       [31:0]   _zz_2374;
  wire       [31:0]   _zz_2375;
  wire       [31:0]   _zz_2376;
  wire       [31:0]   _zz_2377;
  wire       [31:0]   _zz_2378;
  wire       [31:0]   _zz_2379;
  wire       [31:0]   _zz_2380;
  wire       [31:0]   _zz_2381;
  wire       [31:0]   _zz_2382;
  wire       [31:0]   _zz_2383;
  wire       [31:0]   _zz_2384;
  wire       [31:0]   _zz_2385;
  wire       [31:0]   _zz_2386;
  wire       [31:0]   _zz_2387;
  wire       [31:0]   _zz_2388;
  wire       [31:0]   _zz_2389;
  wire       [31:0]   _zz_2390;
  wire       [31:0]   _zz_2391;
  wire       [31:0]   _zz_2392;
  wire       [31:0]   _zz_2393;
  wire       [31:0]   _zz_2394;
  wire       [31:0]   _zz_2395;
  wire       [31:0]   _zz_2396;
  wire       [31:0]   _zz_2397;
  wire       [31:0]   _zz_2398;
  wire       [31:0]   _zz_2399;
  wire       [31:0]   _zz_2400;
  wire       [31:0]   _zz_2401;
  wire       [31:0]   _zz_2402;
  wire       [31:0]   _zz_2403;
  wire       [31:0]   _zz_2404;
  wire       [31:0]   _zz_2405;
  wire       [31:0]   _zz_2406;
  wire       [31:0]   _zz_2407;
  wire       [31:0]   _zz_2408;
  wire       [31:0]   _zz_2409;
  wire       [31:0]   _zz_2410;
  wire       [31:0]   _zz_2411;
  wire       [31:0]   _zz_2412;
  wire       [31:0]   _zz_2413;
  wire       [31:0]   _zz_2414;
  wire       [31:0]   _zz_2415;
  wire       [31:0]   _zz_2416;
  wire       [31:0]   _zz_2417;
  wire       [31:0]   _zz_2418;
  wire       [31:0]   _zz_2419;
  wire       [31:0]   _zz_2420;
  wire       [31:0]   _zz_2421;
  wire       [31:0]   _zz_2422;
  wire       [31:0]   _zz_2423;
  wire       [31:0]   _zz_2424;
  wire       [31:0]   _zz_2425;
  wire       [31:0]   _zz_2426;
  wire       [31:0]   _zz_2427;
  wire       [31:0]   _zz_2428;
  wire       [31:0]   _zz_2429;
  wire       [31:0]   _zz_2430;
  wire       [31:0]   _zz_2431;
  wire       [31:0]   _zz_2432;
  wire       [31:0]   _zz_2433;
  wire       [31:0]   _zz_2434;
  wire       [31:0]   _zz_2435;
  wire       [31:0]   _zz_2436;
  wire       [31:0]   _zz_2437;
  wire       [31:0]   _zz_2438;
  wire       [31:0]   _zz_2439;
  wire       [31:0]   _zz_2440;
  wire       [31:0]   _zz_2441;
  wire       [31:0]   _zz_2442;
  wire       [31:0]   _zz_2443;
  wire       [31:0]   _zz_2444;
  wire       [31:0]   _zz_2445;
  wire       [31:0]   _zz_2446;
  wire       [31:0]   _zz_2447;
  wire       [31:0]   _zz_2448;
  wire       [31:0]   _zz_2449;
  wire       [31:0]   _zz_2450;
  wire       [31:0]   _zz_2451;
  wire       [31:0]   _zz_2452;
  wire       [31:0]   _zz_2453;
  wire       [31:0]   _zz_2454;
  wire       [31:0]   _zz_2455;
  wire       [31:0]   _zz_2456;
  wire       [31:0]   _zz_2457;
  wire       [31:0]   _zz_2458;
  wire       [31:0]   _zz_2459;
  wire       [31:0]   _zz_2460;
  wire       [31:0]   _zz_2461;
  wire       [31:0]   _zz_2462;
  wire       [31:0]   _zz_2463;
  wire       [31:0]   _zz_2464;
  wire       [31:0]   _zz_2465;
  wire       [31:0]   _zz_2466;
  wire       [31:0]   _zz_2467;
  wire       [31:0]   _zz_2468;
  wire       [31:0]   _zz_2469;
  wire       [31:0]   _zz_2470;
  wire       [31:0]   _zz_2471;
  wire       [31:0]   _zz_2472;
  wire       [31:0]   _zz_2473;
  wire       [31:0]   _zz_2474;
  wire       [31:0]   _zz_2475;
  wire       [31:0]   _zz_2476;
  wire       [31:0]   _zz_2477;
  wire       [31:0]   _zz_2478;
  wire       [31:0]   _zz_2479;
  wire       [31:0]   _zz_2480;
  wire       [31:0]   _zz_2481;
  wire       [31:0]   _zz_2482;
  wire       [31:0]   _zz_2483;
  wire       [31:0]   _zz_2484;
  wire       [31:0]   _zz_2485;
  wire       [31:0]   _zz_2486;
  wire       [31:0]   _zz_2487;
  wire       [31:0]   _zz_2488;
  wire       [31:0]   _zz_2489;
  wire       [31:0]   _zz_2490;
  wire       [31:0]   _zz_2491;
  wire       [31:0]   _zz_2492;
  wire       [31:0]   _zz_2493;
  wire       [31:0]   _zz_2494;
  wire       [31:0]   _zz_2495;
  wire       [31:0]   _zz_2496;
  wire       [31:0]   _zz_2497;
  wire       [31:0]   _zz_2498;
  wire       [31:0]   _zz_2499;
  wire       [31:0]   _zz_2500;
  wire       [31:0]   _zz_2501;
  wire       [31:0]   _zz_2502;
  wire       [31:0]   _zz_2503;
  wire       [31:0]   _zz_2504;
  wire       [31:0]   _zz_2505;
  wire       [31:0]   _zz_2506;
  wire       [31:0]   _zz_2507;
  wire       [31:0]   _zz_2508;
  wire       [31:0]   _zz_2509;
  wire       [31:0]   _zz_2510;
  wire       [31:0]   _zz_2511;
  wire       [31:0]   _zz_2512;
  wire       [31:0]   _zz_2513;
  wire       [31:0]   _zz_2514;
  wire       [31:0]   _zz_2515;
  wire       [31:0]   _zz_2516;
  wire       [31:0]   _zz_2517;
  wire       [31:0]   _zz_2518;
  wire       [31:0]   _zz_2519;
  wire       [31:0]   _zz_2520;
  wire       [31:0]   _zz_2521;
  wire       [31:0]   _zz_2522;
  wire       [31:0]   _zz_2523;
  wire       [31:0]   _zz_2524;
  wire       [31:0]   _zz_2525;
  wire       [31:0]   _zz_2526;
  wire       [31:0]   _zz_2527;
  wire       [31:0]   _zz_2528;
  wire       [31:0]   _zz_2529;
  wire       [31:0]   _zz_2530;
  wire       [31:0]   _zz_2531;
  wire       [31:0]   _zz_2532;
  wire       [31:0]   _zz_2533;
  wire       [31:0]   _zz_2534;
  wire       [31:0]   _zz_2535;
  wire       [31:0]   _zz_2536;
  wire       [31:0]   _zz_2537;
  wire       [31:0]   _zz_2538;
  wire       [31:0]   _zz_2539;
  wire       [31:0]   _zz_2540;
  wire       [31:0]   _zz_2541;
  wire       [31:0]   _zz_2542;
  wire       [31:0]   _zz_2543;
  wire       [31:0]   _zz_2544;
  wire       [31:0]   _zz_2545;
  wire       [31:0]   _zz_2546;
  wire       [31:0]   _zz_2547;
  wire       [31:0]   _zz_2548;
  wire       [31:0]   _zz_2549;
  wire       [31:0]   _zz_2550;
  wire       [31:0]   _zz_2551;
  wire       [31:0]   _zz_2552;
  wire       [31:0]   _zz_2553;
  wire       [31:0]   _zz_2554;
  wire       [31:0]   _zz_2555;
  wire       [31:0]   _zz_2556;
  wire       [31:0]   _zz_2557;
  wire       [31:0]   _zz_2558;
  wire       [31:0]   _zz_2559;
  wire       [31:0]   _zz_2560;
  wire       [31:0]   _zz_2561;
  wire       [31:0]   _zz_2562;
  wire       [31:0]   _zz_2563;
  wire       [31:0]   _zz_2564;
  wire       [31:0]   _zz_2565;
  wire       [31:0]   _zz_2566;
  wire       [31:0]   _zz_2567;
  wire       [31:0]   _zz_2568;
  wire       [31:0]   _zz_2569;
  wire       [31:0]   _zz_2570;
  wire       [31:0]   _zz_2571;
  wire       [31:0]   _zz_2572;
  wire       [31:0]   _zz_2573;
  wire       [31:0]   _zz_2574;
  wire       [31:0]   _zz_2575;
  wire       [31:0]   _zz_2576;
  wire       [31:0]   _zz_2577;
  wire       [31:0]   _zz_2578;
  wire       [31:0]   _zz_2579;
  wire       [31:0]   _zz_2580;
  wire       [31:0]   _zz_2581;
  wire       [31:0]   _zz_2582;
  wire       [31:0]   _zz_2583;
  wire       [31:0]   _zz_2584;
  wire       [31:0]   _zz_2585;
  wire       [31:0]   _zz_2586;
  wire       [31:0]   _zz_2587;
  wire       [31:0]   _zz_2588;
  wire       [31:0]   _zz_2589;
  wire       [31:0]   _zz_2590;
  wire       [31:0]   _zz_2591;
  wire       [31:0]   _zz_2592;
  wire       [31:0]   _zz_2593;
  wire       [31:0]   _zz_2594;
  wire       [31:0]   _zz_2595;
  wire       [31:0]   _zz_2596;
  wire       [31:0]   _zz_2597;
  wire       [31:0]   _zz_2598;
  wire       [31:0]   _zz_2599;
  wire       [31:0]   _zz_2600;
  wire       [31:0]   _zz_2601;
  wire       [31:0]   _zz_2602;
  wire       [31:0]   _zz_2603;
  wire       [31:0]   _zz_2604;
  wire       [31:0]   _zz_2605;
  wire       [31:0]   _zz_2606;
  wire       [31:0]   _zz_2607;
  wire       [31:0]   _zz_2608;
  wire       [31:0]   _zz_2609;
  wire       [31:0]   _zz_2610;
  wire       [31:0]   _zz_2611;
  wire       [31:0]   _zz_2612;
  wire       [31:0]   _zz_2613;
  wire       [31:0]   _zz_2614;
  wire       [31:0]   _zz_2615;
  wire       [31:0]   _zz_2616;
  wire       [31:0]   _zz_2617;
  wire       [31:0]   _zz_2618;
  wire       [31:0]   _zz_2619;
  wire       [31:0]   _zz_2620;
  wire       [31:0]   _zz_2621;
  wire       [31:0]   _zz_2622;
  wire       [31:0]   _zz_2623;
  wire       [31:0]   _zz_2624;
  wire       [31:0]   _zz_2625;
  wire       [31:0]   _zz_2626;
  wire       [31:0]   _zz_2627;
  wire       [31:0]   _zz_2628;
  wire       [31:0]   _zz_2629;
  wire       [31:0]   _zz_2630;
  wire       [31:0]   _zz_2631;
  wire       [31:0]   _zz_2632;
  wire       [31:0]   _zz_2633;
  wire       [31:0]   _zz_2634;
  wire       [31:0]   _zz_2635;
  wire       [31:0]   _zz_2636;
  wire       [31:0]   _zz_2637;
  wire       [31:0]   _zz_2638;
  wire       [31:0]   _zz_2639;
  wire       [31:0]   _zz_2640;
  wire       [31:0]   _zz_2641;
  wire       [31:0]   _zz_2642;
  wire       [31:0]   _zz_2643;
  wire       [31:0]   _zz_2644;
  wire       [31:0]   _zz_2645;
  wire       [31:0]   _zz_2646;
  wire       [31:0]   _zz_2647;
  wire       [31:0]   _zz_2648;
  wire       [31:0]   _zz_2649;
  wire       [31:0]   _zz_2650;
  wire       [31:0]   _zz_2651;
  wire       [31:0]   _zz_2652;
  wire       [31:0]   _zz_2653;
  wire       [31:0]   _zz_2654;
  wire       [31:0]   _zz_2655;
  wire       [31:0]   _zz_2656;
  wire       [31:0]   _zz_2657;
  wire       [31:0]   _zz_2658;
  wire       [31:0]   _zz_2659;
  wire       [31:0]   _zz_2660;
  wire       [31:0]   _zz_2661;
  wire       [31:0]   _zz_2662;
  wire       [31:0]   _zz_2663;
  wire       [31:0]   _zz_2664;
  wire       [31:0]   _zz_2665;
  wire       [31:0]   _zz_2666;
  wire       [31:0]   _zz_2667;
  wire       [31:0]   _zz_2668;
  wire       [31:0]   _zz_2669;
  wire       [31:0]   _zz_2670;
  wire       [31:0]   _zz_2671;
  wire       [31:0]   _zz_2672;
  wire       [31:0]   _zz_2673;
  wire       [31:0]   _zz_2674;
  wire       [31:0]   _zz_2675;
  wire       [31:0]   _zz_2676;
  wire       [31:0]   _zz_2677;
  wire       [31:0]   _zz_2678;
  wire       [31:0]   _zz_2679;
  wire       [31:0]   _zz_2680;
  wire       [31:0]   _zz_2681;
  wire       [31:0]   _zz_2682;
  wire       [31:0]   _zz_2683;
  wire       [31:0]   _zz_2684;
  wire       [31:0]   _zz_2685;
  wire       [31:0]   _zz_2686;
  wire       [31:0]   _zz_2687;
  wire       [31:0]   _zz_2688;
  wire       [31:0]   _zz_2689;
  wire       [31:0]   _zz_2690;
  wire       [31:0]   _zz_2691;
  wire       [31:0]   _zz_2692;
  wire       [31:0]   _zz_2693;
  wire       [31:0]   _zz_2694;
  wire       [31:0]   _zz_2695;
  wire       [31:0]   _zz_2696;
  wire       [31:0]   _zz_2697;
  wire       [31:0]   _zz_2698;
  wire       [31:0]   _zz_2699;
  wire       [31:0]   _zz_2700;
  wire       [31:0]   _zz_2701;
  wire       [31:0]   _zz_2702;
  wire       [31:0]   _zz_2703;
  wire       [31:0]   _zz_2704;
  wire       [31:0]   _zz_2705;
  wire       [31:0]   _zz_2706;
  wire       [31:0]   _zz_2707;
  wire       [31:0]   _zz_2708;
  wire       [31:0]   _zz_2709;
  wire       [31:0]   _zz_2710;
  wire       [31:0]   _zz_2711;
  wire       [31:0]   _zz_2712;
  wire       [31:0]   _zz_2713;
  wire       [31:0]   _zz_2714;
  wire       [31:0]   _zz_2715;
  wire       [31:0]   _zz_2716;
  wire       [31:0]   _zz_2717;
  wire       [31:0]   _zz_2718;
  wire       [31:0]   _zz_2719;
  wire       [31:0]   _zz_2720;
  wire       [31:0]   _zz_2721;
  wire       [31:0]   _zz_2722;
  wire       [31:0]   _zz_2723;
  wire       [31:0]   _zz_2724;
  wire       [31:0]   _zz_2725;
  wire       [31:0]   _zz_2726;
  wire       [31:0]   _zz_2727;
  wire       [31:0]   _zz_2728;
  wire       [31:0]   _zz_2729;
  wire       [31:0]   _zz_2730;
  wire       [31:0]   _zz_2731;
  wire       [31:0]   _zz_2732;
  wire       [31:0]   _zz_2733;
  wire       [31:0]   _zz_2734;
  wire       [31:0]   _zz_2735;
  wire       [31:0]   _zz_2736;
  wire       [31:0]   _zz_2737;
  wire       [31:0]   _zz_2738;
  wire       [31:0]   _zz_2739;
  wire       [31:0]   _zz_2740;
  wire       [31:0]   _zz_2741;
  wire       [31:0]   _zz_2742;
  wire       [31:0]   _zz_2743;
  wire       [31:0]   _zz_2744;
  wire       [31:0]   _zz_2745;
  wire       [31:0]   _zz_2746;
  wire       [31:0]   _zz_2747;
  wire       [31:0]   _zz_2748;
  wire       [31:0]   _zz_2749;
  wire       [31:0]   _zz_2750;
  wire       [31:0]   _zz_2751;
  wire       [31:0]   _zz_2752;
  wire       [31:0]   _zz_2753;
  wire       [31:0]   _zz_2754;
  wire       [31:0]   _zz_2755;
  wire       [31:0]   _zz_2756;
  wire       [31:0]   _zz_2757;
  wire       [31:0]   _zz_2758;
  wire       [31:0]   _zz_2759;
  wire       [31:0]   _zz_2760;
  wire       [31:0]   _zz_2761;
  wire       [31:0]   _zz_2762;
  wire       [31:0]   _zz_2763;
  wire       [31:0]   _zz_2764;
  wire       [31:0]   _zz_2765;
  wire       [31:0]   _zz_2766;
  wire       [31:0]   _zz_2767;
  wire       [31:0]   _zz_2768;
  wire       [31:0]   _zz_2769;
  wire       [31:0]   _zz_2770;
  wire       [31:0]   _zz_2771;
  wire       [31:0]   _zz_2772;
  wire       [31:0]   _zz_2773;
  wire       [31:0]   _zz_2774;
  wire       [31:0]   _zz_2775;
  wire       [31:0]   _zz_2776;
  wire       [31:0]   _zz_2777;
  wire       [31:0]   _zz_2778;
  wire       [31:0]   _zz_2779;
  wire       [31:0]   _zz_2780;
  wire       [31:0]   _zz_2781;
  wire       [31:0]   _zz_2782;
  wire       [31:0]   _zz_2783;
  wire       [31:0]   _zz_2784;
  wire       [31:0]   _zz_2785;
  wire       [31:0]   _zz_2786;
  wire       [31:0]   _zz_2787;
  wire       [31:0]   _zz_2788;
  wire       [31:0]   _zz_2789;
  wire       [31:0]   _zz_2790;
  wire       [31:0]   _zz_2791;
  wire       [31:0]   _zz_2792;
  wire       [31:0]   _zz_2793;
  wire       [31:0]   _zz_2794;
  wire       [31:0]   _zz_2795;
  wire       [31:0]   _zz_2796;
  wire       [31:0]   _zz_2797;
  wire       [31:0]   _zz_2798;
  wire       [31:0]   _zz_2799;
  wire       [31:0]   _zz_2800;
  wire       [31:0]   _zz_2801;
  wire       [31:0]   _zz_2802;
  wire       [31:0]   _zz_2803;
  wire       [31:0]   _zz_2804;
  wire       [31:0]   _zz_2805;
  wire       [31:0]   _zz_2806;
  wire       [31:0]   _zz_2807;
  wire       [31:0]   _zz_2808;
  wire       [31:0]   _zz_2809;
  wire       [31:0]   _zz_2810;
  wire       [31:0]   _zz_2811;
  wire       [31:0]   _zz_2812;
  wire       [31:0]   _zz_2813;
  wire       [31:0]   _zz_2814;
  wire       [31:0]   _zz_2815;
  wire       [31:0]   _zz_2816;
  wire       [31:0]   _zz_2817;
  wire       [31:0]   _zz_2818;
  wire       [31:0]   _zz_2819;
  wire       [31:0]   _zz_2820;
  wire       [31:0]   _zz_2821;
  wire       [31:0]   _zz_2822;
  wire       [31:0]   _zz_2823;
  wire       [31:0]   _zz_2824;
  wire       [31:0]   _zz_2825;
  wire       [31:0]   _zz_2826;
  wire       [31:0]   _zz_2827;
  wire       [31:0]   _zz_2828;
  wire       [31:0]   _zz_2829;
  wire       [31:0]   _zz_2830;
  wire       [31:0]   _zz_2831;
  wire       [31:0]   _zz_2832;
  wire       [31:0]   _zz_2833;
  wire       [31:0]   _zz_2834;
  wire       [31:0]   _zz_2835;
  wire       [31:0]   _zz_2836;
  wire       [31:0]   _zz_2837;
  wire       [31:0]   _zz_2838;
  wire       [31:0]   _zz_2839;
  wire       [31:0]   _zz_2840;
  wire       [31:0]   _zz_2841;
  wire       [31:0]   _zz_2842;
  wire       [31:0]   _zz_2843;
  wire       [31:0]   _zz_2844;
  wire       [31:0]   _zz_2845;
  wire       [31:0]   _zz_2846;
  wire       [31:0]   _zz_2847;
  wire       [31:0]   _zz_2848;
  wire       [31:0]   _zz_2849;
  wire       [31:0]   _zz_2850;
  wire       [31:0]   _zz_2851;
  wire       [31:0]   _zz_2852;
  wire       [31:0]   _zz_2853;
  wire       [31:0]   _zz_2854;
  wire       [31:0]   _zz_2855;
  wire       [31:0]   _zz_2856;
  wire       [31:0]   _zz_2857;
  wire       [31:0]   _zz_2858;
  wire       [31:0]   _zz_2859;
  wire       [31:0]   _zz_2860;
  wire       [31:0]   _zz_2861;
  wire       [31:0]   _zz_2862;
  wire       [31:0]   _zz_2863;
  wire       [31:0]   _zz_2864;
  wire       [31:0]   _zz_2865;
  wire       [31:0]   _zz_2866;
  wire       [31:0]   _zz_2867;
  wire       [31:0]   _zz_2868;
  wire       [31:0]   _zz_2869;
  wire       [31:0]   _zz_2870;
  wire       [31:0]   _zz_2871;
  wire       [31:0]   _zz_2872;
  wire       [31:0]   _zz_2873;
  wire       [31:0]   _zz_2874;
  wire       [31:0]   _zz_2875;
  wire       [31:0]   _zz_2876;
  wire       [31:0]   _zz_2877;
  wire       [31:0]   _zz_2878;
  wire       [31:0]   _zz_2879;
  wire       [31:0]   _zz_2880;
  wire       [31:0]   _zz_2881;
  wire       [31:0]   _zz_2882;
  wire       [31:0]   _zz_2883;
  wire       [31:0]   _zz_2884;
  wire       [31:0]   _zz_2885;
  wire       [31:0]   _zz_2886;
  wire       [31:0]   _zz_2887;
  wire       [31:0]   _zz_2888;
  wire       [31:0]   _zz_2889;
  wire       [31:0]   _zz_2890;
  wire       [31:0]   _zz_2891;
  wire       [31:0]   _zz_2892;
  wire       [31:0]   _zz_2893;
  wire       [31:0]   _zz_2894;
  wire       [31:0]   _zz_2895;
  wire       [31:0]   _zz_2896;
  wire       [31:0]   _zz_2897;
  wire       [31:0]   _zz_2898;
  wire       [31:0]   _zz_2899;
  wire       [31:0]   _zz_2900;
  wire       [31:0]   _zz_2901;
  wire       [31:0]   _zz_2902;
  wire       [31:0]   _zz_2903;
  wire       [31:0]   _zz_2904;
  wire       [31:0]   _zz_2905;
  wire       [31:0]   _zz_2906;
  wire       [31:0]   _zz_2907;
  wire       [31:0]   _zz_2908;
  wire       [31:0]   _zz_2909;
  wire       [31:0]   _zz_2910;
  wire       [31:0]   _zz_2911;
  wire       [31:0]   _zz_2912;
  wire       [31:0]   _zz_2913;
  wire       [31:0]   _zz_2914;
  wire       [31:0]   _zz_2915;
  wire       [31:0]   _zz_2916;
  wire       [31:0]   _zz_2917;
  wire       [31:0]   _zz_2918;
  wire       [31:0]   _zz_2919;
  wire       [31:0]   _zz_2920;
  wire       [31:0]   _zz_2921;
  wire       [31:0]   _zz_2922;
  wire       [31:0]   _zz_2923;
  wire       [31:0]   _zz_2924;
  wire       [31:0]   _zz_2925;
  wire       [31:0]   _zz_2926;
  wire       [31:0]   _zz_2927;
  wire       [31:0]   _zz_2928;
  wire       [31:0]   _zz_2929;
  wire       [31:0]   _zz_2930;
  wire       [31:0]   _zz_2931;
  wire       [31:0]   _zz_2932;
  wire       [31:0]   _zz_2933;
  wire       [31:0]   _zz_2934;
  wire       [31:0]   _zz_2935;
  wire       [31:0]   _zz_2936;
  wire       [31:0]   _zz_2937;
  wire       [31:0]   _zz_2938;
  wire       [31:0]   _zz_2939;
  wire       [31:0]   _zz_2940;
  wire       [31:0]   _zz_2941;
  wire       [31:0]   _zz_2942;
  wire       [31:0]   _zz_2943;
  wire       [31:0]   _zz_2944;
  wire       [31:0]   _zz_2945;
  wire       [31:0]   _zz_2946;
  wire       [31:0]   _zz_2947;
  wire       [31:0]   _zz_2948;
  wire       [31:0]   _zz_2949;
  wire       [31:0]   _zz_2950;
  wire       [31:0]   _zz_2951;
  wire       [31:0]   _zz_2952;
  wire       [31:0]   _zz_2953;
  wire       [31:0]   _zz_2954;
  wire       [31:0]   _zz_2955;
  wire       [31:0]   _zz_2956;
  wire       [31:0]   _zz_2957;
  wire       [31:0]   _zz_2958;
  wire       [31:0]   _zz_2959;
  wire       [31:0]   _zz_2960;
  wire       [31:0]   _zz_2961;
  wire       [31:0]   _zz_2962;
  wire       [31:0]   _zz_2963;
  wire       [31:0]   _zz_2964;
  wire       [31:0]   _zz_2965;
  wire       [31:0]   _zz_2966;
  wire       [31:0]   _zz_2967;
  wire       [31:0]   _zz_2968;
  wire       [31:0]   _zz_2969;
  wire       [31:0]   _zz_2970;
  wire       [31:0]   _zz_2971;
  wire       [31:0]   _zz_2972;
  wire       [31:0]   _zz_2973;
  wire       [31:0]   _zz_2974;
  wire       [31:0]   _zz_2975;
  wire       [31:0]   _zz_2976;
  wire       [31:0]   _zz_2977;
  wire       [31:0]   _zz_2978;
  wire       [31:0]   _zz_2979;
  wire       [31:0]   _zz_2980;
  wire       [31:0]   _zz_2981;
  wire       [31:0]   _zz_2982;
  wire       [31:0]   _zz_2983;
  wire       [31:0]   _zz_2984;
  wire       [31:0]   _zz_2985;
  wire       [31:0]   _zz_2986;
  wire       [31:0]   _zz_2987;
  wire       [31:0]   _zz_2988;
  wire       [31:0]   _zz_2989;
  wire       [31:0]   _zz_2990;
  wire       [31:0]   _zz_2991;
  wire       [31:0]   _zz_2992;
  wire       [31:0]   _zz_2993;
  wire       [31:0]   _zz_2994;
  wire       [31:0]   _zz_2995;
  wire       [31:0]   _zz_2996;
  wire       [31:0]   _zz_2997;
  wire       [31:0]   _zz_2998;
  wire       [31:0]   _zz_2999;
  wire       [31:0]   _zz_3000;
  wire       [31:0]   _zz_3001;
  wire       [31:0]   _zz_3002;
  wire       [31:0]   _zz_3003;
  wire       [31:0]   _zz_3004;
  wire       [31:0]   _zz_3005;
  wire       [31:0]   _zz_3006;
  wire       [31:0]   _zz_3007;
  wire       [31:0]   _zz_3008;
  wire       [31:0]   _zz_3009;
  wire       [31:0]   _zz_3010;
  wire       [31:0]   _zz_3011;
  wire       [31:0]   _zz_3012;
  wire       [31:0]   _zz_3013;
  wire       [31:0]   _zz_3014;
  wire       [31:0]   _zz_3015;
  wire       [31:0]   _zz_3016;
  wire       [31:0]   _zz_3017;
  wire       [31:0]   _zz_3018;
  wire       [31:0]   _zz_3019;
  wire       [31:0]   _zz_3020;
  wire       [31:0]   _zz_3021;
  wire       [31:0]   _zz_3022;
  wire       [31:0]   _zz_3023;
  wire       [31:0]   _zz_3024;
  wire       [31:0]   _zz_3025;
  wire       [31:0]   _zz_3026;
  wire       [31:0]   _zz_3027;
  wire       [31:0]   _zz_3028;
  wire       [31:0]   _zz_3029;
  wire       [31:0]   _zz_3030;
  wire       [31:0]   _zz_3031;
  wire       [31:0]   _zz_3032;
  wire       [31:0]   _zz_3033;
  wire       [31:0]   _zz_3034;
  wire       [31:0]   _zz_3035;
  wire       [31:0]   _zz_3036;
  wire       [31:0]   _zz_3037;
  wire       [31:0]   _zz_3038;
  wire       [31:0]   _zz_3039;
  wire       [31:0]   _zz_3040;
  wire       [31:0]   _zz_3041;
  wire       [31:0]   _zz_3042;
  wire       [31:0]   _zz_3043;
  wire       [31:0]   _zz_3044;
  wire       [31:0]   _zz_3045;
  wire       [31:0]   _zz_3046;
  wire       [31:0]   _zz_3047;
  wire       [31:0]   _zz_3048;
  wire       [31:0]   _zz_3049;
  wire       [31:0]   _zz_3050;
  wire       [31:0]   _zz_3051;
  wire       [31:0]   _zz_3052;
  wire       [31:0]   _zz_3053;
  wire       [31:0]   _zz_3054;
  wire       [31:0]   _zz_3055;
  wire       [31:0]   _zz_3056;
  wire       [31:0]   _zz_3057;
  wire       [31:0]   _zz_3058;
  wire       [31:0]   _zz_3059;
  wire       [31:0]   _zz_3060;
  wire       [31:0]   _zz_3061;
  wire       [31:0]   _zz_3062;
  wire       [31:0]   _zz_3063;
  wire       [31:0]   _zz_3064;
  wire       [31:0]   _zz_3065;
  wire       [31:0]   _zz_3066;
  wire       [31:0]   _zz_3067;
  wire       [31:0]   _zz_3068;
  wire       [31:0]   _zz_3069;
  wire       [31:0]   _zz_3070;
  wire       [31:0]   _zz_3071;
  wire       [31:0]   _zz_3072;
  wire       [31:0]   _zz_3073;
  wire       [31:0]   _zz_3074;
  wire       [31:0]   _zz_3075;
  wire       [31:0]   _zz_3076;
  wire       [31:0]   _zz_3077;
  wire       [31:0]   _zz_3078;
  wire       [31:0]   _zz_3079;
  wire       [31:0]   _zz_3080;
  wire       [31:0]   _zz_3081;
  wire       [31:0]   _zz_3082;
  wire       [31:0]   _zz_3083;
  wire       [31:0]   _zz_3084;
  wire       [31:0]   _zz_3085;
  wire       [31:0]   _zz_3086;
  wire       [31:0]   _zz_3087;
  wire       [31:0]   _zz_3088;
  wire       [31:0]   _zz_3089;
  wire       [31:0]   _zz_3090;
  wire       [31:0]   _zz_3091;
  wire       [31:0]   _zz_3092;
  wire       [31:0]   _zz_3093;
  wire       [31:0]   _zz_3094;
  wire       [31:0]   _zz_3095;
  wire       [31:0]   _zz_3096;
  wire       [31:0]   _zz_3097;
  wire       [31:0]   _zz_3098;
  wire       [31:0]   _zz_3099;
  wire       [31:0]   _zz_3100;
  wire       [31:0]   _zz_3101;
  wire       [31:0]   _zz_3102;
  wire       [31:0]   _zz_3103;
  wire       [31:0]   _zz_3104;
  wire       [31:0]   _zz_3105;
  wire       [31:0]   _zz_3106;
  wire       [31:0]   _zz_3107;
  wire       [31:0]   _zz_3108;
  wire       [31:0]   _zz_3109;
  wire       [31:0]   _zz_3110;
  wire       [31:0]   _zz_3111;
  wire       [31:0]   _zz_3112;
  wire       [31:0]   _zz_3113;
  wire       [31:0]   _zz_3114;
  wire       [31:0]   _zz_3115;
  wire       [31:0]   _zz_3116;
  wire       [31:0]   _zz_3117;
  wire       [31:0]   _zz_3118;
  wire       [31:0]   _zz_3119;
  wire       [31:0]   _zz_3120;
  wire       [31:0]   _zz_3121;
  wire       [31:0]   _zz_3122;
  wire       [31:0]   _zz_3123;
  wire       [31:0]   _zz_3124;
  wire       [31:0]   _zz_3125;
  wire       [31:0]   _zz_3126;
  wire       [31:0]   _zz_3127;
  wire       [31:0]   _zz_3128;
  wire       [31:0]   _zz_3129;
  wire       [31:0]   _zz_3130;
  wire       [31:0]   _zz_3131;
  wire       [31:0]   _zz_3132;
  wire       [31:0]   _zz_3133;
  wire       [31:0]   _zz_3134;
  wire       [31:0]   _zz_3135;
  wire       [31:0]   _zz_3136;
  wire       [31:0]   _zz_3137;
  wire       [31:0]   _zz_3138;
  wire       [31:0]   _zz_3139;
  wire       [31:0]   _zz_3140;
  wire       [31:0]   _zz_3141;
  wire       [31:0]   _zz_3142;
  wire       [31:0]   _zz_3143;
  wire       [31:0]   _zz_3144;
  wire       [31:0]   _zz_3145;
  wire       [31:0]   _zz_3146;
  wire       [31:0]   _zz_3147;
  wire       [31:0]   _zz_3148;
  wire       [31:0]   _zz_3149;
  wire       [31:0]   _zz_3150;
  wire       [31:0]   _zz_3151;
  wire       [31:0]   _zz_3152;
  wire       [31:0]   _zz_3153;
  wire       [31:0]   _zz_3154;
  wire       [31:0]   _zz_3155;
  wire       [31:0]   _zz_3156;
  wire       [31:0]   _zz_3157;
  wire       [31:0]   _zz_3158;
  wire       [31:0]   _zz_3159;
  wire       [31:0]   _zz_3160;
  wire       [31:0]   _zz_3161;
  wire       [31:0]   _zz_3162;
  wire       [31:0]   _zz_3163;
  wire       [31:0]   _zz_3164;
  wire       [31:0]   _zz_3165;
  wire       [31:0]   _zz_3166;
  wire       [31:0]   _zz_3167;
  wire       [31:0]   _zz_3168;
  wire       [31:0]   _zz_3169;
  wire       [31:0]   _zz_3170;
  wire       [31:0]   _zz_3171;
  wire       [31:0]   _zz_3172;
  wire       [31:0]   _zz_3173;
  wire       [31:0]   _zz_3174;
  wire       [31:0]   _zz_3175;
  wire       [31:0]   _zz_3176;
  wire       [31:0]   _zz_3177;
  wire       [31:0]   _zz_3178;
  wire       [31:0]   _zz_3179;
  wire       [31:0]   _zz_3180;
  wire       [31:0]   _zz_3181;
  wire       [31:0]   _zz_3182;
  wire       [31:0]   _zz_3183;
  wire       [31:0]   _zz_3184;
  wire       [31:0]   _zz_3185;
  wire       [31:0]   _zz_3186;
  wire       [31:0]   _zz_3187;
  wire       [31:0]   _zz_3188;
  wire       [31:0]   _zz_3189;
  wire       [31:0]   _zz_3190;
  wire       [31:0]   _zz_3191;
  wire       [31:0]   _zz_3192;
  wire       [31:0]   _zz_3193;
  wire       [31:0]   _zz_3194;
  wire       [31:0]   _zz_3195;
  wire       [31:0]   _zz_3196;
  wire       [31:0]   _zz_3197;
  wire       [31:0]   _zz_3198;
  wire       [31:0]   _zz_3199;
  wire       [31:0]   _zz_3200;
  wire       [31:0]   _zz_3201;
  wire       [31:0]   _zz_3202;
  wire       [31:0]   _zz_3203;
  wire       [31:0]   _zz_3204;
  wire       [31:0]   _zz_3205;
  wire       [31:0]   _zz_3206;
  wire       [31:0]   _zz_3207;
  wire       [31:0]   _zz_3208;
  wire       [31:0]   _zz_3209;
  wire       [31:0]   _zz_3210;
  wire       [31:0]   _zz_3211;
  wire       [31:0]   _zz_3212;
  wire       [31:0]   _zz_3213;
  wire       [31:0]   _zz_3214;
  wire       [31:0]   _zz_3215;
  wire       [31:0]   _zz_3216;
  wire       [31:0]   _zz_3217;
  wire       [31:0]   _zz_3218;
  wire       [31:0]   _zz_3219;
  wire       [31:0]   _zz_3220;
  wire       [31:0]   _zz_3221;
  wire       [31:0]   _zz_3222;
  wire       [31:0]   _zz_3223;
  wire       [31:0]   _zz_3224;
  wire       [31:0]   _zz_3225;
  wire       [31:0]   _zz_3226;
  wire       [31:0]   _zz_3227;
  wire       [31:0]   _zz_3228;
  wire       [31:0]   _zz_3229;
  wire       [31:0]   _zz_3230;
  wire       [31:0]   _zz_3231;
  wire       [31:0]   _zz_3232;
  wire       [31:0]   _zz_3233;
  wire       [31:0]   _zz_3234;
  wire       [31:0]   _zz_3235;
  wire       [31:0]   _zz_3236;
  wire       [31:0]   _zz_3237;
  wire       [31:0]   _zz_3238;
  wire       [31:0]   _zz_3239;
  wire       [31:0]   _zz_3240;
  wire       [31:0]   _zz_3241;
  wire       [31:0]   _zz_3242;
  wire       [31:0]   _zz_3243;
  wire       [31:0]   _zz_3244;
  wire       [31:0]   _zz_3245;
  wire       [31:0]   _zz_3246;
  wire       [31:0]   _zz_3247;
  wire       [31:0]   _zz_3248;
  wire       [31:0]   _zz_3249;
  wire       [31:0]   _zz_3250;
  wire       [31:0]   _zz_3251;
  wire       [31:0]   _zz_3252;
  wire       [31:0]   _zz_3253;
  wire       [31:0]   _zz_3254;
  wire       [31:0]   _zz_3255;
  wire       [31:0]   _zz_3256;
  wire       [31:0]   _zz_3257;
  wire       [31:0]   _zz_3258;
  wire       [31:0]   _zz_3259;
  wire       [31:0]   _zz_3260;
  wire       [31:0]   _zz_3261;
  wire       [31:0]   _zz_3262;
  wire       [31:0]   _zz_3263;
  wire       [31:0]   _zz_3264;
  wire       [31:0]   _zz_3265;
  wire       [31:0]   _zz_3266;
  wire       [31:0]   _zz_3267;
  wire       [31:0]   _zz_3268;
  wire       [31:0]   _zz_3269;
  wire       [31:0]   _zz_3270;
  wire       [31:0]   _zz_3271;
  wire       [31:0]   _zz_3272;
  wire       [31:0]   _zz_3273;
  wire       [31:0]   _zz_3274;
  wire       [31:0]   _zz_3275;
  wire       [31:0]   _zz_3276;
  wire       [31:0]   _zz_3277;
  wire       [31:0]   _zz_3278;
  wire       [31:0]   _zz_3279;
  wire       [31:0]   _zz_3280;
  wire       [31:0]   _zz_3281;
  wire       [31:0]   _zz_3282;
  wire       [31:0]   _zz_3283;
  wire       [31:0]   _zz_3284;
  wire       [31:0]   _zz_3285;
  wire       [31:0]   _zz_3286;
  wire       [31:0]   _zz_3287;
  wire       [31:0]   _zz_3288;
  wire       [31:0]   _zz_3289;
  wire       [31:0]   _zz_3290;
  wire       [31:0]   _zz_3291;
  wire       [31:0]   _zz_3292;
  wire       [31:0]   _zz_3293;
  wire       [31:0]   _zz_3294;
  wire       [31:0]   _zz_3295;
  wire       [31:0]   _zz_3296;
  wire       [31:0]   _zz_3297;
  wire       [31:0]   _zz_3298;
  wire       [31:0]   _zz_3299;
  wire       [31:0]   _zz_3300;
  wire       [31:0]   _zz_3301;
  wire       [31:0]   _zz_3302;
  wire       [31:0]   _zz_3303;
  wire       [31:0]   _zz_3304;
  wire       [31:0]   _zz_3305;
  wire       [31:0]   _zz_3306;
  wire       [31:0]   _zz_3307;
  wire       [31:0]   _zz_3308;
  wire       [31:0]   _zz_3309;
  wire       [31:0]   _zz_3310;
  wire       [31:0]   _zz_3311;
  wire       [31:0]   _zz_3312;
  wire       [31:0]   _zz_3313;
  wire       [31:0]   _zz_3314;
  wire       [31:0]   _zz_3315;
  wire       [31:0]   _zz_3316;
  wire       [31:0]   _zz_3317;
  wire       [31:0]   _zz_3318;
  wire       [31:0]   _zz_3319;
  wire       [31:0]   _zz_3320;
  wire       [31:0]   _zz_3321;
  wire       [31:0]   _zz_3322;
  wire       [31:0]   _zz_3323;
  wire       [31:0]   _zz_3324;
  wire       [31:0]   _zz_3325;
  wire       [31:0]   _zz_3326;
  wire       [31:0]   _zz_3327;
  wire       [31:0]   _zz_3328;
  wire       [31:0]   _zz_3329;
  wire       [31:0]   _zz_3330;
  wire       [31:0]   _zz_3331;
  wire       [31:0]   _zz_3332;
  wire       [31:0]   _zz_3333;
  wire       [31:0]   _zz_3334;
  wire       [31:0]   _zz_3335;
  wire       [31:0]   _zz_3336;
  wire       [31:0]   _zz_3337;
  wire       [31:0]   _zz_3338;
  wire       [31:0]   _zz_3339;
  wire       [31:0]   _zz_3340;
  wire       [31:0]   _zz_3341;
  wire       [31:0]   _zz_3342;
  wire       [31:0]   _zz_3343;
  wire       [31:0]   _zz_3344;
  wire       [31:0]   _zz_3345;
  wire       [31:0]   _zz_3346;
  wire       [31:0]   _zz_3347;
  wire       [31:0]   _zz_3348;
  wire       [31:0]   _zz_3349;
  wire       [31:0]   _zz_3350;
  wire       [31:0]   _zz_3351;
  wire       [31:0]   _zz_3352;
  wire       [31:0]   _zz_3353;
  wire       [31:0]   _zz_3354;
  wire       [31:0]   _zz_3355;
  wire       [31:0]   _zz_3356;
  wire       [31:0]   _zz_3357;
  wire       [31:0]   _zz_3358;
  wire       [31:0]   _zz_3359;
  wire       [31:0]   _zz_3360;
  wire       [31:0]   _zz_3361;
  wire       [31:0]   _zz_3362;
  wire       [31:0]   _zz_3363;
  wire       [31:0]   _zz_3364;
  wire       [31:0]   _zz_3365;
  wire       [31:0]   _zz_3366;
  wire       [31:0]   _zz_3367;
  wire       [31:0]   _zz_3368;
  wire       [31:0]   _zz_3369;
  wire       [31:0]   _zz_3370;
  wire       [31:0]   _zz_3371;
  wire       [31:0]   _zz_3372;
  wire       [31:0]   _zz_3373;
  wire       [31:0]   _zz_3374;
  wire       [31:0]   _zz_3375;
  wire       [31:0]   _zz_3376;
  wire       [31:0]   _zz_3377;
  wire       [31:0]   _zz_3378;
  wire       [31:0]   _zz_3379;
  wire       [31:0]   _zz_3380;
  wire       [31:0]   _zz_3381;
  wire       [31:0]   _zz_3382;
  wire       [31:0]   _zz_3383;
  wire       [31:0]   _zz_3384;
  wire       [31:0]   _zz_3385;
  wire       [31:0]   _zz_3386;
  wire       [31:0]   _zz_3387;
  wire       [31:0]   _zz_3388;
  wire       [31:0]   _zz_3389;
  wire       [31:0]   _zz_3390;
  wire       [31:0]   _zz_3391;
  wire       [31:0]   _zz_3392;
  wire       [31:0]   _zz_3393;
  wire       [31:0]   _zz_3394;
  wire       [31:0]   _zz_3395;
  wire       [31:0]   _zz_3396;
  wire       [31:0]   _zz_3397;
  wire       [31:0]   _zz_3398;
  wire       [31:0]   _zz_3399;
  wire       [31:0]   _zz_3400;
  wire       [31:0]   _zz_3401;
  wire       [31:0]   _zz_3402;
  wire       [31:0]   _zz_3403;
  wire       [31:0]   _zz_3404;
  wire       [31:0]   _zz_3405;
  wire       [31:0]   _zz_3406;
  wire       [31:0]   _zz_3407;
  wire       [31:0]   _zz_3408;
  wire       [31:0]   _zz_3409;
  wire       [31:0]   _zz_3410;
  wire       [31:0]   _zz_3411;
  wire       [31:0]   _zz_3412;
  wire       [31:0]   _zz_3413;
  wire       [31:0]   _zz_3414;
  wire       [31:0]   _zz_3415;
  wire       [31:0]   _zz_3416;
  wire       [31:0]   _zz_3417;
  wire       [31:0]   _zz_3418;
  wire       [31:0]   _zz_3419;
  wire       [31:0]   _zz_3420;
  wire       [31:0]   _zz_3421;
  wire       [31:0]   _zz_3422;
  wire       [31:0]   _zz_3423;
  wire       [31:0]   _zz_3424;
  wire       [31:0]   _zz_3425;
  wire       [31:0]   _zz_3426;
  wire       [31:0]   _zz_3427;
  wire       [31:0]   _zz_3428;
  wire       [31:0]   _zz_3429;
  wire       [31:0]   _zz_3430;
  wire       [31:0]   _zz_3431;
  wire       [31:0]   _zz_3432;
  wire       [31:0]   _zz_3433;
  wire       [31:0]   _zz_3434;
  wire       [31:0]   _zz_3435;
  wire       [31:0]   _zz_3436;
  wire       [31:0]   _zz_3437;
  wire       [31:0]   _zz_3438;
  wire       [31:0]   _zz_3439;
  wire       [31:0]   _zz_3440;
  wire       [31:0]   _zz_3441;
  wire       [31:0]   _zz_3442;
  wire       [31:0]   _zz_3443;
  wire       [31:0]   _zz_3444;
  wire       [31:0]   _zz_3445;
  wire       [31:0]   _zz_3446;
  wire       [31:0]   _zz_3447;
  wire       [31:0]   _zz_3448;
  wire       [31:0]   _zz_3449;
  wire       [31:0]   _zz_3450;
  wire       [31:0]   _zz_3451;
  wire       [31:0]   _zz_3452;
  wire       [31:0]   _zz_3453;
  wire       [31:0]   _zz_3454;
  wire       [31:0]   _zz_3455;
  wire       [31:0]   _zz_3456;
  wire       [31:0]   _zz_3457;
  wire       [31:0]   _zz_3458;
  wire       [31:0]   _zz_3459;
  wire       [31:0]   _zz_3460;
  wire       [31:0]   _zz_3461;
  wire       [31:0]   _zz_3462;
  wire       [31:0]   _zz_3463;
  wire       [31:0]   _zz_3464;
  wire       [31:0]   _zz_3465;
  wire       [31:0]   _zz_3466;
  wire       [31:0]   _zz_3467;
  wire       [31:0]   _zz_3468;
  wire       [31:0]   _zz_3469;
  wire       [31:0]   _zz_3470;
  wire       [31:0]   _zz_3471;
  wire       [31:0]   _zz_3472;
  wire       [31:0]   _zz_3473;
  wire       [31:0]   _zz_3474;
  wire       [31:0]   _zz_3475;
  wire       [31:0]   _zz_3476;
  wire       [31:0]   _zz_3477;
  wire       [31:0]   _zz_3478;
  wire       [31:0]   _zz_3479;
  wire       [31:0]   _zz_3480;
  wire       [31:0]   _zz_3481;
  wire       [31:0]   _zz_3482;
  wire       [31:0]   _zz_3483;
  wire       [31:0]   _zz_3484;
  wire       [31:0]   _zz_3485;
  wire       [31:0]   _zz_3486;
  wire       [31:0]   _zz_3487;
  wire       [31:0]   _zz_3488;
  wire       [31:0]   _zz_3489;
  wire       [31:0]   _zz_3490;
  wire       [31:0]   _zz_3491;
  wire       [31:0]   _zz_3492;
  wire       [31:0]   _zz_3493;
  wire       [31:0]   _zz_3494;
  wire       [31:0]   _zz_3495;
  wire       [31:0]   _zz_3496;
  wire       [31:0]   _zz_3497;
  wire       [31:0]   _zz_3498;
  wire       [31:0]   _zz_3499;
  wire       [31:0]   _zz_3500;
  wire       [31:0]   _zz_3501;
  wire       [31:0]   _zz_3502;
  wire       [31:0]   _zz_3503;
  wire       [31:0]   _zz_3504;
  wire       [31:0]   _zz_3505;
  wire       [31:0]   _zz_3506;
  wire       [31:0]   _zz_3507;
  wire       [31:0]   _zz_3508;
  wire       [31:0]   _zz_3509;
  wire       [31:0]   _zz_3510;
  wire       [31:0]   _zz_3511;
  wire       [31:0]   _zz_3512;
  wire       [31:0]   _zz_3513;
  wire       [31:0]   _zz_3514;
  wire       [31:0]   _zz_3515;
  wire       [31:0]   _zz_3516;
  wire       [31:0]   _zz_3517;
  wire       [31:0]   _zz_3518;
  wire       [31:0]   _zz_3519;
  wire       [31:0]   _zz_3520;
  wire       [31:0]   _zz_3521;
  wire       [31:0]   _zz_3522;
  wire       [31:0]   _zz_3523;
  wire       [31:0]   _zz_3524;
  wire       [31:0]   _zz_3525;
  wire       [31:0]   _zz_3526;
  wire       [31:0]   _zz_3527;
  wire       [31:0]   _zz_3528;
  wire       [31:0]   _zz_3529;
  wire       [31:0]   _zz_3530;
  wire       [31:0]   _zz_3531;
  wire       [31:0]   _zz_3532;
  wire       [31:0]   _zz_3533;
  wire       [31:0]   _zz_3534;
  wire       [31:0]   _zz_3535;
  wire       [31:0]   _zz_3536;
  wire       [31:0]   _zz_3537;
  wire       [31:0]   _zz_3538;
  wire       [31:0]   _zz_3539;
  wire       [31:0]   _zz_3540;
  wire       [31:0]   _zz_3541;
  wire       [31:0]   _zz_3542;
  wire       [31:0]   _zz_3543;
  wire       [31:0]   _zz_3544;
  wire       [31:0]   _zz_3545;
  wire       [31:0]   _zz_3546;
  wire       [31:0]   _zz_3547;
  wire       [31:0]   _zz_3548;
  wire       [31:0]   _zz_3549;
  wire       [31:0]   _zz_3550;
  wire       [31:0]   _zz_3551;
  wire       [31:0]   _zz_3552;
  wire       [31:0]   _zz_3553;
  wire       [31:0]   _zz_3554;
  wire       [31:0]   _zz_3555;
  wire       [31:0]   _zz_3556;
  wire       [31:0]   _zz_3557;
  wire       [31:0]   _zz_3558;
  wire       [31:0]   _zz_3559;
  wire       [31:0]   _zz_3560;
  wire       [31:0]   _zz_3561;
  wire       [31:0]   _zz_3562;
  wire       [31:0]   _zz_3563;
  wire       [31:0]   _zz_3564;
  wire       [31:0]   _zz_3565;
  wire       [31:0]   _zz_3566;
  wire       [31:0]   _zz_3567;
  wire       [31:0]   _zz_3568;
  wire       [31:0]   _zz_3569;
  wire       [31:0]   _zz_3570;
  wire       [31:0]   _zz_3571;
  wire       [31:0]   _zz_3572;
  wire       [31:0]   _zz_3573;
  wire       [31:0]   _zz_3574;
  wire       [31:0]   _zz_3575;
  wire       [31:0]   _zz_3576;
  wire       [31:0]   _zz_3577;
  wire       [31:0]   _zz_3578;
  wire       [31:0]   _zz_3579;
  wire       [31:0]   _zz_3580;
  wire       [31:0]   _zz_3581;
  wire       [31:0]   _zz_3582;
  wire       [31:0]   _zz_3583;
  wire       [31:0]   _zz_3584;
  wire       [31:0]   _zz_3585;
  wire       [31:0]   _zz_3586;
  wire       [31:0]   _zz_3587;
  wire       [31:0]   _zz_3588;
  wire       [31:0]   _zz_3589;
  wire       [31:0]   _zz_3590;
  wire       [31:0]   _zz_3591;
  wire       [31:0]   _zz_3592;
  wire       [31:0]   _zz_3593;
  wire       [31:0]   _zz_3594;
  wire       [31:0]   _zz_3595;
  wire       [31:0]   _zz_3596;
  wire       [31:0]   _zz_3597;
  wire       [31:0]   _zz_3598;
  wire       [31:0]   _zz_3599;
  wire       [31:0]   _zz_3600;
  wire       [31:0]   _zz_3601;
  wire       [31:0]   _zz_3602;
  wire       [31:0]   _zz_3603;
  wire       [31:0]   _zz_3604;
  wire       [31:0]   _zz_3605;
  wire       [31:0]   _zz_3606;
  wire       [31:0]   _zz_3607;
  wire       [31:0]   _zz_3608;
  wire       [31:0]   _zz_3609;
  wire       [31:0]   _zz_3610;
  wire       [31:0]   _zz_3611;
  wire       [31:0]   _zz_3612;
  wire       [31:0]   _zz_3613;
  wire       [31:0]   _zz_3614;
  wire       [31:0]   _zz_3615;
  wire       [31:0]   _zz_3616;
  wire       [31:0]   _zz_3617;
  wire       [31:0]   _zz_3618;
  wire       [31:0]   _zz_3619;
  wire       [31:0]   _zz_3620;
  wire       [31:0]   _zz_3621;
  wire       [31:0]   _zz_3622;
  wire       [31:0]   _zz_3623;
  wire       [31:0]   _zz_3624;
  wire       [31:0]   _zz_3625;
  wire       [31:0]   _zz_3626;
  wire       [31:0]   _zz_3627;
  wire       [31:0]   _zz_3628;
  wire       [31:0]   _zz_3629;
  wire       [31:0]   _zz_3630;
  wire       [31:0]   _zz_3631;
  wire       [31:0]   _zz_3632;
  wire       [31:0]   _zz_3633;
  wire       [31:0]   _zz_3634;
  wire       [31:0]   _zz_3635;
  wire       [31:0]   _zz_3636;
  wire       [31:0]   _zz_3637;
  wire       [31:0]   _zz_3638;
  wire       [31:0]   _zz_3639;
  wire       [31:0]   _zz_3640;
  wire       [31:0]   _zz_3641;
  wire       [31:0]   _zz_3642;
  wire       [31:0]   _zz_3643;
  wire       [31:0]   _zz_3644;
  wire       [31:0]   _zz_3645;
  wire       [31:0]   _zz_3646;
  wire       [31:0]   _zz_3647;
  wire       [31:0]   _zz_3648;
  wire       [31:0]   _zz_3649;
  wire       [31:0]   _zz_3650;
  wire       [31:0]   _zz_3651;
  wire       [31:0]   _zz_3652;
  wire       [31:0]   _zz_3653;
  wire       [31:0]   _zz_3654;
  wire       [31:0]   _zz_3655;
  wire       [31:0]   _zz_3656;
  wire       [31:0]   _zz_3657;
  wire       [31:0]   _zz_3658;
  wire       [31:0]   _zz_3659;
  wire       [31:0]   _zz_3660;
  wire       [31:0]   _zz_3661;
  wire       [31:0]   _zz_3662;
  wire       [31:0]   _zz_3663;
  wire       [31:0]   _zz_3664;
  wire       [31:0]   _zz_3665;
  wire       [31:0]   _zz_3666;
  wire       [31:0]   _zz_3667;
  wire       [31:0]   _zz_3668;
  wire       [31:0]   _zz_3669;
  wire       [31:0]   _zz_3670;
  wire       [31:0]   _zz_3671;
  wire       [31:0]   _zz_3672;
  wire       [31:0]   _zz_3673;
  wire       [31:0]   _zz_3674;
  wire       [31:0]   _zz_3675;
  wire       [31:0]   _zz_3676;
  wire       [31:0]   _zz_3677;
  wire       [31:0]   _zz_3678;
  wire       [31:0]   _zz_3679;
  wire       [31:0]   _zz_3680;
  wire       [31:0]   _zz_3681;
  wire       [31:0]   _zz_3682;
  wire       [31:0]   _zz_3683;
  wire       [31:0]   _zz_3684;
  wire       [31:0]   _zz_3685;
  wire       [31:0]   _zz_3686;
  wire       [31:0]   _zz_3687;
  wire       [31:0]   _zz_3688;
  wire       [31:0]   _zz_3689;
  wire       [31:0]   _zz_3690;
  wire       [31:0]   _zz_3691;
  wire       [31:0]   _zz_3692;
  wire       [31:0]   _zz_3693;
  wire       [31:0]   _zz_3694;
  wire       [31:0]   _zz_3695;
  wire       [31:0]   _zz_3696;
  wire       [31:0]   _zz_3697;
  wire       [31:0]   _zz_3698;
  wire       [31:0]   _zz_3699;
  wire       [31:0]   _zz_3700;
  wire       [31:0]   _zz_3701;
  wire       [31:0]   _zz_3702;
  wire       [31:0]   _zz_3703;
  wire       [31:0]   _zz_3704;
  wire       [31:0]   _zz_3705;
  wire       [31:0]   _zz_3706;
  wire       [31:0]   _zz_3707;
  wire       [31:0]   _zz_3708;
  wire       [31:0]   _zz_3709;
  wire       [31:0]   _zz_3710;
  wire       [31:0]   _zz_3711;
  wire       [31:0]   _zz_3712;
  wire       [31:0]   _zz_3713;
  wire       [31:0]   _zz_3714;
  wire       [31:0]   _zz_3715;
  wire       [31:0]   _zz_3716;
  wire       [31:0]   _zz_3717;
  wire       [31:0]   _zz_3718;
  wire       [31:0]   _zz_3719;
  wire       [31:0]   _zz_3720;
  wire       [31:0]   _zz_3721;
  wire       [31:0]   _zz_3722;
  wire       [31:0]   _zz_3723;
  wire       [31:0]   _zz_3724;
  wire       [31:0]   _zz_3725;
  wire       [31:0]   _zz_3726;
  wire       [31:0]   _zz_3727;
  wire       [31:0]   _zz_3728;
  wire       [31:0]   _zz_3729;
  wire       [31:0]   _zz_3730;
  wire       [31:0]   _zz_3731;
  wire       [31:0]   _zz_3732;
  wire       [31:0]   _zz_3733;
  wire       [31:0]   _zz_3734;
  wire       [31:0]   _zz_3735;
  wire       [31:0]   _zz_3736;
  wire       [31:0]   _zz_3737;
  wire       [31:0]   _zz_3738;
  wire       [31:0]   _zz_3739;
  wire       [31:0]   _zz_3740;
  wire       [31:0]   _zz_3741;
  wire       [31:0]   _zz_3742;
  wire       [31:0]   _zz_3743;
  wire       [31:0]   _zz_3744;
  wire       [31:0]   _zz_3745;
  wire       [31:0]   _zz_3746;
  wire       [31:0]   _zz_3747;
  wire       [31:0]   _zz_3748;
  wire       [31:0]   _zz_3749;
  wire       [31:0]   _zz_3750;
  wire       [31:0]   _zz_3751;
  wire       [31:0]   _zz_3752;
  wire       [31:0]   _zz_3753;
  wire       [31:0]   _zz_3754;
  wire       [31:0]   _zz_3755;
  wire       [31:0]   _zz_3756;
  wire       [31:0]   _zz_3757;
  wire       [31:0]   _zz_3758;
  wire       [31:0]   _zz_3759;
  wire       [31:0]   _zz_3760;
  wire       [31:0]   _zz_3761;
  wire       [31:0]   _zz_3762;
  wire       [31:0]   _zz_3763;
  wire       [31:0]   _zz_3764;
  wire       [31:0]   _zz_3765;
  wire       [31:0]   _zz_3766;
  wire       [31:0]   _zz_3767;
  wire       [31:0]   _zz_3768;
  wire       [31:0]   _zz_3769;
  wire       [31:0]   _zz_3770;
  wire       [31:0]   _zz_3771;
  wire       [31:0]   _zz_3772;
  wire       [31:0]   _zz_3773;
  wire       [31:0]   _zz_3774;
  wire       [31:0]   _zz_3775;
  wire       [31:0]   _zz_3776;
  wire       [31:0]   _zz_3777;
  wire       [31:0]   _zz_3778;
  wire       [31:0]   _zz_3779;
  wire       [31:0]   _zz_3780;
  wire       [31:0]   _zz_3781;
  wire       [31:0]   _zz_3782;
  wire       [31:0]   _zz_3783;
  wire       [31:0]   _zz_3784;
  wire       [31:0]   _zz_3785;
  wire       [31:0]   _zz_3786;
  wire       [31:0]   _zz_3787;
  wire       [31:0]   _zz_3788;
  wire       [31:0]   _zz_3789;
  wire       [31:0]   _zz_3790;
  wire       [31:0]   _zz_3791;
  wire       [31:0]   _zz_3792;
  wire       [31:0]   _zz_3793;
  wire       [31:0]   _zz_3794;
  wire       [31:0]   _zz_3795;
  wire       [31:0]   _zz_3796;
  wire       [31:0]   _zz_3797;
  wire       [31:0]   _zz_3798;
  wire       [31:0]   _zz_3799;
  wire       [31:0]   _zz_3800;
  wire       [31:0]   _zz_3801;
  wire       [31:0]   _zz_3802;
  wire       [31:0]   _zz_3803;
  wire       [31:0]   _zz_3804;
  wire       [31:0]   _zz_3805;
  wire       [31:0]   _zz_3806;
  wire       [31:0]   _zz_3807;
  wire       [31:0]   _zz_3808;
  wire       [31:0]   _zz_3809;
  wire       [31:0]   _zz_3810;
  wire       [31:0]   _zz_3811;
  wire       [31:0]   _zz_3812;
  wire       [31:0]   _zz_3813;
  wire       [31:0]   _zz_3814;
  wire       [31:0]   _zz_3815;
  wire       [31:0]   _zz_3816;
  wire       [31:0]   _zz_3817;
  wire       [31:0]   _zz_3818;
  wire       [31:0]   _zz_3819;
  wire       [31:0]   _zz_3820;
  wire       [31:0]   _zz_3821;
  wire       [31:0]   _zz_3822;
  wire       [31:0]   _zz_3823;
  wire       [31:0]   _zz_3824;
  wire       [31:0]   _zz_3825;
  wire       [31:0]   _zz_3826;
  wire       [31:0]   _zz_3827;
  wire       [31:0]   _zz_3828;
  wire       [31:0]   _zz_3829;
  wire       [31:0]   _zz_3830;
  wire       [31:0]   _zz_3831;
  wire       [31:0]   _zz_3832;
  wire       [31:0]   _zz_3833;
  wire       [31:0]   _zz_3834;
  wire       [31:0]   _zz_3835;
  wire       [31:0]   _zz_3836;
  wire       [31:0]   _zz_3837;
  wire       [31:0]   _zz_3838;
  wire       [31:0]   _zz_3839;
  wire       [31:0]   _zz_3840;
  wire       [31:0]   _zz_3841;
  wire       [31:0]   _zz_3842;
  wire       [31:0]   _zz_3843;
  wire       [31:0]   _zz_3844;
  wire       [31:0]   _zz_3845;
  wire       [31:0]   _zz_3846;
  wire       [31:0]   _zz_3847;
  wire       [31:0]   _zz_3848;
  wire       [31:0]   _zz_3849;
  wire       [31:0]   _zz_3850;
  wire       [31:0]   _zz_3851;
  wire       [31:0]   _zz_3852;
  wire       [31:0]   _zz_3853;
  wire       [31:0]   _zz_3854;
  wire       [31:0]   _zz_3855;
  wire       [31:0]   _zz_3856;
  wire       [31:0]   _zz_3857;
  wire       [31:0]   _zz_3858;
  wire       [31:0]   _zz_3859;
  wire       [31:0]   _zz_3860;
  wire       [31:0]   _zz_3861;
  wire       [31:0]   _zz_3862;
  wire       [31:0]   _zz_3863;
  wire       [31:0]   _zz_3864;
  wire       [31:0]   _zz_3865;
  wire       [31:0]   _zz_3866;
  wire       [31:0]   _zz_3867;
  wire       [31:0]   _zz_3868;
  wire       [31:0]   _zz_3869;
  wire       [31:0]   _zz_3870;
  wire       [31:0]   _zz_3871;
  wire       [31:0]   _zz_3872;
  wire       [31:0]   _zz_3873;
  wire       [31:0]   _zz_3874;
  wire       [31:0]   _zz_3875;
  wire       [31:0]   _zz_3876;
  wire       [31:0]   _zz_3877;
  wire       [31:0]   _zz_3878;
  wire       [31:0]   _zz_3879;
  wire       [31:0]   _zz_3880;
  wire       [31:0]   _zz_3881;
  wire       [31:0]   _zz_3882;
  wire       [31:0]   _zz_3883;
  wire       [31:0]   _zz_3884;
  wire       [31:0]   _zz_3885;
  wire       [31:0]   _zz_3886;
  wire       [31:0]   _zz_3887;
  wire       [31:0]   _zz_3888;
  wire       [31:0]   _zz_3889;
  wire       [31:0]   _zz_3890;
  wire       [31:0]   _zz_3891;
  wire       [31:0]   _zz_3892;
  wire       [31:0]   _zz_3893;
  wire       [31:0]   _zz_3894;
  wire       [31:0]   _zz_3895;
  wire       [31:0]   _zz_3896;
  wire       [31:0]   _zz_3897;
  wire       [31:0]   _zz_3898;
  wire       [31:0]   _zz_3899;
  wire       [31:0]   _zz_3900;
  wire       [31:0]   _zz_3901;
  wire       [31:0]   _zz_3902;
  wire       [31:0]   _zz_3903;
  wire       [31:0]   _zz_3904;
  wire       [31:0]   _zz_3905;
  wire       [31:0]   _zz_3906;
  wire       [31:0]   _zz_3907;
  wire       [31:0]   _zz_3908;
  wire       [31:0]   _zz_3909;
  wire       [31:0]   _zz_3910;
  wire       [31:0]   _zz_3911;
  wire       [31:0]   _zz_3912;
  wire       [31:0]   _zz_3913;
  wire       [31:0]   _zz_3914;
  wire       [31:0]   _zz_3915;
  wire       [31:0]   _zz_3916;
  wire       [31:0]   _zz_3917;
  wire       [31:0]   _zz_3918;
  wire       [31:0]   _zz_3919;
  wire       [31:0]   _zz_3920;
  wire       [31:0]   _zz_3921;
  wire       [31:0]   _zz_3922;
  wire       [31:0]   _zz_3923;
  wire       [31:0]   _zz_3924;
  wire       [31:0]   _zz_3925;
  wire       [31:0]   _zz_3926;
  wire       [31:0]   _zz_3927;
  wire       [31:0]   _zz_3928;
  wire       [31:0]   _zz_3929;
  wire       [31:0]   _zz_3930;
  wire       [31:0]   _zz_3931;
  wire       [31:0]   _zz_3932;
  wire       [31:0]   _zz_3933;
  wire       [31:0]   _zz_3934;
  wire       [31:0]   _zz_3935;
  wire       [31:0]   _zz_3936;
  wire       [31:0]   _zz_3937;
  wire       [31:0]   _zz_3938;
  wire       [31:0]   _zz_3939;
  wire       [31:0]   _zz_3940;
  wire       [31:0]   _zz_3941;
  wire       [31:0]   _zz_3942;
  wire       [31:0]   _zz_3943;
  wire       [31:0]   _zz_3944;
  wire       [31:0]   _zz_3945;
  wire       [31:0]   _zz_3946;
  wire       [31:0]   _zz_3947;
  wire       [31:0]   _zz_3948;
  wire       [31:0]   _zz_3949;
  wire       [31:0]   _zz_3950;
  wire       [31:0]   _zz_3951;
  wire       [31:0]   _zz_3952;
  wire       [31:0]   _zz_3953;
  wire       [31:0]   _zz_3954;
  wire       [31:0]   _zz_3955;
  wire       [31:0]   _zz_3956;
  wire       [31:0]   _zz_3957;
  wire       [31:0]   _zz_3958;
  wire       [31:0]   _zz_3959;
  wire       [31:0]   _zz_3960;
  wire       [31:0]   _zz_3961;
  wire       [31:0]   _zz_3962;
  wire       [31:0]   _zz_3963;
  wire       [31:0]   _zz_3964;
  wire       [31:0]   _zz_3965;
  wire       [31:0]   _zz_3966;
  wire       [31:0]   _zz_3967;
  wire       [31:0]   _zz_3968;
  wire       [31:0]   _zz_3969;
  wire       [31:0]   _zz_3970;
  wire       [31:0]   _zz_3971;
  wire       [31:0]   _zz_3972;
  wire       [31:0]   _zz_3973;
  wire       [31:0]   _zz_3974;
  wire       [31:0]   _zz_3975;
  wire       [31:0]   _zz_3976;
  wire       [31:0]   _zz_3977;
  wire       [31:0]   _zz_3978;
  wire       [31:0]   _zz_3979;
  wire       [31:0]   _zz_3980;
  wire       [31:0]   _zz_3981;
  wire       [31:0]   _zz_3982;
  wire       [31:0]   _zz_3983;
  wire       [31:0]   _zz_3984;
  wire       [31:0]   _zz_3985;
  wire       [31:0]   _zz_3986;
  wire       [31:0]   _zz_3987;
  wire       [31:0]   _zz_3988;
  wire       [31:0]   _zz_3989;
  wire       [31:0]   _zz_3990;
  wire       [31:0]   _zz_3991;
  wire       [31:0]   _zz_3992;
  wire       [31:0]   _zz_3993;
  wire       [31:0]   _zz_3994;
  wire       [31:0]   _zz_3995;
  wire       [31:0]   _zz_3996;
  wire       [31:0]   _zz_3997;
  wire       [31:0]   _zz_3998;
  wire       [31:0]   _zz_3999;
  wire       [31:0]   _zz_4000;
  wire       [31:0]   _zz_4001;
  wire       [31:0]   _zz_4002;
  wire       [31:0]   _zz_4003;
  wire       [31:0]   _zz_4004;
  wire       [31:0]   _zz_4005;
  wire       [31:0]   _zz_4006;
  wire       [31:0]   _zz_4007;
  wire       [31:0]   _zz_4008;
  wire       [31:0]   _zz_4009;
  wire       [31:0]   _zz_4010;
  wire       [31:0]   _zz_4011;
  wire       [31:0]   _zz_4012;
  wire       [31:0]   _zz_4013;
  wire       [31:0]   _zz_4014;
  wire       [31:0]   _zz_4015;
  wire       [31:0]   _zz_4016;
  wire       [31:0]   _zz_4017;
  wire       [31:0]   _zz_4018;
  wire       [31:0]   _zz_4019;
  wire       [31:0]   _zz_4020;
  wire       [31:0]   _zz_4021;
  wire       [31:0]   _zz_4022;
  wire       [31:0]   _zz_4023;
  wire       [31:0]   _zz_4024;
  wire       [31:0]   _zz_4025;
  wire       [31:0]   _zz_4026;
  wire       [31:0]   _zz_4027;
  wire       [31:0]   _zz_4028;
  wire       [31:0]   _zz_4029;
  wire       [31:0]   _zz_4030;
  wire       [31:0]   _zz_4031;
  wire       [31:0]   _zz_4032;
  wire       [31:0]   _zz_4033;
  wire       [31:0]   _zz_4034;
  wire       [31:0]   _zz_4035;
  wire       [31:0]   _zz_4036;
  wire       [31:0]   _zz_4037;
  wire       [31:0]   _zz_4038;
  wire       [31:0]   _zz_4039;
  wire       [31:0]   _zz_4040;
  wire       [31:0]   _zz_4041;
  wire       [31:0]   _zz_4042;
  wire       [31:0]   _zz_4043;
  wire       [31:0]   _zz_4044;
  wire       [31:0]   _zz_4045;
  wire       [31:0]   _zz_4046;
  wire       [31:0]   _zz_4047;
  wire       [31:0]   _zz_4048;
  wire       [31:0]   _zz_4049;
  wire       [31:0]   _zz_4050;
  wire       [31:0]   _zz_4051;
  wire       [31:0]   _zz_4052;
  wire       [31:0]   _zz_4053;
  wire       [31:0]   _zz_4054;
  wire       [31:0]   _zz_4055;
  wire       [31:0]   _zz_4056;
  wire       [31:0]   _zz_4057;
  wire       [31:0]   _zz_4058;
  wire       [31:0]   _zz_4059;
  wire       [31:0]   _zz_4060;
  wire       [31:0]   _zz_4061;
  wire       [31:0]   _zz_4062;
  wire       [31:0]   _zz_4063;
  wire       [31:0]   _zz_4064;
  wire       [31:0]   _zz_4065;
  wire       [31:0]   _zz_4066;
  wire       [31:0]   _zz_4067;
  wire       [31:0]   _zz_4068;
  wire       [31:0]   _zz_4069;
  wire       [31:0]   _zz_4070;
  wire       [31:0]   _zz_4071;
  wire       [31:0]   _zz_4072;
  wire       [31:0]   _zz_4073;
  wire       [31:0]   _zz_4074;
  wire       [31:0]   _zz_4075;
  wire       [31:0]   _zz_4076;
  wire       [31:0]   _zz_4077;
  wire       [31:0]   _zz_4078;
  wire       [31:0]   _zz_4079;
  wire       [31:0]   _zz_4080;
  wire       [31:0]   _zz_4081;
  wire       [31:0]   _zz_4082;
  wire       [31:0]   _zz_4083;
  wire       [31:0]   _zz_4084;
  wire       [31:0]   _zz_4085;
  wire       [31:0]   _zz_4086;
  wire       [31:0]   _zz_4087;
  wire       [31:0]   _zz_4088;
  wire       [31:0]   _zz_4089;
  wire       [31:0]   _zz_4090;
  wire       [31:0]   _zz_4091;
  wire       [31:0]   _zz_4092;
  wire       [31:0]   _zz_4093;
  wire       [31:0]   _zz_4094;
  wire       [31:0]   _zz_4095;
  wire       [31:0]   _zz_4096;
  wire       [31:0]   _zz_4097;
  wire       [31:0]   _zz_4098;
  wire       [31:0]   _zz_4099;
  wire       [31:0]   _zz_4100;
  wire       [31:0]   _zz_4101;
  wire       [31:0]   _zz_4102;
  wire       [31:0]   _zz_4103;
  wire       [31:0]   _zz_4104;
  wire       [31:0]   _zz_4105;
  wire       [31:0]   _zz_4106;
  wire       [31:0]   _zz_4107;
  wire       [31:0]   _zz_4108;
  wire       [31:0]   _zz_4109;
  wire       [31:0]   _zz_4110;
  wire       [31:0]   _zz_4111;
  wire       [31:0]   _zz_4112;
  wire       [31:0]   _zz_4113;
  wire       [31:0]   _zz_4114;
  wire       [31:0]   _zz_4115;
  wire       [31:0]   _zz_4116;
  wire       [31:0]   _zz_4117;
  wire       [31:0]   _zz_4118;
  wire       [31:0]   _zz_4119;
  wire       [31:0]   _zz_4120;
  wire       [31:0]   _zz_4121;
  wire       [31:0]   _zz_4122;
  wire       [31:0]   _zz_4123;
  wire       [31:0]   _zz_4124;
  wire       [31:0]   _zz_4125;
  wire       [31:0]   _zz_4126;
  wire       [31:0]   _zz_4127;
  wire       [31:0]   _zz_4128;
  wire       [31:0]   _zz_4129;
  wire       [31:0]   _zz_4130;
  wire       [31:0]   _zz_4131;
  wire       [31:0]   _zz_4132;
  wire       [31:0]   _zz_4133;
  wire       [31:0]   _zz_4134;
  wire       [31:0]   _zz_4135;
  wire       [31:0]   _zz_4136;
  wire       [31:0]   _zz_4137;
  wire       [31:0]   _zz_4138;
  wire       [31:0]   _zz_4139;
  wire       [31:0]   _zz_4140;
  wire       [31:0]   _zz_4141;
  wire       [31:0]   _zz_4142;
  wire       [31:0]   _zz_4143;
  wire       [31:0]   _zz_4144;
  wire       [31:0]   _zz_4145;
  wire       [31:0]   _zz_4146;
  wire       [31:0]   _zz_4147;
  wire       [31:0]   _zz_4148;
  wire       [31:0]   _zz_4149;
  wire       [31:0]   _zz_4150;
  wire       [31:0]   _zz_4151;
  wire       [31:0]   _zz_4152;
  wire       [31:0]   _zz_4153;
  wire       [31:0]   _zz_4154;
  wire       [31:0]   _zz_4155;
  wire       [31:0]   _zz_4156;
  wire       [31:0]   _zz_4157;
  wire       [31:0]   _zz_4158;
  wire       [31:0]   _zz_4159;
  wire       [31:0]   _zz_4160;
  wire       [31:0]   _zz_4161;
  wire       [31:0]   _zz_4162;
  wire       [31:0]   _zz_4163;
  wire       [31:0]   _zz_4164;
  wire       [31:0]   _zz_4165;
  wire       [31:0]   _zz_4166;
  wire       [31:0]   _zz_4167;
  wire       [31:0]   _zz_4168;
  wire       [31:0]   _zz_4169;
  wire       [31:0]   _zz_4170;
  wire       [31:0]   _zz_4171;
  wire       [31:0]   _zz_4172;
  wire       [31:0]   _zz_4173;
  wire       [31:0]   _zz_4174;
  wire       [31:0]   _zz_4175;
  wire       [31:0]   _zz_4176;
  wire       [31:0]   _zz_4177;
  wire       [31:0]   _zz_4178;
  wire       [31:0]   _zz_4179;
  wire       [31:0]   _zz_4180;
  wire       [31:0]   _zz_4181;
  wire       [31:0]   _zz_4182;
  wire       [31:0]   _zz_4183;
  wire       [31:0]   _zz_4184;
  wire       [31:0]   _zz_4185;
  wire       [31:0]   _zz_4186;
  wire       [31:0]   _zz_4187;
  wire       [31:0]   _zz_4188;
  wire       [31:0]   _zz_4189;
  wire       [31:0]   _zz_4190;
  wire       [31:0]   _zz_4191;
  wire       [31:0]   _zz_4192;
  wire       [31:0]   _zz_4193;
  wire       [31:0]   _zz_4194;
  wire       [31:0]   _zz_4195;
  wire       [31:0]   _zz_4196;
  wire       [31:0]   _zz_4197;
  wire       [31:0]   _zz_4198;
  wire       [31:0]   _zz_4199;
  wire       [31:0]   _zz_4200;
  wire       [31:0]   _zz_4201;
  wire       [31:0]   _zz_4202;
  wire       [31:0]   _zz_4203;
  wire       [31:0]   _zz_4204;
  wire       [31:0]   _zz_4205;
  wire       [31:0]   _zz_4206;
  wire       [31:0]   _zz_4207;
  wire       [31:0]   _zz_4208;
  wire       [31:0]   _zz_4209;
  wire       [31:0]   _zz_4210;
  wire       [31:0]   _zz_4211;
  wire       [31:0]   _zz_4212;
  wire       [31:0]   _zz_4213;
  wire       [31:0]   _zz_4214;
  wire       [31:0]   _zz_4215;
  wire       [31:0]   _zz_4216;
  wire       [31:0]   _zz_4217;
  wire       [31:0]   _zz_4218;
  wire       [31:0]   _zz_4219;
  wire       [31:0]   _zz_4220;
  wire       [31:0]   _zz_4221;
  wire       [31:0]   _zz_4222;
  wire       [31:0]   _zz_4223;
  wire       [31:0]   _zz_4224;
  wire       [31:0]   _zz_4225;
  wire       [31:0]   _zz_4226;
  wire       [31:0]   _zz_4227;
  wire       [31:0]   _zz_4228;
  wire       [31:0]   _zz_4229;
  wire       [31:0]   _zz_4230;
  wire       [31:0]   _zz_4231;
  wire       [31:0]   _zz_4232;
  wire       [31:0]   _zz_4233;
  wire       [31:0]   _zz_4234;
  wire       [31:0]   _zz_4235;
  wire       [31:0]   _zz_4236;
  wire       [31:0]   _zz_4237;
  wire       [31:0]   _zz_4238;
  wire       [31:0]   _zz_4239;
  wire       [31:0]   _zz_4240;
  wire       [31:0]   _zz_4241;
  wire       [31:0]   _zz_4242;
  wire       [31:0]   _zz_4243;
  wire       [31:0]   _zz_4244;
  wire       [31:0]   _zz_4245;
  wire       [31:0]   _zz_4246;
  wire       [31:0]   _zz_4247;
  wire       [31:0]   _zz_4248;
  wire       [31:0]   _zz_4249;
  wire       [31:0]   _zz_4250;
  wire       [31:0]   _zz_4251;
  wire       [31:0]   _zz_4252;
  wire       [31:0]   _zz_4253;
  wire       [31:0]   _zz_4254;
  wire       [31:0]   _zz_4255;
  wire       [31:0]   _zz_4256;
  wire       [31:0]   _zz_4257;
  wire       [31:0]   _zz_4258;
  wire       [31:0]   _zz_4259;
  wire       [31:0]   _zz_4260;
  wire       [31:0]   _zz_4261;
  wire       [31:0]   _zz_4262;
  wire       [31:0]   _zz_4263;
  wire       [31:0]   _zz_4264;
  wire       [31:0]   _zz_4265;
  wire       [31:0]   _zz_4266;
  wire       [31:0]   _zz_4267;
  wire       [31:0]   _zz_4268;
  wire       [31:0]   _zz_4269;
  wire       [31:0]   _zz_4270;
  wire       [31:0]   _zz_4271;
  wire       [31:0]   _zz_4272;
  wire       [31:0]   _zz_4273;
  wire       [31:0]   _zz_4274;
  wire       [31:0]   _zz_4275;
  wire       [31:0]   _zz_4276;
  wire       [31:0]   _zz_4277;
  wire       [31:0]   _zz_4278;
  wire       [31:0]   _zz_4279;
  wire       [31:0]   _zz_4280;
  wire       [31:0]   _zz_4281;
  wire       [31:0]   _zz_4282;
  wire       [31:0]   _zz_4283;
  wire       [31:0]   _zz_4284;
  wire       [31:0]   _zz_4285;
  wire       [31:0]   _zz_4286;
  wire       [31:0]   _zz_4287;
  wire       [31:0]   _zz_4288;
  wire       [31:0]   _zz_4289;
  wire       [31:0]   _zz_4290;
  wire       [31:0]   _zz_4291;
  wire       [31:0]   _zz_4292;
  wire       [31:0]   _zz_4293;
  wire       [31:0]   _zz_4294;
  wire       [31:0]   _zz_4295;
  wire       [31:0]   _zz_4296;
  wire       [31:0]   _zz_4297;
  wire       [31:0]   _zz_4298;
  wire       [31:0]   _zz_4299;
  wire       [31:0]   _zz_4300;
  wire       [31:0]   _zz_4301;
  wire       [31:0]   _zz_4302;
  wire       [31:0]   _zz_4303;
  wire       [31:0]   _zz_4304;
  wire       [31:0]   _zz_4305;
  wire       [31:0]   _zz_4306;
  wire       [31:0]   _zz_4307;
  wire       [31:0]   _zz_4308;
  wire       [31:0]   _zz_4309;
  wire       [31:0]   _zz_4310;
  wire       [31:0]   _zz_4311;
  wire       [31:0]   _zz_4312;
  wire       [31:0]   _zz_4313;
  wire       [31:0]   _zz_4314;
  wire       [31:0]   _zz_4315;
  wire       [31:0]   _zz_4316;
  wire       [31:0]   _zz_4317;
  wire       [31:0]   _zz_4318;
  wire       [31:0]   _zz_4319;
  wire       [31:0]   _zz_4320;
  wire       [31:0]   _zz_4321;
  wire       [31:0]   _zz_4322;
  wire       [31:0]   _zz_4323;
  wire       [31:0]   _zz_4324;
  wire       [31:0]   _zz_4325;
  wire       [31:0]   _zz_4326;
  wire       [31:0]   _zz_4327;
  wire       [31:0]   _zz_4328;
  wire       [31:0]   _zz_4329;
  wire       [31:0]   _zz_4330;
  wire       [31:0]   _zz_4331;
  wire       [31:0]   _zz_4332;
  wire       [31:0]   _zz_4333;
  wire       [31:0]   _zz_4334;
  wire       [31:0]   _zz_4335;
  wire       [31:0]   _zz_4336;
  wire       [31:0]   _zz_4337;
  wire       [31:0]   _zz_4338;
  wire       [31:0]   _zz_4339;
  wire       [31:0]   _zz_4340;
  wire       [31:0]   _zz_4341;
  wire       [31:0]   _zz_4342;
  wire       [31:0]   _zz_4343;
  wire       [31:0]   _zz_4344;
  wire       [31:0]   _zz_4345;
  wire       [31:0]   _zz_4346;
  wire       [31:0]   _zz_4347;
  wire       [31:0]   _zz_4348;
  wire       [31:0]   _zz_4349;
  wire       [31:0]   _zz_4350;
  wire       [31:0]   _zz_4351;
  wire       [31:0]   _zz_4352;
  wire       [31:0]   _zz_4353;
  wire       [31:0]   _zz_4354;
  wire       [31:0]   _zz_4355;
  wire       [31:0]   _zz_4356;
  wire       [31:0]   _zz_4357;
  wire       [31:0]   _zz_4358;
  wire       [31:0]   _zz_4359;
  wire       [31:0]   _zz_4360;
  wire       [31:0]   _zz_4361;
  wire       [31:0]   _zz_4362;
  wire       [31:0]   _zz_4363;
  wire       [31:0]   _zz_4364;
  wire       [31:0]   _zz_4365;
  wire       [31:0]   _zz_4366;
  wire       [31:0]   _zz_4367;
  wire       [31:0]   _zz_4368;
  wire       [31:0]   _zz_4369;
  wire       [31:0]   _zz_4370;
  wire       [31:0]   _zz_4371;
  wire       [31:0]   _zz_4372;
  wire       [31:0]   _zz_4373;
  wire       [31:0]   _zz_4374;
  wire       [31:0]   _zz_4375;
  wire       [31:0]   _zz_4376;
  wire       [31:0]   _zz_4377;
  wire       [31:0]   _zz_4378;
  wire       [31:0]   _zz_4379;
  wire       [31:0]   _zz_4380;
  wire       [31:0]   _zz_4381;
  wire       [31:0]   _zz_4382;
  wire       [31:0]   _zz_4383;
  wire       [31:0]   _zz_4384;
  wire       [31:0]   _zz_4385;
  wire       [31:0]   _zz_4386;
  wire       [31:0]   _zz_4387;
  wire       [31:0]   _zz_4388;
  wire       [31:0]   _zz_4389;
  wire       [31:0]   _zz_4390;
  wire       [31:0]   _zz_4391;
  wire       [31:0]   _zz_4392;
  wire       [31:0]   _zz_4393;
  wire       [31:0]   _zz_4394;
  wire       [31:0]   _zz_4395;
  wire       [31:0]   _zz_4396;
  wire       [31:0]   _zz_4397;
  wire       [31:0]   _zz_4398;
  wire       [31:0]   _zz_4399;
  wire       [31:0]   _zz_4400;
  wire       [31:0]   _zz_4401;
  wire       [31:0]   _zz_4402;
  wire       [31:0]   _zz_4403;
  wire       [31:0]   _zz_4404;
  wire       [31:0]   _zz_4405;
  wire       [31:0]   _zz_4406;
  wire       [31:0]   _zz_4407;
  wire       [31:0]   _zz_4408;
  wire       [31:0]   _zz_4409;
  wire       [31:0]   _zz_4410;
  wire       [31:0]   _zz_4411;
  wire       [31:0]   _zz_4412;
  wire       [31:0]   _zz_4413;
  wire       [31:0]   _zz_4414;
  wire       [31:0]   _zz_4415;
  wire       [31:0]   _zz_4416;
  wire       [31:0]   _zz_4417;
  wire       [31:0]   _zz_4418;
  wire       [31:0]   _zz_4419;
  wire       [31:0]   _zz_4420;
  wire       [31:0]   _zz_4421;
  wire       [31:0]   _zz_4422;
  wire       [31:0]   _zz_4423;
  wire       [31:0]   _zz_4424;
  wire       [31:0]   _zz_4425;
  wire       [31:0]   _zz_4426;
  wire       [31:0]   _zz_4427;
  wire       [31:0]   _zz_4428;
  wire       [31:0]   _zz_4429;
  wire       [31:0]   _zz_4430;
  wire       [31:0]   _zz_4431;
  wire       [31:0]   _zz_4432;
  wire       [31:0]   _zz_4433;
  wire       [31:0]   _zz_4434;
  wire       [31:0]   _zz_4435;
  wire       [31:0]   _zz_4436;
  wire       [31:0]   _zz_4437;
  wire       [31:0]   _zz_4438;
  wire       [31:0]   _zz_4439;
  wire       [31:0]   _zz_4440;
  wire       [31:0]   _zz_4441;
  wire       [31:0]   _zz_4442;
  wire       [31:0]   _zz_4443;
  wire       [31:0]   _zz_4444;
  wire       [31:0]   _zz_4445;
  wire       [31:0]   _zz_4446;
  wire       [31:0]   _zz_4447;
  wire       [31:0]   _zz_4448;
  wire       [31:0]   _zz_4449;
  wire       [31:0]   _zz_4450;
  wire       [31:0]   _zz_4451;
  wire       [31:0]   _zz_4452;
  wire       [31:0]   _zz_4453;
  wire       [31:0]   _zz_4454;
  wire       [31:0]   _zz_4455;
  wire       [31:0]   _zz_4456;
  wire       [31:0]   _zz_4457;
  wire       [31:0]   _zz_4458;
  wire       [31:0]   _zz_4459;
  wire       [31:0]   _zz_4460;
  wire       [31:0]   _zz_4461;
  wire       [31:0]   _zz_4462;
  wire       [31:0]   _zz_4463;
  wire       [31:0]   _zz_4464;
  wire       [31:0]   _zz_4465;
  wire       [31:0]   _zz_4466;
  wire       [31:0]   _zz_4467;
  wire       [31:0]   _zz_4468;
  wire       [31:0]   _zz_4469;
  wire       [31:0]   _zz_4470;
  wire       [31:0]   _zz_4471;
  wire       [31:0]   _zz_4472;
  wire       [31:0]   _zz_4473;
  wire       [31:0]   _zz_4474;
  wire       [31:0]   _zz_4475;
  wire       [31:0]   _zz_4476;
  wire       [31:0]   _zz_4477;
  wire       [31:0]   _zz_4478;
  wire       [31:0]   _zz_4479;
  wire       [31:0]   _zz_4480;
  wire       [31:0]   _zz_4481;
  wire       [31:0]   _zz_4482;
  wire       [31:0]   _zz_4483;
  wire       [31:0]   _zz_4484;
  wire       [31:0]   _zz_4485;
  wire       [31:0]   _zz_4486;
  wire       [31:0]   _zz_4487;
  wire       [31:0]   _zz_4488;
  wire       [31:0]   _zz_4489;
  wire       [31:0]   _zz_4490;
  wire       [31:0]   _zz_4491;
  wire       [31:0]   _zz_4492;
  wire       [31:0]   _zz_4493;
  wire       [31:0]   _zz_4494;
  wire       [31:0]   _zz_4495;
  wire       [31:0]   _zz_4496;
  wire       [31:0]   _zz_4497;
  wire       [31:0]   _zz_4498;
  wire       [31:0]   _zz_4499;
  wire       [31:0]   _zz_4500;
  wire       [31:0]   _zz_4501;
  wire       [31:0]   _zz_4502;
  wire       [31:0]   _zz_4503;
  wire       [31:0]   _zz_4504;
  wire       [31:0]   _zz_4505;
  wire       [31:0]   _zz_4506;
  wire       [31:0]   _zz_4507;
  wire       [31:0]   _zz_4508;
  wire       [31:0]   _zz_4509;
  wire       [31:0]   _zz_4510;
  wire       [31:0]   _zz_4511;
  wire       [31:0]   _zz_4512;
  wire       [31:0]   _zz_4513;
  wire       [31:0]   _zz_4514;
  wire       [31:0]   _zz_4515;
  wire       [31:0]   _zz_4516;
  wire       [31:0]   _zz_4517;
  wire       [31:0]   _zz_4518;
  wire       [31:0]   _zz_4519;
  wire       [31:0]   _zz_4520;
  wire       [31:0]   _zz_4521;
  wire       [31:0]   _zz_4522;
  wire       [31:0]   _zz_4523;
  wire       [31:0]   _zz_4524;
  wire       [31:0]   _zz_4525;
  wire       [31:0]   _zz_4526;
  wire       [31:0]   _zz_4527;
  wire       [31:0]   _zz_4528;
  wire       [31:0]   _zz_4529;
  wire       [31:0]   _zz_4530;
  wire       [31:0]   _zz_4531;
  wire       [31:0]   _zz_4532;
  wire       [31:0]   _zz_4533;
  wire       [31:0]   _zz_4534;
  wire       [31:0]   _zz_4535;
  wire       [31:0]   _zz_4536;
  wire       [31:0]   _zz_4537;
  wire       [31:0]   _zz_4538;
  wire       [31:0]   _zz_4539;
  wire       [31:0]   _zz_4540;
  wire       [31:0]   _zz_4541;
  wire       [31:0]   _zz_4542;
  wire       [31:0]   _zz_4543;
  wire       [31:0]   _zz_4544;
  wire       [31:0]   _zz_4545;
  wire       [31:0]   _zz_4546;
  wire       [31:0]   _zz_4547;
  wire       [31:0]   _zz_4548;
  wire       [31:0]   _zz_4549;
  wire       [31:0]   _zz_4550;
  wire       [31:0]   _zz_4551;
  wire       [31:0]   _zz_4552;
  wire       [31:0]   _zz_4553;
  wire       [31:0]   _zz_4554;
  wire       [31:0]   _zz_4555;
  wire       [31:0]   _zz_4556;
  wire       [31:0]   _zz_4557;
  wire       [31:0]   _zz_4558;
  wire       [31:0]   _zz_4559;
  wire       [31:0]   _zz_4560;
  wire       [31:0]   _zz_4561;
  wire       [31:0]   _zz_4562;
  wire       [31:0]   _zz_4563;
  wire       [31:0]   _zz_4564;
  wire       [31:0]   _zz_4565;
  wire       [31:0]   _zz_4566;
  wire       [31:0]   _zz_4567;
  wire       [31:0]   _zz_4568;
  wire       [31:0]   _zz_4569;
  wire       [31:0]   _zz_4570;
  wire       [31:0]   _zz_4571;
  wire       [31:0]   _zz_4572;
  wire       [31:0]   _zz_4573;
  wire       [31:0]   _zz_4574;
  wire       [31:0]   _zz_4575;
  wire       [31:0]   _zz_4576;
  wire       [31:0]   _zz_4577;
  wire       [31:0]   _zz_4578;
  wire       [31:0]   _zz_4579;
  wire       [31:0]   _zz_4580;
  wire       [31:0]   _zz_4581;
  wire       [31:0]   _zz_4582;
  wire       [31:0]   _zz_4583;
  wire       [31:0]   _zz_4584;
  wire       [31:0]   _zz_4585;
  wire       [31:0]   _zz_4586;
  wire       [31:0]   _zz_4587;
  wire       [31:0]   _zz_4588;
  wire       [31:0]   _zz_4589;
  wire       [31:0]   _zz_4590;
  wire       [31:0]   _zz_4591;
  wire       [31:0]   _zz_4592;
  wire       [31:0]   _zz_4593;
  wire       [31:0]   _zz_4594;
  wire       [31:0]   _zz_4595;
  wire       [31:0]   _zz_4596;
  wire       [31:0]   _zz_4597;
  wire       [31:0]   _zz_4598;
  wire       [31:0]   _zz_4599;
  wire       [31:0]   _zz_4600;
  wire       [31:0]   _zz_4601;
  wire       [31:0]   _zz_4602;
  wire       [31:0]   _zz_4603;
  wire       [31:0]   _zz_4604;
  wire       [31:0]   _zz_4605;
  wire       [31:0]   _zz_4606;
  wire       [31:0]   _zz_4607;
  wire       [31:0]   _zz_4608;
  wire       [31:0]   _zz_4609;
  wire       [31:0]   _zz_4610;
  wire       [31:0]   _zz_4611;
  wire       [31:0]   _zz_4612;
  wire       [31:0]   _zz_4613;
  wire       [31:0]   _zz_4614;
  wire       [31:0]   _zz_4615;
  wire       [31:0]   _zz_4616;
  wire       [31:0]   _zz_4617;
  wire       [31:0]   _zz_4618;
  wire       [31:0]   _zz_4619;
  wire       [31:0]   _zz_4620;
  wire       [31:0]   _zz_4621;
  wire       [31:0]   _zz_4622;
  wire       [31:0]   _zz_4623;
  wire       [31:0]   _zz_4624;
  wire       [31:0]   _zz_4625;
  wire       [31:0]   _zz_4626;
  wire       [31:0]   _zz_4627;
  wire       [31:0]   _zz_4628;
  wire       [31:0]   _zz_4629;
  wire       [31:0]   _zz_4630;
  wire       [31:0]   _zz_4631;
  wire       [31:0]   _zz_4632;
  wire       [31:0]   _zz_4633;
  wire       [31:0]   _zz_4634;
  wire       [31:0]   _zz_4635;
  wire       [31:0]   _zz_4636;
  wire       [31:0]   _zz_4637;
  wire       [31:0]   _zz_4638;
  wire       [31:0]   _zz_4639;
  wire       [31:0]   _zz_4640;
  wire       [31:0]   _zz_4641;
  wire       [31:0]   _zz_4642;
  wire       [31:0]   _zz_4643;
  wire       [31:0]   _zz_4644;
  wire       [31:0]   _zz_4645;
  wire       [31:0]   _zz_4646;
  wire       [31:0]   _zz_4647;
  wire       [31:0]   _zz_4648;
  wire       [31:0]   _zz_4649;
  wire       [31:0]   _zz_4650;
  wire       [31:0]   _zz_4651;
  wire       [31:0]   _zz_4652;
  wire       [31:0]   _zz_4653;
  wire       [31:0]   _zz_4654;
  wire       [31:0]   _zz_4655;
  wire       [31:0]   _zz_4656;
  wire       [31:0]   _zz_4657;
  wire       [31:0]   _zz_4658;
  wire       [31:0]   _zz_4659;
  wire       [31:0]   _zz_4660;
  wire       [31:0]   _zz_4661;
  wire       [31:0]   _zz_4662;
  wire       [31:0]   _zz_4663;
  wire       [31:0]   _zz_4664;
  wire       [31:0]   _zz_4665;
  wire       [31:0]   _zz_4666;
  wire       [31:0]   _zz_4667;
  wire       [31:0]   _zz_4668;
  wire       [31:0]   _zz_4669;
  wire       [31:0]   _zz_4670;
  wire       [31:0]   _zz_4671;
  wire       [31:0]   _zz_4672;
  wire       [31:0]   _zz_4673;
  wire       [31:0]   _zz_4674;
  wire       [31:0]   _zz_4675;
  wire       [31:0]   _zz_4676;
  wire       [31:0]   _zz_4677;
  wire       [31:0]   _zz_4678;
  wire       [31:0]   _zz_4679;
  wire       [31:0]   _zz_4680;
  wire       [31:0]   _zz_4681;
  wire       [31:0]   _zz_4682;
  wire       [31:0]   _zz_4683;
  wire       [31:0]   _zz_4684;
  wire       [31:0]   _zz_4685;
  wire       [31:0]   _zz_4686;
  wire       [31:0]   _zz_4687;
  wire       [31:0]   _zz_4688;
  wire       [31:0]   _zz_4689;
  wire       [31:0]   _zz_4690;
  wire       [31:0]   _zz_4691;
  wire       [31:0]   _zz_4692;
  wire       [31:0]   _zz_4693;
  wire       [31:0]   _zz_4694;
  wire       [31:0]   _zz_4695;
  wire       [31:0]   _zz_4696;
  wire       [31:0]   _zz_4697;
  wire       [31:0]   _zz_4698;
  wire       [31:0]   _zz_4699;
  wire       [31:0]   _zz_4700;
  wire       [31:0]   _zz_4701;
  wire       [31:0]   _zz_4702;
  wire       [31:0]   _zz_4703;
  wire       [31:0]   _zz_4704;
  wire       [31:0]   _zz_4705;
  wire       [31:0]   _zz_4706;
  wire       [31:0]   _zz_4707;
  wire       [31:0]   _zz_4708;
  wire       [31:0]   _zz_4709;
  wire       [31:0]   _zz_4710;
  wire       [31:0]   _zz_4711;
  wire       [31:0]   _zz_4712;
  wire       [31:0]   _zz_4713;
  wire       [31:0]   _zz_4714;
  wire       [31:0]   _zz_4715;
  wire       [31:0]   _zz_4716;
  wire       [31:0]   _zz_4717;
  wire       [31:0]   _zz_4718;
  wire       [31:0]   _zz_4719;
  wire       [31:0]   _zz_4720;
  wire       [31:0]   _zz_4721;
  wire       [31:0]   _zz_4722;
  wire       [31:0]   _zz_4723;
  wire       [31:0]   _zz_4724;
  wire       [31:0]   _zz_4725;
  wire       [31:0]   _zz_4726;
  wire       [31:0]   _zz_4727;
  wire       [31:0]   _zz_4728;
  wire       [31:0]   _zz_4729;
  wire       [31:0]   _zz_4730;
  wire       [31:0]   _zz_4731;
  wire       [31:0]   _zz_4732;
  wire       [31:0]   _zz_4733;
  wire       [31:0]   _zz_4734;
  wire       [31:0]   _zz_4735;
  wire       [31:0]   _zz_4736;
  wire       [31:0]   _zz_4737;
  wire       [31:0]   _zz_4738;
  wire       [31:0]   _zz_4739;
  wire       [31:0]   _zz_4740;
  wire       [31:0]   _zz_4741;
  wire       [31:0]   _zz_4742;
  wire       [31:0]   _zz_4743;
  wire       [31:0]   _zz_4744;
  wire       [31:0]   _zz_4745;
  wire       [31:0]   _zz_4746;
  wire       [31:0]   _zz_4747;
  wire       [31:0]   _zz_4748;
  wire       [31:0]   _zz_4749;
  wire       [31:0]   _zz_4750;
  wire       [31:0]   _zz_4751;
  wire       [31:0]   _zz_4752;
  wire       [31:0]   _zz_4753;
  wire       [31:0]   _zz_4754;
  wire       [31:0]   _zz_4755;
  wire       [31:0]   _zz_4756;
  wire       [31:0]   _zz_4757;
  wire       [31:0]   _zz_4758;
  wire       [31:0]   _zz_4759;
  wire       [31:0]   _zz_4760;
  wire       [31:0]   _zz_4761;
  wire       [31:0]   _zz_4762;
  wire       [31:0]   _zz_4763;
  wire       [31:0]   _zz_4764;
  wire       [31:0]   _zz_4765;
  wire       [31:0]   _zz_4766;
  wire       [31:0]   _zz_4767;
  wire       [31:0]   _zz_4768;
  wire       [31:0]   _zz_4769;
  wire       [31:0]   _zz_4770;
  wire       [31:0]   _zz_4771;
  wire       [31:0]   _zz_4772;
  wire       [31:0]   _zz_4773;
  wire       [31:0]   _zz_4774;
  wire       [31:0]   _zz_4775;
  wire       [31:0]   _zz_4776;
  wire       [31:0]   _zz_4777;
  wire       [31:0]   _zz_4778;
  wire       [31:0]   _zz_4779;
  wire       [31:0]   _zz_4780;
  wire       [31:0]   _zz_4781;
  wire       [31:0]   _zz_4782;
  wire       [31:0]   _zz_4783;
  wire       [31:0]   _zz_4784;
  wire       [31:0]   _zz_4785;
  wire       [31:0]   _zz_4786;
  wire       [31:0]   _zz_4787;
  wire       [31:0]   _zz_4788;
  wire       [31:0]   _zz_4789;
  wire       [31:0]   _zz_4790;
  wire       [31:0]   _zz_4791;
  wire       [31:0]   _zz_4792;
  wire       [31:0]   _zz_4793;
  wire       [31:0]   _zz_4794;
  wire       [31:0]   _zz_4795;
  wire       [31:0]   _zz_4796;
  wire       [31:0]   _zz_4797;
  wire       [31:0]   _zz_4798;
  wire       [31:0]   _zz_4799;
  wire       [31:0]   _zz_4800;
  wire       [31:0]   _zz_4801;
  wire       [31:0]   _zz_4802;
  wire       [31:0]   _zz_4803;
  wire       [31:0]   _zz_4804;
  wire       [31:0]   _zz_4805;
  wire       [31:0]   _zz_4806;
  wire       [31:0]   _zz_4807;
  wire       [31:0]   _zz_4808;
  wire       [31:0]   _zz_4809;
  wire       [31:0]   _zz_4810;
  wire       [31:0]   _zz_4811;
  wire       [31:0]   _zz_4812;
  wire       [31:0]   _zz_4813;
  wire       [31:0]   _zz_4814;
  wire       [31:0]   _zz_4815;
  wire       [31:0]   _zz_4816;
  wire       [31:0]   _zz_4817;
  wire       [31:0]   _zz_4818;
  wire       [31:0]   _zz_4819;
  wire       [31:0]   _zz_4820;
  wire       [31:0]   _zz_4821;
  wire       [31:0]   _zz_4822;
  wire       [31:0]   _zz_4823;
  wire       [31:0]   _zz_4824;
  wire       [31:0]   _zz_4825;
  wire       [31:0]   _zz_4826;
  wire       [31:0]   _zz_4827;
  wire       [31:0]   _zz_4828;
  wire       [31:0]   _zz_4829;
  wire       [31:0]   _zz_4830;
  wire       [31:0]   _zz_4831;
  wire       [31:0]   _zz_4832;
  wire       [31:0]   _zz_4833;
  wire       [31:0]   _zz_4834;
  wire       [31:0]   _zz_4835;
  wire       [31:0]   _zz_4836;
  wire       [31:0]   _zz_4837;
  wire       [31:0]   _zz_4838;
  wire       [31:0]   _zz_4839;
  wire       [31:0]   _zz_4840;
  wire       [31:0]   _zz_4841;
  wire       [31:0]   _zz_4842;
  wire       [31:0]   _zz_4843;
  wire       [31:0]   _zz_4844;
  wire       [31:0]   _zz_4845;
  wire       [31:0]   _zz_4846;
  wire       [31:0]   _zz_4847;
  wire       [31:0]   _zz_4848;
  wire       [31:0]   _zz_4849;
  wire       [31:0]   _zz_4850;
  wire       [31:0]   _zz_4851;
  wire       [31:0]   _zz_4852;
  wire       [31:0]   _zz_4853;
  wire       [31:0]   _zz_4854;
  wire       [31:0]   _zz_4855;
  wire       [31:0]   _zz_4856;
  wire       [31:0]   _zz_4857;
  wire       [31:0]   _zz_4858;
  wire       [31:0]   _zz_4859;
  wire       [31:0]   _zz_4860;
  wire       [31:0]   _zz_4861;
  wire       [31:0]   _zz_4862;
  wire       [31:0]   _zz_4863;
  wire       [31:0]   _zz_4864;
  wire       [31:0]   _zz_4865;
  wire       [31:0]   _zz_4866;
  wire       [31:0]   _zz_4867;
  wire       [31:0]   _zz_4868;
  wire       [31:0]   _zz_4869;
  wire       [31:0]   _zz_4870;
  wire       [31:0]   _zz_4871;
  wire       [31:0]   _zz_4872;
  wire       [31:0]   _zz_4873;
  wire       [31:0]   _zz_4874;
  wire       [31:0]   _zz_4875;
  wire       [31:0]   _zz_4876;
  wire       [31:0]   _zz_4877;
  wire       [31:0]   _zz_4878;
  wire       [31:0]   _zz_4879;
  wire       [31:0]   _zz_4880;
  wire       [31:0]   _zz_4881;
  wire       [31:0]   _zz_4882;
  wire       [31:0]   _zz_4883;
  wire       [31:0]   _zz_4884;
  wire       [31:0]   _zz_4885;
  wire       [31:0]   _zz_4886;
  wire       [31:0]   _zz_4887;
  wire       [31:0]   _zz_4888;
  wire       [31:0]   _zz_4889;
  wire       [31:0]   _zz_4890;
  wire       [31:0]   _zz_4891;
  wire       [31:0]   _zz_4892;
  wire       [31:0]   _zz_4893;
  wire       [31:0]   _zz_4894;
  wire       [31:0]   _zz_4895;
  wire       [31:0]   _zz_4896;
  wire       [31:0]   _zz_4897;
  wire       [31:0]   _zz_4898;
  wire       [31:0]   _zz_4899;
  wire       [31:0]   _zz_4900;
  wire       [31:0]   _zz_4901;
  wire       [31:0]   _zz_4902;
  wire       [31:0]   _zz_4903;
  wire       [31:0]   _zz_4904;
  wire       [31:0]   _zz_4905;
  wire       [31:0]   _zz_4906;
  wire       [31:0]   _zz_4907;
  wire       [31:0]   _zz_4908;
  wire       [31:0]   _zz_4909;
  wire       [31:0]   _zz_4910;
  wire       [31:0]   _zz_4911;
  wire       [31:0]   _zz_4912;
  wire       [31:0]   _zz_4913;
  wire       [31:0]   _zz_4914;
  wire       [31:0]   _zz_4915;
  wire       [31:0]   _zz_4916;
  wire       [31:0]   _zz_4917;
  wire       [31:0]   _zz_4918;
  wire       [31:0]   _zz_4919;
  wire       [31:0]   _zz_4920;
  wire       [31:0]   _zz_4921;
  wire       [31:0]   _zz_4922;
  wire       [31:0]   _zz_4923;
  wire       [31:0]   _zz_4924;
  wire       [31:0]   _zz_4925;
  wire       [31:0]   _zz_4926;
  wire       [31:0]   _zz_4927;
  wire       [31:0]   _zz_4928;
  wire       [31:0]   fixTo_dout;
  wire       [31:0]   fixTo_1_dout;
  wire       [15:0]   fixTo_2_dout;
  wire       [15:0]   fixTo_3_dout;
  wire       [15:0]   fixTo_4_dout;
  wire       [15:0]   fixTo_5_dout;
  wire       [31:0]   fixTo_6_dout;
  wire       [31:0]   fixTo_7_dout;
  wire       [15:0]   fixTo_8_dout;
  wire       [15:0]   fixTo_9_dout;
  wire       [15:0]   fixTo_10_dout;
  wire       [15:0]   fixTo_11_dout;
  wire       [31:0]   fixTo_12_dout;
  wire       [31:0]   fixTo_13_dout;
  wire       [15:0]   fixTo_14_dout;
  wire       [15:0]   fixTo_15_dout;
  wire       [15:0]   fixTo_16_dout;
  wire       [15:0]   fixTo_17_dout;
  wire       [31:0]   fixTo_18_dout;
  wire       [31:0]   fixTo_19_dout;
  wire       [15:0]   fixTo_20_dout;
  wire       [15:0]   fixTo_21_dout;
  wire       [15:0]   fixTo_22_dout;
  wire       [15:0]   fixTo_23_dout;
  wire       [31:0]   fixTo_24_dout;
  wire       [31:0]   fixTo_25_dout;
  wire       [15:0]   fixTo_26_dout;
  wire       [15:0]   fixTo_27_dout;
  wire       [15:0]   fixTo_28_dout;
  wire       [15:0]   fixTo_29_dout;
  wire       [31:0]   fixTo_30_dout;
  wire       [31:0]   fixTo_31_dout;
  wire       [15:0]   fixTo_32_dout;
  wire       [15:0]   fixTo_33_dout;
  wire       [15:0]   fixTo_34_dout;
  wire       [15:0]   fixTo_35_dout;
  wire       [31:0]   fixTo_36_dout;
  wire       [31:0]   fixTo_37_dout;
  wire       [15:0]   fixTo_38_dout;
  wire       [15:0]   fixTo_39_dout;
  wire       [15:0]   fixTo_40_dout;
  wire       [15:0]   fixTo_41_dout;
  wire       [31:0]   fixTo_42_dout;
  wire       [31:0]   fixTo_43_dout;
  wire       [15:0]   fixTo_44_dout;
  wire       [15:0]   fixTo_45_dout;
  wire       [15:0]   fixTo_46_dout;
  wire       [15:0]   fixTo_47_dout;
  wire       [31:0]   fixTo_48_dout;
  wire       [31:0]   fixTo_49_dout;
  wire       [15:0]   fixTo_50_dout;
  wire       [15:0]   fixTo_51_dout;
  wire       [15:0]   fixTo_52_dout;
  wire       [15:0]   fixTo_53_dout;
  wire       [31:0]   fixTo_54_dout;
  wire       [31:0]   fixTo_55_dout;
  wire       [15:0]   fixTo_56_dout;
  wire       [15:0]   fixTo_57_dout;
  wire       [15:0]   fixTo_58_dout;
  wire       [15:0]   fixTo_59_dout;
  wire       [31:0]   fixTo_60_dout;
  wire       [31:0]   fixTo_61_dout;
  wire       [15:0]   fixTo_62_dout;
  wire       [15:0]   fixTo_63_dout;
  wire       [15:0]   fixTo_64_dout;
  wire       [15:0]   fixTo_65_dout;
  wire       [31:0]   fixTo_66_dout;
  wire       [31:0]   fixTo_67_dout;
  wire       [15:0]   fixTo_68_dout;
  wire       [15:0]   fixTo_69_dout;
  wire       [15:0]   fixTo_70_dout;
  wire       [15:0]   fixTo_71_dout;
  wire       [31:0]   fixTo_72_dout;
  wire       [31:0]   fixTo_73_dout;
  wire       [15:0]   fixTo_74_dout;
  wire       [15:0]   fixTo_75_dout;
  wire       [15:0]   fixTo_76_dout;
  wire       [15:0]   fixTo_77_dout;
  wire       [31:0]   fixTo_78_dout;
  wire       [31:0]   fixTo_79_dout;
  wire       [15:0]   fixTo_80_dout;
  wire       [15:0]   fixTo_81_dout;
  wire       [15:0]   fixTo_82_dout;
  wire       [15:0]   fixTo_83_dout;
  wire       [31:0]   fixTo_84_dout;
  wire       [31:0]   fixTo_85_dout;
  wire       [15:0]   fixTo_86_dout;
  wire       [15:0]   fixTo_87_dout;
  wire       [15:0]   fixTo_88_dout;
  wire       [15:0]   fixTo_89_dout;
  wire       [31:0]   fixTo_90_dout;
  wire       [31:0]   fixTo_91_dout;
  wire       [15:0]   fixTo_92_dout;
  wire       [15:0]   fixTo_93_dout;
  wire       [15:0]   fixTo_94_dout;
  wire       [15:0]   fixTo_95_dout;
  wire       [31:0]   fixTo_96_dout;
  wire       [31:0]   fixTo_97_dout;
  wire       [15:0]   fixTo_98_dout;
  wire       [15:0]   fixTo_99_dout;
  wire       [15:0]   fixTo_100_dout;
  wire       [15:0]   fixTo_101_dout;
  wire       [31:0]   fixTo_102_dout;
  wire       [31:0]   fixTo_103_dout;
  wire       [15:0]   fixTo_104_dout;
  wire       [15:0]   fixTo_105_dout;
  wire       [15:0]   fixTo_106_dout;
  wire       [15:0]   fixTo_107_dout;
  wire       [31:0]   fixTo_108_dout;
  wire       [31:0]   fixTo_109_dout;
  wire       [15:0]   fixTo_110_dout;
  wire       [15:0]   fixTo_111_dout;
  wire       [15:0]   fixTo_112_dout;
  wire       [15:0]   fixTo_113_dout;
  wire       [31:0]   fixTo_114_dout;
  wire       [31:0]   fixTo_115_dout;
  wire       [15:0]   fixTo_116_dout;
  wire       [15:0]   fixTo_117_dout;
  wire       [15:0]   fixTo_118_dout;
  wire       [15:0]   fixTo_119_dout;
  wire       [31:0]   fixTo_120_dout;
  wire       [31:0]   fixTo_121_dout;
  wire       [15:0]   fixTo_122_dout;
  wire       [15:0]   fixTo_123_dout;
  wire       [15:0]   fixTo_124_dout;
  wire       [15:0]   fixTo_125_dout;
  wire       [31:0]   fixTo_126_dout;
  wire       [31:0]   fixTo_127_dout;
  wire       [15:0]   fixTo_128_dout;
  wire       [15:0]   fixTo_129_dout;
  wire       [15:0]   fixTo_130_dout;
  wire       [15:0]   fixTo_131_dout;
  wire       [31:0]   fixTo_132_dout;
  wire       [31:0]   fixTo_133_dout;
  wire       [15:0]   fixTo_134_dout;
  wire       [15:0]   fixTo_135_dout;
  wire       [15:0]   fixTo_136_dout;
  wire       [15:0]   fixTo_137_dout;
  wire       [31:0]   fixTo_138_dout;
  wire       [31:0]   fixTo_139_dout;
  wire       [15:0]   fixTo_140_dout;
  wire       [15:0]   fixTo_141_dout;
  wire       [15:0]   fixTo_142_dout;
  wire       [15:0]   fixTo_143_dout;
  wire       [31:0]   fixTo_144_dout;
  wire       [31:0]   fixTo_145_dout;
  wire       [15:0]   fixTo_146_dout;
  wire       [15:0]   fixTo_147_dout;
  wire       [15:0]   fixTo_148_dout;
  wire       [15:0]   fixTo_149_dout;
  wire       [31:0]   fixTo_150_dout;
  wire       [31:0]   fixTo_151_dout;
  wire       [15:0]   fixTo_152_dout;
  wire       [15:0]   fixTo_153_dout;
  wire       [15:0]   fixTo_154_dout;
  wire       [15:0]   fixTo_155_dout;
  wire       [31:0]   fixTo_156_dout;
  wire       [31:0]   fixTo_157_dout;
  wire       [15:0]   fixTo_158_dout;
  wire       [15:0]   fixTo_159_dout;
  wire       [15:0]   fixTo_160_dout;
  wire       [15:0]   fixTo_161_dout;
  wire       [31:0]   fixTo_162_dout;
  wire       [31:0]   fixTo_163_dout;
  wire       [15:0]   fixTo_164_dout;
  wire       [15:0]   fixTo_165_dout;
  wire       [15:0]   fixTo_166_dout;
  wire       [15:0]   fixTo_167_dout;
  wire       [31:0]   fixTo_168_dout;
  wire       [31:0]   fixTo_169_dout;
  wire       [15:0]   fixTo_170_dout;
  wire       [15:0]   fixTo_171_dout;
  wire       [15:0]   fixTo_172_dout;
  wire       [15:0]   fixTo_173_dout;
  wire       [31:0]   fixTo_174_dout;
  wire       [31:0]   fixTo_175_dout;
  wire       [15:0]   fixTo_176_dout;
  wire       [15:0]   fixTo_177_dout;
  wire       [15:0]   fixTo_178_dout;
  wire       [15:0]   fixTo_179_dout;
  wire       [31:0]   fixTo_180_dout;
  wire       [31:0]   fixTo_181_dout;
  wire       [15:0]   fixTo_182_dout;
  wire       [15:0]   fixTo_183_dout;
  wire       [15:0]   fixTo_184_dout;
  wire       [15:0]   fixTo_185_dout;
  wire       [31:0]   fixTo_186_dout;
  wire       [31:0]   fixTo_187_dout;
  wire       [15:0]   fixTo_188_dout;
  wire       [15:0]   fixTo_189_dout;
  wire       [15:0]   fixTo_190_dout;
  wire       [15:0]   fixTo_191_dout;
  wire       [31:0]   fixTo_192_dout;
  wire       [31:0]   fixTo_193_dout;
  wire       [15:0]   fixTo_194_dout;
  wire       [15:0]   fixTo_195_dout;
  wire       [15:0]   fixTo_196_dout;
  wire       [15:0]   fixTo_197_dout;
  wire       [31:0]   fixTo_198_dout;
  wire       [31:0]   fixTo_199_dout;
  wire       [15:0]   fixTo_200_dout;
  wire       [15:0]   fixTo_201_dout;
  wire       [15:0]   fixTo_202_dout;
  wire       [15:0]   fixTo_203_dout;
  wire       [31:0]   fixTo_204_dout;
  wire       [31:0]   fixTo_205_dout;
  wire       [15:0]   fixTo_206_dout;
  wire       [15:0]   fixTo_207_dout;
  wire       [15:0]   fixTo_208_dout;
  wire       [15:0]   fixTo_209_dout;
  wire       [31:0]   fixTo_210_dout;
  wire       [31:0]   fixTo_211_dout;
  wire       [15:0]   fixTo_212_dout;
  wire       [15:0]   fixTo_213_dout;
  wire       [15:0]   fixTo_214_dout;
  wire       [15:0]   fixTo_215_dout;
  wire       [31:0]   fixTo_216_dout;
  wire       [31:0]   fixTo_217_dout;
  wire       [15:0]   fixTo_218_dout;
  wire       [15:0]   fixTo_219_dout;
  wire       [15:0]   fixTo_220_dout;
  wire       [15:0]   fixTo_221_dout;
  wire       [31:0]   fixTo_222_dout;
  wire       [31:0]   fixTo_223_dout;
  wire       [15:0]   fixTo_224_dout;
  wire       [15:0]   fixTo_225_dout;
  wire       [15:0]   fixTo_226_dout;
  wire       [15:0]   fixTo_227_dout;
  wire       [31:0]   fixTo_228_dout;
  wire       [31:0]   fixTo_229_dout;
  wire       [15:0]   fixTo_230_dout;
  wire       [15:0]   fixTo_231_dout;
  wire       [15:0]   fixTo_232_dout;
  wire       [15:0]   fixTo_233_dout;
  wire       [31:0]   fixTo_234_dout;
  wire       [31:0]   fixTo_235_dout;
  wire       [15:0]   fixTo_236_dout;
  wire       [15:0]   fixTo_237_dout;
  wire       [15:0]   fixTo_238_dout;
  wire       [15:0]   fixTo_239_dout;
  wire       [31:0]   fixTo_240_dout;
  wire       [31:0]   fixTo_241_dout;
  wire       [15:0]   fixTo_242_dout;
  wire       [15:0]   fixTo_243_dout;
  wire       [15:0]   fixTo_244_dout;
  wire       [15:0]   fixTo_245_dout;
  wire       [31:0]   fixTo_246_dout;
  wire       [31:0]   fixTo_247_dout;
  wire       [15:0]   fixTo_248_dout;
  wire       [15:0]   fixTo_249_dout;
  wire       [15:0]   fixTo_250_dout;
  wire       [15:0]   fixTo_251_dout;
  wire       [31:0]   fixTo_252_dout;
  wire       [31:0]   fixTo_253_dout;
  wire       [15:0]   fixTo_254_dout;
  wire       [15:0]   fixTo_255_dout;
  wire       [15:0]   fixTo_256_dout;
  wire       [15:0]   fixTo_257_dout;
  wire       [31:0]   fixTo_258_dout;
  wire       [31:0]   fixTo_259_dout;
  wire       [15:0]   fixTo_260_dout;
  wire       [15:0]   fixTo_261_dout;
  wire       [15:0]   fixTo_262_dout;
  wire       [15:0]   fixTo_263_dout;
  wire       [31:0]   fixTo_264_dout;
  wire       [31:0]   fixTo_265_dout;
  wire       [15:0]   fixTo_266_dout;
  wire       [15:0]   fixTo_267_dout;
  wire       [15:0]   fixTo_268_dout;
  wire       [15:0]   fixTo_269_dout;
  wire       [31:0]   fixTo_270_dout;
  wire       [31:0]   fixTo_271_dout;
  wire       [15:0]   fixTo_272_dout;
  wire       [15:0]   fixTo_273_dout;
  wire       [15:0]   fixTo_274_dout;
  wire       [15:0]   fixTo_275_dout;
  wire       [31:0]   fixTo_276_dout;
  wire       [31:0]   fixTo_277_dout;
  wire       [15:0]   fixTo_278_dout;
  wire       [15:0]   fixTo_279_dout;
  wire       [15:0]   fixTo_280_dout;
  wire       [15:0]   fixTo_281_dout;
  wire       [31:0]   fixTo_282_dout;
  wire       [31:0]   fixTo_283_dout;
  wire       [15:0]   fixTo_284_dout;
  wire       [15:0]   fixTo_285_dout;
  wire       [15:0]   fixTo_286_dout;
  wire       [15:0]   fixTo_287_dout;
  wire       [31:0]   fixTo_288_dout;
  wire       [31:0]   fixTo_289_dout;
  wire       [15:0]   fixTo_290_dout;
  wire       [15:0]   fixTo_291_dout;
  wire       [15:0]   fixTo_292_dout;
  wire       [15:0]   fixTo_293_dout;
  wire       [31:0]   fixTo_294_dout;
  wire       [31:0]   fixTo_295_dout;
  wire       [15:0]   fixTo_296_dout;
  wire       [15:0]   fixTo_297_dout;
  wire       [15:0]   fixTo_298_dout;
  wire       [15:0]   fixTo_299_dout;
  wire       [31:0]   fixTo_300_dout;
  wire       [31:0]   fixTo_301_dout;
  wire       [15:0]   fixTo_302_dout;
  wire       [15:0]   fixTo_303_dout;
  wire       [15:0]   fixTo_304_dout;
  wire       [15:0]   fixTo_305_dout;
  wire       [31:0]   fixTo_306_dout;
  wire       [31:0]   fixTo_307_dout;
  wire       [15:0]   fixTo_308_dout;
  wire       [15:0]   fixTo_309_dout;
  wire       [15:0]   fixTo_310_dout;
  wire       [15:0]   fixTo_311_dout;
  wire       [31:0]   fixTo_312_dout;
  wire       [31:0]   fixTo_313_dout;
  wire       [15:0]   fixTo_314_dout;
  wire       [15:0]   fixTo_315_dout;
  wire       [15:0]   fixTo_316_dout;
  wire       [15:0]   fixTo_317_dout;
  wire       [31:0]   fixTo_318_dout;
  wire       [31:0]   fixTo_319_dout;
  wire       [15:0]   fixTo_320_dout;
  wire       [15:0]   fixTo_321_dout;
  wire       [15:0]   fixTo_322_dout;
  wire       [15:0]   fixTo_323_dout;
  wire       [31:0]   fixTo_324_dout;
  wire       [31:0]   fixTo_325_dout;
  wire       [15:0]   fixTo_326_dout;
  wire       [15:0]   fixTo_327_dout;
  wire       [15:0]   fixTo_328_dout;
  wire       [15:0]   fixTo_329_dout;
  wire       [31:0]   fixTo_330_dout;
  wire       [31:0]   fixTo_331_dout;
  wire       [15:0]   fixTo_332_dout;
  wire       [15:0]   fixTo_333_dout;
  wire       [15:0]   fixTo_334_dout;
  wire       [15:0]   fixTo_335_dout;
  wire       [31:0]   fixTo_336_dout;
  wire       [31:0]   fixTo_337_dout;
  wire       [15:0]   fixTo_338_dout;
  wire       [15:0]   fixTo_339_dout;
  wire       [15:0]   fixTo_340_dout;
  wire       [15:0]   fixTo_341_dout;
  wire       [31:0]   fixTo_342_dout;
  wire       [31:0]   fixTo_343_dout;
  wire       [15:0]   fixTo_344_dout;
  wire       [15:0]   fixTo_345_dout;
  wire       [15:0]   fixTo_346_dout;
  wire       [15:0]   fixTo_347_dout;
  wire       [31:0]   fixTo_348_dout;
  wire       [31:0]   fixTo_349_dout;
  wire       [15:0]   fixTo_350_dout;
  wire       [15:0]   fixTo_351_dout;
  wire       [15:0]   fixTo_352_dout;
  wire       [15:0]   fixTo_353_dout;
  wire       [31:0]   fixTo_354_dout;
  wire       [31:0]   fixTo_355_dout;
  wire       [15:0]   fixTo_356_dout;
  wire       [15:0]   fixTo_357_dout;
  wire       [15:0]   fixTo_358_dout;
  wire       [15:0]   fixTo_359_dout;
  wire       [31:0]   fixTo_360_dout;
  wire       [31:0]   fixTo_361_dout;
  wire       [15:0]   fixTo_362_dout;
  wire       [15:0]   fixTo_363_dout;
  wire       [15:0]   fixTo_364_dout;
  wire       [15:0]   fixTo_365_dout;
  wire       [31:0]   fixTo_366_dout;
  wire       [31:0]   fixTo_367_dout;
  wire       [15:0]   fixTo_368_dout;
  wire       [15:0]   fixTo_369_dout;
  wire       [15:0]   fixTo_370_dout;
  wire       [15:0]   fixTo_371_dout;
  wire       [31:0]   fixTo_372_dout;
  wire       [31:0]   fixTo_373_dout;
  wire       [15:0]   fixTo_374_dout;
  wire       [15:0]   fixTo_375_dout;
  wire       [15:0]   fixTo_376_dout;
  wire       [15:0]   fixTo_377_dout;
  wire       [31:0]   fixTo_378_dout;
  wire       [31:0]   fixTo_379_dout;
  wire       [15:0]   fixTo_380_dout;
  wire       [15:0]   fixTo_381_dout;
  wire       [15:0]   fixTo_382_dout;
  wire       [15:0]   fixTo_383_dout;
  wire       [31:0]   fixTo_384_dout;
  wire       [31:0]   fixTo_385_dout;
  wire       [15:0]   fixTo_386_dout;
  wire       [15:0]   fixTo_387_dout;
  wire       [15:0]   fixTo_388_dout;
  wire       [15:0]   fixTo_389_dout;
  wire       [31:0]   fixTo_390_dout;
  wire       [31:0]   fixTo_391_dout;
  wire       [15:0]   fixTo_392_dout;
  wire       [15:0]   fixTo_393_dout;
  wire       [15:0]   fixTo_394_dout;
  wire       [15:0]   fixTo_395_dout;
  wire       [31:0]   fixTo_396_dout;
  wire       [31:0]   fixTo_397_dout;
  wire       [15:0]   fixTo_398_dout;
  wire       [15:0]   fixTo_399_dout;
  wire       [15:0]   fixTo_400_dout;
  wire       [15:0]   fixTo_401_dout;
  wire       [31:0]   fixTo_402_dout;
  wire       [31:0]   fixTo_403_dout;
  wire       [15:0]   fixTo_404_dout;
  wire       [15:0]   fixTo_405_dout;
  wire       [15:0]   fixTo_406_dout;
  wire       [15:0]   fixTo_407_dout;
  wire       [31:0]   fixTo_408_dout;
  wire       [31:0]   fixTo_409_dout;
  wire       [15:0]   fixTo_410_dout;
  wire       [15:0]   fixTo_411_dout;
  wire       [15:0]   fixTo_412_dout;
  wire       [15:0]   fixTo_413_dout;
  wire       [31:0]   fixTo_414_dout;
  wire       [31:0]   fixTo_415_dout;
  wire       [15:0]   fixTo_416_dout;
  wire       [15:0]   fixTo_417_dout;
  wire       [15:0]   fixTo_418_dout;
  wire       [15:0]   fixTo_419_dout;
  wire       [31:0]   fixTo_420_dout;
  wire       [31:0]   fixTo_421_dout;
  wire       [15:0]   fixTo_422_dout;
  wire       [15:0]   fixTo_423_dout;
  wire       [15:0]   fixTo_424_dout;
  wire       [15:0]   fixTo_425_dout;
  wire       [31:0]   fixTo_426_dout;
  wire       [31:0]   fixTo_427_dout;
  wire       [15:0]   fixTo_428_dout;
  wire       [15:0]   fixTo_429_dout;
  wire       [15:0]   fixTo_430_dout;
  wire       [15:0]   fixTo_431_dout;
  wire       [31:0]   fixTo_432_dout;
  wire       [31:0]   fixTo_433_dout;
  wire       [15:0]   fixTo_434_dout;
  wire       [15:0]   fixTo_435_dout;
  wire       [15:0]   fixTo_436_dout;
  wire       [15:0]   fixTo_437_dout;
  wire       [31:0]   fixTo_438_dout;
  wire       [31:0]   fixTo_439_dout;
  wire       [15:0]   fixTo_440_dout;
  wire       [15:0]   fixTo_441_dout;
  wire       [15:0]   fixTo_442_dout;
  wire       [15:0]   fixTo_443_dout;
  wire       [31:0]   fixTo_444_dout;
  wire       [31:0]   fixTo_445_dout;
  wire       [15:0]   fixTo_446_dout;
  wire       [15:0]   fixTo_447_dout;
  wire       [15:0]   fixTo_448_dout;
  wire       [15:0]   fixTo_449_dout;
  wire       [31:0]   fixTo_450_dout;
  wire       [31:0]   fixTo_451_dout;
  wire       [15:0]   fixTo_452_dout;
  wire       [15:0]   fixTo_453_dout;
  wire       [15:0]   fixTo_454_dout;
  wire       [15:0]   fixTo_455_dout;
  wire       [31:0]   fixTo_456_dout;
  wire       [31:0]   fixTo_457_dout;
  wire       [15:0]   fixTo_458_dout;
  wire       [15:0]   fixTo_459_dout;
  wire       [15:0]   fixTo_460_dout;
  wire       [15:0]   fixTo_461_dout;
  wire       [31:0]   fixTo_462_dout;
  wire       [31:0]   fixTo_463_dout;
  wire       [15:0]   fixTo_464_dout;
  wire       [15:0]   fixTo_465_dout;
  wire       [15:0]   fixTo_466_dout;
  wire       [15:0]   fixTo_467_dout;
  wire       [31:0]   fixTo_468_dout;
  wire       [31:0]   fixTo_469_dout;
  wire       [15:0]   fixTo_470_dout;
  wire       [15:0]   fixTo_471_dout;
  wire       [15:0]   fixTo_472_dout;
  wire       [15:0]   fixTo_473_dout;
  wire       [31:0]   fixTo_474_dout;
  wire       [31:0]   fixTo_475_dout;
  wire       [15:0]   fixTo_476_dout;
  wire       [15:0]   fixTo_477_dout;
  wire       [15:0]   fixTo_478_dout;
  wire       [15:0]   fixTo_479_dout;
  wire       [31:0]   fixTo_480_dout;
  wire       [31:0]   fixTo_481_dout;
  wire       [15:0]   fixTo_482_dout;
  wire       [15:0]   fixTo_483_dout;
  wire       [15:0]   fixTo_484_dout;
  wire       [15:0]   fixTo_485_dout;
  wire       [31:0]   fixTo_486_dout;
  wire       [31:0]   fixTo_487_dout;
  wire       [15:0]   fixTo_488_dout;
  wire       [15:0]   fixTo_489_dout;
  wire       [15:0]   fixTo_490_dout;
  wire       [15:0]   fixTo_491_dout;
  wire       [31:0]   fixTo_492_dout;
  wire       [31:0]   fixTo_493_dout;
  wire       [15:0]   fixTo_494_dout;
  wire       [15:0]   fixTo_495_dout;
  wire       [15:0]   fixTo_496_dout;
  wire       [15:0]   fixTo_497_dout;
  wire       [31:0]   fixTo_498_dout;
  wire       [31:0]   fixTo_499_dout;
  wire       [15:0]   fixTo_500_dout;
  wire       [15:0]   fixTo_501_dout;
  wire       [15:0]   fixTo_502_dout;
  wire       [15:0]   fixTo_503_dout;
  wire       [31:0]   fixTo_504_dout;
  wire       [31:0]   fixTo_505_dout;
  wire       [15:0]   fixTo_506_dout;
  wire       [15:0]   fixTo_507_dout;
  wire       [15:0]   fixTo_508_dout;
  wire       [15:0]   fixTo_509_dout;
  wire       [31:0]   fixTo_510_dout;
  wire       [31:0]   fixTo_511_dout;
  wire       [15:0]   fixTo_512_dout;
  wire       [15:0]   fixTo_513_dout;
  wire       [15:0]   fixTo_514_dout;
  wire       [15:0]   fixTo_515_dout;
  wire       [31:0]   fixTo_516_dout;
  wire       [31:0]   fixTo_517_dout;
  wire       [15:0]   fixTo_518_dout;
  wire       [15:0]   fixTo_519_dout;
  wire       [15:0]   fixTo_520_dout;
  wire       [15:0]   fixTo_521_dout;
  wire       [31:0]   fixTo_522_dout;
  wire       [31:0]   fixTo_523_dout;
  wire       [15:0]   fixTo_524_dout;
  wire       [15:0]   fixTo_525_dout;
  wire       [15:0]   fixTo_526_dout;
  wire       [15:0]   fixTo_527_dout;
  wire       [31:0]   fixTo_528_dout;
  wire       [31:0]   fixTo_529_dout;
  wire       [15:0]   fixTo_530_dout;
  wire       [15:0]   fixTo_531_dout;
  wire       [15:0]   fixTo_532_dout;
  wire       [15:0]   fixTo_533_dout;
  wire       [31:0]   fixTo_534_dout;
  wire       [31:0]   fixTo_535_dout;
  wire       [15:0]   fixTo_536_dout;
  wire       [15:0]   fixTo_537_dout;
  wire       [15:0]   fixTo_538_dout;
  wire       [15:0]   fixTo_539_dout;
  wire       [31:0]   fixTo_540_dout;
  wire       [31:0]   fixTo_541_dout;
  wire       [15:0]   fixTo_542_dout;
  wire       [15:0]   fixTo_543_dout;
  wire       [15:0]   fixTo_544_dout;
  wire       [15:0]   fixTo_545_dout;
  wire       [31:0]   fixTo_546_dout;
  wire       [31:0]   fixTo_547_dout;
  wire       [15:0]   fixTo_548_dout;
  wire       [15:0]   fixTo_549_dout;
  wire       [15:0]   fixTo_550_dout;
  wire       [15:0]   fixTo_551_dout;
  wire       [31:0]   fixTo_552_dout;
  wire       [31:0]   fixTo_553_dout;
  wire       [15:0]   fixTo_554_dout;
  wire       [15:0]   fixTo_555_dout;
  wire       [15:0]   fixTo_556_dout;
  wire       [15:0]   fixTo_557_dout;
  wire       [31:0]   fixTo_558_dout;
  wire       [31:0]   fixTo_559_dout;
  wire       [15:0]   fixTo_560_dout;
  wire       [15:0]   fixTo_561_dout;
  wire       [15:0]   fixTo_562_dout;
  wire       [15:0]   fixTo_563_dout;
  wire       [31:0]   fixTo_564_dout;
  wire       [31:0]   fixTo_565_dout;
  wire       [15:0]   fixTo_566_dout;
  wire       [15:0]   fixTo_567_dout;
  wire       [15:0]   fixTo_568_dout;
  wire       [15:0]   fixTo_569_dout;
  wire       [31:0]   fixTo_570_dout;
  wire       [31:0]   fixTo_571_dout;
  wire       [15:0]   fixTo_572_dout;
  wire       [15:0]   fixTo_573_dout;
  wire       [15:0]   fixTo_574_dout;
  wire       [15:0]   fixTo_575_dout;
  wire       [31:0]   fixTo_576_dout;
  wire       [31:0]   fixTo_577_dout;
  wire       [15:0]   fixTo_578_dout;
  wire       [15:0]   fixTo_579_dout;
  wire       [15:0]   fixTo_580_dout;
  wire       [15:0]   fixTo_581_dout;
  wire       [31:0]   fixTo_582_dout;
  wire       [31:0]   fixTo_583_dout;
  wire       [15:0]   fixTo_584_dout;
  wire       [15:0]   fixTo_585_dout;
  wire       [15:0]   fixTo_586_dout;
  wire       [15:0]   fixTo_587_dout;
  wire       [31:0]   fixTo_588_dout;
  wire       [31:0]   fixTo_589_dout;
  wire       [15:0]   fixTo_590_dout;
  wire       [15:0]   fixTo_591_dout;
  wire       [15:0]   fixTo_592_dout;
  wire       [15:0]   fixTo_593_dout;
  wire       [31:0]   fixTo_594_dout;
  wire       [31:0]   fixTo_595_dout;
  wire       [15:0]   fixTo_596_dout;
  wire       [15:0]   fixTo_597_dout;
  wire       [15:0]   fixTo_598_dout;
  wire       [15:0]   fixTo_599_dout;
  wire       [31:0]   fixTo_600_dout;
  wire       [31:0]   fixTo_601_dout;
  wire       [15:0]   fixTo_602_dout;
  wire       [15:0]   fixTo_603_dout;
  wire       [15:0]   fixTo_604_dout;
  wire       [15:0]   fixTo_605_dout;
  wire       [31:0]   fixTo_606_dout;
  wire       [31:0]   fixTo_607_dout;
  wire       [15:0]   fixTo_608_dout;
  wire       [15:0]   fixTo_609_dout;
  wire       [15:0]   fixTo_610_dout;
  wire       [15:0]   fixTo_611_dout;
  wire       [31:0]   fixTo_612_dout;
  wire       [31:0]   fixTo_613_dout;
  wire       [15:0]   fixTo_614_dout;
  wire       [15:0]   fixTo_615_dout;
  wire       [15:0]   fixTo_616_dout;
  wire       [15:0]   fixTo_617_dout;
  wire       [31:0]   fixTo_618_dout;
  wire       [31:0]   fixTo_619_dout;
  wire       [15:0]   fixTo_620_dout;
  wire       [15:0]   fixTo_621_dout;
  wire       [15:0]   fixTo_622_dout;
  wire       [15:0]   fixTo_623_dout;
  wire       [31:0]   fixTo_624_dout;
  wire       [31:0]   fixTo_625_dout;
  wire       [15:0]   fixTo_626_dout;
  wire       [15:0]   fixTo_627_dout;
  wire       [15:0]   fixTo_628_dout;
  wire       [15:0]   fixTo_629_dout;
  wire       [31:0]   fixTo_630_dout;
  wire       [31:0]   fixTo_631_dout;
  wire       [15:0]   fixTo_632_dout;
  wire       [15:0]   fixTo_633_dout;
  wire       [15:0]   fixTo_634_dout;
  wire       [15:0]   fixTo_635_dout;
  wire       [31:0]   fixTo_636_dout;
  wire       [31:0]   fixTo_637_dout;
  wire       [15:0]   fixTo_638_dout;
  wire       [15:0]   fixTo_639_dout;
  wire       [15:0]   fixTo_640_dout;
  wire       [15:0]   fixTo_641_dout;
  wire       [31:0]   fixTo_642_dout;
  wire       [31:0]   fixTo_643_dout;
  wire       [15:0]   fixTo_644_dout;
  wire       [15:0]   fixTo_645_dout;
  wire       [15:0]   fixTo_646_dout;
  wire       [15:0]   fixTo_647_dout;
  wire       [31:0]   fixTo_648_dout;
  wire       [31:0]   fixTo_649_dout;
  wire       [15:0]   fixTo_650_dout;
  wire       [15:0]   fixTo_651_dout;
  wire       [15:0]   fixTo_652_dout;
  wire       [15:0]   fixTo_653_dout;
  wire       [31:0]   fixTo_654_dout;
  wire       [31:0]   fixTo_655_dout;
  wire       [15:0]   fixTo_656_dout;
  wire       [15:0]   fixTo_657_dout;
  wire       [15:0]   fixTo_658_dout;
  wire       [15:0]   fixTo_659_dout;
  wire       [31:0]   fixTo_660_dout;
  wire       [31:0]   fixTo_661_dout;
  wire       [15:0]   fixTo_662_dout;
  wire       [15:0]   fixTo_663_dout;
  wire       [15:0]   fixTo_664_dout;
  wire       [15:0]   fixTo_665_dout;
  wire       [31:0]   fixTo_666_dout;
  wire       [31:0]   fixTo_667_dout;
  wire       [15:0]   fixTo_668_dout;
  wire       [15:0]   fixTo_669_dout;
  wire       [15:0]   fixTo_670_dout;
  wire       [15:0]   fixTo_671_dout;
  wire       [31:0]   fixTo_672_dout;
  wire       [31:0]   fixTo_673_dout;
  wire       [15:0]   fixTo_674_dout;
  wire       [15:0]   fixTo_675_dout;
  wire       [15:0]   fixTo_676_dout;
  wire       [15:0]   fixTo_677_dout;
  wire       [31:0]   fixTo_678_dout;
  wire       [31:0]   fixTo_679_dout;
  wire       [15:0]   fixTo_680_dout;
  wire       [15:0]   fixTo_681_dout;
  wire       [15:0]   fixTo_682_dout;
  wire       [15:0]   fixTo_683_dout;
  wire       [31:0]   fixTo_684_dout;
  wire       [31:0]   fixTo_685_dout;
  wire       [15:0]   fixTo_686_dout;
  wire       [15:0]   fixTo_687_dout;
  wire       [15:0]   fixTo_688_dout;
  wire       [15:0]   fixTo_689_dout;
  wire       [31:0]   fixTo_690_dout;
  wire       [31:0]   fixTo_691_dout;
  wire       [15:0]   fixTo_692_dout;
  wire       [15:0]   fixTo_693_dout;
  wire       [15:0]   fixTo_694_dout;
  wire       [15:0]   fixTo_695_dout;
  wire       [31:0]   fixTo_696_dout;
  wire       [31:0]   fixTo_697_dout;
  wire       [15:0]   fixTo_698_dout;
  wire       [15:0]   fixTo_699_dout;
  wire       [15:0]   fixTo_700_dout;
  wire       [15:0]   fixTo_701_dout;
  wire       [31:0]   fixTo_702_dout;
  wire       [31:0]   fixTo_703_dout;
  wire       [15:0]   fixTo_704_dout;
  wire       [15:0]   fixTo_705_dout;
  wire       [15:0]   fixTo_706_dout;
  wire       [15:0]   fixTo_707_dout;
  wire       [31:0]   fixTo_708_dout;
  wire       [31:0]   fixTo_709_dout;
  wire       [15:0]   fixTo_710_dout;
  wire       [15:0]   fixTo_711_dout;
  wire       [15:0]   fixTo_712_dout;
  wire       [15:0]   fixTo_713_dout;
  wire       [31:0]   fixTo_714_dout;
  wire       [31:0]   fixTo_715_dout;
  wire       [15:0]   fixTo_716_dout;
  wire       [15:0]   fixTo_717_dout;
  wire       [15:0]   fixTo_718_dout;
  wire       [15:0]   fixTo_719_dout;
  wire       [31:0]   fixTo_720_dout;
  wire       [31:0]   fixTo_721_dout;
  wire       [15:0]   fixTo_722_dout;
  wire       [15:0]   fixTo_723_dout;
  wire       [15:0]   fixTo_724_dout;
  wire       [15:0]   fixTo_725_dout;
  wire       [31:0]   fixTo_726_dout;
  wire       [31:0]   fixTo_727_dout;
  wire       [15:0]   fixTo_728_dout;
  wire       [15:0]   fixTo_729_dout;
  wire       [15:0]   fixTo_730_dout;
  wire       [15:0]   fixTo_731_dout;
  wire       [31:0]   fixTo_732_dout;
  wire       [31:0]   fixTo_733_dout;
  wire       [15:0]   fixTo_734_dout;
  wire       [15:0]   fixTo_735_dout;
  wire       [15:0]   fixTo_736_dout;
  wire       [15:0]   fixTo_737_dout;
  wire       [31:0]   fixTo_738_dout;
  wire       [31:0]   fixTo_739_dout;
  wire       [15:0]   fixTo_740_dout;
  wire       [15:0]   fixTo_741_dout;
  wire       [15:0]   fixTo_742_dout;
  wire       [15:0]   fixTo_743_dout;
  wire       [31:0]   fixTo_744_dout;
  wire       [31:0]   fixTo_745_dout;
  wire       [15:0]   fixTo_746_dout;
  wire       [15:0]   fixTo_747_dout;
  wire       [15:0]   fixTo_748_dout;
  wire       [15:0]   fixTo_749_dout;
  wire       [31:0]   fixTo_750_dout;
  wire       [31:0]   fixTo_751_dout;
  wire       [15:0]   fixTo_752_dout;
  wire       [15:0]   fixTo_753_dout;
  wire       [15:0]   fixTo_754_dout;
  wire       [15:0]   fixTo_755_dout;
  wire       [31:0]   fixTo_756_dout;
  wire       [31:0]   fixTo_757_dout;
  wire       [15:0]   fixTo_758_dout;
  wire       [15:0]   fixTo_759_dout;
  wire       [15:0]   fixTo_760_dout;
  wire       [15:0]   fixTo_761_dout;
  wire       [31:0]   fixTo_762_dout;
  wire       [31:0]   fixTo_763_dout;
  wire       [15:0]   fixTo_764_dout;
  wire       [15:0]   fixTo_765_dout;
  wire       [15:0]   fixTo_766_dout;
  wire       [15:0]   fixTo_767_dout;
  wire       [31:0]   fixTo_768_dout;
  wire       [31:0]   fixTo_769_dout;
  wire       [15:0]   fixTo_770_dout;
  wire       [15:0]   fixTo_771_dout;
  wire       [15:0]   fixTo_772_dout;
  wire       [15:0]   fixTo_773_dout;
  wire       [31:0]   fixTo_774_dout;
  wire       [31:0]   fixTo_775_dout;
  wire       [15:0]   fixTo_776_dout;
  wire       [15:0]   fixTo_777_dout;
  wire       [15:0]   fixTo_778_dout;
  wire       [15:0]   fixTo_779_dout;
  wire       [31:0]   fixTo_780_dout;
  wire       [31:0]   fixTo_781_dout;
  wire       [15:0]   fixTo_782_dout;
  wire       [15:0]   fixTo_783_dout;
  wire       [15:0]   fixTo_784_dout;
  wire       [15:0]   fixTo_785_dout;
  wire       [31:0]   fixTo_786_dout;
  wire       [31:0]   fixTo_787_dout;
  wire       [15:0]   fixTo_788_dout;
  wire       [15:0]   fixTo_789_dout;
  wire       [15:0]   fixTo_790_dout;
  wire       [15:0]   fixTo_791_dout;
  wire       [31:0]   fixTo_792_dout;
  wire       [31:0]   fixTo_793_dout;
  wire       [15:0]   fixTo_794_dout;
  wire       [15:0]   fixTo_795_dout;
  wire       [15:0]   fixTo_796_dout;
  wire       [15:0]   fixTo_797_dout;
  wire       [31:0]   fixTo_798_dout;
  wire       [31:0]   fixTo_799_dout;
  wire       [15:0]   fixTo_800_dout;
  wire       [15:0]   fixTo_801_dout;
  wire       [15:0]   fixTo_802_dout;
  wire       [15:0]   fixTo_803_dout;
  wire       [31:0]   fixTo_804_dout;
  wire       [31:0]   fixTo_805_dout;
  wire       [15:0]   fixTo_806_dout;
  wire       [15:0]   fixTo_807_dout;
  wire       [15:0]   fixTo_808_dout;
  wire       [15:0]   fixTo_809_dout;
  wire       [31:0]   fixTo_810_dout;
  wire       [31:0]   fixTo_811_dout;
  wire       [15:0]   fixTo_812_dout;
  wire       [15:0]   fixTo_813_dout;
  wire       [15:0]   fixTo_814_dout;
  wire       [15:0]   fixTo_815_dout;
  wire       [31:0]   fixTo_816_dout;
  wire       [31:0]   fixTo_817_dout;
  wire       [15:0]   fixTo_818_dout;
  wire       [15:0]   fixTo_819_dout;
  wire       [15:0]   fixTo_820_dout;
  wire       [15:0]   fixTo_821_dout;
  wire       [31:0]   fixTo_822_dout;
  wire       [31:0]   fixTo_823_dout;
  wire       [15:0]   fixTo_824_dout;
  wire       [15:0]   fixTo_825_dout;
  wire       [15:0]   fixTo_826_dout;
  wire       [15:0]   fixTo_827_dout;
  wire       [31:0]   fixTo_828_dout;
  wire       [31:0]   fixTo_829_dout;
  wire       [15:0]   fixTo_830_dout;
  wire       [15:0]   fixTo_831_dout;
  wire       [15:0]   fixTo_832_dout;
  wire       [15:0]   fixTo_833_dout;
  wire       [31:0]   fixTo_834_dout;
  wire       [31:0]   fixTo_835_dout;
  wire       [15:0]   fixTo_836_dout;
  wire       [15:0]   fixTo_837_dout;
  wire       [15:0]   fixTo_838_dout;
  wire       [15:0]   fixTo_839_dout;
  wire       [31:0]   fixTo_840_dout;
  wire       [31:0]   fixTo_841_dout;
  wire       [15:0]   fixTo_842_dout;
  wire       [15:0]   fixTo_843_dout;
  wire       [15:0]   fixTo_844_dout;
  wire       [15:0]   fixTo_845_dout;
  wire       [31:0]   fixTo_846_dout;
  wire       [31:0]   fixTo_847_dout;
  wire       [15:0]   fixTo_848_dout;
  wire       [15:0]   fixTo_849_dout;
  wire       [15:0]   fixTo_850_dout;
  wire       [15:0]   fixTo_851_dout;
  wire       [31:0]   fixTo_852_dout;
  wire       [31:0]   fixTo_853_dout;
  wire       [15:0]   fixTo_854_dout;
  wire       [15:0]   fixTo_855_dout;
  wire       [15:0]   fixTo_856_dout;
  wire       [15:0]   fixTo_857_dout;
  wire       [31:0]   fixTo_858_dout;
  wire       [31:0]   fixTo_859_dout;
  wire       [15:0]   fixTo_860_dout;
  wire       [15:0]   fixTo_861_dout;
  wire       [15:0]   fixTo_862_dout;
  wire       [15:0]   fixTo_863_dout;
  wire       [31:0]   fixTo_864_dout;
  wire       [31:0]   fixTo_865_dout;
  wire       [15:0]   fixTo_866_dout;
  wire       [15:0]   fixTo_867_dout;
  wire       [15:0]   fixTo_868_dout;
  wire       [15:0]   fixTo_869_dout;
  wire       [31:0]   fixTo_870_dout;
  wire       [31:0]   fixTo_871_dout;
  wire       [15:0]   fixTo_872_dout;
  wire       [15:0]   fixTo_873_dout;
  wire       [15:0]   fixTo_874_dout;
  wire       [15:0]   fixTo_875_dout;
  wire       [31:0]   fixTo_876_dout;
  wire       [31:0]   fixTo_877_dout;
  wire       [15:0]   fixTo_878_dout;
  wire       [15:0]   fixTo_879_dout;
  wire       [15:0]   fixTo_880_dout;
  wire       [15:0]   fixTo_881_dout;
  wire       [31:0]   fixTo_882_dout;
  wire       [31:0]   fixTo_883_dout;
  wire       [15:0]   fixTo_884_dout;
  wire       [15:0]   fixTo_885_dout;
  wire       [15:0]   fixTo_886_dout;
  wire       [15:0]   fixTo_887_dout;
  wire       [31:0]   fixTo_888_dout;
  wire       [31:0]   fixTo_889_dout;
  wire       [15:0]   fixTo_890_dout;
  wire       [15:0]   fixTo_891_dout;
  wire       [15:0]   fixTo_892_dout;
  wire       [15:0]   fixTo_893_dout;
  wire       [31:0]   fixTo_894_dout;
  wire       [31:0]   fixTo_895_dout;
  wire       [15:0]   fixTo_896_dout;
  wire       [15:0]   fixTo_897_dout;
  wire       [15:0]   fixTo_898_dout;
  wire       [15:0]   fixTo_899_dout;
  wire       [31:0]   fixTo_900_dout;
  wire       [31:0]   fixTo_901_dout;
  wire       [15:0]   fixTo_902_dout;
  wire       [15:0]   fixTo_903_dout;
  wire       [15:0]   fixTo_904_dout;
  wire       [15:0]   fixTo_905_dout;
  wire       [31:0]   fixTo_906_dout;
  wire       [31:0]   fixTo_907_dout;
  wire       [15:0]   fixTo_908_dout;
  wire       [15:0]   fixTo_909_dout;
  wire       [15:0]   fixTo_910_dout;
  wire       [15:0]   fixTo_911_dout;
  wire       [31:0]   fixTo_912_dout;
  wire       [31:0]   fixTo_913_dout;
  wire       [15:0]   fixTo_914_dout;
  wire       [15:0]   fixTo_915_dout;
  wire       [15:0]   fixTo_916_dout;
  wire       [15:0]   fixTo_917_dout;
  wire       [31:0]   fixTo_918_dout;
  wire       [31:0]   fixTo_919_dout;
  wire       [15:0]   fixTo_920_dout;
  wire       [15:0]   fixTo_921_dout;
  wire       [15:0]   fixTo_922_dout;
  wire       [15:0]   fixTo_923_dout;
  wire       [31:0]   fixTo_924_dout;
  wire       [31:0]   fixTo_925_dout;
  wire       [15:0]   fixTo_926_dout;
  wire       [15:0]   fixTo_927_dout;
  wire       [15:0]   fixTo_928_dout;
  wire       [15:0]   fixTo_929_dout;
  wire       [31:0]   fixTo_930_dout;
  wire       [31:0]   fixTo_931_dout;
  wire       [15:0]   fixTo_932_dout;
  wire       [15:0]   fixTo_933_dout;
  wire       [15:0]   fixTo_934_dout;
  wire       [15:0]   fixTo_935_dout;
  wire       [31:0]   fixTo_936_dout;
  wire       [31:0]   fixTo_937_dout;
  wire       [15:0]   fixTo_938_dout;
  wire       [15:0]   fixTo_939_dout;
  wire       [15:0]   fixTo_940_dout;
  wire       [15:0]   fixTo_941_dout;
  wire       [31:0]   fixTo_942_dout;
  wire       [31:0]   fixTo_943_dout;
  wire       [15:0]   fixTo_944_dout;
  wire       [15:0]   fixTo_945_dout;
  wire       [15:0]   fixTo_946_dout;
  wire       [15:0]   fixTo_947_dout;
  wire       [31:0]   fixTo_948_dout;
  wire       [31:0]   fixTo_949_dout;
  wire       [15:0]   fixTo_950_dout;
  wire       [15:0]   fixTo_951_dout;
  wire       [15:0]   fixTo_952_dout;
  wire       [15:0]   fixTo_953_dout;
  wire       [31:0]   fixTo_954_dout;
  wire       [31:0]   fixTo_955_dout;
  wire       [15:0]   fixTo_956_dout;
  wire       [15:0]   fixTo_957_dout;
  wire       [15:0]   fixTo_958_dout;
  wire       [15:0]   fixTo_959_dout;
  wire       [31:0]   fixTo_960_dout;
  wire       [31:0]   fixTo_961_dout;
  wire       [15:0]   fixTo_962_dout;
  wire       [15:0]   fixTo_963_dout;
  wire       [15:0]   fixTo_964_dout;
  wire       [15:0]   fixTo_965_dout;
  wire       [31:0]   fixTo_966_dout;
  wire       [31:0]   fixTo_967_dout;
  wire       [15:0]   fixTo_968_dout;
  wire       [15:0]   fixTo_969_dout;
  wire       [15:0]   fixTo_970_dout;
  wire       [15:0]   fixTo_971_dout;
  wire       [31:0]   fixTo_972_dout;
  wire       [31:0]   fixTo_973_dout;
  wire       [15:0]   fixTo_974_dout;
  wire       [15:0]   fixTo_975_dout;
  wire       [15:0]   fixTo_976_dout;
  wire       [15:0]   fixTo_977_dout;
  wire       [31:0]   fixTo_978_dout;
  wire       [31:0]   fixTo_979_dout;
  wire       [15:0]   fixTo_980_dout;
  wire       [15:0]   fixTo_981_dout;
  wire       [15:0]   fixTo_982_dout;
  wire       [15:0]   fixTo_983_dout;
  wire       [31:0]   fixTo_984_dout;
  wire       [31:0]   fixTo_985_dout;
  wire       [15:0]   fixTo_986_dout;
  wire       [15:0]   fixTo_987_dout;
  wire       [15:0]   fixTo_988_dout;
  wire       [15:0]   fixTo_989_dout;
  wire       [31:0]   fixTo_990_dout;
  wire       [31:0]   fixTo_991_dout;
  wire       [15:0]   fixTo_992_dout;
  wire       [15:0]   fixTo_993_dout;
  wire       [15:0]   fixTo_994_dout;
  wire       [15:0]   fixTo_995_dout;
  wire       [31:0]   fixTo_996_dout;
  wire       [31:0]   fixTo_997_dout;
  wire       [15:0]   fixTo_998_dout;
  wire       [15:0]   fixTo_999_dout;
  wire       [15:0]   fixTo_1000_dout;
  wire       [15:0]   fixTo_1001_dout;
  wire       [31:0]   fixTo_1002_dout;
  wire       [31:0]   fixTo_1003_dout;
  wire       [15:0]   fixTo_1004_dout;
  wire       [15:0]   fixTo_1005_dout;
  wire       [15:0]   fixTo_1006_dout;
  wire       [15:0]   fixTo_1007_dout;
  wire       [31:0]   fixTo_1008_dout;
  wire       [31:0]   fixTo_1009_dout;
  wire       [15:0]   fixTo_1010_dout;
  wire       [15:0]   fixTo_1011_dout;
  wire       [15:0]   fixTo_1012_dout;
  wire       [15:0]   fixTo_1013_dout;
  wire       [31:0]   fixTo_1014_dout;
  wire       [31:0]   fixTo_1015_dout;
  wire       [15:0]   fixTo_1016_dout;
  wire       [15:0]   fixTo_1017_dout;
  wire       [15:0]   fixTo_1018_dout;
  wire       [15:0]   fixTo_1019_dout;
  wire       [31:0]   fixTo_1020_dout;
  wire       [31:0]   fixTo_1021_dout;
  wire       [15:0]   fixTo_1022_dout;
  wire       [15:0]   fixTo_1023_dout;
  wire       [15:0]   fixTo_1024_dout;
  wire       [15:0]   fixTo_1025_dout;
  wire       [31:0]   fixTo_1026_dout;
  wire       [31:0]   fixTo_1027_dout;
  wire       [15:0]   fixTo_1028_dout;
  wire       [15:0]   fixTo_1029_dout;
  wire       [15:0]   fixTo_1030_dout;
  wire       [15:0]   fixTo_1031_dout;
  wire       [31:0]   fixTo_1032_dout;
  wire       [31:0]   fixTo_1033_dout;
  wire       [15:0]   fixTo_1034_dout;
  wire       [15:0]   fixTo_1035_dout;
  wire       [15:0]   fixTo_1036_dout;
  wire       [15:0]   fixTo_1037_dout;
  wire       [31:0]   fixTo_1038_dout;
  wire       [31:0]   fixTo_1039_dout;
  wire       [15:0]   fixTo_1040_dout;
  wire       [15:0]   fixTo_1041_dout;
  wire       [15:0]   fixTo_1042_dout;
  wire       [15:0]   fixTo_1043_dout;
  wire       [31:0]   fixTo_1044_dout;
  wire       [31:0]   fixTo_1045_dout;
  wire       [15:0]   fixTo_1046_dout;
  wire       [15:0]   fixTo_1047_dout;
  wire       [15:0]   fixTo_1048_dout;
  wire       [15:0]   fixTo_1049_dout;
  wire       [31:0]   fixTo_1050_dout;
  wire       [31:0]   fixTo_1051_dout;
  wire       [15:0]   fixTo_1052_dout;
  wire       [15:0]   fixTo_1053_dout;
  wire       [15:0]   fixTo_1054_dout;
  wire       [15:0]   fixTo_1055_dout;
  wire       [31:0]   fixTo_1056_dout;
  wire       [31:0]   fixTo_1057_dout;
  wire       [15:0]   fixTo_1058_dout;
  wire       [15:0]   fixTo_1059_dout;
  wire       [15:0]   fixTo_1060_dout;
  wire       [15:0]   fixTo_1061_dout;
  wire       [31:0]   fixTo_1062_dout;
  wire       [31:0]   fixTo_1063_dout;
  wire       [15:0]   fixTo_1064_dout;
  wire       [15:0]   fixTo_1065_dout;
  wire       [15:0]   fixTo_1066_dout;
  wire       [15:0]   fixTo_1067_dout;
  wire       [31:0]   fixTo_1068_dout;
  wire       [31:0]   fixTo_1069_dout;
  wire       [15:0]   fixTo_1070_dout;
  wire       [15:0]   fixTo_1071_dout;
  wire       [15:0]   fixTo_1072_dout;
  wire       [15:0]   fixTo_1073_dout;
  wire       [31:0]   fixTo_1074_dout;
  wire       [31:0]   fixTo_1075_dout;
  wire       [15:0]   fixTo_1076_dout;
  wire       [15:0]   fixTo_1077_dout;
  wire       [15:0]   fixTo_1078_dout;
  wire       [15:0]   fixTo_1079_dout;
  wire       [31:0]   fixTo_1080_dout;
  wire       [31:0]   fixTo_1081_dout;
  wire       [15:0]   fixTo_1082_dout;
  wire       [15:0]   fixTo_1083_dout;
  wire       [15:0]   fixTo_1084_dout;
  wire       [15:0]   fixTo_1085_dout;
  wire       [31:0]   fixTo_1086_dout;
  wire       [31:0]   fixTo_1087_dout;
  wire       [15:0]   fixTo_1088_dout;
  wire       [15:0]   fixTo_1089_dout;
  wire       [15:0]   fixTo_1090_dout;
  wire       [15:0]   fixTo_1091_dout;
  wire       [31:0]   fixTo_1092_dout;
  wire       [31:0]   fixTo_1093_dout;
  wire       [15:0]   fixTo_1094_dout;
  wire       [15:0]   fixTo_1095_dout;
  wire       [15:0]   fixTo_1096_dout;
  wire       [15:0]   fixTo_1097_dout;
  wire       [31:0]   fixTo_1098_dout;
  wire       [31:0]   fixTo_1099_dout;
  wire       [15:0]   fixTo_1100_dout;
  wire       [15:0]   fixTo_1101_dout;
  wire       [15:0]   fixTo_1102_dout;
  wire       [15:0]   fixTo_1103_dout;
  wire       [31:0]   fixTo_1104_dout;
  wire       [31:0]   fixTo_1105_dout;
  wire       [15:0]   fixTo_1106_dout;
  wire       [15:0]   fixTo_1107_dout;
  wire       [15:0]   fixTo_1108_dout;
  wire       [15:0]   fixTo_1109_dout;
  wire       [31:0]   fixTo_1110_dout;
  wire       [31:0]   fixTo_1111_dout;
  wire       [15:0]   fixTo_1112_dout;
  wire       [15:0]   fixTo_1113_dout;
  wire       [15:0]   fixTo_1114_dout;
  wire       [15:0]   fixTo_1115_dout;
  wire       [31:0]   fixTo_1116_dout;
  wire       [31:0]   fixTo_1117_dout;
  wire       [15:0]   fixTo_1118_dout;
  wire       [15:0]   fixTo_1119_dout;
  wire       [15:0]   fixTo_1120_dout;
  wire       [15:0]   fixTo_1121_dout;
  wire       [31:0]   fixTo_1122_dout;
  wire       [31:0]   fixTo_1123_dout;
  wire       [15:0]   fixTo_1124_dout;
  wire       [15:0]   fixTo_1125_dout;
  wire       [15:0]   fixTo_1126_dout;
  wire       [15:0]   fixTo_1127_dout;
  wire       [31:0]   fixTo_1128_dout;
  wire       [31:0]   fixTo_1129_dout;
  wire       [15:0]   fixTo_1130_dout;
  wire       [15:0]   fixTo_1131_dout;
  wire       [15:0]   fixTo_1132_dout;
  wire       [15:0]   fixTo_1133_dout;
  wire       [31:0]   fixTo_1134_dout;
  wire       [31:0]   fixTo_1135_dout;
  wire       [15:0]   fixTo_1136_dout;
  wire       [15:0]   fixTo_1137_dout;
  wire       [15:0]   fixTo_1138_dout;
  wire       [15:0]   fixTo_1139_dout;
  wire       [31:0]   fixTo_1140_dout;
  wire       [31:0]   fixTo_1141_dout;
  wire       [15:0]   fixTo_1142_dout;
  wire       [15:0]   fixTo_1143_dout;
  wire       [15:0]   fixTo_1144_dout;
  wire       [15:0]   fixTo_1145_dout;
  wire       [31:0]   fixTo_1146_dout;
  wire       [31:0]   fixTo_1147_dout;
  wire       [15:0]   fixTo_1148_dout;
  wire       [15:0]   fixTo_1149_dout;
  wire       [15:0]   fixTo_1150_dout;
  wire       [15:0]   fixTo_1151_dout;
  wire       [31:0]   fixTo_1152_dout;
  wire       [31:0]   fixTo_1153_dout;
  wire       [15:0]   fixTo_1154_dout;
  wire       [15:0]   fixTo_1155_dout;
  wire       [15:0]   fixTo_1156_dout;
  wire       [15:0]   fixTo_1157_dout;
  wire       [31:0]   fixTo_1158_dout;
  wire       [31:0]   fixTo_1159_dout;
  wire       [15:0]   fixTo_1160_dout;
  wire       [15:0]   fixTo_1161_dout;
  wire       [15:0]   fixTo_1162_dout;
  wire       [15:0]   fixTo_1163_dout;
  wire       [31:0]   fixTo_1164_dout;
  wire       [31:0]   fixTo_1165_dout;
  wire       [15:0]   fixTo_1166_dout;
  wire       [15:0]   fixTo_1167_dout;
  wire       [15:0]   fixTo_1168_dout;
  wire       [15:0]   fixTo_1169_dout;
  wire       [31:0]   fixTo_1170_dout;
  wire       [31:0]   fixTo_1171_dout;
  wire       [15:0]   fixTo_1172_dout;
  wire       [15:0]   fixTo_1173_dout;
  wire       [15:0]   fixTo_1174_dout;
  wire       [15:0]   fixTo_1175_dout;
  wire       [31:0]   fixTo_1176_dout;
  wire       [31:0]   fixTo_1177_dout;
  wire       [15:0]   fixTo_1178_dout;
  wire       [15:0]   fixTo_1179_dout;
  wire       [15:0]   fixTo_1180_dout;
  wire       [15:0]   fixTo_1181_dout;
  wire       [31:0]   fixTo_1182_dout;
  wire       [31:0]   fixTo_1183_dout;
  wire       [15:0]   fixTo_1184_dout;
  wire       [15:0]   fixTo_1185_dout;
  wire       [15:0]   fixTo_1186_dout;
  wire       [15:0]   fixTo_1187_dout;
  wire       [31:0]   fixTo_1188_dout;
  wire       [31:0]   fixTo_1189_dout;
  wire       [15:0]   fixTo_1190_dout;
  wire       [15:0]   fixTo_1191_dout;
  wire       [15:0]   fixTo_1192_dout;
  wire       [15:0]   fixTo_1193_dout;
  wire       [31:0]   fixTo_1194_dout;
  wire       [31:0]   fixTo_1195_dout;
  wire       [15:0]   fixTo_1196_dout;
  wire       [15:0]   fixTo_1197_dout;
  wire       [15:0]   fixTo_1198_dout;
  wire       [15:0]   fixTo_1199_dout;
  wire       [31:0]   fixTo_1200_dout;
  wire       [31:0]   fixTo_1201_dout;
  wire       [15:0]   fixTo_1202_dout;
  wire       [15:0]   fixTo_1203_dout;
  wire       [15:0]   fixTo_1204_dout;
  wire       [15:0]   fixTo_1205_dout;
  wire       [31:0]   fixTo_1206_dout;
  wire       [31:0]   fixTo_1207_dout;
  wire       [15:0]   fixTo_1208_dout;
  wire       [15:0]   fixTo_1209_dout;
  wire       [15:0]   fixTo_1210_dout;
  wire       [15:0]   fixTo_1211_dout;
  wire       [31:0]   fixTo_1212_dout;
  wire       [31:0]   fixTo_1213_dout;
  wire       [15:0]   fixTo_1214_dout;
  wire       [15:0]   fixTo_1215_dout;
  wire       [15:0]   fixTo_1216_dout;
  wire       [15:0]   fixTo_1217_dout;
  wire       [31:0]   fixTo_1218_dout;
  wire       [31:0]   fixTo_1219_dout;
  wire       [15:0]   fixTo_1220_dout;
  wire       [15:0]   fixTo_1221_dout;
  wire       [15:0]   fixTo_1222_dout;
  wire       [15:0]   fixTo_1223_dout;
  wire       [31:0]   fixTo_1224_dout;
  wire       [31:0]   fixTo_1225_dout;
  wire       [15:0]   fixTo_1226_dout;
  wire       [15:0]   fixTo_1227_dout;
  wire       [15:0]   fixTo_1228_dout;
  wire       [15:0]   fixTo_1229_dout;
  wire       [31:0]   fixTo_1230_dout;
  wire       [31:0]   fixTo_1231_dout;
  wire       [15:0]   fixTo_1232_dout;
  wire       [15:0]   fixTo_1233_dout;
  wire       [15:0]   fixTo_1234_dout;
  wire       [15:0]   fixTo_1235_dout;
  wire       [31:0]   fixTo_1236_dout;
  wire       [31:0]   fixTo_1237_dout;
  wire       [15:0]   fixTo_1238_dout;
  wire       [15:0]   fixTo_1239_dout;
  wire       [15:0]   fixTo_1240_dout;
  wire       [15:0]   fixTo_1241_dout;
  wire       [31:0]   fixTo_1242_dout;
  wire       [31:0]   fixTo_1243_dout;
  wire       [15:0]   fixTo_1244_dout;
  wire       [15:0]   fixTo_1245_dout;
  wire       [15:0]   fixTo_1246_dout;
  wire       [15:0]   fixTo_1247_dout;
  wire       [31:0]   fixTo_1248_dout;
  wire       [31:0]   fixTo_1249_dout;
  wire       [15:0]   fixTo_1250_dout;
  wire       [15:0]   fixTo_1251_dout;
  wire       [15:0]   fixTo_1252_dout;
  wire       [15:0]   fixTo_1253_dout;
  wire       [31:0]   fixTo_1254_dout;
  wire       [31:0]   fixTo_1255_dout;
  wire       [15:0]   fixTo_1256_dout;
  wire       [15:0]   fixTo_1257_dout;
  wire       [15:0]   fixTo_1258_dout;
  wire       [15:0]   fixTo_1259_dout;
  wire       [31:0]   fixTo_1260_dout;
  wire       [31:0]   fixTo_1261_dout;
  wire       [15:0]   fixTo_1262_dout;
  wire       [15:0]   fixTo_1263_dout;
  wire       [15:0]   fixTo_1264_dout;
  wire       [15:0]   fixTo_1265_dout;
  wire       [31:0]   fixTo_1266_dout;
  wire       [31:0]   fixTo_1267_dout;
  wire       [15:0]   fixTo_1268_dout;
  wire       [15:0]   fixTo_1269_dout;
  wire       [15:0]   fixTo_1270_dout;
  wire       [15:0]   fixTo_1271_dout;
  wire       [31:0]   fixTo_1272_dout;
  wire       [31:0]   fixTo_1273_dout;
  wire       [15:0]   fixTo_1274_dout;
  wire       [15:0]   fixTo_1275_dout;
  wire       [15:0]   fixTo_1276_dout;
  wire       [15:0]   fixTo_1277_dout;
  wire       [31:0]   fixTo_1278_dout;
  wire       [31:0]   fixTo_1279_dout;
  wire       [15:0]   fixTo_1280_dout;
  wire       [15:0]   fixTo_1281_dout;
  wire       [15:0]   fixTo_1282_dout;
  wire       [15:0]   fixTo_1283_dout;
  wire       [31:0]   fixTo_1284_dout;
  wire       [31:0]   fixTo_1285_dout;
  wire       [15:0]   fixTo_1286_dout;
  wire       [15:0]   fixTo_1287_dout;
  wire       [15:0]   fixTo_1288_dout;
  wire       [15:0]   fixTo_1289_dout;
  wire       [31:0]   fixTo_1290_dout;
  wire       [31:0]   fixTo_1291_dout;
  wire       [15:0]   fixTo_1292_dout;
  wire       [15:0]   fixTo_1293_dout;
  wire       [15:0]   fixTo_1294_dout;
  wire       [15:0]   fixTo_1295_dout;
  wire       [31:0]   fixTo_1296_dout;
  wire       [31:0]   fixTo_1297_dout;
  wire       [15:0]   fixTo_1298_dout;
  wire       [15:0]   fixTo_1299_dout;
  wire       [15:0]   fixTo_1300_dout;
  wire       [15:0]   fixTo_1301_dout;
  wire       [31:0]   fixTo_1302_dout;
  wire       [31:0]   fixTo_1303_dout;
  wire       [15:0]   fixTo_1304_dout;
  wire       [15:0]   fixTo_1305_dout;
  wire       [15:0]   fixTo_1306_dout;
  wire       [15:0]   fixTo_1307_dout;
  wire       [31:0]   fixTo_1308_dout;
  wire       [31:0]   fixTo_1309_dout;
  wire       [15:0]   fixTo_1310_dout;
  wire       [15:0]   fixTo_1311_dout;
  wire       [15:0]   fixTo_1312_dout;
  wire       [15:0]   fixTo_1313_dout;
  wire       [31:0]   fixTo_1314_dout;
  wire       [31:0]   fixTo_1315_dout;
  wire       [15:0]   fixTo_1316_dout;
  wire       [15:0]   fixTo_1317_dout;
  wire       [15:0]   fixTo_1318_dout;
  wire       [15:0]   fixTo_1319_dout;
  wire       [31:0]   fixTo_1320_dout;
  wire       [31:0]   fixTo_1321_dout;
  wire       [15:0]   fixTo_1322_dout;
  wire       [15:0]   fixTo_1323_dout;
  wire       [15:0]   fixTo_1324_dout;
  wire       [15:0]   fixTo_1325_dout;
  wire       [31:0]   fixTo_1326_dout;
  wire       [31:0]   fixTo_1327_dout;
  wire       [15:0]   fixTo_1328_dout;
  wire       [15:0]   fixTo_1329_dout;
  wire       [15:0]   fixTo_1330_dout;
  wire       [15:0]   fixTo_1331_dout;
  wire       [31:0]   fixTo_1332_dout;
  wire       [31:0]   fixTo_1333_dout;
  wire       [15:0]   fixTo_1334_dout;
  wire       [15:0]   fixTo_1335_dout;
  wire       [15:0]   fixTo_1336_dout;
  wire       [15:0]   fixTo_1337_dout;
  wire       [31:0]   fixTo_1338_dout;
  wire       [31:0]   fixTo_1339_dout;
  wire       [15:0]   fixTo_1340_dout;
  wire       [15:0]   fixTo_1341_dout;
  wire       [15:0]   fixTo_1342_dout;
  wire       [15:0]   fixTo_1343_dout;
  wire       [31:0]   fixTo_1344_dout;
  wire       [31:0]   fixTo_1345_dout;
  wire       [15:0]   fixTo_1346_dout;
  wire       [15:0]   fixTo_1347_dout;
  wire       [15:0]   fixTo_1348_dout;
  wire       [15:0]   fixTo_1349_dout;
  wire       [31:0]   fixTo_1350_dout;
  wire       [31:0]   fixTo_1351_dout;
  wire       [15:0]   fixTo_1352_dout;
  wire       [15:0]   fixTo_1353_dout;
  wire       [15:0]   fixTo_1354_dout;
  wire       [15:0]   fixTo_1355_dout;
  wire       [31:0]   fixTo_1356_dout;
  wire       [31:0]   fixTo_1357_dout;
  wire       [15:0]   fixTo_1358_dout;
  wire       [15:0]   fixTo_1359_dout;
  wire       [15:0]   fixTo_1360_dout;
  wire       [15:0]   fixTo_1361_dout;
  wire       [31:0]   fixTo_1362_dout;
  wire       [31:0]   fixTo_1363_dout;
  wire       [15:0]   fixTo_1364_dout;
  wire       [15:0]   fixTo_1365_dout;
  wire       [15:0]   fixTo_1366_dout;
  wire       [15:0]   fixTo_1367_dout;
  wire       [31:0]   fixTo_1368_dout;
  wire       [31:0]   fixTo_1369_dout;
  wire       [15:0]   fixTo_1370_dout;
  wire       [15:0]   fixTo_1371_dout;
  wire       [15:0]   fixTo_1372_dout;
  wire       [15:0]   fixTo_1373_dout;
  wire       [31:0]   fixTo_1374_dout;
  wire       [31:0]   fixTo_1375_dout;
  wire       [15:0]   fixTo_1376_dout;
  wire       [15:0]   fixTo_1377_dout;
  wire       [15:0]   fixTo_1378_dout;
  wire       [15:0]   fixTo_1379_dout;
  wire       [31:0]   fixTo_1380_dout;
  wire       [31:0]   fixTo_1381_dout;
  wire       [15:0]   fixTo_1382_dout;
  wire       [15:0]   fixTo_1383_dout;
  wire       [15:0]   fixTo_1384_dout;
  wire       [15:0]   fixTo_1385_dout;
  wire       [31:0]   fixTo_1386_dout;
  wire       [31:0]   fixTo_1387_dout;
  wire       [15:0]   fixTo_1388_dout;
  wire       [15:0]   fixTo_1389_dout;
  wire       [15:0]   fixTo_1390_dout;
  wire       [15:0]   fixTo_1391_dout;
  wire       [31:0]   fixTo_1392_dout;
  wire       [31:0]   fixTo_1393_dout;
  wire       [15:0]   fixTo_1394_dout;
  wire       [15:0]   fixTo_1395_dout;
  wire       [15:0]   fixTo_1396_dout;
  wire       [15:0]   fixTo_1397_dout;
  wire       [31:0]   fixTo_1398_dout;
  wire       [31:0]   fixTo_1399_dout;
  wire       [15:0]   fixTo_1400_dout;
  wire       [15:0]   fixTo_1401_dout;
  wire       [15:0]   fixTo_1402_dout;
  wire       [15:0]   fixTo_1403_dout;
  wire       [31:0]   fixTo_1404_dout;
  wire       [31:0]   fixTo_1405_dout;
  wire       [15:0]   fixTo_1406_dout;
  wire       [15:0]   fixTo_1407_dout;
  wire       [15:0]   fixTo_1408_dout;
  wire       [15:0]   fixTo_1409_dout;
  wire       [31:0]   fixTo_1410_dout;
  wire       [31:0]   fixTo_1411_dout;
  wire       [15:0]   fixTo_1412_dout;
  wire       [15:0]   fixTo_1413_dout;
  wire       [15:0]   fixTo_1414_dout;
  wire       [15:0]   fixTo_1415_dout;
  wire       [31:0]   fixTo_1416_dout;
  wire       [31:0]   fixTo_1417_dout;
  wire       [15:0]   fixTo_1418_dout;
  wire       [15:0]   fixTo_1419_dout;
  wire       [15:0]   fixTo_1420_dout;
  wire       [15:0]   fixTo_1421_dout;
  wire       [31:0]   fixTo_1422_dout;
  wire       [31:0]   fixTo_1423_dout;
  wire       [15:0]   fixTo_1424_dout;
  wire       [15:0]   fixTo_1425_dout;
  wire       [15:0]   fixTo_1426_dout;
  wire       [15:0]   fixTo_1427_dout;
  wire       [31:0]   fixTo_1428_dout;
  wire       [31:0]   fixTo_1429_dout;
  wire       [15:0]   fixTo_1430_dout;
  wire       [15:0]   fixTo_1431_dout;
  wire       [15:0]   fixTo_1432_dout;
  wire       [15:0]   fixTo_1433_dout;
  wire       [31:0]   fixTo_1434_dout;
  wire       [31:0]   fixTo_1435_dout;
  wire       [15:0]   fixTo_1436_dout;
  wire       [15:0]   fixTo_1437_dout;
  wire       [15:0]   fixTo_1438_dout;
  wire       [15:0]   fixTo_1439_dout;
  wire       [31:0]   fixTo_1440_dout;
  wire       [31:0]   fixTo_1441_dout;
  wire       [15:0]   fixTo_1442_dout;
  wire       [15:0]   fixTo_1443_dout;
  wire       [15:0]   fixTo_1444_dout;
  wire       [15:0]   fixTo_1445_dout;
  wire       [31:0]   fixTo_1446_dout;
  wire       [31:0]   fixTo_1447_dout;
  wire       [15:0]   fixTo_1448_dout;
  wire       [15:0]   fixTo_1449_dout;
  wire       [15:0]   fixTo_1450_dout;
  wire       [15:0]   fixTo_1451_dout;
  wire       [31:0]   fixTo_1452_dout;
  wire       [31:0]   fixTo_1453_dout;
  wire       [15:0]   fixTo_1454_dout;
  wire       [15:0]   fixTo_1455_dout;
  wire       [15:0]   fixTo_1456_dout;
  wire       [15:0]   fixTo_1457_dout;
  wire       [31:0]   fixTo_1458_dout;
  wire       [31:0]   fixTo_1459_dout;
  wire       [15:0]   fixTo_1460_dout;
  wire       [15:0]   fixTo_1461_dout;
  wire       [15:0]   fixTo_1462_dout;
  wire       [15:0]   fixTo_1463_dout;
  wire       [31:0]   fixTo_1464_dout;
  wire       [31:0]   fixTo_1465_dout;
  wire       [15:0]   fixTo_1466_dout;
  wire       [15:0]   fixTo_1467_dout;
  wire       [15:0]   fixTo_1468_dout;
  wire       [15:0]   fixTo_1469_dout;
  wire       [31:0]   fixTo_1470_dout;
  wire       [31:0]   fixTo_1471_dout;
  wire       [15:0]   fixTo_1472_dout;
  wire       [15:0]   fixTo_1473_dout;
  wire       [15:0]   fixTo_1474_dout;
  wire       [15:0]   fixTo_1475_dout;
  wire       [31:0]   fixTo_1476_dout;
  wire       [31:0]   fixTo_1477_dout;
  wire       [15:0]   fixTo_1478_dout;
  wire       [15:0]   fixTo_1479_dout;
  wire       [15:0]   fixTo_1480_dout;
  wire       [15:0]   fixTo_1481_dout;
  wire       [31:0]   fixTo_1482_dout;
  wire       [31:0]   fixTo_1483_dout;
  wire       [15:0]   fixTo_1484_dout;
  wire       [15:0]   fixTo_1485_dout;
  wire       [15:0]   fixTo_1486_dout;
  wire       [15:0]   fixTo_1487_dout;
  wire       [31:0]   fixTo_1488_dout;
  wire       [31:0]   fixTo_1489_dout;
  wire       [15:0]   fixTo_1490_dout;
  wire       [15:0]   fixTo_1491_dout;
  wire       [15:0]   fixTo_1492_dout;
  wire       [15:0]   fixTo_1493_dout;
  wire       [31:0]   fixTo_1494_dout;
  wire       [31:0]   fixTo_1495_dout;
  wire       [15:0]   fixTo_1496_dout;
  wire       [15:0]   fixTo_1497_dout;
  wire       [15:0]   fixTo_1498_dout;
  wire       [15:0]   fixTo_1499_dout;
  wire       [31:0]   fixTo_1500_dout;
  wire       [31:0]   fixTo_1501_dout;
  wire       [15:0]   fixTo_1502_dout;
  wire       [15:0]   fixTo_1503_dout;
  wire       [15:0]   fixTo_1504_dout;
  wire       [15:0]   fixTo_1505_dout;
  wire       [31:0]   fixTo_1506_dout;
  wire       [31:0]   fixTo_1507_dout;
  wire       [15:0]   fixTo_1508_dout;
  wire       [15:0]   fixTo_1509_dout;
  wire       [15:0]   fixTo_1510_dout;
  wire       [15:0]   fixTo_1511_dout;
  wire       [31:0]   fixTo_1512_dout;
  wire       [31:0]   fixTo_1513_dout;
  wire       [15:0]   fixTo_1514_dout;
  wire       [15:0]   fixTo_1515_dout;
  wire       [15:0]   fixTo_1516_dout;
  wire       [15:0]   fixTo_1517_dout;
  wire       [31:0]   fixTo_1518_dout;
  wire       [31:0]   fixTo_1519_dout;
  wire       [15:0]   fixTo_1520_dout;
  wire       [15:0]   fixTo_1521_dout;
  wire       [15:0]   fixTo_1522_dout;
  wire       [15:0]   fixTo_1523_dout;
  wire       [31:0]   fixTo_1524_dout;
  wire       [31:0]   fixTo_1525_dout;
  wire       [15:0]   fixTo_1526_dout;
  wire       [15:0]   fixTo_1527_dout;
  wire       [15:0]   fixTo_1528_dout;
  wire       [15:0]   fixTo_1529_dout;
  wire       [31:0]   fixTo_1530_dout;
  wire       [31:0]   fixTo_1531_dout;
  wire       [15:0]   fixTo_1532_dout;
  wire       [15:0]   fixTo_1533_dout;
  wire       [15:0]   fixTo_1534_dout;
  wire       [15:0]   fixTo_1535_dout;
  wire       [31:0]   fixTo_1536_dout;
  wire       [31:0]   fixTo_1537_dout;
  wire       [15:0]   fixTo_1538_dout;
  wire       [15:0]   fixTo_1539_dout;
  wire       [15:0]   fixTo_1540_dout;
  wire       [15:0]   fixTo_1541_dout;
  wire       [31:0]   fixTo_1542_dout;
  wire       [31:0]   fixTo_1543_dout;
  wire       [15:0]   fixTo_1544_dout;
  wire       [15:0]   fixTo_1545_dout;
  wire       [15:0]   fixTo_1546_dout;
  wire       [15:0]   fixTo_1547_dout;
  wire       [31:0]   fixTo_1548_dout;
  wire       [31:0]   fixTo_1549_dout;
  wire       [15:0]   fixTo_1550_dout;
  wire       [15:0]   fixTo_1551_dout;
  wire       [15:0]   fixTo_1552_dout;
  wire       [15:0]   fixTo_1553_dout;
  wire       [31:0]   fixTo_1554_dout;
  wire       [31:0]   fixTo_1555_dout;
  wire       [15:0]   fixTo_1556_dout;
  wire       [15:0]   fixTo_1557_dout;
  wire       [15:0]   fixTo_1558_dout;
  wire       [15:0]   fixTo_1559_dout;
  wire       [31:0]   fixTo_1560_dout;
  wire       [31:0]   fixTo_1561_dout;
  wire       [15:0]   fixTo_1562_dout;
  wire       [15:0]   fixTo_1563_dout;
  wire       [15:0]   fixTo_1564_dout;
  wire       [15:0]   fixTo_1565_dout;
  wire       [31:0]   fixTo_1566_dout;
  wire       [31:0]   fixTo_1567_dout;
  wire       [15:0]   fixTo_1568_dout;
  wire       [15:0]   fixTo_1569_dout;
  wire       [15:0]   fixTo_1570_dout;
  wire       [15:0]   fixTo_1571_dout;
  wire       [31:0]   fixTo_1572_dout;
  wire       [31:0]   fixTo_1573_dout;
  wire       [15:0]   fixTo_1574_dout;
  wire       [15:0]   fixTo_1575_dout;
  wire       [15:0]   fixTo_1576_dout;
  wire       [15:0]   fixTo_1577_dout;
  wire       [31:0]   fixTo_1578_dout;
  wire       [31:0]   fixTo_1579_dout;
  wire       [15:0]   fixTo_1580_dout;
  wire       [15:0]   fixTo_1581_dout;
  wire       [15:0]   fixTo_1582_dout;
  wire       [15:0]   fixTo_1583_dout;
  wire       [31:0]   fixTo_1584_dout;
  wire       [31:0]   fixTo_1585_dout;
  wire       [15:0]   fixTo_1586_dout;
  wire       [15:0]   fixTo_1587_dout;
  wire       [15:0]   fixTo_1588_dout;
  wire       [15:0]   fixTo_1589_dout;
  wire       [31:0]   fixTo_1590_dout;
  wire       [31:0]   fixTo_1591_dout;
  wire       [15:0]   fixTo_1592_dout;
  wire       [15:0]   fixTo_1593_dout;
  wire       [15:0]   fixTo_1594_dout;
  wire       [15:0]   fixTo_1595_dout;
  wire       [31:0]   fixTo_1596_dout;
  wire       [31:0]   fixTo_1597_dout;
  wire       [15:0]   fixTo_1598_dout;
  wire       [15:0]   fixTo_1599_dout;
  wire       [15:0]   fixTo_1600_dout;
  wire       [15:0]   fixTo_1601_dout;
  wire       [31:0]   fixTo_1602_dout;
  wire       [31:0]   fixTo_1603_dout;
  wire       [15:0]   fixTo_1604_dout;
  wire       [15:0]   fixTo_1605_dout;
  wire       [15:0]   fixTo_1606_dout;
  wire       [15:0]   fixTo_1607_dout;
  wire       [31:0]   fixTo_1608_dout;
  wire       [31:0]   fixTo_1609_dout;
  wire       [15:0]   fixTo_1610_dout;
  wire       [15:0]   fixTo_1611_dout;
  wire       [15:0]   fixTo_1612_dout;
  wire       [15:0]   fixTo_1613_dout;
  wire       [31:0]   fixTo_1614_dout;
  wire       [31:0]   fixTo_1615_dout;
  wire       [15:0]   fixTo_1616_dout;
  wire       [15:0]   fixTo_1617_dout;
  wire       [15:0]   fixTo_1618_dout;
  wire       [15:0]   fixTo_1619_dout;
  wire       [31:0]   fixTo_1620_dout;
  wire       [31:0]   fixTo_1621_dout;
  wire       [15:0]   fixTo_1622_dout;
  wire       [15:0]   fixTo_1623_dout;
  wire       [15:0]   fixTo_1624_dout;
  wire       [15:0]   fixTo_1625_dout;
  wire       [31:0]   fixTo_1626_dout;
  wire       [31:0]   fixTo_1627_dout;
  wire       [15:0]   fixTo_1628_dout;
  wire       [15:0]   fixTo_1629_dout;
  wire       [15:0]   fixTo_1630_dout;
  wire       [15:0]   fixTo_1631_dout;
  wire       [31:0]   fixTo_1632_dout;
  wire       [31:0]   fixTo_1633_dout;
  wire       [15:0]   fixTo_1634_dout;
  wire       [15:0]   fixTo_1635_dout;
  wire       [15:0]   fixTo_1636_dout;
  wire       [15:0]   fixTo_1637_dout;
  wire       [31:0]   fixTo_1638_dout;
  wire       [31:0]   fixTo_1639_dout;
  wire       [15:0]   fixTo_1640_dout;
  wire       [15:0]   fixTo_1641_dout;
  wire       [15:0]   fixTo_1642_dout;
  wire       [15:0]   fixTo_1643_dout;
  wire       [31:0]   fixTo_1644_dout;
  wire       [31:0]   fixTo_1645_dout;
  wire       [15:0]   fixTo_1646_dout;
  wire       [15:0]   fixTo_1647_dout;
  wire       [15:0]   fixTo_1648_dout;
  wire       [15:0]   fixTo_1649_dout;
  wire       [31:0]   fixTo_1650_dout;
  wire       [31:0]   fixTo_1651_dout;
  wire       [15:0]   fixTo_1652_dout;
  wire       [15:0]   fixTo_1653_dout;
  wire       [15:0]   fixTo_1654_dout;
  wire       [15:0]   fixTo_1655_dout;
  wire       [31:0]   fixTo_1656_dout;
  wire       [31:0]   fixTo_1657_dout;
  wire       [15:0]   fixTo_1658_dout;
  wire       [15:0]   fixTo_1659_dout;
  wire       [15:0]   fixTo_1660_dout;
  wire       [15:0]   fixTo_1661_dout;
  wire       [31:0]   fixTo_1662_dout;
  wire       [31:0]   fixTo_1663_dout;
  wire       [15:0]   fixTo_1664_dout;
  wire       [15:0]   fixTo_1665_dout;
  wire       [15:0]   fixTo_1666_dout;
  wire       [15:0]   fixTo_1667_dout;
  wire       [31:0]   fixTo_1668_dout;
  wire       [31:0]   fixTo_1669_dout;
  wire       [15:0]   fixTo_1670_dout;
  wire       [15:0]   fixTo_1671_dout;
  wire       [15:0]   fixTo_1672_dout;
  wire       [15:0]   fixTo_1673_dout;
  wire       [31:0]   fixTo_1674_dout;
  wire       [31:0]   fixTo_1675_dout;
  wire       [15:0]   fixTo_1676_dout;
  wire       [15:0]   fixTo_1677_dout;
  wire       [15:0]   fixTo_1678_dout;
  wire       [15:0]   fixTo_1679_dout;
  wire       [31:0]   fixTo_1680_dout;
  wire       [31:0]   fixTo_1681_dout;
  wire       [15:0]   fixTo_1682_dout;
  wire       [15:0]   fixTo_1683_dout;
  wire       [15:0]   fixTo_1684_dout;
  wire       [15:0]   fixTo_1685_dout;
  wire       [31:0]   fixTo_1686_dout;
  wire       [31:0]   fixTo_1687_dout;
  wire       [15:0]   fixTo_1688_dout;
  wire       [15:0]   fixTo_1689_dout;
  wire       [15:0]   fixTo_1690_dout;
  wire       [15:0]   fixTo_1691_dout;
  wire       [31:0]   fixTo_1692_dout;
  wire       [31:0]   fixTo_1693_dout;
  wire       [15:0]   fixTo_1694_dout;
  wire       [15:0]   fixTo_1695_dout;
  wire       [15:0]   fixTo_1696_dout;
  wire       [15:0]   fixTo_1697_dout;
  wire       [31:0]   fixTo_1698_dout;
  wire       [31:0]   fixTo_1699_dout;
  wire       [15:0]   fixTo_1700_dout;
  wire       [15:0]   fixTo_1701_dout;
  wire       [15:0]   fixTo_1702_dout;
  wire       [15:0]   fixTo_1703_dout;
  wire       [31:0]   fixTo_1704_dout;
  wire       [31:0]   fixTo_1705_dout;
  wire       [15:0]   fixTo_1706_dout;
  wire       [15:0]   fixTo_1707_dout;
  wire       [15:0]   fixTo_1708_dout;
  wire       [15:0]   fixTo_1709_dout;
  wire       [31:0]   fixTo_1710_dout;
  wire       [31:0]   fixTo_1711_dout;
  wire       [15:0]   fixTo_1712_dout;
  wire       [15:0]   fixTo_1713_dout;
  wire       [15:0]   fixTo_1714_dout;
  wire       [15:0]   fixTo_1715_dout;
  wire       [31:0]   fixTo_1716_dout;
  wire       [31:0]   fixTo_1717_dout;
  wire       [15:0]   fixTo_1718_dout;
  wire       [15:0]   fixTo_1719_dout;
  wire       [15:0]   fixTo_1720_dout;
  wire       [15:0]   fixTo_1721_dout;
  wire       [31:0]   fixTo_1722_dout;
  wire       [31:0]   fixTo_1723_dout;
  wire       [15:0]   fixTo_1724_dout;
  wire       [15:0]   fixTo_1725_dout;
  wire       [15:0]   fixTo_1726_dout;
  wire       [15:0]   fixTo_1727_dout;
  wire       [31:0]   fixTo_1728_dout;
  wire       [31:0]   fixTo_1729_dout;
  wire       [15:0]   fixTo_1730_dout;
  wire       [15:0]   fixTo_1731_dout;
  wire       [15:0]   fixTo_1732_dout;
  wire       [15:0]   fixTo_1733_dout;
  wire       [31:0]   fixTo_1734_dout;
  wire       [31:0]   fixTo_1735_dout;
  wire       [15:0]   fixTo_1736_dout;
  wire       [15:0]   fixTo_1737_dout;
  wire       [15:0]   fixTo_1738_dout;
  wire       [15:0]   fixTo_1739_dout;
  wire       [31:0]   fixTo_1740_dout;
  wire       [31:0]   fixTo_1741_dout;
  wire       [15:0]   fixTo_1742_dout;
  wire       [15:0]   fixTo_1743_dout;
  wire       [15:0]   fixTo_1744_dout;
  wire       [15:0]   fixTo_1745_dout;
  wire       [31:0]   fixTo_1746_dout;
  wire       [31:0]   fixTo_1747_dout;
  wire       [15:0]   fixTo_1748_dout;
  wire       [15:0]   fixTo_1749_dout;
  wire       [15:0]   fixTo_1750_dout;
  wire       [15:0]   fixTo_1751_dout;
  wire       [31:0]   fixTo_1752_dout;
  wire       [31:0]   fixTo_1753_dout;
  wire       [15:0]   fixTo_1754_dout;
  wire       [15:0]   fixTo_1755_dout;
  wire       [15:0]   fixTo_1756_dout;
  wire       [15:0]   fixTo_1757_dout;
  wire       [31:0]   fixTo_1758_dout;
  wire       [31:0]   fixTo_1759_dout;
  wire       [15:0]   fixTo_1760_dout;
  wire       [15:0]   fixTo_1761_dout;
  wire       [15:0]   fixTo_1762_dout;
  wire       [15:0]   fixTo_1763_dout;
  wire       [31:0]   fixTo_1764_dout;
  wire       [31:0]   fixTo_1765_dout;
  wire       [15:0]   fixTo_1766_dout;
  wire       [15:0]   fixTo_1767_dout;
  wire       [15:0]   fixTo_1768_dout;
  wire       [15:0]   fixTo_1769_dout;
  wire       [31:0]   fixTo_1770_dout;
  wire       [31:0]   fixTo_1771_dout;
  wire       [15:0]   fixTo_1772_dout;
  wire       [15:0]   fixTo_1773_dout;
  wire       [15:0]   fixTo_1774_dout;
  wire       [15:0]   fixTo_1775_dout;
  wire       [31:0]   fixTo_1776_dout;
  wire       [31:0]   fixTo_1777_dout;
  wire       [15:0]   fixTo_1778_dout;
  wire       [15:0]   fixTo_1779_dout;
  wire       [15:0]   fixTo_1780_dout;
  wire       [15:0]   fixTo_1781_dout;
  wire       [31:0]   fixTo_1782_dout;
  wire       [31:0]   fixTo_1783_dout;
  wire       [15:0]   fixTo_1784_dout;
  wire       [15:0]   fixTo_1785_dout;
  wire       [15:0]   fixTo_1786_dout;
  wire       [15:0]   fixTo_1787_dout;
  wire       [31:0]   fixTo_1788_dout;
  wire       [31:0]   fixTo_1789_dout;
  wire       [15:0]   fixTo_1790_dout;
  wire       [15:0]   fixTo_1791_dout;
  wire       [15:0]   fixTo_1792_dout;
  wire       [15:0]   fixTo_1793_dout;
  wire       [31:0]   fixTo_1794_dout;
  wire       [31:0]   fixTo_1795_dout;
  wire       [15:0]   fixTo_1796_dout;
  wire       [15:0]   fixTo_1797_dout;
  wire       [15:0]   fixTo_1798_dout;
  wire       [15:0]   fixTo_1799_dout;
  wire       [31:0]   fixTo_1800_dout;
  wire       [31:0]   fixTo_1801_dout;
  wire       [15:0]   fixTo_1802_dout;
  wire       [15:0]   fixTo_1803_dout;
  wire       [15:0]   fixTo_1804_dout;
  wire       [15:0]   fixTo_1805_dout;
  wire       [31:0]   fixTo_1806_dout;
  wire       [31:0]   fixTo_1807_dout;
  wire       [15:0]   fixTo_1808_dout;
  wire       [15:0]   fixTo_1809_dout;
  wire       [15:0]   fixTo_1810_dout;
  wire       [15:0]   fixTo_1811_dout;
  wire       [31:0]   fixTo_1812_dout;
  wire       [31:0]   fixTo_1813_dout;
  wire       [15:0]   fixTo_1814_dout;
  wire       [15:0]   fixTo_1815_dout;
  wire       [15:0]   fixTo_1816_dout;
  wire       [15:0]   fixTo_1817_dout;
  wire       [31:0]   fixTo_1818_dout;
  wire       [31:0]   fixTo_1819_dout;
  wire       [15:0]   fixTo_1820_dout;
  wire       [15:0]   fixTo_1821_dout;
  wire       [15:0]   fixTo_1822_dout;
  wire       [15:0]   fixTo_1823_dout;
  wire       [31:0]   fixTo_1824_dout;
  wire       [31:0]   fixTo_1825_dout;
  wire       [15:0]   fixTo_1826_dout;
  wire       [15:0]   fixTo_1827_dout;
  wire       [15:0]   fixTo_1828_dout;
  wire       [15:0]   fixTo_1829_dout;
  wire       [31:0]   fixTo_1830_dout;
  wire       [31:0]   fixTo_1831_dout;
  wire       [15:0]   fixTo_1832_dout;
  wire       [15:0]   fixTo_1833_dout;
  wire       [15:0]   fixTo_1834_dout;
  wire       [15:0]   fixTo_1835_dout;
  wire       [31:0]   fixTo_1836_dout;
  wire       [31:0]   fixTo_1837_dout;
  wire       [15:0]   fixTo_1838_dout;
  wire       [15:0]   fixTo_1839_dout;
  wire       [15:0]   fixTo_1840_dout;
  wire       [15:0]   fixTo_1841_dout;
  wire       [31:0]   fixTo_1842_dout;
  wire       [31:0]   fixTo_1843_dout;
  wire       [15:0]   fixTo_1844_dout;
  wire       [15:0]   fixTo_1845_dout;
  wire       [15:0]   fixTo_1846_dout;
  wire       [15:0]   fixTo_1847_dout;
  wire       [31:0]   fixTo_1848_dout;
  wire       [31:0]   fixTo_1849_dout;
  wire       [15:0]   fixTo_1850_dout;
  wire       [15:0]   fixTo_1851_dout;
  wire       [15:0]   fixTo_1852_dout;
  wire       [15:0]   fixTo_1853_dout;
  wire       [31:0]   fixTo_1854_dout;
  wire       [31:0]   fixTo_1855_dout;
  wire       [15:0]   fixTo_1856_dout;
  wire       [15:0]   fixTo_1857_dout;
  wire       [15:0]   fixTo_1858_dout;
  wire       [15:0]   fixTo_1859_dout;
  wire       [31:0]   fixTo_1860_dout;
  wire       [31:0]   fixTo_1861_dout;
  wire       [15:0]   fixTo_1862_dout;
  wire       [15:0]   fixTo_1863_dout;
  wire       [15:0]   fixTo_1864_dout;
  wire       [15:0]   fixTo_1865_dout;
  wire       [31:0]   fixTo_1866_dout;
  wire       [31:0]   fixTo_1867_dout;
  wire       [15:0]   fixTo_1868_dout;
  wire       [15:0]   fixTo_1869_dout;
  wire       [15:0]   fixTo_1870_dout;
  wire       [15:0]   fixTo_1871_dout;
  wire       [31:0]   fixTo_1872_dout;
  wire       [31:0]   fixTo_1873_dout;
  wire       [15:0]   fixTo_1874_dout;
  wire       [15:0]   fixTo_1875_dout;
  wire       [15:0]   fixTo_1876_dout;
  wire       [15:0]   fixTo_1877_dout;
  wire       [31:0]   fixTo_1878_dout;
  wire       [31:0]   fixTo_1879_dout;
  wire       [15:0]   fixTo_1880_dout;
  wire       [15:0]   fixTo_1881_dout;
  wire       [15:0]   fixTo_1882_dout;
  wire       [15:0]   fixTo_1883_dout;
  wire       [31:0]   fixTo_1884_dout;
  wire       [31:0]   fixTo_1885_dout;
  wire       [15:0]   fixTo_1886_dout;
  wire       [15:0]   fixTo_1887_dout;
  wire       [15:0]   fixTo_1888_dout;
  wire       [15:0]   fixTo_1889_dout;
  wire       [31:0]   fixTo_1890_dout;
  wire       [31:0]   fixTo_1891_dout;
  wire       [15:0]   fixTo_1892_dout;
  wire       [15:0]   fixTo_1893_dout;
  wire       [15:0]   fixTo_1894_dout;
  wire       [15:0]   fixTo_1895_dout;
  wire       [31:0]   fixTo_1896_dout;
  wire       [31:0]   fixTo_1897_dout;
  wire       [15:0]   fixTo_1898_dout;
  wire       [15:0]   fixTo_1899_dout;
  wire       [15:0]   fixTo_1900_dout;
  wire       [15:0]   fixTo_1901_dout;
  wire       [31:0]   fixTo_1902_dout;
  wire       [31:0]   fixTo_1903_dout;
  wire       [15:0]   fixTo_1904_dout;
  wire       [15:0]   fixTo_1905_dout;
  wire       [15:0]   fixTo_1906_dout;
  wire       [15:0]   fixTo_1907_dout;
  wire       [31:0]   fixTo_1908_dout;
  wire       [31:0]   fixTo_1909_dout;
  wire       [15:0]   fixTo_1910_dout;
  wire       [15:0]   fixTo_1911_dout;
  wire       [15:0]   fixTo_1912_dout;
  wire       [15:0]   fixTo_1913_dout;
  wire       [31:0]   fixTo_1914_dout;
  wire       [31:0]   fixTo_1915_dout;
  wire       [15:0]   fixTo_1916_dout;
  wire       [15:0]   fixTo_1917_dout;
  wire       [15:0]   fixTo_1918_dout;
  wire       [15:0]   fixTo_1919_dout;
  wire       [31:0]   fixTo_1920_dout;
  wire       [31:0]   fixTo_1921_dout;
  wire       [15:0]   fixTo_1922_dout;
  wire       [15:0]   fixTo_1923_dout;
  wire       [15:0]   fixTo_1924_dout;
  wire       [15:0]   fixTo_1925_dout;
  wire       [31:0]   fixTo_1926_dout;
  wire       [31:0]   fixTo_1927_dout;
  wire       [15:0]   fixTo_1928_dout;
  wire       [15:0]   fixTo_1929_dout;
  wire       [15:0]   fixTo_1930_dout;
  wire       [15:0]   fixTo_1931_dout;
  wire       [31:0]   fixTo_1932_dout;
  wire       [31:0]   fixTo_1933_dout;
  wire       [15:0]   fixTo_1934_dout;
  wire       [15:0]   fixTo_1935_dout;
  wire       [15:0]   fixTo_1936_dout;
  wire       [15:0]   fixTo_1937_dout;
  wire       [31:0]   fixTo_1938_dout;
  wire       [31:0]   fixTo_1939_dout;
  wire       [15:0]   fixTo_1940_dout;
  wire       [15:0]   fixTo_1941_dout;
  wire       [15:0]   fixTo_1942_dout;
  wire       [15:0]   fixTo_1943_dout;
  wire       [31:0]   fixTo_1944_dout;
  wire       [31:0]   fixTo_1945_dout;
  wire       [15:0]   fixTo_1946_dout;
  wire       [15:0]   fixTo_1947_dout;
  wire       [15:0]   fixTo_1948_dout;
  wire       [15:0]   fixTo_1949_dout;
  wire       [31:0]   fixTo_1950_dout;
  wire       [31:0]   fixTo_1951_dout;
  wire       [15:0]   fixTo_1952_dout;
  wire       [15:0]   fixTo_1953_dout;
  wire       [15:0]   fixTo_1954_dout;
  wire       [15:0]   fixTo_1955_dout;
  wire       [31:0]   fixTo_1956_dout;
  wire       [31:0]   fixTo_1957_dout;
  wire       [15:0]   fixTo_1958_dout;
  wire       [15:0]   fixTo_1959_dout;
  wire       [15:0]   fixTo_1960_dout;
  wire       [15:0]   fixTo_1961_dout;
  wire       [31:0]   fixTo_1962_dout;
  wire       [31:0]   fixTo_1963_dout;
  wire       [15:0]   fixTo_1964_dout;
  wire       [15:0]   fixTo_1965_dout;
  wire       [15:0]   fixTo_1966_dout;
  wire       [15:0]   fixTo_1967_dout;
  wire       [31:0]   fixTo_1968_dout;
  wire       [31:0]   fixTo_1969_dout;
  wire       [15:0]   fixTo_1970_dout;
  wire       [15:0]   fixTo_1971_dout;
  wire       [15:0]   fixTo_1972_dout;
  wire       [15:0]   fixTo_1973_dout;
  wire       [31:0]   fixTo_1974_dout;
  wire       [31:0]   fixTo_1975_dout;
  wire       [15:0]   fixTo_1976_dout;
  wire       [15:0]   fixTo_1977_dout;
  wire       [15:0]   fixTo_1978_dout;
  wire       [15:0]   fixTo_1979_dout;
  wire       [31:0]   fixTo_1980_dout;
  wire       [31:0]   fixTo_1981_dout;
  wire       [15:0]   fixTo_1982_dout;
  wire       [15:0]   fixTo_1983_dout;
  wire       [15:0]   fixTo_1984_dout;
  wire       [15:0]   fixTo_1985_dout;
  wire       [31:0]   fixTo_1986_dout;
  wire       [31:0]   fixTo_1987_dout;
  wire       [15:0]   fixTo_1988_dout;
  wire       [15:0]   fixTo_1989_dout;
  wire       [15:0]   fixTo_1990_dout;
  wire       [15:0]   fixTo_1991_dout;
  wire       [31:0]   fixTo_1992_dout;
  wire       [31:0]   fixTo_1993_dout;
  wire       [15:0]   fixTo_1994_dout;
  wire       [15:0]   fixTo_1995_dout;
  wire       [15:0]   fixTo_1996_dout;
  wire       [15:0]   fixTo_1997_dout;
  wire       [31:0]   fixTo_1998_dout;
  wire       [31:0]   fixTo_1999_dout;
  wire       [15:0]   fixTo_2000_dout;
  wire       [15:0]   fixTo_2001_dout;
  wire       [15:0]   fixTo_2002_dout;
  wire       [15:0]   fixTo_2003_dout;
  wire       [31:0]   fixTo_2004_dout;
  wire       [31:0]   fixTo_2005_dout;
  wire       [15:0]   fixTo_2006_dout;
  wire       [15:0]   fixTo_2007_dout;
  wire       [15:0]   fixTo_2008_dout;
  wire       [15:0]   fixTo_2009_dout;
  wire       [31:0]   fixTo_2010_dout;
  wire       [31:0]   fixTo_2011_dout;
  wire       [15:0]   fixTo_2012_dout;
  wire       [15:0]   fixTo_2013_dout;
  wire       [15:0]   fixTo_2014_dout;
  wire       [15:0]   fixTo_2015_dout;
  wire       [31:0]   fixTo_2016_dout;
  wire       [31:0]   fixTo_2017_dout;
  wire       [15:0]   fixTo_2018_dout;
  wire       [15:0]   fixTo_2019_dout;
  wire       [15:0]   fixTo_2020_dout;
  wire       [15:0]   fixTo_2021_dout;
  wire       [31:0]   fixTo_2022_dout;
  wire       [31:0]   fixTo_2023_dout;
  wire       [15:0]   fixTo_2024_dout;
  wire       [15:0]   fixTo_2025_dout;
  wire       [15:0]   fixTo_2026_dout;
  wire       [15:0]   fixTo_2027_dout;
  wire       [31:0]   fixTo_2028_dout;
  wire       [31:0]   fixTo_2029_dout;
  wire       [15:0]   fixTo_2030_dout;
  wire       [15:0]   fixTo_2031_dout;
  wire       [15:0]   fixTo_2032_dout;
  wire       [15:0]   fixTo_2033_dout;
  wire       [31:0]   fixTo_2034_dout;
  wire       [31:0]   fixTo_2035_dout;
  wire       [15:0]   fixTo_2036_dout;
  wire       [15:0]   fixTo_2037_dout;
  wire       [15:0]   fixTo_2038_dout;
  wire       [15:0]   fixTo_2039_dout;
  wire       [31:0]   fixTo_2040_dout;
  wire       [31:0]   fixTo_2041_dout;
  wire       [15:0]   fixTo_2042_dout;
  wire       [15:0]   fixTo_2043_dout;
  wire       [15:0]   fixTo_2044_dout;
  wire       [15:0]   fixTo_2045_dout;
  wire       [31:0]   fixTo_2046_dout;
  wire       [31:0]   fixTo_2047_dout;
  wire       [15:0]   fixTo_2048_dout;
  wire       [15:0]   fixTo_2049_dout;
  wire       [15:0]   fixTo_2050_dout;
  wire       [15:0]   fixTo_2051_dout;
  wire       [31:0]   fixTo_2052_dout;
  wire       [31:0]   fixTo_2053_dout;
  wire       [15:0]   fixTo_2054_dout;
  wire       [15:0]   fixTo_2055_dout;
  wire       [15:0]   fixTo_2056_dout;
  wire       [15:0]   fixTo_2057_dout;
  wire       [31:0]   fixTo_2058_dout;
  wire       [31:0]   fixTo_2059_dout;
  wire       [15:0]   fixTo_2060_dout;
  wire       [15:0]   fixTo_2061_dout;
  wire       [15:0]   fixTo_2062_dout;
  wire       [15:0]   fixTo_2063_dout;
  wire       [31:0]   fixTo_2064_dout;
  wire       [31:0]   fixTo_2065_dout;
  wire       [15:0]   fixTo_2066_dout;
  wire       [15:0]   fixTo_2067_dout;
  wire       [15:0]   fixTo_2068_dout;
  wire       [15:0]   fixTo_2069_dout;
  wire       [31:0]   fixTo_2070_dout;
  wire       [31:0]   fixTo_2071_dout;
  wire       [15:0]   fixTo_2072_dout;
  wire       [15:0]   fixTo_2073_dout;
  wire       [15:0]   fixTo_2074_dout;
  wire       [15:0]   fixTo_2075_dout;
  wire       [31:0]   fixTo_2076_dout;
  wire       [31:0]   fixTo_2077_dout;
  wire       [15:0]   fixTo_2078_dout;
  wire       [15:0]   fixTo_2079_dout;
  wire       [15:0]   fixTo_2080_dout;
  wire       [15:0]   fixTo_2081_dout;
  wire       [31:0]   fixTo_2082_dout;
  wire       [31:0]   fixTo_2083_dout;
  wire       [15:0]   fixTo_2084_dout;
  wire       [15:0]   fixTo_2085_dout;
  wire       [15:0]   fixTo_2086_dout;
  wire       [15:0]   fixTo_2087_dout;
  wire       [31:0]   fixTo_2088_dout;
  wire       [31:0]   fixTo_2089_dout;
  wire       [15:0]   fixTo_2090_dout;
  wire       [15:0]   fixTo_2091_dout;
  wire       [15:0]   fixTo_2092_dout;
  wire       [15:0]   fixTo_2093_dout;
  wire       [31:0]   fixTo_2094_dout;
  wire       [31:0]   fixTo_2095_dout;
  wire       [15:0]   fixTo_2096_dout;
  wire       [15:0]   fixTo_2097_dout;
  wire       [15:0]   fixTo_2098_dout;
  wire       [15:0]   fixTo_2099_dout;
  wire       [31:0]   fixTo_2100_dout;
  wire       [31:0]   fixTo_2101_dout;
  wire       [15:0]   fixTo_2102_dout;
  wire       [15:0]   fixTo_2103_dout;
  wire       [15:0]   fixTo_2104_dout;
  wire       [15:0]   fixTo_2105_dout;
  wire       [31:0]   fixTo_2106_dout;
  wire       [31:0]   fixTo_2107_dout;
  wire       [15:0]   fixTo_2108_dout;
  wire       [15:0]   fixTo_2109_dout;
  wire       [15:0]   fixTo_2110_dout;
  wire       [15:0]   fixTo_2111_dout;
  wire       [31:0]   fixTo_2112_dout;
  wire       [31:0]   fixTo_2113_dout;
  wire       [15:0]   fixTo_2114_dout;
  wire       [15:0]   fixTo_2115_dout;
  wire       [15:0]   fixTo_2116_dout;
  wire       [15:0]   fixTo_2117_dout;
  wire       [31:0]   fixTo_2118_dout;
  wire       [31:0]   fixTo_2119_dout;
  wire       [15:0]   fixTo_2120_dout;
  wire       [15:0]   fixTo_2121_dout;
  wire       [15:0]   fixTo_2122_dout;
  wire       [15:0]   fixTo_2123_dout;
  wire       [31:0]   fixTo_2124_dout;
  wire       [31:0]   fixTo_2125_dout;
  wire       [15:0]   fixTo_2126_dout;
  wire       [15:0]   fixTo_2127_dout;
  wire       [15:0]   fixTo_2128_dout;
  wire       [15:0]   fixTo_2129_dout;
  wire       [31:0]   fixTo_2130_dout;
  wire       [31:0]   fixTo_2131_dout;
  wire       [15:0]   fixTo_2132_dout;
  wire       [15:0]   fixTo_2133_dout;
  wire       [15:0]   fixTo_2134_dout;
  wire       [15:0]   fixTo_2135_dout;
  wire       [31:0]   fixTo_2136_dout;
  wire       [31:0]   fixTo_2137_dout;
  wire       [15:0]   fixTo_2138_dout;
  wire       [15:0]   fixTo_2139_dout;
  wire       [15:0]   fixTo_2140_dout;
  wire       [15:0]   fixTo_2141_dout;
  wire       [31:0]   fixTo_2142_dout;
  wire       [31:0]   fixTo_2143_dout;
  wire       [15:0]   fixTo_2144_dout;
  wire       [15:0]   fixTo_2145_dout;
  wire       [15:0]   fixTo_2146_dout;
  wire       [15:0]   fixTo_2147_dout;
  wire       [31:0]   fixTo_2148_dout;
  wire       [31:0]   fixTo_2149_dout;
  wire       [15:0]   fixTo_2150_dout;
  wire       [15:0]   fixTo_2151_dout;
  wire       [15:0]   fixTo_2152_dout;
  wire       [15:0]   fixTo_2153_dout;
  wire       [31:0]   fixTo_2154_dout;
  wire       [31:0]   fixTo_2155_dout;
  wire       [15:0]   fixTo_2156_dout;
  wire       [15:0]   fixTo_2157_dout;
  wire       [15:0]   fixTo_2158_dout;
  wire       [15:0]   fixTo_2159_dout;
  wire       [31:0]   fixTo_2160_dout;
  wire       [31:0]   fixTo_2161_dout;
  wire       [15:0]   fixTo_2162_dout;
  wire       [15:0]   fixTo_2163_dout;
  wire       [15:0]   fixTo_2164_dout;
  wire       [15:0]   fixTo_2165_dout;
  wire       [31:0]   fixTo_2166_dout;
  wire       [31:0]   fixTo_2167_dout;
  wire       [15:0]   fixTo_2168_dout;
  wire       [15:0]   fixTo_2169_dout;
  wire       [15:0]   fixTo_2170_dout;
  wire       [15:0]   fixTo_2171_dout;
  wire       [31:0]   fixTo_2172_dout;
  wire       [31:0]   fixTo_2173_dout;
  wire       [15:0]   fixTo_2174_dout;
  wire       [15:0]   fixTo_2175_dout;
  wire       [15:0]   fixTo_2176_dout;
  wire       [15:0]   fixTo_2177_dout;
  wire       [31:0]   fixTo_2178_dout;
  wire       [31:0]   fixTo_2179_dout;
  wire       [15:0]   fixTo_2180_dout;
  wire       [15:0]   fixTo_2181_dout;
  wire       [15:0]   fixTo_2182_dout;
  wire       [15:0]   fixTo_2183_dout;
  wire       [31:0]   fixTo_2184_dout;
  wire       [31:0]   fixTo_2185_dout;
  wire       [15:0]   fixTo_2186_dout;
  wire       [15:0]   fixTo_2187_dout;
  wire       [15:0]   fixTo_2188_dout;
  wire       [15:0]   fixTo_2189_dout;
  wire       [31:0]   fixTo_2190_dout;
  wire       [31:0]   fixTo_2191_dout;
  wire       [15:0]   fixTo_2192_dout;
  wire       [15:0]   fixTo_2193_dout;
  wire       [15:0]   fixTo_2194_dout;
  wire       [15:0]   fixTo_2195_dout;
  wire       [31:0]   fixTo_2196_dout;
  wire       [31:0]   fixTo_2197_dout;
  wire       [15:0]   fixTo_2198_dout;
  wire       [15:0]   fixTo_2199_dout;
  wire       [15:0]   fixTo_2200_dout;
  wire       [15:0]   fixTo_2201_dout;
  wire       [31:0]   fixTo_2202_dout;
  wire       [31:0]   fixTo_2203_dout;
  wire       [15:0]   fixTo_2204_dout;
  wire       [15:0]   fixTo_2205_dout;
  wire       [15:0]   fixTo_2206_dout;
  wire       [15:0]   fixTo_2207_dout;
  wire       [31:0]   fixTo_2208_dout;
  wire       [31:0]   fixTo_2209_dout;
  wire       [15:0]   fixTo_2210_dout;
  wire       [15:0]   fixTo_2211_dout;
  wire       [15:0]   fixTo_2212_dout;
  wire       [15:0]   fixTo_2213_dout;
  wire       [31:0]   fixTo_2214_dout;
  wire       [31:0]   fixTo_2215_dout;
  wire       [15:0]   fixTo_2216_dout;
  wire       [15:0]   fixTo_2217_dout;
  wire       [15:0]   fixTo_2218_dout;
  wire       [15:0]   fixTo_2219_dout;
  wire       [31:0]   fixTo_2220_dout;
  wire       [31:0]   fixTo_2221_dout;
  wire       [15:0]   fixTo_2222_dout;
  wire       [15:0]   fixTo_2223_dout;
  wire       [15:0]   fixTo_2224_dout;
  wire       [15:0]   fixTo_2225_dout;
  wire       [31:0]   fixTo_2226_dout;
  wire       [31:0]   fixTo_2227_dout;
  wire       [15:0]   fixTo_2228_dout;
  wire       [15:0]   fixTo_2229_dout;
  wire       [15:0]   fixTo_2230_dout;
  wire       [15:0]   fixTo_2231_dout;
  wire       [31:0]   fixTo_2232_dout;
  wire       [31:0]   fixTo_2233_dout;
  wire       [15:0]   fixTo_2234_dout;
  wire       [15:0]   fixTo_2235_dout;
  wire       [15:0]   fixTo_2236_dout;
  wire       [15:0]   fixTo_2237_dout;
  wire       [31:0]   fixTo_2238_dout;
  wire       [31:0]   fixTo_2239_dout;
  wire       [15:0]   fixTo_2240_dout;
  wire       [15:0]   fixTo_2241_dout;
  wire       [15:0]   fixTo_2242_dout;
  wire       [15:0]   fixTo_2243_dout;
  wire       [31:0]   fixTo_2244_dout;
  wire       [31:0]   fixTo_2245_dout;
  wire       [15:0]   fixTo_2246_dout;
  wire       [15:0]   fixTo_2247_dout;
  wire       [15:0]   fixTo_2248_dout;
  wire       [15:0]   fixTo_2249_dout;
  wire       [31:0]   fixTo_2250_dout;
  wire       [31:0]   fixTo_2251_dout;
  wire       [15:0]   fixTo_2252_dout;
  wire       [15:0]   fixTo_2253_dout;
  wire       [15:0]   fixTo_2254_dout;
  wire       [15:0]   fixTo_2255_dout;
  wire       [31:0]   fixTo_2256_dout;
  wire       [31:0]   fixTo_2257_dout;
  wire       [15:0]   fixTo_2258_dout;
  wire       [15:0]   fixTo_2259_dout;
  wire       [15:0]   fixTo_2260_dout;
  wire       [15:0]   fixTo_2261_dout;
  wire       [31:0]   fixTo_2262_dout;
  wire       [31:0]   fixTo_2263_dout;
  wire       [15:0]   fixTo_2264_dout;
  wire       [15:0]   fixTo_2265_dout;
  wire       [15:0]   fixTo_2266_dout;
  wire       [15:0]   fixTo_2267_dout;
  wire       [31:0]   fixTo_2268_dout;
  wire       [31:0]   fixTo_2269_dout;
  wire       [15:0]   fixTo_2270_dout;
  wire       [15:0]   fixTo_2271_dout;
  wire       [15:0]   fixTo_2272_dout;
  wire       [15:0]   fixTo_2273_dout;
  wire       [31:0]   fixTo_2274_dout;
  wire       [31:0]   fixTo_2275_dout;
  wire       [15:0]   fixTo_2276_dout;
  wire       [15:0]   fixTo_2277_dout;
  wire       [15:0]   fixTo_2278_dout;
  wire       [15:0]   fixTo_2279_dout;
  wire       [31:0]   fixTo_2280_dout;
  wire       [31:0]   fixTo_2281_dout;
  wire       [15:0]   fixTo_2282_dout;
  wire       [15:0]   fixTo_2283_dout;
  wire       [15:0]   fixTo_2284_dout;
  wire       [15:0]   fixTo_2285_dout;
  wire       [31:0]   fixTo_2286_dout;
  wire       [31:0]   fixTo_2287_dout;
  wire       [15:0]   fixTo_2288_dout;
  wire       [15:0]   fixTo_2289_dout;
  wire       [15:0]   fixTo_2290_dout;
  wire       [15:0]   fixTo_2291_dout;
  wire       [31:0]   fixTo_2292_dout;
  wire       [31:0]   fixTo_2293_dout;
  wire       [15:0]   fixTo_2294_dout;
  wire       [15:0]   fixTo_2295_dout;
  wire       [15:0]   fixTo_2296_dout;
  wire       [15:0]   fixTo_2297_dout;
  wire       [31:0]   fixTo_2298_dout;
  wire       [31:0]   fixTo_2299_dout;
  wire       [15:0]   fixTo_2300_dout;
  wire       [15:0]   fixTo_2301_dout;
  wire       [15:0]   fixTo_2302_dout;
  wire       [15:0]   fixTo_2303_dout;
  wire       [31:0]   fixTo_2304_dout;
  wire       [31:0]   fixTo_2305_dout;
  wire       [15:0]   fixTo_2306_dout;
  wire       [15:0]   fixTo_2307_dout;
  wire       [15:0]   fixTo_2308_dout;
  wire       [15:0]   fixTo_2309_dout;
  wire       [31:0]   fixTo_2310_dout;
  wire       [31:0]   fixTo_2311_dout;
  wire       [15:0]   fixTo_2312_dout;
  wire       [15:0]   fixTo_2313_dout;
  wire       [15:0]   fixTo_2314_dout;
  wire       [15:0]   fixTo_2315_dout;
  wire       [31:0]   fixTo_2316_dout;
  wire       [31:0]   fixTo_2317_dout;
  wire       [15:0]   fixTo_2318_dout;
  wire       [15:0]   fixTo_2319_dout;
  wire       [15:0]   fixTo_2320_dout;
  wire       [15:0]   fixTo_2321_dout;
  wire       [31:0]   fixTo_2322_dout;
  wire       [31:0]   fixTo_2323_dout;
  wire       [15:0]   fixTo_2324_dout;
  wire       [15:0]   fixTo_2325_dout;
  wire       [15:0]   fixTo_2326_dout;
  wire       [15:0]   fixTo_2327_dout;
  wire       [31:0]   fixTo_2328_dout;
  wire       [31:0]   fixTo_2329_dout;
  wire       [15:0]   fixTo_2330_dout;
  wire       [15:0]   fixTo_2331_dout;
  wire       [15:0]   fixTo_2332_dout;
  wire       [15:0]   fixTo_2333_dout;
  wire       [31:0]   fixTo_2334_dout;
  wire       [31:0]   fixTo_2335_dout;
  wire       [15:0]   fixTo_2336_dout;
  wire       [15:0]   fixTo_2337_dout;
  wire       [15:0]   fixTo_2338_dout;
  wire       [15:0]   fixTo_2339_dout;
  wire       [31:0]   fixTo_2340_dout;
  wire       [31:0]   fixTo_2341_dout;
  wire       [15:0]   fixTo_2342_dout;
  wire       [15:0]   fixTo_2343_dout;
  wire       [15:0]   fixTo_2344_dout;
  wire       [15:0]   fixTo_2345_dout;
  wire       [31:0]   fixTo_2346_dout;
  wire       [31:0]   fixTo_2347_dout;
  wire       [15:0]   fixTo_2348_dout;
  wire       [15:0]   fixTo_2349_dout;
  wire       [15:0]   fixTo_2350_dout;
  wire       [15:0]   fixTo_2351_dout;
  wire       [31:0]   fixTo_2352_dout;
  wire       [31:0]   fixTo_2353_dout;
  wire       [15:0]   fixTo_2354_dout;
  wire       [15:0]   fixTo_2355_dout;
  wire       [15:0]   fixTo_2356_dout;
  wire       [15:0]   fixTo_2357_dout;
  wire       [31:0]   fixTo_2358_dout;
  wire       [31:0]   fixTo_2359_dout;
  wire       [15:0]   fixTo_2360_dout;
  wire       [15:0]   fixTo_2361_dout;
  wire       [15:0]   fixTo_2362_dout;
  wire       [15:0]   fixTo_2363_dout;
  wire       [31:0]   fixTo_2364_dout;
  wire       [31:0]   fixTo_2365_dout;
  wire       [15:0]   fixTo_2366_dout;
  wire       [15:0]   fixTo_2367_dout;
  wire       [15:0]   fixTo_2368_dout;
  wire       [15:0]   fixTo_2369_dout;
  wire       [31:0]   fixTo_2370_dout;
  wire       [31:0]   fixTo_2371_dout;
  wire       [15:0]   fixTo_2372_dout;
  wire       [15:0]   fixTo_2373_dout;
  wire       [15:0]   fixTo_2374_dout;
  wire       [15:0]   fixTo_2375_dout;
  wire       [31:0]   fixTo_2376_dout;
  wire       [31:0]   fixTo_2377_dout;
  wire       [15:0]   fixTo_2378_dout;
  wire       [15:0]   fixTo_2379_dout;
  wire       [15:0]   fixTo_2380_dout;
  wire       [15:0]   fixTo_2381_dout;
  wire       [31:0]   fixTo_2382_dout;
  wire       [31:0]   fixTo_2383_dout;
  wire       [15:0]   fixTo_2384_dout;
  wire       [15:0]   fixTo_2385_dout;
  wire       [15:0]   fixTo_2386_dout;
  wire       [15:0]   fixTo_2387_dout;
  wire       [31:0]   fixTo_2388_dout;
  wire       [31:0]   fixTo_2389_dout;
  wire       [15:0]   fixTo_2390_dout;
  wire       [15:0]   fixTo_2391_dout;
  wire       [15:0]   fixTo_2392_dout;
  wire       [15:0]   fixTo_2393_dout;
  wire       [31:0]   fixTo_2394_dout;
  wire       [31:0]   fixTo_2395_dout;
  wire       [15:0]   fixTo_2396_dout;
  wire       [15:0]   fixTo_2397_dout;
  wire       [15:0]   fixTo_2398_dout;
  wire       [15:0]   fixTo_2399_dout;
  wire       [31:0]   fixTo_2400_dout;
  wire       [31:0]   fixTo_2401_dout;
  wire       [15:0]   fixTo_2402_dout;
  wire       [15:0]   fixTo_2403_dout;
  wire       [15:0]   fixTo_2404_dout;
  wire       [15:0]   fixTo_2405_dout;
  wire       [31:0]   fixTo_2406_dout;
  wire       [31:0]   fixTo_2407_dout;
  wire       [15:0]   fixTo_2408_dout;
  wire       [15:0]   fixTo_2409_dout;
  wire       [15:0]   fixTo_2410_dout;
  wire       [15:0]   fixTo_2411_dout;
  wire       [31:0]   fixTo_2412_dout;
  wire       [31:0]   fixTo_2413_dout;
  wire       [15:0]   fixTo_2414_dout;
  wire       [15:0]   fixTo_2415_dout;
  wire       [15:0]   fixTo_2416_dout;
  wire       [15:0]   fixTo_2417_dout;
  wire       [31:0]   fixTo_2418_dout;
  wire       [31:0]   fixTo_2419_dout;
  wire       [15:0]   fixTo_2420_dout;
  wire       [15:0]   fixTo_2421_dout;
  wire       [15:0]   fixTo_2422_dout;
  wire       [15:0]   fixTo_2423_dout;
  wire       [31:0]   fixTo_2424_dout;
  wire       [31:0]   fixTo_2425_dout;
  wire       [15:0]   fixTo_2426_dout;
  wire       [15:0]   fixTo_2427_dout;
  wire       [15:0]   fixTo_2428_dout;
  wire       [15:0]   fixTo_2429_dout;
  wire       [31:0]   fixTo_2430_dout;
  wire       [31:0]   fixTo_2431_dout;
  wire       [15:0]   fixTo_2432_dout;
  wire       [15:0]   fixTo_2433_dout;
  wire       [15:0]   fixTo_2434_dout;
  wire       [15:0]   fixTo_2435_dout;
  wire       [31:0]   fixTo_2436_dout;
  wire       [31:0]   fixTo_2437_dout;
  wire       [15:0]   fixTo_2438_dout;
  wire       [15:0]   fixTo_2439_dout;
  wire       [15:0]   fixTo_2440_dout;
  wire       [15:0]   fixTo_2441_dout;
  wire       [31:0]   fixTo_2442_dout;
  wire       [31:0]   fixTo_2443_dout;
  wire       [15:0]   fixTo_2444_dout;
  wire       [15:0]   fixTo_2445_dout;
  wire       [15:0]   fixTo_2446_dout;
  wire       [15:0]   fixTo_2447_dout;
  wire       [31:0]   fixTo_2448_dout;
  wire       [31:0]   fixTo_2449_dout;
  wire       [15:0]   fixTo_2450_dout;
  wire       [15:0]   fixTo_2451_dout;
  wire       [15:0]   fixTo_2452_dout;
  wire       [15:0]   fixTo_2453_dout;
  wire       [31:0]   fixTo_2454_dout;
  wire       [31:0]   fixTo_2455_dout;
  wire       [15:0]   fixTo_2456_dout;
  wire       [15:0]   fixTo_2457_dout;
  wire       [15:0]   fixTo_2458_dout;
  wire       [15:0]   fixTo_2459_dout;
  wire       [31:0]   fixTo_2460_dout;
  wire       [31:0]   fixTo_2461_dout;
  wire       [15:0]   fixTo_2462_dout;
  wire       [15:0]   fixTo_2463_dout;
  wire       [15:0]   fixTo_2464_dout;
  wire       [15:0]   fixTo_2465_dout;
  wire       [31:0]   fixTo_2466_dout;
  wire       [31:0]   fixTo_2467_dout;
  wire       [15:0]   fixTo_2468_dout;
  wire       [15:0]   fixTo_2469_dout;
  wire       [15:0]   fixTo_2470_dout;
  wire       [15:0]   fixTo_2471_dout;
  wire       [31:0]   fixTo_2472_dout;
  wire       [31:0]   fixTo_2473_dout;
  wire       [15:0]   fixTo_2474_dout;
  wire       [15:0]   fixTo_2475_dout;
  wire       [15:0]   fixTo_2476_dout;
  wire       [15:0]   fixTo_2477_dout;
  wire       [31:0]   fixTo_2478_dout;
  wire       [31:0]   fixTo_2479_dout;
  wire       [15:0]   fixTo_2480_dout;
  wire       [15:0]   fixTo_2481_dout;
  wire       [15:0]   fixTo_2482_dout;
  wire       [15:0]   fixTo_2483_dout;
  wire       [31:0]   fixTo_2484_dout;
  wire       [31:0]   fixTo_2485_dout;
  wire       [15:0]   fixTo_2486_dout;
  wire       [15:0]   fixTo_2487_dout;
  wire       [15:0]   fixTo_2488_dout;
  wire       [15:0]   fixTo_2489_dout;
  wire       [31:0]   fixTo_2490_dout;
  wire       [31:0]   fixTo_2491_dout;
  wire       [15:0]   fixTo_2492_dout;
  wire       [15:0]   fixTo_2493_dout;
  wire       [15:0]   fixTo_2494_dout;
  wire       [15:0]   fixTo_2495_dout;
  wire       [31:0]   fixTo_2496_dout;
  wire       [31:0]   fixTo_2497_dout;
  wire       [15:0]   fixTo_2498_dout;
  wire       [15:0]   fixTo_2499_dout;
  wire       [15:0]   fixTo_2500_dout;
  wire       [15:0]   fixTo_2501_dout;
  wire       [31:0]   fixTo_2502_dout;
  wire       [31:0]   fixTo_2503_dout;
  wire       [15:0]   fixTo_2504_dout;
  wire       [15:0]   fixTo_2505_dout;
  wire       [15:0]   fixTo_2506_dout;
  wire       [15:0]   fixTo_2507_dout;
  wire       [31:0]   fixTo_2508_dout;
  wire       [31:0]   fixTo_2509_dout;
  wire       [15:0]   fixTo_2510_dout;
  wire       [15:0]   fixTo_2511_dout;
  wire       [15:0]   fixTo_2512_dout;
  wire       [15:0]   fixTo_2513_dout;
  wire       [31:0]   fixTo_2514_dout;
  wire       [31:0]   fixTo_2515_dout;
  wire       [15:0]   fixTo_2516_dout;
  wire       [15:0]   fixTo_2517_dout;
  wire       [15:0]   fixTo_2518_dout;
  wire       [15:0]   fixTo_2519_dout;
  wire       [31:0]   fixTo_2520_dout;
  wire       [31:0]   fixTo_2521_dout;
  wire       [15:0]   fixTo_2522_dout;
  wire       [15:0]   fixTo_2523_dout;
  wire       [15:0]   fixTo_2524_dout;
  wire       [15:0]   fixTo_2525_dout;
  wire       [31:0]   fixTo_2526_dout;
  wire       [31:0]   fixTo_2527_dout;
  wire       [15:0]   fixTo_2528_dout;
  wire       [15:0]   fixTo_2529_dout;
  wire       [15:0]   fixTo_2530_dout;
  wire       [15:0]   fixTo_2531_dout;
  wire       [31:0]   fixTo_2532_dout;
  wire       [31:0]   fixTo_2533_dout;
  wire       [15:0]   fixTo_2534_dout;
  wire       [15:0]   fixTo_2535_dout;
  wire       [15:0]   fixTo_2536_dout;
  wire       [15:0]   fixTo_2537_dout;
  wire       [31:0]   fixTo_2538_dout;
  wire       [31:0]   fixTo_2539_dout;
  wire       [15:0]   fixTo_2540_dout;
  wire       [15:0]   fixTo_2541_dout;
  wire       [15:0]   fixTo_2542_dout;
  wire       [15:0]   fixTo_2543_dout;
  wire       [31:0]   fixTo_2544_dout;
  wire       [31:0]   fixTo_2545_dout;
  wire       [15:0]   fixTo_2546_dout;
  wire       [15:0]   fixTo_2547_dout;
  wire       [15:0]   fixTo_2548_dout;
  wire       [15:0]   fixTo_2549_dout;
  wire       [31:0]   fixTo_2550_dout;
  wire       [31:0]   fixTo_2551_dout;
  wire       [15:0]   fixTo_2552_dout;
  wire       [15:0]   fixTo_2553_dout;
  wire       [15:0]   fixTo_2554_dout;
  wire       [15:0]   fixTo_2555_dout;
  wire       [31:0]   fixTo_2556_dout;
  wire       [31:0]   fixTo_2557_dout;
  wire       [15:0]   fixTo_2558_dout;
  wire       [15:0]   fixTo_2559_dout;
  wire       [15:0]   fixTo_2560_dout;
  wire       [15:0]   fixTo_2561_dout;
  wire       [31:0]   fixTo_2562_dout;
  wire       [31:0]   fixTo_2563_dout;
  wire       [15:0]   fixTo_2564_dout;
  wire       [15:0]   fixTo_2565_dout;
  wire       [15:0]   fixTo_2566_dout;
  wire       [15:0]   fixTo_2567_dout;
  wire       [31:0]   fixTo_2568_dout;
  wire       [31:0]   fixTo_2569_dout;
  wire       [15:0]   fixTo_2570_dout;
  wire       [15:0]   fixTo_2571_dout;
  wire       [15:0]   fixTo_2572_dout;
  wire       [15:0]   fixTo_2573_dout;
  wire       [31:0]   fixTo_2574_dout;
  wire       [31:0]   fixTo_2575_dout;
  wire       [15:0]   fixTo_2576_dout;
  wire       [15:0]   fixTo_2577_dout;
  wire       [15:0]   fixTo_2578_dout;
  wire       [15:0]   fixTo_2579_dout;
  wire       [31:0]   fixTo_2580_dout;
  wire       [31:0]   fixTo_2581_dout;
  wire       [15:0]   fixTo_2582_dout;
  wire       [15:0]   fixTo_2583_dout;
  wire       [15:0]   fixTo_2584_dout;
  wire       [15:0]   fixTo_2585_dout;
  wire       [31:0]   fixTo_2586_dout;
  wire       [31:0]   fixTo_2587_dout;
  wire       [15:0]   fixTo_2588_dout;
  wire       [15:0]   fixTo_2589_dout;
  wire       [15:0]   fixTo_2590_dout;
  wire       [15:0]   fixTo_2591_dout;
  wire       [31:0]   fixTo_2592_dout;
  wire       [31:0]   fixTo_2593_dout;
  wire       [15:0]   fixTo_2594_dout;
  wire       [15:0]   fixTo_2595_dout;
  wire       [15:0]   fixTo_2596_dout;
  wire       [15:0]   fixTo_2597_dout;
  wire       [31:0]   fixTo_2598_dout;
  wire       [31:0]   fixTo_2599_dout;
  wire       [15:0]   fixTo_2600_dout;
  wire       [15:0]   fixTo_2601_dout;
  wire       [15:0]   fixTo_2602_dout;
  wire       [15:0]   fixTo_2603_dout;
  wire       [31:0]   fixTo_2604_dout;
  wire       [31:0]   fixTo_2605_dout;
  wire       [15:0]   fixTo_2606_dout;
  wire       [15:0]   fixTo_2607_dout;
  wire       [15:0]   fixTo_2608_dout;
  wire       [15:0]   fixTo_2609_dout;
  wire       [31:0]   fixTo_2610_dout;
  wire       [31:0]   fixTo_2611_dout;
  wire       [15:0]   fixTo_2612_dout;
  wire       [15:0]   fixTo_2613_dout;
  wire       [15:0]   fixTo_2614_dout;
  wire       [15:0]   fixTo_2615_dout;
  wire       [31:0]   fixTo_2616_dout;
  wire       [31:0]   fixTo_2617_dout;
  wire       [15:0]   fixTo_2618_dout;
  wire       [15:0]   fixTo_2619_dout;
  wire       [15:0]   fixTo_2620_dout;
  wire       [15:0]   fixTo_2621_dout;
  wire       [31:0]   fixTo_2622_dout;
  wire       [31:0]   fixTo_2623_dout;
  wire       [15:0]   fixTo_2624_dout;
  wire       [15:0]   fixTo_2625_dout;
  wire       [15:0]   fixTo_2626_dout;
  wire       [15:0]   fixTo_2627_dout;
  wire       [31:0]   fixTo_2628_dout;
  wire       [31:0]   fixTo_2629_dout;
  wire       [15:0]   fixTo_2630_dout;
  wire       [15:0]   fixTo_2631_dout;
  wire       [15:0]   fixTo_2632_dout;
  wire       [15:0]   fixTo_2633_dout;
  wire       [31:0]   fixTo_2634_dout;
  wire       [31:0]   fixTo_2635_dout;
  wire       [15:0]   fixTo_2636_dout;
  wire       [15:0]   fixTo_2637_dout;
  wire       [15:0]   fixTo_2638_dout;
  wire       [15:0]   fixTo_2639_dout;
  wire       [31:0]   fixTo_2640_dout;
  wire       [31:0]   fixTo_2641_dout;
  wire       [15:0]   fixTo_2642_dout;
  wire       [15:0]   fixTo_2643_dout;
  wire       [15:0]   fixTo_2644_dout;
  wire       [15:0]   fixTo_2645_dout;
  wire       [31:0]   fixTo_2646_dout;
  wire       [31:0]   fixTo_2647_dout;
  wire       [15:0]   fixTo_2648_dout;
  wire       [15:0]   fixTo_2649_dout;
  wire       [15:0]   fixTo_2650_dout;
  wire       [15:0]   fixTo_2651_dout;
  wire       [31:0]   fixTo_2652_dout;
  wire       [31:0]   fixTo_2653_dout;
  wire       [15:0]   fixTo_2654_dout;
  wire       [15:0]   fixTo_2655_dout;
  wire       [15:0]   fixTo_2656_dout;
  wire       [15:0]   fixTo_2657_dout;
  wire       [31:0]   fixTo_2658_dout;
  wire       [31:0]   fixTo_2659_dout;
  wire       [15:0]   fixTo_2660_dout;
  wire       [15:0]   fixTo_2661_dout;
  wire       [15:0]   fixTo_2662_dout;
  wire       [15:0]   fixTo_2663_dout;
  wire       [31:0]   fixTo_2664_dout;
  wire       [31:0]   fixTo_2665_dout;
  wire       [15:0]   fixTo_2666_dout;
  wire       [15:0]   fixTo_2667_dout;
  wire       [15:0]   fixTo_2668_dout;
  wire       [15:0]   fixTo_2669_dout;
  wire       [31:0]   fixTo_2670_dout;
  wire       [31:0]   fixTo_2671_dout;
  wire       [15:0]   fixTo_2672_dout;
  wire       [15:0]   fixTo_2673_dout;
  wire       [15:0]   fixTo_2674_dout;
  wire       [15:0]   fixTo_2675_dout;
  wire       [31:0]   fixTo_2676_dout;
  wire       [31:0]   fixTo_2677_dout;
  wire       [15:0]   fixTo_2678_dout;
  wire       [15:0]   fixTo_2679_dout;
  wire       [15:0]   fixTo_2680_dout;
  wire       [15:0]   fixTo_2681_dout;
  wire       [31:0]   fixTo_2682_dout;
  wire       [31:0]   fixTo_2683_dout;
  wire       [15:0]   fixTo_2684_dout;
  wire       [15:0]   fixTo_2685_dout;
  wire       [15:0]   fixTo_2686_dout;
  wire       [15:0]   fixTo_2687_dout;
  wire       [0:0]    _zz_4929;
  wire       [2:0]    _zz_4930;
  wire       [15:0]   _zz_4931;
  wire       [31:0]   _zz_4932;
  wire       [31:0]   _zz_4933;
  wire       [15:0]   _zz_4934;
  wire       [31:0]   _zz_4935;
  wire       [31:0]   _zz_4936;
  wire       [31:0]   _zz_4937;
  wire       [15:0]   _zz_4938;
  wire       [31:0]   _zz_4939;
  wire       [31:0]   _zz_4940;
  wire       [31:0]   _zz_4941;
  wire       [31:0]   _zz_4942;
  wire       [31:0]   _zz_4943;
  wire       [31:0]   _zz_4944;
  wire       [23:0]   _zz_4945;
  wire       [31:0]   _zz_4946;
  wire       [15:0]   _zz_4947;
  wire       [31:0]   _zz_4948;
  wire       [31:0]   _zz_4949;
  wire       [31:0]   _zz_4950;
  wire       [31:0]   _zz_4951;
  wire       [31:0]   _zz_4952;
  wire       [23:0]   _zz_4953;
  wire       [31:0]   _zz_4954;
  wire       [15:0]   _zz_4955;
  wire       [31:0]   _zz_4956;
  wire       [31:0]   _zz_4957;
  wire       [31:0]   _zz_4958;
  wire       [31:0]   _zz_4959;
  wire       [31:0]   _zz_4960;
  wire       [23:0]   _zz_4961;
  wire       [31:0]   _zz_4962;
  wire       [15:0]   _zz_4963;
  wire       [31:0]   _zz_4964;
  wire       [31:0]   _zz_4965;
  wire       [31:0]   _zz_4966;
  wire       [31:0]   _zz_4967;
  wire       [31:0]   _zz_4968;
  wire       [23:0]   _zz_4969;
  wire       [31:0]   _zz_4970;
  wire       [15:0]   _zz_4971;
  wire       [15:0]   _zz_4972;
  wire       [31:0]   _zz_4973;
  wire       [31:0]   _zz_4974;
  wire       [15:0]   _zz_4975;
  wire       [31:0]   _zz_4976;
  wire       [31:0]   _zz_4977;
  wire       [31:0]   _zz_4978;
  wire       [15:0]   _zz_4979;
  wire       [31:0]   _zz_4980;
  wire       [31:0]   _zz_4981;
  wire       [31:0]   _zz_4982;
  wire       [31:0]   _zz_4983;
  wire       [31:0]   _zz_4984;
  wire       [31:0]   _zz_4985;
  wire       [23:0]   _zz_4986;
  wire       [31:0]   _zz_4987;
  wire       [15:0]   _zz_4988;
  wire       [31:0]   _zz_4989;
  wire       [31:0]   _zz_4990;
  wire       [31:0]   _zz_4991;
  wire       [31:0]   _zz_4992;
  wire       [31:0]   _zz_4993;
  wire       [23:0]   _zz_4994;
  wire       [31:0]   _zz_4995;
  wire       [15:0]   _zz_4996;
  wire       [31:0]   _zz_4997;
  wire       [31:0]   _zz_4998;
  wire       [31:0]   _zz_4999;
  wire       [31:0]   _zz_5000;
  wire       [31:0]   _zz_5001;
  wire       [23:0]   _zz_5002;
  wire       [31:0]   _zz_5003;
  wire       [15:0]   _zz_5004;
  wire       [31:0]   _zz_5005;
  wire       [31:0]   _zz_5006;
  wire       [31:0]   _zz_5007;
  wire       [31:0]   _zz_5008;
  wire       [31:0]   _zz_5009;
  wire       [23:0]   _zz_5010;
  wire       [31:0]   _zz_5011;
  wire       [15:0]   _zz_5012;
  wire       [15:0]   _zz_5013;
  wire       [31:0]   _zz_5014;
  wire       [31:0]   _zz_5015;
  wire       [15:0]   _zz_5016;
  wire       [31:0]   _zz_5017;
  wire       [31:0]   _zz_5018;
  wire       [31:0]   _zz_5019;
  wire       [15:0]   _zz_5020;
  wire       [31:0]   _zz_5021;
  wire       [31:0]   _zz_5022;
  wire       [31:0]   _zz_5023;
  wire       [31:0]   _zz_5024;
  wire       [31:0]   _zz_5025;
  wire       [31:0]   _zz_5026;
  wire       [23:0]   _zz_5027;
  wire       [31:0]   _zz_5028;
  wire       [15:0]   _zz_5029;
  wire       [31:0]   _zz_5030;
  wire       [31:0]   _zz_5031;
  wire       [31:0]   _zz_5032;
  wire       [31:0]   _zz_5033;
  wire       [31:0]   _zz_5034;
  wire       [23:0]   _zz_5035;
  wire       [31:0]   _zz_5036;
  wire       [15:0]   _zz_5037;
  wire       [31:0]   _zz_5038;
  wire       [31:0]   _zz_5039;
  wire       [31:0]   _zz_5040;
  wire       [31:0]   _zz_5041;
  wire       [31:0]   _zz_5042;
  wire       [23:0]   _zz_5043;
  wire       [31:0]   _zz_5044;
  wire       [15:0]   _zz_5045;
  wire       [31:0]   _zz_5046;
  wire       [31:0]   _zz_5047;
  wire       [31:0]   _zz_5048;
  wire       [31:0]   _zz_5049;
  wire       [31:0]   _zz_5050;
  wire       [23:0]   _zz_5051;
  wire       [31:0]   _zz_5052;
  wire       [15:0]   _zz_5053;
  wire       [15:0]   _zz_5054;
  wire       [31:0]   _zz_5055;
  wire       [31:0]   _zz_5056;
  wire       [15:0]   _zz_5057;
  wire       [31:0]   _zz_5058;
  wire       [31:0]   _zz_5059;
  wire       [31:0]   _zz_5060;
  wire       [15:0]   _zz_5061;
  wire       [31:0]   _zz_5062;
  wire       [31:0]   _zz_5063;
  wire       [31:0]   _zz_5064;
  wire       [31:0]   _zz_5065;
  wire       [31:0]   _zz_5066;
  wire       [31:0]   _zz_5067;
  wire       [23:0]   _zz_5068;
  wire       [31:0]   _zz_5069;
  wire       [15:0]   _zz_5070;
  wire       [31:0]   _zz_5071;
  wire       [31:0]   _zz_5072;
  wire       [31:0]   _zz_5073;
  wire       [31:0]   _zz_5074;
  wire       [31:0]   _zz_5075;
  wire       [23:0]   _zz_5076;
  wire       [31:0]   _zz_5077;
  wire       [15:0]   _zz_5078;
  wire       [31:0]   _zz_5079;
  wire       [31:0]   _zz_5080;
  wire       [31:0]   _zz_5081;
  wire       [31:0]   _zz_5082;
  wire       [31:0]   _zz_5083;
  wire       [23:0]   _zz_5084;
  wire       [31:0]   _zz_5085;
  wire       [15:0]   _zz_5086;
  wire       [31:0]   _zz_5087;
  wire       [31:0]   _zz_5088;
  wire       [31:0]   _zz_5089;
  wire       [31:0]   _zz_5090;
  wire       [31:0]   _zz_5091;
  wire       [23:0]   _zz_5092;
  wire       [31:0]   _zz_5093;
  wire       [15:0]   _zz_5094;
  wire       [15:0]   _zz_5095;
  wire       [31:0]   _zz_5096;
  wire       [31:0]   _zz_5097;
  wire       [15:0]   _zz_5098;
  wire       [31:0]   _zz_5099;
  wire       [31:0]   _zz_5100;
  wire       [31:0]   _zz_5101;
  wire       [15:0]   _zz_5102;
  wire       [31:0]   _zz_5103;
  wire       [31:0]   _zz_5104;
  wire       [31:0]   _zz_5105;
  wire       [31:0]   _zz_5106;
  wire       [31:0]   _zz_5107;
  wire       [31:0]   _zz_5108;
  wire       [23:0]   _zz_5109;
  wire       [31:0]   _zz_5110;
  wire       [15:0]   _zz_5111;
  wire       [31:0]   _zz_5112;
  wire       [31:0]   _zz_5113;
  wire       [31:0]   _zz_5114;
  wire       [31:0]   _zz_5115;
  wire       [31:0]   _zz_5116;
  wire       [23:0]   _zz_5117;
  wire       [31:0]   _zz_5118;
  wire       [15:0]   _zz_5119;
  wire       [31:0]   _zz_5120;
  wire       [31:0]   _zz_5121;
  wire       [31:0]   _zz_5122;
  wire       [31:0]   _zz_5123;
  wire       [31:0]   _zz_5124;
  wire       [23:0]   _zz_5125;
  wire       [31:0]   _zz_5126;
  wire       [15:0]   _zz_5127;
  wire       [31:0]   _zz_5128;
  wire       [31:0]   _zz_5129;
  wire       [31:0]   _zz_5130;
  wire       [31:0]   _zz_5131;
  wire       [31:0]   _zz_5132;
  wire       [23:0]   _zz_5133;
  wire       [31:0]   _zz_5134;
  wire       [15:0]   _zz_5135;
  wire       [15:0]   _zz_5136;
  wire       [31:0]   _zz_5137;
  wire       [31:0]   _zz_5138;
  wire       [15:0]   _zz_5139;
  wire       [31:0]   _zz_5140;
  wire       [31:0]   _zz_5141;
  wire       [31:0]   _zz_5142;
  wire       [15:0]   _zz_5143;
  wire       [31:0]   _zz_5144;
  wire       [31:0]   _zz_5145;
  wire       [31:0]   _zz_5146;
  wire       [31:0]   _zz_5147;
  wire       [31:0]   _zz_5148;
  wire       [31:0]   _zz_5149;
  wire       [23:0]   _zz_5150;
  wire       [31:0]   _zz_5151;
  wire       [15:0]   _zz_5152;
  wire       [31:0]   _zz_5153;
  wire       [31:0]   _zz_5154;
  wire       [31:0]   _zz_5155;
  wire       [31:0]   _zz_5156;
  wire       [31:0]   _zz_5157;
  wire       [23:0]   _zz_5158;
  wire       [31:0]   _zz_5159;
  wire       [15:0]   _zz_5160;
  wire       [31:0]   _zz_5161;
  wire       [31:0]   _zz_5162;
  wire       [31:0]   _zz_5163;
  wire       [31:0]   _zz_5164;
  wire       [31:0]   _zz_5165;
  wire       [23:0]   _zz_5166;
  wire       [31:0]   _zz_5167;
  wire       [15:0]   _zz_5168;
  wire       [31:0]   _zz_5169;
  wire       [31:0]   _zz_5170;
  wire       [31:0]   _zz_5171;
  wire       [31:0]   _zz_5172;
  wire       [31:0]   _zz_5173;
  wire       [23:0]   _zz_5174;
  wire       [31:0]   _zz_5175;
  wire       [15:0]   _zz_5176;
  wire       [15:0]   _zz_5177;
  wire       [31:0]   _zz_5178;
  wire       [31:0]   _zz_5179;
  wire       [15:0]   _zz_5180;
  wire       [31:0]   _zz_5181;
  wire       [31:0]   _zz_5182;
  wire       [31:0]   _zz_5183;
  wire       [15:0]   _zz_5184;
  wire       [31:0]   _zz_5185;
  wire       [31:0]   _zz_5186;
  wire       [31:0]   _zz_5187;
  wire       [31:0]   _zz_5188;
  wire       [31:0]   _zz_5189;
  wire       [31:0]   _zz_5190;
  wire       [23:0]   _zz_5191;
  wire       [31:0]   _zz_5192;
  wire       [15:0]   _zz_5193;
  wire       [31:0]   _zz_5194;
  wire       [31:0]   _zz_5195;
  wire       [31:0]   _zz_5196;
  wire       [31:0]   _zz_5197;
  wire       [31:0]   _zz_5198;
  wire       [23:0]   _zz_5199;
  wire       [31:0]   _zz_5200;
  wire       [15:0]   _zz_5201;
  wire       [31:0]   _zz_5202;
  wire       [31:0]   _zz_5203;
  wire       [31:0]   _zz_5204;
  wire       [31:0]   _zz_5205;
  wire       [31:0]   _zz_5206;
  wire       [23:0]   _zz_5207;
  wire       [31:0]   _zz_5208;
  wire       [15:0]   _zz_5209;
  wire       [31:0]   _zz_5210;
  wire       [31:0]   _zz_5211;
  wire       [31:0]   _zz_5212;
  wire       [31:0]   _zz_5213;
  wire       [31:0]   _zz_5214;
  wire       [23:0]   _zz_5215;
  wire       [31:0]   _zz_5216;
  wire       [15:0]   _zz_5217;
  wire       [15:0]   _zz_5218;
  wire       [31:0]   _zz_5219;
  wire       [31:0]   _zz_5220;
  wire       [15:0]   _zz_5221;
  wire       [31:0]   _zz_5222;
  wire       [31:0]   _zz_5223;
  wire       [31:0]   _zz_5224;
  wire       [15:0]   _zz_5225;
  wire       [31:0]   _zz_5226;
  wire       [31:0]   _zz_5227;
  wire       [31:0]   _zz_5228;
  wire       [31:0]   _zz_5229;
  wire       [31:0]   _zz_5230;
  wire       [31:0]   _zz_5231;
  wire       [23:0]   _zz_5232;
  wire       [31:0]   _zz_5233;
  wire       [15:0]   _zz_5234;
  wire       [31:0]   _zz_5235;
  wire       [31:0]   _zz_5236;
  wire       [31:0]   _zz_5237;
  wire       [31:0]   _zz_5238;
  wire       [31:0]   _zz_5239;
  wire       [23:0]   _zz_5240;
  wire       [31:0]   _zz_5241;
  wire       [15:0]   _zz_5242;
  wire       [31:0]   _zz_5243;
  wire       [31:0]   _zz_5244;
  wire       [31:0]   _zz_5245;
  wire       [31:0]   _zz_5246;
  wire       [31:0]   _zz_5247;
  wire       [23:0]   _zz_5248;
  wire       [31:0]   _zz_5249;
  wire       [15:0]   _zz_5250;
  wire       [31:0]   _zz_5251;
  wire       [31:0]   _zz_5252;
  wire       [31:0]   _zz_5253;
  wire       [31:0]   _zz_5254;
  wire       [31:0]   _zz_5255;
  wire       [23:0]   _zz_5256;
  wire       [31:0]   _zz_5257;
  wire       [15:0]   _zz_5258;
  wire       [15:0]   _zz_5259;
  wire       [31:0]   _zz_5260;
  wire       [31:0]   _zz_5261;
  wire       [15:0]   _zz_5262;
  wire       [31:0]   _zz_5263;
  wire       [31:0]   _zz_5264;
  wire       [31:0]   _zz_5265;
  wire       [15:0]   _zz_5266;
  wire       [31:0]   _zz_5267;
  wire       [31:0]   _zz_5268;
  wire       [31:0]   _zz_5269;
  wire       [31:0]   _zz_5270;
  wire       [31:0]   _zz_5271;
  wire       [31:0]   _zz_5272;
  wire       [23:0]   _zz_5273;
  wire       [31:0]   _zz_5274;
  wire       [15:0]   _zz_5275;
  wire       [31:0]   _zz_5276;
  wire       [31:0]   _zz_5277;
  wire       [31:0]   _zz_5278;
  wire       [31:0]   _zz_5279;
  wire       [31:0]   _zz_5280;
  wire       [23:0]   _zz_5281;
  wire       [31:0]   _zz_5282;
  wire       [15:0]   _zz_5283;
  wire       [31:0]   _zz_5284;
  wire       [31:0]   _zz_5285;
  wire       [31:0]   _zz_5286;
  wire       [31:0]   _zz_5287;
  wire       [31:0]   _zz_5288;
  wire       [23:0]   _zz_5289;
  wire       [31:0]   _zz_5290;
  wire       [15:0]   _zz_5291;
  wire       [31:0]   _zz_5292;
  wire       [31:0]   _zz_5293;
  wire       [31:0]   _zz_5294;
  wire       [31:0]   _zz_5295;
  wire       [31:0]   _zz_5296;
  wire       [23:0]   _zz_5297;
  wire       [31:0]   _zz_5298;
  wire       [15:0]   _zz_5299;
  wire       [15:0]   _zz_5300;
  wire       [31:0]   _zz_5301;
  wire       [31:0]   _zz_5302;
  wire       [15:0]   _zz_5303;
  wire       [31:0]   _zz_5304;
  wire       [31:0]   _zz_5305;
  wire       [31:0]   _zz_5306;
  wire       [15:0]   _zz_5307;
  wire       [31:0]   _zz_5308;
  wire       [31:0]   _zz_5309;
  wire       [31:0]   _zz_5310;
  wire       [31:0]   _zz_5311;
  wire       [31:0]   _zz_5312;
  wire       [31:0]   _zz_5313;
  wire       [23:0]   _zz_5314;
  wire       [31:0]   _zz_5315;
  wire       [15:0]   _zz_5316;
  wire       [31:0]   _zz_5317;
  wire       [31:0]   _zz_5318;
  wire       [31:0]   _zz_5319;
  wire       [31:0]   _zz_5320;
  wire       [31:0]   _zz_5321;
  wire       [23:0]   _zz_5322;
  wire       [31:0]   _zz_5323;
  wire       [15:0]   _zz_5324;
  wire       [31:0]   _zz_5325;
  wire       [31:0]   _zz_5326;
  wire       [31:0]   _zz_5327;
  wire       [31:0]   _zz_5328;
  wire       [31:0]   _zz_5329;
  wire       [23:0]   _zz_5330;
  wire       [31:0]   _zz_5331;
  wire       [15:0]   _zz_5332;
  wire       [31:0]   _zz_5333;
  wire       [31:0]   _zz_5334;
  wire       [31:0]   _zz_5335;
  wire       [31:0]   _zz_5336;
  wire       [31:0]   _zz_5337;
  wire       [23:0]   _zz_5338;
  wire       [31:0]   _zz_5339;
  wire       [15:0]   _zz_5340;
  wire       [15:0]   _zz_5341;
  wire       [31:0]   _zz_5342;
  wire       [31:0]   _zz_5343;
  wire       [15:0]   _zz_5344;
  wire       [31:0]   _zz_5345;
  wire       [31:0]   _zz_5346;
  wire       [31:0]   _zz_5347;
  wire       [15:0]   _zz_5348;
  wire       [31:0]   _zz_5349;
  wire       [31:0]   _zz_5350;
  wire       [31:0]   _zz_5351;
  wire       [31:0]   _zz_5352;
  wire       [31:0]   _zz_5353;
  wire       [31:0]   _zz_5354;
  wire       [23:0]   _zz_5355;
  wire       [31:0]   _zz_5356;
  wire       [15:0]   _zz_5357;
  wire       [31:0]   _zz_5358;
  wire       [31:0]   _zz_5359;
  wire       [31:0]   _zz_5360;
  wire       [31:0]   _zz_5361;
  wire       [31:0]   _zz_5362;
  wire       [23:0]   _zz_5363;
  wire       [31:0]   _zz_5364;
  wire       [15:0]   _zz_5365;
  wire       [31:0]   _zz_5366;
  wire       [31:0]   _zz_5367;
  wire       [31:0]   _zz_5368;
  wire       [31:0]   _zz_5369;
  wire       [31:0]   _zz_5370;
  wire       [23:0]   _zz_5371;
  wire       [31:0]   _zz_5372;
  wire       [15:0]   _zz_5373;
  wire       [31:0]   _zz_5374;
  wire       [31:0]   _zz_5375;
  wire       [31:0]   _zz_5376;
  wire       [31:0]   _zz_5377;
  wire       [31:0]   _zz_5378;
  wire       [23:0]   _zz_5379;
  wire       [31:0]   _zz_5380;
  wire       [15:0]   _zz_5381;
  wire       [15:0]   _zz_5382;
  wire       [31:0]   _zz_5383;
  wire       [31:0]   _zz_5384;
  wire       [15:0]   _zz_5385;
  wire       [31:0]   _zz_5386;
  wire       [31:0]   _zz_5387;
  wire       [31:0]   _zz_5388;
  wire       [15:0]   _zz_5389;
  wire       [31:0]   _zz_5390;
  wire       [31:0]   _zz_5391;
  wire       [31:0]   _zz_5392;
  wire       [31:0]   _zz_5393;
  wire       [31:0]   _zz_5394;
  wire       [31:0]   _zz_5395;
  wire       [23:0]   _zz_5396;
  wire       [31:0]   _zz_5397;
  wire       [15:0]   _zz_5398;
  wire       [31:0]   _zz_5399;
  wire       [31:0]   _zz_5400;
  wire       [31:0]   _zz_5401;
  wire       [31:0]   _zz_5402;
  wire       [31:0]   _zz_5403;
  wire       [23:0]   _zz_5404;
  wire       [31:0]   _zz_5405;
  wire       [15:0]   _zz_5406;
  wire       [31:0]   _zz_5407;
  wire       [31:0]   _zz_5408;
  wire       [31:0]   _zz_5409;
  wire       [31:0]   _zz_5410;
  wire       [31:0]   _zz_5411;
  wire       [23:0]   _zz_5412;
  wire       [31:0]   _zz_5413;
  wire       [15:0]   _zz_5414;
  wire       [31:0]   _zz_5415;
  wire       [31:0]   _zz_5416;
  wire       [31:0]   _zz_5417;
  wire       [31:0]   _zz_5418;
  wire       [31:0]   _zz_5419;
  wire       [23:0]   _zz_5420;
  wire       [31:0]   _zz_5421;
  wire       [15:0]   _zz_5422;
  wire       [15:0]   _zz_5423;
  wire       [31:0]   _zz_5424;
  wire       [31:0]   _zz_5425;
  wire       [15:0]   _zz_5426;
  wire       [31:0]   _zz_5427;
  wire       [31:0]   _zz_5428;
  wire       [31:0]   _zz_5429;
  wire       [15:0]   _zz_5430;
  wire       [31:0]   _zz_5431;
  wire       [31:0]   _zz_5432;
  wire       [31:0]   _zz_5433;
  wire       [31:0]   _zz_5434;
  wire       [31:0]   _zz_5435;
  wire       [31:0]   _zz_5436;
  wire       [23:0]   _zz_5437;
  wire       [31:0]   _zz_5438;
  wire       [15:0]   _zz_5439;
  wire       [31:0]   _zz_5440;
  wire       [31:0]   _zz_5441;
  wire       [31:0]   _zz_5442;
  wire       [31:0]   _zz_5443;
  wire       [31:0]   _zz_5444;
  wire       [23:0]   _zz_5445;
  wire       [31:0]   _zz_5446;
  wire       [15:0]   _zz_5447;
  wire       [31:0]   _zz_5448;
  wire       [31:0]   _zz_5449;
  wire       [31:0]   _zz_5450;
  wire       [31:0]   _zz_5451;
  wire       [31:0]   _zz_5452;
  wire       [23:0]   _zz_5453;
  wire       [31:0]   _zz_5454;
  wire       [15:0]   _zz_5455;
  wire       [31:0]   _zz_5456;
  wire       [31:0]   _zz_5457;
  wire       [31:0]   _zz_5458;
  wire       [31:0]   _zz_5459;
  wire       [31:0]   _zz_5460;
  wire       [23:0]   _zz_5461;
  wire       [31:0]   _zz_5462;
  wire       [15:0]   _zz_5463;
  wire       [15:0]   _zz_5464;
  wire       [31:0]   _zz_5465;
  wire       [31:0]   _zz_5466;
  wire       [15:0]   _zz_5467;
  wire       [31:0]   _zz_5468;
  wire       [31:0]   _zz_5469;
  wire       [31:0]   _zz_5470;
  wire       [15:0]   _zz_5471;
  wire       [31:0]   _zz_5472;
  wire       [31:0]   _zz_5473;
  wire       [31:0]   _zz_5474;
  wire       [31:0]   _zz_5475;
  wire       [31:0]   _zz_5476;
  wire       [31:0]   _zz_5477;
  wire       [23:0]   _zz_5478;
  wire       [31:0]   _zz_5479;
  wire       [15:0]   _zz_5480;
  wire       [31:0]   _zz_5481;
  wire       [31:0]   _zz_5482;
  wire       [31:0]   _zz_5483;
  wire       [31:0]   _zz_5484;
  wire       [31:0]   _zz_5485;
  wire       [23:0]   _zz_5486;
  wire       [31:0]   _zz_5487;
  wire       [15:0]   _zz_5488;
  wire       [31:0]   _zz_5489;
  wire       [31:0]   _zz_5490;
  wire       [31:0]   _zz_5491;
  wire       [31:0]   _zz_5492;
  wire       [31:0]   _zz_5493;
  wire       [23:0]   _zz_5494;
  wire       [31:0]   _zz_5495;
  wire       [15:0]   _zz_5496;
  wire       [31:0]   _zz_5497;
  wire       [31:0]   _zz_5498;
  wire       [31:0]   _zz_5499;
  wire       [31:0]   _zz_5500;
  wire       [31:0]   _zz_5501;
  wire       [23:0]   _zz_5502;
  wire       [31:0]   _zz_5503;
  wire       [15:0]   _zz_5504;
  wire       [15:0]   _zz_5505;
  wire       [31:0]   _zz_5506;
  wire       [31:0]   _zz_5507;
  wire       [15:0]   _zz_5508;
  wire       [31:0]   _zz_5509;
  wire       [31:0]   _zz_5510;
  wire       [31:0]   _zz_5511;
  wire       [15:0]   _zz_5512;
  wire       [31:0]   _zz_5513;
  wire       [31:0]   _zz_5514;
  wire       [31:0]   _zz_5515;
  wire       [31:0]   _zz_5516;
  wire       [31:0]   _zz_5517;
  wire       [31:0]   _zz_5518;
  wire       [23:0]   _zz_5519;
  wire       [31:0]   _zz_5520;
  wire       [15:0]   _zz_5521;
  wire       [31:0]   _zz_5522;
  wire       [31:0]   _zz_5523;
  wire       [31:0]   _zz_5524;
  wire       [31:0]   _zz_5525;
  wire       [31:0]   _zz_5526;
  wire       [23:0]   _zz_5527;
  wire       [31:0]   _zz_5528;
  wire       [15:0]   _zz_5529;
  wire       [31:0]   _zz_5530;
  wire       [31:0]   _zz_5531;
  wire       [31:0]   _zz_5532;
  wire       [31:0]   _zz_5533;
  wire       [31:0]   _zz_5534;
  wire       [23:0]   _zz_5535;
  wire       [31:0]   _zz_5536;
  wire       [15:0]   _zz_5537;
  wire       [31:0]   _zz_5538;
  wire       [31:0]   _zz_5539;
  wire       [31:0]   _zz_5540;
  wire       [31:0]   _zz_5541;
  wire       [31:0]   _zz_5542;
  wire       [23:0]   _zz_5543;
  wire       [31:0]   _zz_5544;
  wire       [15:0]   _zz_5545;
  wire       [15:0]   _zz_5546;
  wire       [31:0]   _zz_5547;
  wire       [31:0]   _zz_5548;
  wire       [15:0]   _zz_5549;
  wire       [31:0]   _zz_5550;
  wire       [31:0]   _zz_5551;
  wire       [31:0]   _zz_5552;
  wire       [15:0]   _zz_5553;
  wire       [31:0]   _zz_5554;
  wire       [31:0]   _zz_5555;
  wire       [31:0]   _zz_5556;
  wire       [31:0]   _zz_5557;
  wire       [31:0]   _zz_5558;
  wire       [31:0]   _zz_5559;
  wire       [23:0]   _zz_5560;
  wire       [31:0]   _zz_5561;
  wire       [15:0]   _zz_5562;
  wire       [31:0]   _zz_5563;
  wire       [31:0]   _zz_5564;
  wire       [31:0]   _zz_5565;
  wire       [31:0]   _zz_5566;
  wire       [31:0]   _zz_5567;
  wire       [23:0]   _zz_5568;
  wire       [31:0]   _zz_5569;
  wire       [15:0]   _zz_5570;
  wire       [31:0]   _zz_5571;
  wire       [31:0]   _zz_5572;
  wire       [31:0]   _zz_5573;
  wire       [31:0]   _zz_5574;
  wire       [31:0]   _zz_5575;
  wire       [23:0]   _zz_5576;
  wire       [31:0]   _zz_5577;
  wire       [15:0]   _zz_5578;
  wire       [31:0]   _zz_5579;
  wire       [31:0]   _zz_5580;
  wire       [31:0]   _zz_5581;
  wire       [31:0]   _zz_5582;
  wire       [31:0]   _zz_5583;
  wire       [23:0]   _zz_5584;
  wire       [31:0]   _zz_5585;
  wire       [15:0]   _zz_5586;
  wire       [15:0]   _zz_5587;
  wire       [31:0]   _zz_5588;
  wire       [31:0]   _zz_5589;
  wire       [15:0]   _zz_5590;
  wire       [31:0]   _zz_5591;
  wire       [31:0]   _zz_5592;
  wire       [31:0]   _zz_5593;
  wire       [15:0]   _zz_5594;
  wire       [31:0]   _zz_5595;
  wire       [31:0]   _zz_5596;
  wire       [31:0]   _zz_5597;
  wire       [31:0]   _zz_5598;
  wire       [31:0]   _zz_5599;
  wire       [31:0]   _zz_5600;
  wire       [23:0]   _zz_5601;
  wire       [31:0]   _zz_5602;
  wire       [15:0]   _zz_5603;
  wire       [31:0]   _zz_5604;
  wire       [31:0]   _zz_5605;
  wire       [31:0]   _zz_5606;
  wire       [31:0]   _zz_5607;
  wire       [31:0]   _zz_5608;
  wire       [23:0]   _zz_5609;
  wire       [31:0]   _zz_5610;
  wire       [15:0]   _zz_5611;
  wire       [31:0]   _zz_5612;
  wire       [31:0]   _zz_5613;
  wire       [31:0]   _zz_5614;
  wire       [31:0]   _zz_5615;
  wire       [31:0]   _zz_5616;
  wire       [23:0]   _zz_5617;
  wire       [31:0]   _zz_5618;
  wire       [15:0]   _zz_5619;
  wire       [31:0]   _zz_5620;
  wire       [31:0]   _zz_5621;
  wire       [31:0]   _zz_5622;
  wire       [31:0]   _zz_5623;
  wire       [31:0]   _zz_5624;
  wire       [23:0]   _zz_5625;
  wire       [31:0]   _zz_5626;
  wire       [15:0]   _zz_5627;
  wire       [15:0]   _zz_5628;
  wire       [31:0]   _zz_5629;
  wire       [31:0]   _zz_5630;
  wire       [15:0]   _zz_5631;
  wire       [31:0]   _zz_5632;
  wire       [31:0]   _zz_5633;
  wire       [31:0]   _zz_5634;
  wire       [15:0]   _zz_5635;
  wire       [31:0]   _zz_5636;
  wire       [31:0]   _zz_5637;
  wire       [31:0]   _zz_5638;
  wire       [31:0]   _zz_5639;
  wire       [31:0]   _zz_5640;
  wire       [31:0]   _zz_5641;
  wire       [23:0]   _zz_5642;
  wire       [31:0]   _zz_5643;
  wire       [15:0]   _zz_5644;
  wire       [31:0]   _zz_5645;
  wire       [31:0]   _zz_5646;
  wire       [31:0]   _zz_5647;
  wire       [31:0]   _zz_5648;
  wire       [31:0]   _zz_5649;
  wire       [23:0]   _zz_5650;
  wire       [31:0]   _zz_5651;
  wire       [15:0]   _zz_5652;
  wire       [31:0]   _zz_5653;
  wire       [31:0]   _zz_5654;
  wire       [31:0]   _zz_5655;
  wire       [31:0]   _zz_5656;
  wire       [31:0]   _zz_5657;
  wire       [23:0]   _zz_5658;
  wire       [31:0]   _zz_5659;
  wire       [15:0]   _zz_5660;
  wire       [31:0]   _zz_5661;
  wire       [31:0]   _zz_5662;
  wire       [31:0]   _zz_5663;
  wire       [31:0]   _zz_5664;
  wire       [31:0]   _zz_5665;
  wire       [23:0]   _zz_5666;
  wire       [31:0]   _zz_5667;
  wire       [15:0]   _zz_5668;
  wire       [15:0]   _zz_5669;
  wire       [31:0]   _zz_5670;
  wire       [31:0]   _zz_5671;
  wire       [15:0]   _zz_5672;
  wire       [31:0]   _zz_5673;
  wire       [31:0]   _zz_5674;
  wire       [31:0]   _zz_5675;
  wire       [15:0]   _zz_5676;
  wire       [31:0]   _zz_5677;
  wire       [31:0]   _zz_5678;
  wire       [31:0]   _zz_5679;
  wire       [31:0]   _zz_5680;
  wire       [31:0]   _zz_5681;
  wire       [31:0]   _zz_5682;
  wire       [23:0]   _zz_5683;
  wire       [31:0]   _zz_5684;
  wire       [15:0]   _zz_5685;
  wire       [31:0]   _zz_5686;
  wire       [31:0]   _zz_5687;
  wire       [31:0]   _zz_5688;
  wire       [31:0]   _zz_5689;
  wire       [31:0]   _zz_5690;
  wire       [23:0]   _zz_5691;
  wire       [31:0]   _zz_5692;
  wire       [15:0]   _zz_5693;
  wire       [31:0]   _zz_5694;
  wire       [31:0]   _zz_5695;
  wire       [31:0]   _zz_5696;
  wire       [31:0]   _zz_5697;
  wire       [31:0]   _zz_5698;
  wire       [23:0]   _zz_5699;
  wire       [31:0]   _zz_5700;
  wire       [15:0]   _zz_5701;
  wire       [31:0]   _zz_5702;
  wire       [31:0]   _zz_5703;
  wire       [31:0]   _zz_5704;
  wire       [31:0]   _zz_5705;
  wire       [31:0]   _zz_5706;
  wire       [23:0]   _zz_5707;
  wire       [31:0]   _zz_5708;
  wire       [15:0]   _zz_5709;
  wire       [15:0]   _zz_5710;
  wire       [31:0]   _zz_5711;
  wire       [31:0]   _zz_5712;
  wire       [15:0]   _zz_5713;
  wire       [31:0]   _zz_5714;
  wire       [31:0]   _zz_5715;
  wire       [31:0]   _zz_5716;
  wire       [15:0]   _zz_5717;
  wire       [31:0]   _zz_5718;
  wire       [31:0]   _zz_5719;
  wire       [31:0]   _zz_5720;
  wire       [31:0]   _zz_5721;
  wire       [31:0]   _zz_5722;
  wire       [31:0]   _zz_5723;
  wire       [23:0]   _zz_5724;
  wire       [31:0]   _zz_5725;
  wire       [15:0]   _zz_5726;
  wire       [31:0]   _zz_5727;
  wire       [31:0]   _zz_5728;
  wire       [31:0]   _zz_5729;
  wire       [31:0]   _zz_5730;
  wire       [31:0]   _zz_5731;
  wire       [23:0]   _zz_5732;
  wire       [31:0]   _zz_5733;
  wire       [15:0]   _zz_5734;
  wire       [31:0]   _zz_5735;
  wire       [31:0]   _zz_5736;
  wire       [31:0]   _zz_5737;
  wire       [31:0]   _zz_5738;
  wire       [31:0]   _zz_5739;
  wire       [23:0]   _zz_5740;
  wire       [31:0]   _zz_5741;
  wire       [15:0]   _zz_5742;
  wire       [31:0]   _zz_5743;
  wire       [31:0]   _zz_5744;
  wire       [31:0]   _zz_5745;
  wire       [31:0]   _zz_5746;
  wire       [31:0]   _zz_5747;
  wire       [23:0]   _zz_5748;
  wire       [31:0]   _zz_5749;
  wire       [15:0]   _zz_5750;
  wire       [15:0]   _zz_5751;
  wire       [31:0]   _zz_5752;
  wire       [31:0]   _zz_5753;
  wire       [15:0]   _zz_5754;
  wire       [31:0]   _zz_5755;
  wire       [31:0]   _zz_5756;
  wire       [31:0]   _zz_5757;
  wire       [15:0]   _zz_5758;
  wire       [31:0]   _zz_5759;
  wire       [31:0]   _zz_5760;
  wire       [31:0]   _zz_5761;
  wire       [31:0]   _zz_5762;
  wire       [31:0]   _zz_5763;
  wire       [31:0]   _zz_5764;
  wire       [23:0]   _zz_5765;
  wire       [31:0]   _zz_5766;
  wire       [15:0]   _zz_5767;
  wire       [31:0]   _zz_5768;
  wire       [31:0]   _zz_5769;
  wire       [31:0]   _zz_5770;
  wire       [31:0]   _zz_5771;
  wire       [31:0]   _zz_5772;
  wire       [23:0]   _zz_5773;
  wire       [31:0]   _zz_5774;
  wire       [15:0]   _zz_5775;
  wire       [31:0]   _zz_5776;
  wire       [31:0]   _zz_5777;
  wire       [31:0]   _zz_5778;
  wire       [31:0]   _zz_5779;
  wire       [31:0]   _zz_5780;
  wire       [23:0]   _zz_5781;
  wire       [31:0]   _zz_5782;
  wire       [15:0]   _zz_5783;
  wire       [31:0]   _zz_5784;
  wire       [31:0]   _zz_5785;
  wire       [31:0]   _zz_5786;
  wire       [31:0]   _zz_5787;
  wire       [31:0]   _zz_5788;
  wire       [23:0]   _zz_5789;
  wire       [31:0]   _zz_5790;
  wire       [15:0]   _zz_5791;
  wire       [15:0]   _zz_5792;
  wire       [31:0]   _zz_5793;
  wire       [31:0]   _zz_5794;
  wire       [15:0]   _zz_5795;
  wire       [31:0]   _zz_5796;
  wire       [31:0]   _zz_5797;
  wire       [31:0]   _zz_5798;
  wire       [15:0]   _zz_5799;
  wire       [31:0]   _zz_5800;
  wire       [31:0]   _zz_5801;
  wire       [31:0]   _zz_5802;
  wire       [31:0]   _zz_5803;
  wire       [31:0]   _zz_5804;
  wire       [31:0]   _zz_5805;
  wire       [23:0]   _zz_5806;
  wire       [31:0]   _zz_5807;
  wire       [15:0]   _zz_5808;
  wire       [31:0]   _zz_5809;
  wire       [31:0]   _zz_5810;
  wire       [31:0]   _zz_5811;
  wire       [31:0]   _zz_5812;
  wire       [31:0]   _zz_5813;
  wire       [23:0]   _zz_5814;
  wire       [31:0]   _zz_5815;
  wire       [15:0]   _zz_5816;
  wire       [31:0]   _zz_5817;
  wire       [31:0]   _zz_5818;
  wire       [31:0]   _zz_5819;
  wire       [31:0]   _zz_5820;
  wire       [31:0]   _zz_5821;
  wire       [23:0]   _zz_5822;
  wire       [31:0]   _zz_5823;
  wire       [15:0]   _zz_5824;
  wire       [31:0]   _zz_5825;
  wire       [31:0]   _zz_5826;
  wire       [31:0]   _zz_5827;
  wire       [31:0]   _zz_5828;
  wire       [31:0]   _zz_5829;
  wire       [23:0]   _zz_5830;
  wire       [31:0]   _zz_5831;
  wire       [15:0]   _zz_5832;
  wire       [15:0]   _zz_5833;
  wire       [31:0]   _zz_5834;
  wire       [31:0]   _zz_5835;
  wire       [15:0]   _zz_5836;
  wire       [31:0]   _zz_5837;
  wire       [31:0]   _zz_5838;
  wire       [31:0]   _zz_5839;
  wire       [15:0]   _zz_5840;
  wire       [31:0]   _zz_5841;
  wire       [31:0]   _zz_5842;
  wire       [31:0]   _zz_5843;
  wire       [31:0]   _zz_5844;
  wire       [31:0]   _zz_5845;
  wire       [31:0]   _zz_5846;
  wire       [23:0]   _zz_5847;
  wire       [31:0]   _zz_5848;
  wire       [15:0]   _zz_5849;
  wire       [31:0]   _zz_5850;
  wire       [31:0]   _zz_5851;
  wire       [31:0]   _zz_5852;
  wire       [31:0]   _zz_5853;
  wire       [31:0]   _zz_5854;
  wire       [23:0]   _zz_5855;
  wire       [31:0]   _zz_5856;
  wire       [15:0]   _zz_5857;
  wire       [31:0]   _zz_5858;
  wire       [31:0]   _zz_5859;
  wire       [31:0]   _zz_5860;
  wire       [31:0]   _zz_5861;
  wire       [31:0]   _zz_5862;
  wire       [23:0]   _zz_5863;
  wire       [31:0]   _zz_5864;
  wire       [15:0]   _zz_5865;
  wire       [31:0]   _zz_5866;
  wire       [31:0]   _zz_5867;
  wire       [31:0]   _zz_5868;
  wire       [31:0]   _zz_5869;
  wire       [31:0]   _zz_5870;
  wire       [23:0]   _zz_5871;
  wire       [31:0]   _zz_5872;
  wire       [15:0]   _zz_5873;
  wire       [15:0]   _zz_5874;
  wire       [31:0]   _zz_5875;
  wire       [31:0]   _zz_5876;
  wire       [15:0]   _zz_5877;
  wire       [31:0]   _zz_5878;
  wire       [31:0]   _zz_5879;
  wire       [31:0]   _zz_5880;
  wire       [15:0]   _zz_5881;
  wire       [31:0]   _zz_5882;
  wire       [31:0]   _zz_5883;
  wire       [31:0]   _zz_5884;
  wire       [31:0]   _zz_5885;
  wire       [31:0]   _zz_5886;
  wire       [31:0]   _zz_5887;
  wire       [23:0]   _zz_5888;
  wire       [31:0]   _zz_5889;
  wire       [15:0]   _zz_5890;
  wire       [31:0]   _zz_5891;
  wire       [31:0]   _zz_5892;
  wire       [31:0]   _zz_5893;
  wire       [31:0]   _zz_5894;
  wire       [31:0]   _zz_5895;
  wire       [23:0]   _zz_5896;
  wire       [31:0]   _zz_5897;
  wire       [15:0]   _zz_5898;
  wire       [31:0]   _zz_5899;
  wire       [31:0]   _zz_5900;
  wire       [31:0]   _zz_5901;
  wire       [31:0]   _zz_5902;
  wire       [31:0]   _zz_5903;
  wire       [23:0]   _zz_5904;
  wire       [31:0]   _zz_5905;
  wire       [15:0]   _zz_5906;
  wire       [31:0]   _zz_5907;
  wire       [31:0]   _zz_5908;
  wire       [31:0]   _zz_5909;
  wire       [31:0]   _zz_5910;
  wire       [31:0]   _zz_5911;
  wire       [23:0]   _zz_5912;
  wire       [31:0]   _zz_5913;
  wire       [15:0]   _zz_5914;
  wire       [15:0]   _zz_5915;
  wire       [31:0]   _zz_5916;
  wire       [31:0]   _zz_5917;
  wire       [15:0]   _zz_5918;
  wire       [31:0]   _zz_5919;
  wire       [31:0]   _zz_5920;
  wire       [31:0]   _zz_5921;
  wire       [15:0]   _zz_5922;
  wire       [31:0]   _zz_5923;
  wire       [31:0]   _zz_5924;
  wire       [31:0]   _zz_5925;
  wire       [31:0]   _zz_5926;
  wire       [31:0]   _zz_5927;
  wire       [31:0]   _zz_5928;
  wire       [23:0]   _zz_5929;
  wire       [31:0]   _zz_5930;
  wire       [15:0]   _zz_5931;
  wire       [31:0]   _zz_5932;
  wire       [31:0]   _zz_5933;
  wire       [31:0]   _zz_5934;
  wire       [31:0]   _zz_5935;
  wire       [31:0]   _zz_5936;
  wire       [23:0]   _zz_5937;
  wire       [31:0]   _zz_5938;
  wire       [15:0]   _zz_5939;
  wire       [31:0]   _zz_5940;
  wire       [31:0]   _zz_5941;
  wire       [31:0]   _zz_5942;
  wire       [31:0]   _zz_5943;
  wire       [31:0]   _zz_5944;
  wire       [23:0]   _zz_5945;
  wire       [31:0]   _zz_5946;
  wire       [15:0]   _zz_5947;
  wire       [31:0]   _zz_5948;
  wire       [31:0]   _zz_5949;
  wire       [31:0]   _zz_5950;
  wire       [31:0]   _zz_5951;
  wire       [31:0]   _zz_5952;
  wire       [23:0]   _zz_5953;
  wire       [31:0]   _zz_5954;
  wire       [15:0]   _zz_5955;
  wire       [15:0]   _zz_5956;
  wire       [31:0]   _zz_5957;
  wire       [31:0]   _zz_5958;
  wire       [15:0]   _zz_5959;
  wire       [31:0]   _zz_5960;
  wire       [31:0]   _zz_5961;
  wire       [31:0]   _zz_5962;
  wire       [15:0]   _zz_5963;
  wire       [31:0]   _zz_5964;
  wire       [31:0]   _zz_5965;
  wire       [31:0]   _zz_5966;
  wire       [31:0]   _zz_5967;
  wire       [31:0]   _zz_5968;
  wire       [31:0]   _zz_5969;
  wire       [23:0]   _zz_5970;
  wire       [31:0]   _zz_5971;
  wire       [15:0]   _zz_5972;
  wire       [31:0]   _zz_5973;
  wire       [31:0]   _zz_5974;
  wire       [31:0]   _zz_5975;
  wire       [31:0]   _zz_5976;
  wire       [31:0]   _zz_5977;
  wire       [23:0]   _zz_5978;
  wire       [31:0]   _zz_5979;
  wire       [15:0]   _zz_5980;
  wire       [31:0]   _zz_5981;
  wire       [31:0]   _zz_5982;
  wire       [31:0]   _zz_5983;
  wire       [31:0]   _zz_5984;
  wire       [31:0]   _zz_5985;
  wire       [23:0]   _zz_5986;
  wire       [31:0]   _zz_5987;
  wire       [15:0]   _zz_5988;
  wire       [31:0]   _zz_5989;
  wire       [31:0]   _zz_5990;
  wire       [31:0]   _zz_5991;
  wire       [31:0]   _zz_5992;
  wire       [31:0]   _zz_5993;
  wire       [23:0]   _zz_5994;
  wire       [31:0]   _zz_5995;
  wire       [15:0]   _zz_5996;
  wire       [15:0]   _zz_5997;
  wire       [31:0]   _zz_5998;
  wire       [31:0]   _zz_5999;
  wire       [15:0]   _zz_6000;
  wire       [31:0]   _zz_6001;
  wire       [31:0]   _zz_6002;
  wire       [31:0]   _zz_6003;
  wire       [15:0]   _zz_6004;
  wire       [31:0]   _zz_6005;
  wire       [31:0]   _zz_6006;
  wire       [31:0]   _zz_6007;
  wire       [31:0]   _zz_6008;
  wire       [31:0]   _zz_6009;
  wire       [31:0]   _zz_6010;
  wire       [23:0]   _zz_6011;
  wire       [31:0]   _zz_6012;
  wire       [15:0]   _zz_6013;
  wire       [31:0]   _zz_6014;
  wire       [31:0]   _zz_6015;
  wire       [31:0]   _zz_6016;
  wire       [31:0]   _zz_6017;
  wire       [31:0]   _zz_6018;
  wire       [23:0]   _zz_6019;
  wire       [31:0]   _zz_6020;
  wire       [15:0]   _zz_6021;
  wire       [31:0]   _zz_6022;
  wire       [31:0]   _zz_6023;
  wire       [31:0]   _zz_6024;
  wire       [31:0]   _zz_6025;
  wire       [31:0]   _zz_6026;
  wire       [23:0]   _zz_6027;
  wire       [31:0]   _zz_6028;
  wire       [15:0]   _zz_6029;
  wire       [31:0]   _zz_6030;
  wire       [31:0]   _zz_6031;
  wire       [31:0]   _zz_6032;
  wire       [31:0]   _zz_6033;
  wire       [31:0]   _zz_6034;
  wire       [23:0]   _zz_6035;
  wire       [31:0]   _zz_6036;
  wire       [15:0]   _zz_6037;
  wire       [15:0]   _zz_6038;
  wire       [31:0]   _zz_6039;
  wire       [31:0]   _zz_6040;
  wire       [15:0]   _zz_6041;
  wire       [31:0]   _zz_6042;
  wire       [31:0]   _zz_6043;
  wire       [31:0]   _zz_6044;
  wire       [15:0]   _zz_6045;
  wire       [31:0]   _zz_6046;
  wire       [31:0]   _zz_6047;
  wire       [31:0]   _zz_6048;
  wire       [31:0]   _zz_6049;
  wire       [31:0]   _zz_6050;
  wire       [31:0]   _zz_6051;
  wire       [23:0]   _zz_6052;
  wire       [31:0]   _zz_6053;
  wire       [15:0]   _zz_6054;
  wire       [31:0]   _zz_6055;
  wire       [31:0]   _zz_6056;
  wire       [31:0]   _zz_6057;
  wire       [31:0]   _zz_6058;
  wire       [31:0]   _zz_6059;
  wire       [23:0]   _zz_6060;
  wire       [31:0]   _zz_6061;
  wire       [15:0]   _zz_6062;
  wire       [31:0]   _zz_6063;
  wire       [31:0]   _zz_6064;
  wire       [31:0]   _zz_6065;
  wire       [31:0]   _zz_6066;
  wire       [31:0]   _zz_6067;
  wire       [23:0]   _zz_6068;
  wire       [31:0]   _zz_6069;
  wire       [15:0]   _zz_6070;
  wire       [31:0]   _zz_6071;
  wire       [31:0]   _zz_6072;
  wire       [31:0]   _zz_6073;
  wire       [31:0]   _zz_6074;
  wire       [31:0]   _zz_6075;
  wire       [23:0]   _zz_6076;
  wire       [31:0]   _zz_6077;
  wire       [15:0]   _zz_6078;
  wire       [15:0]   _zz_6079;
  wire       [31:0]   _zz_6080;
  wire       [31:0]   _zz_6081;
  wire       [15:0]   _zz_6082;
  wire       [31:0]   _zz_6083;
  wire       [31:0]   _zz_6084;
  wire       [31:0]   _zz_6085;
  wire       [15:0]   _zz_6086;
  wire       [31:0]   _zz_6087;
  wire       [31:0]   _zz_6088;
  wire       [31:0]   _zz_6089;
  wire       [31:0]   _zz_6090;
  wire       [31:0]   _zz_6091;
  wire       [31:0]   _zz_6092;
  wire       [23:0]   _zz_6093;
  wire       [31:0]   _zz_6094;
  wire       [15:0]   _zz_6095;
  wire       [31:0]   _zz_6096;
  wire       [31:0]   _zz_6097;
  wire       [31:0]   _zz_6098;
  wire       [31:0]   _zz_6099;
  wire       [31:0]   _zz_6100;
  wire       [23:0]   _zz_6101;
  wire       [31:0]   _zz_6102;
  wire       [15:0]   _zz_6103;
  wire       [31:0]   _zz_6104;
  wire       [31:0]   _zz_6105;
  wire       [31:0]   _zz_6106;
  wire       [31:0]   _zz_6107;
  wire       [31:0]   _zz_6108;
  wire       [23:0]   _zz_6109;
  wire       [31:0]   _zz_6110;
  wire       [15:0]   _zz_6111;
  wire       [31:0]   _zz_6112;
  wire       [31:0]   _zz_6113;
  wire       [31:0]   _zz_6114;
  wire       [31:0]   _zz_6115;
  wire       [31:0]   _zz_6116;
  wire       [23:0]   _zz_6117;
  wire       [31:0]   _zz_6118;
  wire       [15:0]   _zz_6119;
  wire       [15:0]   _zz_6120;
  wire       [31:0]   _zz_6121;
  wire       [31:0]   _zz_6122;
  wire       [15:0]   _zz_6123;
  wire       [31:0]   _zz_6124;
  wire       [31:0]   _zz_6125;
  wire       [31:0]   _zz_6126;
  wire       [15:0]   _zz_6127;
  wire       [31:0]   _zz_6128;
  wire       [31:0]   _zz_6129;
  wire       [31:0]   _zz_6130;
  wire       [31:0]   _zz_6131;
  wire       [31:0]   _zz_6132;
  wire       [31:0]   _zz_6133;
  wire       [23:0]   _zz_6134;
  wire       [31:0]   _zz_6135;
  wire       [15:0]   _zz_6136;
  wire       [31:0]   _zz_6137;
  wire       [31:0]   _zz_6138;
  wire       [31:0]   _zz_6139;
  wire       [31:0]   _zz_6140;
  wire       [31:0]   _zz_6141;
  wire       [23:0]   _zz_6142;
  wire       [31:0]   _zz_6143;
  wire       [15:0]   _zz_6144;
  wire       [31:0]   _zz_6145;
  wire       [31:0]   _zz_6146;
  wire       [31:0]   _zz_6147;
  wire       [31:0]   _zz_6148;
  wire       [31:0]   _zz_6149;
  wire       [23:0]   _zz_6150;
  wire       [31:0]   _zz_6151;
  wire       [15:0]   _zz_6152;
  wire       [31:0]   _zz_6153;
  wire       [31:0]   _zz_6154;
  wire       [31:0]   _zz_6155;
  wire       [31:0]   _zz_6156;
  wire       [31:0]   _zz_6157;
  wire       [23:0]   _zz_6158;
  wire       [31:0]   _zz_6159;
  wire       [15:0]   _zz_6160;
  wire       [15:0]   _zz_6161;
  wire       [31:0]   _zz_6162;
  wire       [31:0]   _zz_6163;
  wire       [15:0]   _zz_6164;
  wire       [31:0]   _zz_6165;
  wire       [31:0]   _zz_6166;
  wire       [31:0]   _zz_6167;
  wire       [15:0]   _zz_6168;
  wire       [31:0]   _zz_6169;
  wire       [31:0]   _zz_6170;
  wire       [31:0]   _zz_6171;
  wire       [31:0]   _zz_6172;
  wire       [31:0]   _zz_6173;
  wire       [31:0]   _zz_6174;
  wire       [23:0]   _zz_6175;
  wire       [31:0]   _zz_6176;
  wire       [15:0]   _zz_6177;
  wire       [31:0]   _zz_6178;
  wire       [31:0]   _zz_6179;
  wire       [31:0]   _zz_6180;
  wire       [31:0]   _zz_6181;
  wire       [31:0]   _zz_6182;
  wire       [23:0]   _zz_6183;
  wire       [31:0]   _zz_6184;
  wire       [15:0]   _zz_6185;
  wire       [31:0]   _zz_6186;
  wire       [31:0]   _zz_6187;
  wire       [31:0]   _zz_6188;
  wire       [31:0]   _zz_6189;
  wire       [31:0]   _zz_6190;
  wire       [23:0]   _zz_6191;
  wire       [31:0]   _zz_6192;
  wire       [15:0]   _zz_6193;
  wire       [31:0]   _zz_6194;
  wire       [31:0]   _zz_6195;
  wire       [31:0]   _zz_6196;
  wire       [31:0]   _zz_6197;
  wire       [31:0]   _zz_6198;
  wire       [23:0]   _zz_6199;
  wire       [31:0]   _zz_6200;
  wire       [15:0]   _zz_6201;
  wire       [15:0]   _zz_6202;
  wire       [31:0]   _zz_6203;
  wire       [31:0]   _zz_6204;
  wire       [15:0]   _zz_6205;
  wire       [31:0]   _zz_6206;
  wire       [31:0]   _zz_6207;
  wire       [31:0]   _zz_6208;
  wire       [15:0]   _zz_6209;
  wire       [31:0]   _zz_6210;
  wire       [31:0]   _zz_6211;
  wire       [31:0]   _zz_6212;
  wire       [31:0]   _zz_6213;
  wire       [31:0]   _zz_6214;
  wire       [31:0]   _zz_6215;
  wire       [23:0]   _zz_6216;
  wire       [31:0]   _zz_6217;
  wire       [15:0]   _zz_6218;
  wire       [31:0]   _zz_6219;
  wire       [31:0]   _zz_6220;
  wire       [31:0]   _zz_6221;
  wire       [31:0]   _zz_6222;
  wire       [31:0]   _zz_6223;
  wire       [23:0]   _zz_6224;
  wire       [31:0]   _zz_6225;
  wire       [15:0]   _zz_6226;
  wire       [31:0]   _zz_6227;
  wire       [31:0]   _zz_6228;
  wire       [31:0]   _zz_6229;
  wire       [31:0]   _zz_6230;
  wire       [31:0]   _zz_6231;
  wire       [23:0]   _zz_6232;
  wire       [31:0]   _zz_6233;
  wire       [15:0]   _zz_6234;
  wire       [31:0]   _zz_6235;
  wire       [31:0]   _zz_6236;
  wire       [31:0]   _zz_6237;
  wire       [31:0]   _zz_6238;
  wire       [31:0]   _zz_6239;
  wire       [23:0]   _zz_6240;
  wire       [31:0]   _zz_6241;
  wire       [15:0]   _zz_6242;
  wire       [15:0]   _zz_6243;
  wire       [31:0]   _zz_6244;
  wire       [31:0]   _zz_6245;
  wire       [15:0]   _zz_6246;
  wire       [31:0]   _zz_6247;
  wire       [31:0]   _zz_6248;
  wire       [31:0]   _zz_6249;
  wire       [15:0]   _zz_6250;
  wire       [31:0]   _zz_6251;
  wire       [31:0]   _zz_6252;
  wire       [31:0]   _zz_6253;
  wire       [31:0]   _zz_6254;
  wire       [31:0]   _zz_6255;
  wire       [31:0]   _zz_6256;
  wire       [23:0]   _zz_6257;
  wire       [31:0]   _zz_6258;
  wire       [15:0]   _zz_6259;
  wire       [31:0]   _zz_6260;
  wire       [31:0]   _zz_6261;
  wire       [31:0]   _zz_6262;
  wire       [31:0]   _zz_6263;
  wire       [31:0]   _zz_6264;
  wire       [23:0]   _zz_6265;
  wire       [31:0]   _zz_6266;
  wire       [15:0]   _zz_6267;
  wire       [31:0]   _zz_6268;
  wire       [31:0]   _zz_6269;
  wire       [31:0]   _zz_6270;
  wire       [31:0]   _zz_6271;
  wire       [31:0]   _zz_6272;
  wire       [23:0]   _zz_6273;
  wire       [31:0]   _zz_6274;
  wire       [15:0]   _zz_6275;
  wire       [31:0]   _zz_6276;
  wire       [31:0]   _zz_6277;
  wire       [31:0]   _zz_6278;
  wire       [31:0]   _zz_6279;
  wire       [31:0]   _zz_6280;
  wire       [23:0]   _zz_6281;
  wire       [31:0]   _zz_6282;
  wire       [15:0]   _zz_6283;
  wire       [15:0]   _zz_6284;
  wire       [31:0]   _zz_6285;
  wire       [31:0]   _zz_6286;
  wire       [15:0]   _zz_6287;
  wire       [31:0]   _zz_6288;
  wire       [31:0]   _zz_6289;
  wire       [31:0]   _zz_6290;
  wire       [15:0]   _zz_6291;
  wire       [31:0]   _zz_6292;
  wire       [31:0]   _zz_6293;
  wire       [31:0]   _zz_6294;
  wire       [31:0]   _zz_6295;
  wire       [31:0]   _zz_6296;
  wire       [31:0]   _zz_6297;
  wire       [23:0]   _zz_6298;
  wire       [31:0]   _zz_6299;
  wire       [15:0]   _zz_6300;
  wire       [31:0]   _zz_6301;
  wire       [31:0]   _zz_6302;
  wire       [31:0]   _zz_6303;
  wire       [31:0]   _zz_6304;
  wire       [31:0]   _zz_6305;
  wire       [23:0]   _zz_6306;
  wire       [31:0]   _zz_6307;
  wire       [15:0]   _zz_6308;
  wire       [31:0]   _zz_6309;
  wire       [31:0]   _zz_6310;
  wire       [31:0]   _zz_6311;
  wire       [31:0]   _zz_6312;
  wire       [31:0]   _zz_6313;
  wire       [23:0]   _zz_6314;
  wire       [31:0]   _zz_6315;
  wire       [15:0]   _zz_6316;
  wire       [31:0]   _zz_6317;
  wire       [31:0]   _zz_6318;
  wire       [31:0]   _zz_6319;
  wire       [31:0]   _zz_6320;
  wire       [31:0]   _zz_6321;
  wire       [23:0]   _zz_6322;
  wire       [31:0]   _zz_6323;
  wire       [15:0]   _zz_6324;
  wire       [15:0]   _zz_6325;
  wire       [31:0]   _zz_6326;
  wire       [31:0]   _zz_6327;
  wire       [15:0]   _zz_6328;
  wire       [31:0]   _zz_6329;
  wire       [31:0]   _zz_6330;
  wire       [31:0]   _zz_6331;
  wire       [15:0]   _zz_6332;
  wire       [31:0]   _zz_6333;
  wire       [31:0]   _zz_6334;
  wire       [31:0]   _zz_6335;
  wire       [31:0]   _zz_6336;
  wire       [31:0]   _zz_6337;
  wire       [31:0]   _zz_6338;
  wire       [23:0]   _zz_6339;
  wire       [31:0]   _zz_6340;
  wire       [15:0]   _zz_6341;
  wire       [31:0]   _zz_6342;
  wire       [31:0]   _zz_6343;
  wire       [31:0]   _zz_6344;
  wire       [31:0]   _zz_6345;
  wire       [31:0]   _zz_6346;
  wire       [23:0]   _zz_6347;
  wire       [31:0]   _zz_6348;
  wire       [15:0]   _zz_6349;
  wire       [31:0]   _zz_6350;
  wire       [31:0]   _zz_6351;
  wire       [31:0]   _zz_6352;
  wire       [31:0]   _zz_6353;
  wire       [31:0]   _zz_6354;
  wire       [23:0]   _zz_6355;
  wire       [31:0]   _zz_6356;
  wire       [15:0]   _zz_6357;
  wire       [31:0]   _zz_6358;
  wire       [31:0]   _zz_6359;
  wire       [31:0]   _zz_6360;
  wire       [31:0]   _zz_6361;
  wire       [31:0]   _zz_6362;
  wire       [23:0]   _zz_6363;
  wire       [31:0]   _zz_6364;
  wire       [15:0]   _zz_6365;
  wire       [15:0]   _zz_6366;
  wire       [31:0]   _zz_6367;
  wire       [31:0]   _zz_6368;
  wire       [15:0]   _zz_6369;
  wire       [31:0]   _zz_6370;
  wire       [31:0]   _zz_6371;
  wire       [31:0]   _zz_6372;
  wire       [15:0]   _zz_6373;
  wire       [31:0]   _zz_6374;
  wire       [31:0]   _zz_6375;
  wire       [31:0]   _zz_6376;
  wire       [31:0]   _zz_6377;
  wire       [31:0]   _zz_6378;
  wire       [31:0]   _zz_6379;
  wire       [23:0]   _zz_6380;
  wire       [31:0]   _zz_6381;
  wire       [15:0]   _zz_6382;
  wire       [31:0]   _zz_6383;
  wire       [31:0]   _zz_6384;
  wire       [31:0]   _zz_6385;
  wire       [31:0]   _zz_6386;
  wire       [31:0]   _zz_6387;
  wire       [23:0]   _zz_6388;
  wire       [31:0]   _zz_6389;
  wire       [15:0]   _zz_6390;
  wire       [31:0]   _zz_6391;
  wire       [31:0]   _zz_6392;
  wire       [31:0]   _zz_6393;
  wire       [31:0]   _zz_6394;
  wire       [31:0]   _zz_6395;
  wire       [23:0]   _zz_6396;
  wire       [31:0]   _zz_6397;
  wire       [15:0]   _zz_6398;
  wire       [31:0]   _zz_6399;
  wire       [31:0]   _zz_6400;
  wire       [31:0]   _zz_6401;
  wire       [31:0]   _zz_6402;
  wire       [31:0]   _zz_6403;
  wire       [23:0]   _zz_6404;
  wire       [31:0]   _zz_6405;
  wire       [15:0]   _zz_6406;
  wire       [15:0]   _zz_6407;
  wire       [31:0]   _zz_6408;
  wire       [31:0]   _zz_6409;
  wire       [15:0]   _zz_6410;
  wire       [31:0]   _zz_6411;
  wire       [31:0]   _zz_6412;
  wire       [31:0]   _zz_6413;
  wire       [15:0]   _zz_6414;
  wire       [31:0]   _zz_6415;
  wire       [31:0]   _zz_6416;
  wire       [31:0]   _zz_6417;
  wire       [31:0]   _zz_6418;
  wire       [31:0]   _zz_6419;
  wire       [31:0]   _zz_6420;
  wire       [23:0]   _zz_6421;
  wire       [31:0]   _zz_6422;
  wire       [15:0]   _zz_6423;
  wire       [31:0]   _zz_6424;
  wire       [31:0]   _zz_6425;
  wire       [31:0]   _zz_6426;
  wire       [31:0]   _zz_6427;
  wire       [31:0]   _zz_6428;
  wire       [23:0]   _zz_6429;
  wire       [31:0]   _zz_6430;
  wire       [15:0]   _zz_6431;
  wire       [31:0]   _zz_6432;
  wire       [31:0]   _zz_6433;
  wire       [31:0]   _zz_6434;
  wire       [31:0]   _zz_6435;
  wire       [31:0]   _zz_6436;
  wire       [23:0]   _zz_6437;
  wire       [31:0]   _zz_6438;
  wire       [15:0]   _zz_6439;
  wire       [31:0]   _zz_6440;
  wire       [31:0]   _zz_6441;
  wire       [31:0]   _zz_6442;
  wire       [31:0]   _zz_6443;
  wire       [31:0]   _zz_6444;
  wire       [23:0]   _zz_6445;
  wire       [31:0]   _zz_6446;
  wire       [15:0]   _zz_6447;
  wire       [15:0]   _zz_6448;
  wire       [31:0]   _zz_6449;
  wire       [31:0]   _zz_6450;
  wire       [15:0]   _zz_6451;
  wire       [31:0]   _zz_6452;
  wire       [31:0]   _zz_6453;
  wire       [31:0]   _zz_6454;
  wire       [15:0]   _zz_6455;
  wire       [31:0]   _zz_6456;
  wire       [31:0]   _zz_6457;
  wire       [31:0]   _zz_6458;
  wire       [31:0]   _zz_6459;
  wire       [31:0]   _zz_6460;
  wire       [31:0]   _zz_6461;
  wire       [23:0]   _zz_6462;
  wire       [31:0]   _zz_6463;
  wire       [15:0]   _zz_6464;
  wire       [31:0]   _zz_6465;
  wire       [31:0]   _zz_6466;
  wire       [31:0]   _zz_6467;
  wire       [31:0]   _zz_6468;
  wire       [31:0]   _zz_6469;
  wire       [23:0]   _zz_6470;
  wire       [31:0]   _zz_6471;
  wire       [15:0]   _zz_6472;
  wire       [31:0]   _zz_6473;
  wire       [31:0]   _zz_6474;
  wire       [31:0]   _zz_6475;
  wire       [31:0]   _zz_6476;
  wire       [31:0]   _zz_6477;
  wire       [23:0]   _zz_6478;
  wire       [31:0]   _zz_6479;
  wire       [15:0]   _zz_6480;
  wire       [31:0]   _zz_6481;
  wire       [31:0]   _zz_6482;
  wire       [31:0]   _zz_6483;
  wire       [31:0]   _zz_6484;
  wire       [31:0]   _zz_6485;
  wire       [23:0]   _zz_6486;
  wire       [31:0]   _zz_6487;
  wire       [15:0]   _zz_6488;
  wire       [15:0]   _zz_6489;
  wire       [31:0]   _zz_6490;
  wire       [31:0]   _zz_6491;
  wire       [15:0]   _zz_6492;
  wire       [31:0]   _zz_6493;
  wire       [31:0]   _zz_6494;
  wire       [31:0]   _zz_6495;
  wire       [15:0]   _zz_6496;
  wire       [31:0]   _zz_6497;
  wire       [31:0]   _zz_6498;
  wire       [31:0]   _zz_6499;
  wire       [31:0]   _zz_6500;
  wire       [31:0]   _zz_6501;
  wire       [31:0]   _zz_6502;
  wire       [23:0]   _zz_6503;
  wire       [31:0]   _zz_6504;
  wire       [15:0]   _zz_6505;
  wire       [31:0]   _zz_6506;
  wire       [31:0]   _zz_6507;
  wire       [31:0]   _zz_6508;
  wire       [31:0]   _zz_6509;
  wire       [31:0]   _zz_6510;
  wire       [23:0]   _zz_6511;
  wire       [31:0]   _zz_6512;
  wire       [15:0]   _zz_6513;
  wire       [31:0]   _zz_6514;
  wire       [31:0]   _zz_6515;
  wire       [31:0]   _zz_6516;
  wire       [31:0]   _zz_6517;
  wire       [31:0]   _zz_6518;
  wire       [23:0]   _zz_6519;
  wire       [31:0]   _zz_6520;
  wire       [15:0]   _zz_6521;
  wire       [31:0]   _zz_6522;
  wire       [31:0]   _zz_6523;
  wire       [31:0]   _zz_6524;
  wire       [31:0]   _zz_6525;
  wire       [31:0]   _zz_6526;
  wire       [23:0]   _zz_6527;
  wire       [31:0]   _zz_6528;
  wire       [15:0]   _zz_6529;
  wire       [15:0]   _zz_6530;
  wire       [31:0]   _zz_6531;
  wire       [31:0]   _zz_6532;
  wire       [15:0]   _zz_6533;
  wire       [31:0]   _zz_6534;
  wire       [31:0]   _zz_6535;
  wire       [31:0]   _zz_6536;
  wire       [15:0]   _zz_6537;
  wire       [31:0]   _zz_6538;
  wire       [31:0]   _zz_6539;
  wire       [31:0]   _zz_6540;
  wire       [31:0]   _zz_6541;
  wire       [31:0]   _zz_6542;
  wire       [31:0]   _zz_6543;
  wire       [23:0]   _zz_6544;
  wire       [31:0]   _zz_6545;
  wire       [15:0]   _zz_6546;
  wire       [31:0]   _zz_6547;
  wire       [31:0]   _zz_6548;
  wire       [31:0]   _zz_6549;
  wire       [31:0]   _zz_6550;
  wire       [31:0]   _zz_6551;
  wire       [23:0]   _zz_6552;
  wire       [31:0]   _zz_6553;
  wire       [15:0]   _zz_6554;
  wire       [31:0]   _zz_6555;
  wire       [31:0]   _zz_6556;
  wire       [31:0]   _zz_6557;
  wire       [31:0]   _zz_6558;
  wire       [31:0]   _zz_6559;
  wire       [23:0]   _zz_6560;
  wire       [31:0]   _zz_6561;
  wire       [15:0]   _zz_6562;
  wire       [31:0]   _zz_6563;
  wire       [31:0]   _zz_6564;
  wire       [31:0]   _zz_6565;
  wire       [31:0]   _zz_6566;
  wire       [31:0]   _zz_6567;
  wire       [23:0]   _zz_6568;
  wire       [31:0]   _zz_6569;
  wire       [15:0]   _zz_6570;
  wire       [15:0]   _zz_6571;
  wire       [31:0]   _zz_6572;
  wire       [31:0]   _zz_6573;
  wire       [15:0]   _zz_6574;
  wire       [31:0]   _zz_6575;
  wire       [31:0]   _zz_6576;
  wire       [31:0]   _zz_6577;
  wire       [15:0]   _zz_6578;
  wire       [31:0]   _zz_6579;
  wire       [31:0]   _zz_6580;
  wire       [31:0]   _zz_6581;
  wire       [31:0]   _zz_6582;
  wire       [31:0]   _zz_6583;
  wire       [31:0]   _zz_6584;
  wire       [23:0]   _zz_6585;
  wire       [31:0]   _zz_6586;
  wire       [15:0]   _zz_6587;
  wire       [31:0]   _zz_6588;
  wire       [31:0]   _zz_6589;
  wire       [31:0]   _zz_6590;
  wire       [31:0]   _zz_6591;
  wire       [31:0]   _zz_6592;
  wire       [23:0]   _zz_6593;
  wire       [31:0]   _zz_6594;
  wire       [15:0]   _zz_6595;
  wire       [31:0]   _zz_6596;
  wire       [31:0]   _zz_6597;
  wire       [31:0]   _zz_6598;
  wire       [31:0]   _zz_6599;
  wire       [31:0]   _zz_6600;
  wire       [23:0]   _zz_6601;
  wire       [31:0]   _zz_6602;
  wire       [15:0]   _zz_6603;
  wire       [31:0]   _zz_6604;
  wire       [31:0]   _zz_6605;
  wire       [31:0]   _zz_6606;
  wire       [31:0]   _zz_6607;
  wire       [31:0]   _zz_6608;
  wire       [23:0]   _zz_6609;
  wire       [31:0]   _zz_6610;
  wire       [15:0]   _zz_6611;
  wire       [15:0]   _zz_6612;
  wire       [31:0]   _zz_6613;
  wire       [31:0]   _zz_6614;
  wire       [15:0]   _zz_6615;
  wire       [31:0]   _zz_6616;
  wire       [31:0]   _zz_6617;
  wire       [31:0]   _zz_6618;
  wire       [15:0]   _zz_6619;
  wire       [31:0]   _zz_6620;
  wire       [31:0]   _zz_6621;
  wire       [31:0]   _zz_6622;
  wire       [31:0]   _zz_6623;
  wire       [31:0]   _zz_6624;
  wire       [31:0]   _zz_6625;
  wire       [23:0]   _zz_6626;
  wire       [31:0]   _zz_6627;
  wire       [15:0]   _zz_6628;
  wire       [31:0]   _zz_6629;
  wire       [31:0]   _zz_6630;
  wire       [31:0]   _zz_6631;
  wire       [31:0]   _zz_6632;
  wire       [31:0]   _zz_6633;
  wire       [23:0]   _zz_6634;
  wire       [31:0]   _zz_6635;
  wire       [15:0]   _zz_6636;
  wire       [31:0]   _zz_6637;
  wire       [31:0]   _zz_6638;
  wire       [31:0]   _zz_6639;
  wire       [31:0]   _zz_6640;
  wire       [31:0]   _zz_6641;
  wire       [23:0]   _zz_6642;
  wire       [31:0]   _zz_6643;
  wire       [15:0]   _zz_6644;
  wire       [31:0]   _zz_6645;
  wire       [31:0]   _zz_6646;
  wire       [31:0]   _zz_6647;
  wire       [31:0]   _zz_6648;
  wire       [31:0]   _zz_6649;
  wire       [23:0]   _zz_6650;
  wire       [31:0]   _zz_6651;
  wire       [15:0]   _zz_6652;
  wire       [15:0]   _zz_6653;
  wire       [31:0]   _zz_6654;
  wire       [31:0]   _zz_6655;
  wire       [15:0]   _zz_6656;
  wire       [31:0]   _zz_6657;
  wire       [31:0]   _zz_6658;
  wire       [31:0]   _zz_6659;
  wire       [15:0]   _zz_6660;
  wire       [31:0]   _zz_6661;
  wire       [31:0]   _zz_6662;
  wire       [31:0]   _zz_6663;
  wire       [31:0]   _zz_6664;
  wire       [31:0]   _zz_6665;
  wire       [31:0]   _zz_6666;
  wire       [23:0]   _zz_6667;
  wire       [31:0]   _zz_6668;
  wire       [15:0]   _zz_6669;
  wire       [31:0]   _zz_6670;
  wire       [31:0]   _zz_6671;
  wire       [31:0]   _zz_6672;
  wire       [31:0]   _zz_6673;
  wire       [31:0]   _zz_6674;
  wire       [23:0]   _zz_6675;
  wire       [31:0]   _zz_6676;
  wire       [15:0]   _zz_6677;
  wire       [31:0]   _zz_6678;
  wire       [31:0]   _zz_6679;
  wire       [31:0]   _zz_6680;
  wire       [31:0]   _zz_6681;
  wire       [31:0]   _zz_6682;
  wire       [23:0]   _zz_6683;
  wire       [31:0]   _zz_6684;
  wire       [15:0]   _zz_6685;
  wire       [31:0]   _zz_6686;
  wire       [31:0]   _zz_6687;
  wire       [31:0]   _zz_6688;
  wire       [31:0]   _zz_6689;
  wire       [31:0]   _zz_6690;
  wire       [23:0]   _zz_6691;
  wire       [31:0]   _zz_6692;
  wire       [15:0]   _zz_6693;
  wire       [15:0]   _zz_6694;
  wire       [31:0]   _zz_6695;
  wire       [31:0]   _zz_6696;
  wire       [15:0]   _zz_6697;
  wire       [31:0]   _zz_6698;
  wire       [31:0]   _zz_6699;
  wire       [31:0]   _zz_6700;
  wire       [15:0]   _zz_6701;
  wire       [31:0]   _zz_6702;
  wire       [31:0]   _zz_6703;
  wire       [31:0]   _zz_6704;
  wire       [31:0]   _zz_6705;
  wire       [31:0]   _zz_6706;
  wire       [31:0]   _zz_6707;
  wire       [23:0]   _zz_6708;
  wire       [31:0]   _zz_6709;
  wire       [15:0]   _zz_6710;
  wire       [31:0]   _zz_6711;
  wire       [31:0]   _zz_6712;
  wire       [31:0]   _zz_6713;
  wire       [31:0]   _zz_6714;
  wire       [31:0]   _zz_6715;
  wire       [23:0]   _zz_6716;
  wire       [31:0]   _zz_6717;
  wire       [15:0]   _zz_6718;
  wire       [31:0]   _zz_6719;
  wire       [31:0]   _zz_6720;
  wire       [31:0]   _zz_6721;
  wire       [31:0]   _zz_6722;
  wire       [31:0]   _zz_6723;
  wire       [23:0]   _zz_6724;
  wire       [31:0]   _zz_6725;
  wire       [15:0]   _zz_6726;
  wire       [31:0]   _zz_6727;
  wire       [31:0]   _zz_6728;
  wire       [31:0]   _zz_6729;
  wire       [31:0]   _zz_6730;
  wire       [31:0]   _zz_6731;
  wire       [23:0]   _zz_6732;
  wire       [31:0]   _zz_6733;
  wire       [15:0]   _zz_6734;
  wire       [15:0]   _zz_6735;
  wire       [31:0]   _zz_6736;
  wire       [31:0]   _zz_6737;
  wire       [15:0]   _zz_6738;
  wire       [31:0]   _zz_6739;
  wire       [31:0]   _zz_6740;
  wire       [31:0]   _zz_6741;
  wire       [15:0]   _zz_6742;
  wire       [31:0]   _zz_6743;
  wire       [31:0]   _zz_6744;
  wire       [31:0]   _zz_6745;
  wire       [31:0]   _zz_6746;
  wire       [31:0]   _zz_6747;
  wire       [31:0]   _zz_6748;
  wire       [23:0]   _zz_6749;
  wire       [31:0]   _zz_6750;
  wire       [15:0]   _zz_6751;
  wire       [31:0]   _zz_6752;
  wire       [31:0]   _zz_6753;
  wire       [31:0]   _zz_6754;
  wire       [31:0]   _zz_6755;
  wire       [31:0]   _zz_6756;
  wire       [23:0]   _zz_6757;
  wire       [31:0]   _zz_6758;
  wire       [15:0]   _zz_6759;
  wire       [31:0]   _zz_6760;
  wire       [31:0]   _zz_6761;
  wire       [31:0]   _zz_6762;
  wire       [31:0]   _zz_6763;
  wire       [31:0]   _zz_6764;
  wire       [23:0]   _zz_6765;
  wire       [31:0]   _zz_6766;
  wire       [15:0]   _zz_6767;
  wire       [31:0]   _zz_6768;
  wire       [31:0]   _zz_6769;
  wire       [31:0]   _zz_6770;
  wire       [31:0]   _zz_6771;
  wire       [31:0]   _zz_6772;
  wire       [23:0]   _zz_6773;
  wire       [31:0]   _zz_6774;
  wire       [15:0]   _zz_6775;
  wire       [15:0]   _zz_6776;
  wire       [31:0]   _zz_6777;
  wire       [31:0]   _zz_6778;
  wire       [15:0]   _zz_6779;
  wire       [31:0]   _zz_6780;
  wire       [31:0]   _zz_6781;
  wire       [31:0]   _zz_6782;
  wire       [15:0]   _zz_6783;
  wire       [31:0]   _zz_6784;
  wire       [31:0]   _zz_6785;
  wire       [31:0]   _zz_6786;
  wire       [31:0]   _zz_6787;
  wire       [31:0]   _zz_6788;
  wire       [31:0]   _zz_6789;
  wire       [23:0]   _zz_6790;
  wire       [31:0]   _zz_6791;
  wire       [15:0]   _zz_6792;
  wire       [31:0]   _zz_6793;
  wire       [31:0]   _zz_6794;
  wire       [31:0]   _zz_6795;
  wire       [31:0]   _zz_6796;
  wire       [31:0]   _zz_6797;
  wire       [23:0]   _zz_6798;
  wire       [31:0]   _zz_6799;
  wire       [15:0]   _zz_6800;
  wire       [31:0]   _zz_6801;
  wire       [31:0]   _zz_6802;
  wire       [31:0]   _zz_6803;
  wire       [31:0]   _zz_6804;
  wire       [31:0]   _zz_6805;
  wire       [23:0]   _zz_6806;
  wire       [31:0]   _zz_6807;
  wire       [15:0]   _zz_6808;
  wire       [31:0]   _zz_6809;
  wire       [31:0]   _zz_6810;
  wire       [31:0]   _zz_6811;
  wire       [31:0]   _zz_6812;
  wire       [31:0]   _zz_6813;
  wire       [23:0]   _zz_6814;
  wire       [31:0]   _zz_6815;
  wire       [15:0]   _zz_6816;
  wire       [15:0]   _zz_6817;
  wire       [31:0]   _zz_6818;
  wire       [31:0]   _zz_6819;
  wire       [15:0]   _zz_6820;
  wire       [31:0]   _zz_6821;
  wire       [31:0]   _zz_6822;
  wire       [31:0]   _zz_6823;
  wire       [15:0]   _zz_6824;
  wire       [31:0]   _zz_6825;
  wire       [31:0]   _zz_6826;
  wire       [31:0]   _zz_6827;
  wire       [31:0]   _zz_6828;
  wire       [31:0]   _zz_6829;
  wire       [31:0]   _zz_6830;
  wire       [23:0]   _zz_6831;
  wire       [31:0]   _zz_6832;
  wire       [15:0]   _zz_6833;
  wire       [31:0]   _zz_6834;
  wire       [31:0]   _zz_6835;
  wire       [31:0]   _zz_6836;
  wire       [31:0]   _zz_6837;
  wire       [31:0]   _zz_6838;
  wire       [23:0]   _zz_6839;
  wire       [31:0]   _zz_6840;
  wire       [15:0]   _zz_6841;
  wire       [31:0]   _zz_6842;
  wire       [31:0]   _zz_6843;
  wire       [31:0]   _zz_6844;
  wire       [31:0]   _zz_6845;
  wire       [31:0]   _zz_6846;
  wire       [23:0]   _zz_6847;
  wire       [31:0]   _zz_6848;
  wire       [15:0]   _zz_6849;
  wire       [31:0]   _zz_6850;
  wire       [31:0]   _zz_6851;
  wire       [31:0]   _zz_6852;
  wire       [31:0]   _zz_6853;
  wire       [31:0]   _zz_6854;
  wire       [23:0]   _zz_6855;
  wire       [31:0]   _zz_6856;
  wire       [15:0]   _zz_6857;
  wire       [15:0]   _zz_6858;
  wire       [31:0]   _zz_6859;
  wire       [31:0]   _zz_6860;
  wire       [15:0]   _zz_6861;
  wire       [31:0]   _zz_6862;
  wire       [31:0]   _zz_6863;
  wire       [31:0]   _zz_6864;
  wire       [15:0]   _zz_6865;
  wire       [31:0]   _zz_6866;
  wire       [31:0]   _zz_6867;
  wire       [31:0]   _zz_6868;
  wire       [31:0]   _zz_6869;
  wire       [31:0]   _zz_6870;
  wire       [31:0]   _zz_6871;
  wire       [23:0]   _zz_6872;
  wire       [31:0]   _zz_6873;
  wire       [15:0]   _zz_6874;
  wire       [31:0]   _zz_6875;
  wire       [31:0]   _zz_6876;
  wire       [31:0]   _zz_6877;
  wire       [31:0]   _zz_6878;
  wire       [31:0]   _zz_6879;
  wire       [23:0]   _zz_6880;
  wire       [31:0]   _zz_6881;
  wire       [15:0]   _zz_6882;
  wire       [31:0]   _zz_6883;
  wire       [31:0]   _zz_6884;
  wire       [31:0]   _zz_6885;
  wire       [31:0]   _zz_6886;
  wire       [31:0]   _zz_6887;
  wire       [23:0]   _zz_6888;
  wire       [31:0]   _zz_6889;
  wire       [15:0]   _zz_6890;
  wire       [31:0]   _zz_6891;
  wire       [31:0]   _zz_6892;
  wire       [31:0]   _zz_6893;
  wire       [31:0]   _zz_6894;
  wire       [31:0]   _zz_6895;
  wire       [23:0]   _zz_6896;
  wire       [31:0]   _zz_6897;
  wire       [15:0]   _zz_6898;
  wire       [15:0]   _zz_6899;
  wire       [31:0]   _zz_6900;
  wire       [31:0]   _zz_6901;
  wire       [15:0]   _zz_6902;
  wire       [31:0]   _zz_6903;
  wire       [31:0]   _zz_6904;
  wire       [31:0]   _zz_6905;
  wire       [15:0]   _zz_6906;
  wire       [31:0]   _zz_6907;
  wire       [31:0]   _zz_6908;
  wire       [31:0]   _zz_6909;
  wire       [31:0]   _zz_6910;
  wire       [31:0]   _zz_6911;
  wire       [31:0]   _zz_6912;
  wire       [23:0]   _zz_6913;
  wire       [31:0]   _zz_6914;
  wire       [15:0]   _zz_6915;
  wire       [31:0]   _zz_6916;
  wire       [31:0]   _zz_6917;
  wire       [31:0]   _zz_6918;
  wire       [31:0]   _zz_6919;
  wire       [31:0]   _zz_6920;
  wire       [23:0]   _zz_6921;
  wire       [31:0]   _zz_6922;
  wire       [15:0]   _zz_6923;
  wire       [31:0]   _zz_6924;
  wire       [31:0]   _zz_6925;
  wire       [31:0]   _zz_6926;
  wire       [31:0]   _zz_6927;
  wire       [31:0]   _zz_6928;
  wire       [23:0]   _zz_6929;
  wire       [31:0]   _zz_6930;
  wire       [15:0]   _zz_6931;
  wire       [31:0]   _zz_6932;
  wire       [31:0]   _zz_6933;
  wire       [31:0]   _zz_6934;
  wire       [31:0]   _zz_6935;
  wire       [31:0]   _zz_6936;
  wire       [23:0]   _zz_6937;
  wire       [31:0]   _zz_6938;
  wire       [15:0]   _zz_6939;
  wire       [15:0]   _zz_6940;
  wire       [31:0]   _zz_6941;
  wire       [31:0]   _zz_6942;
  wire       [15:0]   _zz_6943;
  wire       [31:0]   _zz_6944;
  wire       [31:0]   _zz_6945;
  wire       [31:0]   _zz_6946;
  wire       [15:0]   _zz_6947;
  wire       [31:0]   _zz_6948;
  wire       [31:0]   _zz_6949;
  wire       [31:0]   _zz_6950;
  wire       [31:0]   _zz_6951;
  wire       [31:0]   _zz_6952;
  wire       [31:0]   _zz_6953;
  wire       [23:0]   _zz_6954;
  wire       [31:0]   _zz_6955;
  wire       [15:0]   _zz_6956;
  wire       [31:0]   _zz_6957;
  wire       [31:0]   _zz_6958;
  wire       [31:0]   _zz_6959;
  wire       [31:0]   _zz_6960;
  wire       [31:0]   _zz_6961;
  wire       [23:0]   _zz_6962;
  wire       [31:0]   _zz_6963;
  wire       [15:0]   _zz_6964;
  wire       [31:0]   _zz_6965;
  wire       [31:0]   _zz_6966;
  wire       [31:0]   _zz_6967;
  wire       [31:0]   _zz_6968;
  wire       [31:0]   _zz_6969;
  wire       [23:0]   _zz_6970;
  wire       [31:0]   _zz_6971;
  wire       [15:0]   _zz_6972;
  wire       [31:0]   _zz_6973;
  wire       [31:0]   _zz_6974;
  wire       [31:0]   _zz_6975;
  wire       [31:0]   _zz_6976;
  wire       [31:0]   _zz_6977;
  wire       [23:0]   _zz_6978;
  wire       [31:0]   _zz_6979;
  wire       [15:0]   _zz_6980;
  wire       [15:0]   _zz_6981;
  wire       [31:0]   _zz_6982;
  wire       [31:0]   _zz_6983;
  wire       [15:0]   _zz_6984;
  wire       [31:0]   _zz_6985;
  wire       [31:0]   _zz_6986;
  wire       [31:0]   _zz_6987;
  wire       [15:0]   _zz_6988;
  wire       [31:0]   _zz_6989;
  wire       [31:0]   _zz_6990;
  wire       [31:0]   _zz_6991;
  wire       [31:0]   _zz_6992;
  wire       [31:0]   _zz_6993;
  wire       [31:0]   _zz_6994;
  wire       [23:0]   _zz_6995;
  wire       [31:0]   _zz_6996;
  wire       [15:0]   _zz_6997;
  wire       [31:0]   _zz_6998;
  wire       [31:0]   _zz_6999;
  wire       [31:0]   _zz_7000;
  wire       [31:0]   _zz_7001;
  wire       [31:0]   _zz_7002;
  wire       [23:0]   _zz_7003;
  wire       [31:0]   _zz_7004;
  wire       [15:0]   _zz_7005;
  wire       [31:0]   _zz_7006;
  wire       [31:0]   _zz_7007;
  wire       [31:0]   _zz_7008;
  wire       [31:0]   _zz_7009;
  wire       [31:0]   _zz_7010;
  wire       [23:0]   _zz_7011;
  wire       [31:0]   _zz_7012;
  wire       [15:0]   _zz_7013;
  wire       [31:0]   _zz_7014;
  wire       [31:0]   _zz_7015;
  wire       [31:0]   _zz_7016;
  wire       [31:0]   _zz_7017;
  wire       [31:0]   _zz_7018;
  wire       [23:0]   _zz_7019;
  wire       [31:0]   _zz_7020;
  wire       [15:0]   _zz_7021;
  wire       [15:0]   _zz_7022;
  wire       [31:0]   _zz_7023;
  wire       [31:0]   _zz_7024;
  wire       [15:0]   _zz_7025;
  wire       [31:0]   _zz_7026;
  wire       [31:0]   _zz_7027;
  wire       [31:0]   _zz_7028;
  wire       [15:0]   _zz_7029;
  wire       [31:0]   _zz_7030;
  wire       [31:0]   _zz_7031;
  wire       [31:0]   _zz_7032;
  wire       [31:0]   _zz_7033;
  wire       [31:0]   _zz_7034;
  wire       [31:0]   _zz_7035;
  wire       [23:0]   _zz_7036;
  wire       [31:0]   _zz_7037;
  wire       [15:0]   _zz_7038;
  wire       [31:0]   _zz_7039;
  wire       [31:0]   _zz_7040;
  wire       [31:0]   _zz_7041;
  wire       [31:0]   _zz_7042;
  wire       [31:0]   _zz_7043;
  wire       [23:0]   _zz_7044;
  wire       [31:0]   _zz_7045;
  wire       [15:0]   _zz_7046;
  wire       [31:0]   _zz_7047;
  wire       [31:0]   _zz_7048;
  wire       [31:0]   _zz_7049;
  wire       [31:0]   _zz_7050;
  wire       [31:0]   _zz_7051;
  wire       [23:0]   _zz_7052;
  wire       [31:0]   _zz_7053;
  wire       [15:0]   _zz_7054;
  wire       [31:0]   _zz_7055;
  wire       [31:0]   _zz_7056;
  wire       [31:0]   _zz_7057;
  wire       [31:0]   _zz_7058;
  wire       [31:0]   _zz_7059;
  wire       [23:0]   _zz_7060;
  wire       [31:0]   _zz_7061;
  wire       [15:0]   _zz_7062;
  wire       [15:0]   _zz_7063;
  wire       [31:0]   _zz_7064;
  wire       [31:0]   _zz_7065;
  wire       [15:0]   _zz_7066;
  wire       [31:0]   _zz_7067;
  wire       [31:0]   _zz_7068;
  wire       [31:0]   _zz_7069;
  wire       [15:0]   _zz_7070;
  wire       [31:0]   _zz_7071;
  wire       [31:0]   _zz_7072;
  wire       [31:0]   _zz_7073;
  wire       [31:0]   _zz_7074;
  wire       [31:0]   _zz_7075;
  wire       [31:0]   _zz_7076;
  wire       [23:0]   _zz_7077;
  wire       [31:0]   _zz_7078;
  wire       [15:0]   _zz_7079;
  wire       [31:0]   _zz_7080;
  wire       [31:0]   _zz_7081;
  wire       [31:0]   _zz_7082;
  wire       [31:0]   _zz_7083;
  wire       [31:0]   _zz_7084;
  wire       [23:0]   _zz_7085;
  wire       [31:0]   _zz_7086;
  wire       [15:0]   _zz_7087;
  wire       [31:0]   _zz_7088;
  wire       [31:0]   _zz_7089;
  wire       [31:0]   _zz_7090;
  wire       [31:0]   _zz_7091;
  wire       [31:0]   _zz_7092;
  wire       [23:0]   _zz_7093;
  wire       [31:0]   _zz_7094;
  wire       [15:0]   _zz_7095;
  wire       [31:0]   _zz_7096;
  wire       [31:0]   _zz_7097;
  wire       [31:0]   _zz_7098;
  wire       [31:0]   _zz_7099;
  wire       [31:0]   _zz_7100;
  wire       [23:0]   _zz_7101;
  wire       [31:0]   _zz_7102;
  wire       [15:0]   _zz_7103;
  wire       [15:0]   _zz_7104;
  wire       [31:0]   _zz_7105;
  wire       [31:0]   _zz_7106;
  wire       [15:0]   _zz_7107;
  wire       [31:0]   _zz_7108;
  wire       [31:0]   _zz_7109;
  wire       [31:0]   _zz_7110;
  wire       [15:0]   _zz_7111;
  wire       [31:0]   _zz_7112;
  wire       [31:0]   _zz_7113;
  wire       [31:0]   _zz_7114;
  wire       [31:0]   _zz_7115;
  wire       [31:0]   _zz_7116;
  wire       [31:0]   _zz_7117;
  wire       [23:0]   _zz_7118;
  wire       [31:0]   _zz_7119;
  wire       [15:0]   _zz_7120;
  wire       [31:0]   _zz_7121;
  wire       [31:0]   _zz_7122;
  wire       [31:0]   _zz_7123;
  wire       [31:0]   _zz_7124;
  wire       [31:0]   _zz_7125;
  wire       [23:0]   _zz_7126;
  wire       [31:0]   _zz_7127;
  wire       [15:0]   _zz_7128;
  wire       [31:0]   _zz_7129;
  wire       [31:0]   _zz_7130;
  wire       [31:0]   _zz_7131;
  wire       [31:0]   _zz_7132;
  wire       [31:0]   _zz_7133;
  wire       [23:0]   _zz_7134;
  wire       [31:0]   _zz_7135;
  wire       [15:0]   _zz_7136;
  wire       [31:0]   _zz_7137;
  wire       [31:0]   _zz_7138;
  wire       [31:0]   _zz_7139;
  wire       [31:0]   _zz_7140;
  wire       [31:0]   _zz_7141;
  wire       [23:0]   _zz_7142;
  wire       [31:0]   _zz_7143;
  wire       [15:0]   _zz_7144;
  wire       [15:0]   _zz_7145;
  wire       [31:0]   _zz_7146;
  wire       [31:0]   _zz_7147;
  wire       [15:0]   _zz_7148;
  wire       [31:0]   _zz_7149;
  wire       [31:0]   _zz_7150;
  wire       [31:0]   _zz_7151;
  wire       [15:0]   _zz_7152;
  wire       [31:0]   _zz_7153;
  wire       [31:0]   _zz_7154;
  wire       [31:0]   _zz_7155;
  wire       [31:0]   _zz_7156;
  wire       [31:0]   _zz_7157;
  wire       [31:0]   _zz_7158;
  wire       [23:0]   _zz_7159;
  wire       [31:0]   _zz_7160;
  wire       [15:0]   _zz_7161;
  wire       [31:0]   _zz_7162;
  wire       [31:0]   _zz_7163;
  wire       [31:0]   _zz_7164;
  wire       [31:0]   _zz_7165;
  wire       [31:0]   _zz_7166;
  wire       [23:0]   _zz_7167;
  wire       [31:0]   _zz_7168;
  wire       [15:0]   _zz_7169;
  wire       [31:0]   _zz_7170;
  wire       [31:0]   _zz_7171;
  wire       [31:0]   _zz_7172;
  wire       [31:0]   _zz_7173;
  wire       [31:0]   _zz_7174;
  wire       [23:0]   _zz_7175;
  wire       [31:0]   _zz_7176;
  wire       [15:0]   _zz_7177;
  wire       [31:0]   _zz_7178;
  wire       [31:0]   _zz_7179;
  wire       [31:0]   _zz_7180;
  wire       [31:0]   _zz_7181;
  wire       [31:0]   _zz_7182;
  wire       [23:0]   _zz_7183;
  wire       [31:0]   _zz_7184;
  wire       [15:0]   _zz_7185;
  wire       [15:0]   _zz_7186;
  wire       [31:0]   _zz_7187;
  wire       [31:0]   _zz_7188;
  wire       [15:0]   _zz_7189;
  wire       [31:0]   _zz_7190;
  wire       [31:0]   _zz_7191;
  wire       [31:0]   _zz_7192;
  wire       [15:0]   _zz_7193;
  wire       [31:0]   _zz_7194;
  wire       [31:0]   _zz_7195;
  wire       [31:0]   _zz_7196;
  wire       [31:0]   _zz_7197;
  wire       [31:0]   _zz_7198;
  wire       [31:0]   _zz_7199;
  wire       [23:0]   _zz_7200;
  wire       [31:0]   _zz_7201;
  wire       [15:0]   _zz_7202;
  wire       [31:0]   _zz_7203;
  wire       [31:0]   _zz_7204;
  wire       [31:0]   _zz_7205;
  wire       [31:0]   _zz_7206;
  wire       [31:0]   _zz_7207;
  wire       [23:0]   _zz_7208;
  wire       [31:0]   _zz_7209;
  wire       [15:0]   _zz_7210;
  wire       [31:0]   _zz_7211;
  wire       [31:0]   _zz_7212;
  wire       [31:0]   _zz_7213;
  wire       [31:0]   _zz_7214;
  wire       [31:0]   _zz_7215;
  wire       [23:0]   _zz_7216;
  wire       [31:0]   _zz_7217;
  wire       [15:0]   _zz_7218;
  wire       [31:0]   _zz_7219;
  wire       [31:0]   _zz_7220;
  wire       [31:0]   _zz_7221;
  wire       [31:0]   _zz_7222;
  wire       [31:0]   _zz_7223;
  wire       [23:0]   _zz_7224;
  wire       [31:0]   _zz_7225;
  wire       [15:0]   _zz_7226;
  wire       [15:0]   _zz_7227;
  wire       [31:0]   _zz_7228;
  wire       [31:0]   _zz_7229;
  wire       [15:0]   _zz_7230;
  wire       [31:0]   _zz_7231;
  wire       [31:0]   _zz_7232;
  wire       [31:0]   _zz_7233;
  wire       [15:0]   _zz_7234;
  wire       [31:0]   _zz_7235;
  wire       [31:0]   _zz_7236;
  wire       [31:0]   _zz_7237;
  wire       [31:0]   _zz_7238;
  wire       [31:0]   _zz_7239;
  wire       [31:0]   _zz_7240;
  wire       [23:0]   _zz_7241;
  wire       [31:0]   _zz_7242;
  wire       [15:0]   _zz_7243;
  wire       [31:0]   _zz_7244;
  wire       [31:0]   _zz_7245;
  wire       [31:0]   _zz_7246;
  wire       [31:0]   _zz_7247;
  wire       [31:0]   _zz_7248;
  wire       [23:0]   _zz_7249;
  wire       [31:0]   _zz_7250;
  wire       [15:0]   _zz_7251;
  wire       [31:0]   _zz_7252;
  wire       [31:0]   _zz_7253;
  wire       [31:0]   _zz_7254;
  wire       [31:0]   _zz_7255;
  wire       [31:0]   _zz_7256;
  wire       [23:0]   _zz_7257;
  wire       [31:0]   _zz_7258;
  wire       [15:0]   _zz_7259;
  wire       [31:0]   _zz_7260;
  wire       [31:0]   _zz_7261;
  wire       [31:0]   _zz_7262;
  wire       [31:0]   _zz_7263;
  wire       [31:0]   _zz_7264;
  wire       [23:0]   _zz_7265;
  wire       [31:0]   _zz_7266;
  wire       [15:0]   _zz_7267;
  wire       [15:0]   _zz_7268;
  wire       [31:0]   _zz_7269;
  wire       [31:0]   _zz_7270;
  wire       [15:0]   _zz_7271;
  wire       [31:0]   _zz_7272;
  wire       [31:0]   _zz_7273;
  wire       [31:0]   _zz_7274;
  wire       [15:0]   _zz_7275;
  wire       [31:0]   _zz_7276;
  wire       [31:0]   _zz_7277;
  wire       [31:0]   _zz_7278;
  wire       [31:0]   _zz_7279;
  wire       [31:0]   _zz_7280;
  wire       [31:0]   _zz_7281;
  wire       [23:0]   _zz_7282;
  wire       [31:0]   _zz_7283;
  wire       [15:0]   _zz_7284;
  wire       [31:0]   _zz_7285;
  wire       [31:0]   _zz_7286;
  wire       [31:0]   _zz_7287;
  wire       [31:0]   _zz_7288;
  wire       [31:0]   _zz_7289;
  wire       [23:0]   _zz_7290;
  wire       [31:0]   _zz_7291;
  wire       [15:0]   _zz_7292;
  wire       [31:0]   _zz_7293;
  wire       [31:0]   _zz_7294;
  wire       [31:0]   _zz_7295;
  wire       [31:0]   _zz_7296;
  wire       [31:0]   _zz_7297;
  wire       [23:0]   _zz_7298;
  wire       [31:0]   _zz_7299;
  wire       [15:0]   _zz_7300;
  wire       [31:0]   _zz_7301;
  wire       [31:0]   _zz_7302;
  wire       [31:0]   _zz_7303;
  wire       [31:0]   _zz_7304;
  wire       [31:0]   _zz_7305;
  wire       [23:0]   _zz_7306;
  wire       [31:0]   _zz_7307;
  wire       [15:0]   _zz_7308;
  wire       [15:0]   _zz_7309;
  wire       [31:0]   _zz_7310;
  wire       [31:0]   _zz_7311;
  wire       [15:0]   _zz_7312;
  wire       [31:0]   _zz_7313;
  wire       [31:0]   _zz_7314;
  wire       [31:0]   _zz_7315;
  wire       [15:0]   _zz_7316;
  wire       [31:0]   _zz_7317;
  wire       [31:0]   _zz_7318;
  wire       [31:0]   _zz_7319;
  wire       [31:0]   _zz_7320;
  wire       [31:0]   _zz_7321;
  wire       [31:0]   _zz_7322;
  wire       [23:0]   _zz_7323;
  wire       [31:0]   _zz_7324;
  wire       [15:0]   _zz_7325;
  wire       [31:0]   _zz_7326;
  wire       [31:0]   _zz_7327;
  wire       [31:0]   _zz_7328;
  wire       [31:0]   _zz_7329;
  wire       [31:0]   _zz_7330;
  wire       [23:0]   _zz_7331;
  wire       [31:0]   _zz_7332;
  wire       [15:0]   _zz_7333;
  wire       [31:0]   _zz_7334;
  wire       [31:0]   _zz_7335;
  wire       [31:0]   _zz_7336;
  wire       [31:0]   _zz_7337;
  wire       [31:0]   _zz_7338;
  wire       [23:0]   _zz_7339;
  wire       [31:0]   _zz_7340;
  wire       [15:0]   _zz_7341;
  wire       [31:0]   _zz_7342;
  wire       [31:0]   _zz_7343;
  wire       [31:0]   _zz_7344;
  wire       [31:0]   _zz_7345;
  wire       [31:0]   _zz_7346;
  wire       [23:0]   _zz_7347;
  wire       [31:0]   _zz_7348;
  wire       [15:0]   _zz_7349;
  wire       [15:0]   _zz_7350;
  wire       [31:0]   _zz_7351;
  wire       [31:0]   _zz_7352;
  wire       [15:0]   _zz_7353;
  wire       [31:0]   _zz_7354;
  wire       [31:0]   _zz_7355;
  wire       [31:0]   _zz_7356;
  wire       [15:0]   _zz_7357;
  wire       [31:0]   _zz_7358;
  wire       [31:0]   _zz_7359;
  wire       [31:0]   _zz_7360;
  wire       [31:0]   _zz_7361;
  wire       [31:0]   _zz_7362;
  wire       [31:0]   _zz_7363;
  wire       [23:0]   _zz_7364;
  wire       [31:0]   _zz_7365;
  wire       [15:0]   _zz_7366;
  wire       [31:0]   _zz_7367;
  wire       [31:0]   _zz_7368;
  wire       [31:0]   _zz_7369;
  wire       [31:0]   _zz_7370;
  wire       [31:0]   _zz_7371;
  wire       [23:0]   _zz_7372;
  wire       [31:0]   _zz_7373;
  wire       [15:0]   _zz_7374;
  wire       [31:0]   _zz_7375;
  wire       [31:0]   _zz_7376;
  wire       [31:0]   _zz_7377;
  wire       [31:0]   _zz_7378;
  wire       [31:0]   _zz_7379;
  wire       [23:0]   _zz_7380;
  wire       [31:0]   _zz_7381;
  wire       [15:0]   _zz_7382;
  wire       [31:0]   _zz_7383;
  wire       [31:0]   _zz_7384;
  wire       [31:0]   _zz_7385;
  wire       [31:0]   _zz_7386;
  wire       [31:0]   _zz_7387;
  wire       [23:0]   _zz_7388;
  wire       [31:0]   _zz_7389;
  wire       [15:0]   _zz_7390;
  wire       [15:0]   _zz_7391;
  wire       [31:0]   _zz_7392;
  wire       [31:0]   _zz_7393;
  wire       [15:0]   _zz_7394;
  wire       [31:0]   _zz_7395;
  wire       [31:0]   _zz_7396;
  wire       [31:0]   _zz_7397;
  wire       [15:0]   _zz_7398;
  wire       [31:0]   _zz_7399;
  wire       [31:0]   _zz_7400;
  wire       [31:0]   _zz_7401;
  wire       [31:0]   _zz_7402;
  wire       [31:0]   _zz_7403;
  wire       [31:0]   _zz_7404;
  wire       [23:0]   _zz_7405;
  wire       [31:0]   _zz_7406;
  wire       [15:0]   _zz_7407;
  wire       [31:0]   _zz_7408;
  wire       [31:0]   _zz_7409;
  wire       [31:0]   _zz_7410;
  wire       [31:0]   _zz_7411;
  wire       [31:0]   _zz_7412;
  wire       [23:0]   _zz_7413;
  wire       [31:0]   _zz_7414;
  wire       [15:0]   _zz_7415;
  wire       [31:0]   _zz_7416;
  wire       [31:0]   _zz_7417;
  wire       [31:0]   _zz_7418;
  wire       [31:0]   _zz_7419;
  wire       [31:0]   _zz_7420;
  wire       [23:0]   _zz_7421;
  wire       [31:0]   _zz_7422;
  wire       [15:0]   _zz_7423;
  wire       [31:0]   _zz_7424;
  wire       [31:0]   _zz_7425;
  wire       [31:0]   _zz_7426;
  wire       [31:0]   _zz_7427;
  wire       [31:0]   _zz_7428;
  wire       [23:0]   _zz_7429;
  wire       [31:0]   _zz_7430;
  wire       [15:0]   _zz_7431;
  wire       [15:0]   _zz_7432;
  wire       [31:0]   _zz_7433;
  wire       [31:0]   _zz_7434;
  wire       [15:0]   _zz_7435;
  wire       [31:0]   _zz_7436;
  wire       [31:0]   _zz_7437;
  wire       [31:0]   _zz_7438;
  wire       [15:0]   _zz_7439;
  wire       [31:0]   _zz_7440;
  wire       [31:0]   _zz_7441;
  wire       [31:0]   _zz_7442;
  wire       [31:0]   _zz_7443;
  wire       [31:0]   _zz_7444;
  wire       [31:0]   _zz_7445;
  wire       [23:0]   _zz_7446;
  wire       [31:0]   _zz_7447;
  wire       [15:0]   _zz_7448;
  wire       [31:0]   _zz_7449;
  wire       [31:0]   _zz_7450;
  wire       [31:0]   _zz_7451;
  wire       [31:0]   _zz_7452;
  wire       [31:0]   _zz_7453;
  wire       [23:0]   _zz_7454;
  wire       [31:0]   _zz_7455;
  wire       [15:0]   _zz_7456;
  wire       [31:0]   _zz_7457;
  wire       [31:0]   _zz_7458;
  wire       [31:0]   _zz_7459;
  wire       [31:0]   _zz_7460;
  wire       [31:0]   _zz_7461;
  wire       [23:0]   _zz_7462;
  wire       [31:0]   _zz_7463;
  wire       [15:0]   _zz_7464;
  wire       [31:0]   _zz_7465;
  wire       [31:0]   _zz_7466;
  wire       [31:0]   _zz_7467;
  wire       [31:0]   _zz_7468;
  wire       [31:0]   _zz_7469;
  wire       [23:0]   _zz_7470;
  wire       [31:0]   _zz_7471;
  wire       [15:0]   _zz_7472;
  wire       [15:0]   _zz_7473;
  wire       [31:0]   _zz_7474;
  wire       [31:0]   _zz_7475;
  wire       [15:0]   _zz_7476;
  wire       [31:0]   _zz_7477;
  wire       [31:0]   _zz_7478;
  wire       [31:0]   _zz_7479;
  wire       [15:0]   _zz_7480;
  wire       [31:0]   _zz_7481;
  wire       [31:0]   _zz_7482;
  wire       [31:0]   _zz_7483;
  wire       [31:0]   _zz_7484;
  wire       [31:0]   _zz_7485;
  wire       [31:0]   _zz_7486;
  wire       [23:0]   _zz_7487;
  wire       [31:0]   _zz_7488;
  wire       [15:0]   _zz_7489;
  wire       [31:0]   _zz_7490;
  wire       [31:0]   _zz_7491;
  wire       [31:0]   _zz_7492;
  wire       [31:0]   _zz_7493;
  wire       [31:0]   _zz_7494;
  wire       [23:0]   _zz_7495;
  wire       [31:0]   _zz_7496;
  wire       [15:0]   _zz_7497;
  wire       [31:0]   _zz_7498;
  wire       [31:0]   _zz_7499;
  wire       [31:0]   _zz_7500;
  wire       [31:0]   _zz_7501;
  wire       [31:0]   _zz_7502;
  wire       [23:0]   _zz_7503;
  wire       [31:0]   _zz_7504;
  wire       [15:0]   _zz_7505;
  wire       [31:0]   _zz_7506;
  wire       [31:0]   _zz_7507;
  wire       [31:0]   _zz_7508;
  wire       [31:0]   _zz_7509;
  wire       [31:0]   _zz_7510;
  wire       [23:0]   _zz_7511;
  wire       [31:0]   _zz_7512;
  wire       [15:0]   _zz_7513;
  wire       [15:0]   _zz_7514;
  wire       [31:0]   _zz_7515;
  wire       [31:0]   _zz_7516;
  wire       [15:0]   _zz_7517;
  wire       [31:0]   _zz_7518;
  wire       [31:0]   _zz_7519;
  wire       [31:0]   _zz_7520;
  wire       [15:0]   _zz_7521;
  wire       [31:0]   _zz_7522;
  wire       [31:0]   _zz_7523;
  wire       [31:0]   _zz_7524;
  wire       [31:0]   _zz_7525;
  wire       [31:0]   _zz_7526;
  wire       [31:0]   _zz_7527;
  wire       [23:0]   _zz_7528;
  wire       [31:0]   _zz_7529;
  wire       [15:0]   _zz_7530;
  wire       [31:0]   _zz_7531;
  wire       [31:0]   _zz_7532;
  wire       [31:0]   _zz_7533;
  wire       [31:0]   _zz_7534;
  wire       [31:0]   _zz_7535;
  wire       [23:0]   _zz_7536;
  wire       [31:0]   _zz_7537;
  wire       [15:0]   _zz_7538;
  wire       [31:0]   _zz_7539;
  wire       [31:0]   _zz_7540;
  wire       [31:0]   _zz_7541;
  wire       [31:0]   _zz_7542;
  wire       [31:0]   _zz_7543;
  wire       [23:0]   _zz_7544;
  wire       [31:0]   _zz_7545;
  wire       [15:0]   _zz_7546;
  wire       [31:0]   _zz_7547;
  wire       [31:0]   _zz_7548;
  wire       [31:0]   _zz_7549;
  wire       [31:0]   _zz_7550;
  wire       [31:0]   _zz_7551;
  wire       [23:0]   _zz_7552;
  wire       [31:0]   _zz_7553;
  wire       [15:0]   _zz_7554;
  wire       [15:0]   _zz_7555;
  wire       [31:0]   _zz_7556;
  wire       [31:0]   _zz_7557;
  wire       [15:0]   _zz_7558;
  wire       [31:0]   _zz_7559;
  wire       [31:0]   _zz_7560;
  wire       [31:0]   _zz_7561;
  wire       [15:0]   _zz_7562;
  wire       [31:0]   _zz_7563;
  wire       [31:0]   _zz_7564;
  wire       [31:0]   _zz_7565;
  wire       [31:0]   _zz_7566;
  wire       [31:0]   _zz_7567;
  wire       [31:0]   _zz_7568;
  wire       [23:0]   _zz_7569;
  wire       [31:0]   _zz_7570;
  wire       [15:0]   _zz_7571;
  wire       [31:0]   _zz_7572;
  wire       [31:0]   _zz_7573;
  wire       [31:0]   _zz_7574;
  wire       [31:0]   _zz_7575;
  wire       [31:0]   _zz_7576;
  wire       [23:0]   _zz_7577;
  wire       [31:0]   _zz_7578;
  wire       [15:0]   _zz_7579;
  wire       [31:0]   _zz_7580;
  wire       [31:0]   _zz_7581;
  wire       [31:0]   _zz_7582;
  wire       [31:0]   _zz_7583;
  wire       [31:0]   _zz_7584;
  wire       [23:0]   _zz_7585;
  wire       [31:0]   _zz_7586;
  wire       [15:0]   _zz_7587;
  wire       [31:0]   _zz_7588;
  wire       [31:0]   _zz_7589;
  wire       [31:0]   _zz_7590;
  wire       [31:0]   _zz_7591;
  wire       [31:0]   _zz_7592;
  wire       [23:0]   _zz_7593;
  wire       [31:0]   _zz_7594;
  wire       [15:0]   _zz_7595;
  wire       [15:0]   _zz_7596;
  wire       [31:0]   _zz_7597;
  wire       [31:0]   _zz_7598;
  wire       [15:0]   _zz_7599;
  wire       [31:0]   _zz_7600;
  wire       [31:0]   _zz_7601;
  wire       [31:0]   _zz_7602;
  wire       [15:0]   _zz_7603;
  wire       [31:0]   _zz_7604;
  wire       [31:0]   _zz_7605;
  wire       [31:0]   _zz_7606;
  wire       [31:0]   _zz_7607;
  wire       [31:0]   _zz_7608;
  wire       [31:0]   _zz_7609;
  wire       [23:0]   _zz_7610;
  wire       [31:0]   _zz_7611;
  wire       [15:0]   _zz_7612;
  wire       [31:0]   _zz_7613;
  wire       [31:0]   _zz_7614;
  wire       [31:0]   _zz_7615;
  wire       [31:0]   _zz_7616;
  wire       [31:0]   _zz_7617;
  wire       [23:0]   _zz_7618;
  wire       [31:0]   _zz_7619;
  wire       [15:0]   _zz_7620;
  wire       [31:0]   _zz_7621;
  wire       [31:0]   _zz_7622;
  wire       [31:0]   _zz_7623;
  wire       [31:0]   _zz_7624;
  wire       [31:0]   _zz_7625;
  wire       [23:0]   _zz_7626;
  wire       [31:0]   _zz_7627;
  wire       [15:0]   _zz_7628;
  wire       [31:0]   _zz_7629;
  wire       [31:0]   _zz_7630;
  wire       [31:0]   _zz_7631;
  wire       [31:0]   _zz_7632;
  wire       [31:0]   _zz_7633;
  wire       [23:0]   _zz_7634;
  wire       [31:0]   _zz_7635;
  wire       [15:0]   _zz_7636;
  wire       [15:0]   _zz_7637;
  wire       [31:0]   _zz_7638;
  wire       [31:0]   _zz_7639;
  wire       [15:0]   _zz_7640;
  wire       [31:0]   _zz_7641;
  wire       [31:0]   _zz_7642;
  wire       [31:0]   _zz_7643;
  wire       [15:0]   _zz_7644;
  wire       [31:0]   _zz_7645;
  wire       [31:0]   _zz_7646;
  wire       [31:0]   _zz_7647;
  wire       [31:0]   _zz_7648;
  wire       [31:0]   _zz_7649;
  wire       [31:0]   _zz_7650;
  wire       [23:0]   _zz_7651;
  wire       [31:0]   _zz_7652;
  wire       [15:0]   _zz_7653;
  wire       [31:0]   _zz_7654;
  wire       [31:0]   _zz_7655;
  wire       [31:0]   _zz_7656;
  wire       [31:0]   _zz_7657;
  wire       [31:0]   _zz_7658;
  wire       [23:0]   _zz_7659;
  wire       [31:0]   _zz_7660;
  wire       [15:0]   _zz_7661;
  wire       [31:0]   _zz_7662;
  wire       [31:0]   _zz_7663;
  wire       [31:0]   _zz_7664;
  wire       [31:0]   _zz_7665;
  wire       [31:0]   _zz_7666;
  wire       [23:0]   _zz_7667;
  wire       [31:0]   _zz_7668;
  wire       [15:0]   _zz_7669;
  wire       [31:0]   _zz_7670;
  wire       [31:0]   _zz_7671;
  wire       [31:0]   _zz_7672;
  wire       [31:0]   _zz_7673;
  wire       [31:0]   _zz_7674;
  wire       [23:0]   _zz_7675;
  wire       [31:0]   _zz_7676;
  wire       [15:0]   _zz_7677;
  wire       [15:0]   _zz_7678;
  wire       [31:0]   _zz_7679;
  wire       [31:0]   _zz_7680;
  wire       [15:0]   _zz_7681;
  wire       [31:0]   _zz_7682;
  wire       [31:0]   _zz_7683;
  wire       [31:0]   _zz_7684;
  wire       [15:0]   _zz_7685;
  wire       [31:0]   _zz_7686;
  wire       [31:0]   _zz_7687;
  wire       [31:0]   _zz_7688;
  wire       [31:0]   _zz_7689;
  wire       [31:0]   _zz_7690;
  wire       [31:0]   _zz_7691;
  wire       [23:0]   _zz_7692;
  wire       [31:0]   _zz_7693;
  wire       [15:0]   _zz_7694;
  wire       [31:0]   _zz_7695;
  wire       [31:0]   _zz_7696;
  wire       [31:0]   _zz_7697;
  wire       [31:0]   _zz_7698;
  wire       [31:0]   _zz_7699;
  wire       [23:0]   _zz_7700;
  wire       [31:0]   _zz_7701;
  wire       [15:0]   _zz_7702;
  wire       [31:0]   _zz_7703;
  wire       [31:0]   _zz_7704;
  wire       [31:0]   _zz_7705;
  wire       [31:0]   _zz_7706;
  wire       [31:0]   _zz_7707;
  wire       [23:0]   _zz_7708;
  wire       [31:0]   _zz_7709;
  wire       [15:0]   _zz_7710;
  wire       [31:0]   _zz_7711;
  wire       [31:0]   _zz_7712;
  wire       [31:0]   _zz_7713;
  wire       [31:0]   _zz_7714;
  wire       [31:0]   _zz_7715;
  wire       [23:0]   _zz_7716;
  wire       [31:0]   _zz_7717;
  wire       [15:0]   _zz_7718;
  wire       [15:0]   _zz_7719;
  wire       [31:0]   _zz_7720;
  wire       [31:0]   _zz_7721;
  wire       [15:0]   _zz_7722;
  wire       [31:0]   _zz_7723;
  wire       [31:0]   _zz_7724;
  wire       [31:0]   _zz_7725;
  wire       [15:0]   _zz_7726;
  wire       [31:0]   _zz_7727;
  wire       [31:0]   _zz_7728;
  wire       [31:0]   _zz_7729;
  wire       [31:0]   _zz_7730;
  wire       [31:0]   _zz_7731;
  wire       [31:0]   _zz_7732;
  wire       [23:0]   _zz_7733;
  wire       [31:0]   _zz_7734;
  wire       [15:0]   _zz_7735;
  wire       [31:0]   _zz_7736;
  wire       [31:0]   _zz_7737;
  wire       [31:0]   _zz_7738;
  wire       [31:0]   _zz_7739;
  wire       [31:0]   _zz_7740;
  wire       [23:0]   _zz_7741;
  wire       [31:0]   _zz_7742;
  wire       [15:0]   _zz_7743;
  wire       [31:0]   _zz_7744;
  wire       [31:0]   _zz_7745;
  wire       [31:0]   _zz_7746;
  wire       [31:0]   _zz_7747;
  wire       [31:0]   _zz_7748;
  wire       [23:0]   _zz_7749;
  wire       [31:0]   _zz_7750;
  wire       [15:0]   _zz_7751;
  wire       [31:0]   _zz_7752;
  wire       [31:0]   _zz_7753;
  wire       [31:0]   _zz_7754;
  wire       [31:0]   _zz_7755;
  wire       [31:0]   _zz_7756;
  wire       [23:0]   _zz_7757;
  wire       [31:0]   _zz_7758;
  wire       [15:0]   _zz_7759;
  wire       [15:0]   _zz_7760;
  wire       [31:0]   _zz_7761;
  wire       [31:0]   _zz_7762;
  wire       [15:0]   _zz_7763;
  wire       [31:0]   _zz_7764;
  wire       [31:0]   _zz_7765;
  wire       [31:0]   _zz_7766;
  wire       [15:0]   _zz_7767;
  wire       [31:0]   _zz_7768;
  wire       [31:0]   _zz_7769;
  wire       [31:0]   _zz_7770;
  wire       [31:0]   _zz_7771;
  wire       [31:0]   _zz_7772;
  wire       [31:0]   _zz_7773;
  wire       [23:0]   _zz_7774;
  wire       [31:0]   _zz_7775;
  wire       [15:0]   _zz_7776;
  wire       [31:0]   _zz_7777;
  wire       [31:0]   _zz_7778;
  wire       [31:0]   _zz_7779;
  wire       [31:0]   _zz_7780;
  wire       [31:0]   _zz_7781;
  wire       [23:0]   _zz_7782;
  wire       [31:0]   _zz_7783;
  wire       [15:0]   _zz_7784;
  wire       [31:0]   _zz_7785;
  wire       [31:0]   _zz_7786;
  wire       [31:0]   _zz_7787;
  wire       [31:0]   _zz_7788;
  wire       [31:0]   _zz_7789;
  wire       [23:0]   _zz_7790;
  wire       [31:0]   _zz_7791;
  wire       [15:0]   _zz_7792;
  wire       [31:0]   _zz_7793;
  wire       [31:0]   _zz_7794;
  wire       [31:0]   _zz_7795;
  wire       [31:0]   _zz_7796;
  wire       [31:0]   _zz_7797;
  wire       [23:0]   _zz_7798;
  wire       [31:0]   _zz_7799;
  wire       [15:0]   _zz_7800;
  wire       [15:0]   _zz_7801;
  wire       [31:0]   _zz_7802;
  wire       [31:0]   _zz_7803;
  wire       [15:0]   _zz_7804;
  wire       [31:0]   _zz_7805;
  wire       [31:0]   _zz_7806;
  wire       [31:0]   _zz_7807;
  wire       [15:0]   _zz_7808;
  wire       [31:0]   _zz_7809;
  wire       [31:0]   _zz_7810;
  wire       [31:0]   _zz_7811;
  wire       [31:0]   _zz_7812;
  wire       [31:0]   _zz_7813;
  wire       [31:0]   _zz_7814;
  wire       [23:0]   _zz_7815;
  wire       [31:0]   _zz_7816;
  wire       [15:0]   _zz_7817;
  wire       [31:0]   _zz_7818;
  wire       [31:0]   _zz_7819;
  wire       [31:0]   _zz_7820;
  wire       [31:0]   _zz_7821;
  wire       [31:0]   _zz_7822;
  wire       [23:0]   _zz_7823;
  wire       [31:0]   _zz_7824;
  wire       [15:0]   _zz_7825;
  wire       [31:0]   _zz_7826;
  wire       [31:0]   _zz_7827;
  wire       [31:0]   _zz_7828;
  wire       [31:0]   _zz_7829;
  wire       [31:0]   _zz_7830;
  wire       [23:0]   _zz_7831;
  wire       [31:0]   _zz_7832;
  wire       [15:0]   _zz_7833;
  wire       [31:0]   _zz_7834;
  wire       [31:0]   _zz_7835;
  wire       [31:0]   _zz_7836;
  wire       [31:0]   _zz_7837;
  wire       [31:0]   _zz_7838;
  wire       [23:0]   _zz_7839;
  wire       [31:0]   _zz_7840;
  wire       [15:0]   _zz_7841;
  wire       [15:0]   _zz_7842;
  wire       [31:0]   _zz_7843;
  wire       [31:0]   _zz_7844;
  wire       [15:0]   _zz_7845;
  wire       [31:0]   _zz_7846;
  wire       [31:0]   _zz_7847;
  wire       [31:0]   _zz_7848;
  wire       [15:0]   _zz_7849;
  wire       [31:0]   _zz_7850;
  wire       [31:0]   _zz_7851;
  wire       [31:0]   _zz_7852;
  wire       [31:0]   _zz_7853;
  wire       [31:0]   _zz_7854;
  wire       [31:0]   _zz_7855;
  wire       [23:0]   _zz_7856;
  wire       [31:0]   _zz_7857;
  wire       [15:0]   _zz_7858;
  wire       [31:0]   _zz_7859;
  wire       [31:0]   _zz_7860;
  wire       [31:0]   _zz_7861;
  wire       [31:0]   _zz_7862;
  wire       [31:0]   _zz_7863;
  wire       [23:0]   _zz_7864;
  wire       [31:0]   _zz_7865;
  wire       [15:0]   _zz_7866;
  wire       [31:0]   _zz_7867;
  wire       [31:0]   _zz_7868;
  wire       [31:0]   _zz_7869;
  wire       [31:0]   _zz_7870;
  wire       [31:0]   _zz_7871;
  wire       [23:0]   _zz_7872;
  wire       [31:0]   _zz_7873;
  wire       [15:0]   _zz_7874;
  wire       [31:0]   _zz_7875;
  wire       [31:0]   _zz_7876;
  wire       [31:0]   _zz_7877;
  wire       [31:0]   _zz_7878;
  wire       [31:0]   _zz_7879;
  wire       [23:0]   _zz_7880;
  wire       [31:0]   _zz_7881;
  wire       [15:0]   _zz_7882;
  wire       [15:0]   _zz_7883;
  wire       [31:0]   _zz_7884;
  wire       [31:0]   _zz_7885;
  wire       [15:0]   _zz_7886;
  wire       [31:0]   _zz_7887;
  wire       [31:0]   _zz_7888;
  wire       [31:0]   _zz_7889;
  wire       [15:0]   _zz_7890;
  wire       [31:0]   _zz_7891;
  wire       [31:0]   _zz_7892;
  wire       [31:0]   _zz_7893;
  wire       [31:0]   _zz_7894;
  wire       [31:0]   _zz_7895;
  wire       [31:0]   _zz_7896;
  wire       [23:0]   _zz_7897;
  wire       [31:0]   _zz_7898;
  wire       [15:0]   _zz_7899;
  wire       [31:0]   _zz_7900;
  wire       [31:0]   _zz_7901;
  wire       [31:0]   _zz_7902;
  wire       [31:0]   _zz_7903;
  wire       [31:0]   _zz_7904;
  wire       [23:0]   _zz_7905;
  wire       [31:0]   _zz_7906;
  wire       [15:0]   _zz_7907;
  wire       [31:0]   _zz_7908;
  wire       [31:0]   _zz_7909;
  wire       [31:0]   _zz_7910;
  wire       [31:0]   _zz_7911;
  wire       [31:0]   _zz_7912;
  wire       [23:0]   _zz_7913;
  wire       [31:0]   _zz_7914;
  wire       [15:0]   _zz_7915;
  wire       [31:0]   _zz_7916;
  wire       [31:0]   _zz_7917;
  wire       [31:0]   _zz_7918;
  wire       [31:0]   _zz_7919;
  wire       [31:0]   _zz_7920;
  wire       [23:0]   _zz_7921;
  wire       [31:0]   _zz_7922;
  wire       [15:0]   _zz_7923;
  wire       [15:0]   _zz_7924;
  wire       [31:0]   _zz_7925;
  wire       [31:0]   _zz_7926;
  wire       [15:0]   _zz_7927;
  wire       [31:0]   _zz_7928;
  wire       [31:0]   _zz_7929;
  wire       [31:0]   _zz_7930;
  wire       [15:0]   _zz_7931;
  wire       [31:0]   _zz_7932;
  wire       [31:0]   _zz_7933;
  wire       [31:0]   _zz_7934;
  wire       [31:0]   _zz_7935;
  wire       [31:0]   _zz_7936;
  wire       [31:0]   _zz_7937;
  wire       [23:0]   _zz_7938;
  wire       [31:0]   _zz_7939;
  wire       [15:0]   _zz_7940;
  wire       [31:0]   _zz_7941;
  wire       [31:0]   _zz_7942;
  wire       [31:0]   _zz_7943;
  wire       [31:0]   _zz_7944;
  wire       [31:0]   _zz_7945;
  wire       [23:0]   _zz_7946;
  wire       [31:0]   _zz_7947;
  wire       [15:0]   _zz_7948;
  wire       [31:0]   _zz_7949;
  wire       [31:0]   _zz_7950;
  wire       [31:0]   _zz_7951;
  wire       [31:0]   _zz_7952;
  wire       [31:0]   _zz_7953;
  wire       [23:0]   _zz_7954;
  wire       [31:0]   _zz_7955;
  wire       [15:0]   _zz_7956;
  wire       [31:0]   _zz_7957;
  wire       [31:0]   _zz_7958;
  wire       [31:0]   _zz_7959;
  wire       [31:0]   _zz_7960;
  wire       [31:0]   _zz_7961;
  wire       [23:0]   _zz_7962;
  wire       [31:0]   _zz_7963;
  wire       [15:0]   _zz_7964;
  wire       [15:0]   _zz_7965;
  wire       [31:0]   _zz_7966;
  wire       [31:0]   _zz_7967;
  wire       [15:0]   _zz_7968;
  wire       [31:0]   _zz_7969;
  wire       [31:0]   _zz_7970;
  wire       [31:0]   _zz_7971;
  wire       [15:0]   _zz_7972;
  wire       [31:0]   _zz_7973;
  wire       [31:0]   _zz_7974;
  wire       [31:0]   _zz_7975;
  wire       [31:0]   _zz_7976;
  wire       [31:0]   _zz_7977;
  wire       [31:0]   _zz_7978;
  wire       [23:0]   _zz_7979;
  wire       [31:0]   _zz_7980;
  wire       [15:0]   _zz_7981;
  wire       [31:0]   _zz_7982;
  wire       [31:0]   _zz_7983;
  wire       [31:0]   _zz_7984;
  wire       [31:0]   _zz_7985;
  wire       [31:0]   _zz_7986;
  wire       [23:0]   _zz_7987;
  wire       [31:0]   _zz_7988;
  wire       [15:0]   _zz_7989;
  wire       [31:0]   _zz_7990;
  wire       [31:0]   _zz_7991;
  wire       [31:0]   _zz_7992;
  wire       [31:0]   _zz_7993;
  wire       [31:0]   _zz_7994;
  wire       [23:0]   _zz_7995;
  wire       [31:0]   _zz_7996;
  wire       [15:0]   _zz_7997;
  wire       [31:0]   _zz_7998;
  wire       [31:0]   _zz_7999;
  wire       [31:0]   _zz_8000;
  wire       [31:0]   _zz_8001;
  wire       [31:0]   _zz_8002;
  wire       [23:0]   _zz_8003;
  wire       [31:0]   _zz_8004;
  wire       [15:0]   _zz_8005;
  wire       [15:0]   _zz_8006;
  wire       [31:0]   _zz_8007;
  wire       [31:0]   _zz_8008;
  wire       [15:0]   _zz_8009;
  wire       [31:0]   _zz_8010;
  wire       [31:0]   _zz_8011;
  wire       [31:0]   _zz_8012;
  wire       [15:0]   _zz_8013;
  wire       [31:0]   _zz_8014;
  wire       [31:0]   _zz_8015;
  wire       [31:0]   _zz_8016;
  wire       [31:0]   _zz_8017;
  wire       [31:0]   _zz_8018;
  wire       [31:0]   _zz_8019;
  wire       [23:0]   _zz_8020;
  wire       [31:0]   _zz_8021;
  wire       [15:0]   _zz_8022;
  wire       [31:0]   _zz_8023;
  wire       [31:0]   _zz_8024;
  wire       [31:0]   _zz_8025;
  wire       [31:0]   _zz_8026;
  wire       [31:0]   _zz_8027;
  wire       [23:0]   _zz_8028;
  wire       [31:0]   _zz_8029;
  wire       [15:0]   _zz_8030;
  wire       [31:0]   _zz_8031;
  wire       [31:0]   _zz_8032;
  wire       [31:0]   _zz_8033;
  wire       [31:0]   _zz_8034;
  wire       [31:0]   _zz_8035;
  wire       [23:0]   _zz_8036;
  wire       [31:0]   _zz_8037;
  wire       [15:0]   _zz_8038;
  wire       [31:0]   _zz_8039;
  wire       [31:0]   _zz_8040;
  wire       [31:0]   _zz_8041;
  wire       [31:0]   _zz_8042;
  wire       [31:0]   _zz_8043;
  wire       [23:0]   _zz_8044;
  wire       [31:0]   _zz_8045;
  wire       [15:0]   _zz_8046;
  wire       [15:0]   _zz_8047;
  wire       [31:0]   _zz_8048;
  wire       [31:0]   _zz_8049;
  wire       [15:0]   _zz_8050;
  wire       [31:0]   _zz_8051;
  wire       [31:0]   _zz_8052;
  wire       [31:0]   _zz_8053;
  wire       [15:0]   _zz_8054;
  wire       [31:0]   _zz_8055;
  wire       [31:0]   _zz_8056;
  wire       [31:0]   _zz_8057;
  wire       [31:0]   _zz_8058;
  wire       [31:0]   _zz_8059;
  wire       [31:0]   _zz_8060;
  wire       [23:0]   _zz_8061;
  wire       [31:0]   _zz_8062;
  wire       [15:0]   _zz_8063;
  wire       [31:0]   _zz_8064;
  wire       [31:0]   _zz_8065;
  wire       [31:0]   _zz_8066;
  wire       [31:0]   _zz_8067;
  wire       [31:0]   _zz_8068;
  wire       [23:0]   _zz_8069;
  wire       [31:0]   _zz_8070;
  wire       [15:0]   _zz_8071;
  wire       [31:0]   _zz_8072;
  wire       [31:0]   _zz_8073;
  wire       [31:0]   _zz_8074;
  wire       [31:0]   _zz_8075;
  wire       [31:0]   _zz_8076;
  wire       [23:0]   _zz_8077;
  wire       [31:0]   _zz_8078;
  wire       [15:0]   _zz_8079;
  wire       [31:0]   _zz_8080;
  wire       [31:0]   _zz_8081;
  wire       [31:0]   _zz_8082;
  wire       [31:0]   _zz_8083;
  wire       [31:0]   _zz_8084;
  wire       [23:0]   _zz_8085;
  wire       [31:0]   _zz_8086;
  wire       [15:0]   _zz_8087;
  wire       [15:0]   _zz_8088;
  wire       [31:0]   _zz_8089;
  wire       [31:0]   _zz_8090;
  wire       [15:0]   _zz_8091;
  wire       [31:0]   _zz_8092;
  wire       [31:0]   _zz_8093;
  wire       [31:0]   _zz_8094;
  wire       [15:0]   _zz_8095;
  wire       [31:0]   _zz_8096;
  wire       [31:0]   _zz_8097;
  wire       [31:0]   _zz_8098;
  wire       [31:0]   _zz_8099;
  wire       [31:0]   _zz_8100;
  wire       [31:0]   _zz_8101;
  wire       [23:0]   _zz_8102;
  wire       [31:0]   _zz_8103;
  wire       [15:0]   _zz_8104;
  wire       [31:0]   _zz_8105;
  wire       [31:0]   _zz_8106;
  wire       [31:0]   _zz_8107;
  wire       [31:0]   _zz_8108;
  wire       [31:0]   _zz_8109;
  wire       [23:0]   _zz_8110;
  wire       [31:0]   _zz_8111;
  wire       [15:0]   _zz_8112;
  wire       [31:0]   _zz_8113;
  wire       [31:0]   _zz_8114;
  wire       [31:0]   _zz_8115;
  wire       [31:0]   _zz_8116;
  wire       [31:0]   _zz_8117;
  wire       [23:0]   _zz_8118;
  wire       [31:0]   _zz_8119;
  wire       [15:0]   _zz_8120;
  wire       [31:0]   _zz_8121;
  wire       [31:0]   _zz_8122;
  wire       [31:0]   _zz_8123;
  wire       [31:0]   _zz_8124;
  wire       [31:0]   _zz_8125;
  wire       [23:0]   _zz_8126;
  wire       [31:0]   _zz_8127;
  wire       [15:0]   _zz_8128;
  wire       [15:0]   _zz_8129;
  wire       [31:0]   _zz_8130;
  wire       [31:0]   _zz_8131;
  wire       [15:0]   _zz_8132;
  wire       [31:0]   _zz_8133;
  wire       [31:0]   _zz_8134;
  wire       [31:0]   _zz_8135;
  wire       [15:0]   _zz_8136;
  wire       [31:0]   _zz_8137;
  wire       [31:0]   _zz_8138;
  wire       [31:0]   _zz_8139;
  wire       [31:0]   _zz_8140;
  wire       [31:0]   _zz_8141;
  wire       [31:0]   _zz_8142;
  wire       [23:0]   _zz_8143;
  wire       [31:0]   _zz_8144;
  wire       [15:0]   _zz_8145;
  wire       [31:0]   _zz_8146;
  wire       [31:0]   _zz_8147;
  wire       [31:0]   _zz_8148;
  wire       [31:0]   _zz_8149;
  wire       [31:0]   _zz_8150;
  wire       [23:0]   _zz_8151;
  wire       [31:0]   _zz_8152;
  wire       [15:0]   _zz_8153;
  wire       [31:0]   _zz_8154;
  wire       [31:0]   _zz_8155;
  wire       [31:0]   _zz_8156;
  wire       [31:0]   _zz_8157;
  wire       [31:0]   _zz_8158;
  wire       [23:0]   _zz_8159;
  wire       [31:0]   _zz_8160;
  wire       [15:0]   _zz_8161;
  wire       [31:0]   _zz_8162;
  wire       [31:0]   _zz_8163;
  wire       [31:0]   _zz_8164;
  wire       [31:0]   _zz_8165;
  wire       [31:0]   _zz_8166;
  wire       [23:0]   _zz_8167;
  wire       [31:0]   _zz_8168;
  wire       [15:0]   _zz_8169;
  wire       [15:0]   _zz_8170;
  wire       [31:0]   _zz_8171;
  wire       [31:0]   _zz_8172;
  wire       [15:0]   _zz_8173;
  wire       [31:0]   _zz_8174;
  wire       [31:0]   _zz_8175;
  wire       [31:0]   _zz_8176;
  wire       [15:0]   _zz_8177;
  wire       [31:0]   _zz_8178;
  wire       [31:0]   _zz_8179;
  wire       [31:0]   _zz_8180;
  wire       [31:0]   _zz_8181;
  wire       [31:0]   _zz_8182;
  wire       [31:0]   _zz_8183;
  wire       [23:0]   _zz_8184;
  wire       [31:0]   _zz_8185;
  wire       [15:0]   _zz_8186;
  wire       [31:0]   _zz_8187;
  wire       [31:0]   _zz_8188;
  wire       [31:0]   _zz_8189;
  wire       [31:0]   _zz_8190;
  wire       [31:0]   _zz_8191;
  wire       [23:0]   _zz_8192;
  wire       [31:0]   _zz_8193;
  wire       [15:0]   _zz_8194;
  wire       [31:0]   _zz_8195;
  wire       [31:0]   _zz_8196;
  wire       [31:0]   _zz_8197;
  wire       [31:0]   _zz_8198;
  wire       [31:0]   _zz_8199;
  wire       [23:0]   _zz_8200;
  wire       [31:0]   _zz_8201;
  wire       [15:0]   _zz_8202;
  wire       [31:0]   _zz_8203;
  wire       [31:0]   _zz_8204;
  wire       [31:0]   _zz_8205;
  wire       [31:0]   _zz_8206;
  wire       [31:0]   _zz_8207;
  wire       [23:0]   _zz_8208;
  wire       [31:0]   _zz_8209;
  wire       [15:0]   _zz_8210;
  wire       [15:0]   _zz_8211;
  wire       [31:0]   _zz_8212;
  wire       [31:0]   _zz_8213;
  wire       [15:0]   _zz_8214;
  wire       [31:0]   _zz_8215;
  wire       [31:0]   _zz_8216;
  wire       [31:0]   _zz_8217;
  wire       [15:0]   _zz_8218;
  wire       [31:0]   _zz_8219;
  wire       [31:0]   _zz_8220;
  wire       [31:0]   _zz_8221;
  wire       [31:0]   _zz_8222;
  wire       [31:0]   _zz_8223;
  wire       [31:0]   _zz_8224;
  wire       [23:0]   _zz_8225;
  wire       [31:0]   _zz_8226;
  wire       [15:0]   _zz_8227;
  wire       [31:0]   _zz_8228;
  wire       [31:0]   _zz_8229;
  wire       [31:0]   _zz_8230;
  wire       [31:0]   _zz_8231;
  wire       [31:0]   _zz_8232;
  wire       [23:0]   _zz_8233;
  wire       [31:0]   _zz_8234;
  wire       [15:0]   _zz_8235;
  wire       [31:0]   _zz_8236;
  wire       [31:0]   _zz_8237;
  wire       [31:0]   _zz_8238;
  wire       [31:0]   _zz_8239;
  wire       [31:0]   _zz_8240;
  wire       [23:0]   _zz_8241;
  wire       [31:0]   _zz_8242;
  wire       [15:0]   _zz_8243;
  wire       [31:0]   _zz_8244;
  wire       [31:0]   _zz_8245;
  wire       [31:0]   _zz_8246;
  wire       [31:0]   _zz_8247;
  wire       [31:0]   _zz_8248;
  wire       [23:0]   _zz_8249;
  wire       [31:0]   _zz_8250;
  wire       [15:0]   _zz_8251;
  wire       [15:0]   _zz_8252;
  wire       [31:0]   _zz_8253;
  wire       [31:0]   _zz_8254;
  wire       [15:0]   _zz_8255;
  wire       [31:0]   _zz_8256;
  wire       [31:0]   _zz_8257;
  wire       [31:0]   _zz_8258;
  wire       [15:0]   _zz_8259;
  wire       [31:0]   _zz_8260;
  wire       [31:0]   _zz_8261;
  wire       [31:0]   _zz_8262;
  wire       [31:0]   _zz_8263;
  wire       [31:0]   _zz_8264;
  wire       [31:0]   _zz_8265;
  wire       [23:0]   _zz_8266;
  wire       [31:0]   _zz_8267;
  wire       [15:0]   _zz_8268;
  wire       [31:0]   _zz_8269;
  wire       [31:0]   _zz_8270;
  wire       [31:0]   _zz_8271;
  wire       [31:0]   _zz_8272;
  wire       [31:0]   _zz_8273;
  wire       [23:0]   _zz_8274;
  wire       [31:0]   _zz_8275;
  wire       [15:0]   _zz_8276;
  wire       [31:0]   _zz_8277;
  wire       [31:0]   _zz_8278;
  wire       [31:0]   _zz_8279;
  wire       [31:0]   _zz_8280;
  wire       [31:0]   _zz_8281;
  wire       [23:0]   _zz_8282;
  wire       [31:0]   _zz_8283;
  wire       [15:0]   _zz_8284;
  wire       [31:0]   _zz_8285;
  wire       [31:0]   _zz_8286;
  wire       [31:0]   _zz_8287;
  wire       [31:0]   _zz_8288;
  wire       [31:0]   _zz_8289;
  wire       [23:0]   _zz_8290;
  wire       [31:0]   _zz_8291;
  wire       [15:0]   _zz_8292;
  wire       [15:0]   _zz_8293;
  wire       [31:0]   _zz_8294;
  wire       [31:0]   _zz_8295;
  wire       [15:0]   _zz_8296;
  wire       [31:0]   _zz_8297;
  wire       [31:0]   _zz_8298;
  wire       [31:0]   _zz_8299;
  wire       [15:0]   _zz_8300;
  wire       [31:0]   _zz_8301;
  wire       [31:0]   _zz_8302;
  wire       [31:0]   _zz_8303;
  wire       [31:0]   _zz_8304;
  wire       [31:0]   _zz_8305;
  wire       [31:0]   _zz_8306;
  wire       [23:0]   _zz_8307;
  wire       [31:0]   _zz_8308;
  wire       [15:0]   _zz_8309;
  wire       [31:0]   _zz_8310;
  wire       [31:0]   _zz_8311;
  wire       [31:0]   _zz_8312;
  wire       [31:0]   _zz_8313;
  wire       [31:0]   _zz_8314;
  wire       [23:0]   _zz_8315;
  wire       [31:0]   _zz_8316;
  wire       [15:0]   _zz_8317;
  wire       [31:0]   _zz_8318;
  wire       [31:0]   _zz_8319;
  wire       [31:0]   _zz_8320;
  wire       [31:0]   _zz_8321;
  wire       [31:0]   _zz_8322;
  wire       [23:0]   _zz_8323;
  wire       [31:0]   _zz_8324;
  wire       [15:0]   _zz_8325;
  wire       [31:0]   _zz_8326;
  wire       [31:0]   _zz_8327;
  wire       [31:0]   _zz_8328;
  wire       [31:0]   _zz_8329;
  wire       [31:0]   _zz_8330;
  wire       [23:0]   _zz_8331;
  wire       [31:0]   _zz_8332;
  wire       [15:0]   _zz_8333;
  wire       [15:0]   _zz_8334;
  wire       [31:0]   _zz_8335;
  wire       [31:0]   _zz_8336;
  wire       [15:0]   _zz_8337;
  wire       [31:0]   _zz_8338;
  wire       [31:0]   _zz_8339;
  wire       [31:0]   _zz_8340;
  wire       [15:0]   _zz_8341;
  wire       [31:0]   _zz_8342;
  wire       [31:0]   _zz_8343;
  wire       [31:0]   _zz_8344;
  wire       [31:0]   _zz_8345;
  wire       [31:0]   _zz_8346;
  wire       [31:0]   _zz_8347;
  wire       [23:0]   _zz_8348;
  wire       [31:0]   _zz_8349;
  wire       [15:0]   _zz_8350;
  wire       [31:0]   _zz_8351;
  wire       [31:0]   _zz_8352;
  wire       [31:0]   _zz_8353;
  wire       [31:0]   _zz_8354;
  wire       [31:0]   _zz_8355;
  wire       [23:0]   _zz_8356;
  wire       [31:0]   _zz_8357;
  wire       [15:0]   _zz_8358;
  wire       [31:0]   _zz_8359;
  wire       [31:0]   _zz_8360;
  wire       [31:0]   _zz_8361;
  wire       [31:0]   _zz_8362;
  wire       [31:0]   _zz_8363;
  wire       [23:0]   _zz_8364;
  wire       [31:0]   _zz_8365;
  wire       [15:0]   _zz_8366;
  wire       [31:0]   _zz_8367;
  wire       [31:0]   _zz_8368;
  wire       [31:0]   _zz_8369;
  wire       [31:0]   _zz_8370;
  wire       [31:0]   _zz_8371;
  wire       [23:0]   _zz_8372;
  wire       [31:0]   _zz_8373;
  wire       [15:0]   _zz_8374;
  wire       [15:0]   _zz_8375;
  wire       [31:0]   _zz_8376;
  wire       [31:0]   _zz_8377;
  wire       [15:0]   _zz_8378;
  wire       [31:0]   _zz_8379;
  wire       [31:0]   _zz_8380;
  wire       [31:0]   _zz_8381;
  wire       [15:0]   _zz_8382;
  wire       [31:0]   _zz_8383;
  wire       [31:0]   _zz_8384;
  wire       [31:0]   _zz_8385;
  wire       [31:0]   _zz_8386;
  wire       [31:0]   _zz_8387;
  wire       [31:0]   _zz_8388;
  wire       [23:0]   _zz_8389;
  wire       [31:0]   _zz_8390;
  wire       [15:0]   _zz_8391;
  wire       [31:0]   _zz_8392;
  wire       [31:0]   _zz_8393;
  wire       [31:0]   _zz_8394;
  wire       [31:0]   _zz_8395;
  wire       [31:0]   _zz_8396;
  wire       [23:0]   _zz_8397;
  wire       [31:0]   _zz_8398;
  wire       [15:0]   _zz_8399;
  wire       [31:0]   _zz_8400;
  wire       [31:0]   _zz_8401;
  wire       [31:0]   _zz_8402;
  wire       [31:0]   _zz_8403;
  wire       [31:0]   _zz_8404;
  wire       [23:0]   _zz_8405;
  wire       [31:0]   _zz_8406;
  wire       [15:0]   _zz_8407;
  wire       [31:0]   _zz_8408;
  wire       [31:0]   _zz_8409;
  wire       [31:0]   _zz_8410;
  wire       [31:0]   _zz_8411;
  wire       [31:0]   _zz_8412;
  wire       [23:0]   _zz_8413;
  wire       [31:0]   _zz_8414;
  wire       [15:0]   _zz_8415;
  wire       [15:0]   _zz_8416;
  wire       [31:0]   _zz_8417;
  wire       [31:0]   _zz_8418;
  wire       [15:0]   _zz_8419;
  wire       [31:0]   _zz_8420;
  wire       [31:0]   _zz_8421;
  wire       [31:0]   _zz_8422;
  wire       [15:0]   _zz_8423;
  wire       [31:0]   _zz_8424;
  wire       [31:0]   _zz_8425;
  wire       [31:0]   _zz_8426;
  wire       [31:0]   _zz_8427;
  wire       [31:0]   _zz_8428;
  wire       [31:0]   _zz_8429;
  wire       [23:0]   _zz_8430;
  wire       [31:0]   _zz_8431;
  wire       [15:0]   _zz_8432;
  wire       [31:0]   _zz_8433;
  wire       [31:0]   _zz_8434;
  wire       [31:0]   _zz_8435;
  wire       [31:0]   _zz_8436;
  wire       [31:0]   _zz_8437;
  wire       [23:0]   _zz_8438;
  wire       [31:0]   _zz_8439;
  wire       [15:0]   _zz_8440;
  wire       [31:0]   _zz_8441;
  wire       [31:0]   _zz_8442;
  wire       [31:0]   _zz_8443;
  wire       [31:0]   _zz_8444;
  wire       [31:0]   _zz_8445;
  wire       [23:0]   _zz_8446;
  wire       [31:0]   _zz_8447;
  wire       [15:0]   _zz_8448;
  wire       [31:0]   _zz_8449;
  wire       [31:0]   _zz_8450;
  wire       [31:0]   _zz_8451;
  wire       [31:0]   _zz_8452;
  wire       [31:0]   _zz_8453;
  wire       [23:0]   _zz_8454;
  wire       [31:0]   _zz_8455;
  wire       [15:0]   _zz_8456;
  wire       [15:0]   _zz_8457;
  wire       [31:0]   _zz_8458;
  wire       [31:0]   _zz_8459;
  wire       [15:0]   _zz_8460;
  wire       [31:0]   _zz_8461;
  wire       [31:0]   _zz_8462;
  wire       [31:0]   _zz_8463;
  wire       [15:0]   _zz_8464;
  wire       [31:0]   _zz_8465;
  wire       [31:0]   _zz_8466;
  wire       [31:0]   _zz_8467;
  wire       [31:0]   _zz_8468;
  wire       [31:0]   _zz_8469;
  wire       [31:0]   _zz_8470;
  wire       [23:0]   _zz_8471;
  wire       [31:0]   _zz_8472;
  wire       [15:0]   _zz_8473;
  wire       [31:0]   _zz_8474;
  wire       [31:0]   _zz_8475;
  wire       [31:0]   _zz_8476;
  wire       [31:0]   _zz_8477;
  wire       [31:0]   _zz_8478;
  wire       [23:0]   _zz_8479;
  wire       [31:0]   _zz_8480;
  wire       [15:0]   _zz_8481;
  wire       [31:0]   _zz_8482;
  wire       [31:0]   _zz_8483;
  wire       [31:0]   _zz_8484;
  wire       [31:0]   _zz_8485;
  wire       [31:0]   _zz_8486;
  wire       [23:0]   _zz_8487;
  wire       [31:0]   _zz_8488;
  wire       [15:0]   _zz_8489;
  wire       [31:0]   _zz_8490;
  wire       [31:0]   _zz_8491;
  wire       [31:0]   _zz_8492;
  wire       [31:0]   _zz_8493;
  wire       [31:0]   _zz_8494;
  wire       [23:0]   _zz_8495;
  wire       [31:0]   _zz_8496;
  wire       [15:0]   _zz_8497;
  wire       [15:0]   _zz_8498;
  wire       [31:0]   _zz_8499;
  wire       [31:0]   _zz_8500;
  wire       [15:0]   _zz_8501;
  wire       [31:0]   _zz_8502;
  wire       [31:0]   _zz_8503;
  wire       [31:0]   _zz_8504;
  wire       [15:0]   _zz_8505;
  wire       [31:0]   _zz_8506;
  wire       [31:0]   _zz_8507;
  wire       [31:0]   _zz_8508;
  wire       [31:0]   _zz_8509;
  wire       [31:0]   _zz_8510;
  wire       [31:0]   _zz_8511;
  wire       [23:0]   _zz_8512;
  wire       [31:0]   _zz_8513;
  wire       [15:0]   _zz_8514;
  wire       [31:0]   _zz_8515;
  wire       [31:0]   _zz_8516;
  wire       [31:0]   _zz_8517;
  wire       [31:0]   _zz_8518;
  wire       [31:0]   _zz_8519;
  wire       [23:0]   _zz_8520;
  wire       [31:0]   _zz_8521;
  wire       [15:0]   _zz_8522;
  wire       [31:0]   _zz_8523;
  wire       [31:0]   _zz_8524;
  wire       [31:0]   _zz_8525;
  wire       [31:0]   _zz_8526;
  wire       [31:0]   _zz_8527;
  wire       [23:0]   _zz_8528;
  wire       [31:0]   _zz_8529;
  wire       [15:0]   _zz_8530;
  wire       [31:0]   _zz_8531;
  wire       [31:0]   _zz_8532;
  wire       [31:0]   _zz_8533;
  wire       [31:0]   _zz_8534;
  wire       [31:0]   _zz_8535;
  wire       [23:0]   _zz_8536;
  wire       [31:0]   _zz_8537;
  wire       [15:0]   _zz_8538;
  wire       [15:0]   _zz_8539;
  wire       [31:0]   _zz_8540;
  wire       [31:0]   _zz_8541;
  wire       [15:0]   _zz_8542;
  wire       [31:0]   _zz_8543;
  wire       [31:0]   _zz_8544;
  wire       [31:0]   _zz_8545;
  wire       [15:0]   _zz_8546;
  wire       [31:0]   _zz_8547;
  wire       [31:0]   _zz_8548;
  wire       [31:0]   _zz_8549;
  wire       [31:0]   _zz_8550;
  wire       [31:0]   _zz_8551;
  wire       [31:0]   _zz_8552;
  wire       [23:0]   _zz_8553;
  wire       [31:0]   _zz_8554;
  wire       [15:0]   _zz_8555;
  wire       [31:0]   _zz_8556;
  wire       [31:0]   _zz_8557;
  wire       [31:0]   _zz_8558;
  wire       [31:0]   _zz_8559;
  wire       [31:0]   _zz_8560;
  wire       [23:0]   _zz_8561;
  wire       [31:0]   _zz_8562;
  wire       [15:0]   _zz_8563;
  wire       [31:0]   _zz_8564;
  wire       [31:0]   _zz_8565;
  wire       [31:0]   _zz_8566;
  wire       [31:0]   _zz_8567;
  wire       [31:0]   _zz_8568;
  wire       [23:0]   _zz_8569;
  wire       [31:0]   _zz_8570;
  wire       [15:0]   _zz_8571;
  wire       [31:0]   _zz_8572;
  wire       [31:0]   _zz_8573;
  wire       [31:0]   _zz_8574;
  wire       [31:0]   _zz_8575;
  wire       [31:0]   _zz_8576;
  wire       [23:0]   _zz_8577;
  wire       [31:0]   _zz_8578;
  wire       [15:0]   _zz_8579;
  wire       [15:0]   _zz_8580;
  wire       [31:0]   _zz_8581;
  wire       [31:0]   _zz_8582;
  wire       [15:0]   _zz_8583;
  wire       [31:0]   _zz_8584;
  wire       [31:0]   _zz_8585;
  wire       [31:0]   _zz_8586;
  wire       [15:0]   _zz_8587;
  wire       [31:0]   _zz_8588;
  wire       [31:0]   _zz_8589;
  wire       [31:0]   _zz_8590;
  wire       [31:0]   _zz_8591;
  wire       [31:0]   _zz_8592;
  wire       [31:0]   _zz_8593;
  wire       [23:0]   _zz_8594;
  wire       [31:0]   _zz_8595;
  wire       [15:0]   _zz_8596;
  wire       [31:0]   _zz_8597;
  wire       [31:0]   _zz_8598;
  wire       [31:0]   _zz_8599;
  wire       [31:0]   _zz_8600;
  wire       [31:0]   _zz_8601;
  wire       [23:0]   _zz_8602;
  wire       [31:0]   _zz_8603;
  wire       [15:0]   _zz_8604;
  wire       [31:0]   _zz_8605;
  wire       [31:0]   _zz_8606;
  wire       [31:0]   _zz_8607;
  wire       [31:0]   _zz_8608;
  wire       [31:0]   _zz_8609;
  wire       [23:0]   _zz_8610;
  wire       [31:0]   _zz_8611;
  wire       [15:0]   _zz_8612;
  wire       [31:0]   _zz_8613;
  wire       [31:0]   _zz_8614;
  wire       [31:0]   _zz_8615;
  wire       [31:0]   _zz_8616;
  wire       [31:0]   _zz_8617;
  wire       [23:0]   _zz_8618;
  wire       [31:0]   _zz_8619;
  wire       [15:0]   _zz_8620;
  wire       [15:0]   _zz_8621;
  wire       [31:0]   _zz_8622;
  wire       [31:0]   _zz_8623;
  wire       [15:0]   _zz_8624;
  wire       [31:0]   _zz_8625;
  wire       [31:0]   _zz_8626;
  wire       [31:0]   _zz_8627;
  wire       [15:0]   _zz_8628;
  wire       [31:0]   _zz_8629;
  wire       [31:0]   _zz_8630;
  wire       [31:0]   _zz_8631;
  wire       [31:0]   _zz_8632;
  wire       [31:0]   _zz_8633;
  wire       [31:0]   _zz_8634;
  wire       [23:0]   _zz_8635;
  wire       [31:0]   _zz_8636;
  wire       [15:0]   _zz_8637;
  wire       [31:0]   _zz_8638;
  wire       [31:0]   _zz_8639;
  wire       [31:0]   _zz_8640;
  wire       [31:0]   _zz_8641;
  wire       [31:0]   _zz_8642;
  wire       [23:0]   _zz_8643;
  wire       [31:0]   _zz_8644;
  wire       [15:0]   _zz_8645;
  wire       [31:0]   _zz_8646;
  wire       [31:0]   _zz_8647;
  wire       [31:0]   _zz_8648;
  wire       [31:0]   _zz_8649;
  wire       [31:0]   _zz_8650;
  wire       [23:0]   _zz_8651;
  wire       [31:0]   _zz_8652;
  wire       [15:0]   _zz_8653;
  wire       [31:0]   _zz_8654;
  wire       [31:0]   _zz_8655;
  wire       [31:0]   _zz_8656;
  wire       [31:0]   _zz_8657;
  wire       [31:0]   _zz_8658;
  wire       [23:0]   _zz_8659;
  wire       [31:0]   _zz_8660;
  wire       [15:0]   _zz_8661;
  wire       [15:0]   _zz_8662;
  wire       [31:0]   _zz_8663;
  wire       [31:0]   _zz_8664;
  wire       [15:0]   _zz_8665;
  wire       [31:0]   _zz_8666;
  wire       [31:0]   _zz_8667;
  wire       [31:0]   _zz_8668;
  wire       [15:0]   _zz_8669;
  wire       [31:0]   _zz_8670;
  wire       [31:0]   _zz_8671;
  wire       [31:0]   _zz_8672;
  wire       [31:0]   _zz_8673;
  wire       [31:0]   _zz_8674;
  wire       [31:0]   _zz_8675;
  wire       [23:0]   _zz_8676;
  wire       [31:0]   _zz_8677;
  wire       [15:0]   _zz_8678;
  wire       [31:0]   _zz_8679;
  wire       [31:0]   _zz_8680;
  wire       [31:0]   _zz_8681;
  wire       [31:0]   _zz_8682;
  wire       [31:0]   _zz_8683;
  wire       [23:0]   _zz_8684;
  wire       [31:0]   _zz_8685;
  wire       [15:0]   _zz_8686;
  wire       [31:0]   _zz_8687;
  wire       [31:0]   _zz_8688;
  wire       [31:0]   _zz_8689;
  wire       [31:0]   _zz_8690;
  wire       [31:0]   _zz_8691;
  wire       [23:0]   _zz_8692;
  wire       [31:0]   _zz_8693;
  wire       [15:0]   _zz_8694;
  wire       [31:0]   _zz_8695;
  wire       [31:0]   _zz_8696;
  wire       [31:0]   _zz_8697;
  wire       [31:0]   _zz_8698;
  wire       [31:0]   _zz_8699;
  wire       [23:0]   _zz_8700;
  wire       [31:0]   _zz_8701;
  wire       [15:0]   _zz_8702;
  wire       [15:0]   _zz_8703;
  wire       [31:0]   _zz_8704;
  wire       [31:0]   _zz_8705;
  wire       [15:0]   _zz_8706;
  wire       [31:0]   _zz_8707;
  wire       [31:0]   _zz_8708;
  wire       [31:0]   _zz_8709;
  wire       [15:0]   _zz_8710;
  wire       [31:0]   _zz_8711;
  wire       [31:0]   _zz_8712;
  wire       [31:0]   _zz_8713;
  wire       [31:0]   _zz_8714;
  wire       [31:0]   _zz_8715;
  wire       [31:0]   _zz_8716;
  wire       [23:0]   _zz_8717;
  wire       [31:0]   _zz_8718;
  wire       [15:0]   _zz_8719;
  wire       [31:0]   _zz_8720;
  wire       [31:0]   _zz_8721;
  wire       [31:0]   _zz_8722;
  wire       [31:0]   _zz_8723;
  wire       [31:0]   _zz_8724;
  wire       [23:0]   _zz_8725;
  wire       [31:0]   _zz_8726;
  wire       [15:0]   _zz_8727;
  wire       [31:0]   _zz_8728;
  wire       [31:0]   _zz_8729;
  wire       [31:0]   _zz_8730;
  wire       [31:0]   _zz_8731;
  wire       [31:0]   _zz_8732;
  wire       [23:0]   _zz_8733;
  wire       [31:0]   _zz_8734;
  wire       [15:0]   _zz_8735;
  wire       [31:0]   _zz_8736;
  wire       [31:0]   _zz_8737;
  wire       [31:0]   _zz_8738;
  wire       [31:0]   _zz_8739;
  wire       [31:0]   _zz_8740;
  wire       [23:0]   _zz_8741;
  wire       [31:0]   _zz_8742;
  wire       [15:0]   _zz_8743;
  wire       [15:0]   _zz_8744;
  wire       [31:0]   _zz_8745;
  wire       [31:0]   _zz_8746;
  wire       [15:0]   _zz_8747;
  wire       [31:0]   _zz_8748;
  wire       [31:0]   _zz_8749;
  wire       [31:0]   _zz_8750;
  wire       [15:0]   _zz_8751;
  wire       [31:0]   _zz_8752;
  wire       [31:0]   _zz_8753;
  wire       [31:0]   _zz_8754;
  wire       [31:0]   _zz_8755;
  wire       [31:0]   _zz_8756;
  wire       [31:0]   _zz_8757;
  wire       [23:0]   _zz_8758;
  wire       [31:0]   _zz_8759;
  wire       [15:0]   _zz_8760;
  wire       [31:0]   _zz_8761;
  wire       [31:0]   _zz_8762;
  wire       [31:0]   _zz_8763;
  wire       [31:0]   _zz_8764;
  wire       [31:0]   _zz_8765;
  wire       [23:0]   _zz_8766;
  wire       [31:0]   _zz_8767;
  wire       [15:0]   _zz_8768;
  wire       [31:0]   _zz_8769;
  wire       [31:0]   _zz_8770;
  wire       [31:0]   _zz_8771;
  wire       [31:0]   _zz_8772;
  wire       [31:0]   _zz_8773;
  wire       [23:0]   _zz_8774;
  wire       [31:0]   _zz_8775;
  wire       [15:0]   _zz_8776;
  wire       [31:0]   _zz_8777;
  wire       [31:0]   _zz_8778;
  wire       [31:0]   _zz_8779;
  wire       [31:0]   _zz_8780;
  wire       [31:0]   _zz_8781;
  wire       [23:0]   _zz_8782;
  wire       [31:0]   _zz_8783;
  wire       [15:0]   _zz_8784;
  wire       [15:0]   _zz_8785;
  wire       [31:0]   _zz_8786;
  wire       [31:0]   _zz_8787;
  wire       [15:0]   _zz_8788;
  wire       [31:0]   _zz_8789;
  wire       [31:0]   _zz_8790;
  wire       [31:0]   _zz_8791;
  wire       [15:0]   _zz_8792;
  wire       [31:0]   _zz_8793;
  wire       [31:0]   _zz_8794;
  wire       [31:0]   _zz_8795;
  wire       [31:0]   _zz_8796;
  wire       [31:0]   _zz_8797;
  wire       [31:0]   _zz_8798;
  wire       [23:0]   _zz_8799;
  wire       [31:0]   _zz_8800;
  wire       [15:0]   _zz_8801;
  wire       [31:0]   _zz_8802;
  wire       [31:0]   _zz_8803;
  wire       [31:0]   _zz_8804;
  wire       [31:0]   _zz_8805;
  wire       [31:0]   _zz_8806;
  wire       [23:0]   _zz_8807;
  wire       [31:0]   _zz_8808;
  wire       [15:0]   _zz_8809;
  wire       [31:0]   _zz_8810;
  wire       [31:0]   _zz_8811;
  wire       [31:0]   _zz_8812;
  wire       [31:0]   _zz_8813;
  wire       [31:0]   _zz_8814;
  wire       [23:0]   _zz_8815;
  wire       [31:0]   _zz_8816;
  wire       [15:0]   _zz_8817;
  wire       [31:0]   _zz_8818;
  wire       [31:0]   _zz_8819;
  wire       [31:0]   _zz_8820;
  wire       [31:0]   _zz_8821;
  wire       [31:0]   _zz_8822;
  wire       [23:0]   _zz_8823;
  wire       [31:0]   _zz_8824;
  wire       [15:0]   _zz_8825;
  wire       [15:0]   _zz_8826;
  wire       [31:0]   _zz_8827;
  wire       [31:0]   _zz_8828;
  wire       [15:0]   _zz_8829;
  wire       [31:0]   _zz_8830;
  wire       [31:0]   _zz_8831;
  wire       [31:0]   _zz_8832;
  wire       [15:0]   _zz_8833;
  wire       [31:0]   _zz_8834;
  wire       [31:0]   _zz_8835;
  wire       [31:0]   _zz_8836;
  wire       [31:0]   _zz_8837;
  wire       [31:0]   _zz_8838;
  wire       [31:0]   _zz_8839;
  wire       [23:0]   _zz_8840;
  wire       [31:0]   _zz_8841;
  wire       [15:0]   _zz_8842;
  wire       [31:0]   _zz_8843;
  wire       [31:0]   _zz_8844;
  wire       [31:0]   _zz_8845;
  wire       [31:0]   _zz_8846;
  wire       [31:0]   _zz_8847;
  wire       [23:0]   _zz_8848;
  wire       [31:0]   _zz_8849;
  wire       [15:0]   _zz_8850;
  wire       [31:0]   _zz_8851;
  wire       [31:0]   _zz_8852;
  wire       [31:0]   _zz_8853;
  wire       [31:0]   _zz_8854;
  wire       [31:0]   _zz_8855;
  wire       [23:0]   _zz_8856;
  wire       [31:0]   _zz_8857;
  wire       [15:0]   _zz_8858;
  wire       [31:0]   _zz_8859;
  wire       [31:0]   _zz_8860;
  wire       [31:0]   _zz_8861;
  wire       [31:0]   _zz_8862;
  wire       [31:0]   _zz_8863;
  wire       [23:0]   _zz_8864;
  wire       [31:0]   _zz_8865;
  wire       [15:0]   _zz_8866;
  wire       [15:0]   _zz_8867;
  wire       [31:0]   _zz_8868;
  wire       [31:0]   _zz_8869;
  wire       [15:0]   _zz_8870;
  wire       [31:0]   _zz_8871;
  wire       [31:0]   _zz_8872;
  wire       [31:0]   _zz_8873;
  wire       [15:0]   _zz_8874;
  wire       [31:0]   _zz_8875;
  wire       [31:0]   _zz_8876;
  wire       [31:0]   _zz_8877;
  wire       [31:0]   _zz_8878;
  wire       [31:0]   _zz_8879;
  wire       [31:0]   _zz_8880;
  wire       [23:0]   _zz_8881;
  wire       [31:0]   _zz_8882;
  wire       [15:0]   _zz_8883;
  wire       [31:0]   _zz_8884;
  wire       [31:0]   _zz_8885;
  wire       [31:0]   _zz_8886;
  wire       [31:0]   _zz_8887;
  wire       [31:0]   _zz_8888;
  wire       [23:0]   _zz_8889;
  wire       [31:0]   _zz_8890;
  wire       [15:0]   _zz_8891;
  wire       [31:0]   _zz_8892;
  wire       [31:0]   _zz_8893;
  wire       [31:0]   _zz_8894;
  wire       [31:0]   _zz_8895;
  wire       [31:0]   _zz_8896;
  wire       [23:0]   _zz_8897;
  wire       [31:0]   _zz_8898;
  wire       [15:0]   _zz_8899;
  wire       [31:0]   _zz_8900;
  wire       [31:0]   _zz_8901;
  wire       [31:0]   _zz_8902;
  wire       [31:0]   _zz_8903;
  wire       [31:0]   _zz_8904;
  wire       [23:0]   _zz_8905;
  wire       [31:0]   _zz_8906;
  wire       [15:0]   _zz_8907;
  wire       [15:0]   _zz_8908;
  wire       [31:0]   _zz_8909;
  wire       [31:0]   _zz_8910;
  wire       [15:0]   _zz_8911;
  wire       [31:0]   _zz_8912;
  wire       [31:0]   _zz_8913;
  wire       [31:0]   _zz_8914;
  wire       [15:0]   _zz_8915;
  wire       [31:0]   _zz_8916;
  wire       [31:0]   _zz_8917;
  wire       [31:0]   _zz_8918;
  wire       [31:0]   _zz_8919;
  wire       [31:0]   _zz_8920;
  wire       [31:0]   _zz_8921;
  wire       [23:0]   _zz_8922;
  wire       [31:0]   _zz_8923;
  wire       [15:0]   _zz_8924;
  wire       [31:0]   _zz_8925;
  wire       [31:0]   _zz_8926;
  wire       [31:0]   _zz_8927;
  wire       [31:0]   _zz_8928;
  wire       [31:0]   _zz_8929;
  wire       [23:0]   _zz_8930;
  wire       [31:0]   _zz_8931;
  wire       [15:0]   _zz_8932;
  wire       [31:0]   _zz_8933;
  wire       [31:0]   _zz_8934;
  wire       [31:0]   _zz_8935;
  wire       [31:0]   _zz_8936;
  wire       [31:0]   _zz_8937;
  wire       [23:0]   _zz_8938;
  wire       [31:0]   _zz_8939;
  wire       [15:0]   _zz_8940;
  wire       [31:0]   _zz_8941;
  wire       [31:0]   _zz_8942;
  wire       [31:0]   _zz_8943;
  wire       [31:0]   _zz_8944;
  wire       [31:0]   _zz_8945;
  wire       [23:0]   _zz_8946;
  wire       [31:0]   _zz_8947;
  wire       [15:0]   _zz_8948;
  wire       [15:0]   _zz_8949;
  wire       [31:0]   _zz_8950;
  wire       [31:0]   _zz_8951;
  wire       [15:0]   _zz_8952;
  wire       [31:0]   _zz_8953;
  wire       [31:0]   _zz_8954;
  wire       [31:0]   _zz_8955;
  wire       [15:0]   _zz_8956;
  wire       [31:0]   _zz_8957;
  wire       [31:0]   _zz_8958;
  wire       [31:0]   _zz_8959;
  wire       [31:0]   _zz_8960;
  wire       [31:0]   _zz_8961;
  wire       [31:0]   _zz_8962;
  wire       [23:0]   _zz_8963;
  wire       [31:0]   _zz_8964;
  wire       [15:0]   _zz_8965;
  wire       [31:0]   _zz_8966;
  wire       [31:0]   _zz_8967;
  wire       [31:0]   _zz_8968;
  wire       [31:0]   _zz_8969;
  wire       [31:0]   _zz_8970;
  wire       [23:0]   _zz_8971;
  wire       [31:0]   _zz_8972;
  wire       [15:0]   _zz_8973;
  wire       [31:0]   _zz_8974;
  wire       [31:0]   _zz_8975;
  wire       [31:0]   _zz_8976;
  wire       [31:0]   _zz_8977;
  wire       [31:0]   _zz_8978;
  wire       [23:0]   _zz_8979;
  wire       [31:0]   _zz_8980;
  wire       [15:0]   _zz_8981;
  wire       [31:0]   _zz_8982;
  wire       [31:0]   _zz_8983;
  wire       [31:0]   _zz_8984;
  wire       [31:0]   _zz_8985;
  wire       [31:0]   _zz_8986;
  wire       [23:0]   _zz_8987;
  wire       [31:0]   _zz_8988;
  wire       [15:0]   _zz_8989;
  wire       [15:0]   _zz_8990;
  wire       [31:0]   _zz_8991;
  wire       [31:0]   _zz_8992;
  wire       [15:0]   _zz_8993;
  wire       [31:0]   _zz_8994;
  wire       [31:0]   _zz_8995;
  wire       [31:0]   _zz_8996;
  wire       [15:0]   _zz_8997;
  wire       [31:0]   _zz_8998;
  wire       [31:0]   _zz_8999;
  wire       [31:0]   _zz_9000;
  wire       [31:0]   _zz_9001;
  wire       [31:0]   _zz_9002;
  wire       [31:0]   _zz_9003;
  wire       [23:0]   _zz_9004;
  wire       [31:0]   _zz_9005;
  wire       [15:0]   _zz_9006;
  wire       [31:0]   _zz_9007;
  wire       [31:0]   _zz_9008;
  wire       [31:0]   _zz_9009;
  wire       [31:0]   _zz_9010;
  wire       [31:0]   _zz_9011;
  wire       [23:0]   _zz_9012;
  wire       [31:0]   _zz_9013;
  wire       [15:0]   _zz_9014;
  wire       [31:0]   _zz_9015;
  wire       [31:0]   _zz_9016;
  wire       [31:0]   _zz_9017;
  wire       [31:0]   _zz_9018;
  wire       [31:0]   _zz_9019;
  wire       [23:0]   _zz_9020;
  wire       [31:0]   _zz_9021;
  wire       [15:0]   _zz_9022;
  wire       [31:0]   _zz_9023;
  wire       [31:0]   _zz_9024;
  wire       [31:0]   _zz_9025;
  wire       [31:0]   _zz_9026;
  wire       [31:0]   _zz_9027;
  wire       [23:0]   _zz_9028;
  wire       [31:0]   _zz_9029;
  wire       [15:0]   _zz_9030;
  wire       [15:0]   _zz_9031;
  wire       [31:0]   _zz_9032;
  wire       [31:0]   _zz_9033;
  wire       [15:0]   _zz_9034;
  wire       [31:0]   _zz_9035;
  wire       [31:0]   _zz_9036;
  wire       [31:0]   _zz_9037;
  wire       [15:0]   _zz_9038;
  wire       [31:0]   _zz_9039;
  wire       [31:0]   _zz_9040;
  wire       [31:0]   _zz_9041;
  wire       [31:0]   _zz_9042;
  wire       [31:0]   _zz_9043;
  wire       [31:0]   _zz_9044;
  wire       [23:0]   _zz_9045;
  wire       [31:0]   _zz_9046;
  wire       [15:0]   _zz_9047;
  wire       [31:0]   _zz_9048;
  wire       [31:0]   _zz_9049;
  wire       [31:0]   _zz_9050;
  wire       [31:0]   _zz_9051;
  wire       [31:0]   _zz_9052;
  wire       [23:0]   _zz_9053;
  wire       [31:0]   _zz_9054;
  wire       [15:0]   _zz_9055;
  wire       [31:0]   _zz_9056;
  wire       [31:0]   _zz_9057;
  wire       [31:0]   _zz_9058;
  wire       [31:0]   _zz_9059;
  wire       [31:0]   _zz_9060;
  wire       [23:0]   _zz_9061;
  wire       [31:0]   _zz_9062;
  wire       [15:0]   _zz_9063;
  wire       [31:0]   _zz_9064;
  wire       [31:0]   _zz_9065;
  wire       [31:0]   _zz_9066;
  wire       [31:0]   _zz_9067;
  wire       [31:0]   _zz_9068;
  wire       [23:0]   _zz_9069;
  wire       [31:0]   _zz_9070;
  wire       [15:0]   _zz_9071;
  wire       [15:0]   _zz_9072;
  wire       [31:0]   _zz_9073;
  wire       [31:0]   _zz_9074;
  wire       [15:0]   _zz_9075;
  wire       [31:0]   _zz_9076;
  wire       [31:0]   _zz_9077;
  wire       [31:0]   _zz_9078;
  wire       [15:0]   _zz_9079;
  wire       [31:0]   _zz_9080;
  wire       [31:0]   _zz_9081;
  wire       [31:0]   _zz_9082;
  wire       [31:0]   _zz_9083;
  wire       [31:0]   _zz_9084;
  wire       [31:0]   _zz_9085;
  wire       [23:0]   _zz_9086;
  wire       [31:0]   _zz_9087;
  wire       [15:0]   _zz_9088;
  wire       [31:0]   _zz_9089;
  wire       [31:0]   _zz_9090;
  wire       [31:0]   _zz_9091;
  wire       [31:0]   _zz_9092;
  wire       [31:0]   _zz_9093;
  wire       [23:0]   _zz_9094;
  wire       [31:0]   _zz_9095;
  wire       [15:0]   _zz_9096;
  wire       [31:0]   _zz_9097;
  wire       [31:0]   _zz_9098;
  wire       [31:0]   _zz_9099;
  wire       [31:0]   _zz_9100;
  wire       [31:0]   _zz_9101;
  wire       [23:0]   _zz_9102;
  wire       [31:0]   _zz_9103;
  wire       [15:0]   _zz_9104;
  wire       [31:0]   _zz_9105;
  wire       [31:0]   _zz_9106;
  wire       [31:0]   _zz_9107;
  wire       [31:0]   _zz_9108;
  wire       [31:0]   _zz_9109;
  wire       [23:0]   _zz_9110;
  wire       [31:0]   _zz_9111;
  wire       [15:0]   _zz_9112;
  wire       [15:0]   _zz_9113;
  wire       [31:0]   _zz_9114;
  wire       [31:0]   _zz_9115;
  wire       [15:0]   _zz_9116;
  wire       [31:0]   _zz_9117;
  wire       [31:0]   _zz_9118;
  wire       [31:0]   _zz_9119;
  wire       [15:0]   _zz_9120;
  wire       [31:0]   _zz_9121;
  wire       [31:0]   _zz_9122;
  wire       [31:0]   _zz_9123;
  wire       [31:0]   _zz_9124;
  wire       [31:0]   _zz_9125;
  wire       [31:0]   _zz_9126;
  wire       [23:0]   _zz_9127;
  wire       [31:0]   _zz_9128;
  wire       [15:0]   _zz_9129;
  wire       [31:0]   _zz_9130;
  wire       [31:0]   _zz_9131;
  wire       [31:0]   _zz_9132;
  wire       [31:0]   _zz_9133;
  wire       [31:0]   _zz_9134;
  wire       [23:0]   _zz_9135;
  wire       [31:0]   _zz_9136;
  wire       [15:0]   _zz_9137;
  wire       [31:0]   _zz_9138;
  wire       [31:0]   _zz_9139;
  wire       [31:0]   _zz_9140;
  wire       [31:0]   _zz_9141;
  wire       [31:0]   _zz_9142;
  wire       [23:0]   _zz_9143;
  wire       [31:0]   _zz_9144;
  wire       [15:0]   _zz_9145;
  wire       [31:0]   _zz_9146;
  wire       [31:0]   _zz_9147;
  wire       [31:0]   _zz_9148;
  wire       [31:0]   _zz_9149;
  wire       [31:0]   _zz_9150;
  wire       [23:0]   _zz_9151;
  wire       [31:0]   _zz_9152;
  wire       [15:0]   _zz_9153;
  wire       [15:0]   _zz_9154;
  wire       [31:0]   _zz_9155;
  wire       [31:0]   _zz_9156;
  wire       [15:0]   _zz_9157;
  wire       [31:0]   _zz_9158;
  wire       [31:0]   _zz_9159;
  wire       [31:0]   _zz_9160;
  wire       [15:0]   _zz_9161;
  wire       [31:0]   _zz_9162;
  wire       [31:0]   _zz_9163;
  wire       [31:0]   _zz_9164;
  wire       [31:0]   _zz_9165;
  wire       [31:0]   _zz_9166;
  wire       [31:0]   _zz_9167;
  wire       [23:0]   _zz_9168;
  wire       [31:0]   _zz_9169;
  wire       [15:0]   _zz_9170;
  wire       [31:0]   _zz_9171;
  wire       [31:0]   _zz_9172;
  wire       [31:0]   _zz_9173;
  wire       [31:0]   _zz_9174;
  wire       [31:0]   _zz_9175;
  wire       [23:0]   _zz_9176;
  wire       [31:0]   _zz_9177;
  wire       [15:0]   _zz_9178;
  wire       [31:0]   _zz_9179;
  wire       [31:0]   _zz_9180;
  wire       [31:0]   _zz_9181;
  wire       [31:0]   _zz_9182;
  wire       [31:0]   _zz_9183;
  wire       [23:0]   _zz_9184;
  wire       [31:0]   _zz_9185;
  wire       [15:0]   _zz_9186;
  wire       [31:0]   _zz_9187;
  wire       [31:0]   _zz_9188;
  wire       [31:0]   _zz_9189;
  wire       [31:0]   _zz_9190;
  wire       [31:0]   _zz_9191;
  wire       [23:0]   _zz_9192;
  wire       [31:0]   _zz_9193;
  wire       [15:0]   _zz_9194;
  wire       [15:0]   _zz_9195;
  wire       [31:0]   _zz_9196;
  wire       [31:0]   _zz_9197;
  wire       [15:0]   _zz_9198;
  wire       [31:0]   _zz_9199;
  wire       [31:0]   _zz_9200;
  wire       [31:0]   _zz_9201;
  wire       [15:0]   _zz_9202;
  wire       [31:0]   _zz_9203;
  wire       [31:0]   _zz_9204;
  wire       [31:0]   _zz_9205;
  wire       [31:0]   _zz_9206;
  wire       [31:0]   _zz_9207;
  wire       [31:0]   _zz_9208;
  wire       [23:0]   _zz_9209;
  wire       [31:0]   _zz_9210;
  wire       [15:0]   _zz_9211;
  wire       [31:0]   _zz_9212;
  wire       [31:0]   _zz_9213;
  wire       [31:0]   _zz_9214;
  wire       [31:0]   _zz_9215;
  wire       [31:0]   _zz_9216;
  wire       [23:0]   _zz_9217;
  wire       [31:0]   _zz_9218;
  wire       [15:0]   _zz_9219;
  wire       [31:0]   _zz_9220;
  wire       [31:0]   _zz_9221;
  wire       [31:0]   _zz_9222;
  wire       [31:0]   _zz_9223;
  wire       [31:0]   _zz_9224;
  wire       [23:0]   _zz_9225;
  wire       [31:0]   _zz_9226;
  wire       [15:0]   _zz_9227;
  wire       [31:0]   _zz_9228;
  wire       [31:0]   _zz_9229;
  wire       [31:0]   _zz_9230;
  wire       [31:0]   _zz_9231;
  wire       [31:0]   _zz_9232;
  wire       [23:0]   _zz_9233;
  wire       [31:0]   _zz_9234;
  wire       [15:0]   _zz_9235;
  wire       [15:0]   _zz_9236;
  wire       [31:0]   _zz_9237;
  wire       [31:0]   _zz_9238;
  wire       [15:0]   _zz_9239;
  wire       [31:0]   _zz_9240;
  wire       [31:0]   _zz_9241;
  wire       [31:0]   _zz_9242;
  wire       [15:0]   _zz_9243;
  wire       [31:0]   _zz_9244;
  wire       [31:0]   _zz_9245;
  wire       [31:0]   _zz_9246;
  wire       [31:0]   _zz_9247;
  wire       [31:0]   _zz_9248;
  wire       [31:0]   _zz_9249;
  wire       [23:0]   _zz_9250;
  wire       [31:0]   _zz_9251;
  wire       [15:0]   _zz_9252;
  wire       [31:0]   _zz_9253;
  wire       [31:0]   _zz_9254;
  wire       [31:0]   _zz_9255;
  wire       [31:0]   _zz_9256;
  wire       [31:0]   _zz_9257;
  wire       [23:0]   _zz_9258;
  wire       [31:0]   _zz_9259;
  wire       [15:0]   _zz_9260;
  wire       [31:0]   _zz_9261;
  wire       [31:0]   _zz_9262;
  wire       [31:0]   _zz_9263;
  wire       [31:0]   _zz_9264;
  wire       [31:0]   _zz_9265;
  wire       [23:0]   _zz_9266;
  wire       [31:0]   _zz_9267;
  wire       [15:0]   _zz_9268;
  wire       [31:0]   _zz_9269;
  wire       [31:0]   _zz_9270;
  wire       [31:0]   _zz_9271;
  wire       [31:0]   _zz_9272;
  wire       [31:0]   _zz_9273;
  wire       [23:0]   _zz_9274;
  wire       [31:0]   _zz_9275;
  wire       [15:0]   _zz_9276;
  wire       [15:0]   _zz_9277;
  wire       [31:0]   _zz_9278;
  wire       [31:0]   _zz_9279;
  wire       [15:0]   _zz_9280;
  wire       [31:0]   _zz_9281;
  wire       [31:0]   _zz_9282;
  wire       [31:0]   _zz_9283;
  wire       [15:0]   _zz_9284;
  wire       [31:0]   _zz_9285;
  wire       [31:0]   _zz_9286;
  wire       [31:0]   _zz_9287;
  wire       [31:0]   _zz_9288;
  wire       [31:0]   _zz_9289;
  wire       [31:0]   _zz_9290;
  wire       [23:0]   _zz_9291;
  wire       [31:0]   _zz_9292;
  wire       [15:0]   _zz_9293;
  wire       [31:0]   _zz_9294;
  wire       [31:0]   _zz_9295;
  wire       [31:0]   _zz_9296;
  wire       [31:0]   _zz_9297;
  wire       [31:0]   _zz_9298;
  wire       [23:0]   _zz_9299;
  wire       [31:0]   _zz_9300;
  wire       [15:0]   _zz_9301;
  wire       [31:0]   _zz_9302;
  wire       [31:0]   _zz_9303;
  wire       [31:0]   _zz_9304;
  wire       [31:0]   _zz_9305;
  wire       [31:0]   _zz_9306;
  wire       [23:0]   _zz_9307;
  wire       [31:0]   _zz_9308;
  wire       [15:0]   _zz_9309;
  wire       [31:0]   _zz_9310;
  wire       [31:0]   _zz_9311;
  wire       [31:0]   _zz_9312;
  wire       [31:0]   _zz_9313;
  wire       [31:0]   _zz_9314;
  wire       [23:0]   _zz_9315;
  wire       [31:0]   _zz_9316;
  wire       [15:0]   _zz_9317;
  wire       [15:0]   _zz_9318;
  wire       [31:0]   _zz_9319;
  wire       [31:0]   _zz_9320;
  wire       [15:0]   _zz_9321;
  wire       [31:0]   _zz_9322;
  wire       [31:0]   _zz_9323;
  wire       [31:0]   _zz_9324;
  wire       [15:0]   _zz_9325;
  wire       [31:0]   _zz_9326;
  wire       [31:0]   _zz_9327;
  wire       [31:0]   _zz_9328;
  wire       [31:0]   _zz_9329;
  wire       [31:0]   _zz_9330;
  wire       [31:0]   _zz_9331;
  wire       [23:0]   _zz_9332;
  wire       [31:0]   _zz_9333;
  wire       [15:0]   _zz_9334;
  wire       [31:0]   _zz_9335;
  wire       [31:0]   _zz_9336;
  wire       [31:0]   _zz_9337;
  wire       [31:0]   _zz_9338;
  wire       [31:0]   _zz_9339;
  wire       [23:0]   _zz_9340;
  wire       [31:0]   _zz_9341;
  wire       [15:0]   _zz_9342;
  wire       [31:0]   _zz_9343;
  wire       [31:0]   _zz_9344;
  wire       [31:0]   _zz_9345;
  wire       [31:0]   _zz_9346;
  wire       [31:0]   _zz_9347;
  wire       [23:0]   _zz_9348;
  wire       [31:0]   _zz_9349;
  wire       [15:0]   _zz_9350;
  wire       [31:0]   _zz_9351;
  wire       [31:0]   _zz_9352;
  wire       [31:0]   _zz_9353;
  wire       [31:0]   _zz_9354;
  wire       [31:0]   _zz_9355;
  wire       [23:0]   _zz_9356;
  wire       [31:0]   _zz_9357;
  wire       [15:0]   _zz_9358;
  wire       [15:0]   _zz_9359;
  wire       [31:0]   _zz_9360;
  wire       [31:0]   _zz_9361;
  wire       [15:0]   _zz_9362;
  wire       [31:0]   _zz_9363;
  wire       [31:0]   _zz_9364;
  wire       [31:0]   _zz_9365;
  wire       [15:0]   _zz_9366;
  wire       [31:0]   _zz_9367;
  wire       [31:0]   _zz_9368;
  wire       [31:0]   _zz_9369;
  wire       [31:0]   _zz_9370;
  wire       [31:0]   _zz_9371;
  wire       [31:0]   _zz_9372;
  wire       [23:0]   _zz_9373;
  wire       [31:0]   _zz_9374;
  wire       [15:0]   _zz_9375;
  wire       [31:0]   _zz_9376;
  wire       [31:0]   _zz_9377;
  wire       [31:0]   _zz_9378;
  wire       [31:0]   _zz_9379;
  wire       [31:0]   _zz_9380;
  wire       [23:0]   _zz_9381;
  wire       [31:0]   _zz_9382;
  wire       [15:0]   _zz_9383;
  wire       [31:0]   _zz_9384;
  wire       [31:0]   _zz_9385;
  wire       [31:0]   _zz_9386;
  wire       [31:0]   _zz_9387;
  wire       [31:0]   _zz_9388;
  wire       [23:0]   _zz_9389;
  wire       [31:0]   _zz_9390;
  wire       [15:0]   _zz_9391;
  wire       [31:0]   _zz_9392;
  wire       [31:0]   _zz_9393;
  wire       [31:0]   _zz_9394;
  wire       [31:0]   _zz_9395;
  wire       [31:0]   _zz_9396;
  wire       [23:0]   _zz_9397;
  wire       [31:0]   _zz_9398;
  wire       [15:0]   _zz_9399;
  wire       [15:0]   _zz_9400;
  wire       [31:0]   _zz_9401;
  wire       [31:0]   _zz_9402;
  wire       [15:0]   _zz_9403;
  wire       [31:0]   _zz_9404;
  wire       [31:0]   _zz_9405;
  wire       [31:0]   _zz_9406;
  wire       [15:0]   _zz_9407;
  wire       [31:0]   _zz_9408;
  wire       [31:0]   _zz_9409;
  wire       [31:0]   _zz_9410;
  wire       [31:0]   _zz_9411;
  wire       [31:0]   _zz_9412;
  wire       [31:0]   _zz_9413;
  wire       [23:0]   _zz_9414;
  wire       [31:0]   _zz_9415;
  wire       [15:0]   _zz_9416;
  wire       [31:0]   _zz_9417;
  wire       [31:0]   _zz_9418;
  wire       [31:0]   _zz_9419;
  wire       [31:0]   _zz_9420;
  wire       [31:0]   _zz_9421;
  wire       [23:0]   _zz_9422;
  wire       [31:0]   _zz_9423;
  wire       [15:0]   _zz_9424;
  wire       [31:0]   _zz_9425;
  wire       [31:0]   _zz_9426;
  wire       [31:0]   _zz_9427;
  wire       [31:0]   _zz_9428;
  wire       [31:0]   _zz_9429;
  wire       [23:0]   _zz_9430;
  wire       [31:0]   _zz_9431;
  wire       [15:0]   _zz_9432;
  wire       [31:0]   _zz_9433;
  wire       [31:0]   _zz_9434;
  wire       [31:0]   _zz_9435;
  wire       [31:0]   _zz_9436;
  wire       [31:0]   _zz_9437;
  wire       [23:0]   _zz_9438;
  wire       [31:0]   _zz_9439;
  wire       [15:0]   _zz_9440;
  wire       [15:0]   _zz_9441;
  wire       [31:0]   _zz_9442;
  wire       [31:0]   _zz_9443;
  wire       [15:0]   _zz_9444;
  wire       [31:0]   _zz_9445;
  wire       [31:0]   _zz_9446;
  wire       [31:0]   _zz_9447;
  wire       [15:0]   _zz_9448;
  wire       [31:0]   _zz_9449;
  wire       [31:0]   _zz_9450;
  wire       [31:0]   _zz_9451;
  wire       [31:0]   _zz_9452;
  wire       [31:0]   _zz_9453;
  wire       [31:0]   _zz_9454;
  wire       [23:0]   _zz_9455;
  wire       [31:0]   _zz_9456;
  wire       [15:0]   _zz_9457;
  wire       [31:0]   _zz_9458;
  wire       [31:0]   _zz_9459;
  wire       [31:0]   _zz_9460;
  wire       [31:0]   _zz_9461;
  wire       [31:0]   _zz_9462;
  wire       [23:0]   _zz_9463;
  wire       [31:0]   _zz_9464;
  wire       [15:0]   _zz_9465;
  wire       [31:0]   _zz_9466;
  wire       [31:0]   _zz_9467;
  wire       [31:0]   _zz_9468;
  wire       [31:0]   _zz_9469;
  wire       [31:0]   _zz_9470;
  wire       [23:0]   _zz_9471;
  wire       [31:0]   _zz_9472;
  wire       [15:0]   _zz_9473;
  wire       [31:0]   _zz_9474;
  wire       [31:0]   _zz_9475;
  wire       [31:0]   _zz_9476;
  wire       [31:0]   _zz_9477;
  wire       [31:0]   _zz_9478;
  wire       [23:0]   _zz_9479;
  wire       [31:0]   _zz_9480;
  wire       [15:0]   _zz_9481;
  wire       [15:0]   _zz_9482;
  wire       [31:0]   _zz_9483;
  wire       [31:0]   _zz_9484;
  wire       [15:0]   _zz_9485;
  wire       [31:0]   _zz_9486;
  wire       [31:0]   _zz_9487;
  wire       [31:0]   _zz_9488;
  wire       [15:0]   _zz_9489;
  wire       [31:0]   _zz_9490;
  wire       [31:0]   _zz_9491;
  wire       [31:0]   _zz_9492;
  wire       [31:0]   _zz_9493;
  wire       [31:0]   _zz_9494;
  wire       [31:0]   _zz_9495;
  wire       [23:0]   _zz_9496;
  wire       [31:0]   _zz_9497;
  wire       [15:0]   _zz_9498;
  wire       [31:0]   _zz_9499;
  wire       [31:0]   _zz_9500;
  wire       [31:0]   _zz_9501;
  wire       [31:0]   _zz_9502;
  wire       [31:0]   _zz_9503;
  wire       [23:0]   _zz_9504;
  wire       [31:0]   _zz_9505;
  wire       [15:0]   _zz_9506;
  wire       [31:0]   _zz_9507;
  wire       [31:0]   _zz_9508;
  wire       [31:0]   _zz_9509;
  wire       [31:0]   _zz_9510;
  wire       [31:0]   _zz_9511;
  wire       [23:0]   _zz_9512;
  wire       [31:0]   _zz_9513;
  wire       [15:0]   _zz_9514;
  wire       [31:0]   _zz_9515;
  wire       [31:0]   _zz_9516;
  wire       [31:0]   _zz_9517;
  wire       [31:0]   _zz_9518;
  wire       [31:0]   _zz_9519;
  wire       [23:0]   _zz_9520;
  wire       [31:0]   _zz_9521;
  wire       [15:0]   _zz_9522;
  wire       [15:0]   _zz_9523;
  wire       [31:0]   _zz_9524;
  wire       [31:0]   _zz_9525;
  wire       [15:0]   _zz_9526;
  wire       [31:0]   _zz_9527;
  wire       [31:0]   _zz_9528;
  wire       [31:0]   _zz_9529;
  wire       [15:0]   _zz_9530;
  wire       [31:0]   _zz_9531;
  wire       [31:0]   _zz_9532;
  wire       [31:0]   _zz_9533;
  wire       [31:0]   _zz_9534;
  wire       [31:0]   _zz_9535;
  wire       [31:0]   _zz_9536;
  wire       [23:0]   _zz_9537;
  wire       [31:0]   _zz_9538;
  wire       [15:0]   _zz_9539;
  wire       [31:0]   _zz_9540;
  wire       [31:0]   _zz_9541;
  wire       [31:0]   _zz_9542;
  wire       [31:0]   _zz_9543;
  wire       [31:0]   _zz_9544;
  wire       [23:0]   _zz_9545;
  wire       [31:0]   _zz_9546;
  wire       [15:0]   _zz_9547;
  wire       [31:0]   _zz_9548;
  wire       [31:0]   _zz_9549;
  wire       [31:0]   _zz_9550;
  wire       [31:0]   _zz_9551;
  wire       [31:0]   _zz_9552;
  wire       [23:0]   _zz_9553;
  wire       [31:0]   _zz_9554;
  wire       [15:0]   _zz_9555;
  wire       [31:0]   _zz_9556;
  wire       [31:0]   _zz_9557;
  wire       [31:0]   _zz_9558;
  wire       [31:0]   _zz_9559;
  wire       [31:0]   _zz_9560;
  wire       [23:0]   _zz_9561;
  wire       [31:0]   _zz_9562;
  wire       [15:0]   _zz_9563;
  wire       [15:0]   _zz_9564;
  wire       [31:0]   _zz_9565;
  wire       [31:0]   _zz_9566;
  wire       [15:0]   _zz_9567;
  wire       [31:0]   _zz_9568;
  wire       [31:0]   _zz_9569;
  wire       [31:0]   _zz_9570;
  wire       [15:0]   _zz_9571;
  wire       [31:0]   _zz_9572;
  wire       [31:0]   _zz_9573;
  wire       [31:0]   _zz_9574;
  wire       [31:0]   _zz_9575;
  wire       [31:0]   _zz_9576;
  wire       [31:0]   _zz_9577;
  wire       [23:0]   _zz_9578;
  wire       [31:0]   _zz_9579;
  wire       [15:0]   _zz_9580;
  wire       [31:0]   _zz_9581;
  wire       [31:0]   _zz_9582;
  wire       [31:0]   _zz_9583;
  wire       [31:0]   _zz_9584;
  wire       [31:0]   _zz_9585;
  wire       [23:0]   _zz_9586;
  wire       [31:0]   _zz_9587;
  wire       [15:0]   _zz_9588;
  wire       [31:0]   _zz_9589;
  wire       [31:0]   _zz_9590;
  wire       [31:0]   _zz_9591;
  wire       [31:0]   _zz_9592;
  wire       [31:0]   _zz_9593;
  wire       [23:0]   _zz_9594;
  wire       [31:0]   _zz_9595;
  wire       [15:0]   _zz_9596;
  wire       [31:0]   _zz_9597;
  wire       [31:0]   _zz_9598;
  wire       [31:0]   _zz_9599;
  wire       [31:0]   _zz_9600;
  wire       [31:0]   _zz_9601;
  wire       [23:0]   _zz_9602;
  wire       [31:0]   _zz_9603;
  wire       [15:0]   _zz_9604;
  wire       [15:0]   _zz_9605;
  wire       [31:0]   _zz_9606;
  wire       [31:0]   _zz_9607;
  wire       [15:0]   _zz_9608;
  wire       [31:0]   _zz_9609;
  wire       [31:0]   _zz_9610;
  wire       [31:0]   _zz_9611;
  wire       [15:0]   _zz_9612;
  wire       [31:0]   _zz_9613;
  wire       [31:0]   _zz_9614;
  wire       [31:0]   _zz_9615;
  wire       [31:0]   _zz_9616;
  wire       [31:0]   _zz_9617;
  wire       [31:0]   _zz_9618;
  wire       [23:0]   _zz_9619;
  wire       [31:0]   _zz_9620;
  wire       [15:0]   _zz_9621;
  wire       [31:0]   _zz_9622;
  wire       [31:0]   _zz_9623;
  wire       [31:0]   _zz_9624;
  wire       [31:0]   _zz_9625;
  wire       [31:0]   _zz_9626;
  wire       [23:0]   _zz_9627;
  wire       [31:0]   _zz_9628;
  wire       [15:0]   _zz_9629;
  wire       [31:0]   _zz_9630;
  wire       [31:0]   _zz_9631;
  wire       [31:0]   _zz_9632;
  wire       [31:0]   _zz_9633;
  wire       [31:0]   _zz_9634;
  wire       [23:0]   _zz_9635;
  wire       [31:0]   _zz_9636;
  wire       [15:0]   _zz_9637;
  wire       [31:0]   _zz_9638;
  wire       [31:0]   _zz_9639;
  wire       [31:0]   _zz_9640;
  wire       [31:0]   _zz_9641;
  wire       [31:0]   _zz_9642;
  wire       [23:0]   _zz_9643;
  wire       [31:0]   _zz_9644;
  wire       [15:0]   _zz_9645;
  wire       [15:0]   _zz_9646;
  wire       [31:0]   _zz_9647;
  wire       [31:0]   _zz_9648;
  wire       [15:0]   _zz_9649;
  wire       [31:0]   _zz_9650;
  wire       [31:0]   _zz_9651;
  wire       [31:0]   _zz_9652;
  wire       [15:0]   _zz_9653;
  wire       [31:0]   _zz_9654;
  wire       [31:0]   _zz_9655;
  wire       [31:0]   _zz_9656;
  wire       [31:0]   _zz_9657;
  wire       [31:0]   _zz_9658;
  wire       [31:0]   _zz_9659;
  wire       [23:0]   _zz_9660;
  wire       [31:0]   _zz_9661;
  wire       [15:0]   _zz_9662;
  wire       [31:0]   _zz_9663;
  wire       [31:0]   _zz_9664;
  wire       [31:0]   _zz_9665;
  wire       [31:0]   _zz_9666;
  wire       [31:0]   _zz_9667;
  wire       [23:0]   _zz_9668;
  wire       [31:0]   _zz_9669;
  wire       [15:0]   _zz_9670;
  wire       [31:0]   _zz_9671;
  wire       [31:0]   _zz_9672;
  wire       [31:0]   _zz_9673;
  wire       [31:0]   _zz_9674;
  wire       [31:0]   _zz_9675;
  wire       [23:0]   _zz_9676;
  wire       [31:0]   _zz_9677;
  wire       [15:0]   _zz_9678;
  wire       [31:0]   _zz_9679;
  wire       [31:0]   _zz_9680;
  wire       [31:0]   _zz_9681;
  wire       [31:0]   _zz_9682;
  wire       [31:0]   _zz_9683;
  wire       [23:0]   _zz_9684;
  wire       [31:0]   _zz_9685;
  wire       [15:0]   _zz_9686;
  wire       [15:0]   _zz_9687;
  wire       [31:0]   _zz_9688;
  wire       [31:0]   _zz_9689;
  wire       [15:0]   _zz_9690;
  wire       [31:0]   _zz_9691;
  wire       [31:0]   _zz_9692;
  wire       [31:0]   _zz_9693;
  wire       [15:0]   _zz_9694;
  wire       [31:0]   _zz_9695;
  wire       [31:0]   _zz_9696;
  wire       [31:0]   _zz_9697;
  wire       [31:0]   _zz_9698;
  wire       [31:0]   _zz_9699;
  wire       [31:0]   _zz_9700;
  wire       [23:0]   _zz_9701;
  wire       [31:0]   _zz_9702;
  wire       [15:0]   _zz_9703;
  wire       [31:0]   _zz_9704;
  wire       [31:0]   _zz_9705;
  wire       [31:0]   _zz_9706;
  wire       [31:0]   _zz_9707;
  wire       [31:0]   _zz_9708;
  wire       [23:0]   _zz_9709;
  wire       [31:0]   _zz_9710;
  wire       [15:0]   _zz_9711;
  wire       [31:0]   _zz_9712;
  wire       [31:0]   _zz_9713;
  wire       [31:0]   _zz_9714;
  wire       [31:0]   _zz_9715;
  wire       [31:0]   _zz_9716;
  wire       [23:0]   _zz_9717;
  wire       [31:0]   _zz_9718;
  wire       [15:0]   _zz_9719;
  wire       [31:0]   _zz_9720;
  wire       [31:0]   _zz_9721;
  wire       [31:0]   _zz_9722;
  wire       [31:0]   _zz_9723;
  wire       [31:0]   _zz_9724;
  wire       [23:0]   _zz_9725;
  wire       [31:0]   _zz_9726;
  wire       [15:0]   _zz_9727;
  wire       [15:0]   _zz_9728;
  wire       [31:0]   _zz_9729;
  wire       [31:0]   _zz_9730;
  wire       [15:0]   _zz_9731;
  wire       [31:0]   _zz_9732;
  wire       [31:0]   _zz_9733;
  wire       [31:0]   _zz_9734;
  wire       [15:0]   _zz_9735;
  wire       [31:0]   _zz_9736;
  wire       [31:0]   _zz_9737;
  wire       [31:0]   _zz_9738;
  wire       [31:0]   _zz_9739;
  wire       [31:0]   _zz_9740;
  wire       [31:0]   _zz_9741;
  wire       [23:0]   _zz_9742;
  wire       [31:0]   _zz_9743;
  wire       [15:0]   _zz_9744;
  wire       [31:0]   _zz_9745;
  wire       [31:0]   _zz_9746;
  wire       [31:0]   _zz_9747;
  wire       [31:0]   _zz_9748;
  wire       [31:0]   _zz_9749;
  wire       [23:0]   _zz_9750;
  wire       [31:0]   _zz_9751;
  wire       [15:0]   _zz_9752;
  wire       [31:0]   _zz_9753;
  wire       [31:0]   _zz_9754;
  wire       [31:0]   _zz_9755;
  wire       [31:0]   _zz_9756;
  wire       [31:0]   _zz_9757;
  wire       [23:0]   _zz_9758;
  wire       [31:0]   _zz_9759;
  wire       [15:0]   _zz_9760;
  wire       [31:0]   _zz_9761;
  wire       [31:0]   _zz_9762;
  wire       [31:0]   _zz_9763;
  wire       [31:0]   _zz_9764;
  wire       [31:0]   _zz_9765;
  wire       [23:0]   _zz_9766;
  wire       [31:0]   _zz_9767;
  wire       [15:0]   _zz_9768;
  wire       [15:0]   _zz_9769;
  wire       [31:0]   _zz_9770;
  wire       [31:0]   _zz_9771;
  wire       [15:0]   _zz_9772;
  wire       [31:0]   _zz_9773;
  wire       [31:0]   _zz_9774;
  wire       [31:0]   _zz_9775;
  wire       [15:0]   _zz_9776;
  wire       [31:0]   _zz_9777;
  wire       [31:0]   _zz_9778;
  wire       [31:0]   _zz_9779;
  wire       [31:0]   _zz_9780;
  wire       [31:0]   _zz_9781;
  wire       [31:0]   _zz_9782;
  wire       [23:0]   _zz_9783;
  wire       [31:0]   _zz_9784;
  wire       [15:0]   _zz_9785;
  wire       [31:0]   _zz_9786;
  wire       [31:0]   _zz_9787;
  wire       [31:0]   _zz_9788;
  wire       [31:0]   _zz_9789;
  wire       [31:0]   _zz_9790;
  wire       [23:0]   _zz_9791;
  wire       [31:0]   _zz_9792;
  wire       [15:0]   _zz_9793;
  wire       [31:0]   _zz_9794;
  wire       [31:0]   _zz_9795;
  wire       [31:0]   _zz_9796;
  wire       [31:0]   _zz_9797;
  wire       [31:0]   _zz_9798;
  wire       [23:0]   _zz_9799;
  wire       [31:0]   _zz_9800;
  wire       [15:0]   _zz_9801;
  wire       [31:0]   _zz_9802;
  wire       [31:0]   _zz_9803;
  wire       [31:0]   _zz_9804;
  wire       [31:0]   _zz_9805;
  wire       [31:0]   _zz_9806;
  wire       [23:0]   _zz_9807;
  wire       [31:0]   _zz_9808;
  wire       [15:0]   _zz_9809;
  wire       [15:0]   _zz_9810;
  wire       [31:0]   _zz_9811;
  wire       [31:0]   _zz_9812;
  wire       [15:0]   _zz_9813;
  wire       [31:0]   _zz_9814;
  wire       [31:0]   _zz_9815;
  wire       [31:0]   _zz_9816;
  wire       [15:0]   _zz_9817;
  wire       [31:0]   _zz_9818;
  wire       [31:0]   _zz_9819;
  wire       [31:0]   _zz_9820;
  wire       [31:0]   _zz_9821;
  wire       [31:0]   _zz_9822;
  wire       [31:0]   _zz_9823;
  wire       [23:0]   _zz_9824;
  wire       [31:0]   _zz_9825;
  wire       [15:0]   _zz_9826;
  wire       [31:0]   _zz_9827;
  wire       [31:0]   _zz_9828;
  wire       [31:0]   _zz_9829;
  wire       [31:0]   _zz_9830;
  wire       [31:0]   _zz_9831;
  wire       [23:0]   _zz_9832;
  wire       [31:0]   _zz_9833;
  wire       [15:0]   _zz_9834;
  wire       [31:0]   _zz_9835;
  wire       [31:0]   _zz_9836;
  wire       [31:0]   _zz_9837;
  wire       [31:0]   _zz_9838;
  wire       [31:0]   _zz_9839;
  wire       [23:0]   _zz_9840;
  wire       [31:0]   _zz_9841;
  wire       [15:0]   _zz_9842;
  wire       [31:0]   _zz_9843;
  wire       [31:0]   _zz_9844;
  wire       [31:0]   _zz_9845;
  wire       [31:0]   _zz_9846;
  wire       [31:0]   _zz_9847;
  wire       [23:0]   _zz_9848;
  wire       [31:0]   _zz_9849;
  wire       [15:0]   _zz_9850;
  wire       [15:0]   _zz_9851;
  wire       [31:0]   _zz_9852;
  wire       [31:0]   _zz_9853;
  wire       [15:0]   _zz_9854;
  wire       [31:0]   _zz_9855;
  wire       [31:0]   _zz_9856;
  wire       [31:0]   _zz_9857;
  wire       [15:0]   _zz_9858;
  wire       [31:0]   _zz_9859;
  wire       [31:0]   _zz_9860;
  wire       [31:0]   _zz_9861;
  wire       [31:0]   _zz_9862;
  wire       [31:0]   _zz_9863;
  wire       [31:0]   _zz_9864;
  wire       [23:0]   _zz_9865;
  wire       [31:0]   _zz_9866;
  wire       [15:0]   _zz_9867;
  wire       [31:0]   _zz_9868;
  wire       [31:0]   _zz_9869;
  wire       [31:0]   _zz_9870;
  wire       [31:0]   _zz_9871;
  wire       [31:0]   _zz_9872;
  wire       [23:0]   _zz_9873;
  wire       [31:0]   _zz_9874;
  wire       [15:0]   _zz_9875;
  wire       [31:0]   _zz_9876;
  wire       [31:0]   _zz_9877;
  wire       [31:0]   _zz_9878;
  wire       [31:0]   _zz_9879;
  wire       [31:0]   _zz_9880;
  wire       [23:0]   _zz_9881;
  wire       [31:0]   _zz_9882;
  wire       [15:0]   _zz_9883;
  wire       [31:0]   _zz_9884;
  wire       [31:0]   _zz_9885;
  wire       [31:0]   _zz_9886;
  wire       [31:0]   _zz_9887;
  wire       [31:0]   _zz_9888;
  wire       [23:0]   _zz_9889;
  wire       [31:0]   _zz_9890;
  wire       [15:0]   _zz_9891;
  wire       [15:0]   _zz_9892;
  wire       [31:0]   _zz_9893;
  wire       [31:0]   _zz_9894;
  wire       [15:0]   _zz_9895;
  wire       [31:0]   _zz_9896;
  wire       [31:0]   _zz_9897;
  wire       [31:0]   _zz_9898;
  wire       [15:0]   _zz_9899;
  wire       [31:0]   _zz_9900;
  wire       [31:0]   _zz_9901;
  wire       [31:0]   _zz_9902;
  wire       [31:0]   _zz_9903;
  wire       [31:0]   _zz_9904;
  wire       [31:0]   _zz_9905;
  wire       [23:0]   _zz_9906;
  wire       [31:0]   _zz_9907;
  wire       [15:0]   _zz_9908;
  wire       [31:0]   _zz_9909;
  wire       [31:0]   _zz_9910;
  wire       [31:0]   _zz_9911;
  wire       [31:0]   _zz_9912;
  wire       [31:0]   _zz_9913;
  wire       [23:0]   _zz_9914;
  wire       [31:0]   _zz_9915;
  wire       [15:0]   _zz_9916;
  wire       [31:0]   _zz_9917;
  wire       [31:0]   _zz_9918;
  wire       [31:0]   _zz_9919;
  wire       [31:0]   _zz_9920;
  wire       [31:0]   _zz_9921;
  wire       [23:0]   _zz_9922;
  wire       [31:0]   _zz_9923;
  wire       [15:0]   _zz_9924;
  wire       [31:0]   _zz_9925;
  wire       [31:0]   _zz_9926;
  wire       [31:0]   _zz_9927;
  wire       [31:0]   _zz_9928;
  wire       [31:0]   _zz_9929;
  wire       [23:0]   _zz_9930;
  wire       [31:0]   _zz_9931;
  wire       [15:0]   _zz_9932;
  wire       [15:0]   _zz_9933;
  wire       [31:0]   _zz_9934;
  wire       [31:0]   _zz_9935;
  wire       [15:0]   _zz_9936;
  wire       [31:0]   _zz_9937;
  wire       [31:0]   _zz_9938;
  wire       [31:0]   _zz_9939;
  wire       [15:0]   _zz_9940;
  wire       [31:0]   _zz_9941;
  wire       [31:0]   _zz_9942;
  wire       [31:0]   _zz_9943;
  wire       [31:0]   _zz_9944;
  wire       [31:0]   _zz_9945;
  wire       [31:0]   _zz_9946;
  wire       [23:0]   _zz_9947;
  wire       [31:0]   _zz_9948;
  wire       [15:0]   _zz_9949;
  wire       [31:0]   _zz_9950;
  wire       [31:0]   _zz_9951;
  wire       [31:0]   _zz_9952;
  wire       [31:0]   _zz_9953;
  wire       [31:0]   _zz_9954;
  wire       [23:0]   _zz_9955;
  wire       [31:0]   _zz_9956;
  wire       [15:0]   _zz_9957;
  wire       [31:0]   _zz_9958;
  wire       [31:0]   _zz_9959;
  wire       [31:0]   _zz_9960;
  wire       [31:0]   _zz_9961;
  wire       [31:0]   _zz_9962;
  wire       [23:0]   _zz_9963;
  wire       [31:0]   _zz_9964;
  wire       [15:0]   _zz_9965;
  wire       [31:0]   _zz_9966;
  wire       [31:0]   _zz_9967;
  wire       [31:0]   _zz_9968;
  wire       [31:0]   _zz_9969;
  wire       [31:0]   _zz_9970;
  wire       [23:0]   _zz_9971;
  wire       [31:0]   _zz_9972;
  wire       [15:0]   _zz_9973;
  wire       [15:0]   _zz_9974;
  wire       [31:0]   _zz_9975;
  wire       [31:0]   _zz_9976;
  wire       [15:0]   _zz_9977;
  wire       [31:0]   _zz_9978;
  wire       [31:0]   _zz_9979;
  wire       [31:0]   _zz_9980;
  wire       [15:0]   _zz_9981;
  wire       [31:0]   _zz_9982;
  wire       [31:0]   _zz_9983;
  wire       [31:0]   _zz_9984;
  wire       [31:0]   _zz_9985;
  wire       [31:0]   _zz_9986;
  wire       [31:0]   _zz_9987;
  wire       [23:0]   _zz_9988;
  wire       [31:0]   _zz_9989;
  wire       [15:0]   _zz_9990;
  wire       [31:0]   _zz_9991;
  wire       [31:0]   _zz_9992;
  wire       [31:0]   _zz_9993;
  wire       [31:0]   _zz_9994;
  wire       [31:0]   _zz_9995;
  wire       [23:0]   _zz_9996;
  wire       [31:0]   _zz_9997;
  wire       [15:0]   _zz_9998;
  wire       [31:0]   _zz_9999;
  wire       [31:0]   _zz_10000;
  wire       [31:0]   _zz_10001;
  wire       [31:0]   _zz_10002;
  wire       [31:0]   _zz_10003;
  wire       [23:0]   _zz_10004;
  wire       [31:0]   _zz_10005;
  wire       [15:0]   _zz_10006;
  wire       [31:0]   _zz_10007;
  wire       [31:0]   _zz_10008;
  wire       [31:0]   _zz_10009;
  wire       [31:0]   _zz_10010;
  wire       [31:0]   _zz_10011;
  wire       [23:0]   _zz_10012;
  wire       [31:0]   _zz_10013;
  wire       [15:0]   _zz_10014;
  wire       [15:0]   _zz_10015;
  wire       [31:0]   _zz_10016;
  wire       [31:0]   _zz_10017;
  wire       [15:0]   _zz_10018;
  wire       [31:0]   _zz_10019;
  wire       [31:0]   _zz_10020;
  wire       [31:0]   _zz_10021;
  wire       [15:0]   _zz_10022;
  wire       [31:0]   _zz_10023;
  wire       [31:0]   _zz_10024;
  wire       [31:0]   _zz_10025;
  wire       [31:0]   _zz_10026;
  wire       [31:0]   _zz_10027;
  wire       [31:0]   _zz_10028;
  wire       [23:0]   _zz_10029;
  wire       [31:0]   _zz_10030;
  wire       [15:0]   _zz_10031;
  wire       [31:0]   _zz_10032;
  wire       [31:0]   _zz_10033;
  wire       [31:0]   _zz_10034;
  wire       [31:0]   _zz_10035;
  wire       [31:0]   _zz_10036;
  wire       [23:0]   _zz_10037;
  wire       [31:0]   _zz_10038;
  wire       [15:0]   _zz_10039;
  wire       [31:0]   _zz_10040;
  wire       [31:0]   _zz_10041;
  wire       [31:0]   _zz_10042;
  wire       [31:0]   _zz_10043;
  wire       [31:0]   _zz_10044;
  wire       [23:0]   _zz_10045;
  wire       [31:0]   _zz_10046;
  wire       [15:0]   _zz_10047;
  wire       [31:0]   _zz_10048;
  wire       [31:0]   _zz_10049;
  wire       [31:0]   _zz_10050;
  wire       [31:0]   _zz_10051;
  wire       [31:0]   _zz_10052;
  wire       [23:0]   _zz_10053;
  wire       [31:0]   _zz_10054;
  wire       [15:0]   _zz_10055;
  wire       [15:0]   _zz_10056;
  wire       [31:0]   _zz_10057;
  wire       [31:0]   _zz_10058;
  wire       [15:0]   _zz_10059;
  wire       [31:0]   _zz_10060;
  wire       [31:0]   _zz_10061;
  wire       [31:0]   _zz_10062;
  wire       [15:0]   _zz_10063;
  wire       [31:0]   _zz_10064;
  wire       [31:0]   _zz_10065;
  wire       [31:0]   _zz_10066;
  wire       [31:0]   _zz_10067;
  wire       [31:0]   _zz_10068;
  wire       [31:0]   _zz_10069;
  wire       [23:0]   _zz_10070;
  wire       [31:0]   _zz_10071;
  wire       [15:0]   _zz_10072;
  wire       [31:0]   _zz_10073;
  wire       [31:0]   _zz_10074;
  wire       [31:0]   _zz_10075;
  wire       [31:0]   _zz_10076;
  wire       [31:0]   _zz_10077;
  wire       [23:0]   _zz_10078;
  wire       [31:0]   _zz_10079;
  wire       [15:0]   _zz_10080;
  wire       [31:0]   _zz_10081;
  wire       [31:0]   _zz_10082;
  wire       [31:0]   _zz_10083;
  wire       [31:0]   _zz_10084;
  wire       [31:0]   _zz_10085;
  wire       [23:0]   _zz_10086;
  wire       [31:0]   _zz_10087;
  wire       [15:0]   _zz_10088;
  wire       [31:0]   _zz_10089;
  wire       [31:0]   _zz_10090;
  wire       [31:0]   _zz_10091;
  wire       [31:0]   _zz_10092;
  wire       [31:0]   _zz_10093;
  wire       [23:0]   _zz_10094;
  wire       [31:0]   _zz_10095;
  wire       [15:0]   _zz_10096;
  wire       [15:0]   _zz_10097;
  wire       [31:0]   _zz_10098;
  wire       [31:0]   _zz_10099;
  wire       [15:0]   _zz_10100;
  wire       [31:0]   _zz_10101;
  wire       [31:0]   _zz_10102;
  wire       [31:0]   _zz_10103;
  wire       [15:0]   _zz_10104;
  wire       [31:0]   _zz_10105;
  wire       [31:0]   _zz_10106;
  wire       [31:0]   _zz_10107;
  wire       [31:0]   _zz_10108;
  wire       [31:0]   _zz_10109;
  wire       [31:0]   _zz_10110;
  wire       [23:0]   _zz_10111;
  wire       [31:0]   _zz_10112;
  wire       [15:0]   _zz_10113;
  wire       [31:0]   _zz_10114;
  wire       [31:0]   _zz_10115;
  wire       [31:0]   _zz_10116;
  wire       [31:0]   _zz_10117;
  wire       [31:0]   _zz_10118;
  wire       [23:0]   _zz_10119;
  wire       [31:0]   _zz_10120;
  wire       [15:0]   _zz_10121;
  wire       [31:0]   _zz_10122;
  wire       [31:0]   _zz_10123;
  wire       [31:0]   _zz_10124;
  wire       [31:0]   _zz_10125;
  wire       [31:0]   _zz_10126;
  wire       [23:0]   _zz_10127;
  wire       [31:0]   _zz_10128;
  wire       [15:0]   _zz_10129;
  wire       [31:0]   _zz_10130;
  wire       [31:0]   _zz_10131;
  wire       [31:0]   _zz_10132;
  wire       [31:0]   _zz_10133;
  wire       [31:0]   _zz_10134;
  wire       [23:0]   _zz_10135;
  wire       [31:0]   _zz_10136;
  wire       [15:0]   _zz_10137;
  wire       [15:0]   _zz_10138;
  wire       [31:0]   _zz_10139;
  wire       [31:0]   _zz_10140;
  wire       [15:0]   _zz_10141;
  wire       [31:0]   _zz_10142;
  wire       [31:0]   _zz_10143;
  wire       [31:0]   _zz_10144;
  wire       [15:0]   _zz_10145;
  wire       [31:0]   _zz_10146;
  wire       [31:0]   _zz_10147;
  wire       [31:0]   _zz_10148;
  wire       [31:0]   _zz_10149;
  wire       [31:0]   _zz_10150;
  wire       [31:0]   _zz_10151;
  wire       [23:0]   _zz_10152;
  wire       [31:0]   _zz_10153;
  wire       [15:0]   _zz_10154;
  wire       [31:0]   _zz_10155;
  wire       [31:0]   _zz_10156;
  wire       [31:0]   _zz_10157;
  wire       [31:0]   _zz_10158;
  wire       [31:0]   _zz_10159;
  wire       [23:0]   _zz_10160;
  wire       [31:0]   _zz_10161;
  wire       [15:0]   _zz_10162;
  wire       [31:0]   _zz_10163;
  wire       [31:0]   _zz_10164;
  wire       [31:0]   _zz_10165;
  wire       [31:0]   _zz_10166;
  wire       [31:0]   _zz_10167;
  wire       [23:0]   _zz_10168;
  wire       [31:0]   _zz_10169;
  wire       [15:0]   _zz_10170;
  wire       [31:0]   _zz_10171;
  wire       [31:0]   _zz_10172;
  wire       [31:0]   _zz_10173;
  wire       [31:0]   _zz_10174;
  wire       [31:0]   _zz_10175;
  wire       [23:0]   _zz_10176;
  wire       [31:0]   _zz_10177;
  wire       [15:0]   _zz_10178;
  wire       [15:0]   _zz_10179;
  wire       [31:0]   _zz_10180;
  wire       [31:0]   _zz_10181;
  wire       [15:0]   _zz_10182;
  wire       [31:0]   _zz_10183;
  wire       [31:0]   _zz_10184;
  wire       [31:0]   _zz_10185;
  wire       [15:0]   _zz_10186;
  wire       [31:0]   _zz_10187;
  wire       [31:0]   _zz_10188;
  wire       [31:0]   _zz_10189;
  wire       [31:0]   _zz_10190;
  wire       [31:0]   _zz_10191;
  wire       [31:0]   _zz_10192;
  wire       [23:0]   _zz_10193;
  wire       [31:0]   _zz_10194;
  wire       [15:0]   _zz_10195;
  wire       [31:0]   _zz_10196;
  wire       [31:0]   _zz_10197;
  wire       [31:0]   _zz_10198;
  wire       [31:0]   _zz_10199;
  wire       [31:0]   _zz_10200;
  wire       [23:0]   _zz_10201;
  wire       [31:0]   _zz_10202;
  wire       [15:0]   _zz_10203;
  wire       [31:0]   _zz_10204;
  wire       [31:0]   _zz_10205;
  wire       [31:0]   _zz_10206;
  wire       [31:0]   _zz_10207;
  wire       [31:0]   _zz_10208;
  wire       [23:0]   _zz_10209;
  wire       [31:0]   _zz_10210;
  wire       [15:0]   _zz_10211;
  wire       [31:0]   _zz_10212;
  wire       [31:0]   _zz_10213;
  wire       [31:0]   _zz_10214;
  wire       [31:0]   _zz_10215;
  wire       [31:0]   _zz_10216;
  wire       [23:0]   _zz_10217;
  wire       [31:0]   _zz_10218;
  wire       [15:0]   _zz_10219;
  wire       [15:0]   _zz_10220;
  wire       [31:0]   _zz_10221;
  wire       [31:0]   _zz_10222;
  wire       [15:0]   _zz_10223;
  wire       [31:0]   _zz_10224;
  wire       [31:0]   _zz_10225;
  wire       [31:0]   _zz_10226;
  wire       [15:0]   _zz_10227;
  wire       [31:0]   _zz_10228;
  wire       [31:0]   _zz_10229;
  wire       [31:0]   _zz_10230;
  wire       [31:0]   _zz_10231;
  wire       [31:0]   _zz_10232;
  wire       [31:0]   _zz_10233;
  wire       [23:0]   _zz_10234;
  wire       [31:0]   _zz_10235;
  wire       [15:0]   _zz_10236;
  wire       [31:0]   _zz_10237;
  wire       [31:0]   _zz_10238;
  wire       [31:0]   _zz_10239;
  wire       [31:0]   _zz_10240;
  wire       [31:0]   _zz_10241;
  wire       [23:0]   _zz_10242;
  wire       [31:0]   _zz_10243;
  wire       [15:0]   _zz_10244;
  wire       [31:0]   _zz_10245;
  wire       [31:0]   _zz_10246;
  wire       [31:0]   _zz_10247;
  wire       [31:0]   _zz_10248;
  wire       [31:0]   _zz_10249;
  wire       [23:0]   _zz_10250;
  wire       [31:0]   _zz_10251;
  wire       [15:0]   _zz_10252;
  wire       [31:0]   _zz_10253;
  wire       [31:0]   _zz_10254;
  wire       [31:0]   _zz_10255;
  wire       [31:0]   _zz_10256;
  wire       [31:0]   _zz_10257;
  wire       [23:0]   _zz_10258;
  wire       [31:0]   _zz_10259;
  wire       [15:0]   _zz_10260;
  wire       [15:0]   _zz_10261;
  wire       [31:0]   _zz_10262;
  wire       [31:0]   _zz_10263;
  wire       [15:0]   _zz_10264;
  wire       [31:0]   _zz_10265;
  wire       [31:0]   _zz_10266;
  wire       [31:0]   _zz_10267;
  wire       [15:0]   _zz_10268;
  wire       [31:0]   _zz_10269;
  wire       [31:0]   _zz_10270;
  wire       [31:0]   _zz_10271;
  wire       [31:0]   _zz_10272;
  wire       [31:0]   _zz_10273;
  wire       [31:0]   _zz_10274;
  wire       [23:0]   _zz_10275;
  wire       [31:0]   _zz_10276;
  wire       [15:0]   _zz_10277;
  wire       [31:0]   _zz_10278;
  wire       [31:0]   _zz_10279;
  wire       [31:0]   _zz_10280;
  wire       [31:0]   _zz_10281;
  wire       [31:0]   _zz_10282;
  wire       [23:0]   _zz_10283;
  wire       [31:0]   _zz_10284;
  wire       [15:0]   _zz_10285;
  wire       [31:0]   _zz_10286;
  wire       [31:0]   _zz_10287;
  wire       [31:0]   _zz_10288;
  wire       [31:0]   _zz_10289;
  wire       [31:0]   _zz_10290;
  wire       [23:0]   _zz_10291;
  wire       [31:0]   _zz_10292;
  wire       [15:0]   _zz_10293;
  wire       [31:0]   _zz_10294;
  wire       [31:0]   _zz_10295;
  wire       [31:0]   _zz_10296;
  wire       [31:0]   _zz_10297;
  wire       [31:0]   _zz_10298;
  wire       [23:0]   _zz_10299;
  wire       [31:0]   _zz_10300;
  wire       [15:0]   _zz_10301;
  wire       [15:0]   _zz_10302;
  wire       [31:0]   _zz_10303;
  wire       [31:0]   _zz_10304;
  wire       [15:0]   _zz_10305;
  wire       [31:0]   _zz_10306;
  wire       [31:0]   _zz_10307;
  wire       [31:0]   _zz_10308;
  wire       [15:0]   _zz_10309;
  wire       [31:0]   _zz_10310;
  wire       [31:0]   _zz_10311;
  wire       [31:0]   _zz_10312;
  wire       [31:0]   _zz_10313;
  wire       [31:0]   _zz_10314;
  wire       [31:0]   _zz_10315;
  wire       [23:0]   _zz_10316;
  wire       [31:0]   _zz_10317;
  wire       [15:0]   _zz_10318;
  wire       [31:0]   _zz_10319;
  wire       [31:0]   _zz_10320;
  wire       [31:0]   _zz_10321;
  wire       [31:0]   _zz_10322;
  wire       [31:0]   _zz_10323;
  wire       [23:0]   _zz_10324;
  wire       [31:0]   _zz_10325;
  wire       [15:0]   _zz_10326;
  wire       [31:0]   _zz_10327;
  wire       [31:0]   _zz_10328;
  wire       [31:0]   _zz_10329;
  wire       [31:0]   _zz_10330;
  wire       [31:0]   _zz_10331;
  wire       [23:0]   _zz_10332;
  wire       [31:0]   _zz_10333;
  wire       [15:0]   _zz_10334;
  wire       [31:0]   _zz_10335;
  wire       [31:0]   _zz_10336;
  wire       [31:0]   _zz_10337;
  wire       [31:0]   _zz_10338;
  wire       [31:0]   _zz_10339;
  wire       [23:0]   _zz_10340;
  wire       [31:0]   _zz_10341;
  wire       [15:0]   _zz_10342;
  wire       [15:0]   _zz_10343;
  wire       [31:0]   _zz_10344;
  wire       [31:0]   _zz_10345;
  wire       [15:0]   _zz_10346;
  wire       [31:0]   _zz_10347;
  wire       [31:0]   _zz_10348;
  wire       [31:0]   _zz_10349;
  wire       [15:0]   _zz_10350;
  wire       [31:0]   _zz_10351;
  wire       [31:0]   _zz_10352;
  wire       [31:0]   _zz_10353;
  wire       [31:0]   _zz_10354;
  wire       [31:0]   _zz_10355;
  wire       [31:0]   _zz_10356;
  wire       [23:0]   _zz_10357;
  wire       [31:0]   _zz_10358;
  wire       [15:0]   _zz_10359;
  wire       [31:0]   _zz_10360;
  wire       [31:0]   _zz_10361;
  wire       [31:0]   _zz_10362;
  wire       [31:0]   _zz_10363;
  wire       [31:0]   _zz_10364;
  wire       [23:0]   _zz_10365;
  wire       [31:0]   _zz_10366;
  wire       [15:0]   _zz_10367;
  wire       [31:0]   _zz_10368;
  wire       [31:0]   _zz_10369;
  wire       [31:0]   _zz_10370;
  wire       [31:0]   _zz_10371;
  wire       [31:0]   _zz_10372;
  wire       [23:0]   _zz_10373;
  wire       [31:0]   _zz_10374;
  wire       [15:0]   _zz_10375;
  wire       [31:0]   _zz_10376;
  wire       [31:0]   _zz_10377;
  wire       [31:0]   _zz_10378;
  wire       [31:0]   _zz_10379;
  wire       [31:0]   _zz_10380;
  wire       [23:0]   _zz_10381;
  wire       [31:0]   _zz_10382;
  wire       [15:0]   _zz_10383;
  wire       [15:0]   _zz_10384;
  wire       [31:0]   _zz_10385;
  wire       [31:0]   _zz_10386;
  wire       [15:0]   _zz_10387;
  wire       [31:0]   _zz_10388;
  wire       [31:0]   _zz_10389;
  wire       [31:0]   _zz_10390;
  wire       [15:0]   _zz_10391;
  wire       [31:0]   _zz_10392;
  wire       [31:0]   _zz_10393;
  wire       [31:0]   _zz_10394;
  wire       [31:0]   _zz_10395;
  wire       [31:0]   _zz_10396;
  wire       [31:0]   _zz_10397;
  wire       [23:0]   _zz_10398;
  wire       [31:0]   _zz_10399;
  wire       [15:0]   _zz_10400;
  wire       [31:0]   _zz_10401;
  wire       [31:0]   _zz_10402;
  wire       [31:0]   _zz_10403;
  wire       [31:0]   _zz_10404;
  wire       [31:0]   _zz_10405;
  wire       [23:0]   _zz_10406;
  wire       [31:0]   _zz_10407;
  wire       [15:0]   _zz_10408;
  wire       [31:0]   _zz_10409;
  wire       [31:0]   _zz_10410;
  wire       [31:0]   _zz_10411;
  wire       [31:0]   _zz_10412;
  wire       [31:0]   _zz_10413;
  wire       [23:0]   _zz_10414;
  wire       [31:0]   _zz_10415;
  wire       [15:0]   _zz_10416;
  wire       [31:0]   _zz_10417;
  wire       [31:0]   _zz_10418;
  wire       [31:0]   _zz_10419;
  wire       [31:0]   _zz_10420;
  wire       [31:0]   _zz_10421;
  wire       [23:0]   _zz_10422;
  wire       [31:0]   _zz_10423;
  wire       [15:0]   _zz_10424;
  wire       [15:0]   _zz_10425;
  wire       [31:0]   _zz_10426;
  wire       [31:0]   _zz_10427;
  wire       [15:0]   _zz_10428;
  wire       [31:0]   _zz_10429;
  wire       [31:0]   _zz_10430;
  wire       [31:0]   _zz_10431;
  wire       [15:0]   _zz_10432;
  wire       [31:0]   _zz_10433;
  wire       [31:0]   _zz_10434;
  wire       [31:0]   _zz_10435;
  wire       [31:0]   _zz_10436;
  wire       [31:0]   _zz_10437;
  wire       [31:0]   _zz_10438;
  wire       [23:0]   _zz_10439;
  wire       [31:0]   _zz_10440;
  wire       [15:0]   _zz_10441;
  wire       [31:0]   _zz_10442;
  wire       [31:0]   _zz_10443;
  wire       [31:0]   _zz_10444;
  wire       [31:0]   _zz_10445;
  wire       [31:0]   _zz_10446;
  wire       [23:0]   _zz_10447;
  wire       [31:0]   _zz_10448;
  wire       [15:0]   _zz_10449;
  wire       [31:0]   _zz_10450;
  wire       [31:0]   _zz_10451;
  wire       [31:0]   _zz_10452;
  wire       [31:0]   _zz_10453;
  wire       [31:0]   _zz_10454;
  wire       [23:0]   _zz_10455;
  wire       [31:0]   _zz_10456;
  wire       [15:0]   _zz_10457;
  wire       [31:0]   _zz_10458;
  wire       [31:0]   _zz_10459;
  wire       [31:0]   _zz_10460;
  wire       [31:0]   _zz_10461;
  wire       [31:0]   _zz_10462;
  wire       [23:0]   _zz_10463;
  wire       [31:0]   _zz_10464;
  wire       [15:0]   _zz_10465;
  wire       [15:0]   _zz_10466;
  wire       [31:0]   _zz_10467;
  wire       [31:0]   _zz_10468;
  wire       [15:0]   _zz_10469;
  wire       [31:0]   _zz_10470;
  wire       [31:0]   _zz_10471;
  wire       [31:0]   _zz_10472;
  wire       [15:0]   _zz_10473;
  wire       [31:0]   _zz_10474;
  wire       [31:0]   _zz_10475;
  wire       [31:0]   _zz_10476;
  wire       [31:0]   _zz_10477;
  wire       [31:0]   _zz_10478;
  wire       [31:0]   _zz_10479;
  wire       [23:0]   _zz_10480;
  wire       [31:0]   _zz_10481;
  wire       [15:0]   _zz_10482;
  wire       [31:0]   _zz_10483;
  wire       [31:0]   _zz_10484;
  wire       [31:0]   _zz_10485;
  wire       [31:0]   _zz_10486;
  wire       [31:0]   _zz_10487;
  wire       [23:0]   _zz_10488;
  wire       [31:0]   _zz_10489;
  wire       [15:0]   _zz_10490;
  wire       [31:0]   _zz_10491;
  wire       [31:0]   _zz_10492;
  wire       [31:0]   _zz_10493;
  wire       [31:0]   _zz_10494;
  wire       [31:0]   _zz_10495;
  wire       [23:0]   _zz_10496;
  wire       [31:0]   _zz_10497;
  wire       [15:0]   _zz_10498;
  wire       [31:0]   _zz_10499;
  wire       [31:0]   _zz_10500;
  wire       [31:0]   _zz_10501;
  wire       [31:0]   _zz_10502;
  wire       [31:0]   _zz_10503;
  wire       [23:0]   _zz_10504;
  wire       [31:0]   _zz_10505;
  wire       [15:0]   _zz_10506;
  wire       [15:0]   _zz_10507;
  wire       [31:0]   _zz_10508;
  wire       [31:0]   _zz_10509;
  wire       [15:0]   _zz_10510;
  wire       [31:0]   _zz_10511;
  wire       [31:0]   _zz_10512;
  wire       [31:0]   _zz_10513;
  wire       [15:0]   _zz_10514;
  wire       [31:0]   _zz_10515;
  wire       [31:0]   _zz_10516;
  wire       [31:0]   _zz_10517;
  wire       [31:0]   _zz_10518;
  wire       [31:0]   _zz_10519;
  wire       [31:0]   _zz_10520;
  wire       [23:0]   _zz_10521;
  wire       [31:0]   _zz_10522;
  wire       [15:0]   _zz_10523;
  wire       [31:0]   _zz_10524;
  wire       [31:0]   _zz_10525;
  wire       [31:0]   _zz_10526;
  wire       [31:0]   _zz_10527;
  wire       [31:0]   _zz_10528;
  wire       [23:0]   _zz_10529;
  wire       [31:0]   _zz_10530;
  wire       [15:0]   _zz_10531;
  wire       [31:0]   _zz_10532;
  wire       [31:0]   _zz_10533;
  wire       [31:0]   _zz_10534;
  wire       [31:0]   _zz_10535;
  wire       [31:0]   _zz_10536;
  wire       [23:0]   _zz_10537;
  wire       [31:0]   _zz_10538;
  wire       [15:0]   _zz_10539;
  wire       [31:0]   _zz_10540;
  wire       [31:0]   _zz_10541;
  wire       [31:0]   _zz_10542;
  wire       [31:0]   _zz_10543;
  wire       [31:0]   _zz_10544;
  wire       [23:0]   _zz_10545;
  wire       [31:0]   _zz_10546;
  wire       [15:0]   _zz_10547;
  wire       [15:0]   _zz_10548;
  wire       [31:0]   _zz_10549;
  wire       [31:0]   _zz_10550;
  wire       [15:0]   _zz_10551;
  wire       [31:0]   _zz_10552;
  wire       [31:0]   _zz_10553;
  wire       [31:0]   _zz_10554;
  wire       [15:0]   _zz_10555;
  wire       [31:0]   _zz_10556;
  wire       [31:0]   _zz_10557;
  wire       [31:0]   _zz_10558;
  wire       [31:0]   _zz_10559;
  wire       [31:0]   _zz_10560;
  wire       [31:0]   _zz_10561;
  wire       [23:0]   _zz_10562;
  wire       [31:0]   _zz_10563;
  wire       [15:0]   _zz_10564;
  wire       [31:0]   _zz_10565;
  wire       [31:0]   _zz_10566;
  wire       [31:0]   _zz_10567;
  wire       [31:0]   _zz_10568;
  wire       [31:0]   _zz_10569;
  wire       [23:0]   _zz_10570;
  wire       [31:0]   _zz_10571;
  wire       [15:0]   _zz_10572;
  wire       [31:0]   _zz_10573;
  wire       [31:0]   _zz_10574;
  wire       [31:0]   _zz_10575;
  wire       [31:0]   _zz_10576;
  wire       [31:0]   _zz_10577;
  wire       [23:0]   _zz_10578;
  wire       [31:0]   _zz_10579;
  wire       [15:0]   _zz_10580;
  wire       [31:0]   _zz_10581;
  wire       [31:0]   _zz_10582;
  wire       [31:0]   _zz_10583;
  wire       [31:0]   _zz_10584;
  wire       [31:0]   _zz_10585;
  wire       [23:0]   _zz_10586;
  wire       [31:0]   _zz_10587;
  wire       [15:0]   _zz_10588;
  wire       [15:0]   _zz_10589;
  wire       [31:0]   _zz_10590;
  wire       [31:0]   _zz_10591;
  wire       [15:0]   _zz_10592;
  wire       [31:0]   _zz_10593;
  wire       [31:0]   _zz_10594;
  wire       [31:0]   _zz_10595;
  wire       [15:0]   _zz_10596;
  wire       [31:0]   _zz_10597;
  wire       [31:0]   _zz_10598;
  wire       [31:0]   _zz_10599;
  wire       [31:0]   _zz_10600;
  wire       [31:0]   _zz_10601;
  wire       [31:0]   _zz_10602;
  wire       [23:0]   _zz_10603;
  wire       [31:0]   _zz_10604;
  wire       [15:0]   _zz_10605;
  wire       [31:0]   _zz_10606;
  wire       [31:0]   _zz_10607;
  wire       [31:0]   _zz_10608;
  wire       [31:0]   _zz_10609;
  wire       [31:0]   _zz_10610;
  wire       [23:0]   _zz_10611;
  wire       [31:0]   _zz_10612;
  wire       [15:0]   _zz_10613;
  wire       [31:0]   _zz_10614;
  wire       [31:0]   _zz_10615;
  wire       [31:0]   _zz_10616;
  wire       [31:0]   _zz_10617;
  wire       [31:0]   _zz_10618;
  wire       [23:0]   _zz_10619;
  wire       [31:0]   _zz_10620;
  wire       [15:0]   _zz_10621;
  wire       [31:0]   _zz_10622;
  wire       [31:0]   _zz_10623;
  wire       [31:0]   _zz_10624;
  wire       [31:0]   _zz_10625;
  wire       [31:0]   _zz_10626;
  wire       [23:0]   _zz_10627;
  wire       [31:0]   _zz_10628;
  wire       [15:0]   _zz_10629;
  wire       [15:0]   _zz_10630;
  wire       [31:0]   _zz_10631;
  wire       [31:0]   _zz_10632;
  wire       [15:0]   _zz_10633;
  wire       [31:0]   _zz_10634;
  wire       [31:0]   _zz_10635;
  wire       [31:0]   _zz_10636;
  wire       [15:0]   _zz_10637;
  wire       [31:0]   _zz_10638;
  wire       [31:0]   _zz_10639;
  wire       [31:0]   _zz_10640;
  wire       [31:0]   _zz_10641;
  wire       [31:0]   _zz_10642;
  wire       [31:0]   _zz_10643;
  wire       [23:0]   _zz_10644;
  wire       [31:0]   _zz_10645;
  wire       [15:0]   _zz_10646;
  wire       [31:0]   _zz_10647;
  wire       [31:0]   _zz_10648;
  wire       [31:0]   _zz_10649;
  wire       [31:0]   _zz_10650;
  wire       [31:0]   _zz_10651;
  wire       [23:0]   _zz_10652;
  wire       [31:0]   _zz_10653;
  wire       [15:0]   _zz_10654;
  wire       [31:0]   _zz_10655;
  wire       [31:0]   _zz_10656;
  wire       [31:0]   _zz_10657;
  wire       [31:0]   _zz_10658;
  wire       [31:0]   _zz_10659;
  wire       [23:0]   _zz_10660;
  wire       [31:0]   _zz_10661;
  wire       [15:0]   _zz_10662;
  wire       [31:0]   _zz_10663;
  wire       [31:0]   _zz_10664;
  wire       [31:0]   _zz_10665;
  wire       [31:0]   _zz_10666;
  wire       [31:0]   _zz_10667;
  wire       [23:0]   _zz_10668;
  wire       [31:0]   _zz_10669;
  wire       [15:0]   _zz_10670;
  wire       [15:0]   _zz_10671;
  wire       [31:0]   _zz_10672;
  wire       [31:0]   _zz_10673;
  wire       [15:0]   _zz_10674;
  wire       [31:0]   _zz_10675;
  wire       [31:0]   _zz_10676;
  wire       [31:0]   _zz_10677;
  wire       [15:0]   _zz_10678;
  wire       [31:0]   _zz_10679;
  wire       [31:0]   _zz_10680;
  wire       [31:0]   _zz_10681;
  wire       [31:0]   _zz_10682;
  wire       [31:0]   _zz_10683;
  wire       [31:0]   _zz_10684;
  wire       [23:0]   _zz_10685;
  wire       [31:0]   _zz_10686;
  wire       [15:0]   _zz_10687;
  wire       [31:0]   _zz_10688;
  wire       [31:0]   _zz_10689;
  wire       [31:0]   _zz_10690;
  wire       [31:0]   _zz_10691;
  wire       [31:0]   _zz_10692;
  wire       [23:0]   _zz_10693;
  wire       [31:0]   _zz_10694;
  wire       [15:0]   _zz_10695;
  wire       [31:0]   _zz_10696;
  wire       [31:0]   _zz_10697;
  wire       [31:0]   _zz_10698;
  wire       [31:0]   _zz_10699;
  wire       [31:0]   _zz_10700;
  wire       [23:0]   _zz_10701;
  wire       [31:0]   _zz_10702;
  wire       [15:0]   _zz_10703;
  wire       [31:0]   _zz_10704;
  wire       [31:0]   _zz_10705;
  wire       [31:0]   _zz_10706;
  wire       [31:0]   _zz_10707;
  wire       [31:0]   _zz_10708;
  wire       [23:0]   _zz_10709;
  wire       [31:0]   _zz_10710;
  wire       [15:0]   _zz_10711;
  wire       [15:0]   _zz_10712;
  wire       [31:0]   _zz_10713;
  wire       [31:0]   _zz_10714;
  wire       [15:0]   _zz_10715;
  wire       [31:0]   _zz_10716;
  wire       [31:0]   _zz_10717;
  wire       [31:0]   _zz_10718;
  wire       [15:0]   _zz_10719;
  wire       [31:0]   _zz_10720;
  wire       [31:0]   _zz_10721;
  wire       [31:0]   _zz_10722;
  wire       [31:0]   _zz_10723;
  wire       [31:0]   _zz_10724;
  wire       [31:0]   _zz_10725;
  wire       [23:0]   _zz_10726;
  wire       [31:0]   _zz_10727;
  wire       [15:0]   _zz_10728;
  wire       [31:0]   _zz_10729;
  wire       [31:0]   _zz_10730;
  wire       [31:0]   _zz_10731;
  wire       [31:0]   _zz_10732;
  wire       [31:0]   _zz_10733;
  wire       [23:0]   _zz_10734;
  wire       [31:0]   _zz_10735;
  wire       [15:0]   _zz_10736;
  wire       [31:0]   _zz_10737;
  wire       [31:0]   _zz_10738;
  wire       [31:0]   _zz_10739;
  wire       [31:0]   _zz_10740;
  wire       [31:0]   _zz_10741;
  wire       [23:0]   _zz_10742;
  wire       [31:0]   _zz_10743;
  wire       [15:0]   _zz_10744;
  wire       [31:0]   _zz_10745;
  wire       [31:0]   _zz_10746;
  wire       [31:0]   _zz_10747;
  wire       [31:0]   _zz_10748;
  wire       [31:0]   _zz_10749;
  wire       [23:0]   _zz_10750;
  wire       [31:0]   _zz_10751;
  wire       [15:0]   _zz_10752;
  wire       [15:0]   _zz_10753;
  wire       [31:0]   _zz_10754;
  wire       [31:0]   _zz_10755;
  wire       [15:0]   _zz_10756;
  wire       [31:0]   _zz_10757;
  wire       [31:0]   _zz_10758;
  wire       [31:0]   _zz_10759;
  wire       [15:0]   _zz_10760;
  wire       [31:0]   _zz_10761;
  wire       [31:0]   _zz_10762;
  wire       [31:0]   _zz_10763;
  wire       [31:0]   _zz_10764;
  wire       [31:0]   _zz_10765;
  wire       [31:0]   _zz_10766;
  wire       [23:0]   _zz_10767;
  wire       [31:0]   _zz_10768;
  wire       [15:0]   _zz_10769;
  wire       [31:0]   _zz_10770;
  wire       [31:0]   _zz_10771;
  wire       [31:0]   _zz_10772;
  wire       [31:0]   _zz_10773;
  wire       [31:0]   _zz_10774;
  wire       [23:0]   _zz_10775;
  wire       [31:0]   _zz_10776;
  wire       [15:0]   _zz_10777;
  wire       [31:0]   _zz_10778;
  wire       [31:0]   _zz_10779;
  wire       [31:0]   _zz_10780;
  wire       [31:0]   _zz_10781;
  wire       [31:0]   _zz_10782;
  wire       [23:0]   _zz_10783;
  wire       [31:0]   _zz_10784;
  wire       [15:0]   _zz_10785;
  wire       [31:0]   _zz_10786;
  wire       [31:0]   _zz_10787;
  wire       [31:0]   _zz_10788;
  wire       [31:0]   _zz_10789;
  wire       [31:0]   _zz_10790;
  wire       [23:0]   _zz_10791;
  wire       [31:0]   _zz_10792;
  wire       [15:0]   _zz_10793;
  wire       [15:0]   _zz_10794;
  wire       [31:0]   _zz_10795;
  wire       [31:0]   _zz_10796;
  wire       [15:0]   _zz_10797;
  wire       [31:0]   _zz_10798;
  wire       [31:0]   _zz_10799;
  wire       [31:0]   _zz_10800;
  wire       [15:0]   _zz_10801;
  wire       [31:0]   _zz_10802;
  wire       [31:0]   _zz_10803;
  wire       [31:0]   _zz_10804;
  wire       [31:0]   _zz_10805;
  wire       [31:0]   _zz_10806;
  wire       [31:0]   _zz_10807;
  wire       [23:0]   _zz_10808;
  wire       [31:0]   _zz_10809;
  wire       [15:0]   _zz_10810;
  wire       [31:0]   _zz_10811;
  wire       [31:0]   _zz_10812;
  wire       [31:0]   _zz_10813;
  wire       [31:0]   _zz_10814;
  wire       [31:0]   _zz_10815;
  wire       [23:0]   _zz_10816;
  wire       [31:0]   _zz_10817;
  wire       [15:0]   _zz_10818;
  wire       [31:0]   _zz_10819;
  wire       [31:0]   _zz_10820;
  wire       [31:0]   _zz_10821;
  wire       [31:0]   _zz_10822;
  wire       [31:0]   _zz_10823;
  wire       [23:0]   _zz_10824;
  wire       [31:0]   _zz_10825;
  wire       [15:0]   _zz_10826;
  wire       [31:0]   _zz_10827;
  wire       [31:0]   _zz_10828;
  wire       [31:0]   _zz_10829;
  wire       [31:0]   _zz_10830;
  wire       [31:0]   _zz_10831;
  wire       [23:0]   _zz_10832;
  wire       [31:0]   _zz_10833;
  wire       [15:0]   _zz_10834;
  wire       [15:0]   _zz_10835;
  wire       [31:0]   _zz_10836;
  wire       [31:0]   _zz_10837;
  wire       [15:0]   _zz_10838;
  wire       [31:0]   _zz_10839;
  wire       [31:0]   _zz_10840;
  wire       [31:0]   _zz_10841;
  wire       [15:0]   _zz_10842;
  wire       [31:0]   _zz_10843;
  wire       [31:0]   _zz_10844;
  wire       [31:0]   _zz_10845;
  wire       [31:0]   _zz_10846;
  wire       [31:0]   _zz_10847;
  wire       [31:0]   _zz_10848;
  wire       [23:0]   _zz_10849;
  wire       [31:0]   _zz_10850;
  wire       [15:0]   _zz_10851;
  wire       [31:0]   _zz_10852;
  wire       [31:0]   _zz_10853;
  wire       [31:0]   _zz_10854;
  wire       [31:0]   _zz_10855;
  wire       [31:0]   _zz_10856;
  wire       [23:0]   _zz_10857;
  wire       [31:0]   _zz_10858;
  wire       [15:0]   _zz_10859;
  wire       [31:0]   _zz_10860;
  wire       [31:0]   _zz_10861;
  wire       [31:0]   _zz_10862;
  wire       [31:0]   _zz_10863;
  wire       [31:0]   _zz_10864;
  wire       [23:0]   _zz_10865;
  wire       [31:0]   _zz_10866;
  wire       [15:0]   _zz_10867;
  wire       [31:0]   _zz_10868;
  wire       [31:0]   _zz_10869;
  wire       [31:0]   _zz_10870;
  wire       [31:0]   _zz_10871;
  wire       [31:0]   _zz_10872;
  wire       [23:0]   _zz_10873;
  wire       [31:0]   _zz_10874;
  wire       [15:0]   _zz_10875;
  wire       [15:0]   _zz_10876;
  wire       [31:0]   _zz_10877;
  wire       [31:0]   _zz_10878;
  wire       [15:0]   _zz_10879;
  wire       [31:0]   _zz_10880;
  wire       [31:0]   _zz_10881;
  wire       [31:0]   _zz_10882;
  wire       [15:0]   _zz_10883;
  wire       [31:0]   _zz_10884;
  wire       [31:0]   _zz_10885;
  wire       [31:0]   _zz_10886;
  wire       [31:0]   _zz_10887;
  wire       [31:0]   _zz_10888;
  wire       [31:0]   _zz_10889;
  wire       [23:0]   _zz_10890;
  wire       [31:0]   _zz_10891;
  wire       [15:0]   _zz_10892;
  wire       [31:0]   _zz_10893;
  wire       [31:0]   _zz_10894;
  wire       [31:0]   _zz_10895;
  wire       [31:0]   _zz_10896;
  wire       [31:0]   _zz_10897;
  wire       [23:0]   _zz_10898;
  wire       [31:0]   _zz_10899;
  wire       [15:0]   _zz_10900;
  wire       [31:0]   _zz_10901;
  wire       [31:0]   _zz_10902;
  wire       [31:0]   _zz_10903;
  wire       [31:0]   _zz_10904;
  wire       [31:0]   _zz_10905;
  wire       [23:0]   _zz_10906;
  wire       [31:0]   _zz_10907;
  wire       [15:0]   _zz_10908;
  wire       [31:0]   _zz_10909;
  wire       [31:0]   _zz_10910;
  wire       [31:0]   _zz_10911;
  wire       [31:0]   _zz_10912;
  wire       [31:0]   _zz_10913;
  wire       [23:0]   _zz_10914;
  wire       [31:0]   _zz_10915;
  wire       [15:0]   _zz_10916;
  wire       [15:0]   _zz_10917;
  wire       [31:0]   _zz_10918;
  wire       [31:0]   _zz_10919;
  wire       [15:0]   _zz_10920;
  wire       [31:0]   _zz_10921;
  wire       [31:0]   _zz_10922;
  wire       [31:0]   _zz_10923;
  wire       [15:0]   _zz_10924;
  wire       [31:0]   _zz_10925;
  wire       [31:0]   _zz_10926;
  wire       [31:0]   _zz_10927;
  wire       [31:0]   _zz_10928;
  wire       [31:0]   _zz_10929;
  wire       [31:0]   _zz_10930;
  wire       [23:0]   _zz_10931;
  wire       [31:0]   _zz_10932;
  wire       [15:0]   _zz_10933;
  wire       [31:0]   _zz_10934;
  wire       [31:0]   _zz_10935;
  wire       [31:0]   _zz_10936;
  wire       [31:0]   _zz_10937;
  wire       [31:0]   _zz_10938;
  wire       [23:0]   _zz_10939;
  wire       [31:0]   _zz_10940;
  wire       [15:0]   _zz_10941;
  wire       [31:0]   _zz_10942;
  wire       [31:0]   _zz_10943;
  wire       [31:0]   _zz_10944;
  wire       [31:0]   _zz_10945;
  wire       [31:0]   _zz_10946;
  wire       [23:0]   _zz_10947;
  wire       [31:0]   _zz_10948;
  wire       [15:0]   _zz_10949;
  wire       [31:0]   _zz_10950;
  wire       [31:0]   _zz_10951;
  wire       [31:0]   _zz_10952;
  wire       [31:0]   _zz_10953;
  wire       [31:0]   _zz_10954;
  wire       [23:0]   _zz_10955;
  wire       [31:0]   _zz_10956;
  wire       [15:0]   _zz_10957;
  wire       [15:0]   _zz_10958;
  wire       [31:0]   _zz_10959;
  wire       [31:0]   _zz_10960;
  wire       [15:0]   _zz_10961;
  wire       [31:0]   _zz_10962;
  wire       [31:0]   _zz_10963;
  wire       [31:0]   _zz_10964;
  wire       [15:0]   _zz_10965;
  wire       [31:0]   _zz_10966;
  wire       [31:0]   _zz_10967;
  wire       [31:0]   _zz_10968;
  wire       [31:0]   _zz_10969;
  wire       [31:0]   _zz_10970;
  wire       [31:0]   _zz_10971;
  wire       [23:0]   _zz_10972;
  wire       [31:0]   _zz_10973;
  wire       [15:0]   _zz_10974;
  wire       [31:0]   _zz_10975;
  wire       [31:0]   _zz_10976;
  wire       [31:0]   _zz_10977;
  wire       [31:0]   _zz_10978;
  wire       [31:0]   _zz_10979;
  wire       [23:0]   _zz_10980;
  wire       [31:0]   _zz_10981;
  wire       [15:0]   _zz_10982;
  wire       [31:0]   _zz_10983;
  wire       [31:0]   _zz_10984;
  wire       [31:0]   _zz_10985;
  wire       [31:0]   _zz_10986;
  wire       [31:0]   _zz_10987;
  wire       [23:0]   _zz_10988;
  wire       [31:0]   _zz_10989;
  wire       [15:0]   _zz_10990;
  wire       [31:0]   _zz_10991;
  wire       [31:0]   _zz_10992;
  wire       [31:0]   _zz_10993;
  wire       [31:0]   _zz_10994;
  wire       [31:0]   _zz_10995;
  wire       [23:0]   _zz_10996;
  wire       [31:0]   _zz_10997;
  wire       [15:0]   _zz_10998;
  wire       [15:0]   _zz_10999;
  wire       [31:0]   _zz_11000;
  wire       [31:0]   _zz_11001;
  wire       [15:0]   _zz_11002;
  wire       [31:0]   _zz_11003;
  wire       [31:0]   _zz_11004;
  wire       [31:0]   _zz_11005;
  wire       [15:0]   _zz_11006;
  wire       [31:0]   _zz_11007;
  wire       [31:0]   _zz_11008;
  wire       [31:0]   _zz_11009;
  wire       [31:0]   _zz_11010;
  wire       [31:0]   _zz_11011;
  wire       [31:0]   _zz_11012;
  wire       [23:0]   _zz_11013;
  wire       [31:0]   _zz_11014;
  wire       [15:0]   _zz_11015;
  wire       [31:0]   _zz_11016;
  wire       [31:0]   _zz_11017;
  wire       [31:0]   _zz_11018;
  wire       [31:0]   _zz_11019;
  wire       [31:0]   _zz_11020;
  wire       [23:0]   _zz_11021;
  wire       [31:0]   _zz_11022;
  wire       [15:0]   _zz_11023;
  wire       [31:0]   _zz_11024;
  wire       [31:0]   _zz_11025;
  wire       [31:0]   _zz_11026;
  wire       [31:0]   _zz_11027;
  wire       [31:0]   _zz_11028;
  wire       [23:0]   _zz_11029;
  wire       [31:0]   _zz_11030;
  wire       [15:0]   _zz_11031;
  wire       [31:0]   _zz_11032;
  wire       [31:0]   _zz_11033;
  wire       [31:0]   _zz_11034;
  wire       [31:0]   _zz_11035;
  wire       [31:0]   _zz_11036;
  wire       [23:0]   _zz_11037;
  wire       [31:0]   _zz_11038;
  wire       [15:0]   _zz_11039;
  wire       [15:0]   _zz_11040;
  wire       [31:0]   _zz_11041;
  wire       [31:0]   _zz_11042;
  wire       [15:0]   _zz_11043;
  wire       [31:0]   _zz_11044;
  wire       [31:0]   _zz_11045;
  wire       [31:0]   _zz_11046;
  wire       [15:0]   _zz_11047;
  wire       [31:0]   _zz_11048;
  wire       [31:0]   _zz_11049;
  wire       [31:0]   _zz_11050;
  wire       [31:0]   _zz_11051;
  wire       [31:0]   _zz_11052;
  wire       [31:0]   _zz_11053;
  wire       [23:0]   _zz_11054;
  wire       [31:0]   _zz_11055;
  wire       [15:0]   _zz_11056;
  wire       [31:0]   _zz_11057;
  wire       [31:0]   _zz_11058;
  wire       [31:0]   _zz_11059;
  wire       [31:0]   _zz_11060;
  wire       [31:0]   _zz_11061;
  wire       [23:0]   _zz_11062;
  wire       [31:0]   _zz_11063;
  wire       [15:0]   _zz_11064;
  wire       [31:0]   _zz_11065;
  wire       [31:0]   _zz_11066;
  wire       [31:0]   _zz_11067;
  wire       [31:0]   _zz_11068;
  wire       [31:0]   _zz_11069;
  wire       [23:0]   _zz_11070;
  wire       [31:0]   _zz_11071;
  wire       [15:0]   _zz_11072;
  wire       [31:0]   _zz_11073;
  wire       [31:0]   _zz_11074;
  wire       [31:0]   _zz_11075;
  wire       [31:0]   _zz_11076;
  wire       [31:0]   _zz_11077;
  wire       [23:0]   _zz_11078;
  wire       [31:0]   _zz_11079;
  wire       [15:0]   _zz_11080;
  wire       [15:0]   _zz_11081;
  wire       [31:0]   _zz_11082;
  wire       [31:0]   _zz_11083;
  wire       [15:0]   _zz_11084;
  wire       [31:0]   _zz_11085;
  wire       [31:0]   _zz_11086;
  wire       [31:0]   _zz_11087;
  wire       [15:0]   _zz_11088;
  wire       [31:0]   _zz_11089;
  wire       [31:0]   _zz_11090;
  wire       [31:0]   _zz_11091;
  wire       [31:0]   _zz_11092;
  wire       [31:0]   _zz_11093;
  wire       [31:0]   _zz_11094;
  wire       [23:0]   _zz_11095;
  wire       [31:0]   _zz_11096;
  wire       [15:0]   _zz_11097;
  wire       [31:0]   _zz_11098;
  wire       [31:0]   _zz_11099;
  wire       [31:0]   _zz_11100;
  wire       [31:0]   _zz_11101;
  wire       [31:0]   _zz_11102;
  wire       [23:0]   _zz_11103;
  wire       [31:0]   _zz_11104;
  wire       [15:0]   _zz_11105;
  wire       [31:0]   _zz_11106;
  wire       [31:0]   _zz_11107;
  wire       [31:0]   _zz_11108;
  wire       [31:0]   _zz_11109;
  wire       [31:0]   _zz_11110;
  wire       [23:0]   _zz_11111;
  wire       [31:0]   _zz_11112;
  wire       [15:0]   _zz_11113;
  wire       [31:0]   _zz_11114;
  wire       [31:0]   _zz_11115;
  wire       [31:0]   _zz_11116;
  wire       [31:0]   _zz_11117;
  wire       [31:0]   _zz_11118;
  wire       [23:0]   _zz_11119;
  wire       [31:0]   _zz_11120;
  wire       [15:0]   _zz_11121;
  wire       [15:0]   _zz_11122;
  wire       [31:0]   _zz_11123;
  wire       [31:0]   _zz_11124;
  wire       [15:0]   _zz_11125;
  wire       [31:0]   _zz_11126;
  wire       [31:0]   _zz_11127;
  wire       [31:0]   _zz_11128;
  wire       [15:0]   _zz_11129;
  wire       [31:0]   _zz_11130;
  wire       [31:0]   _zz_11131;
  wire       [31:0]   _zz_11132;
  wire       [31:0]   _zz_11133;
  wire       [31:0]   _zz_11134;
  wire       [31:0]   _zz_11135;
  wire       [23:0]   _zz_11136;
  wire       [31:0]   _zz_11137;
  wire       [15:0]   _zz_11138;
  wire       [31:0]   _zz_11139;
  wire       [31:0]   _zz_11140;
  wire       [31:0]   _zz_11141;
  wire       [31:0]   _zz_11142;
  wire       [31:0]   _zz_11143;
  wire       [23:0]   _zz_11144;
  wire       [31:0]   _zz_11145;
  wire       [15:0]   _zz_11146;
  wire       [31:0]   _zz_11147;
  wire       [31:0]   _zz_11148;
  wire       [31:0]   _zz_11149;
  wire       [31:0]   _zz_11150;
  wire       [31:0]   _zz_11151;
  wire       [23:0]   _zz_11152;
  wire       [31:0]   _zz_11153;
  wire       [15:0]   _zz_11154;
  wire       [31:0]   _zz_11155;
  wire       [31:0]   _zz_11156;
  wire       [31:0]   _zz_11157;
  wire       [31:0]   _zz_11158;
  wire       [31:0]   _zz_11159;
  wire       [23:0]   _zz_11160;
  wire       [31:0]   _zz_11161;
  wire       [15:0]   _zz_11162;
  wire       [15:0]   _zz_11163;
  wire       [31:0]   _zz_11164;
  wire       [31:0]   _zz_11165;
  wire       [15:0]   _zz_11166;
  wire       [31:0]   _zz_11167;
  wire       [31:0]   _zz_11168;
  wire       [31:0]   _zz_11169;
  wire       [15:0]   _zz_11170;
  wire       [31:0]   _zz_11171;
  wire       [31:0]   _zz_11172;
  wire       [31:0]   _zz_11173;
  wire       [31:0]   _zz_11174;
  wire       [31:0]   _zz_11175;
  wire       [31:0]   _zz_11176;
  wire       [23:0]   _zz_11177;
  wire       [31:0]   _zz_11178;
  wire       [15:0]   _zz_11179;
  wire       [31:0]   _zz_11180;
  wire       [31:0]   _zz_11181;
  wire       [31:0]   _zz_11182;
  wire       [31:0]   _zz_11183;
  wire       [31:0]   _zz_11184;
  wire       [23:0]   _zz_11185;
  wire       [31:0]   _zz_11186;
  wire       [15:0]   _zz_11187;
  wire       [31:0]   _zz_11188;
  wire       [31:0]   _zz_11189;
  wire       [31:0]   _zz_11190;
  wire       [31:0]   _zz_11191;
  wire       [31:0]   _zz_11192;
  wire       [23:0]   _zz_11193;
  wire       [31:0]   _zz_11194;
  wire       [15:0]   _zz_11195;
  wire       [31:0]   _zz_11196;
  wire       [31:0]   _zz_11197;
  wire       [31:0]   _zz_11198;
  wire       [31:0]   _zz_11199;
  wire       [31:0]   _zz_11200;
  wire       [23:0]   _zz_11201;
  wire       [31:0]   _zz_11202;
  wire       [15:0]   _zz_11203;
  wire       [15:0]   _zz_11204;
  wire       [31:0]   _zz_11205;
  wire       [31:0]   _zz_11206;
  wire       [15:0]   _zz_11207;
  wire       [31:0]   _zz_11208;
  wire       [31:0]   _zz_11209;
  wire       [31:0]   _zz_11210;
  wire       [15:0]   _zz_11211;
  wire       [31:0]   _zz_11212;
  wire       [31:0]   _zz_11213;
  wire       [31:0]   _zz_11214;
  wire       [31:0]   _zz_11215;
  wire       [31:0]   _zz_11216;
  wire       [31:0]   _zz_11217;
  wire       [23:0]   _zz_11218;
  wire       [31:0]   _zz_11219;
  wire       [15:0]   _zz_11220;
  wire       [31:0]   _zz_11221;
  wire       [31:0]   _zz_11222;
  wire       [31:0]   _zz_11223;
  wire       [31:0]   _zz_11224;
  wire       [31:0]   _zz_11225;
  wire       [23:0]   _zz_11226;
  wire       [31:0]   _zz_11227;
  wire       [15:0]   _zz_11228;
  wire       [31:0]   _zz_11229;
  wire       [31:0]   _zz_11230;
  wire       [31:0]   _zz_11231;
  wire       [31:0]   _zz_11232;
  wire       [31:0]   _zz_11233;
  wire       [23:0]   _zz_11234;
  wire       [31:0]   _zz_11235;
  wire       [15:0]   _zz_11236;
  wire       [31:0]   _zz_11237;
  wire       [31:0]   _zz_11238;
  wire       [31:0]   _zz_11239;
  wire       [31:0]   _zz_11240;
  wire       [31:0]   _zz_11241;
  wire       [23:0]   _zz_11242;
  wire       [31:0]   _zz_11243;
  wire       [15:0]   _zz_11244;
  wire       [15:0]   _zz_11245;
  wire       [31:0]   _zz_11246;
  wire       [31:0]   _zz_11247;
  wire       [15:0]   _zz_11248;
  wire       [31:0]   _zz_11249;
  wire       [31:0]   _zz_11250;
  wire       [31:0]   _zz_11251;
  wire       [15:0]   _zz_11252;
  wire       [31:0]   _zz_11253;
  wire       [31:0]   _zz_11254;
  wire       [31:0]   _zz_11255;
  wire       [31:0]   _zz_11256;
  wire       [31:0]   _zz_11257;
  wire       [31:0]   _zz_11258;
  wire       [23:0]   _zz_11259;
  wire       [31:0]   _zz_11260;
  wire       [15:0]   _zz_11261;
  wire       [31:0]   _zz_11262;
  wire       [31:0]   _zz_11263;
  wire       [31:0]   _zz_11264;
  wire       [31:0]   _zz_11265;
  wire       [31:0]   _zz_11266;
  wire       [23:0]   _zz_11267;
  wire       [31:0]   _zz_11268;
  wire       [15:0]   _zz_11269;
  wire       [31:0]   _zz_11270;
  wire       [31:0]   _zz_11271;
  wire       [31:0]   _zz_11272;
  wire       [31:0]   _zz_11273;
  wire       [31:0]   _zz_11274;
  wire       [23:0]   _zz_11275;
  wire       [31:0]   _zz_11276;
  wire       [15:0]   _zz_11277;
  wire       [31:0]   _zz_11278;
  wire       [31:0]   _zz_11279;
  wire       [31:0]   _zz_11280;
  wire       [31:0]   _zz_11281;
  wire       [31:0]   _zz_11282;
  wire       [23:0]   _zz_11283;
  wire       [31:0]   _zz_11284;
  wire       [15:0]   _zz_11285;
  wire       [15:0]   _zz_11286;
  wire       [31:0]   _zz_11287;
  wire       [31:0]   _zz_11288;
  wire       [15:0]   _zz_11289;
  wire       [31:0]   _zz_11290;
  wire       [31:0]   _zz_11291;
  wire       [31:0]   _zz_11292;
  wire       [15:0]   _zz_11293;
  wire       [31:0]   _zz_11294;
  wire       [31:0]   _zz_11295;
  wire       [31:0]   _zz_11296;
  wire       [31:0]   _zz_11297;
  wire       [31:0]   _zz_11298;
  wire       [31:0]   _zz_11299;
  wire       [23:0]   _zz_11300;
  wire       [31:0]   _zz_11301;
  wire       [15:0]   _zz_11302;
  wire       [31:0]   _zz_11303;
  wire       [31:0]   _zz_11304;
  wire       [31:0]   _zz_11305;
  wire       [31:0]   _zz_11306;
  wire       [31:0]   _zz_11307;
  wire       [23:0]   _zz_11308;
  wire       [31:0]   _zz_11309;
  wire       [15:0]   _zz_11310;
  wire       [31:0]   _zz_11311;
  wire       [31:0]   _zz_11312;
  wire       [31:0]   _zz_11313;
  wire       [31:0]   _zz_11314;
  wire       [31:0]   _zz_11315;
  wire       [23:0]   _zz_11316;
  wire       [31:0]   _zz_11317;
  wire       [15:0]   _zz_11318;
  wire       [31:0]   _zz_11319;
  wire       [31:0]   _zz_11320;
  wire       [31:0]   _zz_11321;
  wire       [31:0]   _zz_11322;
  wire       [31:0]   _zz_11323;
  wire       [23:0]   _zz_11324;
  wire       [31:0]   _zz_11325;
  wire       [15:0]   _zz_11326;
  wire       [15:0]   _zz_11327;
  wire       [31:0]   _zz_11328;
  wire       [31:0]   _zz_11329;
  wire       [15:0]   _zz_11330;
  wire       [31:0]   _zz_11331;
  wire       [31:0]   _zz_11332;
  wire       [31:0]   _zz_11333;
  wire       [15:0]   _zz_11334;
  wire       [31:0]   _zz_11335;
  wire       [31:0]   _zz_11336;
  wire       [31:0]   _zz_11337;
  wire       [31:0]   _zz_11338;
  wire       [31:0]   _zz_11339;
  wire       [31:0]   _zz_11340;
  wire       [23:0]   _zz_11341;
  wire       [31:0]   _zz_11342;
  wire       [15:0]   _zz_11343;
  wire       [31:0]   _zz_11344;
  wire       [31:0]   _zz_11345;
  wire       [31:0]   _zz_11346;
  wire       [31:0]   _zz_11347;
  wire       [31:0]   _zz_11348;
  wire       [23:0]   _zz_11349;
  wire       [31:0]   _zz_11350;
  wire       [15:0]   _zz_11351;
  wire       [31:0]   _zz_11352;
  wire       [31:0]   _zz_11353;
  wire       [31:0]   _zz_11354;
  wire       [31:0]   _zz_11355;
  wire       [31:0]   _zz_11356;
  wire       [23:0]   _zz_11357;
  wire       [31:0]   _zz_11358;
  wire       [15:0]   _zz_11359;
  wire       [31:0]   _zz_11360;
  wire       [31:0]   _zz_11361;
  wire       [31:0]   _zz_11362;
  wire       [31:0]   _zz_11363;
  wire       [31:0]   _zz_11364;
  wire       [23:0]   _zz_11365;
  wire       [31:0]   _zz_11366;
  wire       [15:0]   _zz_11367;
  wire       [15:0]   _zz_11368;
  wire       [31:0]   _zz_11369;
  wire       [31:0]   _zz_11370;
  wire       [15:0]   _zz_11371;
  wire       [31:0]   _zz_11372;
  wire       [31:0]   _zz_11373;
  wire       [31:0]   _zz_11374;
  wire       [15:0]   _zz_11375;
  wire       [31:0]   _zz_11376;
  wire       [31:0]   _zz_11377;
  wire       [31:0]   _zz_11378;
  wire       [31:0]   _zz_11379;
  wire       [31:0]   _zz_11380;
  wire       [31:0]   _zz_11381;
  wire       [23:0]   _zz_11382;
  wire       [31:0]   _zz_11383;
  wire       [15:0]   _zz_11384;
  wire       [31:0]   _zz_11385;
  wire       [31:0]   _zz_11386;
  wire       [31:0]   _zz_11387;
  wire       [31:0]   _zz_11388;
  wire       [31:0]   _zz_11389;
  wire       [23:0]   _zz_11390;
  wire       [31:0]   _zz_11391;
  wire       [15:0]   _zz_11392;
  wire       [31:0]   _zz_11393;
  wire       [31:0]   _zz_11394;
  wire       [31:0]   _zz_11395;
  wire       [31:0]   _zz_11396;
  wire       [31:0]   _zz_11397;
  wire       [23:0]   _zz_11398;
  wire       [31:0]   _zz_11399;
  wire       [15:0]   _zz_11400;
  wire       [31:0]   _zz_11401;
  wire       [31:0]   _zz_11402;
  wire       [31:0]   _zz_11403;
  wire       [31:0]   _zz_11404;
  wire       [31:0]   _zz_11405;
  wire       [23:0]   _zz_11406;
  wire       [31:0]   _zz_11407;
  wire       [15:0]   _zz_11408;
  wire       [15:0]   _zz_11409;
  wire       [31:0]   _zz_11410;
  wire       [31:0]   _zz_11411;
  wire       [15:0]   _zz_11412;
  wire       [31:0]   _zz_11413;
  wire       [31:0]   _zz_11414;
  wire       [31:0]   _zz_11415;
  wire       [15:0]   _zz_11416;
  wire       [31:0]   _zz_11417;
  wire       [31:0]   _zz_11418;
  wire       [31:0]   _zz_11419;
  wire       [31:0]   _zz_11420;
  wire       [31:0]   _zz_11421;
  wire       [31:0]   _zz_11422;
  wire       [23:0]   _zz_11423;
  wire       [31:0]   _zz_11424;
  wire       [15:0]   _zz_11425;
  wire       [31:0]   _zz_11426;
  wire       [31:0]   _zz_11427;
  wire       [31:0]   _zz_11428;
  wire       [31:0]   _zz_11429;
  wire       [31:0]   _zz_11430;
  wire       [23:0]   _zz_11431;
  wire       [31:0]   _zz_11432;
  wire       [15:0]   _zz_11433;
  wire       [31:0]   _zz_11434;
  wire       [31:0]   _zz_11435;
  wire       [31:0]   _zz_11436;
  wire       [31:0]   _zz_11437;
  wire       [31:0]   _zz_11438;
  wire       [23:0]   _zz_11439;
  wire       [31:0]   _zz_11440;
  wire       [15:0]   _zz_11441;
  wire       [31:0]   _zz_11442;
  wire       [31:0]   _zz_11443;
  wire       [31:0]   _zz_11444;
  wire       [31:0]   _zz_11445;
  wire       [31:0]   _zz_11446;
  wire       [23:0]   _zz_11447;
  wire       [31:0]   _zz_11448;
  wire       [15:0]   _zz_11449;
  wire       [15:0]   _zz_11450;
  wire       [31:0]   _zz_11451;
  wire       [31:0]   _zz_11452;
  wire       [15:0]   _zz_11453;
  wire       [31:0]   _zz_11454;
  wire       [31:0]   _zz_11455;
  wire       [31:0]   _zz_11456;
  wire       [15:0]   _zz_11457;
  wire       [31:0]   _zz_11458;
  wire       [31:0]   _zz_11459;
  wire       [31:0]   _zz_11460;
  wire       [31:0]   _zz_11461;
  wire       [31:0]   _zz_11462;
  wire       [31:0]   _zz_11463;
  wire       [23:0]   _zz_11464;
  wire       [31:0]   _zz_11465;
  wire       [15:0]   _zz_11466;
  wire       [31:0]   _zz_11467;
  wire       [31:0]   _zz_11468;
  wire       [31:0]   _zz_11469;
  wire       [31:0]   _zz_11470;
  wire       [31:0]   _zz_11471;
  wire       [23:0]   _zz_11472;
  wire       [31:0]   _zz_11473;
  wire       [15:0]   _zz_11474;
  wire       [31:0]   _zz_11475;
  wire       [31:0]   _zz_11476;
  wire       [31:0]   _zz_11477;
  wire       [31:0]   _zz_11478;
  wire       [31:0]   _zz_11479;
  wire       [23:0]   _zz_11480;
  wire       [31:0]   _zz_11481;
  wire       [15:0]   _zz_11482;
  wire       [31:0]   _zz_11483;
  wire       [31:0]   _zz_11484;
  wire       [31:0]   _zz_11485;
  wire       [31:0]   _zz_11486;
  wire       [31:0]   _zz_11487;
  wire       [23:0]   _zz_11488;
  wire       [31:0]   _zz_11489;
  wire       [15:0]   _zz_11490;
  wire       [15:0]   _zz_11491;
  wire       [31:0]   _zz_11492;
  wire       [31:0]   _zz_11493;
  wire       [15:0]   _zz_11494;
  wire       [31:0]   _zz_11495;
  wire       [31:0]   _zz_11496;
  wire       [31:0]   _zz_11497;
  wire       [15:0]   _zz_11498;
  wire       [31:0]   _zz_11499;
  wire       [31:0]   _zz_11500;
  wire       [31:0]   _zz_11501;
  wire       [31:0]   _zz_11502;
  wire       [31:0]   _zz_11503;
  wire       [31:0]   _zz_11504;
  wire       [23:0]   _zz_11505;
  wire       [31:0]   _zz_11506;
  wire       [15:0]   _zz_11507;
  wire       [31:0]   _zz_11508;
  wire       [31:0]   _zz_11509;
  wire       [31:0]   _zz_11510;
  wire       [31:0]   _zz_11511;
  wire       [31:0]   _zz_11512;
  wire       [23:0]   _zz_11513;
  wire       [31:0]   _zz_11514;
  wire       [15:0]   _zz_11515;
  wire       [31:0]   _zz_11516;
  wire       [31:0]   _zz_11517;
  wire       [31:0]   _zz_11518;
  wire       [31:0]   _zz_11519;
  wire       [31:0]   _zz_11520;
  wire       [23:0]   _zz_11521;
  wire       [31:0]   _zz_11522;
  wire       [15:0]   _zz_11523;
  wire       [31:0]   _zz_11524;
  wire       [31:0]   _zz_11525;
  wire       [31:0]   _zz_11526;
  wire       [31:0]   _zz_11527;
  wire       [31:0]   _zz_11528;
  wire       [23:0]   _zz_11529;
  wire       [31:0]   _zz_11530;
  wire       [15:0]   _zz_11531;
  wire       [15:0]   _zz_11532;
  wire       [31:0]   _zz_11533;
  wire       [31:0]   _zz_11534;
  wire       [15:0]   _zz_11535;
  wire       [31:0]   _zz_11536;
  wire       [31:0]   _zz_11537;
  wire       [31:0]   _zz_11538;
  wire       [15:0]   _zz_11539;
  wire       [31:0]   _zz_11540;
  wire       [31:0]   _zz_11541;
  wire       [31:0]   _zz_11542;
  wire       [31:0]   _zz_11543;
  wire       [31:0]   _zz_11544;
  wire       [31:0]   _zz_11545;
  wire       [23:0]   _zz_11546;
  wire       [31:0]   _zz_11547;
  wire       [15:0]   _zz_11548;
  wire       [31:0]   _zz_11549;
  wire       [31:0]   _zz_11550;
  wire       [31:0]   _zz_11551;
  wire       [31:0]   _zz_11552;
  wire       [31:0]   _zz_11553;
  wire       [23:0]   _zz_11554;
  wire       [31:0]   _zz_11555;
  wire       [15:0]   _zz_11556;
  wire       [31:0]   _zz_11557;
  wire       [31:0]   _zz_11558;
  wire       [31:0]   _zz_11559;
  wire       [31:0]   _zz_11560;
  wire       [31:0]   _zz_11561;
  wire       [23:0]   _zz_11562;
  wire       [31:0]   _zz_11563;
  wire       [15:0]   _zz_11564;
  wire       [31:0]   _zz_11565;
  wire       [31:0]   _zz_11566;
  wire       [31:0]   _zz_11567;
  wire       [31:0]   _zz_11568;
  wire       [31:0]   _zz_11569;
  wire       [23:0]   _zz_11570;
  wire       [31:0]   _zz_11571;
  wire       [15:0]   _zz_11572;
  wire       [15:0]   _zz_11573;
  wire       [31:0]   _zz_11574;
  wire       [31:0]   _zz_11575;
  wire       [15:0]   _zz_11576;
  wire       [31:0]   _zz_11577;
  wire       [31:0]   _zz_11578;
  wire       [31:0]   _zz_11579;
  wire       [15:0]   _zz_11580;
  wire       [31:0]   _zz_11581;
  wire       [31:0]   _zz_11582;
  wire       [31:0]   _zz_11583;
  wire       [31:0]   _zz_11584;
  wire       [31:0]   _zz_11585;
  wire       [31:0]   _zz_11586;
  wire       [23:0]   _zz_11587;
  wire       [31:0]   _zz_11588;
  wire       [15:0]   _zz_11589;
  wire       [31:0]   _zz_11590;
  wire       [31:0]   _zz_11591;
  wire       [31:0]   _zz_11592;
  wire       [31:0]   _zz_11593;
  wire       [31:0]   _zz_11594;
  wire       [23:0]   _zz_11595;
  wire       [31:0]   _zz_11596;
  wire       [15:0]   _zz_11597;
  wire       [31:0]   _zz_11598;
  wire       [31:0]   _zz_11599;
  wire       [31:0]   _zz_11600;
  wire       [31:0]   _zz_11601;
  wire       [31:0]   _zz_11602;
  wire       [23:0]   _zz_11603;
  wire       [31:0]   _zz_11604;
  wire       [15:0]   _zz_11605;
  wire       [31:0]   _zz_11606;
  wire       [31:0]   _zz_11607;
  wire       [31:0]   _zz_11608;
  wire       [31:0]   _zz_11609;
  wire       [31:0]   _zz_11610;
  wire       [23:0]   _zz_11611;
  wire       [31:0]   _zz_11612;
  wire       [15:0]   _zz_11613;
  wire       [15:0]   _zz_11614;
  wire       [31:0]   _zz_11615;
  wire       [31:0]   _zz_11616;
  wire       [15:0]   _zz_11617;
  wire       [31:0]   _zz_11618;
  wire       [31:0]   _zz_11619;
  wire       [31:0]   _zz_11620;
  wire       [15:0]   _zz_11621;
  wire       [31:0]   _zz_11622;
  wire       [31:0]   _zz_11623;
  wire       [31:0]   _zz_11624;
  wire       [31:0]   _zz_11625;
  wire       [31:0]   _zz_11626;
  wire       [31:0]   _zz_11627;
  wire       [23:0]   _zz_11628;
  wire       [31:0]   _zz_11629;
  wire       [15:0]   _zz_11630;
  wire       [31:0]   _zz_11631;
  wire       [31:0]   _zz_11632;
  wire       [31:0]   _zz_11633;
  wire       [31:0]   _zz_11634;
  wire       [31:0]   _zz_11635;
  wire       [23:0]   _zz_11636;
  wire       [31:0]   _zz_11637;
  wire       [15:0]   _zz_11638;
  wire       [31:0]   _zz_11639;
  wire       [31:0]   _zz_11640;
  wire       [31:0]   _zz_11641;
  wire       [31:0]   _zz_11642;
  wire       [31:0]   _zz_11643;
  wire       [23:0]   _zz_11644;
  wire       [31:0]   _zz_11645;
  wire       [15:0]   _zz_11646;
  wire       [31:0]   _zz_11647;
  wire       [31:0]   _zz_11648;
  wire       [31:0]   _zz_11649;
  wire       [31:0]   _zz_11650;
  wire       [31:0]   _zz_11651;
  wire       [23:0]   _zz_11652;
  wire       [31:0]   _zz_11653;
  wire       [15:0]   _zz_11654;
  wire       [15:0]   _zz_11655;
  wire       [31:0]   _zz_11656;
  wire       [31:0]   _zz_11657;
  wire       [15:0]   _zz_11658;
  wire       [31:0]   _zz_11659;
  wire       [31:0]   _zz_11660;
  wire       [31:0]   _zz_11661;
  wire       [15:0]   _zz_11662;
  wire       [31:0]   _zz_11663;
  wire       [31:0]   _zz_11664;
  wire       [31:0]   _zz_11665;
  wire       [31:0]   _zz_11666;
  wire       [31:0]   _zz_11667;
  wire       [31:0]   _zz_11668;
  wire       [23:0]   _zz_11669;
  wire       [31:0]   _zz_11670;
  wire       [15:0]   _zz_11671;
  wire       [31:0]   _zz_11672;
  wire       [31:0]   _zz_11673;
  wire       [31:0]   _zz_11674;
  wire       [31:0]   _zz_11675;
  wire       [31:0]   _zz_11676;
  wire       [23:0]   _zz_11677;
  wire       [31:0]   _zz_11678;
  wire       [15:0]   _zz_11679;
  wire       [31:0]   _zz_11680;
  wire       [31:0]   _zz_11681;
  wire       [31:0]   _zz_11682;
  wire       [31:0]   _zz_11683;
  wire       [31:0]   _zz_11684;
  wire       [23:0]   _zz_11685;
  wire       [31:0]   _zz_11686;
  wire       [15:0]   _zz_11687;
  wire       [31:0]   _zz_11688;
  wire       [31:0]   _zz_11689;
  wire       [31:0]   _zz_11690;
  wire       [31:0]   _zz_11691;
  wire       [31:0]   _zz_11692;
  wire       [23:0]   _zz_11693;
  wire       [31:0]   _zz_11694;
  wire       [15:0]   _zz_11695;
  wire       [15:0]   _zz_11696;
  wire       [31:0]   _zz_11697;
  wire       [31:0]   _zz_11698;
  wire       [15:0]   _zz_11699;
  wire       [31:0]   _zz_11700;
  wire       [31:0]   _zz_11701;
  wire       [31:0]   _zz_11702;
  wire       [15:0]   _zz_11703;
  wire       [31:0]   _zz_11704;
  wire       [31:0]   _zz_11705;
  wire       [31:0]   _zz_11706;
  wire       [31:0]   _zz_11707;
  wire       [31:0]   _zz_11708;
  wire       [31:0]   _zz_11709;
  wire       [23:0]   _zz_11710;
  wire       [31:0]   _zz_11711;
  wire       [15:0]   _zz_11712;
  wire       [31:0]   _zz_11713;
  wire       [31:0]   _zz_11714;
  wire       [31:0]   _zz_11715;
  wire       [31:0]   _zz_11716;
  wire       [31:0]   _zz_11717;
  wire       [23:0]   _zz_11718;
  wire       [31:0]   _zz_11719;
  wire       [15:0]   _zz_11720;
  wire       [31:0]   _zz_11721;
  wire       [31:0]   _zz_11722;
  wire       [31:0]   _zz_11723;
  wire       [31:0]   _zz_11724;
  wire       [31:0]   _zz_11725;
  wire       [23:0]   _zz_11726;
  wire       [31:0]   _zz_11727;
  wire       [15:0]   _zz_11728;
  wire       [31:0]   _zz_11729;
  wire       [31:0]   _zz_11730;
  wire       [31:0]   _zz_11731;
  wire       [31:0]   _zz_11732;
  wire       [31:0]   _zz_11733;
  wire       [23:0]   _zz_11734;
  wire       [31:0]   _zz_11735;
  wire       [15:0]   _zz_11736;
  wire       [15:0]   _zz_11737;
  wire       [31:0]   _zz_11738;
  wire       [31:0]   _zz_11739;
  wire       [15:0]   _zz_11740;
  wire       [31:0]   _zz_11741;
  wire       [31:0]   _zz_11742;
  wire       [31:0]   _zz_11743;
  wire       [15:0]   _zz_11744;
  wire       [31:0]   _zz_11745;
  wire       [31:0]   _zz_11746;
  wire       [31:0]   _zz_11747;
  wire       [31:0]   _zz_11748;
  wire       [31:0]   _zz_11749;
  wire       [31:0]   _zz_11750;
  wire       [23:0]   _zz_11751;
  wire       [31:0]   _zz_11752;
  wire       [15:0]   _zz_11753;
  wire       [31:0]   _zz_11754;
  wire       [31:0]   _zz_11755;
  wire       [31:0]   _zz_11756;
  wire       [31:0]   _zz_11757;
  wire       [31:0]   _zz_11758;
  wire       [23:0]   _zz_11759;
  wire       [31:0]   _zz_11760;
  wire       [15:0]   _zz_11761;
  wire       [31:0]   _zz_11762;
  wire       [31:0]   _zz_11763;
  wire       [31:0]   _zz_11764;
  wire       [31:0]   _zz_11765;
  wire       [31:0]   _zz_11766;
  wire       [23:0]   _zz_11767;
  wire       [31:0]   _zz_11768;
  wire       [15:0]   _zz_11769;
  wire       [31:0]   _zz_11770;
  wire       [31:0]   _zz_11771;
  wire       [31:0]   _zz_11772;
  wire       [31:0]   _zz_11773;
  wire       [31:0]   _zz_11774;
  wire       [23:0]   _zz_11775;
  wire       [31:0]   _zz_11776;
  wire       [15:0]   _zz_11777;
  wire       [15:0]   _zz_11778;
  wire       [31:0]   _zz_11779;
  wire       [31:0]   _zz_11780;
  wire       [15:0]   _zz_11781;
  wire       [31:0]   _zz_11782;
  wire       [31:0]   _zz_11783;
  wire       [31:0]   _zz_11784;
  wire       [15:0]   _zz_11785;
  wire       [31:0]   _zz_11786;
  wire       [31:0]   _zz_11787;
  wire       [31:0]   _zz_11788;
  wire       [31:0]   _zz_11789;
  wire       [31:0]   _zz_11790;
  wire       [31:0]   _zz_11791;
  wire       [23:0]   _zz_11792;
  wire       [31:0]   _zz_11793;
  wire       [15:0]   _zz_11794;
  wire       [31:0]   _zz_11795;
  wire       [31:0]   _zz_11796;
  wire       [31:0]   _zz_11797;
  wire       [31:0]   _zz_11798;
  wire       [31:0]   _zz_11799;
  wire       [23:0]   _zz_11800;
  wire       [31:0]   _zz_11801;
  wire       [15:0]   _zz_11802;
  wire       [31:0]   _zz_11803;
  wire       [31:0]   _zz_11804;
  wire       [31:0]   _zz_11805;
  wire       [31:0]   _zz_11806;
  wire       [31:0]   _zz_11807;
  wire       [23:0]   _zz_11808;
  wire       [31:0]   _zz_11809;
  wire       [15:0]   _zz_11810;
  wire       [31:0]   _zz_11811;
  wire       [31:0]   _zz_11812;
  wire       [31:0]   _zz_11813;
  wire       [31:0]   _zz_11814;
  wire       [31:0]   _zz_11815;
  wire       [23:0]   _zz_11816;
  wire       [31:0]   _zz_11817;
  wire       [15:0]   _zz_11818;
  wire       [15:0]   _zz_11819;
  wire       [31:0]   _zz_11820;
  wire       [31:0]   _zz_11821;
  wire       [15:0]   _zz_11822;
  wire       [31:0]   _zz_11823;
  wire       [31:0]   _zz_11824;
  wire       [31:0]   _zz_11825;
  wire       [15:0]   _zz_11826;
  wire       [31:0]   _zz_11827;
  wire       [31:0]   _zz_11828;
  wire       [31:0]   _zz_11829;
  wire       [31:0]   _zz_11830;
  wire       [31:0]   _zz_11831;
  wire       [31:0]   _zz_11832;
  wire       [23:0]   _zz_11833;
  wire       [31:0]   _zz_11834;
  wire       [15:0]   _zz_11835;
  wire       [31:0]   _zz_11836;
  wire       [31:0]   _zz_11837;
  wire       [31:0]   _zz_11838;
  wire       [31:0]   _zz_11839;
  wire       [31:0]   _zz_11840;
  wire       [23:0]   _zz_11841;
  wire       [31:0]   _zz_11842;
  wire       [15:0]   _zz_11843;
  wire       [31:0]   _zz_11844;
  wire       [31:0]   _zz_11845;
  wire       [31:0]   _zz_11846;
  wire       [31:0]   _zz_11847;
  wire       [31:0]   _zz_11848;
  wire       [23:0]   _zz_11849;
  wire       [31:0]   _zz_11850;
  wire       [15:0]   _zz_11851;
  wire       [31:0]   _zz_11852;
  wire       [31:0]   _zz_11853;
  wire       [31:0]   _zz_11854;
  wire       [31:0]   _zz_11855;
  wire       [31:0]   _zz_11856;
  wire       [23:0]   _zz_11857;
  wire       [31:0]   _zz_11858;
  wire       [15:0]   _zz_11859;
  wire       [15:0]   _zz_11860;
  wire       [31:0]   _zz_11861;
  wire       [31:0]   _zz_11862;
  wire       [15:0]   _zz_11863;
  wire       [31:0]   _zz_11864;
  wire       [31:0]   _zz_11865;
  wire       [31:0]   _zz_11866;
  wire       [15:0]   _zz_11867;
  wire       [31:0]   _zz_11868;
  wire       [31:0]   _zz_11869;
  wire       [31:0]   _zz_11870;
  wire       [31:0]   _zz_11871;
  wire       [31:0]   _zz_11872;
  wire       [31:0]   _zz_11873;
  wire       [23:0]   _zz_11874;
  wire       [31:0]   _zz_11875;
  wire       [15:0]   _zz_11876;
  wire       [31:0]   _zz_11877;
  wire       [31:0]   _zz_11878;
  wire       [31:0]   _zz_11879;
  wire       [31:0]   _zz_11880;
  wire       [31:0]   _zz_11881;
  wire       [23:0]   _zz_11882;
  wire       [31:0]   _zz_11883;
  wire       [15:0]   _zz_11884;
  wire       [31:0]   _zz_11885;
  wire       [31:0]   _zz_11886;
  wire       [31:0]   _zz_11887;
  wire       [31:0]   _zz_11888;
  wire       [31:0]   _zz_11889;
  wire       [23:0]   _zz_11890;
  wire       [31:0]   _zz_11891;
  wire       [15:0]   _zz_11892;
  wire       [31:0]   _zz_11893;
  wire       [31:0]   _zz_11894;
  wire       [31:0]   _zz_11895;
  wire       [31:0]   _zz_11896;
  wire       [31:0]   _zz_11897;
  wire       [23:0]   _zz_11898;
  wire       [31:0]   _zz_11899;
  wire       [15:0]   _zz_11900;
  wire       [15:0]   _zz_11901;
  wire       [31:0]   _zz_11902;
  wire       [31:0]   _zz_11903;
  wire       [15:0]   _zz_11904;
  wire       [31:0]   _zz_11905;
  wire       [31:0]   _zz_11906;
  wire       [31:0]   _zz_11907;
  wire       [15:0]   _zz_11908;
  wire       [31:0]   _zz_11909;
  wire       [31:0]   _zz_11910;
  wire       [31:0]   _zz_11911;
  wire       [31:0]   _zz_11912;
  wire       [31:0]   _zz_11913;
  wire       [31:0]   _zz_11914;
  wire       [23:0]   _zz_11915;
  wire       [31:0]   _zz_11916;
  wire       [15:0]   _zz_11917;
  wire       [31:0]   _zz_11918;
  wire       [31:0]   _zz_11919;
  wire       [31:0]   _zz_11920;
  wire       [31:0]   _zz_11921;
  wire       [31:0]   _zz_11922;
  wire       [23:0]   _zz_11923;
  wire       [31:0]   _zz_11924;
  wire       [15:0]   _zz_11925;
  wire       [31:0]   _zz_11926;
  wire       [31:0]   _zz_11927;
  wire       [31:0]   _zz_11928;
  wire       [31:0]   _zz_11929;
  wire       [31:0]   _zz_11930;
  wire       [23:0]   _zz_11931;
  wire       [31:0]   _zz_11932;
  wire       [15:0]   _zz_11933;
  wire       [31:0]   _zz_11934;
  wire       [31:0]   _zz_11935;
  wire       [31:0]   _zz_11936;
  wire       [31:0]   _zz_11937;
  wire       [31:0]   _zz_11938;
  wire       [23:0]   _zz_11939;
  wire       [31:0]   _zz_11940;
  wire       [15:0]   _zz_11941;
  wire       [15:0]   _zz_11942;
  wire       [31:0]   _zz_11943;
  wire       [31:0]   _zz_11944;
  wire       [15:0]   _zz_11945;
  wire       [31:0]   _zz_11946;
  wire       [31:0]   _zz_11947;
  wire       [31:0]   _zz_11948;
  wire       [15:0]   _zz_11949;
  wire       [31:0]   _zz_11950;
  wire       [31:0]   _zz_11951;
  wire       [31:0]   _zz_11952;
  wire       [31:0]   _zz_11953;
  wire       [31:0]   _zz_11954;
  wire       [31:0]   _zz_11955;
  wire       [23:0]   _zz_11956;
  wire       [31:0]   _zz_11957;
  wire       [15:0]   _zz_11958;
  wire       [31:0]   _zz_11959;
  wire       [31:0]   _zz_11960;
  wire       [31:0]   _zz_11961;
  wire       [31:0]   _zz_11962;
  wire       [31:0]   _zz_11963;
  wire       [23:0]   _zz_11964;
  wire       [31:0]   _zz_11965;
  wire       [15:0]   _zz_11966;
  wire       [31:0]   _zz_11967;
  wire       [31:0]   _zz_11968;
  wire       [31:0]   _zz_11969;
  wire       [31:0]   _zz_11970;
  wire       [31:0]   _zz_11971;
  wire       [23:0]   _zz_11972;
  wire       [31:0]   _zz_11973;
  wire       [15:0]   _zz_11974;
  wire       [31:0]   _zz_11975;
  wire       [31:0]   _zz_11976;
  wire       [31:0]   _zz_11977;
  wire       [31:0]   _zz_11978;
  wire       [31:0]   _zz_11979;
  wire       [23:0]   _zz_11980;
  wire       [31:0]   _zz_11981;
  wire       [15:0]   _zz_11982;
  wire       [15:0]   _zz_11983;
  wire       [31:0]   _zz_11984;
  wire       [31:0]   _zz_11985;
  wire       [15:0]   _zz_11986;
  wire       [31:0]   _zz_11987;
  wire       [31:0]   _zz_11988;
  wire       [31:0]   _zz_11989;
  wire       [15:0]   _zz_11990;
  wire       [31:0]   _zz_11991;
  wire       [31:0]   _zz_11992;
  wire       [31:0]   _zz_11993;
  wire       [31:0]   _zz_11994;
  wire       [31:0]   _zz_11995;
  wire       [31:0]   _zz_11996;
  wire       [23:0]   _zz_11997;
  wire       [31:0]   _zz_11998;
  wire       [15:0]   _zz_11999;
  wire       [31:0]   _zz_12000;
  wire       [31:0]   _zz_12001;
  wire       [31:0]   _zz_12002;
  wire       [31:0]   _zz_12003;
  wire       [31:0]   _zz_12004;
  wire       [23:0]   _zz_12005;
  wire       [31:0]   _zz_12006;
  wire       [15:0]   _zz_12007;
  wire       [31:0]   _zz_12008;
  wire       [31:0]   _zz_12009;
  wire       [31:0]   _zz_12010;
  wire       [31:0]   _zz_12011;
  wire       [31:0]   _zz_12012;
  wire       [23:0]   _zz_12013;
  wire       [31:0]   _zz_12014;
  wire       [15:0]   _zz_12015;
  wire       [31:0]   _zz_12016;
  wire       [31:0]   _zz_12017;
  wire       [31:0]   _zz_12018;
  wire       [31:0]   _zz_12019;
  wire       [31:0]   _zz_12020;
  wire       [23:0]   _zz_12021;
  wire       [31:0]   _zz_12022;
  wire       [15:0]   _zz_12023;
  wire       [15:0]   _zz_12024;
  wire       [31:0]   _zz_12025;
  wire       [31:0]   _zz_12026;
  wire       [15:0]   _zz_12027;
  wire       [31:0]   _zz_12028;
  wire       [31:0]   _zz_12029;
  wire       [31:0]   _zz_12030;
  wire       [15:0]   _zz_12031;
  wire       [31:0]   _zz_12032;
  wire       [31:0]   _zz_12033;
  wire       [31:0]   _zz_12034;
  wire       [31:0]   _zz_12035;
  wire       [31:0]   _zz_12036;
  wire       [31:0]   _zz_12037;
  wire       [23:0]   _zz_12038;
  wire       [31:0]   _zz_12039;
  wire       [15:0]   _zz_12040;
  wire       [31:0]   _zz_12041;
  wire       [31:0]   _zz_12042;
  wire       [31:0]   _zz_12043;
  wire       [31:0]   _zz_12044;
  wire       [31:0]   _zz_12045;
  wire       [23:0]   _zz_12046;
  wire       [31:0]   _zz_12047;
  wire       [15:0]   _zz_12048;
  wire       [31:0]   _zz_12049;
  wire       [31:0]   _zz_12050;
  wire       [31:0]   _zz_12051;
  wire       [31:0]   _zz_12052;
  wire       [31:0]   _zz_12053;
  wire       [23:0]   _zz_12054;
  wire       [31:0]   _zz_12055;
  wire       [15:0]   _zz_12056;
  wire       [31:0]   _zz_12057;
  wire       [31:0]   _zz_12058;
  wire       [31:0]   _zz_12059;
  wire       [31:0]   _zz_12060;
  wire       [31:0]   _zz_12061;
  wire       [23:0]   _zz_12062;
  wire       [31:0]   _zz_12063;
  wire       [15:0]   _zz_12064;
  wire       [15:0]   _zz_12065;
  wire       [31:0]   _zz_12066;
  wire       [31:0]   _zz_12067;
  wire       [15:0]   _zz_12068;
  wire       [31:0]   _zz_12069;
  wire       [31:0]   _zz_12070;
  wire       [31:0]   _zz_12071;
  wire       [15:0]   _zz_12072;
  wire       [31:0]   _zz_12073;
  wire       [31:0]   _zz_12074;
  wire       [31:0]   _zz_12075;
  wire       [31:0]   _zz_12076;
  wire       [31:0]   _zz_12077;
  wire       [31:0]   _zz_12078;
  wire       [23:0]   _zz_12079;
  wire       [31:0]   _zz_12080;
  wire       [15:0]   _zz_12081;
  wire       [31:0]   _zz_12082;
  wire       [31:0]   _zz_12083;
  wire       [31:0]   _zz_12084;
  wire       [31:0]   _zz_12085;
  wire       [31:0]   _zz_12086;
  wire       [23:0]   _zz_12087;
  wire       [31:0]   _zz_12088;
  wire       [15:0]   _zz_12089;
  wire       [31:0]   _zz_12090;
  wire       [31:0]   _zz_12091;
  wire       [31:0]   _zz_12092;
  wire       [31:0]   _zz_12093;
  wire       [31:0]   _zz_12094;
  wire       [23:0]   _zz_12095;
  wire       [31:0]   _zz_12096;
  wire       [15:0]   _zz_12097;
  wire       [31:0]   _zz_12098;
  wire       [31:0]   _zz_12099;
  wire       [31:0]   _zz_12100;
  wire       [31:0]   _zz_12101;
  wire       [31:0]   _zz_12102;
  wire       [23:0]   _zz_12103;
  wire       [31:0]   _zz_12104;
  wire       [15:0]   _zz_12105;
  wire       [15:0]   _zz_12106;
  wire       [31:0]   _zz_12107;
  wire       [31:0]   _zz_12108;
  wire       [15:0]   _zz_12109;
  wire       [31:0]   _zz_12110;
  wire       [31:0]   _zz_12111;
  wire       [31:0]   _zz_12112;
  wire       [15:0]   _zz_12113;
  wire       [31:0]   _zz_12114;
  wire       [31:0]   _zz_12115;
  wire       [31:0]   _zz_12116;
  wire       [31:0]   _zz_12117;
  wire       [31:0]   _zz_12118;
  wire       [31:0]   _zz_12119;
  wire       [23:0]   _zz_12120;
  wire       [31:0]   _zz_12121;
  wire       [15:0]   _zz_12122;
  wire       [31:0]   _zz_12123;
  wire       [31:0]   _zz_12124;
  wire       [31:0]   _zz_12125;
  wire       [31:0]   _zz_12126;
  wire       [31:0]   _zz_12127;
  wire       [23:0]   _zz_12128;
  wire       [31:0]   _zz_12129;
  wire       [15:0]   _zz_12130;
  wire       [31:0]   _zz_12131;
  wire       [31:0]   _zz_12132;
  wire       [31:0]   _zz_12133;
  wire       [31:0]   _zz_12134;
  wire       [31:0]   _zz_12135;
  wire       [23:0]   _zz_12136;
  wire       [31:0]   _zz_12137;
  wire       [15:0]   _zz_12138;
  wire       [31:0]   _zz_12139;
  wire       [31:0]   _zz_12140;
  wire       [31:0]   _zz_12141;
  wire       [31:0]   _zz_12142;
  wire       [31:0]   _zz_12143;
  wire       [23:0]   _zz_12144;
  wire       [31:0]   _zz_12145;
  wire       [15:0]   _zz_12146;
  wire       [15:0]   _zz_12147;
  wire       [31:0]   _zz_12148;
  wire       [31:0]   _zz_12149;
  wire       [15:0]   _zz_12150;
  wire       [31:0]   _zz_12151;
  wire       [31:0]   _zz_12152;
  wire       [31:0]   _zz_12153;
  wire       [15:0]   _zz_12154;
  wire       [31:0]   _zz_12155;
  wire       [31:0]   _zz_12156;
  wire       [31:0]   _zz_12157;
  wire       [31:0]   _zz_12158;
  wire       [31:0]   _zz_12159;
  wire       [31:0]   _zz_12160;
  wire       [23:0]   _zz_12161;
  wire       [31:0]   _zz_12162;
  wire       [15:0]   _zz_12163;
  wire       [31:0]   _zz_12164;
  wire       [31:0]   _zz_12165;
  wire       [31:0]   _zz_12166;
  wire       [31:0]   _zz_12167;
  wire       [31:0]   _zz_12168;
  wire       [23:0]   _zz_12169;
  wire       [31:0]   _zz_12170;
  wire       [15:0]   _zz_12171;
  wire       [31:0]   _zz_12172;
  wire       [31:0]   _zz_12173;
  wire       [31:0]   _zz_12174;
  wire       [31:0]   _zz_12175;
  wire       [31:0]   _zz_12176;
  wire       [23:0]   _zz_12177;
  wire       [31:0]   _zz_12178;
  wire       [15:0]   _zz_12179;
  wire       [31:0]   _zz_12180;
  wire       [31:0]   _zz_12181;
  wire       [31:0]   _zz_12182;
  wire       [31:0]   _zz_12183;
  wire       [31:0]   _zz_12184;
  wire       [23:0]   _zz_12185;
  wire       [31:0]   _zz_12186;
  wire       [15:0]   _zz_12187;
  wire       [15:0]   _zz_12188;
  wire       [31:0]   _zz_12189;
  wire       [31:0]   _zz_12190;
  wire       [15:0]   _zz_12191;
  wire       [31:0]   _zz_12192;
  wire       [31:0]   _zz_12193;
  wire       [31:0]   _zz_12194;
  wire       [15:0]   _zz_12195;
  wire       [31:0]   _zz_12196;
  wire       [31:0]   _zz_12197;
  wire       [31:0]   _zz_12198;
  wire       [31:0]   _zz_12199;
  wire       [31:0]   _zz_12200;
  wire       [31:0]   _zz_12201;
  wire       [23:0]   _zz_12202;
  wire       [31:0]   _zz_12203;
  wire       [15:0]   _zz_12204;
  wire       [31:0]   _zz_12205;
  wire       [31:0]   _zz_12206;
  wire       [31:0]   _zz_12207;
  wire       [31:0]   _zz_12208;
  wire       [31:0]   _zz_12209;
  wire       [23:0]   _zz_12210;
  wire       [31:0]   _zz_12211;
  wire       [15:0]   _zz_12212;
  wire       [31:0]   _zz_12213;
  wire       [31:0]   _zz_12214;
  wire       [31:0]   _zz_12215;
  wire       [31:0]   _zz_12216;
  wire       [31:0]   _zz_12217;
  wire       [23:0]   _zz_12218;
  wire       [31:0]   _zz_12219;
  wire       [15:0]   _zz_12220;
  wire       [31:0]   _zz_12221;
  wire       [31:0]   _zz_12222;
  wire       [31:0]   _zz_12223;
  wire       [31:0]   _zz_12224;
  wire       [31:0]   _zz_12225;
  wire       [23:0]   _zz_12226;
  wire       [31:0]   _zz_12227;
  wire       [15:0]   _zz_12228;
  wire       [15:0]   _zz_12229;
  wire       [31:0]   _zz_12230;
  wire       [31:0]   _zz_12231;
  wire       [15:0]   _zz_12232;
  wire       [31:0]   _zz_12233;
  wire       [31:0]   _zz_12234;
  wire       [31:0]   _zz_12235;
  wire       [15:0]   _zz_12236;
  wire       [31:0]   _zz_12237;
  wire       [31:0]   _zz_12238;
  wire       [31:0]   _zz_12239;
  wire       [31:0]   _zz_12240;
  wire       [31:0]   _zz_12241;
  wire       [31:0]   _zz_12242;
  wire       [23:0]   _zz_12243;
  wire       [31:0]   _zz_12244;
  wire       [15:0]   _zz_12245;
  wire       [31:0]   _zz_12246;
  wire       [31:0]   _zz_12247;
  wire       [31:0]   _zz_12248;
  wire       [31:0]   _zz_12249;
  wire       [31:0]   _zz_12250;
  wire       [23:0]   _zz_12251;
  wire       [31:0]   _zz_12252;
  wire       [15:0]   _zz_12253;
  wire       [31:0]   _zz_12254;
  wire       [31:0]   _zz_12255;
  wire       [31:0]   _zz_12256;
  wire       [31:0]   _zz_12257;
  wire       [31:0]   _zz_12258;
  wire       [23:0]   _zz_12259;
  wire       [31:0]   _zz_12260;
  wire       [15:0]   _zz_12261;
  wire       [31:0]   _zz_12262;
  wire       [31:0]   _zz_12263;
  wire       [31:0]   _zz_12264;
  wire       [31:0]   _zz_12265;
  wire       [31:0]   _zz_12266;
  wire       [23:0]   _zz_12267;
  wire       [31:0]   _zz_12268;
  wire       [15:0]   _zz_12269;
  wire       [15:0]   _zz_12270;
  wire       [31:0]   _zz_12271;
  wire       [31:0]   _zz_12272;
  wire       [15:0]   _zz_12273;
  wire       [31:0]   _zz_12274;
  wire       [31:0]   _zz_12275;
  wire       [31:0]   _zz_12276;
  wire       [15:0]   _zz_12277;
  wire       [31:0]   _zz_12278;
  wire       [31:0]   _zz_12279;
  wire       [31:0]   _zz_12280;
  wire       [31:0]   _zz_12281;
  wire       [31:0]   _zz_12282;
  wire       [31:0]   _zz_12283;
  wire       [23:0]   _zz_12284;
  wire       [31:0]   _zz_12285;
  wire       [15:0]   _zz_12286;
  wire       [31:0]   _zz_12287;
  wire       [31:0]   _zz_12288;
  wire       [31:0]   _zz_12289;
  wire       [31:0]   _zz_12290;
  wire       [31:0]   _zz_12291;
  wire       [23:0]   _zz_12292;
  wire       [31:0]   _zz_12293;
  wire       [15:0]   _zz_12294;
  wire       [31:0]   _zz_12295;
  wire       [31:0]   _zz_12296;
  wire       [31:0]   _zz_12297;
  wire       [31:0]   _zz_12298;
  wire       [31:0]   _zz_12299;
  wire       [23:0]   _zz_12300;
  wire       [31:0]   _zz_12301;
  wire       [15:0]   _zz_12302;
  wire       [31:0]   _zz_12303;
  wire       [31:0]   _zz_12304;
  wire       [31:0]   _zz_12305;
  wire       [31:0]   _zz_12306;
  wire       [31:0]   _zz_12307;
  wire       [23:0]   _zz_12308;
  wire       [31:0]   _zz_12309;
  wire       [15:0]   _zz_12310;
  wire       [15:0]   _zz_12311;
  wire       [31:0]   _zz_12312;
  wire       [31:0]   _zz_12313;
  wire       [15:0]   _zz_12314;
  wire       [31:0]   _zz_12315;
  wire       [31:0]   _zz_12316;
  wire       [31:0]   _zz_12317;
  wire       [15:0]   _zz_12318;
  wire       [31:0]   _zz_12319;
  wire       [31:0]   _zz_12320;
  wire       [31:0]   _zz_12321;
  wire       [31:0]   _zz_12322;
  wire       [31:0]   _zz_12323;
  wire       [31:0]   _zz_12324;
  wire       [23:0]   _zz_12325;
  wire       [31:0]   _zz_12326;
  wire       [15:0]   _zz_12327;
  wire       [31:0]   _zz_12328;
  wire       [31:0]   _zz_12329;
  wire       [31:0]   _zz_12330;
  wire       [31:0]   _zz_12331;
  wire       [31:0]   _zz_12332;
  wire       [23:0]   _zz_12333;
  wire       [31:0]   _zz_12334;
  wire       [15:0]   _zz_12335;
  wire       [31:0]   _zz_12336;
  wire       [31:0]   _zz_12337;
  wire       [31:0]   _zz_12338;
  wire       [31:0]   _zz_12339;
  wire       [31:0]   _zz_12340;
  wire       [23:0]   _zz_12341;
  wire       [31:0]   _zz_12342;
  wire       [15:0]   _zz_12343;
  wire       [31:0]   _zz_12344;
  wire       [31:0]   _zz_12345;
  wire       [31:0]   _zz_12346;
  wire       [31:0]   _zz_12347;
  wire       [31:0]   _zz_12348;
  wire       [23:0]   _zz_12349;
  wire       [31:0]   _zz_12350;
  wire       [15:0]   _zz_12351;
  wire       [15:0]   _zz_12352;
  wire       [31:0]   _zz_12353;
  wire       [31:0]   _zz_12354;
  wire       [15:0]   _zz_12355;
  wire       [31:0]   _zz_12356;
  wire       [31:0]   _zz_12357;
  wire       [31:0]   _zz_12358;
  wire       [15:0]   _zz_12359;
  wire       [31:0]   _zz_12360;
  wire       [31:0]   _zz_12361;
  wire       [31:0]   _zz_12362;
  wire       [31:0]   _zz_12363;
  wire       [31:0]   _zz_12364;
  wire       [31:0]   _zz_12365;
  wire       [23:0]   _zz_12366;
  wire       [31:0]   _zz_12367;
  wire       [15:0]   _zz_12368;
  wire       [31:0]   _zz_12369;
  wire       [31:0]   _zz_12370;
  wire       [31:0]   _zz_12371;
  wire       [31:0]   _zz_12372;
  wire       [31:0]   _zz_12373;
  wire       [23:0]   _zz_12374;
  wire       [31:0]   _zz_12375;
  wire       [15:0]   _zz_12376;
  wire       [31:0]   _zz_12377;
  wire       [31:0]   _zz_12378;
  wire       [31:0]   _zz_12379;
  wire       [31:0]   _zz_12380;
  wire       [31:0]   _zz_12381;
  wire       [23:0]   _zz_12382;
  wire       [31:0]   _zz_12383;
  wire       [15:0]   _zz_12384;
  wire       [31:0]   _zz_12385;
  wire       [31:0]   _zz_12386;
  wire       [31:0]   _zz_12387;
  wire       [31:0]   _zz_12388;
  wire       [31:0]   _zz_12389;
  wire       [23:0]   _zz_12390;
  wire       [31:0]   _zz_12391;
  wire       [15:0]   _zz_12392;
  wire       [15:0]   _zz_12393;
  wire       [31:0]   _zz_12394;
  wire       [31:0]   _zz_12395;
  wire       [15:0]   _zz_12396;
  wire       [31:0]   _zz_12397;
  wire       [31:0]   _zz_12398;
  wire       [31:0]   _zz_12399;
  wire       [15:0]   _zz_12400;
  wire       [31:0]   _zz_12401;
  wire       [31:0]   _zz_12402;
  wire       [31:0]   _zz_12403;
  wire       [31:0]   _zz_12404;
  wire       [31:0]   _zz_12405;
  wire       [31:0]   _zz_12406;
  wire       [23:0]   _zz_12407;
  wire       [31:0]   _zz_12408;
  wire       [15:0]   _zz_12409;
  wire       [31:0]   _zz_12410;
  wire       [31:0]   _zz_12411;
  wire       [31:0]   _zz_12412;
  wire       [31:0]   _zz_12413;
  wire       [31:0]   _zz_12414;
  wire       [23:0]   _zz_12415;
  wire       [31:0]   _zz_12416;
  wire       [15:0]   _zz_12417;
  wire       [31:0]   _zz_12418;
  wire       [31:0]   _zz_12419;
  wire       [31:0]   _zz_12420;
  wire       [31:0]   _zz_12421;
  wire       [31:0]   _zz_12422;
  wire       [23:0]   _zz_12423;
  wire       [31:0]   _zz_12424;
  wire       [15:0]   _zz_12425;
  wire       [31:0]   _zz_12426;
  wire       [31:0]   _zz_12427;
  wire       [31:0]   _zz_12428;
  wire       [31:0]   _zz_12429;
  wire       [31:0]   _zz_12430;
  wire       [23:0]   _zz_12431;
  wire       [31:0]   _zz_12432;
  wire       [15:0]   _zz_12433;
  wire       [15:0]   _zz_12434;
  wire       [31:0]   _zz_12435;
  wire       [31:0]   _zz_12436;
  wire       [15:0]   _zz_12437;
  wire       [31:0]   _zz_12438;
  wire       [31:0]   _zz_12439;
  wire       [31:0]   _zz_12440;
  wire       [15:0]   _zz_12441;
  wire       [31:0]   _zz_12442;
  wire       [31:0]   _zz_12443;
  wire       [31:0]   _zz_12444;
  wire       [31:0]   _zz_12445;
  wire       [31:0]   _zz_12446;
  wire       [31:0]   _zz_12447;
  wire       [23:0]   _zz_12448;
  wire       [31:0]   _zz_12449;
  wire       [15:0]   _zz_12450;
  wire       [31:0]   _zz_12451;
  wire       [31:0]   _zz_12452;
  wire       [31:0]   _zz_12453;
  wire       [31:0]   _zz_12454;
  wire       [31:0]   _zz_12455;
  wire       [23:0]   _zz_12456;
  wire       [31:0]   _zz_12457;
  wire       [15:0]   _zz_12458;
  wire       [31:0]   _zz_12459;
  wire       [31:0]   _zz_12460;
  wire       [31:0]   _zz_12461;
  wire       [31:0]   _zz_12462;
  wire       [31:0]   _zz_12463;
  wire       [23:0]   _zz_12464;
  wire       [31:0]   _zz_12465;
  wire       [15:0]   _zz_12466;
  wire       [31:0]   _zz_12467;
  wire       [31:0]   _zz_12468;
  wire       [31:0]   _zz_12469;
  wire       [31:0]   _zz_12470;
  wire       [31:0]   _zz_12471;
  wire       [23:0]   _zz_12472;
  wire       [31:0]   _zz_12473;
  wire       [15:0]   _zz_12474;
  wire       [15:0]   _zz_12475;
  wire       [31:0]   _zz_12476;
  wire       [31:0]   _zz_12477;
  wire       [15:0]   _zz_12478;
  wire       [31:0]   _zz_12479;
  wire       [31:0]   _zz_12480;
  wire       [31:0]   _zz_12481;
  wire       [15:0]   _zz_12482;
  wire       [31:0]   _zz_12483;
  wire       [31:0]   _zz_12484;
  wire       [31:0]   _zz_12485;
  wire       [31:0]   _zz_12486;
  wire       [31:0]   _zz_12487;
  wire       [31:0]   _zz_12488;
  wire       [23:0]   _zz_12489;
  wire       [31:0]   _zz_12490;
  wire       [15:0]   _zz_12491;
  wire       [31:0]   _zz_12492;
  wire       [31:0]   _zz_12493;
  wire       [31:0]   _zz_12494;
  wire       [31:0]   _zz_12495;
  wire       [31:0]   _zz_12496;
  wire       [23:0]   _zz_12497;
  wire       [31:0]   _zz_12498;
  wire       [15:0]   _zz_12499;
  wire       [31:0]   _zz_12500;
  wire       [31:0]   _zz_12501;
  wire       [31:0]   _zz_12502;
  wire       [31:0]   _zz_12503;
  wire       [31:0]   _zz_12504;
  wire       [23:0]   _zz_12505;
  wire       [31:0]   _zz_12506;
  wire       [15:0]   _zz_12507;
  wire       [31:0]   _zz_12508;
  wire       [31:0]   _zz_12509;
  wire       [31:0]   _zz_12510;
  wire       [31:0]   _zz_12511;
  wire       [31:0]   _zz_12512;
  wire       [23:0]   _zz_12513;
  wire       [31:0]   _zz_12514;
  wire       [15:0]   _zz_12515;
  wire       [15:0]   _zz_12516;
  wire       [31:0]   _zz_12517;
  wire       [31:0]   _zz_12518;
  wire       [15:0]   _zz_12519;
  wire       [31:0]   _zz_12520;
  wire       [31:0]   _zz_12521;
  wire       [31:0]   _zz_12522;
  wire       [15:0]   _zz_12523;
  wire       [31:0]   _zz_12524;
  wire       [31:0]   _zz_12525;
  wire       [31:0]   _zz_12526;
  wire       [31:0]   _zz_12527;
  wire       [31:0]   _zz_12528;
  wire       [31:0]   _zz_12529;
  wire       [23:0]   _zz_12530;
  wire       [31:0]   _zz_12531;
  wire       [15:0]   _zz_12532;
  wire       [31:0]   _zz_12533;
  wire       [31:0]   _zz_12534;
  wire       [31:0]   _zz_12535;
  wire       [31:0]   _zz_12536;
  wire       [31:0]   _zz_12537;
  wire       [23:0]   _zz_12538;
  wire       [31:0]   _zz_12539;
  wire       [15:0]   _zz_12540;
  wire       [31:0]   _zz_12541;
  wire       [31:0]   _zz_12542;
  wire       [31:0]   _zz_12543;
  wire       [31:0]   _zz_12544;
  wire       [31:0]   _zz_12545;
  wire       [23:0]   _zz_12546;
  wire       [31:0]   _zz_12547;
  wire       [15:0]   _zz_12548;
  wire       [31:0]   _zz_12549;
  wire       [31:0]   _zz_12550;
  wire       [31:0]   _zz_12551;
  wire       [31:0]   _zz_12552;
  wire       [31:0]   _zz_12553;
  wire       [23:0]   _zz_12554;
  wire       [31:0]   _zz_12555;
  wire       [15:0]   _zz_12556;
  wire       [15:0]   _zz_12557;
  wire       [31:0]   _zz_12558;
  wire       [31:0]   _zz_12559;
  wire       [15:0]   _zz_12560;
  wire       [31:0]   _zz_12561;
  wire       [31:0]   _zz_12562;
  wire       [31:0]   _zz_12563;
  wire       [15:0]   _zz_12564;
  wire       [31:0]   _zz_12565;
  wire       [31:0]   _zz_12566;
  wire       [31:0]   _zz_12567;
  wire       [31:0]   _zz_12568;
  wire       [31:0]   _zz_12569;
  wire       [31:0]   _zz_12570;
  wire       [23:0]   _zz_12571;
  wire       [31:0]   _zz_12572;
  wire       [15:0]   _zz_12573;
  wire       [31:0]   _zz_12574;
  wire       [31:0]   _zz_12575;
  wire       [31:0]   _zz_12576;
  wire       [31:0]   _zz_12577;
  wire       [31:0]   _zz_12578;
  wire       [23:0]   _zz_12579;
  wire       [31:0]   _zz_12580;
  wire       [15:0]   _zz_12581;
  wire       [31:0]   _zz_12582;
  wire       [31:0]   _zz_12583;
  wire       [31:0]   _zz_12584;
  wire       [31:0]   _zz_12585;
  wire       [31:0]   _zz_12586;
  wire       [23:0]   _zz_12587;
  wire       [31:0]   _zz_12588;
  wire       [15:0]   _zz_12589;
  wire       [31:0]   _zz_12590;
  wire       [31:0]   _zz_12591;
  wire       [31:0]   _zz_12592;
  wire       [31:0]   _zz_12593;
  wire       [31:0]   _zz_12594;
  wire       [23:0]   _zz_12595;
  wire       [31:0]   _zz_12596;
  wire       [15:0]   _zz_12597;
  wire       [15:0]   _zz_12598;
  wire       [31:0]   _zz_12599;
  wire       [31:0]   _zz_12600;
  wire       [15:0]   _zz_12601;
  wire       [31:0]   _zz_12602;
  wire       [31:0]   _zz_12603;
  wire       [31:0]   _zz_12604;
  wire       [15:0]   _zz_12605;
  wire       [31:0]   _zz_12606;
  wire       [31:0]   _zz_12607;
  wire       [31:0]   _zz_12608;
  wire       [31:0]   _zz_12609;
  wire       [31:0]   _zz_12610;
  wire       [31:0]   _zz_12611;
  wire       [23:0]   _zz_12612;
  wire       [31:0]   _zz_12613;
  wire       [15:0]   _zz_12614;
  wire       [31:0]   _zz_12615;
  wire       [31:0]   _zz_12616;
  wire       [31:0]   _zz_12617;
  wire       [31:0]   _zz_12618;
  wire       [31:0]   _zz_12619;
  wire       [23:0]   _zz_12620;
  wire       [31:0]   _zz_12621;
  wire       [15:0]   _zz_12622;
  wire       [31:0]   _zz_12623;
  wire       [31:0]   _zz_12624;
  wire       [31:0]   _zz_12625;
  wire       [31:0]   _zz_12626;
  wire       [31:0]   _zz_12627;
  wire       [23:0]   _zz_12628;
  wire       [31:0]   _zz_12629;
  wire       [15:0]   _zz_12630;
  wire       [31:0]   _zz_12631;
  wire       [31:0]   _zz_12632;
  wire       [31:0]   _zz_12633;
  wire       [31:0]   _zz_12634;
  wire       [31:0]   _zz_12635;
  wire       [23:0]   _zz_12636;
  wire       [31:0]   _zz_12637;
  wire       [15:0]   _zz_12638;
  wire       [15:0]   _zz_12639;
  wire       [31:0]   _zz_12640;
  wire       [31:0]   _zz_12641;
  wire       [15:0]   _zz_12642;
  wire       [31:0]   _zz_12643;
  wire       [31:0]   _zz_12644;
  wire       [31:0]   _zz_12645;
  wire       [15:0]   _zz_12646;
  wire       [31:0]   _zz_12647;
  wire       [31:0]   _zz_12648;
  wire       [31:0]   _zz_12649;
  wire       [31:0]   _zz_12650;
  wire       [31:0]   _zz_12651;
  wire       [31:0]   _zz_12652;
  wire       [23:0]   _zz_12653;
  wire       [31:0]   _zz_12654;
  wire       [15:0]   _zz_12655;
  wire       [31:0]   _zz_12656;
  wire       [31:0]   _zz_12657;
  wire       [31:0]   _zz_12658;
  wire       [31:0]   _zz_12659;
  wire       [31:0]   _zz_12660;
  wire       [23:0]   _zz_12661;
  wire       [31:0]   _zz_12662;
  wire       [15:0]   _zz_12663;
  wire       [31:0]   _zz_12664;
  wire       [31:0]   _zz_12665;
  wire       [31:0]   _zz_12666;
  wire       [31:0]   _zz_12667;
  wire       [31:0]   _zz_12668;
  wire       [23:0]   _zz_12669;
  wire       [31:0]   _zz_12670;
  wire       [15:0]   _zz_12671;
  wire       [31:0]   _zz_12672;
  wire       [31:0]   _zz_12673;
  wire       [31:0]   _zz_12674;
  wire       [31:0]   _zz_12675;
  wire       [31:0]   _zz_12676;
  wire       [23:0]   _zz_12677;
  wire       [31:0]   _zz_12678;
  wire       [15:0]   _zz_12679;
  wire       [15:0]   _zz_12680;
  wire       [31:0]   _zz_12681;
  wire       [31:0]   _zz_12682;
  wire       [15:0]   _zz_12683;
  wire       [31:0]   _zz_12684;
  wire       [31:0]   _zz_12685;
  wire       [31:0]   _zz_12686;
  wire       [15:0]   _zz_12687;
  wire       [31:0]   _zz_12688;
  wire       [31:0]   _zz_12689;
  wire       [31:0]   _zz_12690;
  wire       [31:0]   _zz_12691;
  wire       [31:0]   _zz_12692;
  wire       [31:0]   _zz_12693;
  wire       [23:0]   _zz_12694;
  wire       [31:0]   _zz_12695;
  wire       [15:0]   _zz_12696;
  wire       [31:0]   _zz_12697;
  wire       [31:0]   _zz_12698;
  wire       [31:0]   _zz_12699;
  wire       [31:0]   _zz_12700;
  wire       [31:0]   _zz_12701;
  wire       [23:0]   _zz_12702;
  wire       [31:0]   _zz_12703;
  wire       [15:0]   _zz_12704;
  wire       [31:0]   _zz_12705;
  wire       [31:0]   _zz_12706;
  wire       [31:0]   _zz_12707;
  wire       [31:0]   _zz_12708;
  wire       [31:0]   _zz_12709;
  wire       [23:0]   _zz_12710;
  wire       [31:0]   _zz_12711;
  wire       [15:0]   _zz_12712;
  wire       [31:0]   _zz_12713;
  wire       [31:0]   _zz_12714;
  wire       [31:0]   _zz_12715;
  wire       [31:0]   _zz_12716;
  wire       [31:0]   _zz_12717;
  wire       [23:0]   _zz_12718;
  wire       [31:0]   _zz_12719;
  wire       [15:0]   _zz_12720;
  wire       [15:0]   _zz_12721;
  wire       [31:0]   _zz_12722;
  wire       [31:0]   _zz_12723;
  wire       [15:0]   _zz_12724;
  wire       [31:0]   _zz_12725;
  wire       [31:0]   _zz_12726;
  wire       [31:0]   _zz_12727;
  wire       [15:0]   _zz_12728;
  wire       [31:0]   _zz_12729;
  wire       [31:0]   _zz_12730;
  wire       [31:0]   _zz_12731;
  wire       [31:0]   _zz_12732;
  wire       [31:0]   _zz_12733;
  wire       [31:0]   _zz_12734;
  wire       [23:0]   _zz_12735;
  wire       [31:0]   _zz_12736;
  wire       [15:0]   _zz_12737;
  wire       [31:0]   _zz_12738;
  wire       [31:0]   _zz_12739;
  wire       [31:0]   _zz_12740;
  wire       [31:0]   _zz_12741;
  wire       [31:0]   _zz_12742;
  wire       [23:0]   _zz_12743;
  wire       [31:0]   _zz_12744;
  wire       [15:0]   _zz_12745;
  wire       [31:0]   _zz_12746;
  wire       [31:0]   _zz_12747;
  wire       [31:0]   _zz_12748;
  wire       [31:0]   _zz_12749;
  wire       [31:0]   _zz_12750;
  wire       [23:0]   _zz_12751;
  wire       [31:0]   _zz_12752;
  wire       [15:0]   _zz_12753;
  wire       [31:0]   _zz_12754;
  wire       [31:0]   _zz_12755;
  wire       [31:0]   _zz_12756;
  wire       [31:0]   _zz_12757;
  wire       [31:0]   _zz_12758;
  wire       [23:0]   _zz_12759;
  wire       [31:0]   _zz_12760;
  wire       [15:0]   _zz_12761;
  wire       [15:0]   _zz_12762;
  wire       [31:0]   _zz_12763;
  wire       [31:0]   _zz_12764;
  wire       [15:0]   _zz_12765;
  wire       [31:0]   _zz_12766;
  wire       [31:0]   _zz_12767;
  wire       [31:0]   _zz_12768;
  wire       [15:0]   _zz_12769;
  wire       [31:0]   _zz_12770;
  wire       [31:0]   _zz_12771;
  wire       [31:0]   _zz_12772;
  wire       [31:0]   _zz_12773;
  wire       [31:0]   _zz_12774;
  wire       [31:0]   _zz_12775;
  wire       [23:0]   _zz_12776;
  wire       [31:0]   _zz_12777;
  wire       [15:0]   _zz_12778;
  wire       [31:0]   _zz_12779;
  wire       [31:0]   _zz_12780;
  wire       [31:0]   _zz_12781;
  wire       [31:0]   _zz_12782;
  wire       [31:0]   _zz_12783;
  wire       [23:0]   _zz_12784;
  wire       [31:0]   _zz_12785;
  wire       [15:0]   _zz_12786;
  wire       [31:0]   _zz_12787;
  wire       [31:0]   _zz_12788;
  wire       [31:0]   _zz_12789;
  wire       [31:0]   _zz_12790;
  wire       [31:0]   _zz_12791;
  wire       [23:0]   _zz_12792;
  wire       [31:0]   _zz_12793;
  wire       [15:0]   _zz_12794;
  wire       [31:0]   _zz_12795;
  wire       [31:0]   _zz_12796;
  wire       [31:0]   _zz_12797;
  wire       [31:0]   _zz_12798;
  wire       [31:0]   _zz_12799;
  wire       [23:0]   _zz_12800;
  wire       [31:0]   _zz_12801;
  wire       [15:0]   _zz_12802;
  wire       [15:0]   _zz_12803;
  wire       [31:0]   _zz_12804;
  wire       [31:0]   _zz_12805;
  wire       [15:0]   _zz_12806;
  wire       [31:0]   _zz_12807;
  wire       [31:0]   _zz_12808;
  wire       [31:0]   _zz_12809;
  wire       [15:0]   _zz_12810;
  wire       [31:0]   _zz_12811;
  wire       [31:0]   _zz_12812;
  wire       [31:0]   _zz_12813;
  wire       [31:0]   _zz_12814;
  wire       [31:0]   _zz_12815;
  wire       [31:0]   _zz_12816;
  wire       [23:0]   _zz_12817;
  wire       [31:0]   _zz_12818;
  wire       [15:0]   _zz_12819;
  wire       [31:0]   _zz_12820;
  wire       [31:0]   _zz_12821;
  wire       [31:0]   _zz_12822;
  wire       [31:0]   _zz_12823;
  wire       [31:0]   _zz_12824;
  wire       [23:0]   _zz_12825;
  wire       [31:0]   _zz_12826;
  wire       [15:0]   _zz_12827;
  wire       [31:0]   _zz_12828;
  wire       [31:0]   _zz_12829;
  wire       [31:0]   _zz_12830;
  wire       [31:0]   _zz_12831;
  wire       [31:0]   _zz_12832;
  wire       [23:0]   _zz_12833;
  wire       [31:0]   _zz_12834;
  wire       [15:0]   _zz_12835;
  wire       [31:0]   _zz_12836;
  wire       [31:0]   _zz_12837;
  wire       [31:0]   _zz_12838;
  wire       [31:0]   _zz_12839;
  wire       [31:0]   _zz_12840;
  wire       [23:0]   _zz_12841;
  wire       [31:0]   _zz_12842;
  wire       [15:0]   _zz_12843;
  wire       [15:0]   _zz_12844;
  wire       [31:0]   _zz_12845;
  wire       [31:0]   _zz_12846;
  wire       [15:0]   _zz_12847;
  wire       [31:0]   _zz_12848;
  wire       [31:0]   _zz_12849;
  wire       [31:0]   _zz_12850;
  wire       [15:0]   _zz_12851;
  wire       [31:0]   _zz_12852;
  wire       [31:0]   _zz_12853;
  wire       [31:0]   _zz_12854;
  wire       [31:0]   _zz_12855;
  wire       [31:0]   _zz_12856;
  wire       [31:0]   _zz_12857;
  wire       [23:0]   _zz_12858;
  wire       [31:0]   _zz_12859;
  wire       [15:0]   _zz_12860;
  wire       [31:0]   _zz_12861;
  wire       [31:0]   _zz_12862;
  wire       [31:0]   _zz_12863;
  wire       [31:0]   _zz_12864;
  wire       [31:0]   _zz_12865;
  wire       [23:0]   _zz_12866;
  wire       [31:0]   _zz_12867;
  wire       [15:0]   _zz_12868;
  wire       [31:0]   _zz_12869;
  wire       [31:0]   _zz_12870;
  wire       [31:0]   _zz_12871;
  wire       [31:0]   _zz_12872;
  wire       [31:0]   _zz_12873;
  wire       [23:0]   _zz_12874;
  wire       [31:0]   _zz_12875;
  wire       [15:0]   _zz_12876;
  wire       [31:0]   _zz_12877;
  wire       [31:0]   _zz_12878;
  wire       [31:0]   _zz_12879;
  wire       [31:0]   _zz_12880;
  wire       [31:0]   _zz_12881;
  wire       [23:0]   _zz_12882;
  wire       [31:0]   _zz_12883;
  wire       [15:0]   _zz_12884;
  wire       [15:0]   _zz_12885;
  wire       [31:0]   _zz_12886;
  wire       [31:0]   _zz_12887;
  wire       [15:0]   _zz_12888;
  wire       [31:0]   _zz_12889;
  wire       [31:0]   _zz_12890;
  wire       [31:0]   _zz_12891;
  wire       [15:0]   _zz_12892;
  wire       [31:0]   _zz_12893;
  wire       [31:0]   _zz_12894;
  wire       [31:0]   _zz_12895;
  wire       [31:0]   _zz_12896;
  wire       [31:0]   _zz_12897;
  wire       [31:0]   _zz_12898;
  wire       [23:0]   _zz_12899;
  wire       [31:0]   _zz_12900;
  wire       [15:0]   _zz_12901;
  wire       [31:0]   _zz_12902;
  wire       [31:0]   _zz_12903;
  wire       [31:0]   _zz_12904;
  wire       [31:0]   _zz_12905;
  wire       [31:0]   _zz_12906;
  wire       [23:0]   _zz_12907;
  wire       [31:0]   _zz_12908;
  wire       [15:0]   _zz_12909;
  wire       [31:0]   _zz_12910;
  wire       [31:0]   _zz_12911;
  wire       [31:0]   _zz_12912;
  wire       [31:0]   _zz_12913;
  wire       [31:0]   _zz_12914;
  wire       [23:0]   _zz_12915;
  wire       [31:0]   _zz_12916;
  wire       [15:0]   _zz_12917;
  wire       [31:0]   _zz_12918;
  wire       [31:0]   _zz_12919;
  wire       [31:0]   _zz_12920;
  wire       [31:0]   _zz_12921;
  wire       [31:0]   _zz_12922;
  wire       [23:0]   _zz_12923;
  wire       [31:0]   _zz_12924;
  wire       [15:0]   _zz_12925;
  wire       [15:0]   _zz_12926;
  wire       [31:0]   _zz_12927;
  wire       [31:0]   _zz_12928;
  wire       [15:0]   _zz_12929;
  wire       [31:0]   _zz_12930;
  wire       [31:0]   _zz_12931;
  wire       [31:0]   _zz_12932;
  wire       [15:0]   _zz_12933;
  wire       [31:0]   _zz_12934;
  wire       [31:0]   _zz_12935;
  wire       [31:0]   _zz_12936;
  wire       [31:0]   _zz_12937;
  wire       [31:0]   _zz_12938;
  wire       [31:0]   _zz_12939;
  wire       [23:0]   _zz_12940;
  wire       [31:0]   _zz_12941;
  wire       [15:0]   _zz_12942;
  wire       [31:0]   _zz_12943;
  wire       [31:0]   _zz_12944;
  wire       [31:0]   _zz_12945;
  wire       [31:0]   _zz_12946;
  wire       [31:0]   _zz_12947;
  wire       [23:0]   _zz_12948;
  wire       [31:0]   _zz_12949;
  wire       [15:0]   _zz_12950;
  wire       [31:0]   _zz_12951;
  wire       [31:0]   _zz_12952;
  wire       [31:0]   _zz_12953;
  wire       [31:0]   _zz_12954;
  wire       [31:0]   _zz_12955;
  wire       [23:0]   _zz_12956;
  wire       [31:0]   _zz_12957;
  wire       [15:0]   _zz_12958;
  wire       [31:0]   _zz_12959;
  wire       [31:0]   _zz_12960;
  wire       [31:0]   _zz_12961;
  wire       [31:0]   _zz_12962;
  wire       [31:0]   _zz_12963;
  wire       [23:0]   _zz_12964;
  wire       [31:0]   _zz_12965;
  wire       [15:0]   _zz_12966;
  wire       [15:0]   _zz_12967;
  wire       [31:0]   _zz_12968;
  wire       [31:0]   _zz_12969;
  wire       [15:0]   _zz_12970;
  wire       [31:0]   _zz_12971;
  wire       [31:0]   _zz_12972;
  wire       [31:0]   _zz_12973;
  wire       [15:0]   _zz_12974;
  wire       [31:0]   _zz_12975;
  wire       [31:0]   _zz_12976;
  wire       [31:0]   _zz_12977;
  wire       [31:0]   _zz_12978;
  wire       [31:0]   _zz_12979;
  wire       [31:0]   _zz_12980;
  wire       [23:0]   _zz_12981;
  wire       [31:0]   _zz_12982;
  wire       [15:0]   _zz_12983;
  wire       [31:0]   _zz_12984;
  wire       [31:0]   _zz_12985;
  wire       [31:0]   _zz_12986;
  wire       [31:0]   _zz_12987;
  wire       [31:0]   _zz_12988;
  wire       [23:0]   _zz_12989;
  wire       [31:0]   _zz_12990;
  wire       [15:0]   _zz_12991;
  wire       [31:0]   _zz_12992;
  wire       [31:0]   _zz_12993;
  wire       [31:0]   _zz_12994;
  wire       [31:0]   _zz_12995;
  wire       [31:0]   _zz_12996;
  wire       [23:0]   _zz_12997;
  wire       [31:0]   _zz_12998;
  wire       [15:0]   _zz_12999;
  wire       [31:0]   _zz_13000;
  wire       [31:0]   _zz_13001;
  wire       [31:0]   _zz_13002;
  wire       [31:0]   _zz_13003;
  wire       [31:0]   _zz_13004;
  wire       [23:0]   _zz_13005;
  wire       [31:0]   _zz_13006;
  wire       [15:0]   _zz_13007;
  wire       [15:0]   _zz_13008;
  wire       [31:0]   _zz_13009;
  wire       [31:0]   _zz_13010;
  wire       [15:0]   _zz_13011;
  wire       [31:0]   _zz_13012;
  wire       [31:0]   _zz_13013;
  wire       [31:0]   _zz_13014;
  wire       [15:0]   _zz_13015;
  wire       [31:0]   _zz_13016;
  wire       [31:0]   _zz_13017;
  wire       [31:0]   _zz_13018;
  wire       [31:0]   _zz_13019;
  wire       [31:0]   _zz_13020;
  wire       [31:0]   _zz_13021;
  wire       [23:0]   _zz_13022;
  wire       [31:0]   _zz_13023;
  wire       [15:0]   _zz_13024;
  wire       [31:0]   _zz_13025;
  wire       [31:0]   _zz_13026;
  wire       [31:0]   _zz_13027;
  wire       [31:0]   _zz_13028;
  wire       [31:0]   _zz_13029;
  wire       [23:0]   _zz_13030;
  wire       [31:0]   _zz_13031;
  wire       [15:0]   _zz_13032;
  wire       [31:0]   _zz_13033;
  wire       [31:0]   _zz_13034;
  wire       [31:0]   _zz_13035;
  wire       [31:0]   _zz_13036;
  wire       [31:0]   _zz_13037;
  wire       [23:0]   _zz_13038;
  wire       [31:0]   _zz_13039;
  wire       [15:0]   _zz_13040;
  wire       [31:0]   _zz_13041;
  wire       [31:0]   _zz_13042;
  wire       [31:0]   _zz_13043;
  wire       [31:0]   _zz_13044;
  wire       [31:0]   _zz_13045;
  wire       [23:0]   _zz_13046;
  wire       [31:0]   _zz_13047;
  wire       [15:0]   _zz_13048;
  wire       [15:0]   _zz_13049;
  wire       [31:0]   _zz_13050;
  wire       [31:0]   _zz_13051;
  wire       [15:0]   _zz_13052;
  wire       [31:0]   _zz_13053;
  wire       [31:0]   _zz_13054;
  wire       [31:0]   _zz_13055;
  wire       [15:0]   _zz_13056;
  wire       [31:0]   _zz_13057;
  wire       [31:0]   _zz_13058;
  wire       [31:0]   _zz_13059;
  wire       [31:0]   _zz_13060;
  wire       [31:0]   _zz_13061;
  wire       [31:0]   _zz_13062;
  wire       [23:0]   _zz_13063;
  wire       [31:0]   _zz_13064;
  wire       [15:0]   _zz_13065;
  wire       [31:0]   _zz_13066;
  wire       [31:0]   _zz_13067;
  wire       [31:0]   _zz_13068;
  wire       [31:0]   _zz_13069;
  wire       [31:0]   _zz_13070;
  wire       [23:0]   _zz_13071;
  wire       [31:0]   _zz_13072;
  wire       [15:0]   _zz_13073;
  wire       [31:0]   _zz_13074;
  wire       [31:0]   _zz_13075;
  wire       [31:0]   _zz_13076;
  wire       [31:0]   _zz_13077;
  wire       [31:0]   _zz_13078;
  wire       [23:0]   _zz_13079;
  wire       [31:0]   _zz_13080;
  wire       [15:0]   _zz_13081;
  wire       [31:0]   _zz_13082;
  wire       [31:0]   _zz_13083;
  wire       [31:0]   _zz_13084;
  wire       [31:0]   _zz_13085;
  wire       [31:0]   _zz_13086;
  wire       [23:0]   _zz_13087;
  wire       [31:0]   _zz_13088;
  wire       [15:0]   _zz_13089;
  wire       [15:0]   _zz_13090;
  wire       [31:0]   _zz_13091;
  wire       [31:0]   _zz_13092;
  wire       [15:0]   _zz_13093;
  wire       [31:0]   _zz_13094;
  wire       [31:0]   _zz_13095;
  wire       [31:0]   _zz_13096;
  wire       [15:0]   _zz_13097;
  wire       [31:0]   _zz_13098;
  wire       [31:0]   _zz_13099;
  wire       [31:0]   _zz_13100;
  wire       [31:0]   _zz_13101;
  wire       [31:0]   _zz_13102;
  wire       [31:0]   _zz_13103;
  wire       [23:0]   _zz_13104;
  wire       [31:0]   _zz_13105;
  wire       [15:0]   _zz_13106;
  wire       [31:0]   _zz_13107;
  wire       [31:0]   _zz_13108;
  wire       [31:0]   _zz_13109;
  wire       [31:0]   _zz_13110;
  wire       [31:0]   _zz_13111;
  wire       [23:0]   _zz_13112;
  wire       [31:0]   _zz_13113;
  wire       [15:0]   _zz_13114;
  wire       [31:0]   _zz_13115;
  wire       [31:0]   _zz_13116;
  wire       [31:0]   _zz_13117;
  wire       [31:0]   _zz_13118;
  wire       [31:0]   _zz_13119;
  wire       [23:0]   _zz_13120;
  wire       [31:0]   _zz_13121;
  wire       [15:0]   _zz_13122;
  wire       [31:0]   _zz_13123;
  wire       [31:0]   _zz_13124;
  wire       [31:0]   _zz_13125;
  wire       [31:0]   _zz_13126;
  wire       [31:0]   _zz_13127;
  wire       [23:0]   _zz_13128;
  wire       [31:0]   _zz_13129;
  wire       [15:0]   _zz_13130;
  wire       [15:0]   _zz_13131;
  wire       [31:0]   _zz_13132;
  wire       [31:0]   _zz_13133;
  wire       [15:0]   _zz_13134;
  wire       [31:0]   _zz_13135;
  wire       [31:0]   _zz_13136;
  wire       [31:0]   _zz_13137;
  wire       [15:0]   _zz_13138;
  wire       [31:0]   _zz_13139;
  wire       [31:0]   _zz_13140;
  wire       [31:0]   _zz_13141;
  wire       [31:0]   _zz_13142;
  wire       [31:0]   _zz_13143;
  wire       [31:0]   _zz_13144;
  wire       [23:0]   _zz_13145;
  wire       [31:0]   _zz_13146;
  wire       [15:0]   _zz_13147;
  wire       [31:0]   _zz_13148;
  wire       [31:0]   _zz_13149;
  wire       [31:0]   _zz_13150;
  wire       [31:0]   _zz_13151;
  wire       [31:0]   _zz_13152;
  wire       [23:0]   _zz_13153;
  wire       [31:0]   _zz_13154;
  wire       [15:0]   _zz_13155;
  wire       [31:0]   _zz_13156;
  wire       [31:0]   _zz_13157;
  wire       [31:0]   _zz_13158;
  wire       [31:0]   _zz_13159;
  wire       [31:0]   _zz_13160;
  wire       [23:0]   _zz_13161;
  wire       [31:0]   _zz_13162;
  wire       [15:0]   _zz_13163;
  wire       [31:0]   _zz_13164;
  wire       [31:0]   _zz_13165;
  wire       [31:0]   _zz_13166;
  wire       [31:0]   _zz_13167;
  wire       [31:0]   _zz_13168;
  wire       [23:0]   _zz_13169;
  wire       [31:0]   _zz_13170;
  wire       [15:0]   _zz_13171;
  wire       [15:0]   _zz_13172;
  wire       [31:0]   _zz_13173;
  wire       [31:0]   _zz_13174;
  wire       [15:0]   _zz_13175;
  wire       [31:0]   _zz_13176;
  wire       [31:0]   _zz_13177;
  wire       [31:0]   _zz_13178;
  wire       [15:0]   _zz_13179;
  wire       [31:0]   _zz_13180;
  wire       [31:0]   _zz_13181;
  wire       [31:0]   _zz_13182;
  wire       [31:0]   _zz_13183;
  wire       [31:0]   _zz_13184;
  wire       [31:0]   _zz_13185;
  wire       [23:0]   _zz_13186;
  wire       [31:0]   _zz_13187;
  wire       [15:0]   _zz_13188;
  wire       [31:0]   _zz_13189;
  wire       [31:0]   _zz_13190;
  wire       [31:0]   _zz_13191;
  wire       [31:0]   _zz_13192;
  wire       [31:0]   _zz_13193;
  wire       [23:0]   _zz_13194;
  wire       [31:0]   _zz_13195;
  wire       [15:0]   _zz_13196;
  wire       [31:0]   _zz_13197;
  wire       [31:0]   _zz_13198;
  wire       [31:0]   _zz_13199;
  wire       [31:0]   _zz_13200;
  wire       [31:0]   _zz_13201;
  wire       [23:0]   _zz_13202;
  wire       [31:0]   _zz_13203;
  wire       [15:0]   _zz_13204;
  wire       [31:0]   _zz_13205;
  wire       [31:0]   _zz_13206;
  wire       [31:0]   _zz_13207;
  wire       [31:0]   _zz_13208;
  wire       [31:0]   _zz_13209;
  wire       [23:0]   _zz_13210;
  wire       [31:0]   _zz_13211;
  wire       [15:0]   _zz_13212;
  wire       [15:0]   _zz_13213;
  wire       [31:0]   _zz_13214;
  wire       [31:0]   _zz_13215;
  wire       [15:0]   _zz_13216;
  wire       [31:0]   _zz_13217;
  wire       [31:0]   _zz_13218;
  wire       [31:0]   _zz_13219;
  wire       [15:0]   _zz_13220;
  wire       [31:0]   _zz_13221;
  wire       [31:0]   _zz_13222;
  wire       [31:0]   _zz_13223;
  wire       [31:0]   _zz_13224;
  wire       [31:0]   _zz_13225;
  wire       [31:0]   _zz_13226;
  wire       [23:0]   _zz_13227;
  wire       [31:0]   _zz_13228;
  wire       [15:0]   _zz_13229;
  wire       [31:0]   _zz_13230;
  wire       [31:0]   _zz_13231;
  wire       [31:0]   _zz_13232;
  wire       [31:0]   _zz_13233;
  wire       [31:0]   _zz_13234;
  wire       [23:0]   _zz_13235;
  wire       [31:0]   _zz_13236;
  wire       [15:0]   _zz_13237;
  wire       [31:0]   _zz_13238;
  wire       [31:0]   _zz_13239;
  wire       [31:0]   _zz_13240;
  wire       [31:0]   _zz_13241;
  wire       [31:0]   _zz_13242;
  wire       [23:0]   _zz_13243;
  wire       [31:0]   _zz_13244;
  wire       [15:0]   _zz_13245;
  wire       [31:0]   _zz_13246;
  wire       [31:0]   _zz_13247;
  wire       [31:0]   _zz_13248;
  wire       [31:0]   _zz_13249;
  wire       [31:0]   _zz_13250;
  wire       [23:0]   _zz_13251;
  wire       [31:0]   _zz_13252;
  wire       [15:0]   _zz_13253;
  wire       [15:0]   _zz_13254;
  wire       [31:0]   _zz_13255;
  wire       [31:0]   _zz_13256;
  wire       [15:0]   _zz_13257;
  wire       [31:0]   _zz_13258;
  wire       [31:0]   _zz_13259;
  wire       [31:0]   _zz_13260;
  wire       [15:0]   _zz_13261;
  wire       [31:0]   _zz_13262;
  wire       [31:0]   _zz_13263;
  wire       [31:0]   _zz_13264;
  wire       [31:0]   _zz_13265;
  wire       [31:0]   _zz_13266;
  wire       [31:0]   _zz_13267;
  wire       [23:0]   _zz_13268;
  wire       [31:0]   _zz_13269;
  wire       [15:0]   _zz_13270;
  wire       [31:0]   _zz_13271;
  wire       [31:0]   _zz_13272;
  wire       [31:0]   _zz_13273;
  wire       [31:0]   _zz_13274;
  wire       [31:0]   _zz_13275;
  wire       [23:0]   _zz_13276;
  wire       [31:0]   _zz_13277;
  wire       [15:0]   _zz_13278;
  wire       [31:0]   _zz_13279;
  wire       [31:0]   _zz_13280;
  wire       [31:0]   _zz_13281;
  wire       [31:0]   _zz_13282;
  wire       [31:0]   _zz_13283;
  wire       [23:0]   _zz_13284;
  wire       [31:0]   _zz_13285;
  wire       [15:0]   _zz_13286;
  wire       [31:0]   _zz_13287;
  wire       [31:0]   _zz_13288;
  wire       [31:0]   _zz_13289;
  wire       [31:0]   _zz_13290;
  wire       [31:0]   _zz_13291;
  wire       [23:0]   _zz_13292;
  wire       [31:0]   _zz_13293;
  wire       [15:0]   _zz_13294;
  wire       [15:0]   _zz_13295;
  wire       [31:0]   _zz_13296;
  wire       [31:0]   _zz_13297;
  wire       [15:0]   _zz_13298;
  wire       [31:0]   _zz_13299;
  wire       [31:0]   _zz_13300;
  wire       [31:0]   _zz_13301;
  wire       [15:0]   _zz_13302;
  wire       [31:0]   _zz_13303;
  wire       [31:0]   _zz_13304;
  wire       [31:0]   _zz_13305;
  wire       [31:0]   _zz_13306;
  wire       [31:0]   _zz_13307;
  wire       [31:0]   _zz_13308;
  wire       [23:0]   _zz_13309;
  wire       [31:0]   _zz_13310;
  wire       [15:0]   _zz_13311;
  wire       [31:0]   _zz_13312;
  wire       [31:0]   _zz_13313;
  wire       [31:0]   _zz_13314;
  wire       [31:0]   _zz_13315;
  wire       [31:0]   _zz_13316;
  wire       [23:0]   _zz_13317;
  wire       [31:0]   _zz_13318;
  wire       [15:0]   _zz_13319;
  wire       [31:0]   _zz_13320;
  wire       [31:0]   _zz_13321;
  wire       [31:0]   _zz_13322;
  wire       [31:0]   _zz_13323;
  wire       [31:0]   _zz_13324;
  wire       [23:0]   _zz_13325;
  wire       [31:0]   _zz_13326;
  wire       [15:0]   _zz_13327;
  wire       [31:0]   _zz_13328;
  wire       [31:0]   _zz_13329;
  wire       [31:0]   _zz_13330;
  wire       [31:0]   _zz_13331;
  wire       [31:0]   _zz_13332;
  wire       [23:0]   _zz_13333;
  wire       [31:0]   _zz_13334;
  wire       [15:0]   _zz_13335;
  wire       [15:0]   _zz_13336;
  wire       [31:0]   _zz_13337;
  wire       [31:0]   _zz_13338;
  wire       [15:0]   _zz_13339;
  wire       [31:0]   _zz_13340;
  wire       [31:0]   _zz_13341;
  wire       [31:0]   _zz_13342;
  wire       [15:0]   _zz_13343;
  wire       [31:0]   _zz_13344;
  wire       [31:0]   _zz_13345;
  wire       [31:0]   _zz_13346;
  wire       [31:0]   _zz_13347;
  wire       [31:0]   _zz_13348;
  wire       [31:0]   _zz_13349;
  wire       [23:0]   _zz_13350;
  wire       [31:0]   _zz_13351;
  wire       [15:0]   _zz_13352;
  wire       [31:0]   _zz_13353;
  wire       [31:0]   _zz_13354;
  wire       [31:0]   _zz_13355;
  wire       [31:0]   _zz_13356;
  wire       [31:0]   _zz_13357;
  wire       [23:0]   _zz_13358;
  wire       [31:0]   _zz_13359;
  wire       [15:0]   _zz_13360;
  wire       [31:0]   _zz_13361;
  wire       [31:0]   _zz_13362;
  wire       [31:0]   _zz_13363;
  wire       [31:0]   _zz_13364;
  wire       [31:0]   _zz_13365;
  wire       [23:0]   _zz_13366;
  wire       [31:0]   _zz_13367;
  wire       [15:0]   _zz_13368;
  wire       [31:0]   _zz_13369;
  wire       [31:0]   _zz_13370;
  wire       [31:0]   _zz_13371;
  wire       [31:0]   _zz_13372;
  wire       [31:0]   _zz_13373;
  wire       [23:0]   _zz_13374;
  wire       [31:0]   _zz_13375;
  wire       [15:0]   _zz_13376;
  wire       [15:0]   _zz_13377;
  wire       [31:0]   _zz_13378;
  wire       [31:0]   _zz_13379;
  wire       [15:0]   _zz_13380;
  wire       [31:0]   _zz_13381;
  wire       [31:0]   _zz_13382;
  wire       [31:0]   _zz_13383;
  wire       [15:0]   _zz_13384;
  wire       [31:0]   _zz_13385;
  wire       [31:0]   _zz_13386;
  wire       [31:0]   _zz_13387;
  wire       [31:0]   _zz_13388;
  wire       [31:0]   _zz_13389;
  wire       [31:0]   _zz_13390;
  wire       [23:0]   _zz_13391;
  wire       [31:0]   _zz_13392;
  wire       [15:0]   _zz_13393;
  wire       [31:0]   _zz_13394;
  wire       [31:0]   _zz_13395;
  wire       [31:0]   _zz_13396;
  wire       [31:0]   _zz_13397;
  wire       [31:0]   _zz_13398;
  wire       [23:0]   _zz_13399;
  wire       [31:0]   _zz_13400;
  wire       [15:0]   _zz_13401;
  wire       [31:0]   _zz_13402;
  wire       [31:0]   _zz_13403;
  wire       [31:0]   _zz_13404;
  wire       [31:0]   _zz_13405;
  wire       [31:0]   _zz_13406;
  wire       [23:0]   _zz_13407;
  wire       [31:0]   _zz_13408;
  wire       [15:0]   _zz_13409;
  wire       [31:0]   _zz_13410;
  wire       [31:0]   _zz_13411;
  wire       [31:0]   _zz_13412;
  wire       [31:0]   _zz_13413;
  wire       [31:0]   _zz_13414;
  wire       [23:0]   _zz_13415;
  wire       [31:0]   _zz_13416;
  wire       [15:0]   _zz_13417;
  wire       [15:0]   _zz_13418;
  wire       [31:0]   _zz_13419;
  wire       [31:0]   _zz_13420;
  wire       [15:0]   _zz_13421;
  wire       [31:0]   _zz_13422;
  wire       [31:0]   _zz_13423;
  wire       [31:0]   _zz_13424;
  wire       [15:0]   _zz_13425;
  wire       [31:0]   _zz_13426;
  wire       [31:0]   _zz_13427;
  wire       [31:0]   _zz_13428;
  wire       [31:0]   _zz_13429;
  wire       [31:0]   _zz_13430;
  wire       [31:0]   _zz_13431;
  wire       [23:0]   _zz_13432;
  wire       [31:0]   _zz_13433;
  wire       [15:0]   _zz_13434;
  wire       [31:0]   _zz_13435;
  wire       [31:0]   _zz_13436;
  wire       [31:0]   _zz_13437;
  wire       [31:0]   _zz_13438;
  wire       [31:0]   _zz_13439;
  wire       [23:0]   _zz_13440;
  wire       [31:0]   _zz_13441;
  wire       [15:0]   _zz_13442;
  wire       [31:0]   _zz_13443;
  wire       [31:0]   _zz_13444;
  wire       [31:0]   _zz_13445;
  wire       [31:0]   _zz_13446;
  wire       [31:0]   _zz_13447;
  wire       [23:0]   _zz_13448;
  wire       [31:0]   _zz_13449;
  wire       [15:0]   _zz_13450;
  wire       [31:0]   _zz_13451;
  wire       [31:0]   _zz_13452;
  wire       [31:0]   _zz_13453;
  wire       [31:0]   _zz_13454;
  wire       [31:0]   _zz_13455;
  wire       [23:0]   _zz_13456;
  wire       [31:0]   _zz_13457;
  wire       [15:0]   _zz_13458;
  wire       [15:0]   _zz_13459;
  wire       [31:0]   _zz_13460;
  wire       [31:0]   _zz_13461;
  wire       [15:0]   _zz_13462;
  wire       [31:0]   _zz_13463;
  wire       [31:0]   _zz_13464;
  wire       [31:0]   _zz_13465;
  wire       [15:0]   _zz_13466;
  wire       [31:0]   _zz_13467;
  wire       [31:0]   _zz_13468;
  wire       [31:0]   _zz_13469;
  wire       [31:0]   _zz_13470;
  wire       [31:0]   _zz_13471;
  wire       [31:0]   _zz_13472;
  wire       [23:0]   _zz_13473;
  wire       [31:0]   _zz_13474;
  wire       [15:0]   _zz_13475;
  wire       [31:0]   _zz_13476;
  wire       [31:0]   _zz_13477;
  wire       [31:0]   _zz_13478;
  wire       [31:0]   _zz_13479;
  wire       [31:0]   _zz_13480;
  wire       [23:0]   _zz_13481;
  wire       [31:0]   _zz_13482;
  wire       [15:0]   _zz_13483;
  wire       [31:0]   _zz_13484;
  wire       [31:0]   _zz_13485;
  wire       [31:0]   _zz_13486;
  wire       [31:0]   _zz_13487;
  wire       [31:0]   _zz_13488;
  wire       [23:0]   _zz_13489;
  wire       [31:0]   _zz_13490;
  wire       [15:0]   _zz_13491;
  wire       [31:0]   _zz_13492;
  wire       [31:0]   _zz_13493;
  wire       [31:0]   _zz_13494;
  wire       [31:0]   _zz_13495;
  wire       [31:0]   _zz_13496;
  wire       [23:0]   _zz_13497;
  wire       [31:0]   _zz_13498;
  wire       [15:0]   _zz_13499;
  wire       [15:0]   _zz_13500;
  wire       [31:0]   _zz_13501;
  wire       [31:0]   _zz_13502;
  wire       [15:0]   _zz_13503;
  wire       [31:0]   _zz_13504;
  wire       [31:0]   _zz_13505;
  wire       [31:0]   _zz_13506;
  wire       [15:0]   _zz_13507;
  wire       [31:0]   _zz_13508;
  wire       [31:0]   _zz_13509;
  wire       [31:0]   _zz_13510;
  wire       [31:0]   _zz_13511;
  wire       [31:0]   _zz_13512;
  wire       [31:0]   _zz_13513;
  wire       [23:0]   _zz_13514;
  wire       [31:0]   _zz_13515;
  wire       [15:0]   _zz_13516;
  wire       [31:0]   _zz_13517;
  wire       [31:0]   _zz_13518;
  wire       [31:0]   _zz_13519;
  wire       [31:0]   _zz_13520;
  wire       [31:0]   _zz_13521;
  wire       [23:0]   _zz_13522;
  wire       [31:0]   _zz_13523;
  wire       [15:0]   _zz_13524;
  wire       [31:0]   _zz_13525;
  wire       [31:0]   _zz_13526;
  wire       [31:0]   _zz_13527;
  wire       [31:0]   _zz_13528;
  wire       [31:0]   _zz_13529;
  wire       [23:0]   _zz_13530;
  wire       [31:0]   _zz_13531;
  wire       [15:0]   _zz_13532;
  wire       [31:0]   _zz_13533;
  wire       [31:0]   _zz_13534;
  wire       [31:0]   _zz_13535;
  wire       [31:0]   _zz_13536;
  wire       [31:0]   _zz_13537;
  wire       [23:0]   _zz_13538;
  wire       [31:0]   _zz_13539;
  wire       [15:0]   _zz_13540;
  wire       [15:0]   _zz_13541;
  wire       [31:0]   _zz_13542;
  wire       [31:0]   _zz_13543;
  wire       [15:0]   _zz_13544;
  wire       [31:0]   _zz_13545;
  wire       [31:0]   _zz_13546;
  wire       [31:0]   _zz_13547;
  wire       [15:0]   _zz_13548;
  wire       [31:0]   _zz_13549;
  wire       [31:0]   _zz_13550;
  wire       [31:0]   _zz_13551;
  wire       [31:0]   _zz_13552;
  wire       [31:0]   _zz_13553;
  wire       [31:0]   _zz_13554;
  wire       [23:0]   _zz_13555;
  wire       [31:0]   _zz_13556;
  wire       [15:0]   _zz_13557;
  wire       [31:0]   _zz_13558;
  wire       [31:0]   _zz_13559;
  wire       [31:0]   _zz_13560;
  wire       [31:0]   _zz_13561;
  wire       [31:0]   _zz_13562;
  wire       [23:0]   _zz_13563;
  wire       [31:0]   _zz_13564;
  wire       [15:0]   _zz_13565;
  wire       [31:0]   _zz_13566;
  wire       [31:0]   _zz_13567;
  wire       [31:0]   _zz_13568;
  wire       [31:0]   _zz_13569;
  wire       [31:0]   _zz_13570;
  wire       [23:0]   _zz_13571;
  wire       [31:0]   _zz_13572;
  wire       [15:0]   _zz_13573;
  wire       [31:0]   _zz_13574;
  wire       [31:0]   _zz_13575;
  wire       [31:0]   _zz_13576;
  wire       [31:0]   _zz_13577;
  wire       [31:0]   _zz_13578;
  wire       [23:0]   _zz_13579;
  wire       [31:0]   _zz_13580;
  wire       [15:0]   _zz_13581;
  wire       [15:0]   _zz_13582;
  wire       [31:0]   _zz_13583;
  wire       [31:0]   _zz_13584;
  wire       [15:0]   _zz_13585;
  wire       [31:0]   _zz_13586;
  wire       [31:0]   _zz_13587;
  wire       [31:0]   _zz_13588;
  wire       [15:0]   _zz_13589;
  wire       [31:0]   _zz_13590;
  wire       [31:0]   _zz_13591;
  wire       [31:0]   _zz_13592;
  wire       [31:0]   _zz_13593;
  wire       [31:0]   _zz_13594;
  wire       [31:0]   _zz_13595;
  wire       [23:0]   _zz_13596;
  wire       [31:0]   _zz_13597;
  wire       [15:0]   _zz_13598;
  wire       [31:0]   _zz_13599;
  wire       [31:0]   _zz_13600;
  wire       [31:0]   _zz_13601;
  wire       [31:0]   _zz_13602;
  wire       [31:0]   _zz_13603;
  wire       [23:0]   _zz_13604;
  wire       [31:0]   _zz_13605;
  wire       [15:0]   _zz_13606;
  wire       [31:0]   _zz_13607;
  wire       [31:0]   _zz_13608;
  wire       [31:0]   _zz_13609;
  wire       [31:0]   _zz_13610;
  wire       [31:0]   _zz_13611;
  wire       [23:0]   _zz_13612;
  wire       [31:0]   _zz_13613;
  wire       [15:0]   _zz_13614;
  wire       [31:0]   _zz_13615;
  wire       [31:0]   _zz_13616;
  wire       [31:0]   _zz_13617;
  wire       [31:0]   _zz_13618;
  wire       [31:0]   _zz_13619;
  wire       [23:0]   _zz_13620;
  wire       [31:0]   _zz_13621;
  wire       [15:0]   _zz_13622;
  wire       [15:0]   _zz_13623;
  wire       [31:0]   _zz_13624;
  wire       [31:0]   _zz_13625;
  wire       [15:0]   _zz_13626;
  wire       [31:0]   _zz_13627;
  wire       [31:0]   _zz_13628;
  wire       [31:0]   _zz_13629;
  wire       [15:0]   _zz_13630;
  wire       [31:0]   _zz_13631;
  wire       [31:0]   _zz_13632;
  wire       [31:0]   _zz_13633;
  wire       [31:0]   _zz_13634;
  wire       [31:0]   _zz_13635;
  wire       [31:0]   _zz_13636;
  wire       [23:0]   _zz_13637;
  wire       [31:0]   _zz_13638;
  wire       [15:0]   _zz_13639;
  wire       [31:0]   _zz_13640;
  wire       [31:0]   _zz_13641;
  wire       [31:0]   _zz_13642;
  wire       [31:0]   _zz_13643;
  wire       [31:0]   _zz_13644;
  wire       [23:0]   _zz_13645;
  wire       [31:0]   _zz_13646;
  wire       [15:0]   _zz_13647;
  wire       [31:0]   _zz_13648;
  wire       [31:0]   _zz_13649;
  wire       [31:0]   _zz_13650;
  wire       [31:0]   _zz_13651;
  wire       [31:0]   _zz_13652;
  wire       [23:0]   _zz_13653;
  wire       [31:0]   _zz_13654;
  wire       [15:0]   _zz_13655;
  wire       [31:0]   _zz_13656;
  wire       [31:0]   _zz_13657;
  wire       [31:0]   _zz_13658;
  wire       [31:0]   _zz_13659;
  wire       [31:0]   _zz_13660;
  wire       [23:0]   _zz_13661;
  wire       [31:0]   _zz_13662;
  wire       [15:0]   _zz_13663;
  wire       [15:0]   _zz_13664;
  wire       [31:0]   _zz_13665;
  wire       [31:0]   _zz_13666;
  wire       [15:0]   _zz_13667;
  wire       [31:0]   _zz_13668;
  wire       [31:0]   _zz_13669;
  wire       [31:0]   _zz_13670;
  wire       [15:0]   _zz_13671;
  wire       [31:0]   _zz_13672;
  wire       [31:0]   _zz_13673;
  wire       [31:0]   _zz_13674;
  wire       [31:0]   _zz_13675;
  wire       [31:0]   _zz_13676;
  wire       [31:0]   _zz_13677;
  wire       [23:0]   _zz_13678;
  wire       [31:0]   _zz_13679;
  wire       [15:0]   _zz_13680;
  wire       [31:0]   _zz_13681;
  wire       [31:0]   _zz_13682;
  wire       [31:0]   _zz_13683;
  wire       [31:0]   _zz_13684;
  wire       [31:0]   _zz_13685;
  wire       [23:0]   _zz_13686;
  wire       [31:0]   _zz_13687;
  wire       [15:0]   _zz_13688;
  wire       [31:0]   _zz_13689;
  wire       [31:0]   _zz_13690;
  wire       [31:0]   _zz_13691;
  wire       [31:0]   _zz_13692;
  wire       [31:0]   _zz_13693;
  wire       [23:0]   _zz_13694;
  wire       [31:0]   _zz_13695;
  wire       [15:0]   _zz_13696;
  wire       [31:0]   _zz_13697;
  wire       [31:0]   _zz_13698;
  wire       [31:0]   _zz_13699;
  wire       [31:0]   _zz_13700;
  wire       [31:0]   _zz_13701;
  wire       [23:0]   _zz_13702;
  wire       [31:0]   _zz_13703;
  wire       [15:0]   _zz_13704;
  wire       [15:0]   _zz_13705;
  wire       [31:0]   _zz_13706;
  wire       [31:0]   _zz_13707;
  wire       [15:0]   _zz_13708;
  wire       [31:0]   _zz_13709;
  wire       [31:0]   _zz_13710;
  wire       [31:0]   _zz_13711;
  wire       [15:0]   _zz_13712;
  wire       [31:0]   _zz_13713;
  wire       [31:0]   _zz_13714;
  wire       [31:0]   _zz_13715;
  wire       [31:0]   _zz_13716;
  wire       [31:0]   _zz_13717;
  wire       [31:0]   _zz_13718;
  wire       [23:0]   _zz_13719;
  wire       [31:0]   _zz_13720;
  wire       [15:0]   _zz_13721;
  wire       [31:0]   _zz_13722;
  wire       [31:0]   _zz_13723;
  wire       [31:0]   _zz_13724;
  wire       [31:0]   _zz_13725;
  wire       [31:0]   _zz_13726;
  wire       [23:0]   _zz_13727;
  wire       [31:0]   _zz_13728;
  wire       [15:0]   _zz_13729;
  wire       [31:0]   _zz_13730;
  wire       [31:0]   _zz_13731;
  wire       [31:0]   _zz_13732;
  wire       [31:0]   _zz_13733;
  wire       [31:0]   _zz_13734;
  wire       [23:0]   _zz_13735;
  wire       [31:0]   _zz_13736;
  wire       [15:0]   _zz_13737;
  wire       [31:0]   _zz_13738;
  wire       [31:0]   _zz_13739;
  wire       [31:0]   _zz_13740;
  wire       [31:0]   _zz_13741;
  wire       [31:0]   _zz_13742;
  wire       [23:0]   _zz_13743;
  wire       [31:0]   _zz_13744;
  wire       [15:0]   _zz_13745;
  wire       [15:0]   _zz_13746;
  wire       [31:0]   _zz_13747;
  wire       [31:0]   _zz_13748;
  wire       [15:0]   _zz_13749;
  wire       [31:0]   _zz_13750;
  wire       [31:0]   _zz_13751;
  wire       [31:0]   _zz_13752;
  wire       [15:0]   _zz_13753;
  wire       [31:0]   _zz_13754;
  wire       [31:0]   _zz_13755;
  wire       [31:0]   _zz_13756;
  wire       [31:0]   _zz_13757;
  wire       [31:0]   _zz_13758;
  wire       [31:0]   _zz_13759;
  wire       [23:0]   _zz_13760;
  wire       [31:0]   _zz_13761;
  wire       [15:0]   _zz_13762;
  wire       [31:0]   _zz_13763;
  wire       [31:0]   _zz_13764;
  wire       [31:0]   _zz_13765;
  wire       [31:0]   _zz_13766;
  wire       [31:0]   _zz_13767;
  wire       [23:0]   _zz_13768;
  wire       [31:0]   _zz_13769;
  wire       [15:0]   _zz_13770;
  wire       [31:0]   _zz_13771;
  wire       [31:0]   _zz_13772;
  wire       [31:0]   _zz_13773;
  wire       [31:0]   _zz_13774;
  wire       [31:0]   _zz_13775;
  wire       [23:0]   _zz_13776;
  wire       [31:0]   _zz_13777;
  wire       [15:0]   _zz_13778;
  wire       [31:0]   _zz_13779;
  wire       [31:0]   _zz_13780;
  wire       [31:0]   _zz_13781;
  wire       [31:0]   _zz_13782;
  wire       [31:0]   _zz_13783;
  wire       [23:0]   _zz_13784;
  wire       [31:0]   _zz_13785;
  wire       [15:0]   _zz_13786;
  wire       [15:0]   _zz_13787;
  wire       [31:0]   _zz_13788;
  wire       [31:0]   _zz_13789;
  wire       [15:0]   _zz_13790;
  wire       [31:0]   _zz_13791;
  wire       [31:0]   _zz_13792;
  wire       [31:0]   _zz_13793;
  wire       [15:0]   _zz_13794;
  wire       [31:0]   _zz_13795;
  wire       [31:0]   _zz_13796;
  wire       [31:0]   _zz_13797;
  wire       [31:0]   _zz_13798;
  wire       [31:0]   _zz_13799;
  wire       [31:0]   _zz_13800;
  wire       [23:0]   _zz_13801;
  wire       [31:0]   _zz_13802;
  wire       [15:0]   _zz_13803;
  wire       [31:0]   _zz_13804;
  wire       [31:0]   _zz_13805;
  wire       [31:0]   _zz_13806;
  wire       [31:0]   _zz_13807;
  wire       [31:0]   _zz_13808;
  wire       [23:0]   _zz_13809;
  wire       [31:0]   _zz_13810;
  wire       [15:0]   _zz_13811;
  wire       [31:0]   _zz_13812;
  wire       [31:0]   _zz_13813;
  wire       [31:0]   _zz_13814;
  wire       [31:0]   _zz_13815;
  wire       [31:0]   _zz_13816;
  wire       [23:0]   _zz_13817;
  wire       [31:0]   _zz_13818;
  wire       [15:0]   _zz_13819;
  wire       [31:0]   _zz_13820;
  wire       [31:0]   _zz_13821;
  wire       [31:0]   _zz_13822;
  wire       [31:0]   _zz_13823;
  wire       [31:0]   _zz_13824;
  wire       [23:0]   _zz_13825;
  wire       [31:0]   _zz_13826;
  wire       [15:0]   _zz_13827;
  wire       [15:0]   _zz_13828;
  wire       [31:0]   _zz_13829;
  wire       [31:0]   _zz_13830;
  wire       [15:0]   _zz_13831;
  wire       [31:0]   _zz_13832;
  wire       [31:0]   _zz_13833;
  wire       [31:0]   _zz_13834;
  wire       [15:0]   _zz_13835;
  wire       [31:0]   _zz_13836;
  wire       [31:0]   _zz_13837;
  wire       [31:0]   _zz_13838;
  wire       [31:0]   _zz_13839;
  wire       [31:0]   _zz_13840;
  wire       [31:0]   _zz_13841;
  wire       [23:0]   _zz_13842;
  wire       [31:0]   _zz_13843;
  wire       [15:0]   _zz_13844;
  wire       [31:0]   _zz_13845;
  wire       [31:0]   _zz_13846;
  wire       [31:0]   _zz_13847;
  wire       [31:0]   _zz_13848;
  wire       [31:0]   _zz_13849;
  wire       [23:0]   _zz_13850;
  wire       [31:0]   _zz_13851;
  wire       [15:0]   _zz_13852;
  wire       [31:0]   _zz_13853;
  wire       [31:0]   _zz_13854;
  wire       [31:0]   _zz_13855;
  wire       [31:0]   _zz_13856;
  wire       [31:0]   _zz_13857;
  wire       [23:0]   _zz_13858;
  wire       [31:0]   _zz_13859;
  wire       [15:0]   _zz_13860;
  wire       [31:0]   _zz_13861;
  wire       [31:0]   _zz_13862;
  wire       [31:0]   _zz_13863;
  wire       [31:0]   _zz_13864;
  wire       [31:0]   _zz_13865;
  wire       [23:0]   _zz_13866;
  wire       [31:0]   _zz_13867;
  wire       [15:0]   _zz_13868;
  wire       [15:0]   _zz_13869;
  wire       [31:0]   _zz_13870;
  wire       [31:0]   _zz_13871;
  wire       [15:0]   _zz_13872;
  wire       [31:0]   _zz_13873;
  wire       [31:0]   _zz_13874;
  wire       [31:0]   _zz_13875;
  wire       [15:0]   _zz_13876;
  wire       [31:0]   _zz_13877;
  wire       [31:0]   _zz_13878;
  wire       [31:0]   _zz_13879;
  wire       [31:0]   _zz_13880;
  wire       [31:0]   _zz_13881;
  wire       [31:0]   _zz_13882;
  wire       [23:0]   _zz_13883;
  wire       [31:0]   _zz_13884;
  wire       [15:0]   _zz_13885;
  wire       [31:0]   _zz_13886;
  wire       [31:0]   _zz_13887;
  wire       [31:0]   _zz_13888;
  wire       [31:0]   _zz_13889;
  wire       [31:0]   _zz_13890;
  wire       [23:0]   _zz_13891;
  wire       [31:0]   _zz_13892;
  wire       [15:0]   _zz_13893;
  wire       [31:0]   _zz_13894;
  wire       [31:0]   _zz_13895;
  wire       [31:0]   _zz_13896;
  wire       [31:0]   _zz_13897;
  wire       [31:0]   _zz_13898;
  wire       [23:0]   _zz_13899;
  wire       [31:0]   _zz_13900;
  wire       [15:0]   _zz_13901;
  wire       [31:0]   _zz_13902;
  wire       [31:0]   _zz_13903;
  wire       [31:0]   _zz_13904;
  wire       [31:0]   _zz_13905;
  wire       [31:0]   _zz_13906;
  wire       [23:0]   _zz_13907;
  wire       [31:0]   _zz_13908;
  wire       [15:0]   _zz_13909;
  wire       [15:0]   _zz_13910;
  wire       [31:0]   _zz_13911;
  wire       [31:0]   _zz_13912;
  wire       [15:0]   _zz_13913;
  wire       [31:0]   _zz_13914;
  wire       [31:0]   _zz_13915;
  wire       [31:0]   _zz_13916;
  wire       [15:0]   _zz_13917;
  wire       [31:0]   _zz_13918;
  wire       [31:0]   _zz_13919;
  wire       [31:0]   _zz_13920;
  wire       [31:0]   _zz_13921;
  wire       [31:0]   _zz_13922;
  wire       [31:0]   _zz_13923;
  wire       [23:0]   _zz_13924;
  wire       [31:0]   _zz_13925;
  wire       [15:0]   _zz_13926;
  wire       [31:0]   _zz_13927;
  wire       [31:0]   _zz_13928;
  wire       [31:0]   _zz_13929;
  wire       [31:0]   _zz_13930;
  wire       [31:0]   _zz_13931;
  wire       [23:0]   _zz_13932;
  wire       [31:0]   _zz_13933;
  wire       [15:0]   _zz_13934;
  wire       [31:0]   _zz_13935;
  wire       [31:0]   _zz_13936;
  wire       [31:0]   _zz_13937;
  wire       [31:0]   _zz_13938;
  wire       [31:0]   _zz_13939;
  wire       [23:0]   _zz_13940;
  wire       [31:0]   _zz_13941;
  wire       [15:0]   _zz_13942;
  wire       [31:0]   _zz_13943;
  wire       [31:0]   _zz_13944;
  wire       [31:0]   _zz_13945;
  wire       [31:0]   _zz_13946;
  wire       [31:0]   _zz_13947;
  wire       [23:0]   _zz_13948;
  wire       [31:0]   _zz_13949;
  wire       [15:0]   _zz_13950;
  wire       [15:0]   _zz_13951;
  wire       [31:0]   _zz_13952;
  wire       [31:0]   _zz_13953;
  wire       [15:0]   _zz_13954;
  wire       [31:0]   _zz_13955;
  wire       [31:0]   _zz_13956;
  wire       [31:0]   _zz_13957;
  wire       [15:0]   _zz_13958;
  wire       [31:0]   _zz_13959;
  wire       [31:0]   _zz_13960;
  wire       [31:0]   _zz_13961;
  wire       [31:0]   _zz_13962;
  wire       [31:0]   _zz_13963;
  wire       [31:0]   _zz_13964;
  wire       [23:0]   _zz_13965;
  wire       [31:0]   _zz_13966;
  wire       [15:0]   _zz_13967;
  wire       [31:0]   _zz_13968;
  wire       [31:0]   _zz_13969;
  wire       [31:0]   _zz_13970;
  wire       [31:0]   _zz_13971;
  wire       [31:0]   _zz_13972;
  wire       [23:0]   _zz_13973;
  wire       [31:0]   _zz_13974;
  wire       [15:0]   _zz_13975;
  wire       [31:0]   _zz_13976;
  wire       [31:0]   _zz_13977;
  wire       [31:0]   _zz_13978;
  wire       [31:0]   _zz_13979;
  wire       [31:0]   _zz_13980;
  wire       [23:0]   _zz_13981;
  wire       [31:0]   _zz_13982;
  wire       [15:0]   _zz_13983;
  wire       [31:0]   _zz_13984;
  wire       [31:0]   _zz_13985;
  wire       [31:0]   _zz_13986;
  wire       [31:0]   _zz_13987;
  wire       [31:0]   _zz_13988;
  wire       [23:0]   _zz_13989;
  wire       [31:0]   _zz_13990;
  wire       [15:0]   _zz_13991;
  wire       [15:0]   _zz_13992;
  wire       [31:0]   _zz_13993;
  wire       [31:0]   _zz_13994;
  wire       [15:0]   _zz_13995;
  wire       [31:0]   _zz_13996;
  wire       [31:0]   _zz_13997;
  wire       [31:0]   _zz_13998;
  wire       [15:0]   _zz_13999;
  wire       [31:0]   _zz_14000;
  wire       [31:0]   _zz_14001;
  wire       [31:0]   _zz_14002;
  wire       [31:0]   _zz_14003;
  wire       [31:0]   _zz_14004;
  wire       [31:0]   _zz_14005;
  wire       [23:0]   _zz_14006;
  wire       [31:0]   _zz_14007;
  wire       [15:0]   _zz_14008;
  wire       [31:0]   _zz_14009;
  wire       [31:0]   _zz_14010;
  wire       [31:0]   _zz_14011;
  wire       [31:0]   _zz_14012;
  wire       [31:0]   _zz_14013;
  wire       [23:0]   _zz_14014;
  wire       [31:0]   _zz_14015;
  wire       [15:0]   _zz_14016;
  wire       [31:0]   _zz_14017;
  wire       [31:0]   _zz_14018;
  wire       [31:0]   _zz_14019;
  wire       [31:0]   _zz_14020;
  wire       [31:0]   _zz_14021;
  wire       [23:0]   _zz_14022;
  wire       [31:0]   _zz_14023;
  wire       [15:0]   _zz_14024;
  wire       [31:0]   _zz_14025;
  wire       [31:0]   _zz_14026;
  wire       [31:0]   _zz_14027;
  wire       [31:0]   _zz_14028;
  wire       [31:0]   _zz_14029;
  wire       [23:0]   _zz_14030;
  wire       [31:0]   _zz_14031;
  wire       [15:0]   _zz_14032;
  wire       [15:0]   _zz_14033;
  wire       [31:0]   _zz_14034;
  wire       [31:0]   _zz_14035;
  wire       [15:0]   _zz_14036;
  wire       [31:0]   _zz_14037;
  wire       [31:0]   _zz_14038;
  wire       [31:0]   _zz_14039;
  wire       [15:0]   _zz_14040;
  wire       [31:0]   _zz_14041;
  wire       [31:0]   _zz_14042;
  wire       [31:0]   _zz_14043;
  wire       [31:0]   _zz_14044;
  wire       [31:0]   _zz_14045;
  wire       [31:0]   _zz_14046;
  wire       [23:0]   _zz_14047;
  wire       [31:0]   _zz_14048;
  wire       [15:0]   _zz_14049;
  wire       [31:0]   _zz_14050;
  wire       [31:0]   _zz_14051;
  wire       [31:0]   _zz_14052;
  wire       [31:0]   _zz_14053;
  wire       [31:0]   _zz_14054;
  wire       [23:0]   _zz_14055;
  wire       [31:0]   _zz_14056;
  wire       [15:0]   _zz_14057;
  wire       [31:0]   _zz_14058;
  wire       [31:0]   _zz_14059;
  wire       [31:0]   _zz_14060;
  wire       [31:0]   _zz_14061;
  wire       [31:0]   _zz_14062;
  wire       [23:0]   _zz_14063;
  wire       [31:0]   _zz_14064;
  wire       [15:0]   _zz_14065;
  wire       [31:0]   _zz_14066;
  wire       [31:0]   _zz_14067;
  wire       [31:0]   _zz_14068;
  wire       [31:0]   _zz_14069;
  wire       [31:0]   _zz_14070;
  wire       [23:0]   _zz_14071;
  wire       [31:0]   _zz_14072;
  wire       [15:0]   _zz_14073;
  wire       [15:0]   _zz_14074;
  wire       [31:0]   _zz_14075;
  wire       [31:0]   _zz_14076;
  wire       [15:0]   _zz_14077;
  wire       [31:0]   _zz_14078;
  wire       [31:0]   _zz_14079;
  wire       [31:0]   _zz_14080;
  wire       [15:0]   _zz_14081;
  wire       [31:0]   _zz_14082;
  wire       [31:0]   _zz_14083;
  wire       [31:0]   _zz_14084;
  wire       [31:0]   _zz_14085;
  wire       [31:0]   _zz_14086;
  wire       [31:0]   _zz_14087;
  wire       [23:0]   _zz_14088;
  wire       [31:0]   _zz_14089;
  wire       [15:0]   _zz_14090;
  wire       [31:0]   _zz_14091;
  wire       [31:0]   _zz_14092;
  wire       [31:0]   _zz_14093;
  wire       [31:0]   _zz_14094;
  wire       [31:0]   _zz_14095;
  wire       [23:0]   _zz_14096;
  wire       [31:0]   _zz_14097;
  wire       [15:0]   _zz_14098;
  wire       [31:0]   _zz_14099;
  wire       [31:0]   _zz_14100;
  wire       [31:0]   _zz_14101;
  wire       [31:0]   _zz_14102;
  wire       [31:0]   _zz_14103;
  wire       [23:0]   _zz_14104;
  wire       [31:0]   _zz_14105;
  wire       [15:0]   _zz_14106;
  wire       [31:0]   _zz_14107;
  wire       [31:0]   _zz_14108;
  wire       [31:0]   _zz_14109;
  wire       [31:0]   _zz_14110;
  wire       [31:0]   _zz_14111;
  wire       [23:0]   _zz_14112;
  wire       [31:0]   _zz_14113;
  wire       [15:0]   _zz_14114;
  wire       [15:0]   _zz_14115;
  wire       [31:0]   _zz_14116;
  wire       [31:0]   _zz_14117;
  wire       [15:0]   _zz_14118;
  wire       [31:0]   _zz_14119;
  wire       [31:0]   _zz_14120;
  wire       [31:0]   _zz_14121;
  wire       [15:0]   _zz_14122;
  wire       [31:0]   _zz_14123;
  wire       [31:0]   _zz_14124;
  wire       [31:0]   _zz_14125;
  wire       [31:0]   _zz_14126;
  wire       [31:0]   _zz_14127;
  wire       [31:0]   _zz_14128;
  wire       [23:0]   _zz_14129;
  wire       [31:0]   _zz_14130;
  wire       [15:0]   _zz_14131;
  wire       [31:0]   _zz_14132;
  wire       [31:0]   _zz_14133;
  wire       [31:0]   _zz_14134;
  wire       [31:0]   _zz_14135;
  wire       [31:0]   _zz_14136;
  wire       [23:0]   _zz_14137;
  wire       [31:0]   _zz_14138;
  wire       [15:0]   _zz_14139;
  wire       [31:0]   _zz_14140;
  wire       [31:0]   _zz_14141;
  wire       [31:0]   _zz_14142;
  wire       [31:0]   _zz_14143;
  wire       [31:0]   _zz_14144;
  wire       [23:0]   _zz_14145;
  wire       [31:0]   _zz_14146;
  wire       [15:0]   _zz_14147;
  wire       [31:0]   _zz_14148;
  wire       [31:0]   _zz_14149;
  wire       [31:0]   _zz_14150;
  wire       [31:0]   _zz_14151;
  wire       [31:0]   _zz_14152;
  wire       [23:0]   _zz_14153;
  wire       [31:0]   _zz_14154;
  wire       [15:0]   _zz_14155;
  wire       [15:0]   _zz_14156;
  wire       [31:0]   _zz_14157;
  wire       [31:0]   _zz_14158;
  wire       [15:0]   _zz_14159;
  wire       [31:0]   _zz_14160;
  wire       [31:0]   _zz_14161;
  wire       [31:0]   _zz_14162;
  wire       [15:0]   _zz_14163;
  wire       [31:0]   _zz_14164;
  wire       [31:0]   _zz_14165;
  wire       [31:0]   _zz_14166;
  wire       [31:0]   _zz_14167;
  wire       [31:0]   _zz_14168;
  wire       [31:0]   _zz_14169;
  wire       [23:0]   _zz_14170;
  wire       [31:0]   _zz_14171;
  wire       [15:0]   _zz_14172;
  wire       [31:0]   _zz_14173;
  wire       [31:0]   _zz_14174;
  wire       [31:0]   _zz_14175;
  wire       [31:0]   _zz_14176;
  wire       [31:0]   _zz_14177;
  wire       [23:0]   _zz_14178;
  wire       [31:0]   _zz_14179;
  wire       [15:0]   _zz_14180;
  wire       [31:0]   _zz_14181;
  wire       [31:0]   _zz_14182;
  wire       [31:0]   _zz_14183;
  wire       [31:0]   _zz_14184;
  wire       [31:0]   _zz_14185;
  wire       [23:0]   _zz_14186;
  wire       [31:0]   _zz_14187;
  wire       [15:0]   _zz_14188;
  wire       [31:0]   _zz_14189;
  wire       [31:0]   _zz_14190;
  wire       [31:0]   _zz_14191;
  wire       [31:0]   _zz_14192;
  wire       [31:0]   _zz_14193;
  wire       [23:0]   _zz_14194;
  wire       [31:0]   _zz_14195;
  wire       [15:0]   _zz_14196;
  wire       [15:0]   _zz_14197;
  wire       [31:0]   _zz_14198;
  wire       [31:0]   _zz_14199;
  wire       [15:0]   _zz_14200;
  wire       [31:0]   _zz_14201;
  wire       [31:0]   _zz_14202;
  wire       [31:0]   _zz_14203;
  wire       [15:0]   _zz_14204;
  wire       [31:0]   _zz_14205;
  wire       [31:0]   _zz_14206;
  wire       [31:0]   _zz_14207;
  wire       [31:0]   _zz_14208;
  wire       [31:0]   _zz_14209;
  wire       [31:0]   _zz_14210;
  wire       [23:0]   _zz_14211;
  wire       [31:0]   _zz_14212;
  wire       [15:0]   _zz_14213;
  wire       [31:0]   _zz_14214;
  wire       [31:0]   _zz_14215;
  wire       [31:0]   _zz_14216;
  wire       [31:0]   _zz_14217;
  wire       [31:0]   _zz_14218;
  wire       [23:0]   _zz_14219;
  wire       [31:0]   _zz_14220;
  wire       [15:0]   _zz_14221;
  wire       [31:0]   _zz_14222;
  wire       [31:0]   _zz_14223;
  wire       [31:0]   _zz_14224;
  wire       [31:0]   _zz_14225;
  wire       [31:0]   _zz_14226;
  wire       [23:0]   _zz_14227;
  wire       [31:0]   _zz_14228;
  wire       [15:0]   _zz_14229;
  wire       [31:0]   _zz_14230;
  wire       [31:0]   _zz_14231;
  wire       [31:0]   _zz_14232;
  wire       [31:0]   _zz_14233;
  wire       [31:0]   _zz_14234;
  wire       [23:0]   _zz_14235;
  wire       [31:0]   _zz_14236;
  wire       [15:0]   _zz_14237;
  wire       [15:0]   _zz_14238;
  wire       [31:0]   _zz_14239;
  wire       [31:0]   _zz_14240;
  wire       [15:0]   _zz_14241;
  wire       [31:0]   _zz_14242;
  wire       [31:0]   _zz_14243;
  wire       [31:0]   _zz_14244;
  wire       [15:0]   _zz_14245;
  wire       [31:0]   _zz_14246;
  wire       [31:0]   _zz_14247;
  wire       [31:0]   _zz_14248;
  wire       [31:0]   _zz_14249;
  wire       [31:0]   _zz_14250;
  wire       [31:0]   _zz_14251;
  wire       [23:0]   _zz_14252;
  wire       [31:0]   _zz_14253;
  wire       [15:0]   _zz_14254;
  wire       [31:0]   _zz_14255;
  wire       [31:0]   _zz_14256;
  wire       [31:0]   _zz_14257;
  wire       [31:0]   _zz_14258;
  wire       [31:0]   _zz_14259;
  wire       [23:0]   _zz_14260;
  wire       [31:0]   _zz_14261;
  wire       [15:0]   _zz_14262;
  wire       [31:0]   _zz_14263;
  wire       [31:0]   _zz_14264;
  wire       [31:0]   _zz_14265;
  wire       [31:0]   _zz_14266;
  wire       [31:0]   _zz_14267;
  wire       [23:0]   _zz_14268;
  wire       [31:0]   _zz_14269;
  wire       [15:0]   _zz_14270;
  wire       [31:0]   _zz_14271;
  wire       [31:0]   _zz_14272;
  wire       [31:0]   _zz_14273;
  wire       [31:0]   _zz_14274;
  wire       [31:0]   _zz_14275;
  wire       [23:0]   _zz_14276;
  wire       [31:0]   _zz_14277;
  wire       [15:0]   _zz_14278;
  wire       [15:0]   _zz_14279;
  wire       [31:0]   _zz_14280;
  wire       [31:0]   _zz_14281;
  wire       [15:0]   _zz_14282;
  wire       [31:0]   _zz_14283;
  wire       [31:0]   _zz_14284;
  wire       [31:0]   _zz_14285;
  wire       [15:0]   _zz_14286;
  wire       [31:0]   _zz_14287;
  wire       [31:0]   _zz_14288;
  wire       [31:0]   _zz_14289;
  wire       [31:0]   _zz_14290;
  wire       [31:0]   _zz_14291;
  wire       [31:0]   _zz_14292;
  wire       [23:0]   _zz_14293;
  wire       [31:0]   _zz_14294;
  wire       [15:0]   _zz_14295;
  wire       [31:0]   _zz_14296;
  wire       [31:0]   _zz_14297;
  wire       [31:0]   _zz_14298;
  wire       [31:0]   _zz_14299;
  wire       [31:0]   _zz_14300;
  wire       [23:0]   _zz_14301;
  wire       [31:0]   _zz_14302;
  wire       [15:0]   _zz_14303;
  wire       [31:0]   _zz_14304;
  wire       [31:0]   _zz_14305;
  wire       [31:0]   _zz_14306;
  wire       [31:0]   _zz_14307;
  wire       [31:0]   _zz_14308;
  wire       [23:0]   _zz_14309;
  wire       [31:0]   _zz_14310;
  wire       [15:0]   _zz_14311;
  wire       [31:0]   _zz_14312;
  wire       [31:0]   _zz_14313;
  wire       [31:0]   _zz_14314;
  wire       [31:0]   _zz_14315;
  wire       [31:0]   _zz_14316;
  wire       [23:0]   _zz_14317;
  wire       [31:0]   _zz_14318;
  wire       [15:0]   _zz_14319;
  wire       [15:0]   _zz_14320;
  wire       [31:0]   _zz_14321;
  wire       [31:0]   _zz_14322;
  wire       [15:0]   _zz_14323;
  wire       [31:0]   _zz_14324;
  wire       [31:0]   _zz_14325;
  wire       [31:0]   _zz_14326;
  wire       [15:0]   _zz_14327;
  wire       [31:0]   _zz_14328;
  wire       [31:0]   _zz_14329;
  wire       [31:0]   _zz_14330;
  wire       [31:0]   _zz_14331;
  wire       [31:0]   _zz_14332;
  wire       [31:0]   _zz_14333;
  wire       [23:0]   _zz_14334;
  wire       [31:0]   _zz_14335;
  wire       [15:0]   _zz_14336;
  wire       [31:0]   _zz_14337;
  wire       [31:0]   _zz_14338;
  wire       [31:0]   _zz_14339;
  wire       [31:0]   _zz_14340;
  wire       [31:0]   _zz_14341;
  wire       [23:0]   _zz_14342;
  wire       [31:0]   _zz_14343;
  wire       [15:0]   _zz_14344;
  wire       [31:0]   _zz_14345;
  wire       [31:0]   _zz_14346;
  wire       [31:0]   _zz_14347;
  wire       [31:0]   _zz_14348;
  wire       [31:0]   _zz_14349;
  wire       [23:0]   _zz_14350;
  wire       [31:0]   _zz_14351;
  wire       [15:0]   _zz_14352;
  wire       [31:0]   _zz_14353;
  wire       [31:0]   _zz_14354;
  wire       [31:0]   _zz_14355;
  wire       [31:0]   _zz_14356;
  wire       [31:0]   _zz_14357;
  wire       [23:0]   _zz_14358;
  wire       [31:0]   _zz_14359;
  wire       [15:0]   _zz_14360;
  wire       [15:0]   _zz_14361;
  wire       [31:0]   _zz_14362;
  wire       [31:0]   _zz_14363;
  wire       [15:0]   _zz_14364;
  wire       [31:0]   _zz_14365;
  wire       [31:0]   _zz_14366;
  wire       [31:0]   _zz_14367;
  wire       [15:0]   _zz_14368;
  wire       [31:0]   _zz_14369;
  wire       [31:0]   _zz_14370;
  wire       [31:0]   _zz_14371;
  wire       [31:0]   _zz_14372;
  wire       [31:0]   _zz_14373;
  wire       [31:0]   _zz_14374;
  wire       [23:0]   _zz_14375;
  wire       [31:0]   _zz_14376;
  wire       [15:0]   _zz_14377;
  wire       [31:0]   _zz_14378;
  wire       [31:0]   _zz_14379;
  wire       [31:0]   _zz_14380;
  wire       [31:0]   _zz_14381;
  wire       [31:0]   _zz_14382;
  wire       [23:0]   _zz_14383;
  wire       [31:0]   _zz_14384;
  wire       [15:0]   _zz_14385;
  wire       [31:0]   _zz_14386;
  wire       [31:0]   _zz_14387;
  wire       [31:0]   _zz_14388;
  wire       [31:0]   _zz_14389;
  wire       [31:0]   _zz_14390;
  wire       [23:0]   _zz_14391;
  wire       [31:0]   _zz_14392;
  wire       [15:0]   _zz_14393;
  wire       [31:0]   _zz_14394;
  wire       [31:0]   _zz_14395;
  wire       [31:0]   _zz_14396;
  wire       [31:0]   _zz_14397;
  wire       [31:0]   _zz_14398;
  wire       [23:0]   _zz_14399;
  wire       [31:0]   _zz_14400;
  wire       [15:0]   _zz_14401;
  wire       [15:0]   _zz_14402;
  wire       [31:0]   _zz_14403;
  wire       [31:0]   _zz_14404;
  wire       [15:0]   _zz_14405;
  wire       [31:0]   _zz_14406;
  wire       [31:0]   _zz_14407;
  wire       [31:0]   _zz_14408;
  wire       [15:0]   _zz_14409;
  wire       [31:0]   _zz_14410;
  wire       [31:0]   _zz_14411;
  wire       [31:0]   _zz_14412;
  wire       [31:0]   _zz_14413;
  wire       [31:0]   _zz_14414;
  wire       [31:0]   _zz_14415;
  wire       [23:0]   _zz_14416;
  wire       [31:0]   _zz_14417;
  wire       [15:0]   _zz_14418;
  wire       [31:0]   _zz_14419;
  wire       [31:0]   _zz_14420;
  wire       [31:0]   _zz_14421;
  wire       [31:0]   _zz_14422;
  wire       [31:0]   _zz_14423;
  wire       [23:0]   _zz_14424;
  wire       [31:0]   _zz_14425;
  wire       [15:0]   _zz_14426;
  wire       [31:0]   _zz_14427;
  wire       [31:0]   _zz_14428;
  wire       [31:0]   _zz_14429;
  wire       [31:0]   _zz_14430;
  wire       [31:0]   _zz_14431;
  wire       [23:0]   _zz_14432;
  wire       [31:0]   _zz_14433;
  wire       [15:0]   _zz_14434;
  wire       [31:0]   _zz_14435;
  wire       [31:0]   _zz_14436;
  wire       [31:0]   _zz_14437;
  wire       [31:0]   _zz_14438;
  wire       [31:0]   _zz_14439;
  wire       [23:0]   _zz_14440;
  wire       [31:0]   _zz_14441;
  wire       [15:0]   _zz_14442;
  wire       [15:0]   _zz_14443;
  wire       [31:0]   _zz_14444;
  wire       [31:0]   _zz_14445;
  wire       [15:0]   _zz_14446;
  wire       [31:0]   _zz_14447;
  wire       [31:0]   _zz_14448;
  wire       [31:0]   _zz_14449;
  wire       [15:0]   _zz_14450;
  wire       [31:0]   _zz_14451;
  wire       [31:0]   _zz_14452;
  wire       [31:0]   _zz_14453;
  wire       [31:0]   _zz_14454;
  wire       [31:0]   _zz_14455;
  wire       [31:0]   _zz_14456;
  wire       [23:0]   _zz_14457;
  wire       [31:0]   _zz_14458;
  wire       [15:0]   _zz_14459;
  wire       [31:0]   _zz_14460;
  wire       [31:0]   _zz_14461;
  wire       [31:0]   _zz_14462;
  wire       [31:0]   _zz_14463;
  wire       [31:0]   _zz_14464;
  wire       [23:0]   _zz_14465;
  wire       [31:0]   _zz_14466;
  wire       [15:0]   _zz_14467;
  wire       [31:0]   _zz_14468;
  wire       [31:0]   _zz_14469;
  wire       [31:0]   _zz_14470;
  wire       [31:0]   _zz_14471;
  wire       [31:0]   _zz_14472;
  wire       [23:0]   _zz_14473;
  wire       [31:0]   _zz_14474;
  wire       [15:0]   _zz_14475;
  wire       [31:0]   _zz_14476;
  wire       [31:0]   _zz_14477;
  wire       [31:0]   _zz_14478;
  wire       [31:0]   _zz_14479;
  wire       [31:0]   _zz_14480;
  wire       [23:0]   _zz_14481;
  wire       [31:0]   _zz_14482;
  wire       [15:0]   _zz_14483;
  wire       [15:0]   _zz_14484;
  wire       [31:0]   _zz_14485;
  wire       [31:0]   _zz_14486;
  wire       [15:0]   _zz_14487;
  wire       [31:0]   _zz_14488;
  wire       [31:0]   _zz_14489;
  wire       [31:0]   _zz_14490;
  wire       [15:0]   _zz_14491;
  wire       [31:0]   _zz_14492;
  wire       [31:0]   _zz_14493;
  wire       [31:0]   _zz_14494;
  wire       [31:0]   _zz_14495;
  wire       [31:0]   _zz_14496;
  wire       [31:0]   _zz_14497;
  wire       [23:0]   _zz_14498;
  wire       [31:0]   _zz_14499;
  wire       [15:0]   _zz_14500;
  wire       [31:0]   _zz_14501;
  wire       [31:0]   _zz_14502;
  wire       [31:0]   _zz_14503;
  wire       [31:0]   _zz_14504;
  wire       [31:0]   _zz_14505;
  wire       [23:0]   _zz_14506;
  wire       [31:0]   _zz_14507;
  wire       [15:0]   _zz_14508;
  wire       [31:0]   _zz_14509;
  wire       [31:0]   _zz_14510;
  wire       [31:0]   _zz_14511;
  wire       [31:0]   _zz_14512;
  wire       [31:0]   _zz_14513;
  wire       [23:0]   _zz_14514;
  wire       [31:0]   _zz_14515;
  wire       [15:0]   _zz_14516;
  wire       [31:0]   _zz_14517;
  wire       [31:0]   _zz_14518;
  wire       [31:0]   _zz_14519;
  wire       [31:0]   _zz_14520;
  wire       [31:0]   _zz_14521;
  wire       [23:0]   _zz_14522;
  wire       [31:0]   _zz_14523;
  wire       [15:0]   _zz_14524;
  wire       [15:0]   _zz_14525;
  wire       [31:0]   _zz_14526;
  wire       [31:0]   _zz_14527;
  wire       [15:0]   _zz_14528;
  wire       [31:0]   _zz_14529;
  wire       [31:0]   _zz_14530;
  wire       [31:0]   _zz_14531;
  wire       [15:0]   _zz_14532;
  wire       [31:0]   _zz_14533;
  wire       [31:0]   _zz_14534;
  wire       [31:0]   _zz_14535;
  wire       [31:0]   _zz_14536;
  wire       [31:0]   _zz_14537;
  wire       [31:0]   _zz_14538;
  wire       [23:0]   _zz_14539;
  wire       [31:0]   _zz_14540;
  wire       [15:0]   _zz_14541;
  wire       [31:0]   _zz_14542;
  wire       [31:0]   _zz_14543;
  wire       [31:0]   _zz_14544;
  wire       [31:0]   _zz_14545;
  wire       [31:0]   _zz_14546;
  wire       [23:0]   _zz_14547;
  wire       [31:0]   _zz_14548;
  wire       [15:0]   _zz_14549;
  wire       [31:0]   _zz_14550;
  wire       [31:0]   _zz_14551;
  wire       [31:0]   _zz_14552;
  wire       [31:0]   _zz_14553;
  wire       [31:0]   _zz_14554;
  wire       [23:0]   _zz_14555;
  wire       [31:0]   _zz_14556;
  wire       [15:0]   _zz_14557;
  wire       [31:0]   _zz_14558;
  wire       [31:0]   _zz_14559;
  wire       [31:0]   _zz_14560;
  wire       [31:0]   _zz_14561;
  wire       [31:0]   _zz_14562;
  wire       [23:0]   _zz_14563;
  wire       [31:0]   _zz_14564;
  wire       [15:0]   _zz_14565;
  wire       [15:0]   _zz_14566;
  wire       [31:0]   _zz_14567;
  wire       [31:0]   _zz_14568;
  wire       [15:0]   _zz_14569;
  wire       [31:0]   _zz_14570;
  wire       [31:0]   _zz_14571;
  wire       [31:0]   _zz_14572;
  wire       [15:0]   _zz_14573;
  wire       [31:0]   _zz_14574;
  wire       [31:0]   _zz_14575;
  wire       [31:0]   _zz_14576;
  wire       [31:0]   _zz_14577;
  wire       [31:0]   _zz_14578;
  wire       [31:0]   _zz_14579;
  wire       [23:0]   _zz_14580;
  wire       [31:0]   _zz_14581;
  wire       [15:0]   _zz_14582;
  wire       [31:0]   _zz_14583;
  wire       [31:0]   _zz_14584;
  wire       [31:0]   _zz_14585;
  wire       [31:0]   _zz_14586;
  wire       [31:0]   _zz_14587;
  wire       [23:0]   _zz_14588;
  wire       [31:0]   _zz_14589;
  wire       [15:0]   _zz_14590;
  wire       [31:0]   _zz_14591;
  wire       [31:0]   _zz_14592;
  wire       [31:0]   _zz_14593;
  wire       [31:0]   _zz_14594;
  wire       [31:0]   _zz_14595;
  wire       [23:0]   _zz_14596;
  wire       [31:0]   _zz_14597;
  wire       [15:0]   _zz_14598;
  wire       [31:0]   _zz_14599;
  wire       [31:0]   _zz_14600;
  wire       [31:0]   _zz_14601;
  wire       [31:0]   _zz_14602;
  wire       [31:0]   _zz_14603;
  wire       [23:0]   _zz_14604;
  wire       [31:0]   _zz_14605;
  wire       [15:0]   _zz_14606;
  wire       [15:0]   _zz_14607;
  wire       [31:0]   _zz_14608;
  wire       [31:0]   _zz_14609;
  wire       [15:0]   _zz_14610;
  wire       [31:0]   _zz_14611;
  wire       [31:0]   _zz_14612;
  wire       [31:0]   _zz_14613;
  wire       [15:0]   _zz_14614;
  wire       [31:0]   _zz_14615;
  wire       [31:0]   _zz_14616;
  wire       [31:0]   _zz_14617;
  wire       [31:0]   _zz_14618;
  wire       [31:0]   _zz_14619;
  wire       [31:0]   _zz_14620;
  wire       [23:0]   _zz_14621;
  wire       [31:0]   _zz_14622;
  wire       [15:0]   _zz_14623;
  wire       [31:0]   _zz_14624;
  wire       [31:0]   _zz_14625;
  wire       [31:0]   _zz_14626;
  wire       [31:0]   _zz_14627;
  wire       [31:0]   _zz_14628;
  wire       [23:0]   _zz_14629;
  wire       [31:0]   _zz_14630;
  wire       [15:0]   _zz_14631;
  wire       [31:0]   _zz_14632;
  wire       [31:0]   _zz_14633;
  wire       [31:0]   _zz_14634;
  wire       [31:0]   _zz_14635;
  wire       [31:0]   _zz_14636;
  wire       [23:0]   _zz_14637;
  wire       [31:0]   _zz_14638;
  wire       [15:0]   _zz_14639;
  wire       [31:0]   _zz_14640;
  wire       [31:0]   _zz_14641;
  wire       [31:0]   _zz_14642;
  wire       [31:0]   _zz_14643;
  wire       [31:0]   _zz_14644;
  wire       [23:0]   _zz_14645;
  wire       [31:0]   _zz_14646;
  wire       [15:0]   _zz_14647;
  wire       [15:0]   _zz_14648;
  wire       [31:0]   _zz_14649;
  wire       [31:0]   _zz_14650;
  wire       [15:0]   _zz_14651;
  wire       [31:0]   _zz_14652;
  wire       [31:0]   _zz_14653;
  wire       [31:0]   _zz_14654;
  wire       [15:0]   _zz_14655;
  wire       [31:0]   _zz_14656;
  wire       [31:0]   _zz_14657;
  wire       [31:0]   _zz_14658;
  wire       [31:0]   _zz_14659;
  wire       [31:0]   _zz_14660;
  wire       [31:0]   _zz_14661;
  wire       [23:0]   _zz_14662;
  wire       [31:0]   _zz_14663;
  wire       [15:0]   _zz_14664;
  wire       [31:0]   _zz_14665;
  wire       [31:0]   _zz_14666;
  wire       [31:0]   _zz_14667;
  wire       [31:0]   _zz_14668;
  wire       [31:0]   _zz_14669;
  wire       [23:0]   _zz_14670;
  wire       [31:0]   _zz_14671;
  wire       [15:0]   _zz_14672;
  wire       [31:0]   _zz_14673;
  wire       [31:0]   _zz_14674;
  wire       [31:0]   _zz_14675;
  wire       [31:0]   _zz_14676;
  wire       [31:0]   _zz_14677;
  wire       [23:0]   _zz_14678;
  wire       [31:0]   _zz_14679;
  wire       [15:0]   _zz_14680;
  wire       [31:0]   _zz_14681;
  wire       [31:0]   _zz_14682;
  wire       [31:0]   _zz_14683;
  wire       [31:0]   _zz_14684;
  wire       [31:0]   _zz_14685;
  wire       [23:0]   _zz_14686;
  wire       [31:0]   _zz_14687;
  wire       [15:0]   _zz_14688;
  wire       [15:0]   _zz_14689;
  wire       [31:0]   _zz_14690;
  wire       [31:0]   _zz_14691;
  wire       [15:0]   _zz_14692;
  wire       [31:0]   _zz_14693;
  wire       [31:0]   _zz_14694;
  wire       [31:0]   _zz_14695;
  wire       [15:0]   _zz_14696;
  wire       [31:0]   _zz_14697;
  wire       [31:0]   _zz_14698;
  wire       [31:0]   _zz_14699;
  wire       [31:0]   _zz_14700;
  wire       [31:0]   _zz_14701;
  wire       [31:0]   _zz_14702;
  wire       [23:0]   _zz_14703;
  wire       [31:0]   _zz_14704;
  wire       [15:0]   _zz_14705;
  wire       [31:0]   _zz_14706;
  wire       [31:0]   _zz_14707;
  wire       [31:0]   _zz_14708;
  wire       [31:0]   _zz_14709;
  wire       [31:0]   _zz_14710;
  wire       [23:0]   _zz_14711;
  wire       [31:0]   _zz_14712;
  wire       [15:0]   _zz_14713;
  wire       [31:0]   _zz_14714;
  wire       [31:0]   _zz_14715;
  wire       [31:0]   _zz_14716;
  wire       [31:0]   _zz_14717;
  wire       [31:0]   _zz_14718;
  wire       [23:0]   _zz_14719;
  wire       [31:0]   _zz_14720;
  wire       [15:0]   _zz_14721;
  wire       [31:0]   _zz_14722;
  wire       [31:0]   _zz_14723;
  wire       [31:0]   _zz_14724;
  wire       [31:0]   _zz_14725;
  wire       [31:0]   _zz_14726;
  wire       [23:0]   _zz_14727;
  wire       [31:0]   _zz_14728;
  wire       [15:0]   _zz_14729;
  wire       [15:0]   _zz_14730;
  wire       [31:0]   _zz_14731;
  wire       [31:0]   _zz_14732;
  wire       [15:0]   _zz_14733;
  wire       [31:0]   _zz_14734;
  wire       [31:0]   _zz_14735;
  wire       [31:0]   _zz_14736;
  wire       [15:0]   _zz_14737;
  wire       [31:0]   _zz_14738;
  wire       [31:0]   _zz_14739;
  wire       [31:0]   _zz_14740;
  wire       [31:0]   _zz_14741;
  wire       [31:0]   _zz_14742;
  wire       [31:0]   _zz_14743;
  wire       [23:0]   _zz_14744;
  wire       [31:0]   _zz_14745;
  wire       [15:0]   _zz_14746;
  wire       [31:0]   _zz_14747;
  wire       [31:0]   _zz_14748;
  wire       [31:0]   _zz_14749;
  wire       [31:0]   _zz_14750;
  wire       [31:0]   _zz_14751;
  wire       [23:0]   _zz_14752;
  wire       [31:0]   _zz_14753;
  wire       [15:0]   _zz_14754;
  wire       [31:0]   _zz_14755;
  wire       [31:0]   _zz_14756;
  wire       [31:0]   _zz_14757;
  wire       [31:0]   _zz_14758;
  wire       [31:0]   _zz_14759;
  wire       [23:0]   _zz_14760;
  wire       [31:0]   _zz_14761;
  wire       [15:0]   _zz_14762;
  wire       [31:0]   _zz_14763;
  wire       [31:0]   _zz_14764;
  wire       [31:0]   _zz_14765;
  wire       [31:0]   _zz_14766;
  wire       [31:0]   _zz_14767;
  wire       [23:0]   _zz_14768;
  wire       [31:0]   _zz_14769;
  wire       [15:0]   _zz_14770;
  wire       [15:0]   _zz_14771;
  wire       [31:0]   _zz_14772;
  wire       [31:0]   _zz_14773;
  wire       [15:0]   _zz_14774;
  wire       [31:0]   _zz_14775;
  wire       [31:0]   _zz_14776;
  wire       [31:0]   _zz_14777;
  wire       [15:0]   _zz_14778;
  wire       [31:0]   _zz_14779;
  wire       [31:0]   _zz_14780;
  wire       [31:0]   _zz_14781;
  wire       [31:0]   _zz_14782;
  wire       [31:0]   _zz_14783;
  wire       [31:0]   _zz_14784;
  wire       [23:0]   _zz_14785;
  wire       [31:0]   _zz_14786;
  wire       [15:0]   _zz_14787;
  wire       [31:0]   _zz_14788;
  wire       [31:0]   _zz_14789;
  wire       [31:0]   _zz_14790;
  wire       [31:0]   _zz_14791;
  wire       [31:0]   _zz_14792;
  wire       [23:0]   _zz_14793;
  wire       [31:0]   _zz_14794;
  wire       [15:0]   _zz_14795;
  wire       [31:0]   _zz_14796;
  wire       [31:0]   _zz_14797;
  wire       [31:0]   _zz_14798;
  wire       [31:0]   _zz_14799;
  wire       [31:0]   _zz_14800;
  wire       [23:0]   _zz_14801;
  wire       [31:0]   _zz_14802;
  wire       [15:0]   _zz_14803;
  wire       [31:0]   _zz_14804;
  wire       [31:0]   _zz_14805;
  wire       [31:0]   _zz_14806;
  wire       [31:0]   _zz_14807;
  wire       [31:0]   _zz_14808;
  wire       [23:0]   _zz_14809;
  wire       [31:0]   _zz_14810;
  wire       [15:0]   _zz_14811;
  wire       [15:0]   _zz_14812;
  wire       [31:0]   _zz_14813;
  wire       [31:0]   _zz_14814;
  wire       [15:0]   _zz_14815;
  wire       [31:0]   _zz_14816;
  wire       [31:0]   _zz_14817;
  wire       [31:0]   _zz_14818;
  wire       [15:0]   _zz_14819;
  wire       [31:0]   _zz_14820;
  wire       [31:0]   _zz_14821;
  wire       [31:0]   _zz_14822;
  wire       [31:0]   _zz_14823;
  wire       [31:0]   _zz_14824;
  wire       [31:0]   _zz_14825;
  wire       [23:0]   _zz_14826;
  wire       [31:0]   _zz_14827;
  wire       [15:0]   _zz_14828;
  wire       [31:0]   _zz_14829;
  wire       [31:0]   _zz_14830;
  wire       [31:0]   _zz_14831;
  wire       [31:0]   _zz_14832;
  wire       [31:0]   _zz_14833;
  wire       [23:0]   _zz_14834;
  wire       [31:0]   _zz_14835;
  wire       [15:0]   _zz_14836;
  wire       [31:0]   _zz_14837;
  wire       [31:0]   _zz_14838;
  wire       [31:0]   _zz_14839;
  wire       [31:0]   _zz_14840;
  wire       [31:0]   _zz_14841;
  wire       [23:0]   _zz_14842;
  wire       [31:0]   _zz_14843;
  wire       [15:0]   _zz_14844;
  wire       [31:0]   _zz_14845;
  wire       [31:0]   _zz_14846;
  wire       [31:0]   _zz_14847;
  wire       [31:0]   _zz_14848;
  wire       [31:0]   _zz_14849;
  wire       [23:0]   _zz_14850;
  wire       [31:0]   _zz_14851;
  wire       [15:0]   _zz_14852;
  wire       [15:0]   _zz_14853;
  wire       [31:0]   _zz_14854;
  wire       [31:0]   _zz_14855;
  wire       [15:0]   _zz_14856;
  wire       [31:0]   _zz_14857;
  wire       [31:0]   _zz_14858;
  wire       [31:0]   _zz_14859;
  wire       [15:0]   _zz_14860;
  wire       [31:0]   _zz_14861;
  wire       [31:0]   _zz_14862;
  wire       [31:0]   _zz_14863;
  wire       [31:0]   _zz_14864;
  wire       [31:0]   _zz_14865;
  wire       [31:0]   _zz_14866;
  wire       [23:0]   _zz_14867;
  wire       [31:0]   _zz_14868;
  wire       [15:0]   _zz_14869;
  wire       [31:0]   _zz_14870;
  wire       [31:0]   _zz_14871;
  wire       [31:0]   _zz_14872;
  wire       [31:0]   _zz_14873;
  wire       [31:0]   _zz_14874;
  wire       [23:0]   _zz_14875;
  wire       [31:0]   _zz_14876;
  wire       [15:0]   _zz_14877;
  wire       [31:0]   _zz_14878;
  wire       [31:0]   _zz_14879;
  wire       [31:0]   _zz_14880;
  wire       [31:0]   _zz_14881;
  wire       [31:0]   _zz_14882;
  wire       [23:0]   _zz_14883;
  wire       [31:0]   _zz_14884;
  wire       [15:0]   _zz_14885;
  wire       [31:0]   _zz_14886;
  wire       [31:0]   _zz_14887;
  wire       [31:0]   _zz_14888;
  wire       [31:0]   _zz_14889;
  wire       [31:0]   _zz_14890;
  wire       [23:0]   _zz_14891;
  wire       [31:0]   _zz_14892;
  wire       [15:0]   _zz_14893;
  wire       [15:0]   _zz_14894;
  wire       [31:0]   _zz_14895;
  wire       [31:0]   _zz_14896;
  wire       [15:0]   _zz_14897;
  wire       [31:0]   _zz_14898;
  wire       [31:0]   _zz_14899;
  wire       [31:0]   _zz_14900;
  wire       [15:0]   _zz_14901;
  wire       [31:0]   _zz_14902;
  wire       [31:0]   _zz_14903;
  wire       [31:0]   _zz_14904;
  wire       [31:0]   _zz_14905;
  wire       [31:0]   _zz_14906;
  wire       [31:0]   _zz_14907;
  wire       [23:0]   _zz_14908;
  wire       [31:0]   _zz_14909;
  wire       [15:0]   _zz_14910;
  wire       [31:0]   _zz_14911;
  wire       [31:0]   _zz_14912;
  wire       [31:0]   _zz_14913;
  wire       [31:0]   _zz_14914;
  wire       [31:0]   _zz_14915;
  wire       [23:0]   _zz_14916;
  wire       [31:0]   _zz_14917;
  wire       [15:0]   _zz_14918;
  wire       [31:0]   _zz_14919;
  wire       [31:0]   _zz_14920;
  wire       [31:0]   _zz_14921;
  wire       [31:0]   _zz_14922;
  wire       [31:0]   _zz_14923;
  wire       [23:0]   _zz_14924;
  wire       [31:0]   _zz_14925;
  wire       [15:0]   _zz_14926;
  wire       [31:0]   _zz_14927;
  wire       [31:0]   _zz_14928;
  wire       [31:0]   _zz_14929;
  wire       [31:0]   _zz_14930;
  wire       [31:0]   _zz_14931;
  wire       [23:0]   _zz_14932;
  wire       [31:0]   _zz_14933;
  wire       [15:0]   _zz_14934;
  wire       [15:0]   _zz_14935;
  wire       [31:0]   _zz_14936;
  wire       [31:0]   _zz_14937;
  wire       [15:0]   _zz_14938;
  wire       [31:0]   _zz_14939;
  wire       [31:0]   _zz_14940;
  wire       [31:0]   _zz_14941;
  wire       [15:0]   _zz_14942;
  wire       [31:0]   _zz_14943;
  wire       [31:0]   _zz_14944;
  wire       [31:0]   _zz_14945;
  wire       [31:0]   _zz_14946;
  wire       [31:0]   _zz_14947;
  wire       [31:0]   _zz_14948;
  wire       [23:0]   _zz_14949;
  wire       [31:0]   _zz_14950;
  wire       [15:0]   _zz_14951;
  wire       [31:0]   _zz_14952;
  wire       [31:0]   _zz_14953;
  wire       [31:0]   _zz_14954;
  wire       [31:0]   _zz_14955;
  wire       [31:0]   _zz_14956;
  wire       [23:0]   _zz_14957;
  wire       [31:0]   _zz_14958;
  wire       [15:0]   _zz_14959;
  wire       [31:0]   _zz_14960;
  wire       [31:0]   _zz_14961;
  wire       [31:0]   _zz_14962;
  wire       [31:0]   _zz_14963;
  wire       [31:0]   _zz_14964;
  wire       [23:0]   _zz_14965;
  wire       [31:0]   _zz_14966;
  wire       [15:0]   _zz_14967;
  wire       [31:0]   _zz_14968;
  wire       [31:0]   _zz_14969;
  wire       [31:0]   _zz_14970;
  wire       [31:0]   _zz_14971;
  wire       [31:0]   _zz_14972;
  wire       [23:0]   _zz_14973;
  wire       [31:0]   _zz_14974;
  wire       [15:0]   _zz_14975;
  wire       [15:0]   _zz_14976;
  wire       [31:0]   _zz_14977;
  wire       [31:0]   _zz_14978;
  wire       [15:0]   _zz_14979;
  wire       [31:0]   _zz_14980;
  wire       [31:0]   _zz_14981;
  wire       [31:0]   _zz_14982;
  wire       [15:0]   _zz_14983;
  wire       [31:0]   _zz_14984;
  wire       [31:0]   _zz_14985;
  wire       [31:0]   _zz_14986;
  wire       [31:0]   _zz_14987;
  wire       [31:0]   _zz_14988;
  wire       [31:0]   _zz_14989;
  wire       [23:0]   _zz_14990;
  wire       [31:0]   _zz_14991;
  wire       [15:0]   _zz_14992;
  wire       [31:0]   _zz_14993;
  wire       [31:0]   _zz_14994;
  wire       [31:0]   _zz_14995;
  wire       [31:0]   _zz_14996;
  wire       [31:0]   _zz_14997;
  wire       [23:0]   _zz_14998;
  wire       [31:0]   _zz_14999;
  wire       [15:0]   _zz_15000;
  wire       [31:0]   _zz_15001;
  wire       [31:0]   _zz_15002;
  wire       [31:0]   _zz_15003;
  wire       [31:0]   _zz_15004;
  wire       [31:0]   _zz_15005;
  wire       [23:0]   _zz_15006;
  wire       [31:0]   _zz_15007;
  wire       [15:0]   _zz_15008;
  wire       [31:0]   _zz_15009;
  wire       [31:0]   _zz_15010;
  wire       [31:0]   _zz_15011;
  wire       [31:0]   _zz_15012;
  wire       [31:0]   _zz_15013;
  wire       [23:0]   _zz_15014;
  wire       [31:0]   _zz_15015;
  wire       [15:0]   _zz_15016;
  wire       [15:0]   _zz_15017;
  wire       [31:0]   _zz_15018;
  wire       [31:0]   _zz_15019;
  wire       [15:0]   _zz_15020;
  wire       [31:0]   _zz_15021;
  wire       [31:0]   _zz_15022;
  wire       [31:0]   _zz_15023;
  wire       [15:0]   _zz_15024;
  wire       [31:0]   _zz_15025;
  wire       [31:0]   _zz_15026;
  wire       [31:0]   _zz_15027;
  wire       [31:0]   _zz_15028;
  wire       [31:0]   _zz_15029;
  wire       [31:0]   _zz_15030;
  wire       [23:0]   _zz_15031;
  wire       [31:0]   _zz_15032;
  wire       [15:0]   _zz_15033;
  wire       [31:0]   _zz_15034;
  wire       [31:0]   _zz_15035;
  wire       [31:0]   _zz_15036;
  wire       [31:0]   _zz_15037;
  wire       [31:0]   _zz_15038;
  wire       [23:0]   _zz_15039;
  wire       [31:0]   _zz_15040;
  wire       [15:0]   _zz_15041;
  wire       [31:0]   _zz_15042;
  wire       [31:0]   _zz_15043;
  wire       [31:0]   _zz_15044;
  wire       [31:0]   _zz_15045;
  wire       [31:0]   _zz_15046;
  wire       [23:0]   _zz_15047;
  wire       [31:0]   _zz_15048;
  wire       [15:0]   _zz_15049;
  wire       [31:0]   _zz_15050;
  wire       [31:0]   _zz_15051;
  wire       [31:0]   _zz_15052;
  wire       [31:0]   _zz_15053;
  wire       [31:0]   _zz_15054;
  wire       [23:0]   _zz_15055;
  wire       [31:0]   _zz_15056;
  wire       [15:0]   _zz_15057;
  wire       [15:0]   _zz_15058;
  wire       [31:0]   _zz_15059;
  wire       [31:0]   _zz_15060;
  wire       [15:0]   _zz_15061;
  wire       [31:0]   _zz_15062;
  wire       [31:0]   _zz_15063;
  wire       [31:0]   _zz_15064;
  wire       [15:0]   _zz_15065;
  wire       [31:0]   _zz_15066;
  wire       [31:0]   _zz_15067;
  wire       [31:0]   _zz_15068;
  wire       [31:0]   _zz_15069;
  wire       [31:0]   _zz_15070;
  wire       [31:0]   _zz_15071;
  wire       [23:0]   _zz_15072;
  wire       [31:0]   _zz_15073;
  wire       [15:0]   _zz_15074;
  wire       [31:0]   _zz_15075;
  wire       [31:0]   _zz_15076;
  wire       [31:0]   _zz_15077;
  wire       [31:0]   _zz_15078;
  wire       [31:0]   _zz_15079;
  wire       [23:0]   _zz_15080;
  wire       [31:0]   _zz_15081;
  wire       [15:0]   _zz_15082;
  wire       [31:0]   _zz_15083;
  wire       [31:0]   _zz_15084;
  wire       [31:0]   _zz_15085;
  wire       [31:0]   _zz_15086;
  wire       [31:0]   _zz_15087;
  wire       [23:0]   _zz_15088;
  wire       [31:0]   _zz_15089;
  wire       [15:0]   _zz_15090;
  wire       [31:0]   _zz_15091;
  wire       [31:0]   _zz_15092;
  wire       [31:0]   _zz_15093;
  wire       [31:0]   _zz_15094;
  wire       [31:0]   _zz_15095;
  wire       [23:0]   _zz_15096;
  wire       [31:0]   _zz_15097;
  wire       [15:0]   _zz_15098;
  wire       [15:0]   _zz_15099;
  wire       [31:0]   _zz_15100;
  wire       [31:0]   _zz_15101;
  wire       [15:0]   _zz_15102;
  wire       [31:0]   _zz_15103;
  wire       [31:0]   _zz_15104;
  wire       [31:0]   _zz_15105;
  wire       [15:0]   _zz_15106;
  wire       [31:0]   _zz_15107;
  wire       [31:0]   _zz_15108;
  wire       [31:0]   _zz_15109;
  wire       [31:0]   _zz_15110;
  wire       [31:0]   _zz_15111;
  wire       [31:0]   _zz_15112;
  wire       [23:0]   _zz_15113;
  wire       [31:0]   _zz_15114;
  wire       [15:0]   _zz_15115;
  wire       [31:0]   _zz_15116;
  wire       [31:0]   _zz_15117;
  wire       [31:0]   _zz_15118;
  wire       [31:0]   _zz_15119;
  wire       [31:0]   _zz_15120;
  wire       [23:0]   _zz_15121;
  wire       [31:0]   _zz_15122;
  wire       [15:0]   _zz_15123;
  wire       [31:0]   _zz_15124;
  wire       [31:0]   _zz_15125;
  wire       [31:0]   _zz_15126;
  wire       [31:0]   _zz_15127;
  wire       [31:0]   _zz_15128;
  wire       [23:0]   _zz_15129;
  wire       [31:0]   _zz_15130;
  wire       [15:0]   _zz_15131;
  wire       [31:0]   _zz_15132;
  wire       [31:0]   _zz_15133;
  wire       [31:0]   _zz_15134;
  wire       [31:0]   _zz_15135;
  wire       [31:0]   _zz_15136;
  wire       [23:0]   _zz_15137;
  wire       [31:0]   _zz_15138;
  wire       [15:0]   _zz_15139;
  wire       [15:0]   _zz_15140;
  wire       [31:0]   _zz_15141;
  wire       [31:0]   _zz_15142;
  wire       [15:0]   _zz_15143;
  wire       [31:0]   _zz_15144;
  wire       [31:0]   _zz_15145;
  wire       [31:0]   _zz_15146;
  wire       [15:0]   _zz_15147;
  wire       [31:0]   _zz_15148;
  wire       [31:0]   _zz_15149;
  wire       [31:0]   _zz_15150;
  wire       [31:0]   _zz_15151;
  wire       [31:0]   _zz_15152;
  wire       [31:0]   _zz_15153;
  wire       [23:0]   _zz_15154;
  wire       [31:0]   _zz_15155;
  wire       [15:0]   _zz_15156;
  wire       [31:0]   _zz_15157;
  wire       [31:0]   _zz_15158;
  wire       [31:0]   _zz_15159;
  wire       [31:0]   _zz_15160;
  wire       [31:0]   _zz_15161;
  wire       [23:0]   _zz_15162;
  wire       [31:0]   _zz_15163;
  wire       [15:0]   _zz_15164;
  wire       [31:0]   _zz_15165;
  wire       [31:0]   _zz_15166;
  wire       [31:0]   _zz_15167;
  wire       [31:0]   _zz_15168;
  wire       [31:0]   _zz_15169;
  wire       [23:0]   _zz_15170;
  wire       [31:0]   _zz_15171;
  wire       [15:0]   _zz_15172;
  wire       [31:0]   _zz_15173;
  wire       [31:0]   _zz_15174;
  wire       [31:0]   _zz_15175;
  wire       [31:0]   _zz_15176;
  wire       [31:0]   _zz_15177;
  wire       [23:0]   _zz_15178;
  wire       [31:0]   _zz_15179;
  wire       [15:0]   _zz_15180;
  wire       [15:0]   _zz_15181;
  wire       [31:0]   _zz_15182;
  wire       [31:0]   _zz_15183;
  wire       [15:0]   _zz_15184;
  wire       [31:0]   _zz_15185;
  wire       [31:0]   _zz_15186;
  wire       [31:0]   _zz_15187;
  wire       [15:0]   _zz_15188;
  wire       [31:0]   _zz_15189;
  wire       [31:0]   _zz_15190;
  wire       [31:0]   _zz_15191;
  wire       [31:0]   _zz_15192;
  wire       [31:0]   _zz_15193;
  wire       [31:0]   _zz_15194;
  wire       [23:0]   _zz_15195;
  wire       [31:0]   _zz_15196;
  wire       [15:0]   _zz_15197;
  wire       [31:0]   _zz_15198;
  wire       [31:0]   _zz_15199;
  wire       [31:0]   _zz_15200;
  wire       [31:0]   _zz_15201;
  wire       [31:0]   _zz_15202;
  wire       [23:0]   _zz_15203;
  wire       [31:0]   _zz_15204;
  wire       [15:0]   _zz_15205;
  wire       [31:0]   _zz_15206;
  wire       [31:0]   _zz_15207;
  wire       [31:0]   _zz_15208;
  wire       [31:0]   _zz_15209;
  wire       [31:0]   _zz_15210;
  wire       [23:0]   _zz_15211;
  wire       [31:0]   _zz_15212;
  wire       [15:0]   _zz_15213;
  wire       [31:0]   _zz_15214;
  wire       [31:0]   _zz_15215;
  wire       [31:0]   _zz_15216;
  wire       [31:0]   _zz_15217;
  wire       [31:0]   _zz_15218;
  wire       [23:0]   _zz_15219;
  wire       [31:0]   _zz_15220;
  wire       [15:0]   _zz_15221;
  wire       [15:0]   _zz_15222;
  wire       [31:0]   _zz_15223;
  wire       [31:0]   _zz_15224;
  wire       [15:0]   _zz_15225;
  wire       [31:0]   _zz_15226;
  wire       [31:0]   _zz_15227;
  wire       [31:0]   _zz_15228;
  wire       [15:0]   _zz_15229;
  wire       [31:0]   _zz_15230;
  wire       [31:0]   _zz_15231;
  wire       [31:0]   _zz_15232;
  wire       [31:0]   _zz_15233;
  wire       [31:0]   _zz_15234;
  wire       [31:0]   _zz_15235;
  wire       [23:0]   _zz_15236;
  wire       [31:0]   _zz_15237;
  wire       [15:0]   _zz_15238;
  wire       [31:0]   _zz_15239;
  wire       [31:0]   _zz_15240;
  wire       [31:0]   _zz_15241;
  wire       [31:0]   _zz_15242;
  wire       [31:0]   _zz_15243;
  wire       [23:0]   _zz_15244;
  wire       [31:0]   _zz_15245;
  wire       [15:0]   _zz_15246;
  wire       [31:0]   _zz_15247;
  wire       [31:0]   _zz_15248;
  wire       [31:0]   _zz_15249;
  wire       [31:0]   _zz_15250;
  wire       [31:0]   _zz_15251;
  wire       [23:0]   _zz_15252;
  wire       [31:0]   _zz_15253;
  wire       [15:0]   _zz_15254;
  wire       [31:0]   _zz_15255;
  wire       [31:0]   _zz_15256;
  wire       [31:0]   _zz_15257;
  wire       [31:0]   _zz_15258;
  wire       [31:0]   _zz_15259;
  wire       [23:0]   _zz_15260;
  wire       [31:0]   _zz_15261;
  wire       [15:0]   _zz_15262;
  wire       [15:0]   _zz_15263;
  wire       [31:0]   _zz_15264;
  wire       [31:0]   _zz_15265;
  wire       [15:0]   _zz_15266;
  wire       [31:0]   _zz_15267;
  wire       [31:0]   _zz_15268;
  wire       [31:0]   _zz_15269;
  wire       [15:0]   _zz_15270;
  wire       [31:0]   _zz_15271;
  wire       [31:0]   _zz_15272;
  wire       [31:0]   _zz_15273;
  wire       [31:0]   _zz_15274;
  wire       [31:0]   _zz_15275;
  wire       [31:0]   _zz_15276;
  wire       [23:0]   _zz_15277;
  wire       [31:0]   _zz_15278;
  wire       [15:0]   _zz_15279;
  wire       [31:0]   _zz_15280;
  wire       [31:0]   _zz_15281;
  wire       [31:0]   _zz_15282;
  wire       [31:0]   _zz_15283;
  wire       [31:0]   _zz_15284;
  wire       [23:0]   _zz_15285;
  wire       [31:0]   _zz_15286;
  wire       [15:0]   _zz_15287;
  wire       [31:0]   _zz_15288;
  wire       [31:0]   _zz_15289;
  wire       [31:0]   _zz_15290;
  wire       [31:0]   _zz_15291;
  wire       [31:0]   _zz_15292;
  wire       [23:0]   _zz_15293;
  wire       [31:0]   _zz_15294;
  wire       [15:0]   _zz_15295;
  wire       [31:0]   _zz_15296;
  wire       [31:0]   _zz_15297;
  wire       [31:0]   _zz_15298;
  wire       [31:0]   _zz_15299;
  wire       [31:0]   _zz_15300;
  wire       [23:0]   _zz_15301;
  wire       [31:0]   _zz_15302;
  wire       [15:0]   _zz_15303;
  wire       [15:0]   _zz_15304;
  wire       [31:0]   _zz_15305;
  wire       [31:0]   _zz_15306;
  wire       [15:0]   _zz_15307;
  wire       [31:0]   _zz_15308;
  wire       [31:0]   _zz_15309;
  wire       [31:0]   _zz_15310;
  wire       [15:0]   _zz_15311;
  wire       [31:0]   _zz_15312;
  wire       [31:0]   _zz_15313;
  wire       [31:0]   _zz_15314;
  wire       [31:0]   _zz_15315;
  wire       [31:0]   _zz_15316;
  wire       [31:0]   _zz_15317;
  wire       [23:0]   _zz_15318;
  wire       [31:0]   _zz_15319;
  wire       [15:0]   _zz_15320;
  wire       [31:0]   _zz_15321;
  wire       [31:0]   _zz_15322;
  wire       [31:0]   _zz_15323;
  wire       [31:0]   _zz_15324;
  wire       [31:0]   _zz_15325;
  wire       [23:0]   _zz_15326;
  wire       [31:0]   _zz_15327;
  wire       [15:0]   _zz_15328;
  wire       [31:0]   _zz_15329;
  wire       [31:0]   _zz_15330;
  wire       [31:0]   _zz_15331;
  wire       [31:0]   _zz_15332;
  wire       [31:0]   _zz_15333;
  wire       [23:0]   _zz_15334;
  wire       [31:0]   _zz_15335;
  wire       [15:0]   _zz_15336;
  wire       [31:0]   _zz_15337;
  wire       [31:0]   _zz_15338;
  wire       [31:0]   _zz_15339;
  wire       [31:0]   _zz_15340;
  wire       [31:0]   _zz_15341;
  wire       [23:0]   _zz_15342;
  wire       [31:0]   _zz_15343;
  wire       [15:0]   _zz_15344;
  wire       [15:0]   _zz_15345;
  wire       [31:0]   _zz_15346;
  wire       [31:0]   _zz_15347;
  wire       [15:0]   _zz_15348;
  wire       [31:0]   _zz_15349;
  wire       [31:0]   _zz_15350;
  wire       [31:0]   _zz_15351;
  wire       [15:0]   _zz_15352;
  wire       [31:0]   _zz_15353;
  wire       [31:0]   _zz_15354;
  wire       [31:0]   _zz_15355;
  wire       [31:0]   _zz_15356;
  wire       [31:0]   _zz_15357;
  wire       [31:0]   _zz_15358;
  wire       [23:0]   _zz_15359;
  wire       [31:0]   _zz_15360;
  wire       [15:0]   _zz_15361;
  wire       [31:0]   _zz_15362;
  wire       [31:0]   _zz_15363;
  wire       [31:0]   _zz_15364;
  wire       [31:0]   _zz_15365;
  wire       [31:0]   _zz_15366;
  wire       [23:0]   _zz_15367;
  wire       [31:0]   _zz_15368;
  wire       [15:0]   _zz_15369;
  wire       [31:0]   _zz_15370;
  wire       [31:0]   _zz_15371;
  wire       [31:0]   _zz_15372;
  wire       [31:0]   _zz_15373;
  wire       [31:0]   _zz_15374;
  wire       [23:0]   _zz_15375;
  wire       [31:0]   _zz_15376;
  wire       [15:0]   _zz_15377;
  wire       [31:0]   _zz_15378;
  wire       [31:0]   _zz_15379;
  wire       [31:0]   _zz_15380;
  wire       [31:0]   _zz_15381;
  wire       [31:0]   _zz_15382;
  wire       [23:0]   _zz_15383;
  wire       [31:0]   _zz_15384;
  wire       [15:0]   _zz_15385;
  wire       [15:0]   _zz_15386;
  wire       [31:0]   _zz_15387;
  wire       [31:0]   _zz_15388;
  wire       [15:0]   _zz_15389;
  wire       [31:0]   _zz_15390;
  wire       [31:0]   _zz_15391;
  wire       [31:0]   _zz_15392;
  wire       [15:0]   _zz_15393;
  wire       [31:0]   _zz_15394;
  wire       [31:0]   _zz_15395;
  wire       [31:0]   _zz_15396;
  wire       [31:0]   _zz_15397;
  wire       [31:0]   _zz_15398;
  wire       [31:0]   _zz_15399;
  wire       [23:0]   _zz_15400;
  wire       [31:0]   _zz_15401;
  wire       [15:0]   _zz_15402;
  wire       [31:0]   _zz_15403;
  wire       [31:0]   _zz_15404;
  wire       [31:0]   _zz_15405;
  wire       [31:0]   _zz_15406;
  wire       [31:0]   _zz_15407;
  wire       [23:0]   _zz_15408;
  wire       [31:0]   _zz_15409;
  wire       [15:0]   _zz_15410;
  wire       [31:0]   _zz_15411;
  wire       [31:0]   _zz_15412;
  wire       [31:0]   _zz_15413;
  wire       [31:0]   _zz_15414;
  wire       [31:0]   _zz_15415;
  wire       [23:0]   _zz_15416;
  wire       [31:0]   _zz_15417;
  wire       [15:0]   _zz_15418;
  wire       [31:0]   _zz_15419;
  wire       [31:0]   _zz_15420;
  wire       [31:0]   _zz_15421;
  wire       [31:0]   _zz_15422;
  wire       [31:0]   _zz_15423;
  wire       [23:0]   _zz_15424;
  wire       [31:0]   _zz_15425;
  wire       [15:0]   _zz_15426;
  wire       [15:0]   _zz_15427;
  wire       [31:0]   _zz_15428;
  wire       [31:0]   _zz_15429;
  wire       [15:0]   _zz_15430;
  wire       [31:0]   _zz_15431;
  wire       [31:0]   _zz_15432;
  wire       [31:0]   _zz_15433;
  wire       [15:0]   _zz_15434;
  wire       [31:0]   _zz_15435;
  wire       [31:0]   _zz_15436;
  wire       [31:0]   _zz_15437;
  wire       [31:0]   _zz_15438;
  wire       [31:0]   _zz_15439;
  wire       [31:0]   _zz_15440;
  wire       [23:0]   _zz_15441;
  wire       [31:0]   _zz_15442;
  wire       [15:0]   _zz_15443;
  wire       [31:0]   _zz_15444;
  wire       [31:0]   _zz_15445;
  wire       [31:0]   _zz_15446;
  wire       [31:0]   _zz_15447;
  wire       [31:0]   _zz_15448;
  wire       [23:0]   _zz_15449;
  wire       [31:0]   _zz_15450;
  wire       [15:0]   _zz_15451;
  wire       [31:0]   _zz_15452;
  wire       [31:0]   _zz_15453;
  wire       [31:0]   _zz_15454;
  wire       [31:0]   _zz_15455;
  wire       [31:0]   _zz_15456;
  wire       [23:0]   _zz_15457;
  wire       [31:0]   _zz_15458;
  wire       [15:0]   _zz_15459;
  wire       [31:0]   _zz_15460;
  wire       [31:0]   _zz_15461;
  wire       [31:0]   _zz_15462;
  wire       [31:0]   _zz_15463;
  wire       [31:0]   _zz_15464;
  wire       [23:0]   _zz_15465;
  wire       [31:0]   _zz_15466;
  wire       [15:0]   _zz_15467;
  wire       [15:0]   _zz_15468;
  wire       [31:0]   _zz_15469;
  wire       [31:0]   _zz_15470;
  wire       [15:0]   _zz_15471;
  wire       [31:0]   _zz_15472;
  wire       [31:0]   _zz_15473;
  wire       [31:0]   _zz_15474;
  wire       [15:0]   _zz_15475;
  wire       [31:0]   _zz_15476;
  wire       [31:0]   _zz_15477;
  wire       [31:0]   _zz_15478;
  wire       [31:0]   _zz_15479;
  wire       [31:0]   _zz_15480;
  wire       [31:0]   _zz_15481;
  wire       [23:0]   _zz_15482;
  wire       [31:0]   _zz_15483;
  wire       [15:0]   _zz_15484;
  wire       [31:0]   _zz_15485;
  wire       [31:0]   _zz_15486;
  wire       [31:0]   _zz_15487;
  wire       [31:0]   _zz_15488;
  wire       [31:0]   _zz_15489;
  wire       [23:0]   _zz_15490;
  wire       [31:0]   _zz_15491;
  wire       [15:0]   _zz_15492;
  wire       [31:0]   _zz_15493;
  wire       [31:0]   _zz_15494;
  wire       [31:0]   _zz_15495;
  wire       [31:0]   _zz_15496;
  wire       [31:0]   _zz_15497;
  wire       [23:0]   _zz_15498;
  wire       [31:0]   _zz_15499;
  wire       [15:0]   _zz_15500;
  wire       [31:0]   _zz_15501;
  wire       [31:0]   _zz_15502;
  wire       [31:0]   _zz_15503;
  wire       [31:0]   _zz_15504;
  wire       [31:0]   _zz_15505;
  wire       [23:0]   _zz_15506;
  wire       [31:0]   _zz_15507;
  wire       [15:0]   _zz_15508;
  wire       [15:0]   _zz_15509;
  wire       [31:0]   _zz_15510;
  wire       [31:0]   _zz_15511;
  wire       [15:0]   _zz_15512;
  wire       [31:0]   _zz_15513;
  wire       [31:0]   _zz_15514;
  wire       [31:0]   _zz_15515;
  wire       [15:0]   _zz_15516;
  wire       [31:0]   _zz_15517;
  wire       [31:0]   _zz_15518;
  wire       [31:0]   _zz_15519;
  wire       [31:0]   _zz_15520;
  wire       [31:0]   _zz_15521;
  wire       [31:0]   _zz_15522;
  wire       [23:0]   _zz_15523;
  wire       [31:0]   _zz_15524;
  wire       [15:0]   _zz_15525;
  wire       [31:0]   _zz_15526;
  wire       [31:0]   _zz_15527;
  wire       [31:0]   _zz_15528;
  wire       [31:0]   _zz_15529;
  wire       [31:0]   _zz_15530;
  wire       [23:0]   _zz_15531;
  wire       [31:0]   _zz_15532;
  wire       [15:0]   _zz_15533;
  wire       [31:0]   _zz_15534;
  wire       [31:0]   _zz_15535;
  wire       [31:0]   _zz_15536;
  wire       [31:0]   _zz_15537;
  wire       [31:0]   _zz_15538;
  wire       [23:0]   _zz_15539;
  wire       [31:0]   _zz_15540;
  wire       [15:0]   _zz_15541;
  wire       [31:0]   _zz_15542;
  wire       [31:0]   _zz_15543;
  wire       [31:0]   _zz_15544;
  wire       [31:0]   _zz_15545;
  wire       [31:0]   _zz_15546;
  wire       [23:0]   _zz_15547;
  wire       [31:0]   _zz_15548;
  wire       [15:0]   _zz_15549;
  wire       [15:0]   _zz_15550;
  wire       [31:0]   _zz_15551;
  wire       [31:0]   _zz_15552;
  wire       [15:0]   _zz_15553;
  wire       [31:0]   _zz_15554;
  wire       [31:0]   _zz_15555;
  wire       [31:0]   _zz_15556;
  wire       [15:0]   _zz_15557;
  wire       [31:0]   _zz_15558;
  wire       [31:0]   _zz_15559;
  wire       [31:0]   _zz_15560;
  wire       [31:0]   _zz_15561;
  wire       [31:0]   _zz_15562;
  wire       [31:0]   _zz_15563;
  wire       [23:0]   _zz_15564;
  wire       [31:0]   _zz_15565;
  wire       [15:0]   _zz_15566;
  wire       [31:0]   _zz_15567;
  wire       [31:0]   _zz_15568;
  wire       [31:0]   _zz_15569;
  wire       [31:0]   _zz_15570;
  wire       [31:0]   _zz_15571;
  wire       [23:0]   _zz_15572;
  wire       [31:0]   _zz_15573;
  wire       [15:0]   _zz_15574;
  wire       [31:0]   _zz_15575;
  wire       [31:0]   _zz_15576;
  wire       [31:0]   _zz_15577;
  wire       [31:0]   _zz_15578;
  wire       [31:0]   _zz_15579;
  wire       [23:0]   _zz_15580;
  wire       [31:0]   _zz_15581;
  wire       [15:0]   _zz_15582;
  wire       [31:0]   _zz_15583;
  wire       [31:0]   _zz_15584;
  wire       [31:0]   _zz_15585;
  wire       [31:0]   _zz_15586;
  wire       [31:0]   _zz_15587;
  wire       [23:0]   _zz_15588;
  wire       [31:0]   _zz_15589;
  wire       [15:0]   _zz_15590;
  wire       [15:0]   _zz_15591;
  wire       [31:0]   _zz_15592;
  wire       [31:0]   _zz_15593;
  wire       [15:0]   _zz_15594;
  wire       [31:0]   _zz_15595;
  wire       [31:0]   _zz_15596;
  wire       [31:0]   _zz_15597;
  wire       [15:0]   _zz_15598;
  wire       [31:0]   _zz_15599;
  wire       [31:0]   _zz_15600;
  wire       [31:0]   _zz_15601;
  wire       [31:0]   _zz_15602;
  wire       [31:0]   _zz_15603;
  wire       [31:0]   _zz_15604;
  wire       [23:0]   _zz_15605;
  wire       [31:0]   _zz_15606;
  wire       [15:0]   _zz_15607;
  wire       [31:0]   _zz_15608;
  wire       [31:0]   _zz_15609;
  wire       [31:0]   _zz_15610;
  wire       [31:0]   _zz_15611;
  wire       [31:0]   _zz_15612;
  wire       [23:0]   _zz_15613;
  wire       [31:0]   _zz_15614;
  wire       [15:0]   _zz_15615;
  wire       [31:0]   _zz_15616;
  wire       [31:0]   _zz_15617;
  wire       [31:0]   _zz_15618;
  wire       [31:0]   _zz_15619;
  wire       [31:0]   _zz_15620;
  wire       [23:0]   _zz_15621;
  wire       [31:0]   _zz_15622;
  wire       [15:0]   _zz_15623;
  wire       [31:0]   _zz_15624;
  wire       [31:0]   _zz_15625;
  wire       [31:0]   _zz_15626;
  wire       [31:0]   _zz_15627;
  wire       [31:0]   _zz_15628;
  wire       [23:0]   _zz_15629;
  wire       [31:0]   _zz_15630;
  wire       [15:0]   _zz_15631;
  wire       [15:0]   _zz_15632;
  wire       [31:0]   _zz_15633;
  wire       [31:0]   _zz_15634;
  wire       [15:0]   _zz_15635;
  wire       [31:0]   _zz_15636;
  wire       [31:0]   _zz_15637;
  wire       [31:0]   _zz_15638;
  wire       [15:0]   _zz_15639;
  wire       [31:0]   _zz_15640;
  wire       [31:0]   _zz_15641;
  wire       [31:0]   _zz_15642;
  wire       [31:0]   _zz_15643;
  wire       [31:0]   _zz_15644;
  wire       [31:0]   _zz_15645;
  wire       [23:0]   _zz_15646;
  wire       [31:0]   _zz_15647;
  wire       [15:0]   _zz_15648;
  wire       [31:0]   _zz_15649;
  wire       [31:0]   _zz_15650;
  wire       [31:0]   _zz_15651;
  wire       [31:0]   _zz_15652;
  wire       [31:0]   _zz_15653;
  wire       [23:0]   _zz_15654;
  wire       [31:0]   _zz_15655;
  wire       [15:0]   _zz_15656;
  wire       [31:0]   _zz_15657;
  wire       [31:0]   _zz_15658;
  wire       [31:0]   _zz_15659;
  wire       [31:0]   _zz_15660;
  wire       [31:0]   _zz_15661;
  wire       [23:0]   _zz_15662;
  wire       [31:0]   _zz_15663;
  wire       [15:0]   _zz_15664;
  wire       [31:0]   _zz_15665;
  wire       [31:0]   _zz_15666;
  wire       [31:0]   _zz_15667;
  wire       [31:0]   _zz_15668;
  wire       [31:0]   _zz_15669;
  wire       [23:0]   _zz_15670;
  wire       [31:0]   _zz_15671;
  wire       [15:0]   _zz_15672;
  wire       [15:0]   _zz_15673;
  wire       [31:0]   _zz_15674;
  wire       [31:0]   _zz_15675;
  wire       [15:0]   _zz_15676;
  wire       [31:0]   _zz_15677;
  wire       [31:0]   _zz_15678;
  wire       [31:0]   _zz_15679;
  wire       [15:0]   _zz_15680;
  wire       [31:0]   _zz_15681;
  wire       [31:0]   _zz_15682;
  wire       [31:0]   _zz_15683;
  wire       [31:0]   _zz_15684;
  wire       [31:0]   _zz_15685;
  wire       [31:0]   _zz_15686;
  wire       [23:0]   _zz_15687;
  wire       [31:0]   _zz_15688;
  wire       [15:0]   _zz_15689;
  wire       [31:0]   _zz_15690;
  wire       [31:0]   _zz_15691;
  wire       [31:0]   _zz_15692;
  wire       [31:0]   _zz_15693;
  wire       [31:0]   _zz_15694;
  wire       [23:0]   _zz_15695;
  wire       [31:0]   _zz_15696;
  wire       [15:0]   _zz_15697;
  wire       [31:0]   _zz_15698;
  wire       [31:0]   _zz_15699;
  wire       [31:0]   _zz_15700;
  wire       [31:0]   _zz_15701;
  wire       [31:0]   _zz_15702;
  wire       [23:0]   _zz_15703;
  wire       [31:0]   _zz_15704;
  wire       [15:0]   _zz_15705;
  wire       [31:0]   _zz_15706;
  wire       [31:0]   _zz_15707;
  wire       [31:0]   _zz_15708;
  wire       [31:0]   _zz_15709;
  wire       [31:0]   _zz_15710;
  wire       [23:0]   _zz_15711;
  wire       [31:0]   _zz_15712;
  wire       [15:0]   _zz_15713;
  wire       [15:0]   _zz_15714;
  wire       [31:0]   _zz_15715;
  wire       [31:0]   _zz_15716;
  wire       [15:0]   _zz_15717;
  wire       [31:0]   _zz_15718;
  wire       [31:0]   _zz_15719;
  wire       [31:0]   _zz_15720;
  wire       [15:0]   _zz_15721;
  wire       [31:0]   _zz_15722;
  wire       [31:0]   _zz_15723;
  wire       [31:0]   _zz_15724;
  wire       [31:0]   _zz_15725;
  wire       [31:0]   _zz_15726;
  wire       [31:0]   _zz_15727;
  wire       [23:0]   _zz_15728;
  wire       [31:0]   _zz_15729;
  wire       [15:0]   _zz_15730;
  wire       [31:0]   _zz_15731;
  wire       [31:0]   _zz_15732;
  wire       [31:0]   _zz_15733;
  wire       [31:0]   _zz_15734;
  wire       [31:0]   _zz_15735;
  wire       [23:0]   _zz_15736;
  wire       [31:0]   _zz_15737;
  wire       [15:0]   _zz_15738;
  wire       [31:0]   _zz_15739;
  wire       [31:0]   _zz_15740;
  wire       [31:0]   _zz_15741;
  wire       [31:0]   _zz_15742;
  wire       [31:0]   _zz_15743;
  wire       [23:0]   _zz_15744;
  wire       [31:0]   _zz_15745;
  wire       [15:0]   _zz_15746;
  wire       [31:0]   _zz_15747;
  wire       [31:0]   _zz_15748;
  wire       [31:0]   _zz_15749;
  wire       [31:0]   _zz_15750;
  wire       [31:0]   _zz_15751;
  wire       [23:0]   _zz_15752;
  wire       [31:0]   _zz_15753;
  wire       [15:0]   _zz_15754;
  wire       [15:0]   _zz_15755;
  wire       [31:0]   _zz_15756;
  wire       [31:0]   _zz_15757;
  wire       [15:0]   _zz_15758;
  wire       [31:0]   _zz_15759;
  wire       [31:0]   _zz_15760;
  wire       [31:0]   _zz_15761;
  wire       [15:0]   _zz_15762;
  wire       [31:0]   _zz_15763;
  wire       [31:0]   _zz_15764;
  wire       [31:0]   _zz_15765;
  wire       [31:0]   _zz_15766;
  wire       [31:0]   _zz_15767;
  wire       [31:0]   _zz_15768;
  wire       [23:0]   _zz_15769;
  wire       [31:0]   _zz_15770;
  wire       [15:0]   _zz_15771;
  wire       [31:0]   _zz_15772;
  wire       [31:0]   _zz_15773;
  wire       [31:0]   _zz_15774;
  wire       [31:0]   _zz_15775;
  wire       [31:0]   _zz_15776;
  wire       [23:0]   _zz_15777;
  wire       [31:0]   _zz_15778;
  wire       [15:0]   _zz_15779;
  wire       [31:0]   _zz_15780;
  wire       [31:0]   _zz_15781;
  wire       [31:0]   _zz_15782;
  wire       [31:0]   _zz_15783;
  wire       [31:0]   _zz_15784;
  wire       [23:0]   _zz_15785;
  wire       [31:0]   _zz_15786;
  wire       [15:0]   _zz_15787;
  wire       [31:0]   _zz_15788;
  wire       [31:0]   _zz_15789;
  wire       [31:0]   _zz_15790;
  wire       [31:0]   _zz_15791;
  wire       [31:0]   _zz_15792;
  wire       [23:0]   _zz_15793;
  wire       [31:0]   _zz_15794;
  wire       [15:0]   _zz_15795;
  wire       [15:0]   _zz_15796;
  wire       [31:0]   _zz_15797;
  wire       [31:0]   _zz_15798;
  wire       [15:0]   _zz_15799;
  wire       [31:0]   _zz_15800;
  wire       [31:0]   _zz_15801;
  wire       [31:0]   _zz_15802;
  wire       [15:0]   _zz_15803;
  wire       [31:0]   _zz_15804;
  wire       [31:0]   _zz_15805;
  wire       [31:0]   _zz_15806;
  wire       [31:0]   _zz_15807;
  wire       [31:0]   _zz_15808;
  wire       [31:0]   _zz_15809;
  wire       [23:0]   _zz_15810;
  wire       [31:0]   _zz_15811;
  wire       [15:0]   _zz_15812;
  wire       [31:0]   _zz_15813;
  wire       [31:0]   _zz_15814;
  wire       [31:0]   _zz_15815;
  wire       [31:0]   _zz_15816;
  wire       [31:0]   _zz_15817;
  wire       [23:0]   _zz_15818;
  wire       [31:0]   _zz_15819;
  wire       [15:0]   _zz_15820;
  wire       [31:0]   _zz_15821;
  wire       [31:0]   _zz_15822;
  wire       [31:0]   _zz_15823;
  wire       [31:0]   _zz_15824;
  wire       [31:0]   _zz_15825;
  wire       [23:0]   _zz_15826;
  wire       [31:0]   _zz_15827;
  wire       [15:0]   _zz_15828;
  wire       [31:0]   _zz_15829;
  wire       [31:0]   _zz_15830;
  wire       [31:0]   _zz_15831;
  wire       [31:0]   _zz_15832;
  wire       [31:0]   _zz_15833;
  wire       [23:0]   _zz_15834;
  wire       [31:0]   _zz_15835;
  wire       [15:0]   _zz_15836;
  wire       [15:0]   _zz_15837;
  wire       [31:0]   _zz_15838;
  wire       [31:0]   _zz_15839;
  wire       [15:0]   _zz_15840;
  wire       [31:0]   _zz_15841;
  wire       [31:0]   _zz_15842;
  wire       [31:0]   _zz_15843;
  wire       [15:0]   _zz_15844;
  wire       [31:0]   _zz_15845;
  wire       [31:0]   _zz_15846;
  wire       [31:0]   _zz_15847;
  wire       [31:0]   _zz_15848;
  wire       [31:0]   _zz_15849;
  wire       [31:0]   _zz_15850;
  wire       [23:0]   _zz_15851;
  wire       [31:0]   _zz_15852;
  wire       [15:0]   _zz_15853;
  wire       [31:0]   _zz_15854;
  wire       [31:0]   _zz_15855;
  wire       [31:0]   _zz_15856;
  wire       [31:0]   _zz_15857;
  wire       [31:0]   _zz_15858;
  wire       [23:0]   _zz_15859;
  wire       [31:0]   _zz_15860;
  wire       [15:0]   _zz_15861;
  wire       [31:0]   _zz_15862;
  wire       [31:0]   _zz_15863;
  wire       [31:0]   _zz_15864;
  wire       [31:0]   _zz_15865;
  wire       [31:0]   _zz_15866;
  wire       [23:0]   _zz_15867;
  wire       [31:0]   _zz_15868;
  wire       [15:0]   _zz_15869;
  wire       [31:0]   _zz_15870;
  wire       [31:0]   _zz_15871;
  wire       [31:0]   _zz_15872;
  wire       [31:0]   _zz_15873;
  wire       [31:0]   _zz_15874;
  wire       [23:0]   _zz_15875;
  wire       [31:0]   _zz_15876;
  wire       [15:0]   _zz_15877;
  wire       [15:0]   _zz_15878;
  wire       [31:0]   _zz_15879;
  wire       [31:0]   _zz_15880;
  wire       [15:0]   _zz_15881;
  wire       [31:0]   _zz_15882;
  wire       [31:0]   _zz_15883;
  wire       [31:0]   _zz_15884;
  wire       [15:0]   _zz_15885;
  wire       [31:0]   _zz_15886;
  wire       [31:0]   _zz_15887;
  wire       [31:0]   _zz_15888;
  wire       [31:0]   _zz_15889;
  wire       [31:0]   _zz_15890;
  wire       [31:0]   _zz_15891;
  wire       [23:0]   _zz_15892;
  wire       [31:0]   _zz_15893;
  wire       [15:0]   _zz_15894;
  wire       [31:0]   _zz_15895;
  wire       [31:0]   _zz_15896;
  wire       [31:0]   _zz_15897;
  wire       [31:0]   _zz_15898;
  wire       [31:0]   _zz_15899;
  wire       [23:0]   _zz_15900;
  wire       [31:0]   _zz_15901;
  wire       [15:0]   _zz_15902;
  wire       [31:0]   _zz_15903;
  wire       [31:0]   _zz_15904;
  wire       [31:0]   _zz_15905;
  wire       [31:0]   _zz_15906;
  wire       [31:0]   _zz_15907;
  wire       [23:0]   _zz_15908;
  wire       [31:0]   _zz_15909;
  wire       [15:0]   _zz_15910;
  wire       [31:0]   _zz_15911;
  wire       [31:0]   _zz_15912;
  wire       [31:0]   _zz_15913;
  wire       [31:0]   _zz_15914;
  wire       [31:0]   _zz_15915;
  wire       [23:0]   _zz_15916;
  wire       [31:0]   _zz_15917;
  wire       [15:0]   _zz_15918;
  wire       [15:0]   _zz_15919;
  wire       [31:0]   _zz_15920;
  wire       [31:0]   _zz_15921;
  wire       [15:0]   _zz_15922;
  wire       [31:0]   _zz_15923;
  wire       [31:0]   _zz_15924;
  wire       [31:0]   _zz_15925;
  wire       [15:0]   _zz_15926;
  wire       [31:0]   _zz_15927;
  wire       [31:0]   _zz_15928;
  wire       [31:0]   _zz_15929;
  wire       [31:0]   _zz_15930;
  wire       [31:0]   _zz_15931;
  wire       [31:0]   _zz_15932;
  wire       [23:0]   _zz_15933;
  wire       [31:0]   _zz_15934;
  wire       [15:0]   _zz_15935;
  wire       [31:0]   _zz_15936;
  wire       [31:0]   _zz_15937;
  wire       [31:0]   _zz_15938;
  wire       [31:0]   _zz_15939;
  wire       [31:0]   _zz_15940;
  wire       [23:0]   _zz_15941;
  wire       [31:0]   _zz_15942;
  wire       [15:0]   _zz_15943;
  wire       [31:0]   _zz_15944;
  wire       [31:0]   _zz_15945;
  wire       [31:0]   _zz_15946;
  wire       [31:0]   _zz_15947;
  wire       [31:0]   _zz_15948;
  wire       [23:0]   _zz_15949;
  wire       [31:0]   _zz_15950;
  wire       [15:0]   _zz_15951;
  wire       [31:0]   _zz_15952;
  wire       [31:0]   _zz_15953;
  wire       [31:0]   _zz_15954;
  wire       [31:0]   _zz_15955;
  wire       [31:0]   _zz_15956;
  wire       [23:0]   _zz_15957;
  wire       [31:0]   _zz_15958;
  wire       [15:0]   _zz_15959;
  wire       [15:0]   _zz_15960;
  wire       [31:0]   _zz_15961;
  wire       [31:0]   _zz_15962;
  wire       [15:0]   _zz_15963;
  wire       [31:0]   _zz_15964;
  wire       [31:0]   _zz_15965;
  wire       [31:0]   _zz_15966;
  wire       [15:0]   _zz_15967;
  wire       [31:0]   _zz_15968;
  wire       [31:0]   _zz_15969;
  wire       [31:0]   _zz_15970;
  wire       [31:0]   _zz_15971;
  wire       [31:0]   _zz_15972;
  wire       [31:0]   _zz_15973;
  wire       [23:0]   _zz_15974;
  wire       [31:0]   _zz_15975;
  wire       [15:0]   _zz_15976;
  wire       [31:0]   _zz_15977;
  wire       [31:0]   _zz_15978;
  wire       [31:0]   _zz_15979;
  wire       [31:0]   _zz_15980;
  wire       [31:0]   _zz_15981;
  wire       [23:0]   _zz_15982;
  wire       [31:0]   _zz_15983;
  wire       [15:0]   _zz_15984;
  wire       [31:0]   _zz_15985;
  wire       [31:0]   _zz_15986;
  wire       [31:0]   _zz_15987;
  wire       [31:0]   _zz_15988;
  wire       [31:0]   _zz_15989;
  wire       [23:0]   _zz_15990;
  wire       [31:0]   _zz_15991;
  wire       [15:0]   _zz_15992;
  wire       [31:0]   _zz_15993;
  wire       [31:0]   _zz_15994;
  wire       [31:0]   _zz_15995;
  wire       [31:0]   _zz_15996;
  wire       [31:0]   _zz_15997;
  wire       [23:0]   _zz_15998;
  wire       [31:0]   _zz_15999;
  wire       [15:0]   _zz_16000;
  wire       [15:0]   _zz_16001;
  wire       [31:0]   _zz_16002;
  wire       [31:0]   _zz_16003;
  wire       [15:0]   _zz_16004;
  wire       [31:0]   _zz_16005;
  wire       [31:0]   _zz_16006;
  wire       [31:0]   _zz_16007;
  wire       [15:0]   _zz_16008;
  wire       [31:0]   _zz_16009;
  wire       [31:0]   _zz_16010;
  wire       [31:0]   _zz_16011;
  wire       [31:0]   _zz_16012;
  wire       [31:0]   _zz_16013;
  wire       [31:0]   _zz_16014;
  wire       [23:0]   _zz_16015;
  wire       [31:0]   _zz_16016;
  wire       [15:0]   _zz_16017;
  wire       [31:0]   _zz_16018;
  wire       [31:0]   _zz_16019;
  wire       [31:0]   _zz_16020;
  wire       [31:0]   _zz_16021;
  wire       [31:0]   _zz_16022;
  wire       [23:0]   _zz_16023;
  wire       [31:0]   _zz_16024;
  wire       [15:0]   _zz_16025;
  wire       [31:0]   _zz_16026;
  wire       [31:0]   _zz_16027;
  wire       [31:0]   _zz_16028;
  wire       [31:0]   _zz_16029;
  wire       [31:0]   _zz_16030;
  wire       [23:0]   _zz_16031;
  wire       [31:0]   _zz_16032;
  wire       [15:0]   _zz_16033;
  wire       [31:0]   _zz_16034;
  wire       [31:0]   _zz_16035;
  wire       [31:0]   _zz_16036;
  wire       [31:0]   _zz_16037;
  wire       [31:0]   _zz_16038;
  wire       [23:0]   _zz_16039;
  wire       [31:0]   _zz_16040;
  wire       [15:0]   _zz_16041;
  wire       [15:0]   _zz_16042;
  wire       [31:0]   _zz_16043;
  wire       [31:0]   _zz_16044;
  wire       [15:0]   _zz_16045;
  wire       [31:0]   _zz_16046;
  wire       [31:0]   _zz_16047;
  wire       [31:0]   _zz_16048;
  wire       [15:0]   _zz_16049;
  wire       [31:0]   _zz_16050;
  wire       [31:0]   _zz_16051;
  wire       [31:0]   _zz_16052;
  wire       [31:0]   _zz_16053;
  wire       [31:0]   _zz_16054;
  wire       [31:0]   _zz_16055;
  wire       [23:0]   _zz_16056;
  wire       [31:0]   _zz_16057;
  wire       [15:0]   _zz_16058;
  wire       [31:0]   _zz_16059;
  wire       [31:0]   _zz_16060;
  wire       [31:0]   _zz_16061;
  wire       [31:0]   _zz_16062;
  wire       [31:0]   _zz_16063;
  wire       [23:0]   _zz_16064;
  wire       [31:0]   _zz_16065;
  wire       [15:0]   _zz_16066;
  wire       [31:0]   _zz_16067;
  wire       [31:0]   _zz_16068;
  wire       [31:0]   _zz_16069;
  wire       [31:0]   _zz_16070;
  wire       [31:0]   _zz_16071;
  wire       [23:0]   _zz_16072;
  wire       [31:0]   _zz_16073;
  wire       [15:0]   _zz_16074;
  wire       [31:0]   _zz_16075;
  wire       [31:0]   _zz_16076;
  wire       [31:0]   _zz_16077;
  wire       [31:0]   _zz_16078;
  wire       [31:0]   _zz_16079;
  wire       [23:0]   _zz_16080;
  wire       [31:0]   _zz_16081;
  wire       [15:0]   _zz_16082;
  wire       [15:0]   _zz_16083;
  wire       [31:0]   _zz_16084;
  wire       [31:0]   _zz_16085;
  wire       [15:0]   _zz_16086;
  wire       [31:0]   _zz_16087;
  wire       [31:0]   _zz_16088;
  wire       [31:0]   _zz_16089;
  wire       [15:0]   _zz_16090;
  wire       [31:0]   _zz_16091;
  wire       [31:0]   _zz_16092;
  wire       [31:0]   _zz_16093;
  wire       [31:0]   _zz_16094;
  wire       [31:0]   _zz_16095;
  wire       [31:0]   _zz_16096;
  wire       [23:0]   _zz_16097;
  wire       [31:0]   _zz_16098;
  wire       [15:0]   _zz_16099;
  wire       [31:0]   _zz_16100;
  wire       [31:0]   _zz_16101;
  wire       [31:0]   _zz_16102;
  wire       [31:0]   _zz_16103;
  wire       [31:0]   _zz_16104;
  wire       [23:0]   _zz_16105;
  wire       [31:0]   _zz_16106;
  wire       [15:0]   _zz_16107;
  wire       [31:0]   _zz_16108;
  wire       [31:0]   _zz_16109;
  wire       [31:0]   _zz_16110;
  wire       [31:0]   _zz_16111;
  wire       [31:0]   _zz_16112;
  wire       [23:0]   _zz_16113;
  wire       [31:0]   _zz_16114;
  wire       [15:0]   _zz_16115;
  wire       [31:0]   _zz_16116;
  wire       [31:0]   _zz_16117;
  wire       [31:0]   _zz_16118;
  wire       [31:0]   _zz_16119;
  wire       [31:0]   _zz_16120;
  wire       [23:0]   _zz_16121;
  wire       [31:0]   _zz_16122;
  wire       [15:0]   _zz_16123;
  wire       [15:0]   _zz_16124;
  wire       [31:0]   _zz_16125;
  wire       [31:0]   _zz_16126;
  wire       [15:0]   _zz_16127;
  wire       [31:0]   _zz_16128;
  wire       [31:0]   _zz_16129;
  wire       [31:0]   _zz_16130;
  wire       [15:0]   _zz_16131;
  wire       [31:0]   _zz_16132;
  wire       [31:0]   _zz_16133;
  wire       [31:0]   _zz_16134;
  wire       [31:0]   _zz_16135;
  wire       [31:0]   _zz_16136;
  wire       [31:0]   _zz_16137;
  wire       [23:0]   _zz_16138;
  wire       [31:0]   _zz_16139;
  wire       [15:0]   _zz_16140;
  wire       [31:0]   _zz_16141;
  wire       [31:0]   _zz_16142;
  wire       [31:0]   _zz_16143;
  wire       [31:0]   _zz_16144;
  wire       [31:0]   _zz_16145;
  wire       [23:0]   _zz_16146;
  wire       [31:0]   _zz_16147;
  wire       [15:0]   _zz_16148;
  wire       [31:0]   _zz_16149;
  wire       [31:0]   _zz_16150;
  wire       [31:0]   _zz_16151;
  wire       [31:0]   _zz_16152;
  wire       [31:0]   _zz_16153;
  wire       [23:0]   _zz_16154;
  wire       [31:0]   _zz_16155;
  wire       [15:0]   _zz_16156;
  wire       [31:0]   _zz_16157;
  wire       [31:0]   _zz_16158;
  wire       [31:0]   _zz_16159;
  wire       [31:0]   _zz_16160;
  wire       [31:0]   _zz_16161;
  wire       [23:0]   _zz_16162;
  wire       [31:0]   _zz_16163;
  wire       [15:0]   _zz_16164;
  wire       [15:0]   _zz_16165;
  wire       [31:0]   _zz_16166;
  wire       [31:0]   _zz_16167;
  wire       [15:0]   _zz_16168;
  wire       [31:0]   _zz_16169;
  wire       [31:0]   _zz_16170;
  wire       [31:0]   _zz_16171;
  wire       [15:0]   _zz_16172;
  wire       [31:0]   _zz_16173;
  wire       [31:0]   _zz_16174;
  wire       [31:0]   _zz_16175;
  wire       [31:0]   _zz_16176;
  wire       [31:0]   _zz_16177;
  wire       [31:0]   _zz_16178;
  wire       [23:0]   _zz_16179;
  wire       [31:0]   _zz_16180;
  wire       [15:0]   _zz_16181;
  wire       [31:0]   _zz_16182;
  wire       [31:0]   _zz_16183;
  wire       [31:0]   _zz_16184;
  wire       [31:0]   _zz_16185;
  wire       [31:0]   _zz_16186;
  wire       [23:0]   _zz_16187;
  wire       [31:0]   _zz_16188;
  wire       [15:0]   _zz_16189;
  wire       [31:0]   _zz_16190;
  wire       [31:0]   _zz_16191;
  wire       [31:0]   _zz_16192;
  wire       [31:0]   _zz_16193;
  wire       [31:0]   _zz_16194;
  wire       [23:0]   _zz_16195;
  wire       [31:0]   _zz_16196;
  wire       [15:0]   _zz_16197;
  wire       [31:0]   _zz_16198;
  wire       [31:0]   _zz_16199;
  wire       [31:0]   _zz_16200;
  wire       [31:0]   _zz_16201;
  wire       [31:0]   _zz_16202;
  wire       [23:0]   _zz_16203;
  wire       [31:0]   _zz_16204;
  wire       [15:0]   _zz_16205;
  wire       [15:0]   _zz_16206;
  wire       [31:0]   _zz_16207;
  wire       [31:0]   _zz_16208;
  wire       [15:0]   _zz_16209;
  wire       [31:0]   _zz_16210;
  wire       [31:0]   _zz_16211;
  wire       [31:0]   _zz_16212;
  wire       [15:0]   _zz_16213;
  wire       [31:0]   _zz_16214;
  wire       [31:0]   _zz_16215;
  wire       [31:0]   _zz_16216;
  wire       [31:0]   _zz_16217;
  wire       [31:0]   _zz_16218;
  wire       [31:0]   _zz_16219;
  wire       [23:0]   _zz_16220;
  wire       [31:0]   _zz_16221;
  wire       [15:0]   _zz_16222;
  wire       [31:0]   _zz_16223;
  wire       [31:0]   _zz_16224;
  wire       [31:0]   _zz_16225;
  wire       [31:0]   _zz_16226;
  wire       [31:0]   _zz_16227;
  wire       [23:0]   _zz_16228;
  wire       [31:0]   _zz_16229;
  wire       [15:0]   _zz_16230;
  wire       [31:0]   _zz_16231;
  wire       [31:0]   _zz_16232;
  wire       [31:0]   _zz_16233;
  wire       [31:0]   _zz_16234;
  wire       [31:0]   _zz_16235;
  wire       [23:0]   _zz_16236;
  wire       [31:0]   _zz_16237;
  wire       [15:0]   _zz_16238;
  wire       [31:0]   _zz_16239;
  wire       [31:0]   _zz_16240;
  wire       [31:0]   _zz_16241;
  wire       [31:0]   _zz_16242;
  wire       [31:0]   _zz_16243;
  wire       [23:0]   _zz_16244;
  wire       [31:0]   _zz_16245;
  wire       [15:0]   _zz_16246;
  wire       [15:0]   _zz_16247;
  wire       [31:0]   _zz_16248;
  wire       [31:0]   _zz_16249;
  wire       [15:0]   _zz_16250;
  wire       [31:0]   _zz_16251;
  wire       [31:0]   _zz_16252;
  wire       [31:0]   _zz_16253;
  wire       [15:0]   _zz_16254;
  wire       [31:0]   _zz_16255;
  wire       [31:0]   _zz_16256;
  wire       [31:0]   _zz_16257;
  wire       [31:0]   _zz_16258;
  wire       [31:0]   _zz_16259;
  wire       [31:0]   _zz_16260;
  wire       [23:0]   _zz_16261;
  wire       [31:0]   _zz_16262;
  wire       [15:0]   _zz_16263;
  wire       [31:0]   _zz_16264;
  wire       [31:0]   _zz_16265;
  wire       [31:0]   _zz_16266;
  wire       [31:0]   _zz_16267;
  wire       [31:0]   _zz_16268;
  wire       [23:0]   _zz_16269;
  wire       [31:0]   _zz_16270;
  wire       [15:0]   _zz_16271;
  wire       [31:0]   _zz_16272;
  wire       [31:0]   _zz_16273;
  wire       [31:0]   _zz_16274;
  wire       [31:0]   _zz_16275;
  wire       [31:0]   _zz_16276;
  wire       [23:0]   _zz_16277;
  wire       [31:0]   _zz_16278;
  wire       [15:0]   _zz_16279;
  wire       [31:0]   _zz_16280;
  wire       [31:0]   _zz_16281;
  wire       [31:0]   _zz_16282;
  wire       [31:0]   _zz_16283;
  wire       [31:0]   _zz_16284;
  wire       [23:0]   _zz_16285;
  wire       [31:0]   _zz_16286;
  wire       [15:0]   _zz_16287;
  wire       [15:0]   _zz_16288;
  wire       [31:0]   _zz_16289;
  wire       [31:0]   _zz_16290;
  wire       [15:0]   _zz_16291;
  wire       [31:0]   _zz_16292;
  wire       [31:0]   _zz_16293;
  wire       [31:0]   _zz_16294;
  wire       [15:0]   _zz_16295;
  wire       [31:0]   _zz_16296;
  wire       [31:0]   _zz_16297;
  wire       [31:0]   _zz_16298;
  wire       [31:0]   _zz_16299;
  wire       [31:0]   _zz_16300;
  wire       [31:0]   _zz_16301;
  wire       [23:0]   _zz_16302;
  wire       [31:0]   _zz_16303;
  wire       [15:0]   _zz_16304;
  wire       [31:0]   _zz_16305;
  wire       [31:0]   _zz_16306;
  wire       [31:0]   _zz_16307;
  wire       [31:0]   _zz_16308;
  wire       [31:0]   _zz_16309;
  wire       [23:0]   _zz_16310;
  wire       [31:0]   _zz_16311;
  wire       [15:0]   _zz_16312;
  wire       [31:0]   _zz_16313;
  wire       [31:0]   _zz_16314;
  wire       [31:0]   _zz_16315;
  wire       [31:0]   _zz_16316;
  wire       [31:0]   _zz_16317;
  wire       [23:0]   _zz_16318;
  wire       [31:0]   _zz_16319;
  wire       [15:0]   _zz_16320;
  wire       [31:0]   _zz_16321;
  wire       [31:0]   _zz_16322;
  wire       [31:0]   _zz_16323;
  wire       [31:0]   _zz_16324;
  wire       [31:0]   _zz_16325;
  wire       [23:0]   _zz_16326;
  wire       [31:0]   _zz_16327;
  wire       [15:0]   _zz_16328;
  wire       [15:0]   _zz_16329;
  wire       [31:0]   _zz_16330;
  wire       [31:0]   _zz_16331;
  wire       [15:0]   _zz_16332;
  wire       [31:0]   _zz_16333;
  wire       [31:0]   _zz_16334;
  wire       [31:0]   _zz_16335;
  wire       [15:0]   _zz_16336;
  wire       [31:0]   _zz_16337;
  wire       [31:0]   _zz_16338;
  wire       [31:0]   _zz_16339;
  wire       [31:0]   _zz_16340;
  wire       [31:0]   _zz_16341;
  wire       [31:0]   _zz_16342;
  wire       [23:0]   _zz_16343;
  wire       [31:0]   _zz_16344;
  wire       [15:0]   _zz_16345;
  wire       [31:0]   _zz_16346;
  wire       [31:0]   _zz_16347;
  wire       [31:0]   _zz_16348;
  wire       [31:0]   _zz_16349;
  wire       [31:0]   _zz_16350;
  wire       [23:0]   _zz_16351;
  wire       [31:0]   _zz_16352;
  wire       [15:0]   _zz_16353;
  wire       [31:0]   _zz_16354;
  wire       [31:0]   _zz_16355;
  wire       [31:0]   _zz_16356;
  wire       [31:0]   _zz_16357;
  wire       [31:0]   _zz_16358;
  wire       [23:0]   _zz_16359;
  wire       [31:0]   _zz_16360;
  wire       [15:0]   _zz_16361;
  wire       [31:0]   _zz_16362;
  wire       [31:0]   _zz_16363;
  wire       [31:0]   _zz_16364;
  wire       [31:0]   _zz_16365;
  wire       [31:0]   _zz_16366;
  wire       [23:0]   _zz_16367;
  wire       [31:0]   _zz_16368;
  wire       [15:0]   _zz_16369;
  wire       [15:0]   _zz_16370;
  wire       [31:0]   _zz_16371;
  wire       [31:0]   _zz_16372;
  wire       [15:0]   _zz_16373;
  wire       [31:0]   _zz_16374;
  wire       [31:0]   _zz_16375;
  wire       [31:0]   _zz_16376;
  wire       [15:0]   _zz_16377;
  wire       [31:0]   _zz_16378;
  wire       [31:0]   _zz_16379;
  wire       [31:0]   _zz_16380;
  wire       [31:0]   _zz_16381;
  wire       [31:0]   _zz_16382;
  wire       [31:0]   _zz_16383;
  wire       [23:0]   _zz_16384;
  wire       [31:0]   _zz_16385;
  wire       [15:0]   _zz_16386;
  wire       [31:0]   _zz_16387;
  wire       [31:0]   _zz_16388;
  wire       [31:0]   _zz_16389;
  wire       [31:0]   _zz_16390;
  wire       [31:0]   _zz_16391;
  wire       [23:0]   _zz_16392;
  wire       [31:0]   _zz_16393;
  wire       [15:0]   _zz_16394;
  wire       [31:0]   _zz_16395;
  wire       [31:0]   _zz_16396;
  wire       [31:0]   _zz_16397;
  wire       [31:0]   _zz_16398;
  wire       [31:0]   _zz_16399;
  wire       [23:0]   _zz_16400;
  wire       [31:0]   _zz_16401;
  wire       [15:0]   _zz_16402;
  wire       [31:0]   _zz_16403;
  wire       [31:0]   _zz_16404;
  wire       [31:0]   _zz_16405;
  wire       [31:0]   _zz_16406;
  wire       [31:0]   _zz_16407;
  wire       [23:0]   _zz_16408;
  wire       [31:0]   _zz_16409;
  wire       [15:0]   _zz_16410;
  wire       [15:0]   _zz_16411;
  wire       [31:0]   _zz_16412;
  wire       [31:0]   _zz_16413;
  wire       [15:0]   _zz_16414;
  wire       [31:0]   _zz_16415;
  wire       [31:0]   _zz_16416;
  wire       [31:0]   _zz_16417;
  wire       [15:0]   _zz_16418;
  wire       [31:0]   _zz_16419;
  wire       [31:0]   _zz_16420;
  wire       [31:0]   _zz_16421;
  wire       [31:0]   _zz_16422;
  wire       [31:0]   _zz_16423;
  wire       [31:0]   _zz_16424;
  wire       [23:0]   _zz_16425;
  wire       [31:0]   _zz_16426;
  wire       [15:0]   _zz_16427;
  wire       [31:0]   _zz_16428;
  wire       [31:0]   _zz_16429;
  wire       [31:0]   _zz_16430;
  wire       [31:0]   _zz_16431;
  wire       [31:0]   _zz_16432;
  wire       [23:0]   _zz_16433;
  wire       [31:0]   _zz_16434;
  wire       [15:0]   _zz_16435;
  wire       [31:0]   _zz_16436;
  wire       [31:0]   _zz_16437;
  wire       [31:0]   _zz_16438;
  wire       [31:0]   _zz_16439;
  wire       [31:0]   _zz_16440;
  wire       [23:0]   _zz_16441;
  wire       [31:0]   _zz_16442;
  wire       [15:0]   _zz_16443;
  wire       [31:0]   _zz_16444;
  wire       [31:0]   _zz_16445;
  wire       [31:0]   _zz_16446;
  wire       [31:0]   _zz_16447;
  wire       [31:0]   _zz_16448;
  wire       [23:0]   _zz_16449;
  wire       [31:0]   _zz_16450;
  wire       [15:0]   _zz_16451;
  wire       [15:0]   _zz_16452;
  wire       [31:0]   _zz_16453;
  wire       [31:0]   _zz_16454;
  wire       [15:0]   _zz_16455;
  wire       [31:0]   _zz_16456;
  wire       [31:0]   _zz_16457;
  wire       [31:0]   _zz_16458;
  wire       [15:0]   _zz_16459;
  wire       [31:0]   _zz_16460;
  wire       [31:0]   _zz_16461;
  wire       [31:0]   _zz_16462;
  wire       [31:0]   _zz_16463;
  wire       [31:0]   _zz_16464;
  wire       [31:0]   _zz_16465;
  wire       [23:0]   _zz_16466;
  wire       [31:0]   _zz_16467;
  wire       [15:0]   _zz_16468;
  wire       [31:0]   _zz_16469;
  wire       [31:0]   _zz_16470;
  wire       [31:0]   _zz_16471;
  wire       [31:0]   _zz_16472;
  wire       [31:0]   _zz_16473;
  wire       [23:0]   _zz_16474;
  wire       [31:0]   _zz_16475;
  wire       [15:0]   _zz_16476;
  wire       [31:0]   _zz_16477;
  wire       [31:0]   _zz_16478;
  wire       [31:0]   _zz_16479;
  wire       [31:0]   _zz_16480;
  wire       [31:0]   _zz_16481;
  wire       [23:0]   _zz_16482;
  wire       [31:0]   _zz_16483;
  wire       [15:0]   _zz_16484;
  wire       [31:0]   _zz_16485;
  wire       [31:0]   _zz_16486;
  wire       [31:0]   _zz_16487;
  wire       [31:0]   _zz_16488;
  wire       [31:0]   _zz_16489;
  wire       [23:0]   _zz_16490;
  wire       [31:0]   _zz_16491;
  wire       [15:0]   _zz_16492;
  wire       [15:0]   _zz_16493;
  wire       [31:0]   _zz_16494;
  wire       [31:0]   _zz_16495;
  wire       [15:0]   _zz_16496;
  wire       [31:0]   _zz_16497;
  wire       [31:0]   _zz_16498;
  wire       [31:0]   _zz_16499;
  wire       [15:0]   _zz_16500;
  wire       [31:0]   _zz_16501;
  wire       [31:0]   _zz_16502;
  wire       [31:0]   _zz_16503;
  wire       [31:0]   _zz_16504;
  wire       [31:0]   _zz_16505;
  wire       [31:0]   _zz_16506;
  wire       [23:0]   _zz_16507;
  wire       [31:0]   _zz_16508;
  wire       [15:0]   _zz_16509;
  wire       [31:0]   _zz_16510;
  wire       [31:0]   _zz_16511;
  wire       [31:0]   _zz_16512;
  wire       [31:0]   _zz_16513;
  wire       [31:0]   _zz_16514;
  wire       [23:0]   _zz_16515;
  wire       [31:0]   _zz_16516;
  wire       [15:0]   _zz_16517;
  wire       [31:0]   _zz_16518;
  wire       [31:0]   _zz_16519;
  wire       [31:0]   _zz_16520;
  wire       [31:0]   _zz_16521;
  wire       [31:0]   _zz_16522;
  wire       [23:0]   _zz_16523;
  wire       [31:0]   _zz_16524;
  wire       [15:0]   _zz_16525;
  wire       [31:0]   _zz_16526;
  wire       [31:0]   _zz_16527;
  wire       [31:0]   _zz_16528;
  wire       [31:0]   _zz_16529;
  wire       [31:0]   _zz_16530;
  wire       [23:0]   _zz_16531;
  wire       [31:0]   _zz_16532;
  wire       [15:0]   _zz_16533;
  wire       [15:0]   _zz_16534;
  wire       [31:0]   _zz_16535;
  wire       [31:0]   _zz_16536;
  wire       [15:0]   _zz_16537;
  wire       [31:0]   _zz_16538;
  wire       [31:0]   _zz_16539;
  wire       [31:0]   _zz_16540;
  wire       [15:0]   _zz_16541;
  wire       [31:0]   _zz_16542;
  wire       [31:0]   _zz_16543;
  wire       [31:0]   _zz_16544;
  wire       [31:0]   _zz_16545;
  wire       [31:0]   _zz_16546;
  wire       [31:0]   _zz_16547;
  wire       [23:0]   _zz_16548;
  wire       [31:0]   _zz_16549;
  wire       [15:0]   _zz_16550;
  wire       [31:0]   _zz_16551;
  wire       [31:0]   _zz_16552;
  wire       [31:0]   _zz_16553;
  wire       [31:0]   _zz_16554;
  wire       [31:0]   _zz_16555;
  wire       [23:0]   _zz_16556;
  wire       [31:0]   _zz_16557;
  wire       [15:0]   _zz_16558;
  wire       [31:0]   _zz_16559;
  wire       [31:0]   _zz_16560;
  wire       [31:0]   _zz_16561;
  wire       [31:0]   _zz_16562;
  wire       [31:0]   _zz_16563;
  wire       [23:0]   _zz_16564;
  wire       [31:0]   _zz_16565;
  wire       [15:0]   _zz_16566;
  wire       [31:0]   _zz_16567;
  wire       [31:0]   _zz_16568;
  wire       [31:0]   _zz_16569;
  wire       [31:0]   _zz_16570;
  wire       [31:0]   _zz_16571;
  wire       [23:0]   _zz_16572;
  wire       [31:0]   _zz_16573;
  wire       [15:0]   _zz_16574;
  wire       [15:0]   _zz_16575;
  wire       [31:0]   _zz_16576;
  wire       [31:0]   _zz_16577;
  wire       [15:0]   _zz_16578;
  wire       [31:0]   _zz_16579;
  wire       [31:0]   _zz_16580;
  wire       [31:0]   _zz_16581;
  wire       [15:0]   _zz_16582;
  wire       [31:0]   _zz_16583;
  wire       [31:0]   _zz_16584;
  wire       [31:0]   _zz_16585;
  wire       [31:0]   _zz_16586;
  wire       [31:0]   _zz_16587;
  wire       [31:0]   _zz_16588;
  wire       [23:0]   _zz_16589;
  wire       [31:0]   _zz_16590;
  wire       [15:0]   _zz_16591;
  wire       [31:0]   _zz_16592;
  wire       [31:0]   _zz_16593;
  wire       [31:0]   _zz_16594;
  wire       [31:0]   _zz_16595;
  wire       [31:0]   _zz_16596;
  wire       [23:0]   _zz_16597;
  wire       [31:0]   _zz_16598;
  wire       [15:0]   _zz_16599;
  wire       [31:0]   _zz_16600;
  wire       [31:0]   _zz_16601;
  wire       [31:0]   _zz_16602;
  wire       [31:0]   _zz_16603;
  wire       [31:0]   _zz_16604;
  wire       [23:0]   _zz_16605;
  wire       [31:0]   _zz_16606;
  wire       [15:0]   _zz_16607;
  wire       [31:0]   _zz_16608;
  wire       [31:0]   _zz_16609;
  wire       [31:0]   _zz_16610;
  wire       [31:0]   _zz_16611;
  wire       [31:0]   _zz_16612;
  wire       [23:0]   _zz_16613;
  wire       [31:0]   _zz_16614;
  wire       [15:0]   _zz_16615;
  wire       [15:0]   _zz_16616;
  wire       [31:0]   _zz_16617;
  wire       [31:0]   _zz_16618;
  wire       [15:0]   _zz_16619;
  wire       [31:0]   _zz_16620;
  wire       [31:0]   _zz_16621;
  wire       [31:0]   _zz_16622;
  wire       [15:0]   _zz_16623;
  wire       [31:0]   _zz_16624;
  wire       [31:0]   _zz_16625;
  wire       [31:0]   _zz_16626;
  wire       [31:0]   _zz_16627;
  wire       [31:0]   _zz_16628;
  wire       [31:0]   _zz_16629;
  wire       [23:0]   _zz_16630;
  wire       [31:0]   _zz_16631;
  wire       [15:0]   _zz_16632;
  wire       [31:0]   _zz_16633;
  wire       [31:0]   _zz_16634;
  wire       [31:0]   _zz_16635;
  wire       [31:0]   _zz_16636;
  wire       [31:0]   _zz_16637;
  wire       [23:0]   _zz_16638;
  wire       [31:0]   _zz_16639;
  wire       [15:0]   _zz_16640;
  wire       [31:0]   _zz_16641;
  wire       [31:0]   _zz_16642;
  wire       [31:0]   _zz_16643;
  wire       [31:0]   _zz_16644;
  wire       [31:0]   _zz_16645;
  wire       [23:0]   _zz_16646;
  wire       [31:0]   _zz_16647;
  wire       [15:0]   _zz_16648;
  wire       [31:0]   _zz_16649;
  wire       [31:0]   _zz_16650;
  wire       [31:0]   _zz_16651;
  wire       [31:0]   _zz_16652;
  wire       [31:0]   _zz_16653;
  wire       [23:0]   _zz_16654;
  wire       [31:0]   _zz_16655;
  wire       [15:0]   _zz_16656;
  wire       [15:0]   _zz_16657;
  wire       [31:0]   _zz_16658;
  wire       [31:0]   _zz_16659;
  wire       [15:0]   _zz_16660;
  wire       [31:0]   _zz_16661;
  wire       [31:0]   _zz_16662;
  wire       [31:0]   _zz_16663;
  wire       [15:0]   _zz_16664;
  wire       [31:0]   _zz_16665;
  wire       [31:0]   _zz_16666;
  wire       [31:0]   _zz_16667;
  wire       [31:0]   _zz_16668;
  wire       [31:0]   _zz_16669;
  wire       [31:0]   _zz_16670;
  wire       [23:0]   _zz_16671;
  wire       [31:0]   _zz_16672;
  wire       [15:0]   _zz_16673;
  wire       [31:0]   _zz_16674;
  wire       [31:0]   _zz_16675;
  wire       [31:0]   _zz_16676;
  wire       [31:0]   _zz_16677;
  wire       [31:0]   _zz_16678;
  wire       [23:0]   _zz_16679;
  wire       [31:0]   _zz_16680;
  wire       [15:0]   _zz_16681;
  wire       [31:0]   _zz_16682;
  wire       [31:0]   _zz_16683;
  wire       [31:0]   _zz_16684;
  wire       [31:0]   _zz_16685;
  wire       [31:0]   _zz_16686;
  wire       [23:0]   _zz_16687;
  wire       [31:0]   _zz_16688;
  wire       [15:0]   _zz_16689;
  wire       [31:0]   _zz_16690;
  wire       [31:0]   _zz_16691;
  wire       [31:0]   _zz_16692;
  wire       [31:0]   _zz_16693;
  wire       [31:0]   _zz_16694;
  wire       [23:0]   _zz_16695;
  wire       [31:0]   _zz_16696;
  wire       [15:0]   _zz_16697;
  wire       [15:0]   _zz_16698;
  wire       [31:0]   _zz_16699;
  wire       [31:0]   _zz_16700;
  wire       [15:0]   _zz_16701;
  wire       [31:0]   _zz_16702;
  wire       [31:0]   _zz_16703;
  wire       [31:0]   _zz_16704;
  wire       [15:0]   _zz_16705;
  wire       [31:0]   _zz_16706;
  wire       [31:0]   _zz_16707;
  wire       [31:0]   _zz_16708;
  wire       [31:0]   _zz_16709;
  wire       [31:0]   _zz_16710;
  wire       [31:0]   _zz_16711;
  wire       [23:0]   _zz_16712;
  wire       [31:0]   _zz_16713;
  wire       [15:0]   _zz_16714;
  wire       [31:0]   _zz_16715;
  wire       [31:0]   _zz_16716;
  wire       [31:0]   _zz_16717;
  wire       [31:0]   _zz_16718;
  wire       [31:0]   _zz_16719;
  wire       [23:0]   _zz_16720;
  wire       [31:0]   _zz_16721;
  wire       [15:0]   _zz_16722;
  wire       [31:0]   _zz_16723;
  wire       [31:0]   _zz_16724;
  wire       [31:0]   _zz_16725;
  wire       [31:0]   _zz_16726;
  wire       [31:0]   _zz_16727;
  wire       [23:0]   _zz_16728;
  wire       [31:0]   _zz_16729;
  wire       [15:0]   _zz_16730;
  wire       [31:0]   _zz_16731;
  wire       [31:0]   _zz_16732;
  wire       [31:0]   _zz_16733;
  wire       [31:0]   _zz_16734;
  wire       [31:0]   _zz_16735;
  wire       [23:0]   _zz_16736;
  wire       [31:0]   _zz_16737;
  wire       [15:0]   _zz_16738;
  wire       [15:0]   _zz_16739;
  wire       [31:0]   _zz_16740;
  wire       [31:0]   _zz_16741;
  wire       [15:0]   _zz_16742;
  wire       [31:0]   _zz_16743;
  wire       [31:0]   _zz_16744;
  wire       [31:0]   _zz_16745;
  wire       [15:0]   _zz_16746;
  wire       [31:0]   _zz_16747;
  wire       [31:0]   _zz_16748;
  wire       [31:0]   _zz_16749;
  wire       [31:0]   _zz_16750;
  wire       [31:0]   _zz_16751;
  wire       [31:0]   _zz_16752;
  wire       [23:0]   _zz_16753;
  wire       [31:0]   _zz_16754;
  wire       [15:0]   _zz_16755;
  wire       [31:0]   _zz_16756;
  wire       [31:0]   _zz_16757;
  wire       [31:0]   _zz_16758;
  wire       [31:0]   _zz_16759;
  wire       [31:0]   _zz_16760;
  wire       [23:0]   _zz_16761;
  wire       [31:0]   _zz_16762;
  wire       [15:0]   _zz_16763;
  wire       [31:0]   _zz_16764;
  wire       [31:0]   _zz_16765;
  wire       [31:0]   _zz_16766;
  wire       [31:0]   _zz_16767;
  wire       [31:0]   _zz_16768;
  wire       [23:0]   _zz_16769;
  wire       [31:0]   _zz_16770;
  wire       [15:0]   _zz_16771;
  wire       [31:0]   _zz_16772;
  wire       [31:0]   _zz_16773;
  wire       [31:0]   _zz_16774;
  wire       [31:0]   _zz_16775;
  wire       [31:0]   _zz_16776;
  wire       [23:0]   _zz_16777;
  wire       [31:0]   _zz_16778;
  wire       [15:0]   _zz_16779;
  wire       [15:0]   _zz_16780;
  wire       [31:0]   _zz_16781;
  wire       [31:0]   _zz_16782;
  wire       [15:0]   _zz_16783;
  wire       [31:0]   _zz_16784;
  wire       [31:0]   _zz_16785;
  wire       [31:0]   _zz_16786;
  wire       [15:0]   _zz_16787;
  wire       [31:0]   _zz_16788;
  wire       [31:0]   _zz_16789;
  wire       [31:0]   _zz_16790;
  wire       [31:0]   _zz_16791;
  wire       [31:0]   _zz_16792;
  wire       [31:0]   _zz_16793;
  wire       [23:0]   _zz_16794;
  wire       [31:0]   _zz_16795;
  wire       [15:0]   _zz_16796;
  wire       [31:0]   _zz_16797;
  wire       [31:0]   _zz_16798;
  wire       [31:0]   _zz_16799;
  wire       [31:0]   _zz_16800;
  wire       [31:0]   _zz_16801;
  wire       [23:0]   _zz_16802;
  wire       [31:0]   _zz_16803;
  wire       [15:0]   _zz_16804;
  wire       [31:0]   _zz_16805;
  wire       [31:0]   _zz_16806;
  wire       [31:0]   _zz_16807;
  wire       [31:0]   _zz_16808;
  wire       [31:0]   _zz_16809;
  wire       [23:0]   _zz_16810;
  wire       [31:0]   _zz_16811;
  wire       [15:0]   _zz_16812;
  wire       [31:0]   _zz_16813;
  wire       [31:0]   _zz_16814;
  wire       [31:0]   _zz_16815;
  wire       [31:0]   _zz_16816;
  wire       [31:0]   _zz_16817;
  wire       [23:0]   _zz_16818;
  wire       [31:0]   _zz_16819;
  wire       [15:0]   _zz_16820;
  wire       [15:0]   _zz_16821;
  wire       [31:0]   _zz_16822;
  wire       [31:0]   _zz_16823;
  wire       [15:0]   _zz_16824;
  wire       [31:0]   _zz_16825;
  wire       [31:0]   _zz_16826;
  wire       [31:0]   _zz_16827;
  wire       [15:0]   _zz_16828;
  wire       [31:0]   _zz_16829;
  wire       [31:0]   _zz_16830;
  wire       [31:0]   _zz_16831;
  wire       [31:0]   _zz_16832;
  wire       [31:0]   _zz_16833;
  wire       [31:0]   _zz_16834;
  wire       [23:0]   _zz_16835;
  wire       [31:0]   _zz_16836;
  wire       [15:0]   _zz_16837;
  wire       [31:0]   _zz_16838;
  wire       [31:0]   _zz_16839;
  wire       [31:0]   _zz_16840;
  wire       [31:0]   _zz_16841;
  wire       [31:0]   _zz_16842;
  wire       [23:0]   _zz_16843;
  wire       [31:0]   _zz_16844;
  wire       [15:0]   _zz_16845;
  wire       [31:0]   _zz_16846;
  wire       [31:0]   _zz_16847;
  wire       [31:0]   _zz_16848;
  wire       [31:0]   _zz_16849;
  wire       [31:0]   _zz_16850;
  wire       [23:0]   _zz_16851;
  wire       [31:0]   _zz_16852;
  wire       [15:0]   _zz_16853;
  wire       [31:0]   _zz_16854;
  wire       [31:0]   _zz_16855;
  wire       [31:0]   _zz_16856;
  wire       [31:0]   _zz_16857;
  wire       [31:0]   _zz_16858;
  wire       [23:0]   _zz_16859;
  wire       [31:0]   _zz_16860;
  wire       [15:0]   _zz_16861;
  wire       [15:0]   _zz_16862;
  wire       [31:0]   _zz_16863;
  wire       [31:0]   _zz_16864;
  wire       [15:0]   _zz_16865;
  wire       [31:0]   _zz_16866;
  wire       [31:0]   _zz_16867;
  wire       [31:0]   _zz_16868;
  wire       [15:0]   _zz_16869;
  wire       [31:0]   _zz_16870;
  wire       [31:0]   _zz_16871;
  wire       [31:0]   _zz_16872;
  wire       [31:0]   _zz_16873;
  wire       [31:0]   _zz_16874;
  wire       [31:0]   _zz_16875;
  wire       [23:0]   _zz_16876;
  wire       [31:0]   _zz_16877;
  wire       [15:0]   _zz_16878;
  wire       [31:0]   _zz_16879;
  wire       [31:0]   _zz_16880;
  wire       [31:0]   _zz_16881;
  wire       [31:0]   _zz_16882;
  wire       [31:0]   _zz_16883;
  wire       [23:0]   _zz_16884;
  wire       [31:0]   _zz_16885;
  wire       [15:0]   _zz_16886;
  wire       [31:0]   _zz_16887;
  wire       [31:0]   _zz_16888;
  wire       [31:0]   _zz_16889;
  wire       [31:0]   _zz_16890;
  wire       [31:0]   _zz_16891;
  wire       [23:0]   _zz_16892;
  wire       [31:0]   _zz_16893;
  wire       [15:0]   _zz_16894;
  wire       [31:0]   _zz_16895;
  wire       [31:0]   _zz_16896;
  wire       [31:0]   _zz_16897;
  wire       [31:0]   _zz_16898;
  wire       [31:0]   _zz_16899;
  wire       [23:0]   _zz_16900;
  wire       [31:0]   _zz_16901;
  wire       [15:0]   _zz_16902;
  wire       [15:0]   _zz_16903;
  wire       [31:0]   _zz_16904;
  wire       [31:0]   _zz_16905;
  wire       [15:0]   _zz_16906;
  wire       [31:0]   _zz_16907;
  wire       [31:0]   _zz_16908;
  wire       [31:0]   _zz_16909;
  wire       [15:0]   _zz_16910;
  wire       [31:0]   _zz_16911;
  wire       [31:0]   _zz_16912;
  wire       [31:0]   _zz_16913;
  wire       [31:0]   _zz_16914;
  wire       [31:0]   _zz_16915;
  wire       [31:0]   _zz_16916;
  wire       [23:0]   _zz_16917;
  wire       [31:0]   _zz_16918;
  wire       [15:0]   _zz_16919;
  wire       [31:0]   _zz_16920;
  wire       [31:0]   _zz_16921;
  wire       [31:0]   _zz_16922;
  wire       [31:0]   _zz_16923;
  wire       [31:0]   _zz_16924;
  wire       [23:0]   _zz_16925;
  wire       [31:0]   _zz_16926;
  wire       [15:0]   _zz_16927;
  wire       [31:0]   _zz_16928;
  wire       [31:0]   _zz_16929;
  wire       [31:0]   _zz_16930;
  wire       [31:0]   _zz_16931;
  wire       [31:0]   _zz_16932;
  wire       [23:0]   _zz_16933;
  wire       [31:0]   _zz_16934;
  wire       [15:0]   _zz_16935;
  wire       [31:0]   _zz_16936;
  wire       [31:0]   _zz_16937;
  wire       [31:0]   _zz_16938;
  wire       [31:0]   _zz_16939;
  wire       [31:0]   _zz_16940;
  wire       [23:0]   _zz_16941;
  wire       [31:0]   _zz_16942;
  wire       [15:0]   _zz_16943;
  wire       [15:0]   _zz_16944;
  wire       [31:0]   _zz_16945;
  wire       [31:0]   _zz_16946;
  wire       [15:0]   _zz_16947;
  wire       [31:0]   _zz_16948;
  wire       [31:0]   _zz_16949;
  wire       [31:0]   _zz_16950;
  wire       [15:0]   _zz_16951;
  wire       [31:0]   _zz_16952;
  wire       [31:0]   _zz_16953;
  wire       [31:0]   _zz_16954;
  wire       [31:0]   _zz_16955;
  wire       [31:0]   _zz_16956;
  wire       [31:0]   _zz_16957;
  wire       [23:0]   _zz_16958;
  wire       [31:0]   _zz_16959;
  wire       [15:0]   _zz_16960;
  wire       [31:0]   _zz_16961;
  wire       [31:0]   _zz_16962;
  wire       [31:0]   _zz_16963;
  wire       [31:0]   _zz_16964;
  wire       [31:0]   _zz_16965;
  wire       [23:0]   _zz_16966;
  wire       [31:0]   _zz_16967;
  wire       [15:0]   _zz_16968;
  wire       [31:0]   _zz_16969;
  wire       [31:0]   _zz_16970;
  wire       [31:0]   _zz_16971;
  wire       [31:0]   _zz_16972;
  wire       [31:0]   _zz_16973;
  wire       [23:0]   _zz_16974;
  wire       [31:0]   _zz_16975;
  wire       [15:0]   _zz_16976;
  wire       [31:0]   _zz_16977;
  wire       [31:0]   _zz_16978;
  wire       [31:0]   _zz_16979;
  wire       [31:0]   _zz_16980;
  wire       [31:0]   _zz_16981;
  wire       [23:0]   _zz_16982;
  wire       [31:0]   _zz_16983;
  wire       [15:0]   _zz_16984;
  wire       [15:0]   _zz_16985;
  wire       [31:0]   _zz_16986;
  wire       [31:0]   _zz_16987;
  wire       [15:0]   _zz_16988;
  wire       [31:0]   _zz_16989;
  wire       [31:0]   _zz_16990;
  wire       [31:0]   _zz_16991;
  wire       [15:0]   _zz_16992;
  wire       [31:0]   _zz_16993;
  wire       [31:0]   _zz_16994;
  wire       [31:0]   _zz_16995;
  wire       [31:0]   _zz_16996;
  wire       [31:0]   _zz_16997;
  wire       [31:0]   _zz_16998;
  wire       [23:0]   _zz_16999;
  wire       [31:0]   _zz_17000;
  wire       [15:0]   _zz_17001;
  wire       [31:0]   _zz_17002;
  wire       [31:0]   _zz_17003;
  wire       [31:0]   _zz_17004;
  wire       [31:0]   _zz_17005;
  wire       [31:0]   _zz_17006;
  wire       [23:0]   _zz_17007;
  wire       [31:0]   _zz_17008;
  wire       [15:0]   _zz_17009;
  wire       [31:0]   _zz_17010;
  wire       [31:0]   _zz_17011;
  wire       [31:0]   _zz_17012;
  wire       [31:0]   _zz_17013;
  wire       [31:0]   _zz_17014;
  wire       [23:0]   _zz_17015;
  wire       [31:0]   _zz_17016;
  wire       [15:0]   _zz_17017;
  wire       [31:0]   _zz_17018;
  wire       [31:0]   _zz_17019;
  wire       [31:0]   _zz_17020;
  wire       [31:0]   _zz_17021;
  wire       [31:0]   _zz_17022;
  wire       [23:0]   _zz_17023;
  wire       [31:0]   _zz_17024;
  wire       [15:0]   _zz_17025;
  wire       [15:0]   _zz_17026;
  wire       [31:0]   _zz_17027;
  wire       [31:0]   _zz_17028;
  wire       [15:0]   _zz_17029;
  wire       [31:0]   _zz_17030;
  wire       [31:0]   _zz_17031;
  wire       [31:0]   _zz_17032;
  wire       [15:0]   _zz_17033;
  wire       [31:0]   _zz_17034;
  wire       [31:0]   _zz_17035;
  wire       [31:0]   _zz_17036;
  wire       [31:0]   _zz_17037;
  wire       [31:0]   _zz_17038;
  wire       [31:0]   _zz_17039;
  wire       [23:0]   _zz_17040;
  wire       [31:0]   _zz_17041;
  wire       [15:0]   _zz_17042;
  wire       [31:0]   _zz_17043;
  wire       [31:0]   _zz_17044;
  wire       [31:0]   _zz_17045;
  wire       [31:0]   _zz_17046;
  wire       [31:0]   _zz_17047;
  wire       [23:0]   _zz_17048;
  wire       [31:0]   _zz_17049;
  wire       [15:0]   _zz_17050;
  wire       [31:0]   _zz_17051;
  wire       [31:0]   _zz_17052;
  wire       [31:0]   _zz_17053;
  wire       [31:0]   _zz_17054;
  wire       [31:0]   _zz_17055;
  wire       [23:0]   _zz_17056;
  wire       [31:0]   _zz_17057;
  wire       [15:0]   _zz_17058;
  wire       [31:0]   _zz_17059;
  wire       [31:0]   _zz_17060;
  wire       [31:0]   _zz_17061;
  wire       [31:0]   _zz_17062;
  wire       [31:0]   _zz_17063;
  wire       [23:0]   _zz_17064;
  wire       [31:0]   _zz_17065;
  wire       [15:0]   _zz_17066;
  wire       [15:0]   _zz_17067;
  wire       [31:0]   _zz_17068;
  wire       [31:0]   _zz_17069;
  wire       [15:0]   _zz_17070;
  wire       [31:0]   _zz_17071;
  wire       [31:0]   _zz_17072;
  wire       [31:0]   _zz_17073;
  wire       [15:0]   _zz_17074;
  wire       [31:0]   _zz_17075;
  wire       [31:0]   _zz_17076;
  wire       [31:0]   _zz_17077;
  wire       [31:0]   _zz_17078;
  wire       [31:0]   _zz_17079;
  wire       [31:0]   _zz_17080;
  wire       [23:0]   _zz_17081;
  wire       [31:0]   _zz_17082;
  wire       [15:0]   _zz_17083;
  wire       [31:0]   _zz_17084;
  wire       [31:0]   _zz_17085;
  wire       [31:0]   _zz_17086;
  wire       [31:0]   _zz_17087;
  wire       [31:0]   _zz_17088;
  wire       [23:0]   _zz_17089;
  wire       [31:0]   _zz_17090;
  wire       [15:0]   _zz_17091;
  wire       [31:0]   _zz_17092;
  wire       [31:0]   _zz_17093;
  wire       [31:0]   _zz_17094;
  wire       [31:0]   _zz_17095;
  wire       [31:0]   _zz_17096;
  wire       [23:0]   _zz_17097;
  wire       [31:0]   _zz_17098;
  wire       [15:0]   _zz_17099;
  wire       [31:0]   _zz_17100;
  wire       [31:0]   _zz_17101;
  wire       [31:0]   _zz_17102;
  wire       [31:0]   _zz_17103;
  wire       [31:0]   _zz_17104;
  wire       [23:0]   _zz_17105;
  wire       [31:0]   _zz_17106;
  wire       [15:0]   _zz_17107;
  wire       [15:0]   _zz_17108;
  wire       [31:0]   _zz_17109;
  wire       [31:0]   _zz_17110;
  wire       [15:0]   _zz_17111;
  wire       [31:0]   _zz_17112;
  wire       [31:0]   _zz_17113;
  wire       [31:0]   _zz_17114;
  wire       [15:0]   _zz_17115;
  wire       [31:0]   _zz_17116;
  wire       [31:0]   _zz_17117;
  wire       [31:0]   _zz_17118;
  wire       [31:0]   _zz_17119;
  wire       [31:0]   _zz_17120;
  wire       [31:0]   _zz_17121;
  wire       [23:0]   _zz_17122;
  wire       [31:0]   _zz_17123;
  wire       [15:0]   _zz_17124;
  wire       [31:0]   _zz_17125;
  wire       [31:0]   _zz_17126;
  wire       [31:0]   _zz_17127;
  wire       [31:0]   _zz_17128;
  wire       [31:0]   _zz_17129;
  wire       [23:0]   _zz_17130;
  wire       [31:0]   _zz_17131;
  wire       [15:0]   _zz_17132;
  wire       [31:0]   _zz_17133;
  wire       [31:0]   _zz_17134;
  wire       [31:0]   _zz_17135;
  wire       [31:0]   _zz_17136;
  wire       [31:0]   _zz_17137;
  wire       [23:0]   _zz_17138;
  wire       [31:0]   _zz_17139;
  wire       [15:0]   _zz_17140;
  wire       [31:0]   _zz_17141;
  wire       [31:0]   _zz_17142;
  wire       [31:0]   _zz_17143;
  wire       [31:0]   _zz_17144;
  wire       [31:0]   _zz_17145;
  wire       [23:0]   _zz_17146;
  wire       [31:0]   _zz_17147;
  wire       [15:0]   _zz_17148;
  wire       [15:0]   _zz_17149;
  wire       [31:0]   _zz_17150;
  wire       [31:0]   _zz_17151;
  wire       [15:0]   _zz_17152;
  wire       [31:0]   _zz_17153;
  wire       [31:0]   _zz_17154;
  wire       [31:0]   _zz_17155;
  wire       [15:0]   _zz_17156;
  wire       [31:0]   _zz_17157;
  wire       [31:0]   _zz_17158;
  wire       [31:0]   _zz_17159;
  wire       [31:0]   _zz_17160;
  wire       [31:0]   _zz_17161;
  wire       [31:0]   _zz_17162;
  wire       [23:0]   _zz_17163;
  wire       [31:0]   _zz_17164;
  wire       [15:0]   _zz_17165;
  wire       [31:0]   _zz_17166;
  wire       [31:0]   _zz_17167;
  wire       [31:0]   _zz_17168;
  wire       [31:0]   _zz_17169;
  wire       [31:0]   _zz_17170;
  wire       [23:0]   _zz_17171;
  wire       [31:0]   _zz_17172;
  wire       [15:0]   _zz_17173;
  wire       [31:0]   _zz_17174;
  wire       [31:0]   _zz_17175;
  wire       [31:0]   _zz_17176;
  wire       [31:0]   _zz_17177;
  wire       [31:0]   _zz_17178;
  wire       [23:0]   _zz_17179;
  wire       [31:0]   _zz_17180;
  wire       [15:0]   _zz_17181;
  wire       [31:0]   _zz_17182;
  wire       [31:0]   _zz_17183;
  wire       [31:0]   _zz_17184;
  wire       [31:0]   _zz_17185;
  wire       [31:0]   _zz_17186;
  wire       [23:0]   _zz_17187;
  wire       [31:0]   _zz_17188;
  wire       [15:0]   _zz_17189;
  wire       [15:0]   _zz_17190;
  wire       [31:0]   _zz_17191;
  wire       [31:0]   _zz_17192;
  wire       [15:0]   _zz_17193;
  wire       [31:0]   _zz_17194;
  wire       [31:0]   _zz_17195;
  wire       [31:0]   _zz_17196;
  wire       [15:0]   _zz_17197;
  wire       [31:0]   _zz_17198;
  wire       [31:0]   _zz_17199;
  wire       [31:0]   _zz_17200;
  wire       [31:0]   _zz_17201;
  wire       [31:0]   _zz_17202;
  wire       [31:0]   _zz_17203;
  wire       [23:0]   _zz_17204;
  wire       [31:0]   _zz_17205;
  wire       [15:0]   _zz_17206;
  wire       [31:0]   _zz_17207;
  wire       [31:0]   _zz_17208;
  wire       [31:0]   _zz_17209;
  wire       [31:0]   _zz_17210;
  wire       [31:0]   _zz_17211;
  wire       [23:0]   _zz_17212;
  wire       [31:0]   _zz_17213;
  wire       [15:0]   _zz_17214;
  wire       [31:0]   _zz_17215;
  wire       [31:0]   _zz_17216;
  wire       [31:0]   _zz_17217;
  wire       [31:0]   _zz_17218;
  wire       [31:0]   _zz_17219;
  wire       [23:0]   _zz_17220;
  wire       [31:0]   _zz_17221;
  wire       [15:0]   _zz_17222;
  wire       [31:0]   _zz_17223;
  wire       [31:0]   _zz_17224;
  wire       [31:0]   _zz_17225;
  wire       [31:0]   _zz_17226;
  wire       [31:0]   _zz_17227;
  wire       [23:0]   _zz_17228;
  wire       [31:0]   _zz_17229;
  wire       [15:0]   _zz_17230;
  wire       [15:0]   _zz_17231;
  wire       [31:0]   _zz_17232;
  wire       [31:0]   _zz_17233;
  wire       [15:0]   _zz_17234;
  wire       [31:0]   _zz_17235;
  wire       [31:0]   _zz_17236;
  wire       [31:0]   _zz_17237;
  wire       [15:0]   _zz_17238;
  wire       [31:0]   _zz_17239;
  wire       [31:0]   _zz_17240;
  wire       [31:0]   _zz_17241;
  wire       [31:0]   _zz_17242;
  wire       [31:0]   _zz_17243;
  wire       [31:0]   _zz_17244;
  wire       [23:0]   _zz_17245;
  wire       [31:0]   _zz_17246;
  wire       [15:0]   _zz_17247;
  wire       [31:0]   _zz_17248;
  wire       [31:0]   _zz_17249;
  wire       [31:0]   _zz_17250;
  wire       [31:0]   _zz_17251;
  wire       [31:0]   _zz_17252;
  wire       [23:0]   _zz_17253;
  wire       [31:0]   _zz_17254;
  wire       [15:0]   _zz_17255;
  wire       [31:0]   _zz_17256;
  wire       [31:0]   _zz_17257;
  wire       [31:0]   _zz_17258;
  wire       [31:0]   _zz_17259;
  wire       [31:0]   _zz_17260;
  wire       [23:0]   _zz_17261;
  wire       [31:0]   _zz_17262;
  wire       [15:0]   _zz_17263;
  wire       [31:0]   _zz_17264;
  wire       [31:0]   _zz_17265;
  wire       [31:0]   _zz_17266;
  wire       [31:0]   _zz_17267;
  wire       [31:0]   _zz_17268;
  wire       [23:0]   _zz_17269;
  wire       [31:0]   _zz_17270;
  wire       [15:0]   _zz_17271;
  wire       [15:0]   _zz_17272;
  wire       [31:0]   _zz_17273;
  wire       [31:0]   _zz_17274;
  wire       [15:0]   _zz_17275;
  wire       [31:0]   _zz_17276;
  wire       [31:0]   _zz_17277;
  wire       [31:0]   _zz_17278;
  wire       [15:0]   _zz_17279;
  wire       [31:0]   _zz_17280;
  wire       [31:0]   _zz_17281;
  wire       [31:0]   _zz_17282;
  wire       [31:0]   _zz_17283;
  wire       [31:0]   _zz_17284;
  wire       [31:0]   _zz_17285;
  wire       [23:0]   _zz_17286;
  wire       [31:0]   _zz_17287;
  wire       [15:0]   _zz_17288;
  wire       [31:0]   _zz_17289;
  wire       [31:0]   _zz_17290;
  wire       [31:0]   _zz_17291;
  wire       [31:0]   _zz_17292;
  wire       [31:0]   _zz_17293;
  wire       [23:0]   _zz_17294;
  wire       [31:0]   _zz_17295;
  wire       [15:0]   _zz_17296;
  wire       [31:0]   _zz_17297;
  wire       [31:0]   _zz_17298;
  wire       [31:0]   _zz_17299;
  wire       [31:0]   _zz_17300;
  wire       [31:0]   _zz_17301;
  wire       [23:0]   _zz_17302;
  wire       [31:0]   _zz_17303;
  wire       [15:0]   _zz_17304;
  wire       [31:0]   _zz_17305;
  wire       [31:0]   _zz_17306;
  wire       [31:0]   _zz_17307;
  wire       [31:0]   _zz_17308;
  wire       [31:0]   _zz_17309;
  wire       [23:0]   _zz_17310;
  wire       [31:0]   _zz_17311;
  wire       [15:0]   _zz_17312;
  wire       [15:0]   _zz_17313;
  wire       [31:0]   _zz_17314;
  wire       [31:0]   _zz_17315;
  wire       [15:0]   _zz_17316;
  wire       [31:0]   _zz_17317;
  wire       [31:0]   _zz_17318;
  wire       [31:0]   _zz_17319;
  wire       [15:0]   _zz_17320;
  wire       [31:0]   _zz_17321;
  wire       [31:0]   _zz_17322;
  wire       [31:0]   _zz_17323;
  wire       [31:0]   _zz_17324;
  wire       [31:0]   _zz_17325;
  wire       [31:0]   _zz_17326;
  wire       [23:0]   _zz_17327;
  wire       [31:0]   _zz_17328;
  wire       [15:0]   _zz_17329;
  wire       [31:0]   _zz_17330;
  wire       [31:0]   _zz_17331;
  wire       [31:0]   _zz_17332;
  wire       [31:0]   _zz_17333;
  wire       [31:0]   _zz_17334;
  wire       [23:0]   _zz_17335;
  wire       [31:0]   _zz_17336;
  wire       [15:0]   _zz_17337;
  wire       [31:0]   _zz_17338;
  wire       [31:0]   _zz_17339;
  wire       [31:0]   _zz_17340;
  wire       [31:0]   _zz_17341;
  wire       [31:0]   _zz_17342;
  wire       [23:0]   _zz_17343;
  wire       [31:0]   _zz_17344;
  wire       [15:0]   _zz_17345;
  wire       [31:0]   _zz_17346;
  wire       [31:0]   _zz_17347;
  wire       [31:0]   _zz_17348;
  wire       [31:0]   _zz_17349;
  wire       [31:0]   _zz_17350;
  wire       [23:0]   _zz_17351;
  wire       [31:0]   _zz_17352;
  wire       [15:0]   _zz_17353;
  wire       [15:0]   _zz_17354;
  wire       [31:0]   _zz_17355;
  wire       [31:0]   _zz_17356;
  wire       [15:0]   _zz_17357;
  wire       [31:0]   _zz_17358;
  wire       [31:0]   _zz_17359;
  wire       [31:0]   _zz_17360;
  wire       [15:0]   _zz_17361;
  wire       [31:0]   _zz_17362;
  wire       [31:0]   _zz_17363;
  wire       [31:0]   _zz_17364;
  wire       [31:0]   _zz_17365;
  wire       [31:0]   _zz_17366;
  wire       [31:0]   _zz_17367;
  wire       [23:0]   _zz_17368;
  wire       [31:0]   _zz_17369;
  wire       [15:0]   _zz_17370;
  wire       [31:0]   _zz_17371;
  wire       [31:0]   _zz_17372;
  wire       [31:0]   _zz_17373;
  wire       [31:0]   _zz_17374;
  wire       [31:0]   _zz_17375;
  wire       [23:0]   _zz_17376;
  wire       [31:0]   _zz_17377;
  wire       [15:0]   _zz_17378;
  wire       [31:0]   _zz_17379;
  wire       [31:0]   _zz_17380;
  wire       [31:0]   _zz_17381;
  wire       [31:0]   _zz_17382;
  wire       [31:0]   _zz_17383;
  wire       [23:0]   _zz_17384;
  wire       [31:0]   _zz_17385;
  wire       [15:0]   _zz_17386;
  wire       [31:0]   _zz_17387;
  wire       [31:0]   _zz_17388;
  wire       [31:0]   _zz_17389;
  wire       [31:0]   _zz_17390;
  wire       [31:0]   _zz_17391;
  wire       [23:0]   _zz_17392;
  wire       [31:0]   _zz_17393;
  wire       [15:0]   _zz_17394;
  wire       [15:0]   _zz_17395;
  wire       [31:0]   _zz_17396;
  wire       [31:0]   _zz_17397;
  wire       [15:0]   _zz_17398;
  wire       [31:0]   _zz_17399;
  wire       [31:0]   _zz_17400;
  wire       [31:0]   _zz_17401;
  wire       [15:0]   _zz_17402;
  wire       [31:0]   _zz_17403;
  wire       [31:0]   _zz_17404;
  wire       [31:0]   _zz_17405;
  wire       [31:0]   _zz_17406;
  wire       [31:0]   _zz_17407;
  wire       [31:0]   _zz_17408;
  wire       [23:0]   _zz_17409;
  wire       [31:0]   _zz_17410;
  wire       [15:0]   _zz_17411;
  wire       [31:0]   _zz_17412;
  wire       [31:0]   _zz_17413;
  wire       [31:0]   _zz_17414;
  wire       [31:0]   _zz_17415;
  wire       [31:0]   _zz_17416;
  wire       [23:0]   _zz_17417;
  wire       [31:0]   _zz_17418;
  wire       [15:0]   _zz_17419;
  wire       [31:0]   _zz_17420;
  wire       [31:0]   _zz_17421;
  wire       [31:0]   _zz_17422;
  wire       [31:0]   _zz_17423;
  wire       [31:0]   _zz_17424;
  wire       [23:0]   _zz_17425;
  wire       [31:0]   _zz_17426;
  wire       [15:0]   _zz_17427;
  wire       [31:0]   _zz_17428;
  wire       [31:0]   _zz_17429;
  wire       [31:0]   _zz_17430;
  wire       [31:0]   _zz_17431;
  wire       [31:0]   _zz_17432;
  wire       [23:0]   _zz_17433;
  wire       [31:0]   _zz_17434;
  wire       [15:0]   _zz_17435;
  wire       [15:0]   _zz_17436;
  wire       [31:0]   _zz_17437;
  wire       [31:0]   _zz_17438;
  wire       [15:0]   _zz_17439;
  wire       [31:0]   _zz_17440;
  wire       [31:0]   _zz_17441;
  wire       [31:0]   _zz_17442;
  wire       [15:0]   _zz_17443;
  wire       [31:0]   _zz_17444;
  wire       [31:0]   _zz_17445;
  wire       [31:0]   _zz_17446;
  wire       [31:0]   _zz_17447;
  wire       [31:0]   _zz_17448;
  wire       [31:0]   _zz_17449;
  wire       [23:0]   _zz_17450;
  wire       [31:0]   _zz_17451;
  wire       [15:0]   _zz_17452;
  wire       [31:0]   _zz_17453;
  wire       [31:0]   _zz_17454;
  wire       [31:0]   _zz_17455;
  wire       [31:0]   _zz_17456;
  wire       [31:0]   _zz_17457;
  wire       [23:0]   _zz_17458;
  wire       [31:0]   _zz_17459;
  wire       [15:0]   _zz_17460;
  wire       [31:0]   _zz_17461;
  wire       [31:0]   _zz_17462;
  wire       [31:0]   _zz_17463;
  wire       [31:0]   _zz_17464;
  wire       [31:0]   _zz_17465;
  wire       [23:0]   _zz_17466;
  wire       [31:0]   _zz_17467;
  wire       [15:0]   _zz_17468;
  wire       [31:0]   _zz_17469;
  wire       [31:0]   _zz_17470;
  wire       [31:0]   _zz_17471;
  wire       [31:0]   _zz_17472;
  wire       [31:0]   _zz_17473;
  wire       [23:0]   _zz_17474;
  wire       [31:0]   _zz_17475;
  wire       [15:0]   _zz_17476;
  wire       [15:0]   _zz_17477;
  wire       [31:0]   _zz_17478;
  wire       [31:0]   _zz_17479;
  wire       [15:0]   _zz_17480;
  wire       [31:0]   _zz_17481;
  wire       [31:0]   _zz_17482;
  wire       [31:0]   _zz_17483;
  wire       [15:0]   _zz_17484;
  wire       [31:0]   _zz_17485;
  wire       [31:0]   _zz_17486;
  wire       [31:0]   _zz_17487;
  wire       [31:0]   _zz_17488;
  wire       [31:0]   _zz_17489;
  wire       [31:0]   _zz_17490;
  wire       [23:0]   _zz_17491;
  wire       [31:0]   _zz_17492;
  wire       [15:0]   _zz_17493;
  wire       [31:0]   _zz_17494;
  wire       [31:0]   _zz_17495;
  wire       [31:0]   _zz_17496;
  wire       [31:0]   _zz_17497;
  wire       [31:0]   _zz_17498;
  wire       [23:0]   _zz_17499;
  wire       [31:0]   _zz_17500;
  wire       [15:0]   _zz_17501;
  wire       [31:0]   _zz_17502;
  wire       [31:0]   _zz_17503;
  wire       [31:0]   _zz_17504;
  wire       [31:0]   _zz_17505;
  wire       [31:0]   _zz_17506;
  wire       [23:0]   _zz_17507;
  wire       [31:0]   _zz_17508;
  wire       [15:0]   _zz_17509;
  wire       [31:0]   _zz_17510;
  wire       [31:0]   _zz_17511;
  wire       [31:0]   _zz_17512;
  wire       [31:0]   _zz_17513;
  wire       [31:0]   _zz_17514;
  wire       [23:0]   _zz_17515;
  wire       [31:0]   _zz_17516;
  wire       [15:0]   _zz_17517;
  wire       [15:0]   _zz_17518;
  wire       [31:0]   _zz_17519;
  wire       [31:0]   _zz_17520;
  wire       [15:0]   _zz_17521;
  wire       [31:0]   _zz_17522;
  wire       [31:0]   _zz_17523;
  wire       [31:0]   _zz_17524;
  wire       [15:0]   _zz_17525;
  wire       [31:0]   _zz_17526;
  wire       [31:0]   _zz_17527;
  wire       [31:0]   _zz_17528;
  wire       [31:0]   _zz_17529;
  wire       [31:0]   _zz_17530;
  wire       [31:0]   _zz_17531;
  wire       [23:0]   _zz_17532;
  wire       [31:0]   _zz_17533;
  wire       [15:0]   _zz_17534;
  wire       [31:0]   _zz_17535;
  wire       [31:0]   _zz_17536;
  wire       [31:0]   _zz_17537;
  wire       [31:0]   _zz_17538;
  wire       [31:0]   _zz_17539;
  wire       [23:0]   _zz_17540;
  wire       [31:0]   _zz_17541;
  wire       [15:0]   _zz_17542;
  wire       [31:0]   _zz_17543;
  wire       [31:0]   _zz_17544;
  wire       [31:0]   _zz_17545;
  wire       [31:0]   _zz_17546;
  wire       [31:0]   _zz_17547;
  wire       [23:0]   _zz_17548;
  wire       [31:0]   _zz_17549;
  wire       [15:0]   _zz_17550;
  wire       [31:0]   _zz_17551;
  wire       [31:0]   _zz_17552;
  wire       [31:0]   _zz_17553;
  wire       [31:0]   _zz_17554;
  wire       [31:0]   _zz_17555;
  wire       [23:0]   _zz_17556;
  wire       [31:0]   _zz_17557;
  wire       [15:0]   _zz_17558;
  wire       [15:0]   _zz_17559;
  wire       [31:0]   _zz_17560;
  wire       [31:0]   _zz_17561;
  wire       [15:0]   _zz_17562;
  wire       [31:0]   _zz_17563;
  wire       [31:0]   _zz_17564;
  wire       [31:0]   _zz_17565;
  wire       [15:0]   _zz_17566;
  wire       [31:0]   _zz_17567;
  wire       [31:0]   _zz_17568;
  wire       [31:0]   _zz_17569;
  wire       [31:0]   _zz_17570;
  wire       [31:0]   _zz_17571;
  wire       [31:0]   _zz_17572;
  wire       [23:0]   _zz_17573;
  wire       [31:0]   _zz_17574;
  wire       [15:0]   _zz_17575;
  wire       [31:0]   _zz_17576;
  wire       [31:0]   _zz_17577;
  wire       [31:0]   _zz_17578;
  wire       [31:0]   _zz_17579;
  wire       [31:0]   _zz_17580;
  wire       [23:0]   _zz_17581;
  wire       [31:0]   _zz_17582;
  wire       [15:0]   _zz_17583;
  wire       [31:0]   _zz_17584;
  wire       [31:0]   _zz_17585;
  wire       [31:0]   _zz_17586;
  wire       [31:0]   _zz_17587;
  wire       [31:0]   _zz_17588;
  wire       [23:0]   _zz_17589;
  wire       [31:0]   _zz_17590;
  wire       [15:0]   _zz_17591;
  wire       [31:0]   _zz_17592;
  wire       [31:0]   _zz_17593;
  wire       [31:0]   _zz_17594;
  wire       [31:0]   _zz_17595;
  wire       [31:0]   _zz_17596;
  wire       [23:0]   _zz_17597;
  wire       [31:0]   _zz_17598;
  wire       [15:0]   _zz_17599;
  wire       [15:0]   _zz_17600;
  wire       [31:0]   _zz_17601;
  wire       [31:0]   _zz_17602;
  wire       [15:0]   _zz_17603;
  wire       [31:0]   _zz_17604;
  wire       [31:0]   _zz_17605;
  wire       [31:0]   _zz_17606;
  wire       [15:0]   _zz_17607;
  wire       [31:0]   _zz_17608;
  wire       [31:0]   _zz_17609;
  wire       [31:0]   _zz_17610;
  wire       [31:0]   _zz_17611;
  wire       [31:0]   _zz_17612;
  wire       [31:0]   _zz_17613;
  wire       [23:0]   _zz_17614;
  wire       [31:0]   _zz_17615;
  wire       [15:0]   _zz_17616;
  wire       [31:0]   _zz_17617;
  wire       [31:0]   _zz_17618;
  wire       [31:0]   _zz_17619;
  wire       [31:0]   _zz_17620;
  wire       [31:0]   _zz_17621;
  wire       [23:0]   _zz_17622;
  wire       [31:0]   _zz_17623;
  wire       [15:0]   _zz_17624;
  wire       [31:0]   _zz_17625;
  wire       [31:0]   _zz_17626;
  wire       [31:0]   _zz_17627;
  wire       [31:0]   _zz_17628;
  wire       [31:0]   _zz_17629;
  wire       [23:0]   _zz_17630;
  wire       [31:0]   _zz_17631;
  wire       [15:0]   _zz_17632;
  wire       [31:0]   _zz_17633;
  wire       [31:0]   _zz_17634;
  wire       [31:0]   _zz_17635;
  wire       [31:0]   _zz_17636;
  wire       [31:0]   _zz_17637;
  wire       [23:0]   _zz_17638;
  wire       [31:0]   _zz_17639;
  wire       [15:0]   _zz_17640;
  wire       [15:0]   _zz_17641;
  wire       [31:0]   _zz_17642;
  wire       [31:0]   _zz_17643;
  wire       [15:0]   _zz_17644;
  wire       [31:0]   _zz_17645;
  wire       [31:0]   _zz_17646;
  wire       [31:0]   _zz_17647;
  wire       [15:0]   _zz_17648;
  wire       [31:0]   _zz_17649;
  wire       [31:0]   _zz_17650;
  wire       [31:0]   _zz_17651;
  wire       [31:0]   _zz_17652;
  wire       [31:0]   _zz_17653;
  wire       [31:0]   _zz_17654;
  wire       [23:0]   _zz_17655;
  wire       [31:0]   _zz_17656;
  wire       [15:0]   _zz_17657;
  wire       [31:0]   _zz_17658;
  wire       [31:0]   _zz_17659;
  wire       [31:0]   _zz_17660;
  wire       [31:0]   _zz_17661;
  wire       [31:0]   _zz_17662;
  wire       [23:0]   _zz_17663;
  wire       [31:0]   _zz_17664;
  wire       [15:0]   _zz_17665;
  wire       [31:0]   _zz_17666;
  wire       [31:0]   _zz_17667;
  wire       [31:0]   _zz_17668;
  wire       [31:0]   _zz_17669;
  wire       [31:0]   _zz_17670;
  wire       [23:0]   _zz_17671;
  wire       [31:0]   _zz_17672;
  wire       [15:0]   _zz_17673;
  wire       [31:0]   _zz_17674;
  wire       [31:0]   _zz_17675;
  wire       [31:0]   _zz_17676;
  wire       [31:0]   _zz_17677;
  wire       [31:0]   _zz_17678;
  wire       [23:0]   _zz_17679;
  wire       [31:0]   _zz_17680;
  wire       [15:0]   _zz_17681;
  wire       [15:0]   _zz_17682;
  wire       [31:0]   _zz_17683;
  wire       [31:0]   _zz_17684;
  wire       [15:0]   _zz_17685;
  wire       [31:0]   _zz_17686;
  wire       [31:0]   _zz_17687;
  wire       [31:0]   _zz_17688;
  wire       [15:0]   _zz_17689;
  wire       [31:0]   _zz_17690;
  wire       [31:0]   _zz_17691;
  wire       [31:0]   _zz_17692;
  wire       [31:0]   _zz_17693;
  wire       [31:0]   _zz_17694;
  wire       [31:0]   _zz_17695;
  wire       [23:0]   _zz_17696;
  wire       [31:0]   _zz_17697;
  wire       [15:0]   _zz_17698;
  wire       [31:0]   _zz_17699;
  wire       [31:0]   _zz_17700;
  wire       [31:0]   _zz_17701;
  wire       [31:0]   _zz_17702;
  wire       [31:0]   _zz_17703;
  wire       [23:0]   _zz_17704;
  wire       [31:0]   _zz_17705;
  wire       [15:0]   _zz_17706;
  wire       [31:0]   _zz_17707;
  wire       [31:0]   _zz_17708;
  wire       [31:0]   _zz_17709;
  wire       [31:0]   _zz_17710;
  wire       [31:0]   _zz_17711;
  wire       [23:0]   _zz_17712;
  wire       [31:0]   _zz_17713;
  wire       [15:0]   _zz_17714;
  wire       [31:0]   _zz_17715;
  wire       [31:0]   _zz_17716;
  wire       [31:0]   _zz_17717;
  wire       [31:0]   _zz_17718;
  wire       [31:0]   _zz_17719;
  wire       [23:0]   _zz_17720;
  wire       [31:0]   _zz_17721;
  wire       [15:0]   _zz_17722;
  wire       [15:0]   _zz_17723;
  wire       [31:0]   _zz_17724;
  wire       [31:0]   _zz_17725;
  wire       [15:0]   _zz_17726;
  wire       [31:0]   _zz_17727;
  wire       [31:0]   _zz_17728;
  wire       [31:0]   _zz_17729;
  wire       [15:0]   _zz_17730;
  wire       [31:0]   _zz_17731;
  wire       [31:0]   _zz_17732;
  wire       [31:0]   _zz_17733;
  wire       [31:0]   _zz_17734;
  wire       [31:0]   _zz_17735;
  wire       [31:0]   _zz_17736;
  wire       [23:0]   _zz_17737;
  wire       [31:0]   _zz_17738;
  wire       [15:0]   _zz_17739;
  wire       [31:0]   _zz_17740;
  wire       [31:0]   _zz_17741;
  wire       [31:0]   _zz_17742;
  wire       [31:0]   _zz_17743;
  wire       [31:0]   _zz_17744;
  wire       [23:0]   _zz_17745;
  wire       [31:0]   _zz_17746;
  wire       [15:0]   _zz_17747;
  wire       [31:0]   _zz_17748;
  wire       [31:0]   _zz_17749;
  wire       [31:0]   _zz_17750;
  wire       [31:0]   _zz_17751;
  wire       [31:0]   _zz_17752;
  wire       [23:0]   _zz_17753;
  wire       [31:0]   _zz_17754;
  wire       [15:0]   _zz_17755;
  wire       [31:0]   _zz_17756;
  wire       [31:0]   _zz_17757;
  wire       [31:0]   _zz_17758;
  wire       [31:0]   _zz_17759;
  wire       [31:0]   _zz_17760;
  wire       [23:0]   _zz_17761;
  wire       [31:0]   _zz_17762;
  wire       [15:0]   _zz_17763;
  wire       [15:0]   _zz_17764;
  wire       [31:0]   _zz_17765;
  wire       [31:0]   _zz_17766;
  wire       [15:0]   _zz_17767;
  wire       [31:0]   _zz_17768;
  wire       [31:0]   _zz_17769;
  wire       [31:0]   _zz_17770;
  wire       [15:0]   _zz_17771;
  wire       [31:0]   _zz_17772;
  wire       [31:0]   _zz_17773;
  wire       [31:0]   _zz_17774;
  wire       [31:0]   _zz_17775;
  wire       [31:0]   _zz_17776;
  wire       [31:0]   _zz_17777;
  wire       [23:0]   _zz_17778;
  wire       [31:0]   _zz_17779;
  wire       [15:0]   _zz_17780;
  wire       [31:0]   _zz_17781;
  wire       [31:0]   _zz_17782;
  wire       [31:0]   _zz_17783;
  wire       [31:0]   _zz_17784;
  wire       [31:0]   _zz_17785;
  wire       [23:0]   _zz_17786;
  wire       [31:0]   _zz_17787;
  wire       [15:0]   _zz_17788;
  wire       [31:0]   _zz_17789;
  wire       [31:0]   _zz_17790;
  wire       [31:0]   _zz_17791;
  wire       [31:0]   _zz_17792;
  wire       [31:0]   _zz_17793;
  wire       [23:0]   _zz_17794;
  wire       [31:0]   _zz_17795;
  wire       [15:0]   _zz_17796;
  wire       [31:0]   _zz_17797;
  wire       [31:0]   _zz_17798;
  wire       [31:0]   _zz_17799;
  wire       [31:0]   _zz_17800;
  wire       [31:0]   _zz_17801;
  wire       [23:0]   _zz_17802;
  wire       [31:0]   _zz_17803;
  wire       [15:0]   _zz_17804;
  wire       [15:0]   _zz_17805;
  wire       [31:0]   _zz_17806;
  wire       [31:0]   _zz_17807;
  wire       [15:0]   _zz_17808;
  wire       [31:0]   _zz_17809;
  wire       [31:0]   _zz_17810;
  wire       [31:0]   _zz_17811;
  wire       [15:0]   _zz_17812;
  wire       [31:0]   _zz_17813;
  wire       [31:0]   _zz_17814;
  wire       [31:0]   _zz_17815;
  wire       [31:0]   _zz_17816;
  wire       [31:0]   _zz_17817;
  wire       [31:0]   _zz_17818;
  wire       [23:0]   _zz_17819;
  wire       [31:0]   _zz_17820;
  wire       [15:0]   _zz_17821;
  wire       [31:0]   _zz_17822;
  wire       [31:0]   _zz_17823;
  wire       [31:0]   _zz_17824;
  wire       [31:0]   _zz_17825;
  wire       [31:0]   _zz_17826;
  wire       [23:0]   _zz_17827;
  wire       [31:0]   _zz_17828;
  wire       [15:0]   _zz_17829;
  wire       [31:0]   _zz_17830;
  wire       [31:0]   _zz_17831;
  wire       [31:0]   _zz_17832;
  wire       [31:0]   _zz_17833;
  wire       [31:0]   _zz_17834;
  wire       [23:0]   _zz_17835;
  wire       [31:0]   _zz_17836;
  wire       [15:0]   _zz_17837;
  wire       [31:0]   _zz_17838;
  wire       [31:0]   _zz_17839;
  wire       [31:0]   _zz_17840;
  wire       [31:0]   _zz_17841;
  wire       [31:0]   _zz_17842;
  wire       [23:0]   _zz_17843;
  wire       [31:0]   _zz_17844;
  wire       [15:0]   _zz_17845;
  wire       [15:0]   _zz_17846;
  wire       [31:0]   _zz_17847;
  wire       [31:0]   _zz_17848;
  wire       [15:0]   _zz_17849;
  wire       [31:0]   _zz_17850;
  wire       [31:0]   _zz_17851;
  wire       [31:0]   _zz_17852;
  wire       [15:0]   _zz_17853;
  wire       [31:0]   _zz_17854;
  wire       [31:0]   _zz_17855;
  wire       [31:0]   _zz_17856;
  wire       [31:0]   _zz_17857;
  wire       [31:0]   _zz_17858;
  wire       [31:0]   _zz_17859;
  wire       [23:0]   _zz_17860;
  wire       [31:0]   _zz_17861;
  wire       [15:0]   _zz_17862;
  wire       [31:0]   _zz_17863;
  wire       [31:0]   _zz_17864;
  wire       [31:0]   _zz_17865;
  wire       [31:0]   _zz_17866;
  wire       [31:0]   _zz_17867;
  wire       [23:0]   _zz_17868;
  wire       [31:0]   _zz_17869;
  wire       [15:0]   _zz_17870;
  wire       [31:0]   _zz_17871;
  wire       [31:0]   _zz_17872;
  wire       [31:0]   _zz_17873;
  wire       [31:0]   _zz_17874;
  wire       [31:0]   _zz_17875;
  wire       [23:0]   _zz_17876;
  wire       [31:0]   _zz_17877;
  wire       [15:0]   _zz_17878;
  wire       [31:0]   _zz_17879;
  wire       [31:0]   _zz_17880;
  wire       [31:0]   _zz_17881;
  wire       [31:0]   _zz_17882;
  wire       [31:0]   _zz_17883;
  wire       [23:0]   _zz_17884;
  wire       [31:0]   _zz_17885;
  wire       [15:0]   _zz_17886;
  wire       [15:0]   _zz_17887;
  wire       [31:0]   _zz_17888;
  wire       [31:0]   _zz_17889;
  wire       [15:0]   _zz_17890;
  wire       [31:0]   _zz_17891;
  wire       [31:0]   _zz_17892;
  wire       [31:0]   _zz_17893;
  wire       [15:0]   _zz_17894;
  wire       [31:0]   _zz_17895;
  wire       [31:0]   _zz_17896;
  wire       [31:0]   _zz_17897;
  wire       [31:0]   _zz_17898;
  wire       [31:0]   _zz_17899;
  wire       [31:0]   _zz_17900;
  wire       [23:0]   _zz_17901;
  wire       [31:0]   _zz_17902;
  wire       [15:0]   _zz_17903;
  wire       [31:0]   _zz_17904;
  wire       [31:0]   _zz_17905;
  wire       [31:0]   _zz_17906;
  wire       [31:0]   _zz_17907;
  wire       [31:0]   _zz_17908;
  wire       [23:0]   _zz_17909;
  wire       [31:0]   _zz_17910;
  wire       [15:0]   _zz_17911;
  wire       [31:0]   _zz_17912;
  wire       [31:0]   _zz_17913;
  wire       [31:0]   _zz_17914;
  wire       [31:0]   _zz_17915;
  wire       [31:0]   _zz_17916;
  wire       [23:0]   _zz_17917;
  wire       [31:0]   _zz_17918;
  wire       [15:0]   _zz_17919;
  wire       [31:0]   _zz_17920;
  wire       [31:0]   _zz_17921;
  wire       [31:0]   _zz_17922;
  wire       [31:0]   _zz_17923;
  wire       [31:0]   _zz_17924;
  wire       [23:0]   _zz_17925;
  wire       [31:0]   _zz_17926;
  wire       [15:0]   _zz_17927;
  wire       [15:0]   _zz_17928;
  wire       [31:0]   _zz_17929;
  wire       [31:0]   _zz_17930;
  wire       [15:0]   _zz_17931;
  wire       [31:0]   _zz_17932;
  wire       [31:0]   _zz_17933;
  wire       [31:0]   _zz_17934;
  wire       [15:0]   _zz_17935;
  wire       [31:0]   _zz_17936;
  wire       [31:0]   _zz_17937;
  wire       [31:0]   _zz_17938;
  wire       [31:0]   _zz_17939;
  wire       [31:0]   _zz_17940;
  wire       [31:0]   _zz_17941;
  wire       [23:0]   _zz_17942;
  wire       [31:0]   _zz_17943;
  wire       [15:0]   _zz_17944;
  wire       [31:0]   _zz_17945;
  wire       [31:0]   _zz_17946;
  wire       [31:0]   _zz_17947;
  wire       [31:0]   _zz_17948;
  wire       [31:0]   _zz_17949;
  wire       [23:0]   _zz_17950;
  wire       [31:0]   _zz_17951;
  wire       [15:0]   _zz_17952;
  wire       [31:0]   _zz_17953;
  wire       [31:0]   _zz_17954;
  wire       [31:0]   _zz_17955;
  wire       [31:0]   _zz_17956;
  wire       [31:0]   _zz_17957;
  wire       [23:0]   _zz_17958;
  wire       [31:0]   _zz_17959;
  wire       [15:0]   _zz_17960;
  wire       [31:0]   _zz_17961;
  wire       [31:0]   _zz_17962;
  wire       [31:0]   _zz_17963;
  wire       [31:0]   _zz_17964;
  wire       [31:0]   _zz_17965;
  wire       [23:0]   _zz_17966;
  wire       [31:0]   _zz_17967;
  wire       [15:0]   _zz_17968;
  wire       [15:0]   _zz_17969;
  wire       [31:0]   _zz_17970;
  wire       [31:0]   _zz_17971;
  wire       [15:0]   _zz_17972;
  wire       [31:0]   _zz_17973;
  wire       [31:0]   _zz_17974;
  wire       [31:0]   _zz_17975;
  wire       [15:0]   _zz_17976;
  wire       [31:0]   _zz_17977;
  wire       [31:0]   _zz_17978;
  wire       [31:0]   _zz_17979;
  wire       [31:0]   _zz_17980;
  wire       [31:0]   _zz_17981;
  wire       [31:0]   _zz_17982;
  wire       [23:0]   _zz_17983;
  wire       [31:0]   _zz_17984;
  wire       [15:0]   _zz_17985;
  wire       [31:0]   _zz_17986;
  wire       [31:0]   _zz_17987;
  wire       [31:0]   _zz_17988;
  wire       [31:0]   _zz_17989;
  wire       [31:0]   _zz_17990;
  wire       [23:0]   _zz_17991;
  wire       [31:0]   _zz_17992;
  wire       [15:0]   _zz_17993;
  wire       [31:0]   _zz_17994;
  wire       [31:0]   _zz_17995;
  wire       [31:0]   _zz_17996;
  wire       [31:0]   _zz_17997;
  wire       [31:0]   _zz_17998;
  wire       [23:0]   _zz_17999;
  wire       [31:0]   _zz_18000;
  wire       [15:0]   _zz_18001;
  wire       [31:0]   _zz_18002;
  wire       [31:0]   _zz_18003;
  wire       [31:0]   _zz_18004;
  wire       [31:0]   _zz_18005;
  wire       [31:0]   _zz_18006;
  wire       [23:0]   _zz_18007;
  wire       [31:0]   _zz_18008;
  wire       [15:0]   _zz_18009;
  wire       [15:0]   _zz_18010;
  wire       [31:0]   _zz_18011;
  wire       [31:0]   _zz_18012;
  wire       [15:0]   _zz_18013;
  wire       [31:0]   _zz_18014;
  wire       [31:0]   _zz_18015;
  wire       [31:0]   _zz_18016;
  wire       [15:0]   _zz_18017;
  wire       [31:0]   _zz_18018;
  wire       [31:0]   _zz_18019;
  wire       [31:0]   _zz_18020;
  wire       [31:0]   _zz_18021;
  wire       [31:0]   _zz_18022;
  wire       [31:0]   _zz_18023;
  wire       [23:0]   _zz_18024;
  wire       [31:0]   _zz_18025;
  wire       [15:0]   _zz_18026;
  wire       [31:0]   _zz_18027;
  wire       [31:0]   _zz_18028;
  wire       [31:0]   _zz_18029;
  wire       [31:0]   _zz_18030;
  wire       [31:0]   _zz_18031;
  wire       [23:0]   _zz_18032;
  wire       [31:0]   _zz_18033;
  wire       [15:0]   _zz_18034;
  wire       [31:0]   _zz_18035;
  wire       [31:0]   _zz_18036;
  wire       [31:0]   _zz_18037;
  wire       [31:0]   _zz_18038;
  wire       [31:0]   _zz_18039;
  wire       [23:0]   _zz_18040;
  wire       [31:0]   _zz_18041;
  wire       [15:0]   _zz_18042;
  wire       [31:0]   _zz_18043;
  wire       [31:0]   _zz_18044;
  wire       [31:0]   _zz_18045;
  wire       [31:0]   _zz_18046;
  wire       [31:0]   _zz_18047;
  wire       [23:0]   _zz_18048;
  wire       [31:0]   _zz_18049;
  wire       [15:0]   _zz_18050;
  wire       [15:0]   _zz_18051;
  wire       [31:0]   _zz_18052;
  wire       [31:0]   _zz_18053;
  wire       [15:0]   _zz_18054;
  wire       [31:0]   _zz_18055;
  wire       [31:0]   _zz_18056;
  wire       [31:0]   _zz_18057;
  wire       [15:0]   _zz_18058;
  wire       [31:0]   _zz_18059;
  wire       [31:0]   _zz_18060;
  wire       [31:0]   _zz_18061;
  wire       [31:0]   _zz_18062;
  wire       [31:0]   _zz_18063;
  wire       [31:0]   _zz_18064;
  wire       [23:0]   _zz_18065;
  wire       [31:0]   _zz_18066;
  wire       [15:0]   _zz_18067;
  wire       [31:0]   _zz_18068;
  wire       [31:0]   _zz_18069;
  wire       [31:0]   _zz_18070;
  wire       [31:0]   _zz_18071;
  wire       [31:0]   _zz_18072;
  wire       [23:0]   _zz_18073;
  wire       [31:0]   _zz_18074;
  wire       [15:0]   _zz_18075;
  wire       [31:0]   _zz_18076;
  wire       [31:0]   _zz_18077;
  wire       [31:0]   _zz_18078;
  wire       [31:0]   _zz_18079;
  wire       [31:0]   _zz_18080;
  wire       [23:0]   _zz_18081;
  wire       [31:0]   _zz_18082;
  wire       [15:0]   _zz_18083;
  wire       [31:0]   _zz_18084;
  wire       [31:0]   _zz_18085;
  wire       [31:0]   _zz_18086;
  wire       [31:0]   _zz_18087;
  wire       [31:0]   _zz_18088;
  wire       [23:0]   _zz_18089;
  wire       [31:0]   _zz_18090;
  wire       [15:0]   _zz_18091;
  wire       [15:0]   _zz_18092;
  wire       [31:0]   _zz_18093;
  wire       [31:0]   _zz_18094;
  wire       [15:0]   _zz_18095;
  wire       [31:0]   _zz_18096;
  wire       [31:0]   _zz_18097;
  wire       [31:0]   _zz_18098;
  wire       [15:0]   _zz_18099;
  wire       [31:0]   _zz_18100;
  wire       [31:0]   _zz_18101;
  wire       [31:0]   _zz_18102;
  wire       [31:0]   _zz_18103;
  wire       [31:0]   _zz_18104;
  wire       [31:0]   _zz_18105;
  wire       [23:0]   _zz_18106;
  wire       [31:0]   _zz_18107;
  wire       [15:0]   _zz_18108;
  wire       [31:0]   _zz_18109;
  wire       [31:0]   _zz_18110;
  wire       [31:0]   _zz_18111;
  wire       [31:0]   _zz_18112;
  wire       [31:0]   _zz_18113;
  wire       [23:0]   _zz_18114;
  wire       [31:0]   _zz_18115;
  wire       [15:0]   _zz_18116;
  wire       [31:0]   _zz_18117;
  wire       [31:0]   _zz_18118;
  wire       [31:0]   _zz_18119;
  wire       [31:0]   _zz_18120;
  wire       [31:0]   _zz_18121;
  wire       [23:0]   _zz_18122;
  wire       [31:0]   _zz_18123;
  wire       [15:0]   _zz_18124;
  wire       [31:0]   _zz_18125;
  wire       [31:0]   _zz_18126;
  wire       [31:0]   _zz_18127;
  wire       [31:0]   _zz_18128;
  wire       [31:0]   _zz_18129;
  wire       [23:0]   _zz_18130;
  wire       [31:0]   _zz_18131;
  wire       [15:0]   _zz_18132;
  wire       [15:0]   _zz_18133;
  wire       [31:0]   _zz_18134;
  wire       [31:0]   _zz_18135;
  wire       [15:0]   _zz_18136;
  wire       [31:0]   _zz_18137;
  wire       [31:0]   _zz_18138;
  wire       [31:0]   _zz_18139;
  wire       [15:0]   _zz_18140;
  wire       [31:0]   _zz_18141;
  wire       [31:0]   _zz_18142;
  wire       [31:0]   _zz_18143;
  wire       [31:0]   _zz_18144;
  wire       [31:0]   _zz_18145;
  wire       [31:0]   _zz_18146;
  wire       [23:0]   _zz_18147;
  wire       [31:0]   _zz_18148;
  wire       [15:0]   _zz_18149;
  wire       [31:0]   _zz_18150;
  wire       [31:0]   _zz_18151;
  wire       [31:0]   _zz_18152;
  wire       [31:0]   _zz_18153;
  wire       [31:0]   _zz_18154;
  wire       [23:0]   _zz_18155;
  wire       [31:0]   _zz_18156;
  wire       [15:0]   _zz_18157;
  wire       [31:0]   _zz_18158;
  wire       [31:0]   _zz_18159;
  wire       [31:0]   _zz_18160;
  wire       [31:0]   _zz_18161;
  wire       [31:0]   _zz_18162;
  wire       [23:0]   _zz_18163;
  wire       [31:0]   _zz_18164;
  wire       [15:0]   _zz_18165;
  wire       [31:0]   _zz_18166;
  wire       [31:0]   _zz_18167;
  wire       [31:0]   _zz_18168;
  wire       [31:0]   _zz_18169;
  wire       [31:0]   _zz_18170;
  wire       [23:0]   _zz_18171;
  wire       [31:0]   _zz_18172;
  wire       [15:0]   _zz_18173;
  wire       [15:0]   _zz_18174;
  wire       [31:0]   _zz_18175;
  wire       [31:0]   _zz_18176;
  wire       [15:0]   _zz_18177;
  wire       [31:0]   _zz_18178;
  wire       [31:0]   _zz_18179;
  wire       [31:0]   _zz_18180;
  wire       [15:0]   _zz_18181;
  wire       [31:0]   _zz_18182;
  wire       [31:0]   _zz_18183;
  wire       [31:0]   _zz_18184;
  wire       [31:0]   _zz_18185;
  wire       [31:0]   _zz_18186;
  wire       [31:0]   _zz_18187;
  wire       [23:0]   _zz_18188;
  wire       [31:0]   _zz_18189;
  wire       [15:0]   _zz_18190;
  wire       [31:0]   _zz_18191;
  wire       [31:0]   _zz_18192;
  wire       [31:0]   _zz_18193;
  wire       [31:0]   _zz_18194;
  wire       [31:0]   _zz_18195;
  wire       [23:0]   _zz_18196;
  wire       [31:0]   _zz_18197;
  wire       [15:0]   _zz_18198;
  wire       [31:0]   _zz_18199;
  wire       [31:0]   _zz_18200;
  wire       [31:0]   _zz_18201;
  wire       [31:0]   _zz_18202;
  wire       [31:0]   _zz_18203;
  wire       [23:0]   _zz_18204;
  wire       [31:0]   _zz_18205;
  wire       [15:0]   _zz_18206;
  wire       [31:0]   _zz_18207;
  wire       [31:0]   _zz_18208;
  wire       [31:0]   _zz_18209;
  wire       [31:0]   _zz_18210;
  wire       [31:0]   _zz_18211;
  wire       [23:0]   _zz_18212;
  wire       [31:0]   _zz_18213;
  wire       [15:0]   _zz_18214;
  wire       [15:0]   _zz_18215;
  wire       [31:0]   _zz_18216;
  wire       [31:0]   _zz_18217;
  wire       [15:0]   _zz_18218;
  wire       [31:0]   _zz_18219;
  wire       [31:0]   _zz_18220;
  wire       [31:0]   _zz_18221;
  wire       [15:0]   _zz_18222;
  wire       [31:0]   _zz_18223;
  wire       [31:0]   _zz_18224;
  wire       [31:0]   _zz_18225;
  wire       [31:0]   _zz_18226;
  wire       [31:0]   _zz_18227;
  wire       [31:0]   _zz_18228;
  wire       [23:0]   _zz_18229;
  wire       [31:0]   _zz_18230;
  wire       [15:0]   _zz_18231;
  wire       [31:0]   _zz_18232;
  wire       [31:0]   _zz_18233;
  wire       [31:0]   _zz_18234;
  wire       [31:0]   _zz_18235;
  wire       [31:0]   _zz_18236;
  wire       [23:0]   _zz_18237;
  wire       [31:0]   _zz_18238;
  wire       [15:0]   _zz_18239;
  wire       [31:0]   _zz_18240;
  wire       [31:0]   _zz_18241;
  wire       [31:0]   _zz_18242;
  wire       [31:0]   _zz_18243;
  wire       [31:0]   _zz_18244;
  wire       [23:0]   _zz_18245;
  wire       [31:0]   _zz_18246;
  wire       [15:0]   _zz_18247;
  wire       [31:0]   _zz_18248;
  wire       [31:0]   _zz_18249;
  wire       [31:0]   _zz_18250;
  wire       [31:0]   _zz_18251;
  wire       [31:0]   _zz_18252;
  wire       [23:0]   _zz_18253;
  wire       [31:0]   _zz_18254;
  wire       [15:0]   _zz_18255;
  wire       [15:0]   _zz_18256;
  wire       [31:0]   _zz_18257;
  wire       [31:0]   _zz_18258;
  wire       [15:0]   _zz_18259;
  wire       [31:0]   _zz_18260;
  wire       [31:0]   _zz_18261;
  wire       [31:0]   _zz_18262;
  wire       [15:0]   _zz_18263;
  wire       [31:0]   _zz_18264;
  wire       [31:0]   _zz_18265;
  wire       [31:0]   _zz_18266;
  wire       [31:0]   _zz_18267;
  wire       [31:0]   _zz_18268;
  wire       [31:0]   _zz_18269;
  wire       [23:0]   _zz_18270;
  wire       [31:0]   _zz_18271;
  wire       [15:0]   _zz_18272;
  wire       [31:0]   _zz_18273;
  wire       [31:0]   _zz_18274;
  wire       [31:0]   _zz_18275;
  wire       [31:0]   _zz_18276;
  wire       [31:0]   _zz_18277;
  wire       [23:0]   _zz_18278;
  wire       [31:0]   _zz_18279;
  wire       [15:0]   _zz_18280;
  wire       [31:0]   _zz_18281;
  wire       [31:0]   _zz_18282;
  wire       [31:0]   _zz_18283;
  wire       [31:0]   _zz_18284;
  wire       [31:0]   _zz_18285;
  wire       [23:0]   _zz_18286;
  wire       [31:0]   _zz_18287;
  wire       [15:0]   _zz_18288;
  wire       [31:0]   _zz_18289;
  wire       [31:0]   _zz_18290;
  wire       [31:0]   _zz_18291;
  wire       [31:0]   _zz_18292;
  wire       [31:0]   _zz_18293;
  wire       [23:0]   _zz_18294;
  wire       [31:0]   _zz_18295;
  wire       [15:0]   _zz_18296;
  wire       [15:0]   _zz_18297;
  wire       [31:0]   _zz_18298;
  wire       [31:0]   _zz_18299;
  wire       [15:0]   _zz_18300;
  wire       [31:0]   _zz_18301;
  wire       [31:0]   _zz_18302;
  wire       [31:0]   _zz_18303;
  wire       [15:0]   _zz_18304;
  wire       [31:0]   _zz_18305;
  wire       [31:0]   _zz_18306;
  wire       [31:0]   _zz_18307;
  wire       [31:0]   _zz_18308;
  wire       [31:0]   _zz_18309;
  wire       [31:0]   _zz_18310;
  wire       [23:0]   _zz_18311;
  wire       [31:0]   _zz_18312;
  wire       [15:0]   _zz_18313;
  wire       [31:0]   _zz_18314;
  wire       [31:0]   _zz_18315;
  wire       [31:0]   _zz_18316;
  wire       [31:0]   _zz_18317;
  wire       [31:0]   _zz_18318;
  wire       [23:0]   _zz_18319;
  wire       [31:0]   _zz_18320;
  wire       [15:0]   _zz_18321;
  wire       [31:0]   _zz_18322;
  wire       [31:0]   _zz_18323;
  wire       [31:0]   _zz_18324;
  wire       [31:0]   _zz_18325;
  wire       [31:0]   _zz_18326;
  wire       [23:0]   _zz_18327;
  wire       [31:0]   _zz_18328;
  wire       [15:0]   _zz_18329;
  wire       [31:0]   _zz_18330;
  wire       [31:0]   _zz_18331;
  wire       [31:0]   _zz_18332;
  wire       [31:0]   _zz_18333;
  wire       [31:0]   _zz_18334;
  wire       [23:0]   _zz_18335;
  wire       [31:0]   _zz_18336;
  wire       [15:0]   _zz_18337;
  wire       [15:0]   _zz_18338;
  wire       [31:0]   _zz_18339;
  wire       [31:0]   _zz_18340;
  wire       [15:0]   _zz_18341;
  wire       [31:0]   _zz_18342;
  wire       [31:0]   _zz_18343;
  wire       [31:0]   _zz_18344;
  wire       [15:0]   _zz_18345;
  wire       [31:0]   _zz_18346;
  wire       [31:0]   _zz_18347;
  wire       [31:0]   _zz_18348;
  wire       [31:0]   _zz_18349;
  wire       [31:0]   _zz_18350;
  wire       [31:0]   _zz_18351;
  wire       [23:0]   _zz_18352;
  wire       [31:0]   _zz_18353;
  wire       [15:0]   _zz_18354;
  wire       [31:0]   _zz_18355;
  wire       [31:0]   _zz_18356;
  wire       [31:0]   _zz_18357;
  wire       [31:0]   _zz_18358;
  wire       [31:0]   _zz_18359;
  wire       [23:0]   _zz_18360;
  wire       [31:0]   _zz_18361;
  wire       [15:0]   _zz_18362;
  wire       [31:0]   _zz_18363;
  wire       [31:0]   _zz_18364;
  wire       [31:0]   _zz_18365;
  wire       [31:0]   _zz_18366;
  wire       [31:0]   _zz_18367;
  wire       [23:0]   _zz_18368;
  wire       [31:0]   _zz_18369;
  wire       [15:0]   _zz_18370;
  wire       [31:0]   _zz_18371;
  wire       [31:0]   _zz_18372;
  wire       [31:0]   _zz_18373;
  wire       [31:0]   _zz_18374;
  wire       [31:0]   _zz_18375;
  wire       [23:0]   _zz_18376;
  wire       [31:0]   _zz_18377;
  wire       [15:0]   _zz_18378;
  wire       [15:0]   _zz_18379;
  wire       [31:0]   _zz_18380;
  wire       [31:0]   _zz_18381;
  wire       [15:0]   _zz_18382;
  wire       [31:0]   _zz_18383;
  wire       [31:0]   _zz_18384;
  wire       [31:0]   _zz_18385;
  wire       [15:0]   _zz_18386;
  wire       [31:0]   _zz_18387;
  wire       [31:0]   _zz_18388;
  wire       [31:0]   _zz_18389;
  wire       [31:0]   _zz_18390;
  wire       [31:0]   _zz_18391;
  wire       [31:0]   _zz_18392;
  wire       [23:0]   _zz_18393;
  wire       [31:0]   _zz_18394;
  wire       [15:0]   _zz_18395;
  wire       [31:0]   _zz_18396;
  wire       [31:0]   _zz_18397;
  wire       [31:0]   _zz_18398;
  wire       [31:0]   _zz_18399;
  wire       [31:0]   _zz_18400;
  wire       [23:0]   _zz_18401;
  wire       [31:0]   _zz_18402;
  wire       [15:0]   _zz_18403;
  wire       [31:0]   _zz_18404;
  wire       [31:0]   _zz_18405;
  wire       [31:0]   _zz_18406;
  wire       [31:0]   _zz_18407;
  wire       [31:0]   _zz_18408;
  wire       [23:0]   _zz_18409;
  wire       [31:0]   _zz_18410;
  wire       [15:0]   _zz_18411;
  wire       [31:0]   _zz_18412;
  wire       [31:0]   _zz_18413;
  wire       [31:0]   _zz_18414;
  wire       [31:0]   _zz_18415;
  wire       [31:0]   _zz_18416;
  wire       [23:0]   _zz_18417;
  wire       [31:0]   _zz_18418;
  wire       [15:0]   _zz_18419;
  wire       [15:0]   _zz_18420;
  wire       [31:0]   _zz_18421;
  wire       [31:0]   _zz_18422;
  wire       [15:0]   _zz_18423;
  wire       [31:0]   _zz_18424;
  wire       [31:0]   _zz_18425;
  wire       [31:0]   _zz_18426;
  wire       [15:0]   _zz_18427;
  wire       [31:0]   _zz_18428;
  wire       [31:0]   _zz_18429;
  wire       [31:0]   _zz_18430;
  wire       [31:0]   _zz_18431;
  wire       [31:0]   _zz_18432;
  wire       [31:0]   _zz_18433;
  wire       [23:0]   _zz_18434;
  wire       [31:0]   _zz_18435;
  wire       [15:0]   _zz_18436;
  wire       [31:0]   _zz_18437;
  wire       [31:0]   _zz_18438;
  wire       [31:0]   _zz_18439;
  wire       [31:0]   _zz_18440;
  wire       [31:0]   _zz_18441;
  wire       [23:0]   _zz_18442;
  wire       [31:0]   _zz_18443;
  wire       [15:0]   _zz_18444;
  wire       [31:0]   _zz_18445;
  wire       [31:0]   _zz_18446;
  wire       [31:0]   _zz_18447;
  wire       [31:0]   _zz_18448;
  wire       [31:0]   _zz_18449;
  wire       [23:0]   _zz_18450;
  wire       [31:0]   _zz_18451;
  wire       [15:0]   _zz_18452;
  wire       [31:0]   _zz_18453;
  wire       [31:0]   _zz_18454;
  wire       [31:0]   _zz_18455;
  wire       [31:0]   _zz_18456;
  wire       [31:0]   _zz_18457;
  wire       [23:0]   _zz_18458;
  wire       [31:0]   _zz_18459;
  wire       [15:0]   _zz_18460;
  wire       [15:0]   _zz_18461;
  wire       [31:0]   _zz_18462;
  wire       [31:0]   _zz_18463;
  wire       [15:0]   _zz_18464;
  wire       [31:0]   _zz_18465;
  wire       [31:0]   _zz_18466;
  wire       [31:0]   _zz_18467;
  wire       [15:0]   _zz_18468;
  wire       [31:0]   _zz_18469;
  wire       [31:0]   _zz_18470;
  wire       [31:0]   _zz_18471;
  wire       [31:0]   _zz_18472;
  wire       [31:0]   _zz_18473;
  wire       [31:0]   _zz_18474;
  wire       [23:0]   _zz_18475;
  wire       [31:0]   _zz_18476;
  wire       [15:0]   _zz_18477;
  wire       [31:0]   _zz_18478;
  wire       [31:0]   _zz_18479;
  wire       [31:0]   _zz_18480;
  wire       [31:0]   _zz_18481;
  wire       [31:0]   _zz_18482;
  wire       [23:0]   _zz_18483;
  wire       [31:0]   _zz_18484;
  wire       [15:0]   _zz_18485;
  wire       [31:0]   _zz_18486;
  wire       [31:0]   _zz_18487;
  wire       [31:0]   _zz_18488;
  wire       [31:0]   _zz_18489;
  wire       [31:0]   _zz_18490;
  wire       [23:0]   _zz_18491;
  wire       [31:0]   _zz_18492;
  wire       [15:0]   _zz_18493;
  wire       [31:0]   _zz_18494;
  wire       [31:0]   _zz_18495;
  wire       [31:0]   _zz_18496;
  wire       [31:0]   _zz_18497;
  wire       [31:0]   _zz_18498;
  wire       [23:0]   _zz_18499;
  wire       [31:0]   _zz_18500;
  wire       [15:0]   _zz_18501;
  wire       [15:0]   _zz_18502;
  wire       [31:0]   _zz_18503;
  wire       [31:0]   _zz_18504;
  wire       [15:0]   _zz_18505;
  wire       [31:0]   _zz_18506;
  wire       [31:0]   _zz_18507;
  wire       [31:0]   _zz_18508;
  wire       [15:0]   _zz_18509;
  wire       [31:0]   _zz_18510;
  wire       [31:0]   _zz_18511;
  wire       [31:0]   _zz_18512;
  wire       [31:0]   _zz_18513;
  wire       [31:0]   _zz_18514;
  wire       [31:0]   _zz_18515;
  wire       [23:0]   _zz_18516;
  wire       [31:0]   _zz_18517;
  wire       [15:0]   _zz_18518;
  wire       [31:0]   _zz_18519;
  wire       [31:0]   _zz_18520;
  wire       [31:0]   _zz_18521;
  wire       [31:0]   _zz_18522;
  wire       [31:0]   _zz_18523;
  wire       [23:0]   _zz_18524;
  wire       [31:0]   _zz_18525;
  wire       [15:0]   _zz_18526;
  wire       [31:0]   _zz_18527;
  wire       [31:0]   _zz_18528;
  wire       [31:0]   _zz_18529;
  wire       [31:0]   _zz_18530;
  wire       [31:0]   _zz_18531;
  wire       [23:0]   _zz_18532;
  wire       [31:0]   _zz_18533;
  wire       [15:0]   _zz_18534;
  wire       [31:0]   _zz_18535;
  wire       [31:0]   _zz_18536;
  wire       [31:0]   _zz_18537;
  wire       [31:0]   _zz_18538;
  wire       [31:0]   _zz_18539;
  wire       [23:0]   _zz_18540;
  wire       [31:0]   _zz_18541;
  wire       [15:0]   _zz_18542;
  wire       [15:0]   _zz_18543;
  wire       [31:0]   _zz_18544;
  wire       [31:0]   _zz_18545;
  wire       [15:0]   _zz_18546;
  wire       [31:0]   _zz_18547;
  wire       [31:0]   _zz_18548;
  wire       [31:0]   _zz_18549;
  wire       [15:0]   _zz_18550;
  wire       [31:0]   _zz_18551;
  wire       [31:0]   _zz_18552;
  wire       [31:0]   _zz_18553;
  wire       [31:0]   _zz_18554;
  wire       [31:0]   _zz_18555;
  wire       [31:0]   _zz_18556;
  wire       [23:0]   _zz_18557;
  wire       [31:0]   _zz_18558;
  wire       [15:0]   _zz_18559;
  wire       [31:0]   _zz_18560;
  wire       [31:0]   _zz_18561;
  wire       [31:0]   _zz_18562;
  wire       [31:0]   _zz_18563;
  wire       [31:0]   _zz_18564;
  wire       [23:0]   _zz_18565;
  wire       [31:0]   _zz_18566;
  wire       [15:0]   _zz_18567;
  wire       [31:0]   _zz_18568;
  wire       [31:0]   _zz_18569;
  wire       [31:0]   _zz_18570;
  wire       [31:0]   _zz_18571;
  wire       [31:0]   _zz_18572;
  wire       [23:0]   _zz_18573;
  wire       [31:0]   _zz_18574;
  wire       [15:0]   _zz_18575;
  wire       [31:0]   _zz_18576;
  wire       [31:0]   _zz_18577;
  wire       [31:0]   _zz_18578;
  wire       [31:0]   _zz_18579;
  wire       [31:0]   _zz_18580;
  wire       [23:0]   _zz_18581;
  wire       [31:0]   _zz_18582;
  wire       [15:0]   _zz_18583;
  wire       [15:0]   _zz_18584;
  wire       [31:0]   _zz_18585;
  wire       [31:0]   _zz_18586;
  wire       [15:0]   _zz_18587;
  wire       [31:0]   _zz_18588;
  wire       [31:0]   _zz_18589;
  wire       [31:0]   _zz_18590;
  wire       [15:0]   _zz_18591;
  wire       [31:0]   _zz_18592;
  wire       [31:0]   _zz_18593;
  wire       [31:0]   _zz_18594;
  wire       [31:0]   _zz_18595;
  wire       [31:0]   _zz_18596;
  wire       [31:0]   _zz_18597;
  wire       [23:0]   _zz_18598;
  wire       [31:0]   _zz_18599;
  wire       [15:0]   _zz_18600;
  wire       [31:0]   _zz_18601;
  wire       [31:0]   _zz_18602;
  wire       [31:0]   _zz_18603;
  wire       [31:0]   _zz_18604;
  wire       [31:0]   _zz_18605;
  wire       [23:0]   _zz_18606;
  wire       [31:0]   _zz_18607;
  wire       [15:0]   _zz_18608;
  wire       [31:0]   _zz_18609;
  wire       [31:0]   _zz_18610;
  wire       [31:0]   _zz_18611;
  wire       [31:0]   _zz_18612;
  wire       [31:0]   _zz_18613;
  wire       [23:0]   _zz_18614;
  wire       [31:0]   _zz_18615;
  wire       [15:0]   _zz_18616;
  wire       [31:0]   _zz_18617;
  wire       [31:0]   _zz_18618;
  wire       [31:0]   _zz_18619;
  wire       [31:0]   _zz_18620;
  wire       [31:0]   _zz_18621;
  wire       [23:0]   _zz_18622;
  wire       [31:0]   _zz_18623;
  wire       [15:0]   _zz_18624;
  wire       [15:0]   _zz_18625;
  wire       [31:0]   _zz_18626;
  wire       [31:0]   _zz_18627;
  wire       [15:0]   _zz_18628;
  wire       [31:0]   _zz_18629;
  wire       [31:0]   _zz_18630;
  wire       [31:0]   _zz_18631;
  wire       [15:0]   _zz_18632;
  wire       [31:0]   _zz_18633;
  wire       [31:0]   _zz_18634;
  wire       [31:0]   _zz_18635;
  wire       [31:0]   _zz_18636;
  wire       [31:0]   _zz_18637;
  wire       [31:0]   _zz_18638;
  wire       [23:0]   _zz_18639;
  wire       [31:0]   _zz_18640;
  wire       [15:0]   _zz_18641;
  wire       [31:0]   _zz_18642;
  wire       [31:0]   _zz_18643;
  wire       [31:0]   _zz_18644;
  wire       [31:0]   _zz_18645;
  wire       [31:0]   _zz_18646;
  wire       [23:0]   _zz_18647;
  wire       [31:0]   _zz_18648;
  wire       [15:0]   _zz_18649;
  wire       [31:0]   _zz_18650;
  wire       [31:0]   _zz_18651;
  wire       [31:0]   _zz_18652;
  wire       [31:0]   _zz_18653;
  wire       [31:0]   _zz_18654;
  wire       [23:0]   _zz_18655;
  wire       [31:0]   _zz_18656;
  wire       [15:0]   _zz_18657;
  wire       [31:0]   _zz_18658;
  wire       [31:0]   _zz_18659;
  wire       [31:0]   _zz_18660;
  wire       [31:0]   _zz_18661;
  wire       [31:0]   _zz_18662;
  wire       [23:0]   _zz_18663;
  wire       [31:0]   _zz_18664;
  wire       [15:0]   _zz_18665;
  wire       [15:0]   _zz_18666;
  wire       [31:0]   _zz_18667;
  wire       [31:0]   _zz_18668;
  wire       [15:0]   _zz_18669;
  wire       [31:0]   _zz_18670;
  wire       [31:0]   _zz_18671;
  wire       [31:0]   _zz_18672;
  wire       [15:0]   _zz_18673;
  wire       [31:0]   _zz_18674;
  wire       [31:0]   _zz_18675;
  wire       [31:0]   _zz_18676;
  wire       [31:0]   _zz_18677;
  wire       [31:0]   _zz_18678;
  wire       [31:0]   _zz_18679;
  wire       [23:0]   _zz_18680;
  wire       [31:0]   _zz_18681;
  wire       [15:0]   _zz_18682;
  wire       [31:0]   _zz_18683;
  wire       [31:0]   _zz_18684;
  wire       [31:0]   _zz_18685;
  wire       [31:0]   _zz_18686;
  wire       [31:0]   _zz_18687;
  wire       [23:0]   _zz_18688;
  wire       [31:0]   _zz_18689;
  wire       [15:0]   _zz_18690;
  wire       [31:0]   _zz_18691;
  wire       [31:0]   _zz_18692;
  wire       [31:0]   _zz_18693;
  wire       [31:0]   _zz_18694;
  wire       [31:0]   _zz_18695;
  wire       [23:0]   _zz_18696;
  wire       [31:0]   _zz_18697;
  wire       [15:0]   _zz_18698;
  wire       [31:0]   _zz_18699;
  wire       [31:0]   _zz_18700;
  wire       [31:0]   _zz_18701;
  wire       [31:0]   _zz_18702;
  wire       [31:0]   _zz_18703;
  wire       [23:0]   _zz_18704;
  wire       [31:0]   _zz_18705;
  wire       [15:0]   _zz_18706;
  wire       [15:0]   _zz_18707;
  wire       [31:0]   _zz_18708;
  wire       [31:0]   _zz_18709;
  wire       [15:0]   _zz_18710;
  wire       [31:0]   _zz_18711;
  wire       [31:0]   _zz_18712;
  wire       [31:0]   _zz_18713;
  wire       [15:0]   _zz_18714;
  wire       [31:0]   _zz_18715;
  wire       [31:0]   _zz_18716;
  wire       [31:0]   _zz_18717;
  wire       [31:0]   _zz_18718;
  wire       [31:0]   _zz_18719;
  wire       [31:0]   _zz_18720;
  wire       [23:0]   _zz_18721;
  wire       [31:0]   _zz_18722;
  wire       [15:0]   _zz_18723;
  wire       [31:0]   _zz_18724;
  wire       [31:0]   _zz_18725;
  wire       [31:0]   _zz_18726;
  wire       [31:0]   _zz_18727;
  wire       [31:0]   _zz_18728;
  wire       [23:0]   _zz_18729;
  wire       [31:0]   _zz_18730;
  wire       [15:0]   _zz_18731;
  wire       [31:0]   _zz_18732;
  wire       [31:0]   _zz_18733;
  wire       [31:0]   _zz_18734;
  wire       [31:0]   _zz_18735;
  wire       [31:0]   _zz_18736;
  wire       [23:0]   _zz_18737;
  wire       [31:0]   _zz_18738;
  wire       [15:0]   _zz_18739;
  wire       [31:0]   _zz_18740;
  wire       [31:0]   _zz_18741;
  wire       [31:0]   _zz_18742;
  wire       [31:0]   _zz_18743;
  wire       [31:0]   _zz_18744;
  wire       [23:0]   _zz_18745;
  wire       [31:0]   _zz_18746;
  wire       [15:0]   _zz_18747;
  wire       [15:0]   _zz_18748;
  wire       [31:0]   _zz_18749;
  wire       [31:0]   _zz_18750;
  wire       [15:0]   _zz_18751;
  wire       [31:0]   _zz_18752;
  wire       [31:0]   _zz_18753;
  wire       [31:0]   _zz_18754;
  wire       [15:0]   _zz_18755;
  wire       [31:0]   _zz_18756;
  wire       [31:0]   _zz_18757;
  wire       [31:0]   _zz_18758;
  wire       [31:0]   _zz_18759;
  wire       [31:0]   _zz_18760;
  wire       [31:0]   _zz_18761;
  wire       [23:0]   _zz_18762;
  wire       [31:0]   _zz_18763;
  wire       [15:0]   _zz_18764;
  wire       [31:0]   _zz_18765;
  wire       [31:0]   _zz_18766;
  wire       [31:0]   _zz_18767;
  wire       [31:0]   _zz_18768;
  wire       [31:0]   _zz_18769;
  wire       [23:0]   _zz_18770;
  wire       [31:0]   _zz_18771;
  wire       [15:0]   _zz_18772;
  wire       [31:0]   _zz_18773;
  wire       [31:0]   _zz_18774;
  wire       [31:0]   _zz_18775;
  wire       [31:0]   _zz_18776;
  wire       [31:0]   _zz_18777;
  wire       [23:0]   _zz_18778;
  wire       [31:0]   _zz_18779;
  wire       [15:0]   _zz_18780;
  wire       [31:0]   _zz_18781;
  wire       [31:0]   _zz_18782;
  wire       [31:0]   _zz_18783;
  wire       [31:0]   _zz_18784;
  wire       [31:0]   _zz_18785;
  wire       [23:0]   _zz_18786;
  wire       [31:0]   _zz_18787;
  wire       [15:0]   _zz_18788;
  wire       [15:0]   _zz_18789;
  wire       [31:0]   _zz_18790;
  wire       [31:0]   _zz_18791;
  wire       [15:0]   _zz_18792;
  wire       [31:0]   _zz_18793;
  wire       [31:0]   _zz_18794;
  wire       [31:0]   _zz_18795;
  wire       [15:0]   _zz_18796;
  wire       [31:0]   _zz_18797;
  wire       [31:0]   _zz_18798;
  wire       [31:0]   _zz_18799;
  wire       [31:0]   _zz_18800;
  wire       [31:0]   _zz_18801;
  wire       [31:0]   _zz_18802;
  wire       [23:0]   _zz_18803;
  wire       [31:0]   _zz_18804;
  wire       [15:0]   _zz_18805;
  wire       [31:0]   _zz_18806;
  wire       [31:0]   _zz_18807;
  wire       [31:0]   _zz_18808;
  wire       [31:0]   _zz_18809;
  wire       [31:0]   _zz_18810;
  wire       [23:0]   _zz_18811;
  wire       [31:0]   _zz_18812;
  wire       [15:0]   _zz_18813;
  wire       [31:0]   _zz_18814;
  wire       [31:0]   _zz_18815;
  wire       [31:0]   _zz_18816;
  wire       [31:0]   _zz_18817;
  wire       [31:0]   _zz_18818;
  wire       [23:0]   _zz_18819;
  wire       [31:0]   _zz_18820;
  wire       [15:0]   _zz_18821;
  wire       [31:0]   _zz_18822;
  wire       [31:0]   _zz_18823;
  wire       [31:0]   _zz_18824;
  wire       [31:0]   _zz_18825;
  wire       [31:0]   _zz_18826;
  wire       [23:0]   _zz_18827;
  wire       [31:0]   _zz_18828;
  wire       [15:0]   _zz_18829;
  wire       [15:0]   _zz_18830;
  wire       [31:0]   _zz_18831;
  wire       [31:0]   _zz_18832;
  wire       [15:0]   _zz_18833;
  wire       [31:0]   _zz_18834;
  wire       [31:0]   _zz_18835;
  wire       [31:0]   _zz_18836;
  wire       [15:0]   _zz_18837;
  wire       [31:0]   _zz_18838;
  wire       [31:0]   _zz_18839;
  wire       [31:0]   _zz_18840;
  wire       [31:0]   _zz_18841;
  wire       [31:0]   _zz_18842;
  wire       [31:0]   _zz_18843;
  wire       [23:0]   _zz_18844;
  wire       [31:0]   _zz_18845;
  wire       [15:0]   _zz_18846;
  wire       [31:0]   _zz_18847;
  wire       [31:0]   _zz_18848;
  wire       [31:0]   _zz_18849;
  wire       [31:0]   _zz_18850;
  wire       [31:0]   _zz_18851;
  wire       [23:0]   _zz_18852;
  wire       [31:0]   _zz_18853;
  wire       [15:0]   _zz_18854;
  wire       [31:0]   _zz_18855;
  wire       [31:0]   _zz_18856;
  wire       [31:0]   _zz_18857;
  wire       [31:0]   _zz_18858;
  wire       [31:0]   _zz_18859;
  wire       [23:0]   _zz_18860;
  wire       [31:0]   _zz_18861;
  wire       [15:0]   _zz_18862;
  wire       [31:0]   _zz_18863;
  wire       [31:0]   _zz_18864;
  wire       [31:0]   _zz_18865;
  wire       [31:0]   _zz_18866;
  wire       [31:0]   _zz_18867;
  wire       [23:0]   _zz_18868;
  wire       [31:0]   _zz_18869;
  wire       [15:0]   _zz_18870;
  wire       [15:0]   _zz_18871;
  wire       [31:0]   _zz_18872;
  wire       [31:0]   _zz_18873;
  wire       [15:0]   _zz_18874;
  wire       [31:0]   _zz_18875;
  wire       [31:0]   _zz_18876;
  wire       [31:0]   _zz_18877;
  wire       [15:0]   _zz_18878;
  wire       [31:0]   _zz_18879;
  wire       [31:0]   _zz_18880;
  wire       [31:0]   _zz_18881;
  wire       [31:0]   _zz_18882;
  wire       [31:0]   _zz_18883;
  wire       [31:0]   _zz_18884;
  wire       [23:0]   _zz_18885;
  wire       [31:0]   _zz_18886;
  wire       [15:0]   _zz_18887;
  wire       [31:0]   _zz_18888;
  wire       [31:0]   _zz_18889;
  wire       [31:0]   _zz_18890;
  wire       [31:0]   _zz_18891;
  wire       [31:0]   _zz_18892;
  wire       [23:0]   _zz_18893;
  wire       [31:0]   _zz_18894;
  wire       [15:0]   _zz_18895;
  wire       [31:0]   _zz_18896;
  wire       [31:0]   _zz_18897;
  wire       [31:0]   _zz_18898;
  wire       [31:0]   _zz_18899;
  wire       [31:0]   _zz_18900;
  wire       [23:0]   _zz_18901;
  wire       [31:0]   _zz_18902;
  wire       [15:0]   _zz_18903;
  wire       [31:0]   _zz_18904;
  wire       [31:0]   _zz_18905;
  wire       [31:0]   _zz_18906;
  wire       [31:0]   _zz_18907;
  wire       [31:0]   _zz_18908;
  wire       [23:0]   _zz_18909;
  wire       [31:0]   _zz_18910;
  wire       [15:0]   _zz_18911;
  wire       [15:0]   _zz_18912;
  wire       [31:0]   _zz_18913;
  wire       [31:0]   _zz_18914;
  wire       [15:0]   _zz_18915;
  wire       [31:0]   _zz_18916;
  wire       [31:0]   _zz_18917;
  wire       [31:0]   _zz_18918;
  wire       [15:0]   _zz_18919;
  wire       [31:0]   _zz_18920;
  wire       [31:0]   _zz_18921;
  wire       [31:0]   _zz_18922;
  wire       [31:0]   _zz_18923;
  wire       [31:0]   _zz_18924;
  wire       [31:0]   _zz_18925;
  wire       [23:0]   _zz_18926;
  wire       [31:0]   _zz_18927;
  wire       [15:0]   _zz_18928;
  wire       [31:0]   _zz_18929;
  wire       [31:0]   _zz_18930;
  wire       [31:0]   _zz_18931;
  wire       [31:0]   _zz_18932;
  wire       [31:0]   _zz_18933;
  wire       [23:0]   _zz_18934;
  wire       [31:0]   _zz_18935;
  wire       [15:0]   _zz_18936;
  wire       [31:0]   _zz_18937;
  wire       [31:0]   _zz_18938;
  wire       [31:0]   _zz_18939;
  wire       [31:0]   _zz_18940;
  wire       [31:0]   _zz_18941;
  wire       [23:0]   _zz_18942;
  wire       [31:0]   _zz_18943;
  wire       [15:0]   _zz_18944;
  wire       [31:0]   _zz_18945;
  wire       [31:0]   _zz_18946;
  wire       [31:0]   _zz_18947;
  wire       [31:0]   _zz_18948;
  wire       [31:0]   _zz_18949;
  wire       [23:0]   _zz_18950;
  wire       [31:0]   _zz_18951;
  wire       [15:0]   _zz_18952;
  wire       [15:0]   _zz_18953;
  wire       [31:0]   _zz_18954;
  wire       [31:0]   _zz_18955;
  wire       [15:0]   _zz_18956;
  wire       [31:0]   _zz_18957;
  wire       [31:0]   _zz_18958;
  wire       [31:0]   _zz_18959;
  wire       [15:0]   _zz_18960;
  wire       [31:0]   _zz_18961;
  wire       [31:0]   _zz_18962;
  wire       [31:0]   _zz_18963;
  wire       [31:0]   _zz_18964;
  wire       [31:0]   _zz_18965;
  wire       [31:0]   _zz_18966;
  wire       [23:0]   _zz_18967;
  wire       [31:0]   _zz_18968;
  wire       [15:0]   _zz_18969;
  wire       [31:0]   _zz_18970;
  wire       [31:0]   _zz_18971;
  wire       [31:0]   _zz_18972;
  wire       [31:0]   _zz_18973;
  wire       [31:0]   _zz_18974;
  wire       [23:0]   _zz_18975;
  wire       [31:0]   _zz_18976;
  wire       [15:0]   _zz_18977;
  wire       [31:0]   _zz_18978;
  wire       [31:0]   _zz_18979;
  wire       [31:0]   _zz_18980;
  wire       [31:0]   _zz_18981;
  wire       [31:0]   _zz_18982;
  wire       [23:0]   _zz_18983;
  wire       [31:0]   _zz_18984;
  wire       [15:0]   _zz_18985;
  wire       [31:0]   _zz_18986;
  wire       [31:0]   _zz_18987;
  wire       [31:0]   _zz_18988;
  wire       [31:0]   _zz_18989;
  wire       [31:0]   _zz_18990;
  wire       [23:0]   _zz_18991;
  wire       [31:0]   _zz_18992;
  wire       [15:0]   _zz_18993;
  wire       [15:0]   _zz_18994;
  wire       [31:0]   _zz_18995;
  wire       [31:0]   _zz_18996;
  wire       [15:0]   _zz_18997;
  wire       [31:0]   _zz_18998;
  wire       [31:0]   _zz_18999;
  wire       [31:0]   _zz_19000;
  wire       [15:0]   _zz_19001;
  wire       [31:0]   _zz_19002;
  wire       [31:0]   _zz_19003;
  wire       [31:0]   _zz_19004;
  wire       [31:0]   _zz_19005;
  wire       [31:0]   _zz_19006;
  wire       [31:0]   _zz_19007;
  wire       [23:0]   _zz_19008;
  wire       [31:0]   _zz_19009;
  wire       [15:0]   _zz_19010;
  wire       [31:0]   _zz_19011;
  wire       [31:0]   _zz_19012;
  wire       [31:0]   _zz_19013;
  wire       [31:0]   _zz_19014;
  wire       [31:0]   _zz_19015;
  wire       [23:0]   _zz_19016;
  wire       [31:0]   _zz_19017;
  wire       [15:0]   _zz_19018;
  wire       [31:0]   _zz_19019;
  wire       [31:0]   _zz_19020;
  wire       [31:0]   _zz_19021;
  wire       [31:0]   _zz_19022;
  wire       [31:0]   _zz_19023;
  wire       [23:0]   _zz_19024;
  wire       [31:0]   _zz_19025;
  wire       [15:0]   _zz_19026;
  wire       [31:0]   _zz_19027;
  wire       [31:0]   _zz_19028;
  wire       [31:0]   _zz_19029;
  wire       [31:0]   _zz_19030;
  wire       [31:0]   _zz_19031;
  wire       [23:0]   _zz_19032;
  wire       [31:0]   _zz_19033;
  wire       [15:0]   _zz_19034;
  wire       [15:0]   _zz_19035;
  wire       [31:0]   _zz_19036;
  wire       [31:0]   _zz_19037;
  wire       [15:0]   _zz_19038;
  wire       [31:0]   _zz_19039;
  wire       [31:0]   _zz_19040;
  wire       [31:0]   _zz_19041;
  wire       [15:0]   _zz_19042;
  wire       [31:0]   _zz_19043;
  wire       [31:0]   _zz_19044;
  wire       [31:0]   _zz_19045;
  wire       [31:0]   _zz_19046;
  wire       [31:0]   _zz_19047;
  wire       [31:0]   _zz_19048;
  wire       [23:0]   _zz_19049;
  wire       [31:0]   _zz_19050;
  wire       [15:0]   _zz_19051;
  wire       [31:0]   _zz_19052;
  wire       [31:0]   _zz_19053;
  wire       [31:0]   _zz_19054;
  wire       [31:0]   _zz_19055;
  wire       [31:0]   _zz_19056;
  wire       [23:0]   _zz_19057;
  wire       [31:0]   _zz_19058;
  wire       [15:0]   _zz_19059;
  wire       [31:0]   _zz_19060;
  wire       [31:0]   _zz_19061;
  wire       [31:0]   _zz_19062;
  wire       [31:0]   _zz_19063;
  wire       [31:0]   _zz_19064;
  wire       [23:0]   _zz_19065;
  wire       [31:0]   _zz_19066;
  wire       [15:0]   _zz_19067;
  wire       [31:0]   _zz_19068;
  wire       [31:0]   _zz_19069;
  wire       [31:0]   _zz_19070;
  wire       [31:0]   _zz_19071;
  wire       [31:0]   _zz_19072;
  wire       [23:0]   _zz_19073;
  wire       [31:0]   _zz_19074;
  wire       [15:0]   _zz_19075;
  wire       [15:0]   _zz_19076;
  wire       [31:0]   _zz_19077;
  wire       [31:0]   _zz_19078;
  wire       [15:0]   _zz_19079;
  wire       [31:0]   _zz_19080;
  wire       [31:0]   _zz_19081;
  wire       [31:0]   _zz_19082;
  wire       [15:0]   _zz_19083;
  wire       [31:0]   _zz_19084;
  wire       [31:0]   _zz_19085;
  wire       [31:0]   _zz_19086;
  wire       [31:0]   _zz_19087;
  wire       [31:0]   _zz_19088;
  wire       [31:0]   _zz_19089;
  wire       [23:0]   _zz_19090;
  wire       [31:0]   _zz_19091;
  wire       [15:0]   _zz_19092;
  wire       [31:0]   _zz_19093;
  wire       [31:0]   _zz_19094;
  wire       [31:0]   _zz_19095;
  wire       [31:0]   _zz_19096;
  wire       [31:0]   _zz_19097;
  wire       [23:0]   _zz_19098;
  wire       [31:0]   _zz_19099;
  wire       [15:0]   _zz_19100;
  wire       [31:0]   _zz_19101;
  wire       [31:0]   _zz_19102;
  wire       [31:0]   _zz_19103;
  wire       [31:0]   _zz_19104;
  wire       [31:0]   _zz_19105;
  wire       [23:0]   _zz_19106;
  wire       [31:0]   _zz_19107;
  wire       [15:0]   _zz_19108;
  wire       [31:0]   _zz_19109;
  wire       [31:0]   _zz_19110;
  wire       [31:0]   _zz_19111;
  wire       [31:0]   _zz_19112;
  wire       [31:0]   _zz_19113;
  wire       [23:0]   _zz_19114;
  wire       [31:0]   _zz_19115;
  wire       [15:0]   _zz_19116;
  wire       [15:0]   _zz_19117;
  wire       [31:0]   _zz_19118;
  wire       [31:0]   _zz_19119;
  wire       [15:0]   _zz_19120;
  wire       [31:0]   _zz_19121;
  wire       [31:0]   _zz_19122;
  wire       [31:0]   _zz_19123;
  wire       [15:0]   _zz_19124;
  wire       [31:0]   _zz_19125;
  wire       [31:0]   _zz_19126;
  wire       [31:0]   _zz_19127;
  wire       [31:0]   _zz_19128;
  wire       [31:0]   _zz_19129;
  wire       [31:0]   _zz_19130;
  wire       [23:0]   _zz_19131;
  wire       [31:0]   _zz_19132;
  wire       [15:0]   _zz_19133;
  wire       [31:0]   _zz_19134;
  wire       [31:0]   _zz_19135;
  wire       [31:0]   _zz_19136;
  wire       [31:0]   _zz_19137;
  wire       [31:0]   _zz_19138;
  wire       [23:0]   _zz_19139;
  wire       [31:0]   _zz_19140;
  wire       [15:0]   _zz_19141;
  wire       [31:0]   _zz_19142;
  wire       [31:0]   _zz_19143;
  wire       [31:0]   _zz_19144;
  wire       [31:0]   _zz_19145;
  wire       [31:0]   _zz_19146;
  wire       [23:0]   _zz_19147;
  wire       [31:0]   _zz_19148;
  wire       [15:0]   _zz_19149;
  wire       [31:0]   _zz_19150;
  wire       [31:0]   _zz_19151;
  wire       [31:0]   _zz_19152;
  wire       [31:0]   _zz_19153;
  wire       [31:0]   _zz_19154;
  wire       [23:0]   _zz_19155;
  wire       [31:0]   _zz_19156;
  wire       [15:0]   _zz_19157;
  wire       [15:0]   _zz_19158;
  wire       [31:0]   _zz_19159;
  wire       [31:0]   _zz_19160;
  wire       [15:0]   _zz_19161;
  wire       [31:0]   _zz_19162;
  wire       [31:0]   _zz_19163;
  wire       [31:0]   _zz_19164;
  wire       [15:0]   _zz_19165;
  wire       [31:0]   _zz_19166;
  wire       [31:0]   _zz_19167;
  wire       [31:0]   _zz_19168;
  wire       [31:0]   _zz_19169;
  wire       [31:0]   _zz_19170;
  wire       [31:0]   _zz_19171;
  wire       [23:0]   _zz_19172;
  wire       [31:0]   _zz_19173;
  wire       [15:0]   _zz_19174;
  wire       [31:0]   _zz_19175;
  wire       [31:0]   _zz_19176;
  wire       [31:0]   _zz_19177;
  wire       [31:0]   _zz_19178;
  wire       [31:0]   _zz_19179;
  wire       [23:0]   _zz_19180;
  wire       [31:0]   _zz_19181;
  wire       [15:0]   _zz_19182;
  wire       [31:0]   _zz_19183;
  wire       [31:0]   _zz_19184;
  wire       [31:0]   _zz_19185;
  wire       [31:0]   _zz_19186;
  wire       [31:0]   _zz_19187;
  wire       [23:0]   _zz_19188;
  wire       [31:0]   _zz_19189;
  wire       [15:0]   _zz_19190;
  wire       [31:0]   _zz_19191;
  wire       [31:0]   _zz_19192;
  wire       [31:0]   _zz_19193;
  wire       [31:0]   _zz_19194;
  wire       [31:0]   _zz_19195;
  wire       [23:0]   _zz_19196;
  wire       [31:0]   _zz_19197;
  wire       [15:0]   _zz_19198;
  wire       [15:0]   _zz_19199;
  wire       [31:0]   _zz_19200;
  wire       [31:0]   _zz_19201;
  wire       [15:0]   _zz_19202;
  wire       [31:0]   _zz_19203;
  wire       [31:0]   _zz_19204;
  wire       [31:0]   _zz_19205;
  wire       [15:0]   _zz_19206;
  wire       [31:0]   _zz_19207;
  wire       [31:0]   _zz_19208;
  wire       [31:0]   _zz_19209;
  wire       [31:0]   _zz_19210;
  wire       [31:0]   _zz_19211;
  wire       [31:0]   _zz_19212;
  wire       [23:0]   _zz_19213;
  wire       [31:0]   _zz_19214;
  wire       [15:0]   _zz_19215;
  wire       [31:0]   _zz_19216;
  wire       [31:0]   _zz_19217;
  wire       [31:0]   _zz_19218;
  wire       [31:0]   _zz_19219;
  wire       [31:0]   _zz_19220;
  wire       [23:0]   _zz_19221;
  wire       [31:0]   _zz_19222;
  wire       [15:0]   _zz_19223;
  wire       [31:0]   _zz_19224;
  wire       [31:0]   _zz_19225;
  wire       [31:0]   _zz_19226;
  wire       [31:0]   _zz_19227;
  wire       [31:0]   _zz_19228;
  wire       [23:0]   _zz_19229;
  wire       [31:0]   _zz_19230;
  wire       [15:0]   _zz_19231;
  wire       [31:0]   _zz_19232;
  wire       [31:0]   _zz_19233;
  wire       [31:0]   _zz_19234;
  wire       [31:0]   _zz_19235;
  wire       [31:0]   _zz_19236;
  wire       [23:0]   _zz_19237;
  wire       [31:0]   _zz_19238;
  wire       [15:0]   _zz_19239;
  wire       [15:0]   _zz_19240;
  wire       [31:0]   _zz_19241;
  wire       [31:0]   _zz_19242;
  wire       [15:0]   _zz_19243;
  wire       [31:0]   _zz_19244;
  wire       [31:0]   _zz_19245;
  wire       [31:0]   _zz_19246;
  wire       [15:0]   _zz_19247;
  wire       [31:0]   _zz_19248;
  wire       [31:0]   _zz_19249;
  wire       [31:0]   _zz_19250;
  wire       [31:0]   _zz_19251;
  wire       [31:0]   _zz_19252;
  wire       [31:0]   _zz_19253;
  wire       [23:0]   _zz_19254;
  wire       [31:0]   _zz_19255;
  wire       [15:0]   _zz_19256;
  wire       [31:0]   _zz_19257;
  wire       [31:0]   _zz_19258;
  wire       [31:0]   _zz_19259;
  wire       [31:0]   _zz_19260;
  wire       [31:0]   _zz_19261;
  wire       [23:0]   _zz_19262;
  wire       [31:0]   _zz_19263;
  wire       [15:0]   _zz_19264;
  wire       [31:0]   _zz_19265;
  wire       [31:0]   _zz_19266;
  wire       [31:0]   _zz_19267;
  wire       [31:0]   _zz_19268;
  wire       [31:0]   _zz_19269;
  wire       [23:0]   _zz_19270;
  wire       [31:0]   _zz_19271;
  wire       [15:0]   _zz_19272;
  wire       [31:0]   _zz_19273;
  wire       [31:0]   _zz_19274;
  wire       [31:0]   _zz_19275;
  wire       [31:0]   _zz_19276;
  wire       [31:0]   _zz_19277;
  wire       [23:0]   _zz_19278;
  wire       [31:0]   _zz_19279;
  wire       [15:0]   _zz_19280;
  wire       [15:0]   _zz_19281;
  wire       [31:0]   _zz_19282;
  wire       [31:0]   _zz_19283;
  wire       [15:0]   _zz_19284;
  wire       [31:0]   _zz_19285;
  wire       [31:0]   _zz_19286;
  wire       [31:0]   _zz_19287;
  wire       [15:0]   _zz_19288;
  wire       [31:0]   _zz_19289;
  wire       [31:0]   _zz_19290;
  wire       [31:0]   _zz_19291;
  wire       [31:0]   _zz_19292;
  wire       [31:0]   _zz_19293;
  wire       [31:0]   _zz_19294;
  wire       [23:0]   _zz_19295;
  wire       [31:0]   _zz_19296;
  wire       [15:0]   _zz_19297;
  wire       [31:0]   _zz_19298;
  wire       [31:0]   _zz_19299;
  wire       [31:0]   _zz_19300;
  wire       [31:0]   _zz_19301;
  wire       [31:0]   _zz_19302;
  wire       [23:0]   _zz_19303;
  wire       [31:0]   _zz_19304;
  wire       [15:0]   _zz_19305;
  wire       [31:0]   _zz_19306;
  wire       [31:0]   _zz_19307;
  wire       [31:0]   _zz_19308;
  wire       [31:0]   _zz_19309;
  wire       [31:0]   _zz_19310;
  wire       [23:0]   _zz_19311;
  wire       [31:0]   _zz_19312;
  wire       [15:0]   _zz_19313;
  wire       [31:0]   _zz_19314;
  wire       [31:0]   _zz_19315;
  wire       [31:0]   _zz_19316;
  wire       [31:0]   _zz_19317;
  wire       [31:0]   _zz_19318;
  wire       [23:0]   _zz_19319;
  wire       [31:0]   _zz_19320;
  wire       [15:0]   _zz_19321;
  wire       [15:0]   _zz_19322;
  wire       [31:0]   _zz_19323;
  wire       [31:0]   _zz_19324;
  wire       [15:0]   _zz_19325;
  wire       [31:0]   _zz_19326;
  wire       [31:0]   _zz_19327;
  wire       [31:0]   _zz_19328;
  wire       [15:0]   _zz_19329;
  wire       [31:0]   _zz_19330;
  wire       [31:0]   _zz_19331;
  wire       [31:0]   _zz_19332;
  wire       [31:0]   _zz_19333;
  wire       [31:0]   _zz_19334;
  wire       [31:0]   _zz_19335;
  wire       [23:0]   _zz_19336;
  wire       [31:0]   _zz_19337;
  wire       [15:0]   _zz_19338;
  wire       [31:0]   _zz_19339;
  wire       [31:0]   _zz_19340;
  wire       [31:0]   _zz_19341;
  wire       [31:0]   _zz_19342;
  wire       [31:0]   _zz_19343;
  wire       [23:0]   _zz_19344;
  wire       [31:0]   _zz_19345;
  wire       [15:0]   _zz_19346;
  wire       [31:0]   _zz_19347;
  wire       [31:0]   _zz_19348;
  wire       [31:0]   _zz_19349;
  wire       [31:0]   _zz_19350;
  wire       [31:0]   _zz_19351;
  wire       [23:0]   _zz_19352;
  wire       [31:0]   _zz_19353;
  wire       [15:0]   _zz_19354;
  wire       [31:0]   _zz_19355;
  wire       [31:0]   _zz_19356;
  wire       [31:0]   _zz_19357;
  wire       [31:0]   _zz_19358;
  wire       [31:0]   _zz_19359;
  wire       [23:0]   _zz_19360;
  wire       [31:0]   _zz_19361;
  wire       [15:0]   _zz_19362;
  wire       [15:0]   _zz_19363;
  wire       [31:0]   _zz_19364;
  wire       [31:0]   _zz_19365;
  wire       [15:0]   _zz_19366;
  wire       [31:0]   _zz_19367;
  wire       [31:0]   _zz_19368;
  wire       [31:0]   _zz_19369;
  wire       [15:0]   _zz_19370;
  wire       [31:0]   _zz_19371;
  wire       [31:0]   _zz_19372;
  wire       [31:0]   _zz_19373;
  wire       [31:0]   _zz_19374;
  wire       [31:0]   _zz_19375;
  wire       [31:0]   _zz_19376;
  wire       [23:0]   _zz_19377;
  wire       [31:0]   _zz_19378;
  wire       [15:0]   _zz_19379;
  wire       [31:0]   _zz_19380;
  wire       [31:0]   _zz_19381;
  wire       [31:0]   _zz_19382;
  wire       [31:0]   _zz_19383;
  wire       [31:0]   _zz_19384;
  wire       [23:0]   _zz_19385;
  wire       [31:0]   _zz_19386;
  wire       [15:0]   _zz_19387;
  wire       [31:0]   _zz_19388;
  wire       [31:0]   _zz_19389;
  wire       [31:0]   _zz_19390;
  wire       [31:0]   _zz_19391;
  wire       [31:0]   _zz_19392;
  wire       [23:0]   _zz_19393;
  wire       [31:0]   _zz_19394;
  wire       [15:0]   _zz_19395;
  wire       [31:0]   _zz_19396;
  wire       [31:0]   _zz_19397;
  wire       [31:0]   _zz_19398;
  wire       [31:0]   _zz_19399;
  wire       [31:0]   _zz_19400;
  wire       [23:0]   _zz_19401;
  wire       [31:0]   _zz_19402;
  wire       [15:0]   _zz_19403;
  wire       [15:0]   _zz_19404;
  wire       [31:0]   _zz_19405;
  wire       [31:0]   _zz_19406;
  wire       [15:0]   _zz_19407;
  wire       [31:0]   _zz_19408;
  wire       [31:0]   _zz_19409;
  wire       [31:0]   _zz_19410;
  wire       [15:0]   _zz_19411;
  wire       [31:0]   _zz_19412;
  wire       [31:0]   _zz_19413;
  wire       [31:0]   _zz_19414;
  wire       [31:0]   _zz_19415;
  wire       [31:0]   _zz_19416;
  wire       [31:0]   _zz_19417;
  wire       [23:0]   _zz_19418;
  wire       [31:0]   _zz_19419;
  wire       [15:0]   _zz_19420;
  wire       [31:0]   _zz_19421;
  wire       [31:0]   _zz_19422;
  wire       [31:0]   _zz_19423;
  wire       [31:0]   _zz_19424;
  wire       [31:0]   _zz_19425;
  wire       [23:0]   _zz_19426;
  wire       [31:0]   _zz_19427;
  wire       [15:0]   _zz_19428;
  wire       [31:0]   _zz_19429;
  wire       [31:0]   _zz_19430;
  wire       [31:0]   _zz_19431;
  wire       [31:0]   _zz_19432;
  wire       [31:0]   _zz_19433;
  wire       [23:0]   _zz_19434;
  wire       [31:0]   _zz_19435;
  wire       [15:0]   _zz_19436;
  wire       [31:0]   _zz_19437;
  wire       [31:0]   _zz_19438;
  wire       [31:0]   _zz_19439;
  wire       [31:0]   _zz_19440;
  wire       [31:0]   _zz_19441;
  wire       [23:0]   _zz_19442;
  wire       [31:0]   _zz_19443;
  wire       [15:0]   _zz_19444;
  wire       [15:0]   _zz_19445;
  wire       [31:0]   _zz_19446;
  wire       [31:0]   _zz_19447;
  wire       [15:0]   _zz_19448;
  wire       [31:0]   _zz_19449;
  wire       [31:0]   _zz_19450;
  wire       [31:0]   _zz_19451;
  wire       [15:0]   _zz_19452;
  wire       [31:0]   _zz_19453;
  wire       [31:0]   _zz_19454;
  wire       [31:0]   _zz_19455;
  wire       [31:0]   _zz_19456;
  wire       [31:0]   _zz_19457;
  wire       [31:0]   _zz_19458;
  wire       [23:0]   _zz_19459;
  wire       [31:0]   _zz_19460;
  wire       [15:0]   _zz_19461;
  wire       [31:0]   _zz_19462;
  wire       [31:0]   _zz_19463;
  wire       [31:0]   _zz_19464;
  wire       [31:0]   _zz_19465;
  wire       [31:0]   _zz_19466;
  wire       [23:0]   _zz_19467;
  wire       [31:0]   _zz_19468;
  wire       [15:0]   _zz_19469;
  wire       [31:0]   _zz_19470;
  wire       [31:0]   _zz_19471;
  wire       [31:0]   _zz_19472;
  wire       [31:0]   _zz_19473;
  wire       [31:0]   _zz_19474;
  wire       [23:0]   _zz_19475;
  wire       [31:0]   _zz_19476;
  wire       [15:0]   _zz_19477;
  wire       [31:0]   _zz_19478;
  wire       [31:0]   _zz_19479;
  wire       [31:0]   _zz_19480;
  wire       [31:0]   _zz_19481;
  wire       [31:0]   _zz_19482;
  wire       [23:0]   _zz_19483;
  wire       [31:0]   _zz_19484;
  wire       [15:0]   _zz_19485;
  wire       [15:0]   _zz_19486;
  wire       [31:0]   _zz_19487;
  wire       [31:0]   _zz_19488;
  wire       [15:0]   _zz_19489;
  wire       [31:0]   _zz_19490;
  wire       [31:0]   _zz_19491;
  wire       [31:0]   _zz_19492;
  wire       [15:0]   _zz_19493;
  wire       [31:0]   _zz_19494;
  wire       [31:0]   _zz_19495;
  wire       [31:0]   _zz_19496;
  wire       [31:0]   _zz_19497;
  wire       [31:0]   _zz_19498;
  wire       [31:0]   _zz_19499;
  wire       [23:0]   _zz_19500;
  wire       [31:0]   _zz_19501;
  wire       [15:0]   _zz_19502;
  wire       [31:0]   _zz_19503;
  wire       [31:0]   _zz_19504;
  wire       [31:0]   _zz_19505;
  wire       [31:0]   _zz_19506;
  wire       [31:0]   _zz_19507;
  wire       [23:0]   _zz_19508;
  wire       [31:0]   _zz_19509;
  wire       [15:0]   _zz_19510;
  wire       [31:0]   _zz_19511;
  wire       [31:0]   _zz_19512;
  wire       [31:0]   _zz_19513;
  wire       [31:0]   _zz_19514;
  wire       [31:0]   _zz_19515;
  wire       [23:0]   _zz_19516;
  wire       [31:0]   _zz_19517;
  wire       [15:0]   _zz_19518;
  wire       [31:0]   _zz_19519;
  wire       [31:0]   _zz_19520;
  wire       [31:0]   _zz_19521;
  wire       [31:0]   _zz_19522;
  wire       [31:0]   _zz_19523;
  wire       [23:0]   _zz_19524;
  wire       [31:0]   _zz_19525;
  wire       [15:0]   _zz_19526;
  wire       [15:0]   _zz_19527;
  wire       [31:0]   _zz_19528;
  wire       [31:0]   _zz_19529;
  wire       [15:0]   _zz_19530;
  wire       [31:0]   _zz_19531;
  wire       [31:0]   _zz_19532;
  wire       [31:0]   _zz_19533;
  wire       [15:0]   _zz_19534;
  wire       [31:0]   _zz_19535;
  wire       [31:0]   _zz_19536;
  wire       [31:0]   _zz_19537;
  wire       [31:0]   _zz_19538;
  wire       [31:0]   _zz_19539;
  wire       [31:0]   _zz_19540;
  wire       [23:0]   _zz_19541;
  wire       [31:0]   _zz_19542;
  wire       [15:0]   _zz_19543;
  wire       [31:0]   _zz_19544;
  wire       [31:0]   _zz_19545;
  wire       [31:0]   _zz_19546;
  wire       [31:0]   _zz_19547;
  wire       [31:0]   _zz_19548;
  wire       [23:0]   _zz_19549;
  wire       [31:0]   _zz_19550;
  wire       [15:0]   _zz_19551;
  wire       [31:0]   _zz_19552;
  wire       [31:0]   _zz_19553;
  wire       [31:0]   _zz_19554;
  wire       [31:0]   _zz_19555;
  wire       [31:0]   _zz_19556;
  wire       [23:0]   _zz_19557;
  wire       [31:0]   _zz_19558;
  wire       [15:0]   _zz_19559;
  wire       [31:0]   _zz_19560;
  wire       [31:0]   _zz_19561;
  wire       [31:0]   _zz_19562;
  wire       [31:0]   _zz_19563;
  wire       [31:0]   _zz_19564;
  wire       [23:0]   _zz_19565;
  wire       [31:0]   _zz_19566;
  wire       [15:0]   _zz_19567;
  wire       [15:0]   _zz_19568;
  wire       [31:0]   _zz_19569;
  wire       [31:0]   _zz_19570;
  wire       [15:0]   _zz_19571;
  wire       [31:0]   _zz_19572;
  wire       [31:0]   _zz_19573;
  wire       [31:0]   _zz_19574;
  wire       [15:0]   _zz_19575;
  wire       [31:0]   _zz_19576;
  wire       [31:0]   _zz_19577;
  wire       [31:0]   _zz_19578;
  wire       [31:0]   _zz_19579;
  wire       [31:0]   _zz_19580;
  wire       [31:0]   _zz_19581;
  wire       [23:0]   _zz_19582;
  wire       [31:0]   _zz_19583;
  wire       [15:0]   _zz_19584;
  wire       [31:0]   _zz_19585;
  wire       [31:0]   _zz_19586;
  wire       [31:0]   _zz_19587;
  wire       [31:0]   _zz_19588;
  wire       [31:0]   _zz_19589;
  wire       [23:0]   _zz_19590;
  wire       [31:0]   _zz_19591;
  wire       [15:0]   _zz_19592;
  wire       [31:0]   _zz_19593;
  wire       [31:0]   _zz_19594;
  wire       [31:0]   _zz_19595;
  wire       [31:0]   _zz_19596;
  wire       [31:0]   _zz_19597;
  wire       [23:0]   _zz_19598;
  wire       [31:0]   _zz_19599;
  wire       [15:0]   _zz_19600;
  wire       [31:0]   _zz_19601;
  wire       [31:0]   _zz_19602;
  wire       [31:0]   _zz_19603;
  wire       [31:0]   _zz_19604;
  wire       [31:0]   _zz_19605;
  wire       [23:0]   _zz_19606;
  wire       [31:0]   _zz_19607;
  wire       [15:0]   _zz_19608;
  wire       [15:0]   _zz_19609;
  wire       [31:0]   _zz_19610;
  wire       [31:0]   _zz_19611;
  wire       [15:0]   _zz_19612;
  wire       [31:0]   _zz_19613;
  wire       [31:0]   _zz_19614;
  wire       [31:0]   _zz_19615;
  wire       [15:0]   _zz_19616;
  wire       [31:0]   _zz_19617;
  wire       [31:0]   _zz_19618;
  wire       [31:0]   _zz_19619;
  wire       [31:0]   _zz_19620;
  wire       [31:0]   _zz_19621;
  wire       [31:0]   _zz_19622;
  wire       [23:0]   _zz_19623;
  wire       [31:0]   _zz_19624;
  wire       [15:0]   _zz_19625;
  wire       [31:0]   _zz_19626;
  wire       [31:0]   _zz_19627;
  wire       [31:0]   _zz_19628;
  wire       [31:0]   _zz_19629;
  wire       [31:0]   _zz_19630;
  wire       [23:0]   _zz_19631;
  wire       [31:0]   _zz_19632;
  wire       [15:0]   _zz_19633;
  wire       [31:0]   _zz_19634;
  wire       [31:0]   _zz_19635;
  wire       [31:0]   _zz_19636;
  wire       [31:0]   _zz_19637;
  wire       [31:0]   _zz_19638;
  wire       [23:0]   _zz_19639;
  wire       [31:0]   _zz_19640;
  wire       [15:0]   _zz_19641;
  wire       [31:0]   _zz_19642;
  wire       [31:0]   _zz_19643;
  wire       [31:0]   _zz_19644;
  wire       [31:0]   _zz_19645;
  wire       [31:0]   _zz_19646;
  wire       [23:0]   _zz_19647;
  wire       [31:0]   _zz_19648;
  wire       [15:0]   _zz_19649;
  wire       [15:0]   _zz_19650;
  wire       [31:0]   _zz_19651;
  wire       [31:0]   _zz_19652;
  wire       [15:0]   _zz_19653;
  wire       [31:0]   _zz_19654;
  wire       [31:0]   _zz_19655;
  wire       [31:0]   _zz_19656;
  wire       [15:0]   _zz_19657;
  wire       [31:0]   _zz_19658;
  wire       [31:0]   _zz_19659;
  wire       [31:0]   _zz_19660;
  wire       [31:0]   _zz_19661;
  wire       [31:0]   _zz_19662;
  wire       [31:0]   _zz_19663;
  wire       [23:0]   _zz_19664;
  wire       [31:0]   _zz_19665;
  wire       [15:0]   _zz_19666;
  wire       [31:0]   _zz_19667;
  wire       [31:0]   _zz_19668;
  wire       [31:0]   _zz_19669;
  wire       [31:0]   _zz_19670;
  wire       [31:0]   _zz_19671;
  wire       [23:0]   _zz_19672;
  wire       [31:0]   _zz_19673;
  wire       [15:0]   _zz_19674;
  wire       [31:0]   _zz_19675;
  wire       [31:0]   _zz_19676;
  wire       [31:0]   _zz_19677;
  wire       [31:0]   _zz_19678;
  wire       [31:0]   _zz_19679;
  wire       [23:0]   _zz_19680;
  wire       [31:0]   _zz_19681;
  wire       [15:0]   _zz_19682;
  wire       [31:0]   _zz_19683;
  wire       [31:0]   _zz_19684;
  wire       [31:0]   _zz_19685;
  wire       [31:0]   _zz_19686;
  wire       [31:0]   _zz_19687;
  wire       [23:0]   _zz_19688;
  wire       [31:0]   _zz_19689;
  wire       [15:0]   _zz_19690;
  wire       [15:0]   _zz_19691;
  wire       [31:0]   _zz_19692;
  wire       [31:0]   _zz_19693;
  wire       [15:0]   _zz_19694;
  wire       [31:0]   _zz_19695;
  wire       [31:0]   _zz_19696;
  wire       [31:0]   _zz_19697;
  wire       [15:0]   _zz_19698;
  wire       [31:0]   _zz_19699;
  wire       [31:0]   _zz_19700;
  wire       [31:0]   _zz_19701;
  wire       [31:0]   _zz_19702;
  wire       [31:0]   _zz_19703;
  wire       [31:0]   _zz_19704;
  wire       [23:0]   _zz_19705;
  wire       [31:0]   _zz_19706;
  wire       [15:0]   _zz_19707;
  wire       [31:0]   _zz_19708;
  wire       [31:0]   _zz_19709;
  wire       [31:0]   _zz_19710;
  wire       [31:0]   _zz_19711;
  wire       [31:0]   _zz_19712;
  wire       [23:0]   _zz_19713;
  wire       [31:0]   _zz_19714;
  wire       [15:0]   _zz_19715;
  wire       [31:0]   _zz_19716;
  wire       [31:0]   _zz_19717;
  wire       [31:0]   _zz_19718;
  wire       [31:0]   _zz_19719;
  wire       [31:0]   _zz_19720;
  wire       [23:0]   _zz_19721;
  wire       [31:0]   _zz_19722;
  wire       [15:0]   _zz_19723;
  wire       [31:0]   _zz_19724;
  wire       [31:0]   _zz_19725;
  wire       [31:0]   _zz_19726;
  wire       [31:0]   _zz_19727;
  wire       [31:0]   _zz_19728;
  wire       [23:0]   _zz_19729;
  wire       [31:0]   _zz_19730;
  wire       [15:0]   _zz_19731;
  wire       [15:0]   _zz_19732;
  wire       [31:0]   _zz_19733;
  wire       [31:0]   _zz_19734;
  wire       [15:0]   _zz_19735;
  wire       [31:0]   _zz_19736;
  wire       [31:0]   _zz_19737;
  wire       [31:0]   _zz_19738;
  wire       [15:0]   _zz_19739;
  wire       [31:0]   _zz_19740;
  wire       [31:0]   _zz_19741;
  wire       [31:0]   _zz_19742;
  wire       [31:0]   _zz_19743;
  wire       [31:0]   _zz_19744;
  wire       [31:0]   _zz_19745;
  wire       [23:0]   _zz_19746;
  wire       [31:0]   _zz_19747;
  wire       [15:0]   _zz_19748;
  wire       [31:0]   _zz_19749;
  wire       [31:0]   _zz_19750;
  wire       [31:0]   _zz_19751;
  wire       [31:0]   _zz_19752;
  wire       [31:0]   _zz_19753;
  wire       [23:0]   _zz_19754;
  wire       [31:0]   _zz_19755;
  wire       [15:0]   _zz_19756;
  wire       [31:0]   _zz_19757;
  wire       [31:0]   _zz_19758;
  wire       [31:0]   _zz_19759;
  wire       [31:0]   _zz_19760;
  wire       [31:0]   _zz_19761;
  wire       [23:0]   _zz_19762;
  wire       [31:0]   _zz_19763;
  wire       [15:0]   _zz_19764;
  wire       [31:0]   _zz_19765;
  wire       [31:0]   _zz_19766;
  wire       [31:0]   _zz_19767;
  wire       [31:0]   _zz_19768;
  wire       [31:0]   _zz_19769;
  wire       [23:0]   _zz_19770;
  wire       [31:0]   _zz_19771;
  wire       [15:0]   _zz_19772;
  wire       [15:0]   _zz_19773;
  wire       [31:0]   _zz_19774;
  wire       [31:0]   _zz_19775;
  wire       [15:0]   _zz_19776;
  wire       [31:0]   _zz_19777;
  wire       [31:0]   _zz_19778;
  wire       [31:0]   _zz_19779;
  wire       [15:0]   _zz_19780;
  wire       [31:0]   _zz_19781;
  wire       [31:0]   _zz_19782;
  wire       [31:0]   _zz_19783;
  wire       [31:0]   _zz_19784;
  wire       [31:0]   _zz_19785;
  wire       [31:0]   _zz_19786;
  wire       [23:0]   _zz_19787;
  wire       [31:0]   _zz_19788;
  wire       [15:0]   _zz_19789;
  wire       [31:0]   _zz_19790;
  wire       [31:0]   _zz_19791;
  wire       [31:0]   _zz_19792;
  wire       [31:0]   _zz_19793;
  wire       [31:0]   _zz_19794;
  wire       [23:0]   _zz_19795;
  wire       [31:0]   _zz_19796;
  wire       [15:0]   _zz_19797;
  wire       [31:0]   _zz_19798;
  wire       [31:0]   _zz_19799;
  wire       [31:0]   _zz_19800;
  wire       [31:0]   _zz_19801;
  wire       [31:0]   _zz_19802;
  wire       [23:0]   _zz_19803;
  wire       [31:0]   _zz_19804;
  wire       [15:0]   _zz_19805;
  wire       [31:0]   _zz_19806;
  wire       [31:0]   _zz_19807;
  wire       [31:0]   _zz_19808;
  wire       [31:0]   _zz_19809;
  wire       [31:0]   _zz_19810;
  wire       [23:0]   _zz_19811;
  wire       [31:0]   _zz_19812;
  wire       [15:0]   _zz_19813;
  wire       [15:0]   _zz_19814;
  wire       [31:0]   _zz_19815;
  wire       [31:0]   _zz_19816;
  wire       [15:0]   _zz_19817;
  wire       [31:0]   _zz_19818;
  wire       [31:0]   _zz_19819;
  wire       [31:0]   _zz_19820;
  wire       [15:0]   _zz_19821;
  wire       [31:0]   _zz_19822;
  wire       [31:0]   _zz_19823;
  wire       [31:0]   _zz_19824;
  wire       [31:0]   _zz_19825;
  wire       [31:0]   _zz_19826;
  wire       [31:0]   _zz_19827;
  wire       [23:0]   _zz_19828;
  wire       [31:0]   _zz_19829;
  wire       [15:0]   _zz_19830;
  wire       [31:0]   _zz_19831;
  wire       [31:0]   _zz_19832;
  wire       [31:0]   _zz_19833;
  wire       [31:0]   _zz_19834;
  wire       [31:0]   _zz_19835;
  wire       [23:0]   _zz_19836;
  wire       [31:0]   _zz_19837;
  wire       [15:0]   _zz_19838;
  wire       [31:0]   _zz_19839;
  wire       [31:0]   _zz_19840;
  wire       [31:0]   _zz_19841;
  wire       [31:0]   _zz_19842;
  wire       [31:0]   _zz_19843;
  wire       [23:0]   _zz_19844;
  wire       [31:0]   _zz_19845;
  wire       [15:0]   _zz_19846;
  wire       [31:0]   _zz_19847;
  wire       [31:0]   _zz_19848;
  wire       [31:0]   _zz_19849;
  wire       [31:0]   _zz_19850;
  wire       [31:0]   _zz_19851;
  wire       [23:0]   _zz_19852;
  wire       [31:0]   _zz_19853;
  wire       [15:0]   _zz_19854;
  wire       [15:0]   _zz_19855;
  wire       [31:0]   _zz_19856;
  wire       [31:0]   _zz_19857;
  wire       [15:0]   _zz_19858;
  wire       [31:0]   _zz_19859;
  wire       [31:0]   _zz_19860;
  wire       [31:0]   _zz_19861;
  wire       [15:0]   _zz_19862;
  wire       [31:0]   _zz_19863;
  wire       [31:0]   _zz_19864;
  wire       [31:0]   _zz_19865;
  wire       [31:0]   _zz_19866;
  wire       [31:0]   _zz_19867;
  wire       [31:0]   _zz_19868;
  wire       [23:0]   _zz_19869;
  wire       [31:0]   _zz_19870;
  wire       [15:0]   _zz_19871;
  wire       [31:0]   _zz_19872;
  wire       [31:0]   _zz_19873;
  wire       [31:0]   _zz_19874;
  wire       [31:0]   _zz_19875;
  wire       [31:0]   _zz_19876;
  wire       [23:0]   _zz_19877;
  wire       [31:0]   _zz_19878;
  wire       [15:0]   _zz_19879;
  wire       [31:0]   _zz_19880;
  wire       [31:0]   _zz_19881;
  wire       [31:0]   _zz_19882;
  wire       [31:0]   _zz_19883;
  wire       [31:0]   _zz_19884;
  wire       [23:0]   _zz_19885;
  wire       [31:0]   _zz_19886;
  wire       [15:0]   _zz_19887;
  wire       [31:0]   _zz_19888;
  wire       [31:0]   _zz_19889;
  wire       [31:0]   _zz_19890;
  wire       [31:0]   _zz_19891;
  wire       [31:0]   _zz_19892;
  wire       [23:0]   _zz_19893;
  wire       [31:0]   _zz_19894;
  wire       [15:0]   _zz_19895;
  wire       [15:0]   _zz_19896;
  wire       [31:0]   _zz_19897;
  wire       [31:0]   _zz_19898;
  wire       [15:0]   _zz_19899;
  wire       [31:0]   _zz_19900;
  wire       [31:0]   _zz_19901;
  wire       [31:0]   _zz_19902;
  wire       [15:0]   _zz_19903;
  wire       [31:0]   _zz_19904;
  wire       [31:0]   _zz_19905;
  wire       [31:0]   _zz_19906;
  wire       [31:0]   _zz_19907;
  wire       [31:0]   _zz_19908;
  wire       [31:0]   _zz_19909;
  wire       [23:0]   _zz_19910;
  wire       [31:0]   _zz_19911;
  wire       [15:0]   _zz_19912;
  wire       [31:0]   _zz_19913;
  wire       [31:0]   _zz_19914;
  wire       [31:0]   _zz_19915;
  wire       [31:0]   _zz_19916;
  wire       [31:0]   _zz_19917;
  wire       [23:0]   _zz_19918;
  wire       [31:0]   _zz_19919;
  wire       [15:0]   _zz_19920;
  wire       [31:0]   _zz_19921;
  wire       [31:0]   _zz_19922;
  wire       [31:0]   _zz_19923;
  wire       [31:0]   _zz_19924;
  wire       [31:0]   _zz_19925;
  wire       [23:0]   _zz_19926;
  wire       [31:0]   _zz_19927;
  wire       [15:0]   _zz_19928;
  wire       [31:0]   _zz_19929;
  wire       [31:0]   _zz_19930;
  wire       [31:0]   _zz_19931;
  wire       [31:0]   _zz_19932;
  wire       [31:0]   _zz_19933;
  wire       [23:0]   _zz_19934;
  wire       [31:0]   _zz_19935;
  wire       [15:0]   _zz_19936;
  wire       [15:0]   _zz_19937;
  wire       [31:0]   _zz_19938;
  wire       [31:0]   _zz_19939;
  wire       [15:0]   _zz_19940;
  wire       [31:0]   _zz_19941;
  wire       [31:0]   _zz_19942;
  wire       [31:0]   _zz_19943;
  wire       [15:0]   _zz_19944;
  wire       [31:0]   _zz_19945;
  wire       [31:0]   _zz_19946;
  wire       [31:0]   _zz_19947;
  wire       [31:0]   _zz_19948;
  wire       [31:0]   _zz_19949;
  wire       [31:0]   _zz_19950;
  wire       [23:0]   _zz_19951;
  wire       [31:0]   _zz_19952;
  wire       [15:0]   _zz_19953;
  wire       [31:0]   _zz_19954;
  wire       [31:0]   _zz_19955;
  wire       [31:0]   _zz_19956;
  wire       [31:0]   _zz_19957;
  wire       [31:0]   _zz_19958;
  wire       [23:0]   _zz_19959;
  wire       [31:0]   _zz_19960;
  wire       [15:0]   _zz_19961;
  wire       [31:0]   _zz_19962;
  wire       [31:0]   _zz_19963;
  wire       [31:0]   _zz_19964;
  wire       [31:0]   _zz_19965;
  wire       [31:0]   _zz_19966;
  wire       [23:0]   _zz_19967;
  wire       [31:0]   _zz_19968;
  wire       [15:0]   _zz_19969;
  wire       [31:0]   _zz_19970;
  wire       [31:0]   _zz_19971;
  wire       [31:0]   _zz_19972;
  wire       [31:0]   _zz_19973;
  wire       [31:0]   _zz_19974;
  wire       [23:0]   _zz_19975;
  wire       [31:0]   _zz_19976;
  wire       [15:0]   _zz_19977;
  wire       [15:0]   _zz_19978;
  wire       [31:0]   _zz_19979;
  wire       [31:0]   _zz_19980;
  wire       [15:0]   _zz_19981;
  wire       [31:0]   _zz_19982;
  wire       [31:0]   _zz_19983;
  wire       [31:0]   _zz_19984;
  wire       [15:0]   _zz_19985;
  wire       [31:0]   _zz_19986;
  wire       [31:0]   _zz_19987;
  wire       [31:0]   _zz_19988;
  wire       [31:0]   _zz_19989;
  wire       [31:0]   _zz_19990;
  wire       [31:0]   _zz_19991;
  wire       [23:0]   _zz_19992;
  wire       [31:0]   _zz_19993;
  wire       [15:0]   _zz_19994;
  wire       [31:0]   _zz_19995;
  wire       [31:0]   _zz_19996;
  wire       [31:0]   _zz_19997;
  wire       [31:0]   _zz_19998;
  wire       [31:0]   _zz_19999;
  wire       [23:0]   _zz_20000;
  wire       [31:0]   _zz_20001;
  wire       [15:0]   _zz_20002;
  wire       [31:0]   _zz_20003;
  wire       [31:0]   _zz_20004;
  wire       [31:0]   _zz_20005;
  wire       [31:0]   _zz_20006;
  wire       [31:0]   _zz_20007;
  wire       [23:0]   _zz_20008;
  wire       [31:0]   _zz_20009;
  wire       [15:0]   _zz_20010;
  wire       [31:0]   _zz_20011;
  wire       [31:0]   _zz_20012;
  wire       [31:0]   _zz_20013;
  wire       [31:0]   _zz_20014;
  wire       [31:0]   _zz_20015;
  wire       [23:0]   _zz_20016;
  wire       [31:0]   _zz_20017;
  wire       [15:0]   _zz_20018;
  wire       [15:0]   _zz_20019;
  wire       [31:0]   _zz_20020;
  wire       [31:0]   _zz_20021;
  wire       [15:0]   _zz_20022;
  wire       [31:0]   _zz_20023;
  wire       [31:0]   _zz_20024;
  wire       [31:0]   _zz_20025;
  wire       [15:0]   _zz_20026;
  wire       [31:0]   _zz_20027;
  wire       [31:0]   _zz_20028;
  wire       [31:0]   _zz_20029;
  wire       [31:0]   _zz_20030;
  wire       [31:0]   _zz_20031;
  wire       [31:0]   _zz_20032;
  wire       [23:0]   _zz_20033;
  wire       [31:0]   _zz_20034;
  wire       [15:0]   _zz_20035;
  wire       [31:0]   _zz_20036;
  wire       [31:0]   _zz_20037;
  wire       [31:0]   _zz_20038;
  wire       [31:0]   _zz_20039;
  wire       [31:0]   _zz_20040;
  wire       [23:0]   _zz_20041;
  wire       [31:0]   _zz_20042;
  wire       [15:0]   _zz_20043;
  wire       [31:0]   _zz_20044;
  wire       [31:0]   _zz_20045;
  wire       [31:0]   _zz_20046;
  wire       [31:0]   _zz_20047;
  wire       [31:0]   _zz_20048;
  wire       [23:0]   _zz_20049;
  wire       [31:0]   _zz_20050;
  wire       [15:0]   _zz_20051;
  wire       [31:0]   _zz_20052;
  wire       [31:0]   _zz_20053;
  wire       [31:0]   _zz_20054;
  wire       [31:0]   _zz_20055;
  wire       [31:0]   _zz_20056;
  wire       [23:0]   _zz_20057;
  wire       [31:0]   _zz_20058;
  wire       [15:0]   _zz_20059;
  wire       [15:0]   _zz_20060;
  wire       [31:0]   _zz_20061;
  wire       [31:0]   _zz_20062;
  wire       [15:0]   _zz_20063;
  wire       [31:0]   _zz_20064;
  wire       [31:0]   _zz_20065;
  wire       [31:0]   _zz_20066;
  wire       [15:0]   _zz_20067;
  wire       [31:0]   _zz_20068;
  wire       [31:0]   _zz_20069;
  wire       [31:0]   _zz_20070;
  wire       [31:0]   _zz_20071;
  wire       [31:0]   _zz_20072;
  wire       [31:0]   _zz_20073;
  wire       [23:0]   _zz_20074;
  wire       [31:0]   _zz_20075;
  wire       [15:0]   _zz_20076;
  wire       [31:0]   _zz_20077;
  wire       [31:0]   _zz_20078;
  wire       [31:0]   _zz_20079;
  wire       [31:0]   _zz_20080;
  wire       [31:0]   _zz_20081;
  wire       [23:0]   _zz_20082;
  wire       [31:0]   _zz_20083;
  wire       [15:0]   _zz_20084;
  wire       [31:0]   _zz_20085;
  wire       [31:0]   _zz_20086;
  wire       [31:0]   _zz_20087;
  wire       [31:0]   _zz_20088;
  wire       [31:0]   _zz_20089;
  wire       [23:0]   _zz_20090;
  wire       [31:0]   _zz_20091;
  wire       [15:0]   _zz_20092;
  wire       [31:0]   _zz_20093;
  wire       [31:0]   _zz_20094;
  wire       [31:0]   _zz_20095;
  wire       [31:0]   _zz_20096;
  wire       [31:0]   _zz_20097;
  wire       [23:0]   _zz_20098;
  wire       [31:0]   _zz_20099;
  wire       [15:0]   _zz_20100;
  wire       [15:0]   _zz_20101;
  wire       [31:0]   _zz_20102;
  wire       [31:0]   _zz_20103;
  wire       [15:0]   _zz_20104;
  wire       [31:0]   _zz_20105;
  wire       [31:0]   _zz_20106;
  wire       [31:0]   _zz_20107;
  wire       [15:0]   _zz_20108;
  wire       [31:0]   _zz_20109;
  wire       [31:0]   _zz_20110;
  wire       [31:0]   _zz_20111;
  wire       [31:0]   _zz_20112;
  wire       [31:0]   _zz_20113;
  wire       [31:0]   _zz_20114;
  wire       [23:0]   _zz_20115;
  wire       [31:0]   _zz_20116;
  wire       [15:0]   _zz_20117;
  wire       [31:0]   _zz_20118;
  wire       [31:0]   _zz_20119;
  wire       [31:0]   _zz_20120;
  wire       [31:0]   _zz_20121;
  wire       [31:0]   _zz_20122;
  wire       [23:0]   _zz_20123;
  wire       [31:0]   _zz_20124;
  wire       [15:0]   _zz_20125;
  wire       [31:0]   _zz_20126;
  wire       [31:0]   _zz_20127;
  wire       [31:0]   _zz_20128;
  wire       [31:0]   _zz_20129;
  wire       [31:0]   _zz_20130;
  wire       [23:0]   _zz_20131;
  wire       [31:0]   _zz_20132;
  wire       [15:0]   _zz_20133;
  wire       [31:0]   _zz_20134;
  wire       [31:0]   _zz_20135;
  wire       [31:0]   _zz_20136;
  wire       [31:0]   _zz_20137;
  wire       [31:0]   _zz_20138;
  wire       [23:0]   _zz_20139;
  wire       [31:0]   _zz_20140;
  wire       [15:0]   _zz_20141;
  wire       [15:0]   _zz_20142;
  wire       [31:0]   _zz_20143;
  wire       [31:0]   _zz_20144;
  wire       [15:0]   _zz_20145;
  wire       [31:0]   _zz_20146;
  wire       [31:0]   _zz_20147;
  wire       [31:0]   _zz_20148;
  wire       [15:0]   _zz_20149;
  wire       [31:0]   _zz_20150;
  wire       [31:0]   _zz_20151;
  wire       [31:0]   _zz_20152;
  wire       [31:0]   _zz_20153;
  wire       [31:0]   _zz_20154;
  wire       [31:0]   _zz_20155;
  wire       [23:0]   _zz_20156;
  wire       [31:0]   _zz_20157;
  wire       [15:0]   _zz_20158;
  wire       [31:0]   _zz_20159;
  wire       [31:0]   _zz_20160;
  wire       [31:0]   _zz_20161;
  wire       [31:0]   _zz_20162;
  wire       [31:0]   _zz_20163;
  wire       [23:0]   _zz_20164;
  wire       [31:0]   _zz_20165;
  wire       [15:0]   _zz_20166;
  wire       [31:0]   _zz_20167;
  wire       [31:0]   _zz_20168;
  wire       [31:0]   _zz_20169;
  wire       [31:0]   _zz_20170;
  wire       [31:0]   _zz_20171;
  wire       [23:0]   _zz_20172;
  wire       [31:0]   _zz_20173;
  wire       [15:0]   _zz_20174;
  wire       [31:0]   _zz_20175;
  wire       [31:0]   _zz_20176;
  wire       [31:0]   _zz_20177;
  wire       [31:0]   _zz_20178;
  wire       [31:0]   _zz_20179;
  wire       [23:0]   _zz_20180;
  wire       [31:0]   _zz_20181;
  wire       [15:0]   _zz_20182;
  wire       [15:0]   _zz_20183;
  wire       [31:0]   _zz_20184;
  wire       [31:0]   _zz_20185;
  wire       [15:0]   _zz_20186;
  wire       [31:0]   _zz_20187;
  wire       [31:0]   _zz_20188;
  wire       [31:0]   _zz_20189;
  wire       [15:0]   _zz_20190;
  wire       [31:0]   _zz_20191;
  wire       [31:0]   _zz_20192;
  wire       [31:0]   _zz_20193;
  wire       [31:0]   _zz_20194;
  wire       [31:0]   _zz_20195;
  wire       [31:0]   _zz_20196;
  wire       [23:0]   _zz_20197;
  wire       [31:0]   _zz_20198;
  wire       [15:0]   _zz_20199;
  wire       [31:0]   _zz_20200;
  wire       [31:0]   _zz_20201;
  wire       [31:0]   _zz_20202;
  wire       [31:0]   _zz_20203;
  wire       [31:0]   _zz_20204;
  wire       [23:0]   _zz_20205;
  wire       [31:0]   _zz_20206;
  wire       [15:0]   _zz_20207;
  wire       [31:0]   _zz_20208;
  wire       [31:0]   _zz_20209;
  wire       [31:0]   _zz_20210;
  wire       [31:0]   _zz_20211;
  wire       [31:0]   _zz_20212;
  wire       [23:0]   _zz_20213;
  wire       [31:0]   _zz_20214;
  wire       [15:0]   _zz_20215;
  wire       [31:0]   _zz_20216;
  wire       [31:0]   _zz_20217;
  wire       [31:0]   _zz_20218;
  wire       [31:0]   _zz_20219;
  wire       [31:0]   _zz_20220;
  wire       [23:0]   _zz_20221;
  wire       [31:0]   _zz_20222;
  wire       [15:0]   _zz_20223;
  wire       [15:0]   _zz_20224;
  wire       [31:0]   _zz_20225;
  wire       [31:0]   _zz_20226;
  wire       [15:0]   _zz_20227;
  wire       [31:0]   _zz_20228;
  wire       [31:0]   _zz_20229;
  wire       [31:0]   _zz_20230;
  wire       [15:0]   _zz_20231;
  wire       [31:0]   _zz_20232;
  wire       [31:0]   _zz_20233;
  wire       [31:0]   _zz_20234;
  wire       [31:0]   _zz_20235;
  wire       [31:0]   _zz_20236;
  wire       [31:0]   _zz_20237;
  wire       [23:0]   _zz_20238;
  wire       [31:0]   _zz_20239;
  wire       [15:0]   _zz_20240;
  wire       [31:0]   _zz_20241;
  wire       [31:0]   _zz_20242;
  wire       [31:0]   _zz_20243;
  wire       [31:0]   _zz_20244;
  wire       [31:0]   _zz_20245;
  wire       [23:0]   _zz_20246;
  wire       [31:0]   _zz_20247;
  wire       [15:0]   _zz_20248;
  wire       [31:0]   _zz_20249;
  wire       [31:0]   _zz_20250;
  wire       [31:0]   _zz_20251;
  wire       [31:0]   _zz_20252;
  wire       [31:0]   _zz_20253;
  wire       [23:0]   _zz_20254;
  wire       [31:0]   _zz_20255;
  wire       [15:0]   _zz_20256;
  wire       [31:0]   _zz_20257;
  wire       [31:0]   _zz_20258;
  wire       [31:0]   _zz_20259;
  wire       [31:0]   _zz_20260;
  wire       [31:0]   _zz_20261;
  wire       [23:0]   _zz_20262;
  wire       [31:0]   _zz_20263;
  wire       [15:0]   _zz_20264;
  wire       [15:0]   _zz_20265;
  wire       [31:0]   _zz_20266;
  wire       [31:0]   _zz_20267;
  wire       [15:0]   _zz_20268;
  wire       [31:0]   _zz_20269;
  wire       [31:0]   _zz_20270;
  wire       [31:0]   _zz_20271;
  wire       [15:0]   _zz_20272;
  wire       [31:0]   _zz_20273;
  wire       [31:0]   _zz_20274;
  wire       [31:0]   _zz_20275;
  wire       [31:0]   _zz_20276;
  wire       [31:0]   _zz_20277;
  wire       [31:0]   _zz_20278;
  wire       [23:0]   _zz_20279;
  wire       [31:0]   _zz_20280;
  wire       [15:0]   _zz_20281;
  wire       [31:0]   _zz_20282;
  wire       [31:0]   _zz_20283;
  wire       [31:0]   _zz_20284;
  wire       [31:0]   _zz_20285;
  wire       [31:0]   _zz_20286;
  wire       [23:0]   _zz_20287;
  wire       [31:0]   _zz_20288;
  wire       [15:0]   _zz_20289;
  wire       [31:0]   _zz_20290;
  wire       [31:0]   _zz_20291;
  wire       [31:0]   _zz_20292;
  wire       [31:0]   _zz_20293;
  wire       [31:0]   _zz_20294;
  wire       [23:0]   _zz_20295;
  wire       [31:0]   _zz_20296;
  wire       [15:0]   _zz_20297;
  wire       [31:0]   _zz_20298;
  wire       [31:0]   _zz_20299;
  wire       [31:0]   _zz_20300;
  wire       [31:0]   _zz_20301;
  wire       [31:0]   _zz_20302;
  wire       [23:0]   _zz_20303;
  wire       [31:0]   _zz_20304;
  wire       [15:0]   _zz_20305;
  wire       [15:0]   _zz_20306;
  wire       [31:0]   _zz_20307;
  wire       [31:0]   _zz_20308;
  wire       [15:0]   _zz_20309;
  wire       [31:0]   _zz_20310;
  wire       [31:0]   _zz_20311;
  wire       [31:0]   _zz_20312;
  wire       [15:0]   _zz_20313;
  wire       [31:0]   _zz_20314;
  wire       [31:0]   _zz_20315;
  wire       [31:0]   _zz_20316;
  wire       [31:0]   _zz_20317;
  wire       [31:0]   _zz_20318;
  wire       [31:0]   _zz_20319;
  wire       [23:0]   _zz_20320;
  wire       [31:0]   _zz_20321;
  wire       [15:0]   _zz_20322;
  wire       [31:0]   _zz_20323;
  wire       [31:0]   _zz_20324;
  wire       [31:0]   _zz_20325;
  wire       [31:0]   _zz_20326;
  wire       [31:0]   _zz_20327;
  wire       [23:0]   _zz_20328;
  wire       [31:0]   _zz_20329;
  wire       [15:0]   _zz_20330;
  wire       [31:0]   _zz_20331;
  wire       [31:0]   _zz_20332;
  wire       [31:0]   _zz_20333;
  wire       [31:0]   _zz_20334;
  wire       [31:0]   _zz_20335;
  wire       [23:0]   _zz_20336;
  wire       [31:0]   _zz_20337;
  wire       [15:0]   _zz_20338;
  wire       [31:0]   _zz_20339;
  wire       [31:0]   _zz_20340;
  wire       [31:0]   _zz_20341;
  wire       [31:0]   _zz_20342;
  wire       [31:0]   _zz_20343;
  wire       [23:0]   _zz_20344;
  wire       [31:0]   _zz_20345;
  wire       [15:0]   _zz_20346;
  wire       [15:0]   _zz_20347;
  wire       [31:0]   _zz_20348;
  wire       [31:0]   _zz_20349;
  wire       [15:0]   _zz_20350;
  wire       [31:0]   _zz_20351;
  wire       [31:0]   _zz_20352;
  wire       [31:0]   _zz_20353;
  wire       [15:0]   _zz_20354;
  wire       [31:0]   _zz_20355;
  wire       [31:0]   _zz_20356;
  wire       [31:0]   _zz_20357;
  wire       [31:0]   _zz_20358;
  wire       [31:0]   _zz_20359;
  wire       [31:0]   _zz_20360;
  wire       [23:0]   _zz_20361;
  wire       [31:0]   _zz_20362;
  wire       [15:0]   _zz_20363;
  wire       [31:0]   _zz_20364;
  wire       [31:0]   _zz_20365;
  wire       [31:0]   _zz_20366;
  wire       [31:0]   _zz_20367;
  wire       [31:0]   _zz_20368;
  wire       [23:0]   _zz_20369;
  wire       [31:0]   _zz_20370;
  wire       [15:0]   _zz_20371;
  wire       [31:0]   _zz_20372;
  wire       [31:0]   _zz_20373;
  wire       [31:0]   _zz_20374;
  wire       [31:0]   _zz_20375;
  wire       [31:0]   _zz_20376;
  wire       [23:0]   _zz_20377;
  wire       [31:0]   _zz_20378;
  wire       [15:0]   _zz_20379;
  wire       [31:0]   _zz_20380;
  wire       [31:0]   _zz_20381;
  wire       [31:0]   _zz_20382;
  wire       [31:0]   _zz_20383;
  wire       [31:0]   _zz_20384;
  wire       [23:0]   _zz_20385;
  wire       [31:0]   _zz_20386;
  wire       [15:0]   _zz_20387;
  wire       [15:0]   _zz_20388;
  wire       [31:0]   _zz_20389;
  wire       [31:0]   _zz_20390;
  wire       [15:0]   _zz_20391;
  wire       [31:0]   _zz_20392;
  wire       [31:0]   _zz_20393;
  wire       [31:0]   _zz_20394;
  wire       [15:0]   _zz_20395;
  wire       [31:0]   _zz_20396;
  wire       [31:0]   _zz_20397;
  wire       [31:0]   _zz_20398;
  wire       [31:0]   _zz_20399;
  wire       [31:0]   _zz_20400;
  wire       [31:0]   _zz_20401;
  wire       [23:0]   _zz_20402;
  wire       [31:0]   _zz_20403;
  wire       [15:0]   _zz_20404;
  wire       [31:0]   _zz_20405;
  wire       [31:0]   _zz_20406;
  wire       [31:0]   _zz_20407;
  wire       [31:0]   _zz_20408;
  wire       [31:0]   _zz_20409;
  wire       [23:0]   _zz_20410;
  wire       [31:0]   _zz_20411;
  wire       [15:0]   _zz_20412;
  wire       [31:0]   _zz_20413;
  wire       [31:0]   _zz_20414;
  wire       [31:0]   _zz_20415;
  wire       [31:0]   _zz_20416;
  wire       [31:0]   _zz_20417;
  wire       [23:0]   _zz_20418;
  wire       [31:0]   _zz_20419;
  wire       [15:0]   _zz_20420;
  wire       [31:0]   _zz_20421;
  wire       [31:0]   _zz_20422;
  wire       [31:0]   _zz_20423;
  wire       [31:0]   _zz_20424;
  wire       [31:0]   _zz_20425;
  wire       [23:0]   _zz_20426;
  wire       [31:0]   _zz_20427;
  wire       [15:0]   _zz_20428;
  wire       [15:0]   _zz_20429;
  wire       [31:0]   _zz_20430;
  wire       [31:0]   _zz_20431;
  wire       [15:0]   _zz_20432;
  wire       [31:0]   _zz_20433;
  wire       [31:0]   _zz_20434;
  wire       [31:0]   _zz_20435;
  wire       [15:0]   _zz_20436;
  wire       [31:0]   _zz_20437;
  wire       [31:0]   _zz_20438;
  wire       [31:0]   _zz_20439;
  wire       [31:0]   _zz_20440;
  wire       [31:0]   _zz_20441;
  wire       [31:0]   _zz_20442;
  wire       [23:0]   _zz_20443;
  wire       [31:0]   _zz_20444;
  wire       [15:0]   _zz_20445;
  wire       [31:0]   _zz_20446;
  wire       [31:0]   _zz_20447;
  wire       [31:0]   _zz_20448;
  wire       [31:0]   _zz_20449;
  wire       [31:0]   _zz_20450;
  wire       [23:0]   _zz_20451;
  wire       [31:0]   _zz_20452;
  wire       [15:0]   _zz_20453;
  wire       [31:0]   _zz_20454;
  wire       [31:0]   _zz_20455;
  wire       [31:0]   _zz_20456;
  wire       [31:0]   _zz_20457;
  wire       [31:0]   _zz_20458;
  wire       [23:0]   _zz_20459;
  wire       [31:0]   _zz_20460;
  wire       [15:0]   _zz_20461;
  wire       [31:0]   _zz_20462;
  wire       [31:0]   _zz_20463;
  wire       [31:0]   _zz_20464;
  wire       [31:0]   _zz_20465;
  wire       [31:0]   _zz_20466;
  wire       [23:0]   _zz_20467;
  wire       [31:0]   _zz_20468;
  wire       [15:0]   _zz_20469;
  wire       [15:0]   _zz_20470;
  wire       [31:0]   _zz_20471;
  wire       [31:0]   _zz_20472;
  wire       [15:0]   _zz_20473;
  wire       [31:0]   _zz_20474;
  wire       [31:0]   _zz_20475;
  wire       [31:0]   _zz_20476;
  wire       [15:0]   _zz_20477;
  wire       [31:0]   _zz_20478;
  wire       [31:0]   _zz_20479;
  wire       [31:0]   _zz_20480;
  wire       [31:0]   _zz_20481;
  wire       [31:0]   _zz_20482;
  wire       [31:0]   _zz_20483;
  wire       [23:0]   _zz_20484;
  wire       [31:0]   _zz_20485;
  wire       [15:0]   _zz_20486;
  wire       [31:0]   _zz_20487;
  wire       [31:0]   _zz_20488;
  wire       [31:0]   _zz_20489;
  wire       [31:0]   _zz_20490;
  wire       [31:0]   _zz_20491;
  wire       [23:0]   _zz_20492;
  wire       [31:0]   _zz_20493;
  wire       [15:0]   _zz_20494;
  wire       [31:0]   _zz_20495;
  wire       [31:0]   _zz_20496;
  wire       [31:0]   _zz_20497;
  wire       [31:0]   _zz_20498;
  wire       [31:0]   _zz_20499;
  wire       [23:0]   _zz_20500;
  wire       [31:0]   _zz_20501;
  wire       [15:0]   _zz_20502;
  wire       [31:0]   _zz_20503;
  wire       [31:0]   _zz_20504;
  wire       [31:0]   _zz_20505;
  wire       [31:0]   _zz_20506;
  wire       [31:0]   _zz_20507;
  wire       [23:0]   _zz_20508;
  wire       [31:0]   _zz_20509;
  wire       [15:0]   _zz_20510;
  wire       [15:0]   _zz_20511;
  wire       [31:0]   _zz_20512;
  wire       [31:0]   _zz_20513;
  wire       [15:0]   _zz_20514;
  wire       [31:0]   _zz_20515;
  wire       [31:0]   _zz_20516;
  wire       [31:0]   _zz_20517;
  wire       [15:0]   _zz_20518;
  wire       [31:0]   _zz_20519;
  wire       [31:0]   _zz_20520;
  wire       [31:0]   _zz_20521;
  wire       [31:0]   _zz_20522;
  wire       [31:0]   _zz_20523;
  wire       [31:0]   _zz_20524;
  wire       [23:0]   _zz_20525;
  wire       [31:0]   _zz_20526;
  wire       [15:0]   _zz_20527;
  wire       [31:0]   _zz_20528;
  wire       [31:0]   _zz_20529;
  wire       [31:0]   _zz_20530;
  wire       [31:0]   _zz_20531;
  wire       [31:0]   _zz_20532;
  wire       [23:0]   _zz_20533;
  wire       [31:0]   _zz_20534;
  wire       [15:0]   _zz_20535;
  wire       [31:0]   _zz_20536;
  wire       [31:0]   _zz_20537;
  wire       [31:0]   _zz_20538;
  wire       [31:0]   _zz_20539;
  wire       [31:0]   _zz_20540;
  wire       [23:0]   _zz_20541;
  wire       [31:0]   _zz_20542;
  wire       [15:0]   _zz_20543;
  wire       [31:0]   _zz_20544;
  wire       [31:0]   _zz_20545;
  wire       [31:0]   _zz_20546;
  wire       [31:0]   _zz_20547;
  wire       [31:0]   _zz_20548;
  wire       [23:0]   _zz_20549;
  wire       [31:0]   _zz_20550;
  wire       [15:0]   _zz_20551;
  wire       [15:0]   _zz_20552;
  wire       [31:0]   _zz_20553;
  wire       [31:0]   _zz_20554;
  wire       [15:0]   _zz_20555;
  wire       [31:0]   _zz_20556;
  wire       [31:0]   _zz_20557;
  wire       [31:0]   _zz_20558;
  wire       [15:0]   _zz_20559;
  wire       [31:0]   _zz_20560;
  wire       [31:0]   _zz_20561;
  wire       [31:0]   _zz_20562;
  wire       [31:0]   _zz_20563;
  wire       [31:0]   _zz_20564;
  wire       [31:0]   _zz_20565;
  wire       [23:0]   _zz_20566;
  wire       [31:0]   _zz_20567;
  wire       [15:0]   _zz_20568;
  wire       [31:0]   _zz_20569;
  wire       [31:0]   _zz_20570;
  wire       [31:0]   _zz_20571;
  wire       [31:0]   _zz_20572;
  wire       [31:0]   _zz_20573;
  wire       [23:0]   _zz_20574;
  wire       [31:0]   _zz_20575;
  wire       [15:0]   _zz_20576;
  wire       [31:0]   _zz_20577;
  wire       [31:0]   _zz_20578;
  wire       [31:0]   _zz_20579;
  wire       [31:0]   _zz_20580;
  wire       [31:0]   _zz_20581;
  wire       [23:0]   _zz_20582;
  wire       [31:0]   _zz_20583;
  wire       [15:0]   _zz_20584;
  wire       [31:0]   _zz_20585;
  wire       [31:0]   _zz_20586;
  wire       [31:0]   _zz_20587;
  wire       [31:0]   _zz_20588;
  wire       [31:0]   _zz_20589;
  wire       [23:0]   _zz_20590;
  wire       [31:0]   _zz_20591;
  wire       [15:0]   _zz_20592;
  wire       [15:0]   _zz_20593;
  wire       [31:0]   _zz_20594;
  wire       [31:0]   _zz_20595;
  wire       [15:0]   _zz_20596;
  wire       [31:0]   _zz_20597;
  wire       [31:0]   _zz_20598;
  wire       [31:0]   _zz_20599;
  wire       [15:0]   _zz_20600;
  wire       [31:0]   _zz_20601;
  wire       [31:0]   _zz_20602;
  wire       [31:0]   _zz_20603;
  wire       [31:0]   _zz_20604;
  wire       [31:0]   _zz_20605;
  wire       [31:0]   _zz_20606;
  wire       [23:0]   _zz_20607;
  wire       [31:0]   _zz_20608;
  wire       [15:0]   _zz_20609;
  wire       [31:0]   _zz_20610;
  wire       [31:0]   _zz_20611;
  wire       [31:0]   _zz_20612;
  wire       [31:0]   _zz_20613;
  wire       [31:0]   _zz_20614;
  wire       [23:0]   _zz_20615;
  wire       [31:0]   _zz_20616;
  wire       [15:0]   _zz_20617;
  wire       [31:0]   _zz_20618;
  wire       [31:0]   _zz_20619;
  wire       [31:0]   _zz_20620;
  wire       [31:0]   _zz_20621;
  wire       [31:0]   _zz_20622;
  wire       [23:0]   _zz_20623;
  wire       [31:0]   _zz_20624;
  wire       [15:0]   _zz_20625;
  wire       [31:0]   _zz_20626;
  wire       [31:0]   _zz_20627;
  wire       [31:0]   _zz_20628;
  wire       [31:0]   _zz_20629;
  wire       [31:0]   _zz_20630;
  wire       [23:0]   _zz_20631;
  wire       [31:0]   _zz_20632;
  wire       [15:0]   _zz_20633;
  wire       [15:0]   _zz_20634;
  wire       [31:0]   _zz_20635;
  wire       [31:0]   _zz_20636;
  wire       [15:0]   _zz_20637;
  wire       [31:0]   _zz_20638;
  wire       [31:0]   _zz_20639;
  wire       [31:0]   _zz_20640;
  wire       [15:0]   _zz_20641;
  wire       [31:0]   _zz_20642;
  wire       [31:0]   _zz_20643;
  wire       [31:0]   _zz_20644;
  wire       [31:0]   _zz_20645;
  wire       [31:0]   _zz_20646;
  wire       [31:0]   _zz_20647;
  wire       [23:0]   _zz_20648;
  wire       [31:0]   _zz_20649;
  wire       [15:0]   _zz_20650;
  wire       [31:0]   _zz_20651;
  wire       [31:0]   _zz_20652;
  wire       [31:0]   _zz_20653;
  wire       [31:0]   _zz_20654;
  wire       [31:0]   _zz_20655;
  wire       [23:0]   _zz_20656;
  wire       [31:0]   _zz_20657;
  wire       [15:0]   _zz_20658;
  wire       [31:0]   _zz_20659;
  wire       [31:0]   _zz_20660;
  wire       [31:0]   _zz_20661;
  wire       [31:0]   _zz_20662;
  wire       [31:0]   _zz_20663;
  wire       [23:0]   _zz_20664;
  wire       [31:0]   _zz_20665;
  wire       [15:0]   _zz_20666;
  wire       [31:0]   _zz_20667;
  wire       [31:0]   _zz_20668;
  wire       [31:0]   _zz_20669;
  wire       [31:0]   _zz_20670;
  wire       [31:0]   _zz_20671;
  wire       [23:0]   _zz_20672;
  wire       [31:0]   _zz_20673;
  wire       [15:0]   _zz_20674;
  wire       [15:0]   _zz_20675;
  wire       [31:0]   _zz_20676;
  wire       [31:0]   _zz_20677;
  wire       [15:0]   _zz_20678;
  wire       [31:0]   _zz_20679;
  wire       [31:0]   _zz_20680;
  wire       [31:0]   _zz_20681;
  wire       [15:0]   _zz_20682;
  wire       [31:0]   _zz_20683;
  wire       [31:0]   _zz_20684;
  wire       [31:0]   _zz_20685;
  wire       [31:0]   _zz_20686;
  wire       [31:0]   _zz_20687;
  wire       [31:0]   _zz_20688;
  wire       [23:0]   _zz_20689;
  wire       [31:0]   _zz_20690;
  wire       [15:0]   _zz_20691;
  wire       [31:0]   _zz_20692;
  wire       [31:0]   _zz_20693;
  wire       [31:0]   _zz_20694;
  wire       [31:0]   _zz_20695;
  wire       [31:0]   _zz_20696;
  wire       [23:0]   _zz_20697;
  wire       [31:0]   _zz_20698;
  wire       [15:0]   _zz_20699;
  wire       [31:0]   _zz_20700;
  wire       [31:0]   _zz_20701;
  wire       [31:0]   _zz_20702;
  wire       [31:0]   _zz_20703;
  wire       [31:0]   _zz_20704;
  wire       [23:0]   _zz_20705;
  wire       [31:0]   _zz_20706;
  wire       [15:0]   _zz_20707;
  wire       [31:0]   _zz_20708;
  wire       [31:0]   _zz_20709;
  wire       [31:0]   _zz_20710;
  wire       [31:0]   _zz_20711;
  wire       [31:0]   _zz_20712;
  wire       [23:0]   _zz_20713;
  wire       [31:0]   _zz_20714;
  wire       [15:0]   _zz_20715;
  wire       [15:0]   _zz_20716;
  wire       [31:0]   _zz_20717;
  wire       [31:0]   _zz_20718;
  wire       [15:0]   _zz_20719;
  wire       [31:0]   _zz_20720;
  wire       [31:0]   _zz_20721;
  wire       [31:0]   _zz_20722;
  wire       [15:0]   _zz_20723;
  wire       [31:0]   _zz_20724;
  wire       [31:0]   _zz_20725;
  wire       [31:0]   _zz_20726;
  wire       [31:0]   _zz_20727;
  wire       [31:0]   _zz_20728;
  wire       [31:0]   _zz_20729;
  wire       [23:0]   _zz_20730;
  wire       [31:0]   _zz_20731;
  wire       [15:0]   _zz_20732;
  wire       [31:0]   _zz_20733;
  wire       [31:0]   _zz_20734;
  wire       [31:0]   _zz_20735;
  wire       [31:0]   _zz_20736;
  wire       [31:0]   _zz_20737;
  wire       [23:0]   _zz_20738;
  wire       [31:0]   _zz_20739;
  wire       [15:0]   _zz_20740;
  wire       [31:0]   _zz_20741;
  wire       [31:0]   _zz_20742;
  wire       [31:0]   _zz_20743;
  wire       [31:0]   _zz_20744;
  wire       [31:0]   _zz_20745;
  wire       [23:0]   _zz_20746;
  wire       [31:0]   _zz_20747;
  wire       [15:0]   _zz_20748;
  wire       [31:0]   _zz_20749;
  wire       [31:0]   _zz_20750;
  wire       [31:0]   _zz_20751;
  wire       [31:0]   _zz_20752;
  wire       [31:0]   _zz_20753;
  wire       [23:0]   _zz_20754;
  wire       [31:0]   _zz_20755;
  wire       [15:0]   _zz_20756;
  wire       [15:0]   _zz_20757;
  wire       [31:0]   _zz_20758;
  wire       [31:0]   _zz_20759;
  wire       [15:0]   _zz_20760;
  wire       [31:0]   _zz_20761;
  wire       [31:0]   _zz_20762;
  wire       [31:0]   _zz_20763;
  wire       [15:0]   _zz_20764;
  wire       [31:0]   _zz_20765;
  wire       [31:0]   _zz_20766;
  wire       [31:0]   _zz_20767;
  wire       [31:0]   _zz_20768;
  wire       [31:0]   _zz_20769;
  wire       [31:0]   _zz_20770;
  wire       [23:0]   _zz_20771;
  wire       [31:0]   _zz_20772;
  wire       [15:0]   _zz_20773;
  wire       [31:0]   _zz_20774;
  wire       [31:0]   _zz_20775;
  wire       [31:0]   _zz_20776;
  wire       [31:0]   _zz_20777;
  wire       [31:0]   _zz_20778;
  wire       [23:0]   _zz_20779;
  wire       [31:0]   _zz_20780;
  wire       [15:0]   _zz_20781;
  wire       [31:0]   _zz_20782;
  wire       [31:0]   _zz_20783;
  wire       [31:0]   _zz_20784;
  wire       [31:0]   _zz_20785;
  wire       [31:0]   _zz_20786;
  wire       [23:0]   _zz_20787;
  wire       [31:0]   _zz_20788;
  wire       [15:0]   _zz_20789;
  wire       [31:0]   _zz_20790;
  wire       [31:0]   _zz_20791;
  wire       [31:0]   _zz_20792;
  wire       [31:0]   _zz_20793;
  wire       [31:0]   _zz_20794;
  wire       [23:0]   _zz_20795;
  wire       [31:0]   _zz_20796;
  wire       [15:0]   _zz_20797;
  wire       [15:0]   _zz_20798;
  wire       [31:0]   _zz_20799;
  wire       [31:0]   _zz_20800;
  wire       [15:0]   _zz_20801;
  wire       [31:0]   _zz_20802;
  wire       [31:0]   _zz_20803;
  wire       [31:0]   _zz_20804;
  wire       [15:0]   _zz_20805;
  wire       [31:0]   _zz_20806;
  wire       [31:0]   _zz_20807;
  wire       [31:0]   _zz_20808;
  wire       [31:0]   _zz_20809;
  wire       [31:0]   _zz_20810;
  wire       [31:0]   _zz_20811;
  wire       [23:0]   _zz_20812;
  wire       [31:0]   _zz_20813;
  wire       [15:0]   _zz_20814;
  wire       [31:0]   _zz_20815;
  wire       [31:0]   _zz_20816;
  wire       [31:0]   _zz_20817;
  wire       [31:0]   _zz_20818;
  wire       [31:0]   _zz_20819;
  wire       [23:0]   _zz_20820;
  wire       [31:0]   _zz_20821;
  wire       [15:0]   _zz_20822;
  wire       [31:0]   _zz_20823;
  wire       [31:0]   _zz_20824;
  wire       [31:0]   _zz_20825;
  wire       [31:0]   _zz_20826;
  wire       [31:0]   _zz_20827;
  wire       [23:0]   _zz_20828;
  wire       [31:0]   _zz_20829;
  wire       [15:0]   _zz_20830;
  wire       [31:0]   _zz_20831;
  wire       [31:0]   _zz_20832;
  wire       [31:0]   _zz_20833;
  wire       [31:0]   _zz_20834;
  wire       [31:0]   _zz_20835;
  wire       [23:0]   _zz_20836;
  wire       [31:0]   _zz_20837;
  wire       [15:0]   _zz_20838;
  wire       [15:0]   _zz_20839;
  wire       [31:0]   _zz_20840;
  wire       [31:0]   _zz_20841;
  wire       [15:0]   _zz_20842;
  wire       [31:0]   _zz_20843;
  wire       [31:0]   _zz_20844;
  wire       [31:0]   _zz_20845;
  wire       [15:0]   _zz_20846;
  wire       [31:0]   _zz_20847;
  wire       [31:0]   _zz_20848;
  wire       [31:0]   _zz_20849;
  wire       [31:0]   _zz_20850;
  wire       [31:0]   _zz_20851;
  wire       [31:0]   _zz_20852;
  wire       [23:0]   _zz_20853;
  wire       [31:0]   _zz_20854;
  wire       [15:0]   _zz_20855;
  wire       [31:0]   _zz_20856;
  wire       [31:0]   _zz_20857;
  wire       [31:0]   _zz_20858;
  wire       [31:0]   _zz_20859;
  wire       [31:0]   _zz_20860;
  wire       [23:0]   _zz_20861;
  wire       [31:0]   _zz_20862;
  wire       [15:0]   _zz_20863;
  wire       [31:0]   _zz_20864;
  wire       [31:0]   _zz_20865;
  wire       [31:0]   _zz_20866;
  wire       [31:0]   _zz_20867;
  wire       [31:0]   _zz_20868;
  wire       [23:0]   _zz_20869;
  wire       [31:0]   _zz_20870;
  wire       [15:0]   _zz_20871;
  wire       [31:0]   _zz_20872;
  wire       [31:0]   _zz_20873;
  wire       [31:0]   _zz_20874;
  wire       [31:0]   _zz_20875;
  wire       [31:0]   _zz_20876;
  wire       [23:0]   _zz_20877;
  wire       [31:0]   _zz_20878;
  wire       [15:0]   _zz_20879;
  wire       [15:0]   _zz_20880;
  wire       [31:0]   _zz_20881;
  wire       [31:0]   _zz_20882;
  wire       [15:0]   _zz_20883;
  wire       [31:0]   _zz_20884;
  wire       [31:0]   _zz_20885;
  wire       [31:0]   _zz_20886;
  wire       [15:0]   _zz_20887;
  wire       [31:0]   _zz_20888;
  wire       [31:0]   _zz_20889;
  wire       [31:0]   _zz_20890;
  wire       [31:0]   _zz_20891;
  wire       [31:0]   _zz_20892;
  wire       [31:0]   _zz_20893;
  wire       [23:0]   _zz_20894;
  wire       [31:0]   _zz_20895;
  wire       [15:0]   _zz_20896;
  wire       [31:0]   _zz_20897;
  wire       [31:0]   _zz_20898;
  wire       [31:0]   _zz_20899;
  wire       [31:0]   _zz_20900;
  wire       [31:0]   _zz_20901;
  wire       [23:0]   _zz_20902;
  wire       [31:0]   _zz_20903;
  wire       [15:0]   _zz_20904;
  wire       [31:0]   _zz_20905;
  wire       [31:0]   _zz_20906;
  wire       [31:0]   _zz_20907;
  wire       [31:0]   _zz_20908;
  wire       [31:0]   _zz_20909;
  wire       [23:0]   _zz_20910;
  wire       [31:0]   _zz_20911;
  wire       [15:0]   _zz_20912;
  wire       [31:0]   _zz_20913;
  wire       [31:0]   _zz_20914;
  wire       [31:0]   _zz_20915;
  wire       [31:0]   _zz_20916;
  wire       [31:0]   _zz_20917;
  wire       [23:0]   _zz_20918;
  wire       [31:0]   _zz_20919;
  wire       [15:0]   _zz_20920;
  wire       [15:0]   _zz_20921;
  wire       [31:0]   _zz_20922;
  wire       [31:0]   _zz_20923;
  wire       [15:0]   _zz_20924;
  wire       [31:0]   _zz_20925;
  wire       [31:0]   _zz_20926;
  wire       [31:0]   _zz_20927;
  wire       [15:0]   _zz_20928;
  wire       [31:0]   _zz_20929;
  wire       [31:0]   _zz_20930;
  wire       [31:0]   _zz_20931;
  wire       [31:0]   _zz_20932;
  wire       [31:0]   _zz_20933;
  wire       [31:0]   _zz_20934;
  wire       [23:0]   _zz_20935;
  wire       [31:0]   _zz_20936;
  wire       [15:0]   _zz_20937;
  wire       [31:0]   _zz_20938;
  wire       [31:0]   _zz_20939;
  wire       [31:0]   _zz_20940;
  wire       [31:0]   _zz_20941;
  wire       [31:0]   _zz_20942;
  wire       [23:0]   _zz_20943;
  wire       [31:0]   _zz_20944;
  wire       [15:0]   _zz_20945;
  wire       [31:0]   _zz_20946;
  wire       [31:0]   _zz_20947;
  wire       [31:0]   _zz_20948;
  wire       [31:0]   _zz_20949;
  wire       [31:0]   _zz_20950;
  wire       [23:0]   _zz_20951;
  wire       [31:0]   _zz_20952;
  wire       [15:0]   _zz_20953;
  wire       [31:0]   _zz_20954;
  wire       [31:0]   _zz_20955;
  wire       [31:0]   _zz_20956;
  wire       [31:0]   _zz_20957;
  wire       [31:0]   _zz_20958;
  wire       [23:0]   _zz_20959;
  wire       [31:0]   _zz_20960;
  wire       [15:0]   _zz_20961;
  wire       [15:0]   _zz_20962;
  wire       [31:0]   _zz_20963;
  wire       [31:0]   _zz_20964;
  wire       [15:0]   _zz_20965;
  wire       [31:0]   _zz_20966;
  wire       [31:0]   _zz_20967;
  wire       [31:0]   _zz_20968;
  wire       [15:0]   _zz_20969;
  wire       [31:0]   _zz_20970;
  wire       [31:0]   _zz_20971;
  wire       [31:0]   _zz_20972;
  wire       [31:0]   _zz_20973;
  wire       [31:0]   _zz_20974;
  wire       [31:0]   _zz_20975;
  wire       [23:0]   _zz_20976;
  wire       [31:0]   _zz_20977;
  wire       [15:0]   _zz_20978;
  wire       [31:0]   _zz_20979;
  wire       [31:0]   _zz_20980;
  wire       [31:0]   _zz_20981;
  wire       [31:0]   _zz_20982;
  wire       [31:0]   _zz_20983;
  wire       [23:0]   _zz_20984;
  wire       [31:0]   _zz_20985;
  wire       [15:0]   _zz_20986;
  wire       [31:0]   _zz_20987;
  wire       [31:0]   _zz_20988;
  wire       [31:0]   _zz_20989;
  wire       [31:0]   _zz_20990;
  wire       [31:0]   _zz_20991;
  wire       [23:0]   _zz_20992;
  wire       [31:0]   _zz_20993;
  wire       [15:0]   _zz_20994;
  wire       [31:0]   _zz_20995;
  wire       [31:0]   _zz_20996;
  wire       [31:0]   _zz_20997;
  wire       [31:0]   _zz_20998;
  wire       [31:0]   _zz_20999;
  wire       [23:0]   _zz_21000;
  wire       [31:0]   _zz_21001;
  wire       [15:0]   _zz_21002;
  wire       [15:0]   _zz_21003;
  wire       [31:0]   _zz_21004;
  wire       [31:0]   _zz_21005;
  wire       [15:0]   _zz_21006;
  wire       [31:0]   _zz_21007;
  wire       [31:0]   _zz_21008;
  wire       [31:0]   _zz_21009;
  wire       [15:0]   _zz_21010;
  wire       [31:0]   _zz_21011;
  wire       [31:0]   _zz_21012;
  wire       [31:0]   _zz_21013;
  wire       [31:0]   _zz_21014;
  wire       [31:0]   _zz_21015;
  wire       [31:0]   _zz_21016;
  wire       [23:0]   _zz_21017;
  wire       [31:0]   _zz_21018;
  wire       [15:0]   _zz_21019;
  wire       [31:0]   _zz_21020;
  wire       [31:0]   _zz_21021;
  wire       [31:0]   _zz_21022;
  wire       [31:0]   _zz_21023;
  wire       [31:0]   _zz_21024;
  wire       [23:0]   _zz_21025;
  wire       [31:0]   _zz_21026;
  wire       [15:0]   _zz_21027;
  wire       [31:0]   _zz_21028;
  wire       [31:0]   _zz_21029;
  wire       [31:0]   _zz_21030;
  wire       [31:0]   _zz_21031;
  wire       [31:0]   _zz_21032;
  wire       [23:0]   _zz_21033;
  wire       [31:0]   _zz_21034;
  wire       [15:0]   _zz_21035;
  wire       [31:0]   _zz_21036;
  wire       [31:0]   _zz_21037;
  wire       [31:0]   _zz_21038;
  wire       [31:0]   _zz_21039;
  wire       [31:0]   _zz_21040;
  wire       [23:0]   _zz_21041;
  wire       [31:0]   _zz_21042;
  wire       [15:0]   _zz_21043;
  wire       [15:0]   _zz_21044;
  wire       [31:0]   _zz_21045;
  wire       [31:0]   _zz_21046;
  wire       [15:0]   _zz_21047;
  wire       [31:0]   _zz_21048;
  wire       [31:0]   _zz_21049;
  wire       [31:0]   _zz_21050;
  wire       [15:0]   _zz_21051;
  wire       [31:0]   _zz_21052;
  wire       [31:0]   _zz_21053;
  wire       [31:0]   _zz_21054;
  wire       [31:0]   _zz_21055;
  wire       [31:0]   _zz_21056;
  wire       [31:0]   _zz_21057;
  wire       [23:0]   _zz_21058;
  wire       [31:0]   _zz_21059;
  wire       [15:0]   _zz_21060;
  wire       [31:0]   _zz_21061;
  wire       [31:0]   _zz_21062;
  wire       [31:0]   _zz_21063;
  wire       [31:0]   _zz_21064;
  wire       [31:0]   _zz_21065;
  wire       [23:0]   _zz_21066;
  wire       [31:0]   _zz_21067;
  wire       [15:0]   _zz_21068;
  wire       [31:0]   _zz_21069;
  wire       [31:0]   _zz_21070;
  wire       [31:0]   _zz_21071;
  wire       [31:0]   _zz_21072;
  wire       [31:0]   _zz_21073;
  wire       [23:0]   _zz_21074;
  wire       [31:0]   _zz_21075;
  wire       [15:0]   _zz_21076;
  wire       [31:0]   _zz_21077;
  wire       [31:0]   _zz_21078;
  wire       [31:0]   _zz_21079;
  wire       [31:0]   _zz_21080;
  wire       [31:0]   _zz_21081;
  wire       [23:0]   _zz_21082;
  wire       [31:0]   _zz_21083;
  wire       [15:0]   _zz_21084;
  wire       [15:0]   _zz_21085;
  wire       [31:0]   _zz_21086;
  wire       [31:0]   _zz_21087;
  wire       [15:0]   _zz_21088;
  wire       [31:0]   _zz_21089;
  wire       [31:0]   _zz_21090;
  wire       [31:0]   _zz_21091;
  wire       [15:0]   _zz_21092;
  wire       [31:0]   _zz_21093;
  wire       [31:0]   _zz_21094;
  wire       [31:0]   _zz_21095;
  wire       [31:0]   _zz_21096;
  wire       [31:0]   _zz_21097;
  wire       [31:0]   _zz_21098;
  wire       [23:0]   _zz_21099;
  wire       [31:0]   _zz_21100;
  wire       [15:0]   _zz_21101;
  wire       [31:0]   _zz_21102;
  wire       [31:0]   _zz_21103;
  wire       [31:0]   _zz_21104;
  wire       [31:0]   _zz_21105;
  wire       [31:0]   _zz_21106;
  wire       [23:0]   _zz_21107;
  wire       [31:0]   _zz_21108;
  wire       [15:0]   _zz_21109;
  wire       [31:0]   _zz_21110;
  wire       [31:0]   _zz_21111;
  wire       [31:0]   _zz_21112;
  wire       [31:0]   _zz_21113;
  wire       [31:0]   _zz_21114;
  wire       [23:0]   _zz_21115;
  wire       [31:0]   _zz_21116;
  wire       [15:0]   _zz_21117;
  wire       [31:0]   _zz_21118;
  wire       [31:0]   _zz_21119;
  wire       [31:0]   _zz_21120;
  wire       [31:0]   _zz_21121;
  wire       [31:0]   _zz_21122;
  wire       [23:0]   _zz_21123;
  wire       [31:0]   _zz_21124;
  wire       [15:0]   _zz_21125;
  wire       [15:0]   _zz_21126;
  wire       [31:0]   _zz_21127;
  wire       [31:0]   _zz_21128;
  wire       [15:0]   _zz_21129;
  wire       [31:0]   _zz_21130;
  wire       [31:0]   _zz_21131;
  wire       [31:0]   _zz_21132;
  wire       [15:0]   _zz_21133;
  wire       [31:0]   _zz_21134;
  wire       [31:0]   _zz_21135;
  wire       [31:0]   _zz_21136;
  wire       [31:0]   _zz_21137;
  wire       [31:0]   _zz_21138;
  wire       [31:0]   _zz_21139;
  wire       [23:0]   _zz_21140;
  wire       [31:0]   _zz_21141;
  wire       [15:0]   _zz_21142;
  wire       [31:0]   _zz_21143;
  wire       [31:0]   _zz_21144;
  wire       [31:0]   _zz_21145;
  wire       [31:0]   _zz_21146;
  wire       [31:0]   _zz_21147;
  wire       [23:0]   _zz_21148;
  wire       [31:0]   _zz_21149;
  wire       [15:0]   _zz_21150;
  wire       [31:0]   _zz_21151;
  wire       [31:0]   _zz_21152;
  wire       [31:0]   _zz_21153;
  wire       [31:0]   _zz_21154;
  wire       [31:0]   _zz_21155;
  wire       [23:0]   _zz_21156;
  wire       [31:0]   _zz_21157;
  wire       [15:0]   _zz_21158;
  wire       [31:0]   _zz_21159;
  wire       [31:0]   _zz_21160;
  wire       [31:0]   _zz_21161;
  wire       [31:0]   _zz_21162;
  wire       [31:0]   _zz_21163;
  wire       [23:0]   _zz_21164;
  wire       [31:0]   _zz_21165;
  wire       [15:0]   _zz_21166;
  wire       [15:0]   _zz_21167;
  wire       [31:0]   _zz_21168;
  wire       [31:0]   _zz_21169;
  wire       [15:0]   _zz_21170;
  wire       [31:0]   _zz_21171;
  wire       [31:0]   _zz_21172;
  wire       [31:0]   _zz_21173;
  wire       [15:0]   _zz_21174;
  wire       [31:0]   _zz_21175;
  wire       [31:0]   _zz_21176;
  wire       [31:0]   _zz_21177;
  wire       [31:0]   _zz_21178;
  wire       [31:0]   _zz_21179;
  wire       [31:0]   _zz_21180;
  wire       [23:0]   _zz_21181;
  wire       [31:0]   _zz_21182;
  wire       [15:0]   _zz_21183;
  wire       [31:0]   _zz_21184;
  wire       [31:0]   _zz_21185;
  wire       [31:0]   _zz_21186;
  wire       [31:0]   _zz_21187;
  wire       [31:0]   _zz_21188;
  wire       [23:0]   _zz_21189;
  wire       [31:0]   _zz_21190;
  wire       [15:0]   _zz_21191;
  wire       [31:0]   _zz_21192;
  wire       [31:0]   _zz_21193;
  wire       [31:0]   _zz_21194;
  wire       [31:0]   _zz_21195;
  wire       [31:0]   _zz_21196;
  wire       [23:0]   _zz_21197;
  wire       [31:0]   _zz_21198;
  wire       [15:0]   _zz_21199;
  wire       [31:0]   _zz_21200;
  wire       [31:0]   _zz_21201;
  wire       [31:0]   _zz_21202;
  wire       [31:0]   _zz_21203;
  wire       [31:0]   _zz_21204;
  wire       [23:0]   _zz_21205;
  wire       [31:0]   _zz_21206;
  wire       [15:0]   _zz_21207;
  wire       [15:0]   _zz_21208;
  wire       [31:0]   _zz_21209;
  wire       [31:0]   _zz_21210;
  wire       [15:0]   _zz_21211;
  wire       [31:0]   _zz_21212;
  wire       [31:0]   _zz_21213;
  wire       [31:0]   _zz_21214;
  wire       [15:0]   _zz_21215;
  wire       [31:0]   _zz_21216;
  wire       [31:0]   _zz_21217;
  wire       [31:0]   _zz_21218;
  wire       [31:0]   _zz_21219;
  wire       [31:0]   _zz_21220;
  wire       [31:0]   _zz_21221;
  wire       [23:0]   _zz_21222;
  wire       [31:0]   _zz_21223;
  wire       [15:0]   _zz_21224;
  wire       [31:0]   _zz_21225;
  wire       [31:0]   _zz_21226;
  wire       [31:0]   _zz_21227;
  wire       [31:0]   _zz_21228;
  wire       [31:0]   _zz_21229;
  wire       [23:0]   _zz_21230;
  wire       [31:0]   _zz_21231;
  wire       [15:0]   _zz_21232;
  wire       [31:0]   _zz_21233;
  wire       [31:0]   _zz_21234;
  wire       [31:0]   _zz_21235;
  wire       [31:0]   _zz_21236;
  wire       [31:0]   _zz_21237;
  wire       [23:0]   _zz_21238;
  wire       [31:0]   _zz_21239;
  wire       [15:0]   _zz_21240;
  wire       [31:0]   _zz_21241;
  wire       [31:0]   _zz_21242;
  wire       [31:0]   _zz_21243;
  wire       [31:0]   _zz_21244;
  wire       [31:0]   _zz_21245;
  wire       [23:0]   _zz_21246;
  wire       [31:0]   _zz_21247;
  wire       [15:0]   _zz_21248;
  wire       [15:0]   _zz_21249;
  wire       [31:0]   _zz_21250;
  wire       [31:0]   _zz_21251;
  wire       [15:0]   _zz_21252;
  wire       [31:0]   _zz_21253;
  wire       [31:0]   _zz_21254;
  wire       [31:0]   _zz_21255;
  wire       [15:0]   _zz_21256;
  wire       [31:0]   _zz_21257;
  wire       [31:0]   _zz_21258;
  wire       [31:0]   _zz_21259;
  wire       [31:0]   _zz_21260;
  wire       [31:0]   _zz_21261;
  wire       [31:0]   _zz_21262;
  wire       [23:0]   _zz_21263;
  wire       [31:0]   _zz_21264;
  wire       [15:0]   _zz_21265;
  wire       [31:0]   _zz_21266;
  wire       [31:0]   _zz_21267;
  wire       [31:0]   _zz_21268;
  wire       [31:0]   _zz_21269;
  wire       [31:0]   _zz_21270;
  wire       [23:0]   _zz_21271;
  wire       [31:0]   _zz_21272;
  wire       [15:0]   _zz_21273;
  wire       [31:0]   _zz_21274;
  wire       [31:0]   _zz_21275;
  wire       [31:0]   _zz_21276;
  wire       [31:0]   _zz_21277;
  wire       [31:0]   _zz_21278;
  wire       [23:0]   _zz_21279;
  wire       [31:0]   _zz_21280;
  wire       [15:0]   _zz_21281;
  wire       [31:0]   _zz_21282;
  wire       [31:0]   _zz_21283;
  wire       [31:0]   _zz_21284;
  wire       [31:0]   _zz_21285;
  wire       [31:0]   _zz_21286;
  wire       [23:0]   _zz_21287;
  wire       [31:0]   _zz_21288;
  wire       [15:0]   _zz_21289;
  wire       [15:0]   _zz_21290;
  wire       [31:0]   _zz_21291;
  wire       [31:0]   _zz_21292;
  wire       [15:0]   _zz_21293;
  wire       [31:0]   _zz_21294;
  wire       [31:0]   _zz_21295;
  wire       [31:0]   _zz_21296;
  wire       [15:0]   _zz_21297;
  wire       [31:0]   _zz_21298;
  wire       [31:0]   _zz_21299;
  wire       [31:0]   _zz_21300;
  wire       [31:0]   _zz_21301;
  wire       [31:0]   _zz_21302;
  wire       [31:0]   _zz_21303;
  wire       [23:0]   _zz_21304;
  wire       [31:0]   _zz_21305;
  wire       [15:0]   _zz_21306;
  wire       [31:0]   _zz_21307;
  wire       [31:0]   _zz_21308;
  wire       [31:0]   _zz_21309;
  wire       [31:0]   _zz_21310;
  wire       [31:0]   _zz_21311;
  wire       [23:0]   _zz_21312;
  wire       [31:0]   _zz_21313;
  wire       [15:0]   _zz_21314;
  wire       [31:0]   _zz_21315;
  wire       [31:0]   _zz_21316;
  wire       [31:0]   _zz_21317;
  wire       [31:0]   _zz_21318;
  wire       [31:0]   _zz_21319;
  wire       [23:0]   _zz_21320;
  wire       [31:0]   _zz_21321;
  wire       [15:0]   _zz_21322;
  wire       [31:0]   _zz_21323;
  wire       [31:0]   _zz_21324;
  wire       [31:0]   _zz_21325;
  wire       [31:0]   _zz_21326;
  wire       [31:0]   _zz_21327;
  wire       [23:0]   _zz_21328;
  wire       [31:0]   _zz_21329;
  wire       [15:0]   _zz_21330;
  wire       [15:0]   _zz_21331;
  wire       [31:0]   _zz_21332;
  wire       [31:0]   _zz_21333;
  wire       [15:0]   _zz_21334;
  wire       [31:0]   _zz_21335;
  wire       [31:0]   _zz_21336;
  wire       [31:0]   _zz_21337;
  wire       [15:0]   _zz_21338;
  wire       [31:0]   _zz_21339;
  wire       [31:0]   _zz_21340;
  wire       [31:0]   _zz_21341;
  wire       [31:0]   _zz_21342;
  wire       [31:0]   _zz_21343;
  wire       [31:0]   _zz_21344;
  wire       [23:0]   _zz_21345;
  wire       [31:0]   _zz_21346;
  wire       [15:0]   _zz_21347;
  wire       [31:0]   _zz_21348;
  wire       [31:0]   _zz_21349;
  wire       [31:0]   _zz_21350;
  wire       [31:0]   _zz_21351;
  wire       [31:0]   _zz_21352;
  wire       [23:0]   _zz_21353;
  wire       [31:0]   _zz_21354;
  wire       [15:0]   _zz_21355;
  wire       [31:0]   _zz_21356;
  wire       [31:0]   _zz_21357;
  wire       [31:0]   _zz_21358;
  wire       [31:0]   _zz_21359;
  wire       [31:0]   _zz_21360;
  wire       [23:0]   _zz_21361;
  wire       [31:0]   _zz_21362;
  wire       [15:0]   _zz_21363;
  wire       [31:0]   _zz_21364;
  wire       [31:0]   _zz_21365;
  wire       [31:0]   _zz_21366;
  wire       [31:0]   _zz_21367;
  wire       [31:0]   _zz_21368;
  wire       [23:0]   _zz_21369;
  wire       [31:0]   _zz_21370;
  wire       [15:0]   _zz_21371;
  wire       [15:0]   _zz_21372;
  wire       [31:0]   _zz_21373;
  wire       [31:0]   _zz_21374;
  wire       [15:0]   _zz_21375;
  wire       [31:0]   _zz_21376;
  wire       [31:0]   _zz_21377;
  wire       [31:0]   _zz_21378;
  wire       [15:0]   _zz_21379;
  wire       [31:0]   _zz_21380;
  wire       [31:0]   _zz_21381;
  wire       [31:0]   _zz_21382;
  wire       [31:0]   _zz_21383;
  wire       [31:0]   _zz_21384;
  wire       [31:0]   _zz_21385;
  wire       [23:0]   _zz_21386;
  wire       [31:0]   _zz_21387;
  wire       [15:0]   _zz_21388;
  wire       [31:0]   _zz_21389;
  wire       [31:0]   _zz_21390;
  wire       [31:0]   _zz_21391;
  wire       [31:0]   _zz_21392;
  wire       [31:0]   _zz_21393;
  wire       [23:0]   _zz_21394;
  wire       [31:0]   _zz_21395;
  wire       [15:0]   _zz_21396;
  wire       [31:0]   _zz_21397;
  wire       [31:0]   _zz_21398;
  wire       [31:0]   _zz_21399;
  wire       [31:0]   _zz_21400;
  wire       [31:0]   _zz_21401;
  wire       [23:0]   _zz_21402;
  wire       [31:0]   _zz_21403;
  wire       [15:0]   _zz_21404;
  wire       [31:0]   _zz_21405;
  wire       [31:0]   _zz_21406;
  wire       [31:0]   _zz_21407;
  wire       [31:0]   _zz_21408;
  wire       [31:0]   _zz_21409;
  wire       [23:0]   _zz_21410;
  wire       [31:0]   _zz_21411;
  wire       [15:0]   _zz_21412;
  wire       [15:0]   _zz_21413;
  wire       [31:0]   _zz_21414;
  wire       [31:0]   _zz_21415;
  wire       [15:0]   _zz_21416;
  wire       [31:0]   _zz_21417;
  wire       [31:0]   _zz_21418;
  wire       [31:0]   _zz_21419;
  wire       [15:0]   _zz_21420;
  wire       [31:0]   _zz_21421;
  wire       [31:0]   _zz_21422;
  wire       [31:0]   _zz_21423;
  wire       [31:0]   _zz_21424;
  wire       [31:0]   _zz_21425;
  wire       [31:0]   _zz_21426;
  wire       [23:0]   _zz_21427;
  wire       [31:0]   _zz_21428;
  wire       [15:0]   _zz_21429;
  wire       [31:0]   _zz_21430;
  wire       [31:0]   _zz_21431;
  wire       [31:0]   _zz_21432;
  wire       [31:0]   _zz_21433;
  wire       [31:0]   _zz_21434;
  wire       [23:0]   _zz_21435;
  wire       [31:0]   _zz_21436;
  wire       [15:0]   _zz_21437;
  wire       [31:0]   _zz_21438;
  wire       [31:0]   _zz_21439;
  wire       [31:0]   _zz_21440;
  wire       [31:0]   _zz_21441;
  wire       [31:0]   _zz_21442;
  wire       [23:0]   _zz_21443;
  wire       [31:0]   _zz_21444;
  wire       [15:0]   _zz_21445;
  wire       [31:0]   _zz_21446;
  wire       [31:0]   _zz_21447;
  wire       [31:0]   _zz_21448;
  wire       [31:0]   _zz_21449;
  wire       [31:0]   _zz_21450;
  wire       [23:0]   _zz_21451;
  wire       [31:0]   _zz_21452;
  wire       [15:0]   _zz_21453;
  wire       [15:0]   _zz_21454;
  wire       [31:0]   _zz_21455;
  wire       [31:0]   _zz_21456;
  wire       [15:0]   _zz_21457;
  wire       [31:0]   _zz_21458;
  wire       [31:0]   _zz_21459;
  wire       [31:0]   _zz_21460;
  wire       [15:0]   _zz_21461;
  wire       [31:0]   _zz_21462;
  wire       [31:0]   _zz_21463;
  wire       [31:0]   _zz_21464;
  wire       [31:0]   _zz_21465;
  wire       [31:0]   _zz_21466;
  wire       [31:0]   _zz_21467;
  wire       [23:0]   _zz_21468;
  wire       [31:0]   _zz_21469;
  wire       [15:0]   _zz_21470;
  wire       [31:0]   _zz_21471;
  wire       [31:0]   _zz_21472;
  wire       [31:0]   _zz_21473;
  wire       [31:0]   _zz_21474;
  wire       [31:0]   _zz_21475;
  wire       [23:0]   _zz_21476;
  wire       [31:0]   _zz_21477;
  wire       [15:0]   _zz_21478;
  wire       [31:0]   _zz_21479;
  wire       [31:0]   _zz_21480;
  wire       [31:0]   _zz_21481;
  wire       [31:0]   _zz_21482;
  wire       [31:0]   _zz_21483;
  wire       [23:0]   _zz_21484;
  wire       [31:0]   _zz_21485;
  wire       [15:0]   _zz_21486;
  wire       [31:0]   _zz_21487;
  wire       [31:0]   _zz_21488;
  wire       [31:0]   _zz_21489;
  wire       [31:0]   _zz_21490;
  wire       [31:0]   _zz_21491;
  wire       [23:0]   _zz_21492;
  wire       [31:0]   _zz_21493;
  wire       [15:0]   _zz_21494;
  wire       [15:0]   _zz_21495;
  wire       [31:0]   _zz_21496;
  wire       [31:0]   _zz_21497;
  wire       [15:0]   _zz_21498;
  wire       [31:0]   _zz_21499;
  wire       [31:0]   _zz_21500;
  wire       [31:0]   _zz_21501;
  wire       [15:0]   _zz_21502;
  wire       [31:0]   _zz_21503;
  wire       [31:0]   _zz_21504;
  wire       [31:0]   _zz_21505;
  wire       [31:0]   _zz_21506;
  wire       [31:0]   _zz_21507;
  wire       [31:0]   _zz_21508;
  wire       [23:0]   _zz_21509;
  wire       [31:0]   _zz_21510;
  wire       [15:0]   _zz_21511;
  wire       [31:0]   _zz_21512;
  wire       [31:0]   _zz_21513;
  wire       [31:0]   _zz_21514;
  wire       [31:0]   _zz_21515;
  wire       [31:0]   _zz_21516;
  wire       [23:0]   _zz_21517;
  wire       [31:0]   _zz_21518;
  wire       [15:0]   _zz_21519;
  wire       [31:0]   _zz_21520;
  wire       [31:0]   _zz_21521;
  wire       [31:0]   _zz_21522;
  wire       [31:0]   _zz_21523;
  wire       [31:0]   _zz_21524;
  wire       [23:0]   _zz_21525;
  wire       [31:0]   _zz_21526;
  wire       [15:0]   _zz_21527;
  wire       [31:0]   _zz_21528;
  wire       [31:0]   _zz_21529;
  wire       [31:0]   _zz_21530;
  wire       [31:0]   _zz_21531;
  wire       [31:0]   _zz_21532;
  wire       [23:0]   _zz_21533;
  wire       [31:0]   _zz_21534;
  wire       [15:0]   _zz_21535;
  wire       [15:0]   _zz_21536;
  wire       [31:0]   _zz_21537;
  wire       [31:0]   _zz_21538;
  wire       [15:0]   _zz_21539;
  wire       [31:0]   _zz_21540;
  wire       [31:0]   _zz_21541;
  wire       [31:0]   _zz_21542;
  wire       [15:0]   _zz_21543;
  wire       [31:0]   _zz_21544;
  wire       [31:0]   _zz_21545;
  wire       [31:0]   _zz_21546;
  wire       [31:0]   _zz_21547;
  wire       [31:0]   _zz_21548;
  wire       [31:0]   _zz_21549;
  wire       [23:0]   _zz_21550;
  wire       [31:0]   _zz_21551;
  wire       [15:0]   _zz_21552;
  wire       [31:0]   _zz_21553;
  wire       [31:0]   _zz_21554;
  wire       [31:0]   _zz_21555;
  wire       [31:0]   _zz_21556;
  wire       [31:0]   _zz_21557;
  wire       [23:0]   _zz_21558;
  wire       [31:0]   _zz_21559;
  wire       [15:0]   _zz_21560;
  wire       [31:0]   _zz_21561;
  wire       [31:0]   _zz_21562;
  wire       [31:0]   _zz_21563;
  wire       [31:0]   _zz_21564;
  wire       [31:0]   _zz_21565;
  wire       [23:0]   _zz_21566;
  wire       [31:0]   _zz_21567;
  wire       [15:0]   _zz_21568;
  wire       [31:0]   _zz_21569;
  wire       [31:0]   _zz_21570;
  wire       [31:0]   _zz_21571;
  wire       [31:0]   _zz_21572;
  wire       [31:0]   _zz_21573;
  wire       [23:0]   _zz_21574;
  wire       [31:0]   _zz_21575;
  wire       [15:0]   _zz_21576;
  wire       [15:0]   _zz_21577;
  wire       [31:0]   _zz_21578;
  wire       [31:0]   _zz_21579;
  wire       [15:0]   _zz_21580;
  wire       [31:0]   _zz_21581;
  wire       [31:0]   _zz_21582;
  wire       [31:0]   _zz_21583;
  wire       [15:0]   _zz_21584;
  wire       [31:0]   _zz_21585;
  wire       [31:0]   _zz_21586;
  wire       [31:0]   _zz_21587;
  wire       [31:0]   _zz_21588;
  wire       [31:0]   _zz_21589;
  wire       [31:0]   _zz_21590;
  wire       [23:0]   _zz_21591;
  wire       [31:0]   _zz_21592;
  wire       [15:0]   _zz_21593;
  wire       [31:0]   _zz_21594;
  wire       [31:0]   _zz_21595;
  wire       [31:0]   _zz_21596;
  wire       [31:0]   _zz_21597;
  wire       [31:0]   _zz_21598;
  wire       [23:0]   _zz_21599;
  wire       [31:0]   _zz_21600;
  wire       [15:0]   _zz_21601;
  wire       [31:0]   _zz_21602;
  wire       [31:0]   _zz_21603;
  wire       [31:0]   _zz_21604;
  wire       [31:0]   _zz_21605;
  wire       [31:0]   _zz_21606;
  wire       [23:0]   _zz_21607;
  wire       [31:0]   _zz_21608;
  wire       [15:0]   _zz_21609;
  wire       [31:0]   _zz_21610;
  wire       [31:0]   _zz_21611;
  wire       [31:0]   _zz_21612;
  wire       [31:0]   _zz_21613;
  wire       [31:0]   _zz_21614;
  wire       [23:0]   _zz_21615;
  wire       [31:0]   _zz_21616;
  wire       [15:0]   _zz_21617;
  wire       [15:0]   _zz_21618;
  wire       [31:0]   _zz_21619;
  wire       [31:0]   _zz_21620;
  wire       [15:0]   _zz_21621;
  wire       [31:0]   _zz_21622;
  wire       [31:0]   _zz_21623;
  wire       [31:0]   _zz_21624;
  wire       [15:0]   _zz_21625;
  wire       [31:0]   _zz_21626;
  wire       [31:0]   _zz_21627;
  wire       [31:0]   _zz_21628;
  wire       [31:0]   _zz_21629;
  wire       [31:0]   _zz_21630;
  wire       [31:0]   _zz_21631;
  wire       [23:0]   _zz_21632;
  wire       [31:0]   _zz_21633;
  wire       [15:0]   _zz_21634;
  wire       [31:0]   _zz_21635;
  wire       [31:0]   _zz_21636;
  wire       [31:0]   _zz_21637;
  wire       [31:0]   _zz_21638;
  wire       [31:0]   _zz_21639;
  wire       [23:0]   _zz_21640;
  wire       [31:0]   _zz_21641;
  wire       [15:0]   _zz_21642;
  wire       [31:0]   _zz_21643;
  wire       [31:0]   _zz_21644;
  wire       [31:0]   _zz_21645;
  wire       [31:0]   _zz_21646;
  wire       [31:0]   _zz_21647;
  wire       [23:0]   _zz_21648;
  wire       [31:0]   _zz_21649;
  wire       [15:0]   _zz_21650;
  wire       [31:0]   _zz_21651;
  wire       [31:0]   _zz_21652;
  wire       [31:0]   _zz_21653;
  wire       [31:0]   _zz_21654;
  wire       [31:0]   _zz_21655;
  wire       [23:0]   _zz_21656;
  wire       [31:0]   _zz_21657;
  wire       [15:0]   _zz_21658;
  wire       [15:0]   _zz_21659;
  wire       [31:0]   _zz_21660;
  wire       [31:0]   _zz_21661;
  wire       [15:0]   _zz_21662;
  wire       [31:0]   _zz_21663;
  wire       [31:0]   _zz_21664;
  wire       [31:0]   _zz_21665;
  wire       [15:0]   _zz_21666;
  wire       [31:0]   _zz_21667;
  wire       [31:0]   _zz_21668;
  wire       [31:0]   _zz_21669;
  wire       [31:0]   _zz_21670;
  wire       [31:0]   _zz_21671;
  wire       [31:0]   _zz_21672;
  wire       [23:0]   _zz_21673;
  wire       [31:0]   _zz_21674;
  wire       [15:0]   _zz_21675;
  wire       [31:0]   _zz_21676;
  wire       [31:0]   _zz_21677;
  wire       [31:0]   _zz_21678;
  wire       [31:0]   _zz_21679;
  wire       [31:0]   _zz_21680;
  wire       [23:0]   _zz_21681;
  wire       [31:0]   _zz_21682;
  wire       [15:0]   _zz_21683;
  wire       [31:0]   _zz_21684;
  wire       [31:0]   _zz_21685;
  wire       [31:0]   _zz_21686;
  wire       [31:0]   _zz_21687;
  wire       [31:0]   _zz_21688;
  wire       [23:0]   _zz_21689;
  wire       [31:0]   _zz_21690;
  wire       [15:0]   _zz_21691;
  wire       [31:0]   _zz_21692;
  wire       [31:0]   _zz_21693;
  wire       [31:0]   _zz_21694;
  wire       [31:0]   _zz_21695;
  wire       [31:0]   _zz_21696;
  wire       [23:0]   _zz_21697;
  wire       [31:0]   _zz_21698;
  wire       [15:0]   _zz_21699;
  wire       [15:0]   _zz_21700;
  wire       [31:0]   _zz_21701;
  wire       [31:0]   _zz_21702;
  wire       [15:0]   _zz_21703;
  wire       [31:0]   _zz_21704;
  wire       [31:0]   _zz_21705;
  wire       [31:0]   _zz_21706;
  wire       [15:0]   _zz_21707;
  wire       [31:0]   _zz_21708;
  wire       [31:0]   _zz_21709;
  wire       [31:0]   _zz_21710;
  wire       [31:0]   _zz_21711;
  wire       [31:0]   _zz_21712;
  wire       [31:0]   _zz_21713;
  wire       [23:0]   _zz_21714;
  wire       [31:0]   _zz_21715;
  wire       [15:0]   _zz_21716;
  wire       [31:0]   _zz_21717;
  wire       [31:0]   _zz_21718;
  wire       [31:0]   _zz_21719;
  wire       [31:0]   _zz_21720;
  wire       [31:0]   _zz_21721;
  wire       [23:0]   _zz_21722;
  wire       [31:0]   _zz_21723;
  wire       [15:0]   _zz_21724;
  wire       [31:0]   _zz_21725;
  wire       [31:0]   _zz_21726;
  wire       [31:0]   _zz_21727;
  wire       [31:0]   _zz_21728;
  wire       [31:0]   _zz_21729;
  wire       [23:0]   _zz_21730;
  wire       [31:0]   _zz_21731;
  wire       [15:0]   _zz_21732;
  wire       [31:0]   _zz_21733;
  wire       [31:0]   _zz_21734;
  wire       [31:0]   _zz_21735;
  wire       [31:0]   _zz_21736;
  wire       [31:0]   _zz_21737;
  wire       [23:0]   _zz_21738;
  wire       [31:0]   _zz_21739;
  wire       [15:0]   _zz_21740;
  wire       [15:0]   _zz_21741;
  wire       [31:0]   _zz_21742;
  wire       [31:0]   _zz_21743;
  wire       [15:0]   _zz_21744;
  wire       [31:0]   _zz_21745;
  wire       [31:0]   _zz_21746;
  wire       [31:0]   _zz_21747;
  wire       [15:0]   _zz_21748;
  wire       [31:0]   _zz_21749;
  wire       [31:0]   _zz_21750;
  wire       [31:0]   _zz_21751;
  wire       [31:0]   _zz_21752;
  wire       [31:0]   _zz_21753;
  wire       [31:0]   _zz_21754;
  wire       [23:0]   _zz_21755;
  wire       [31:0]   _zz_21756;
  wire       [15:0]   _zz_21757;
  wire       [31:0]   _zz_21758;
  wire       [31:0]   _zz_21759;
  wire       [31:0]   _zz_21760;
  wire       [31:0]   _zz_21761;
  wire       [31:0]   _zz_21762;
  wire       [23:0]   _zz_21763;
  wire       [31:0]   _zz_21764;
  wire       [15:0]   _zz_21765;
  wire       [31:0]   _zz_21766;
  wire       [31:0]   _zz_21767;
  wire       [31:0]   _zz_21768;
  wire       [31:0]   _zz_21769;
  wire       [31:0]   _zz_21770;
  wire       [23:0]   _zz_21771;
  wire       [31:0]   _zz_21772;
  wire       [15:0]   _zz_21773;
  wire       [31:0]   _zz_21774;
  wire       [31:0]   _zz_21775;
  wire       [31:0]   _zz_21776;
  wire       [31:0]   _zz_21777;
  wire       [31:0]   _zz_21778;
  wire       [23:0]   _zz_21779;
  wire       [31:0]   _zz_21780;
  wire       [15:0]   _zz_21781;
  wire       [15:0]   _zz_21782;
  wire       [31:0]   _zz_21783;
  wire       [31:0]   _zz_21784;
  wire       [15:0]   _zz_21785;
  wire       [31:0]   _zz_21786;
  wire       [31:0]   _zz_21787;
  wire       [31:0]   _zz_21788;
  wire       [15:0]   _zz_21789;
  wire       [31:0]   _zz_21790;
  wire       [31:0]   _zz_21791;
  wire       [31:0]   _zz_21792;
  wire       [31:0]   _zz_21793;
  wire       [31:0]   _zz_21794;
  wire       [31:0]   _zz_21795;
  wire       [23:0]   _zz_21796;
  wire       [31:0]   _zz_21797;
  wire       [15:0]   _zz_21798;
  wire       [31:0]   _zz_21799;
  wire       [31:0]   _zz_21800;
  wire       [31:0]   _zz_21801;
  wire       [31:0]   _zz_21802;
  wire       [31:0]   _zz_21803;
  wire       [23:0]   _zz_21804;
  wire       [31:0]   _zz_21805;
  wire       [15:0]   _zz_21806;
  wire       [31:0]   _zz_21807;
  wire       [31:0]   _zz_21808;
  wire       [31:0]   _zz_21809;
  wire       [31:0]   _zz_21810;
  wire       [31:0]   _zz_21811;
  wire       [23:0]   _zz_21812;
  wire       [31:0]   _zz_21813;
  wire       [15:0]   _zz_21814;
  wire       [31:0]   _zz_21815;
  wire       [31:0]   _zz_21816;
  wire       [31:0]   _zz_21817;
  wire       [31:0]   _zz_21818;
  wire       [31:0]   _zz_21819;
  wire       [23:0]   _zz_21820;
  wire       [31:0]   _zz_21821;
  wire       [15:0]   _zz_21822;
  wire       [15:0]   _zz_21823;
  wire       [31:0]   _zz_21824;
  wire       [31:0]   _zz_21825;
  wire       [15:0]   _zz_21826;
  wire       [31:0]   _zz_21827;
  wire       [31:0]   _zz_21828;
  wire       [31:0]   _zz_21829;
  wire       [15:0]   _zz_21830;
  wire       [31:0]   _zz_21831;
  wire       [31:0]   _zz_21832;
  wire       [31:0]   _zz_21833;
  wire       [31:0]   _zz_21834;
  wire       [31:0]   _zz_21835;
  wire       [31:0]   _zz_21836;
  wire       [23:0]   _zz_21837;
  wire       [31:0]   _zz_21838;
  wire       [15:0]   _zz_21839;
  wire       [31:0]   _zz_21840;
  wire       [31:0]   _zz_21841;
  wire       [31:0]   _zz_21842;
  wire       [31:0]   _zz_21843;
  wire       [31:0]   _zz_21844;
  wire       [23:0]   _zz_21845;
  wire       [31:0]   _zz_21846;
  wire       [15:0]   _zz_21847;
  wire       [31:0]   _zz_21848;
  wire       [31:0]   _zz_21849;
  wire       [31:0]   _zz_21850;
  wire       [31:0]   _zz_21851;
  wire       [31:0]   _zz_21852;
  wire       [23:0]   _zz_21853;
  wire       [31:0]   _zz_21854;
  wire       [15:0]   _zz_21855;
  wire       [31:0]   _zz_21856;
  wire       [31:0]   _zz_21857;
  wire       [31:0]   _zz_21858;
  wire       [31:0]   _zz_21859;
  wire       [31:0]   _zz_21860;
  wire       [23:0]   _zz_21861;
  wire       [31:0]   _zz_21862;
  wire       [15:0]   _zz_21863;
  wire       [15:0]   _zz_21864;
  wire       [31:0]   _zz_21865;
  wire       [31:0]   _zz_21866;
  wire       [15:0]   _zz_21867;
  wire       [31:0]   _zz_21868;
  wire       [31:0]   _zz_21869;
  wire       [31:0]   _zz_21870;
  wire       [15:0]   _zz_21871;
  wire       [31:0]   _zz_21872;
  wire       [31:0]   _zz_21873;
  wire       [31:0]   _zz_21874;
  wire       [31:0]   _zz_21875;
  wire       [31:0]   _zz_21876;
  wire       [31:0]   _zz_21877;
  wire       [23:0]   _zz_21878;
  wire       [31:0]   _zz_21879;
  wire       [15:0]   _zz_21880;
  wire       [31:0]   _zz_21881;
  wire       [31:0]   _zz_21882;
  wire       [31:0]   _zz_21883;
  wire       [31:0]   _zz_21884;
  wire       [31:0]   _zz_21885;
  wire       [23:0]   _zz_21886;
  wire       [31:0]   _zz_21887;
  wire       [15:0]   _zz_21888;
  wire       [31:0]   _zz_21889;
  wire       [31:0]   _zz_21890;
  wire       [31:0]   _zz_21891;
  wire       [31:0]   _zz_21892;
  wire       [31:0]   _zz_21893;
  wire       [23:0]   _zz_21894;
  wire       [31:0]   _zz_21895;
  wire       [15:0]   _zz_21896;
  wire       [31:0]   _zz_21897;
  wire       [31:0]   _zz_21898;
  wire       [31:0]   _zz_21899;
  wire       [31:0]   _zz_21900;
  wire       [31:0]   _zz_21901;
  wire       [23:0]   _zz_21902;
  wire       [31:0]   _zz_21903;
  wire       [15:0]   _zz_21904;
  wire       [15:0]   _zz_21905;
  wire       [31:0]   _zz_21906;
  wire       [31:0]   _zz_21907;
  wire       [15:0]   _zz_21908;
  wire       [31:0]   _zz_21909;
  wire       [31:0]   _zz_21910;
  wire       [31:0]   _zz_21911;
  wire       [15:0]   _zz_21912;
  wire       [31:0]   _zz_21913;
  wire       [31:0]   _zz_21914;
  wire       [31:0]   _zz_21915;
  wire       [31:0]   _zz_21916;
  wire       [31:0]   _zz_21917;
  wire       [31:0]   _zz_21918;
  wire       [23:0]   _zz_21919;
  wire       [31:0]   _zz_21920;
  wire       [15:0]   _zz_21921;
  wire       [31:0]   _zz_21922;
  wire       [31:0]   _zz_21923;
  wire       [31:0]   _zz_21924;
  wire       [31:0]   _zz_21925;
  wire       [31:0]   _zz_21926;
  wire       [23:0]   _zz_21927;
  wire       [31:0]   _zz_21928;
  wire       [15:0]   _zz_21929;
  wire       [31:0]   _zz_21930;
  wire       [31:0]   _zz_21931;
  wire       [31:0]   _zz_21932;
  wire       [31:0]   _zz_21933;
  wire       [31:0]   _zz_21934;
  wire       [23:0]   _zz_21935;
  wire       [31:0]   _zz_21936;
  wire       [15:0]   _zz_21937;
  wire       [31:0]   _zz_21938;
  wire       [31:0]   _zz_21939;
  wire       [31:0]   _zz_21940;
  wire       [31:0]   _zz_21941;
  wire       [31:0]   _zz_21942;
  wire       [23:0]   _zz_21943;
  wire       [31:0]   _zz_21944;
  wire       [15:0]   _zz_21945;
  wire       [15:0]   _zz_21946;
  wire       [31:0]   _zz_21947;
  wire       [31:0]   _zz_21948;
  wire       [15:0]   _zz_21949;
  wire       [31:0]   _zz_21950;
  wire       [31:0]   _zz_21951;
  wire       [31:0]   _zz_21952;
  wire       [15:0]   _zz_21953;
  wire       [31:0]   _zz_21954;
  wire       [31:0]   _zz_21955;
  wire       [31:0]   _zz_21956;
  wire       [31:0]   _zz_21957;
  wire       [31:0]   _zz_21958;
  wire       [31:0]   _zz_21959;
  wire       [23:0]   _zz_21960;
  wire       [31:0]   _zz_21961;
  wire       [15:0]   _zz_21962;
  wire       [31:0]   _zz_21963;
  wire       [31:0]   _zz_21964;
  wire       [31:0]   _zz_21965;
  wire       [31:0]   _zz_21966;
  wire       [31:0]   _zz_21967;
  wire       [23:0]   _zz_21968;
  wire       [31:0]   _zz_21969;
  wire       [15:0]   _zz_21970;
  wire       [31:0]   _zz_21971;
  wire       [31:0]   _zz_21972;
  wire       [31:0]   _zz_21973;
  wire       [31:0]   _zz_21974;
  wire       [31:0]   _zz_21975;
  wire       [23:0]   _zz_21976;
  wire       [31:0]   _zz_21977;
  wire       [15:0]   _zz_21978;
  wire       [31:0]   _zz_21979;
  wire       [31:0]   _zz_21980;
  wire       [31:0]   _zz_21981;
  wire       [31:0]   _zz_21982;
  wire       [31:0]   _zz_21983;
  wire       [23:0]   _zz_21984;
  wire       [31:0]   _zz_21985;
  wire       [15:0]   _zz_21986;
  wire       [15:0]   _zz_21987;
  wire       [31:0]   _zz_21988;
  wire       [31:0]   _zz_21989;
  wire       [15:0]   _zz_21990;
  wire       [31:0]   _zz_21991;
  wire       [31:0]   _zz_21992;
  wire       [31:0]   _zz_21993;
  wire       [15:0]   _zz_21994;
  wire       [31:0]   _zz_21995;
  wire       [31:0]   _zz_21996;
  wire       [31:0]   _zz_21997;
  wire       [31:0]   _zz_21998;
  wire       [31:0]   _zz_21999;
  wire       [31:0]   _zz_22000;
  wire       [23:0]   _zz_22001;
  wire       [31:0]   _zz_22002;
  wire       [15:0]   _zz_22003;
  wire       [31:0]   _zz_22004;
  wire       [31:0]   _zz_22005;
  wire       [31:0]   _zz_22006;
  wire       [31:0]   _zz_22007;
  wire       [31:0]   _zz_22008;
  wire       [23:0]   _zz_22009;
  wire       [31:0]   _zz_22010;
  wire       [15:0]   _zz_22011;
  wire       [31:0]   _zz_22012;
  wire       [31:0]   _zz_22013;
  wire       [31:0]   _zz_22014;
  wire       [31:0]   _zz_22015;
  wire       [31:0]   _zz_22016;
  wire       [23:0]   _zz_22017;
  wire       [31:0]   _zz_22018;
  wire       [15:0]   _zz_22019;
  wire       [31:0]   _zz_22020;
  wire       [31:0]   _zz_22021;
  wire       [31:0]   _zz_22022;
  wire       [31:0]   _zz_22023;
  wire       [31:0]   _zz_22024;
  wire       [23:0]   _zz_22025;
  wire       [31:0]   _zz_22026;
  wire       [15:0]   _zz_22027;
  wire       [15:0]   _zz_22028;
  wire       [31:0]   _zz_22029;
  wire       [31:0]   _zz_22030;
  wire       [15:0]   _zz_22031;
  wire       [31:0]   _zz_22032;
  wire       [31:0]   _zz_22033;
  wire       [31:0]   _zz_22034;
  wire       [15:0]   _zz_22035;
  wire       [31:0]   _zz_22036;
  wire       [31:0]   _zz_22037;
  wire       [31:0]   _zz_22038;
  wire       [31:0]   _zz_22039;
  wire       [31:0]   _zz_22040;
  wire       [31:0]   _zz_22041;
  wire       [23:0]   _zz_22042;
  wire       [31:0]   _zz_22043;
  wire       [15:0]   _zz_22044;
  wire       [31:0]   _zz_22045;
  wire       [31:0]   _zz_22046;
  wire       [31:0]   _zz_22047;
  wire       [31:0]   _zz_22048;
  wire       [31:0]   _zz_22049;
  wire       [23:0]   _zz_22050;
  wire       [31:0]   _zz_22051;
  wire       [15:0]   _zz_22052;
  wire       [31:0]   _zz_22053;
  wire       [31:0]   _zz_22054;
  wire       [31:0]   _zz_22055;
  wire       [31:0]   _zz_22056;
  wire       [31:0]   _zz_22057;
  wire       [23:0]   _zz_22058;
  wire       [31:0]   _zz_22059;
  wire       [15:0]   _zz_22060;
  wire       [31:0]   _zz_22061;
  wire       [31:0]   _zz_22062;
  wire       [31:0]   _zz_22063;
  wire       [31:0]   _zz_22064;
  wire       [31:0]   _zz_22065;
  wire       [23:0]   _zz_22066;
  wire       [31:0]   _zz_22067;
  wire       [15:0]   _zz_22068;
  wire       [15:0]   _zz_22069;
  wire       [31:0]   _zz_22070;
  wire       [31:0]   _zz_22071;
  wire       [15:0]   _zz_22072;
  wire       [31:0]   _zz_22073;
  wire       [31:0]   _zz_22074;
  wire       [31:0]   _zz_22075;
  wire       [15:0]   _zz_22076;
  wire       [31:0]   _zz_22077;
  wire       [31:0]   _zz_22078;
  wire       [31:0]   _zz_22079;
  wire       [31:0]   _zz_22080;
  wire       [31:0]   _zz_22081;
  wire       [31:0]   _zz_22082;
  wire       [23:0]   _zz_22083;
  wire       [31:0]   _zz_22084;
  wire       [15:0]   _zz_22085;
  wire       [31:0]   _zz_22086;
  wire       [31:0]   _zz_22087;
  wire       [31:0]   _zz_22088;
  wire       [31:0]   _zz_22089;
  wire       [31:0]   _zz_22090;
  wire       [23:0]   _zz_22091;
  wire       [31:0]   _zz_22092;
  wire       [15:0]   _zz_22093;
  wire       [31:0]   _zz_22094;
  wire       [31:0]   _zz_22095;
  wire       [31:0]   _zz_22096;
  wire       [31:0]   _zz_22097;
  wire       [31:0]   _zz_22098;
  wire       [23:0]   _zz_22099;
  wire       [31:0]   _zz_22100;
  wire       [15:0]   _zz_22101;
  wire       [31:0]   _zz_22102;
  wire       [31:0]   _zz_22103;
  wire       [31:0]   _zz_22104;
  wire       [31:0]   _zz_22105;
  wire       [31:0]   _zz_22106;
  wire       [23:0]   _zz_22107;
  wire       [31:0]   _zz_22108;
  wire       [15:0]   _zz_22109;
  wire       [15:0]   _zz_22110;
  wire       [31:0]   _zz_22111;
  wire       [31:0]   _zz_22112;
  wire       [15:0]   _zz_22113;
  wire       [31:0]   _zz_22114;
  wire       [31:0]   _zz_22115;
  wire       [31:0]   _zz_22116;
  wire       [15:0]   _zz_22117;
  wire       [31:0]   _zz_22118;
  wire       [31:0]   _zz_22119;
  wire       [31:0]   _zz_22120;
  wire       [31:0]   _zz_22121;
  wire       [31:0]   _zz_22122;
  wire       [31:0]   _zz_22123;
  wire       [23:0]   _zz_22124;
  wire       [31:0]   _zz_22125;
  wire       [15:0]   _zz_22126;
  wire       [31:0]   _zz_22127;
  wire       [31:0]   _zz_22128;
  wire       [31:0]   _zz_22129;
  wire       [31:0]   _zz_22130;
  wire       [31:0]   _zz_22131;
  wire       [23:0]   _zz_22132;
  wire       [31:0]   _zz_22133;
  wire       [15:0]   _zz_22134;
  wire       [31:0]   _zz_22135;
  wire       [31:0]   _zz_22136;
  wire       [31:0]   _zz_22137;
  wire       [31:0]   _zz_22138;
  wire       [31:0]   _zz_22139;
  wire       [23:0]   _zz_22140;
  wire       [31:0]   _zz_22141;
  wire       [15:0]   _zz_22142;
  wire       [31:0]   _zz_22143;
  wire       [31:0]   _zz_22144;
  wire       [31:0]   _zz_22145;
  wire       [31:0]   _zz_22146;
  wire       [31:0]   _zz_22147;
  wire       [23:0]   _zz_22148;
  wire       [31:0]   _zz_22149;
  wire       [15:0]   _zz_22150;
  wire       [15:0]   _zz_22151;
  wire       [31:0]   _zz_22152;
  wire       [31:0]   _zz_22153;
  wire       [15:0]   _zz_22154;
  wire       [31:0]   _zz_22155;
  wire       [31:0]   _zz_22156;
  wire       [31:0]   _zz_22157;
  wire       [15:0]   _zz_22158;
  wire       [31:0]   _zz_22159;
  wire       [31:0]   _zz_22160;
  wire       [31:0]   _zz_22161;
  wire       [31:0]   _zz_22162;
  wire       [31:0]   _zz_22163;
  wire       [31:0]   _zz_22164;
  wire       [23:0]   _zz_22165;
  wire       [31:0]   _zz_22166;
  wire       [15:0]   _zz_22167;
  wire       [31:0]   _zz_22168;
  wire       [31:0]   _zz_22169;
  wire       [31:0]   _zz_22170;
  wire       [31:0]   _zz_22171;
  wire       [31:0]   _zz_22172;
  wire       [23:0]   _zz_22173;
  wire       [31:0]   _zz_22174;
  wire       [15:0]   _zz_22175;
  wire       [31:0]   _zz_22176;
  wire       [31:0]   _zz_22177;
  wire       [31:0]   _zz_22178;
  wire       [31:0]   _zz_22179;
  wire       [31:0]   _zz_22180;
  wire       [23:0]   _zz_22181;
  wire       [31:0]   _zz_22182;
  wire       [15:0]   _zz_22183;
  wire       [31:0]   _zz_22184;
  wire       [31:0]   _zz_22185;
  wire       [31:0]   _zz_22186;
  wire       [31:0]   _zz_22187;
  wire       [31:0]   _zz_22188;
  wire       [23:0]   _zz_22189;
  wire       [31:0]   _zz_22190;
  wire       [15:0]   _zz_22191;
  wire       [15:0]   _zz_22192;
  wire       [31:0]   _zz_22193;
  wire       [31:0]   _zz_22194;
  wire       [15:0]   _zz_22195;
  wire       [31:0]   _zz_22196;
  wire       [31:0]   _zz_22197;
  wire       [31:0]   _zz_22198;
  wire       [15:0]   _zz_22199;
  wire       [31:0]   _zz_22200;
  wire       [31:0]   _zz_22201;
  wire       [31:0]   _zz_22202;
  wire       [31:0]   _zz_22203;
  wire       [31:0]   _zz_22204;
  wire       [31:0]   _zz_22205;
  wire       [23:0]   _zz_22206;
  wire       [31:0]   _zz_22207;
  wire       [15:0]   _zz_22208;
  wire       [31:0]   _zz_22209;
  wire       [31:0]   _zz_22210;
  wire       [31:0]   _zz_22211;
  wire       [31:0]   _zz_22212;
  wire       [31:0]   _zz_22213;
  wire       [23:0]   _zz_22214;
  wire       [31:0]   _zz_22215;
  wire       [15:0]   _zz_22216;
  wire       [31:0]   _zz_22217;
  wire       [31:0]   _zz_22218;
  wire       [31:0]   _zz_22219;
  wire       [31:0]   _zz_22220;
  wire       [31:0]   _zz_22221;
  wire       [23:0]   _zz_22222;
  wire       [31:0]   _zz_22223;
  wire       [15:0]   _zz_22224;
  wire       [31:0]   _zz_22225;
  wire       [31:0]   _zz_22226;
  wire       [31:0]   _zz_22227;
  wire       [31:0]   _zz_22228;
  wire       [31:0]   _zz_22229;
  wire       [23:0]   _zz_22230;
  wire       [31:0]   _zz_22231;
  wire       [15:0]   _zz_22232;
  wire       [15:0]   _zz_22233;
  wire       [31:0]   _zz_22234;
  wire       [31:0]   _zz_22235;
  wire       [15:0]   _zz_22236;
  wire       [31:0]   _zz_22237;
  wire       [31:0]   _zz_22238;
  wire       [31:0]   _zz_22239;
  wire       [15:0]   _zz_22240;
  wire       [31:0]   _zz_22241;
  wire       [31:0]   _zz_22242;
  wire       [31:0]   _zz_22243;
  wire       [31:0]   _zz_22244;
  wire       [31:0]   _zz_22245;
  wire       [31:0]   _zz_22246;
  wire       [23:0]   _zz_22247;
  wire       [31:0]   _zz_22248;
  wire       [15:0]   _zz_22249;
  wire       [31:0]   _zz_22250;
  wire       [31:0]   _zz_22251;
  wire       [31:0]   _zz_22252;
  wire       [31:0]   _zz_22253;
  wire       [31:0]   _zz_22254;
  wire       [23:0]   _zz_22255;
  wire       [31:0]   _zz_22256;
  wire       [15:0]   _zz_22257;
  wire       [31:0]   _zz_22258;
  wire       [31:0]   _zz_22259;
  wire       [31:0]   _zz_22260;
  wire       [31:0]   _zz_22261;
  wire       [31:0]   _zz_22262;
  wire       [23:0]   _zz_22263;
  wire       [31:0]   _zz_22264;
  wire       [15:0]   _zz_22265;
  wire       [31:0]   _zz_22266;
  wire       [31:0]   _zz_22267;
  wire       [31:0]   _zz_22268;
  wire       [31:0]   _zz_22269;
  wire       [31:0]   _zz_22270;
  wire       [23:0]   _zz_22271;
  wire       [31:0]   _zz_22272;
  wire       [15:0]   _zz_22273;
  wire       [15:0]   _zz_22274;
  wire       [31:0]   _zz_22275;
  wire       [31:0]   _zz_22276;
  wire       [15:0]   _zz_22277;
  wire       [31:0]   _zz_22278;
  wire       [31:0]   _zz_22279;
  wire       [31:0]   _zz_22280;
  wire       [15:0]   _zz_22281;
  wire       [31:0]   _zz_22282;
  wire       [31:0]   _zz_22283;
  wire       [31:0]   _zz_22284;
  wire       [31:0]   _zz_22285;
  wire       [31:0]   _zz_22286;
  wire       [31:0]   _zz_22287;
  wire       [23:0]   _zz_22288;
  wire       [31:0]   _zz_22289;
  wire       [15:0]   _zz_22290;
  wire       [31:0]   _zz_22291;
  wire       [31:0]   _zz_22292;
  wire       [31:0]   _zz_22293;
  wire       [31:0]   _zz_22294;
  wire       [31:0]   _zz_22295;
  wire       [23:0]   _zz_22296;
  wire       [31:0]   _zz_22297;
  wire       [15:0]   _zz_22298;
  wire       [31:0]   _zz_22299;
  wire       [31:0]   _zz_22300;
  wire       [31:0]   _zz_22301;
  wire       [31:0]   _zz_22302;
  wire       [31:0]   _zz_22303;
  wire       [23:0]   _zz_22304;
  wire       [31:0]   _zz_22305;
  wire       [15:0]   _zz_22306;
  wire       [31:0]   _zz_22307;
  wire       [31:0]   _zz_22308;
  wire       [31:0]   _zz_22309;
  wire       [31:0]   _zz_22310;
  wire       [31:0]   _zz_22311;
  wire       [23:0]   _zz_22312;
  wire       [31:0]   _zz_22313;
  wire       [15:0]   _zz_22314;
  wire       [15:0]   _zz_22315;
  wire       [31:0]   _zz_22316;
  wire       [31:0]   _zz_22317;
  wire       [15:0]   _zz_22318;
  wire       [31:0]   _zz_22319;
  wire       [31:0]   _zz_22320;
  wire       [31:0]   _zz_22321;
  wire       [15:0]   _zz_22322;
  wire       [31:0]   _zz_22323;
  wire       [31:0]   _zz_22324;
  wire       [31:0]   _zz_22325;
  wire       [31:0]   _zz_22326;
  wire       [31:0]   _zz_22327;
  wire       [31:0]   _zz_22328;
  wire       [23:0]   _zz_22329;
  wire       [31:0]   _zz_22330;
  wire       [15:0]   _zz_22331;
  wire       [31:0]   _zz_22332;
  wire       [31:0]   _zz_22333;
  wire       [31:0]   _zz_22334;
  wire       [31:0]   _zz_22335;
  wire       [31:0]   _zz_22336;
  wire       [23:0]   _zz_22337;
  wire       [31:0]   _zz_22338;
  wire       [15:0]   _zz_22339;
  wire       [31:0]   _zz_22340;
  wire       [31:0]   _zz_22341;
  wire       [31:0]   _zz_22342;
  wire       [31:0]   _zz_22343;
  wire       [31:0]   _zz_22344;
  wire       [23:0]   _zz_22345;
  wire       [31:0]   _zz_22346;
  wire       [15:0]   _zz_22347;
  wire       [31:0]   _zz_22348;
  wire       [31:0]   _zz_22349;
  wire       [31:0]   _zz_22350;
  wire       [31:0]   _zz_22351;
  wire       [31:0]   _zz_22352;
  wire       [23:0]   _zz_22353;
  wire       [31:0]   _zz_22354;
  wire       [15:0]   _zz_22355;
  wire       [15:0]   _zz_22356;
  wire       [31:0]   _zz_22357;
  wire       [31:0]   _zz_22358;
  wire       [15:0]   _zz_22359;
  wire       [31:0]   _zz_22360;
  wire       [31:0]   _zz_22361;
  wire       [31:0]   _zz_22362;
  wire       [15:0]   _zz_22363;
  wire       [31:0]   _zz_22364;
  wire       [31:0]   _zz_22365;
  wire       [31:0]   _zz_22366;
  wire       [31:0]   _zz_22367;
  wire       [31:0]   _zz_22368;
  wire       [31:0]   _zz_22369;
  wire       [23:0]   _zz_22370;
  wire       [31:0]   _zz_22371;
  wire       [15:0]   _zz_22372;
  wire       [31:0]   _zz_22373;
  wire       [31:0]   _zz_22374;
  wire       [31:0]   _zz_22375;
  wire       [31:0]   _zz_22376;
  wire       [31:0]   _zz_22377;
  wire       [23:0]   _zz_22378;
  wire       [31:0]   _zz_22379;
  wire       [15:0]   _zz_22380;
  wire       [31:0]   _zz_22381;
  wire       [31:0]   _zz_22382;
  wire       [31:0]   _zz_22383;
  wire       [31:0]   _zz_22384;
  wire       [31:0]   _zz_22385;
  wire       [23:0]   _zz_22386;
  wire       [31:0]   _zz_22387;
  wire       [15:0]   _zz_22388;
  wire       [31:0]   _zz_22389;
  wire       [31:0]   _zz_22390;
  wire       [31:0]   _zz_22391;
  wire       [31:0]   _zz_22392;
  wire       [31:0]   _zz_22393;
  wire       [23:0]   _zz_22394;
  wire       [31:0]   _zz_22395;
  wire       [15:0]   _zz_22396;
  wire       [15:0]   _zz_22397;
  wire       [31:0]   _zz_22398;
  wire       [31:0]   _zz_22399;
  wire       [15:0]   _zz_22400;
  wire       [31:0]   _zz_22401;
  wire       [31:0]   _zz_22402;
  wire       [31:0]   _zz_22403;
  wire       [15:0]   _zz_22404;
  wire       [31:0]   _zz_22405;
  wire       [31:0]   _zz_22406;
  wire       [31:0]   _zz_22407;
  wire       [31:0]   _zz_22408;
  wire       [31:0]   _zz_22409;
  wire       [31:0]   _zz_22410;
  wire       [23:0]   _zz_22411;
  wire       [31:0]   _zz_22412;
  wire       [15:0]   _zz_22413;
  wire       [31:0]   _zz_22414;
  wire       [31:0]   _zz_22415;
  wire       [31:0]   _zz_22416;
  wire       [31:0]   _zz_22417;
  wire       [31:0]   _zz_22418;
  wire       [23:0]   _zz_22419;
  wire       [31:0]   _zz_22420;
  wire       [15:0]   _zz_22421;
  wire       [31:0]   _zz_22422;
  wire       [31:0]   _zz_22423;
  wire       [31:0]   _zz_22424;
  wire       [31:0]   _zz_22425;
  wire       [31:0]   _zz_22426;
  wire       [23:0]   _zz_22427;
  wire       [31:0]   _zz_22428;
  wire       [15:0]   _zz_22429;
  wire       [31:0]   _zz_22430;
  wire       [31:0]   _zz_22431;
  wire       [31:0]   _zz_22432;
  wire       [31:0]   _zz_22433;
  wire       [31:0]   _zz_22434;
  wire       [23:0]   _zz_22435;
  wire       [31:0]   _zz_22436;
  wire       [15:0]   _zz_22437;
  wire       [15:0]   _zz_22438;
  wire       [31:0]   _zz_22439;
  wire       [31:0]   _zz_22440;
  wire       [15:0]   _zz_22441;
  wire       [31:0]   _zz_22442;
  wire       [31:0]   _zz_22443;
  wire       [31:0]   _zz_22444;
  wire       [15:0]   _zz_22445;
  wire       [31:0]   _zz_22446;
  wire       [31:0]   _zz_22447;
  wire       [31:0]   _zz_22448;
  wire       [31:0]   _zz_22449;
  wire       [31:0]   _zz_22450;
  wire       [31:0]   _zz_22451;
  wire       [23:0]   _zz_22452;
  wire       [31:0]   _zz_22453;
  wire       [15:0]   _zz_22454;
  wire       [31:0]   _zz_22455;
  wire       [31:0]   _zz_22456;
  wire       [31:0]   _zz_22457;
  wire       [31:0]   _zz_22458;
  wire       [31:0]   _zz_22459;
  wire       [23:0]   _zz_22460;
  wire       [31:0]   _zz_22461;
  wire       [15:0]   _zz_22462;
  wire       [31:0]   _zz_22463;
  wire       [31:0]   _zz_22464;
  wire       [31:0]   _zz_22465;
  wire       [31:0]   _zz_22466;
  wire       [31:0]   _zz_22467;
  wire       [23:0]   _zz_22468;
  wire       [31:0]   _zz_22469;
  wire       [15:0]   _zz_22470;
  wire       [31:0]   _zz_22471;
  wire       [31:0]   _zz_22472;
  wire       [31:0]   _zz_22473;
  wire       [31:0]   _zz_22474;
  wire       [31:0]   _zz_22475;
  wire       [23:0]   _zz_22476;
  wire       [31:0]   _zz_22477;
  wire       [15:0]   _zz_22478;
  wire       [15:0]   _zz_22479;
  wire       [31:0]   _zz_22480;
  wire       [31:0]   _zz_22481;
  wire       [15:0]   _zz_22482;
  wire       [31:0]   _zz_22483;
  wire       [31:0]   _zz_22484;
  wire       [31:0]   _zz_22485;
  wire       [15:0]   _zz_22486;
  wire       [31:0]   _zz_22487;
  wire       [31:0]   _zz_22488;
  wire       [31:0]   _zz_22489;
  wire       [31:0]   _zz_22490;
  wire       [31:0]   _zz_22491;
  wire       [31:0]   _zz_22492;
  wire       [23:0]   _zz_22493;
  wire       [31:0]   _zz_22494;
  wire       [15:0]   _zz_22495;
  wire       [31:0]   _zz_22496;
  wire       [31:0]   _zz_22497;
  wire       [31:0]   _zz_22498;
  wire       [31:0]   _zz_22499;
  wire       [31:0]   _zz_22500;
  wire       [23:0]   _zz_22501;
  wire       [31:0]   _zz_22502;
  wire       [15:0]   _zz_22503;
  wire       [31:0]   _zz_22504;
  wire       [31:0]   _zz_22505;
  wire       [31:0]   _zz_22506;
  wire       [31:0]   _zz_22507;
  wire       [31:0]   _zz_22508;
  wire       [23:0]   _zz_22509;
  wire       [31:0]   _zz_22510;
  wire       [15:0]   _zz_22511;
  wire       [31:0]   _zz_22512;
  wire       [31:0]   _zz_22513;
  wire       [31:0]   _zz_22514;
  wire       [31:0]   _zz_22515;
  wire       [31:0]   _zz_22516;
  wire       [23:0]   _zz_22517;
  wire       [31:0]   _zz_22518;
  wire       [15:0]   _zz_22519;
  wire       [15:0]   _zz_22520;
  wire       [31:0]   _zz_22521;
  wire       [31:0]   _zz_22522;
  wire       [15:0]   _zz_22523;
  wire       [31:0]   _zz_22524;
  wire       [31:0]   _zz_22525;
  wire       [31:0]   _zz_22526;
  wire       [15:0]   _zz_22527;
  wire       [31:0]   _zz_22528;
  wire       [31:0]   _zz_22529;
  wire       [31:0]   _zz_22530;
  wire       [31:0]   _zz_22531;
  wire       [31:0]   _zz_22532;
  wire       [31:0]   _zz_22533;
  wire       [23:0]   _zz_22534;
  wire       [31:0]   _zz_22535;
  wire       [15:0]   _zz_22536;
  wire       [31:0]   _zz_22537;
  wire       [31:0]   _zz_22538;
  wire       [31:0]   _zz_22539;
  wire       [31:0]   _zz_22540;
  wire       [31:0]   _zz_22541;
  wire       [23:0]   _zz_22542;
  wire       [31:0]   _zz_22543;
  wire       [15:0]   _zz_22544;
  wire       [31:0]   _zz_22545;
  wire       [31:0]   _zz_22546;
  wire       [31:0]   _zz_22547;
  wire       [31:0]   _zz_22548;
  wire       [31:0]   _zz_22549;
  wire       [23:0]   _zz_22550;
  wire       [31:0]   _zz_22551;
  wire       [15:0]   _zz_22552;
  wire       [31:0]   _zz_22553;
  wire       [31:0]   _zz_22554;
  wire       [31:0]   _zz_22555;
  wire       [31:0]   _zz_22556;
  wire       [31:0]   _zz_22557;
  wire       [23:0]   _zz_22558;
  wire       [31:0]   _zz_22559;
  wire       [15:0]   _zz_22560;
  wire       [15:0]   _zz_22561;
  wire       [31:0]   _zz_22562;
  wire       [31:0]   _zz_22563;
  wire       [15:0]   _zz_22564;
  wire       [31:0]   _zz_22565;
  wire       [31:0]   _zz_22566;
  wire       [31:0]   _zz_22567;
  wire       [15:0]   _zz_22568;
  wire       [31:0]   _zz_22569;
  wire       [31:0]   _zz_22570;
  wire       [31:0]   _zz_22571;
  wire       [31:0]   _zz_22572;
  wire       [31:0]   _zz_22573;
  wire       [31:0]   _zz_22574;
  wire       [23:0]   _zz_22575;
  wire       [31:0]   _zz_22576;
  wire       [15:0]   _zz_22577;
  wire       [31:0]   _zz_22578;
  wire       [31:0]   _zz_22579;
  wire       [31:0]   _zz_22580;
  wire       [31:0]   _zz_22581;
  wire       [31:0]   _zz_22582;
  wire       [23:0]   _zz_22583;
  wire       [31:0]   _zz_22584;
  wire       [15:0]   _zz_22585;
  wire       [31:0]   _zz_22586;
  wire       [31:0]   _zz_22587;
  wire       [31:0]   _zz_22588;
  wire       [31:0]   _zz_22589;
  wire       [31:0]   _zz_22590;
  wire       [23:0]   _zz_22591;
  wire       [31:0]   _zz_22592;
  wire       [15:0]   _zz_22593;
  wire       [31:0]   _zz_22594;
  wire       [31:0]   _zz_22595;
  wire       [31:0]   _zz_22596;
  wire       [31:0]   _zz_22597;
  wire       [31:0]   _zz_22598;
  wire       [23:0]   _zz_22599;
  wire       [31:0]   _zz_22600;
  wire       [15:0]   _zz_22601;
  wire       [15:0]   _zz_22602;
  wire       [31:0]   _zz_22603;
  wire       [31:0]   _zz_22604;
  wire       [15:0]   _zz_22605;
  wire       [31:0]   _zz_22606;
  wire       [31:0]   _zz_22607;
  wire       [31:0]   _zz_22608;
  wire       [15:0]   _zz_22609;
  wire       [31:0]   _zz_22610;
  wire       [31:0]   _zz_22611;
  wire       [31:0]   _zz_22612;
  wire       [31:0]   _zz_22613;
  wire       [31:0]   _zz_22614;
  wire       [31:0]   _zz_22615;
  wire       [23:0]   _zz_22616;
  wire       [31:0]   _zz_22617;
  wire       [15:0]   _zz_22618;
  wire       [31:0]   _zz_22619;
  wire       [31:0]   _zz_22620;
  wire       [31:0]   _zz_22621;
  wire       [31:0]   _zz_22622;
  wire       [31:0]   _zz_22623;
  wire       [23:0]   _zz_22624;
  wire       [31:0]   _zz_22625;
  wire       [15:0]   _zz_22626;
  wire       [31:0]   _zz_22627;
  wire       [31:0]   _zz_22628;
  wire       [31:0]   _zz_22629;
  wire       [31:0]   _zz_22630;
  wire       [31:0]   _zz_22631;
  wire       [23:0]   _zz_22632;
  wire       [31:0]   _zz_22633;
  wire       [15:0]   _zz_22634;
  wire       [31:0]   _zz_22635;
  wire       [31:0]   _zz_22636;
  wire       [31:0]   _zz_22637;
  wire       [31:0]   _zz_22638;
  wire       [31:0]   _zz_22639;
  wire       [23:0]   _zz_22640;
  wire       [31:0]   _zz_22641;
  wire       [15:0]   _zz_22642;
  wire       [15:0]   _zz_22643;
  wire       [31:0]   _zz_22644;
  wire       [31:0]   _zz_22645;
  wire       [15:0]   _zz_22646;
  wire       [31:0]   _zz_22647;
  wire       [31:0]   _zz_22648;
  wire       [31:0]   _zz_22649;
  wire       [15:0]   _zz_22650;
  wire       [31:0]   _zz_22651;
  wire       [31:0]   _zz_22652;
  wire       [31:0]   _zz_22653;
  wire       [31:0]   _zz_22654;
  wire       [31:0]   _zz_22655;
  wire       [31:0]   _zz_22656;
  wire       [23:0]   _zz_22657;
  wire       [31:0]   _zz_22658;
  wire       [15:0]   _zz_22659;
  wire       [31:0]   _zz_22660;
  wire       [31:0]   _zz_22661;
  wire       [31:0]   _zz_22662;
  wire       [31:0]   _zz_22663;
  wire       [31:0]   _zz_22664;
  wire       [23:0]   _zz_22665;
  wire       [31:0]   _zz_22666;
  wire       [15:0]   _zz_22667;
  wire       [31:0]   _zz_22668;
  wire       [31:0]   _zz_22669;
  wire       [31:0]   _zz_22670;
  wire       [31:0]   _zz_22671;
  wire       [31:0]   _zz_22672;
  wire       [23:0]   _zz_22673;
  wire       [31:0]   _zz_22674;
  wire       [15:0]   _zz_22675;
  wire       [31:0]   _zz_22676;
  wire       [31:0]   _zz_22677;
  wire       [31:0]   _zz_22678;
  wire       [31:0]   _zz_22679;
  wire       [31:0]   _zz_22680;
  wire       [23:0]   _zz_22681;
  wire       [31:0]   _zz_22682;
  wire       [15:0]   _zz_22683;
  wire       [15:0]   _zz_22684;
  wire       [31:0]   _zz_22685;
  wire       [31:0]   _zz_22686;
  wire       [15:0]   _zz_22687;
  wire       [31:0]   _zz_22688;
  wire       [31:0]   _zz_22689;
  wire       [31:0]   _zz_22690;
  wire       [15:0]   _zz_22691;
  wire       [31:0]   _zz_22692;
  wire       [31:0]   _zz_22693;
  wire       [31:0]   _zz_22694;
  wire       [31:0]   _zz_22695;
  wire       [31:0]   _zz_22696;
  wire       [31:0]   _zz_22697;
  wire       [23:0]   _zz_22698;
  wire       [31:0]   _zz_22699;
  wire       [15:0]   _zz_22700;
  wire       [31:0]   _zz_22701;
  wire       [31:0]   _zz_22702;
  wire       [31:0]   _zz_22703;
  wire       [31:0]   _zz_22704;
  wire       [31:0]   _zz_22705;
  wire       [23:0]   _zz_22706;
  wire       [31:0]   _zz_22707;
  wire       [15:0]   _zz_22708;
  wire       [31:0]   _zz_22709;
  wire       [31:0]   _zz_22710;
  wire       [31:0]   _zz_22711;
  wire       [31:0]   _zz_22712;
  wire       [31:0]   _zz_22713;
  wire       [23:0]   _zz_22714;
  wire       [31:0]   _zz_22715;
  wire       [15:0]   _zz_22716;
  wire       [31:0]   _zz_22717;
  wire       [31:0]   _zz_22718;
  wire       [31:0]   _zz_22719;
  wire       [31:0]   _zz_22720;
  wire       [31:0]   _zz_22721;
  wire       [23:0]   _zz_22722;
  wire       [31:0]   _zz_22723;
  wire       [15:0]   _zz_22724;
  wire       [15:0]   _zz_22725;
  wire       [31:0]   _zz_22726;
  wire       [31:0]   _zz_22727;
  wire       [15:0]   _zz_22728;
  wire       [31:0]   _zz_22729;
  wire       [31:0]   _zz_22730;
  wire       [31:0]   _zz_22731;
  wire       [15:0]   _zz_22732;
  wire       [31:0]   _zz_22733;
  wire       [31:0]   _zz_22734;
  wire       [31:0]   _zz_22735;
  wire       [31:0]   _zz_22736;
  wire       [31:0]   _zz_22737;
  wire       [31:0]   _zz_22738;
  wire       [23:0]   _zz_22739;
  wire       [31:0]   _zz_22740;
  wire       [15:0]   _zz_22741;
  wire       [31:0]   _zz_22742;
  wire       [31:0]   _zz_22743;
  wire       [31:0]   _zz_22744;
  wire       [31:0]   _zz_22745;
  wire       [31:0]   _zz_22746;
  wire       [23:0]   _zz_22747;
  wire       [31:0]   _zz_22748;
  wire       [15:0]   _zz_22749;
  wire       [31:0]   _zz_22750;
  wire       [31:0]   _zz_22751;
  wire       [31:0]   _zz_22752;
  wire       [31:0]   _zz_22753;
  wire       [31:0]   _zz_22754;
  wire       [23:0]   _zz_22755;
  wire       [31:0]   _zz_22756;
  wire       [15:0]   _zz_22757;
  wire       [31:0]   _zz_22758;
  wire       [31:0]   _zz_22759;
  wire       [31:0]   _zz_22760;
  wire       [31:0]   _zz_22761;
  wire       [31:0]   _zz_22762;
  wire       [23:0]   _zz_22763;
  wire       [31:0]   _zz_22764;
  wire       [15:0]   _zz_22765;
  wire       [15:0]   _zz_22766;
  wire       [31:0]   _zz_22767;
  wire       [31:0]   _zz_22768;
  wire       [15:0]   _zz_22769;
  wire       [31:0]   _zz_22770;
  wire       [31:0]   _zz_22771;
  wire       [31:0]   _zz_22772;
  wire       [15:0]   _zz_22773;
  wire       [31:0]   _zz_22774;
  wire       [31:0]   _zz_22775;
  wire       [31:0]   _zz_22776;
  wire       [31:0]   _zz_22777;
  wire       [31:0]   _zz_22778;
  wire       [31:0]   _zz_22779;
  wire       [23:0]   _zz_22780;
  wire       [31:0]   _zz_22781;
  wire       [15:0]   _zz_22782;
  wire       [31:0]   _zz_22783;
  wire       [31:0]   _zz_22784;
  wire       [31:0]   _zz_22785;
  wire       [31:0]   _zz_22786;
  wire       [31:0]   _zz_22787;
  wire       [23:0]   _zz_22788;
  wire       [31:0]   _zz_22789;
  wire       [15:0]   _zz_22790;
  wire       [31:0]   _zz_22791;
  wire       [31:0]   _zz_22792;
  wire       [31:0]   _zz_22793;
  wire       [31:0]   _zz_22794;
  wire       [31:0]   _zz_22795;
  wire       [23:0]   _zz_22796;
  wire       [31:0]   _zz_22797;
  wire       [15:0]   _zz_22798;
  wire       [31:0]   _zz_22799;
  wire       [31:0]   _zz_22800;
  wire       [31:0]   _zz_22801;
  wire       [31:0]   _zz_22802;
  wire       [31:0]   _zz_22803;
  wire       [23:0]   _zz_22804;
  wire       [31:0]   _zz_22805;
  wire       [15:0]   _zz_22806;
  wire       [15:0]   _zz_22807;
  wire       [31:0]   _zz_22808;
  wire       [31:0]   _zz_22809;
  wire       [15:0]   _zz_22810;
  wire       [31:0]   _zz_22811;
  wire       [31:0]   _zz_22812;
  wire       [31:0]   _zz_22813;
  wire       [15:0]   _zz_22814;
  wire       [31:0]   _zz_22815;
  wire       [31:0]   _zz_22816;
  wire       [31:0]   _zz_22817;
  wire       [31:0]   _zz_22818;
  wire       [31:0]   _zz_22819;
  wire       [31:0]   _zz_22820;
  wire       [23:0]   _zz_22821;
  wire       [31:0]   _zz_22822;
  wire       [15:0]   _zz_22823;
  wire       [31:0]   _zz_22824;
  wire       [31:0]   _zz_22825;
  wire       [31:0]   _zz_22826;
  wire       [31:0]   _zz_22827;
  wire       [31:0]   _zz_22828;
  wire       [23:0]   _zz_22829;
  wire       [31:0]   _zz_22830;
  wire       [15:0]   _zz_22831;
  wire       [31:0]   _zz_22832;
  wire       [31:0]   _zz_22833;
  wire       [31:0]   _zz_22834;
  wire       [31:0]   _zz_22835;
  wire       [31:0]   _zz_22836;
  wire       [23:0]   _zz_22837;
  wire       [31:0]   _zz_22838;
  wire       [15:0]   _zz_22839;
  wire       [31:0]   _zz_22840;
  wire       [31:0]   _zz_22841;
  wire       [31:0]   _zz_22842;
  wire       [31:0]   _zz_22843;
  wire       [31:0]   _zz_22844;
  wire       [23:0]   _zz_22845;
  wire       [31:0]   _zz_22846;
  wire       [15:0]   _zz_22847;
  wire       [15:0]   _zz_22848;
  wire       [31:0]   _zz_22849;
  wire       [31:0]   _zz_22850;
  wire       [15:0]   _zz_22851;
  wire       [31:0]   _zz_22852;
  wire       [31:0]   _zz_22853;
  wire       [31:0]   _zz_22854;
  wire       [15:0]   _zz_22855;
  wire       [31:0]   _zz_22856;
  wire       [31:0]   _zz_22857;
  wire       [31:0]   _zz_22858;
  wire       [31:0]   _zz_22859;
  wire       [31:0]   _zz_22860;
  wire       [31:0]   _zz_22861;
  wire       [23:0]   _zz_22862;
  wire       [31:0]   _zz_22863;
  wire       [15:0]   _zz_22864;
  wire       [31:0]   _zz_22865;
  wire       [31:0]   _zz_22866;
  wire       [31:0]   _zz_22867;
  wire       [31:0]   _zz_22868;
  wire       [31:0]   _zz_22869;
  wire       [23:0]   _zz_22870;
  wire       [31:0]   _zz_22871;
  wire       [15:0]   _zz_22872;
  wire       [31:0]   _zz_22873;
  wire       [31:0]   _zz_22874;
  wire       [31:0]   _zz_22875;
  wire       [31:0]   _zz_22876;
  wire       [31:0]   _zz_22877;
  wire       [23:0]   _zz_22878;
  wire       [31:0]   _zz_22879;
  wire       [15:0]   _zz_22880;
  wire       [31:0]   _zz_22881;
  wire       [31:0]   _zz_22882;
  wire       [31:0]   _zz_22883;
  wire       [31:0]   _zz_22884;
  wire       [31:0]   _zz_22885;
  wire       [23:0]   _zz_22886;
  wire       [31:0]   _zz_22887;
  wire       [15:0]   _zz_22888;
  wire       [15:0]   _zz_22889;
  wire       [31:0]   _zz_22890;
  wire       [31:0]   _zz_22891;
  wire       [15:0]   _zz_22892;
  wire       [31:0]   _zz_22893;
  wire       [31:0]   _zz_22894;
  wire       [31:0]   _zz_22895;
  wire       [15:0]   _zz_22896;
  wire       [31:0]   _zz_22897;
  wire       [31:0]   _zz_22898;
  wire       [31:0]   _zz_22899;
  wire       [31:0]   _zz_22900;
  wire       [31:0]   _zz_22901;
  wire       [31:0]   _zz_22902;
  wire       [23:0]   _zz_22903;
  wire       [31:0]   _zz_22904;
  wire       [15:0]   _zz_22905;
  wire       [31:0]   _zz_22906;
  wire       [31:0]   _zz_22907;
  wire       [31:0]   _zz_22908;
  wire       [31:0]   _zz_22909;
  wire       [31:0]   _zz_22910;
  wire       [23:0]   _zz_22911;
  wire       [31:0]   _zz_22912;
  wire       [15:0]   _zz_22913;
  wire       [31:0]   _zz_22914;
  wire       [31:0]   _zz_22915;
  wire       [31:0]   _zz_22916;
  wire       [31:0]   _zz_22917;
  wire       [31:0]   _zz_22918;
  wire       [23:0]   _zz_22919;
  wire       [31:0]   _zz_22920;
  wire       [15:0]   _zz_22921;
  wire       [31:0]   _zz_22922;
  wire       [31:0]   _zz_22923;
  wire       [31:0]   _zz_22924;
  wire       [31:0]   _zz_22925;
  wire       [31:0]   _zz_22926;
  wire       [23:0]   _zz_22927;
  wire       [31:0]   _zz_22928;
  wire       [15:0]   _zz_22929;
  wire       [15:0]   _zz_22930;
  wire       [31:0]   _zz_22931;
  wire       [31:0]   _zz_22932;
  wire       [15:0]   _zz_22933;
  wire       [31:0]   _zz_22934;
  wire       [31:0]   _zz_22935;
  wire       [31:0]   _zz_22936;
  wire       [15:0]   _zz_22937;
  wire       [31:0]   _zz_22938;
  wire       [31:0]   _zz_22939;
  wire       [31:0]   _zz_22940;
  wire       [31:0]   _zz_22941;
  wire       [31:0]   _zz_22942;
  wire       [31:0]   _zz_22943;
  wire       [23:0]   _zz_22944;
  wire       [31:0]   _zz_22945;
  wire       [15:0]   _zz_22946;
  wire       [31:0]   _zz_22947;
  wire       [31:0]   _zz_22948;
  wire       [31:0]   _zz_22949;
  wire       [31:0]   _zz_22950;
  wire       [31:0]   _zz_22951;
  wire       [23:0]   _zz_22952;
  wire       [31:0]   _zz_22953;
  wire       [15:0]   _zz_22954;
  wire       [31:0]   _zz_22955;
  wire       [31:0]   _zz_22956;
  wire       [31:0]   _zz_22957;
  wire       [31:0]   _zz_22958;
  wire       [31:0]   _zz_22959;
  wire       [23:0]   _zz_22960;
  wire       [31:0]   _zz_22961;
  wire       [15:0]   _zz_22962;
  wire       [31:0]   _zz_22963;
  wire       [31:0]   _zz_22964;
  wire       [31:0]   _zz_22965;
  wire       [31:0]   _zz_22966;
  wire       [31:0]   _zz_22967;
  wire       [23:0]   _zz_22968;
  wire       [31:0]   _zz_22969;
  wire       [15:0]   _zz_22970;
  wire       [15:0]   _zz_22971;
  wire       [31:0]   _zz_22972;
  wire       [31:0]   _zz_22973;
  wire       [15:0]   _zz_22974;
  wire       [31:0]   _zz_22975;
  wire       [31:0]   _zz_22976;
  wire       [31:0]   _zz_22977;
  wire       [15:0]   _zz_22978;
  wire       [31:0]   _zz_22979;
  wire       [31:0]   _zz_22980;
  wire       [31:0]   _zz_22981;
  wire       [31:0]   _zz_22982;
  wire       [31:0]   _zz_22983;
  wire       [31:0]   _zz_22984;
  wire       [23:0]   _zz_22985;
  wire       [31:0]   _zz_22986;
  wire       [15:0]   _zz_22987;
  wire       [31:0]   _zz_22988;
  wire       [31:0]   _zz_22989;
  wire       [31:0]   _zz_22990;
  wire       [31:0]   _zz_22991;
  wire       [31:0]   _zz_22992;
  wire       [23:0]   _zz_22993;
  wire       [31:0]   _zz_22994;
  wire       [15:0]   _zz_22995;
  wire       [31:0]   _zz_22996;
  wire       [31:0]   _zz_22997;
  wire       [31:0]   _zz_22998;
  wire       [31:0]   _zz_22999;
  wire       [31:0]   _zz_23000;
  wire       [23:0]   _zz_23001;
  wire       [31:0]   _zz_23002;
  wire       [15:0]   _zz_23003;
  wire       [31:0]   _zz_23004;
  wire       [31:0]   _zz_23005;
  wire       [31:0]   _zz_23006;
  wire       [31:0]   _zz_23007;
  wire       [31:0]   _zz_23008;
  wire       [23:0]   _zz_23009;
  wire       [31:0]   _zz_23010;
  wire       [15:0]   _zz_23011;
  wire       [15:0]   _zz_23012;
  wire       [31:0]   _zz_23013;
  wire       [31:0]   _zz_23014;
  wire       [15:0]   _zz_23015;
  wire       [31:0]   _zz_23016;
  wire       [31:0]   _zz_23017;
  wire       [31:0]   _zz_23018;
  wire       [15:0]   _zz_23019;
  wire       [31:0]   _zz_23020;
  wire       [31:0]   _zz_23021;
  wire       [31:0]   _zz_23022;
  wire       [31:0]   _zz_23023;
  wire       [31:0]   _zz_23024;
  wire       [31:0]   _zz_23025;
  wire       [23:0]   _zz_23026;
  wire       [31:0]   _zz_23027;
  wire       [15:0]   _zz_23028;
  wire       [31:0]   _zz_23029;
  wire       [31:0]   _zz_23030;
  wire       [31:0]   _zz_23031;
  wire       [31:0]   _zz_23032;
  wire       [31:0]   _zz_23033;
  wire       [23:0]   _zz_23034;
  wire       [31:0]   _zz_23035;
  wire       [15:0]   _zz_23036;
  wire       [31:0]   _zz_23037;
  wire       [31:0]   _zz_23038;
  wire       [31:0]   _zz_23039;
  wire       [31:0]   _zz_23040;
  wire       [31:0]   _zz_23041;
  wire       [23:0]   _zz_23042;
  wire       [31:0]   _zz_23043;
  wire       [15:0]   _zz_23044;
  wire       [31:0]   _zz_23045;
  wire       [31:0]   _zz_23046;
  wire       [31:0]   _zz_23047;
  wire       [31:0]   _zz_23048;
  wire       [31:0]   _zz_23049;
  wire       [23:0]   _zz_23050;
  wire       [31:0]   _zz_23051;
  wire       [15:0]   _zz_23052;
  wire       [15:0]   _zz_23053;
  wire       [31:0]   _zz_23054;
  wire       [31:0]   _zz_23055;
  wire       [15:0]   _zz_23056;
  wire       [31:0]   _zz_23057;
  wire       [31:0]   _zz_23058;
  wire       [31:0]   _zz_23059;
  wire       [15:0]   _zz_23060;
  wire       [31:0]   _zz_23061;
  wire       [31:0]   _zz_23062;
  wire       [31:0]   _zz_23063;
  wire       [31:0]   _zz_23064;
  wire       [31:0]   _zz_23065;
  wire       [31:0]   _zz_23066;
  wire       [23:0]   _zz_23067;
  wire       [31:0]   _zz_23068;
  wire       [15:0]   _zz_23069;
  wire       [31:0]   _zz_23070;
  wire       [31:0]   _zz_23071;
  wire       [31:0]   _zz_23072;
  wire       [31:0]   _zz_23073;
  wire       [31:0]   _zz_23074;
  wire       [23:0]   _zz_23075;
  wire       [31:0]   _zz_23076;
  wire       [15:0]   _zz_23077;
  wire       [31:0]   _zz_23078;
  wire       [31:0]   _zz_23079;
  wire       [31:0]   _zz_23080;
  wire       [31:0]   _zz_23081;
  wire       [31:0]   _zz_23082;
  wire       [23:0]   _zz_23083;
  wire       [31:0]   _zz_23084;
  wire       [15:0]   _zz_23085;
  wire       [31:0]   _zz_23086;
  wire       [31:0]   _zz_23087;
  wire       [31:0]   _zz_23088;
  wire       [31:0]   _zz_23089;
  wire       [31:0]   _zz_23090;
  wire       [23:0]   _zz_23091;
  wire       [31:0]   _zz_23092;
  wire       [15:0]   _zz_23093;
  wire       [15:0]   _zz_23094;
  wire       [31:0]   _zz_23095;
  wire       [31:0]   _zz_23096;
  wire       [15:0]   _zz_23097;
  wire       [31:0]   _zz_23098;
  wire       [31:0]   _zz_23099;
  wire       [31:0]   _zz_23100;
  wire       [15:0]   _zz_23101;
  wire       [31:0]   _zz_23102;
  wire       [31:0]   _zz_23103;
  wire       [31:0]   _zz_23104;
  wire       [31:0]   _zz_23105;
  wire       [31:0]   _zz_23106;
  wire       [31:0]   _zz_23107;
  wire       [23:0]   _zz_23108;
  wire       [31:0]   _zz_23109;
  wire       [15:0]   _zz_23110;
  wire       [31:0]   _zz_23111;
  wire       [31:0]   _zz_23112;
  wire       [31:0]   _zz_23113;
  wire       [31:0]   _zz_23114;
  wire       [31:0]   _zz_23115;
  wire       [23:0]   _zz_23116;
  wire       [31:0]   _zz_23117;
  wire       [15:0]   _zz_23118;
  wire       [31:0]   _zz_23119;
  wire       [31:0]   _zz_23120;
  wire       [31:0]   _zz_23121;
  wire       [31:0]   _zz_23122;
  wire       [31:0]   _zz_23123;
  wire       [23:0]   _zz_23124;
  wire       [31:0]   _zz_23125;
  wire       [15:0]   _zz_23126;
  wire       [31:0]   _zz_23127;
  wire       [31:0]   _zz_23128;
  wire       [31:0]   _zz_23129;
  wire       [31:0]   _zz_23130;
  wire       [31:0]   _zz_23131;
  wire       [23:0]   _zz_23132;
  wire       [31:0]   _zz_23133;
  wire       [15:0]   _zz_23134;
  wire       [15:0]   _zz_23135;
  wire       [31:0]   _zz_23136;
  wire       [31:0]   _zz_23137;
  wire       [15:0]   _zz_23138;
  wire       [31:0]   _zz_23139;
  wire       [31:0]   _zz_23140;
  wire       [31:0]   _zz_23141;
  wire       [15:0]   _zz_23142;
  wire       [31:0]   _zz_23143;
  wire       [31:0]   _zz_23144;
  wire       [31:0]   _zz_23145;
  wire       [31:0]   _zz_23146;
  wire       [31:0]   _zz_23147;
  wire       [31:0]   _zz_23148;
  wire       [23:0]   _zz_23149;
  wire       [31:0]   _zz_23150;
  wire       [15:0]   _zz_23151;
  wire       [31:0]   _zz_23152;
  wire       [31:0]   _zz_23153;
  wire       [31:0]   _zz_23154;
  wire       [31:0]   _zz_23155;
  wire       [31:0]   _zz_23156;
  wire       [23:0]   _zz_23157;
  wire       [31:0]   _zz_23158;
  wire       [15:0]   _zz_23159;
  wire       [31:0]   _zz_23160;
  wire       [31:0]   _zz_23161;
  wire       [31:0]   _zz_23162;
  wire       [31:0]   _zz_23163;
  wire       [31:0]   _zz_23164;
  wire       [23:0]   _zz_23165;
  wire       [31:0]   _zz_23166;
  wire       [15:0]   _zz_23167;
  wire       [31:0]   _zz_23168;
  wire       [31:0]   _zz_23169;
  wire       [31:0]   _zz_23170;
  wire       [31:0]   _zz_23171;
  wire       [31:0]   _zz_23172;
  wire       [23:0]   _zz_23173;
  wire       [31:0]   _zz_23174;
  wire       [15:0]   _zz_23175;
  wire       [15:0]   _zz_23176;
  wire       [31:0]   _zz_23177;
  wire       [31:0]   _zz_23178;
  wire       [15:0]   _zz_23179;
  wire       [31:0]   _zz_23180;
  wire       [31:0]   _zz_23181;
  wire       [31:0]   _zz_23182;
  wire       [15:0]   _zz_23183;
  wire       [31:0]   _zz_23184;
  wire       [31:0]   _zz_23185;
  wire       [31:0]   _zz_23186;
  wire       [31:0]   _zz_23187;
  wire       [31:0]   _zz_23188;
  wire       [31:0]   _zz_23189;
  wire       [23:0]   _zz_23190;
  wire       [31:0]   _zz_23191;
  wire       [15:0]   _zz_23192;
  wire       [31:0]   _zz_23193;
  wire       [31:0]   _zz_23194;
  wire       [31:0]   _zz_23195;
  wire       [31:0]   _zz_23196;
  wire       [31:0]   _zz_23197;
  wire       [23:0]   _zz_23198;
  wire       [31:0]   _zz_23199;
  wire       [15:0]   _zz_23200;
  wire       [31:0]   _zz_23201;
  wire       [31:0]   _zz_23202;
  wire       [31:0]   _zz_23203;
  wire       [31:0]   _zz_23204;
  wire       [31:0]   _zz_23205;
  wire       [23:0]   _zz_23206;
  wire       [31:0]   _zz_23207;
  wire       [15:0]   _zz_23208;
  wire       [31:0]   _zz_23209;
  wire       [31:0]   _zz_23210;
  wire       [31:0]   _zz_23211;
  wire       [31:0]   _zz_23212;
  wire       [31:0]   _zz_23213;
  wire       [23:0]   _zz_23214;
  wire       [31:0]   _zz_23215;
  wire       [15:0]   _zz_23216;
  wire       [15:0]   _zz_23217;
  wire       [31:0]   _zz_23218;
  wire       [31:0]   _zz_23219;
  wire       [15:0]   _zz_23220;
  wire       [31:0]   _zz_23221;
  wire       [31:0]   _zz_23222;
  wire       [31:0]   _zz_23223;
  wire       [15:0]   _zz_23224;
  wire       [31:0]   _zz_23225;
  wire       [31:0]   _zz_23226;
  wire       [31:0]   _zz_23227;
  wire       [31:0]   _zz_23228;
  wire       [31:0]   _zz_23229;
  wire       [31:0]   _zz_23230;
  wire       [23:0]   _zz_23231;
  wire       [31:0]   _zz_23232;
  wire       [15:0]   _zz_23233;
  wire       [31:0]   _zz_23234;
  wire       [31:0]   _zz_23235;
  wire       [31:0]   _zz_23236;
  wire       [31:0]   _zz_23237;
  wire       [31:0]   _zz_23238;
  wire       [23:0]   _zz_23239;
  wire       [31:0]   _zz_23240;
  wire       [15:0]   _zz_23241;
  wire       [31:0]   _zz_23242;
  wire       [31:0]   _zz_23243;
  wire       [31:0]   _zz_23244;
  wire       [31:0]   _zz_23245;
  wire       [31:0]   _zz_23246;
  wire       [23:0]   _zz_23247;
  wire       [31:0]   _zz_23248;
  wire       [15:0]   _zz_23249;
  wire       [31:0]   _zz_23250;
  wire       [31:0]   _zz_23251;
  wire       [31:0]   _zz_23252;
  wire       [31:0]   _zz_23253;
  wire       [31:0]   _zz_23254;
  wire       [23:0]   _zz_23255;
  wire       [31:0]   _zz_23256;
  wire       [15:0]   _zz_23257;
  wire       [15:0]   _zz_23258;
  wire       [31:0]   _zz_23259;
  wire       [31:0]   _zz_23260;
  wire       [15:0]   _zz_23261;
  wire       [31:0]   _zz_23262;
  wire       [31:0]   _zz_23263;
  wire       [31:0]   _zz_23264;
  wire       [15:0]   _zz_23265;
  wire       [31:0]   _zz_23266;
  wire       [31:0]   _zz_23267;
  wire       [31:0]   _zz_23268;
  wire       [31:0]   _zz_23269;
  wire       [31:0]   _zz_23270;
  wire       [31:0]   _zz_23271;
  wire       [23:0]   _zz_23272;
  wire       [31:0]   _zz_23273;
  wire       [15:0]   _zz_23274;
  wire       [31:0]   _zz_23275;
  wire       [31:0]   _zz_23276;
  wire       [31:0]   _zz_23277;
  wire       [31:0]   _zz_23278;
  wire       [31:0]   _zz_23279;
  wire       [23:0]   _zz_23280;
  wire       [31:0]   _zz_23281;
  wire       [15:0]   _zz_23282;
  wire       [31:0]   _zz_23283;
  wire       [31:0]   _zz_23284;
  wire       [31:0]   _zz_23285;
  wire       [31:0]   _zz_23286;
  wire       [31:0]   _zz_23287;
  wire       [23:0]   _zz_23288;
  wire       [31:0]   _zz_23289;
  wire       [15:0]   _zz_23290;
  wire       [31:0]   _zz_23291;
  wire       [31:0]   _zz_23292;
  wire       [31:0]   _zz_23293;
  wire       [31:0]   _zz_23294;
  wire       [31:0]   _zz_23295;
  wire       [23:0]   _zz_23296;
  wire       [31:0]   _zz_23297;
  wire       [15:0]   _zz_23298;
  reg        [15:0]   data_in_0_real;
  reg        [15:0]   data_in_0_imag;
  reg        [15:0]   data_in_1_real;
  reg        [15:0]   data_in_1_imag;
  reg        [15:0]   data_in_2_real;
  reg        [15:0]   data_in_2_imag;
  reg        [15:0]   data_in_3_real;
  reg        [15:0]   data_in_3_imag;
  reg        [15:0]   data_in_4_real;
  reg        [15:0]   data_in_4_imag;
  reg        [15:0]   data_in_5_real;
  reg        [15:0]   data_in_5_imag;
  reg        [15:0]   data_in_6_real;
  reg        [15:0]   data_in_6_imag;
  reg        [15:0]   data_in_7_real;
  reg        [15:0]   data_in_7_imag;
  reg        [15:0]   data_in_8_real;
  reg        [15:0]   data_in_8_imag;
  reg        [15:0]   data_in_9_real;
  reg        [15:0]   data_in_9_imag;
  reg        [15:0]   data_in_10_real;
  reg        [15:0]   data_in_10_imag;
  reg        [15:0]   data_in_11_real;
  reg        [15:0]   data_in_11_imag;
  reg        [15:0]   data_in_12_real;
  reg        [15:0]   data_in_12_imag;
  reg        [15:0]   data_in_13_real;
  reg        [15:0]   data_in_13_imag;
  reg        [15:0]   data_in_14_real;
  reg        [15:0]   data_in_14_imag;
  reg        [15:0]   data_in_15_real;
  reg        [15:0]   data_in_15_imag;
  reg        [15:0]   data_in_16_real;
  reg        [15:0]   data_in_16_imag;
  reg        [15:0]   data_in_17_real;
  reg        [15:0]   data_in_17_imag;
  reg        [15:0]   data_in_18_real;
  reg        [15:0]   data_in_18_imag;
  reg        [15:0]   data_in_19_real;
  reg        [15:0]   data_in_19_imag;
  reg        [15:0]   data_in_20_real;
  reg        [15:0]   data_in_20_imag;
  reg        [15:0]   data_in_21_real;
  reg        [15:0]   data_in_21_imag;
  reg        [15:0]   data_in_22_real;
  reg        [15:0]   data_in_22_imag;
  reg        [15:0]   data_in_23_real;
  reg        [15:0]   data_in_23_imag;
  reg        [15:0]   data_in_24_real;
  reg        [15:0]   data_in_24_imag;
  reg        [15:0]   data_in_25_real;
  reg        [15:0]   data_in_25_imag;
  reg        [15:0]   data_in_26_real;
  reg        [15:0]   data_in_26_imag;
  reg        [15:0]   data_in_27_real;
  reg        [15:0]   data_in_27_imag;
  reg        [15:0]   data_in_28_real;
  reg        [15:0]   data_in_28_imag;
  reg        [15:0]   data_in_29_real;
  reg        [15:0]   data_in_29_imag;
  reg        [15:0]   data_in_30_real;
  reg        [15:0]   data_in_30_imag;
  reg        [15:0]   data_in_31_real;
  reg        [15:0]   data_in_31_imag;
  reg        [15:0]   data_in_32_real;
  reg        [15:0]   data_in_32_imag;
  reg        [15:0]   data_in_33_real;
  reg        [15:0]   data_in_33_imag;
  reg        [15:0]   data_in_34_real;
  reg        [15:0]   data_in_34_imag;
  reg        [15:0]   data_in_35_real;
  reg        [15:0]   data_in_35_imag;
  reg        [15:0]   data_in_36_real;
  reg        [15:0]   data_in_36_imag;
  reg        [15:0]   data_in_37_real;
  reg        [15:0]   data_in_37_imag;
  reg        [15:0]   data_in_38_real;
  reg        [15:0]   data_in_38_imag;
  reg        [15:0]   data_in_39_real;
  reg        [15:0]   data_in_39_imag;
  reg        [15:0]   data_in_40_real;
  reg        [15:0]   data_in_40_imag;
  reg        [15:0]   data_in_41_real;
  reg        [15:0]   data_in_41_imag;
  reg        [15:0]   data_in_42_real;
  reg        [15:0]   data_in_42_imag;
  reg        [15:0]   data_in_43_real;
  reg        [15:0]   data_in_43_imag;
  reg        [15:0]   data_in_44_real;
  reg        [15:0]   data_in_44_imag;
  reg        [15:0]   data_in_45_real;
  reg        [15:0]   data_in_45_imag;
  reg        [15:0]   data_in_46_real;
  reg        [15:0]   data_in_46_imag;
  reg        [15:0]   data_in_47_real;
  reg        [15:0]   data_in_47_imag;
  reg        [15:0]   data_in_48_real;
  reg        [15:0]   data_in_48_imag;
  reg        [15:0]   data_in_49_real;
  reg        [15:0]   data_in_49_imag;
  reg        [15:0]   data_in_50_real;
  reg        [15:0]   data_in_50_imag;
  reg        [15:0]   data_in_51_real;
  reg        [15:0]   data_in_51_imag;
  reg        [15:0]   data_in_52_real;
  reg        [15:0]   data_in_52_imag;
  reg        [15:0]   data_in_53_real;
  reg        [15:0]   data_in_53_imag;
  reg        [15:0]   data_in_54_real;
  reg        [15:0]   data_in_54_imag;
  reg        [15:0]   data_in_55_real;
  reg        [15:0]   data_in_55_imag;
  reg        [15:0]   data_in_56_real;
  reg        [15:0]   data_in_56_imag;
  reg        [15:0]   data_in_57_real;
  reg        [15:0]   data_in_57_imag;
  reg        [15:0]   data_in_58_real;
  reg        [15:0]   data_in_58_imag;
  reg        [15:0]   data_in_59_real;
  reg        [15:0]   data_in_59_imag;
  reg        [15:0]   data_in_60_real;
  reg        [15:0]   data_in_60_imag;
  reg        [15:0]   data_in_61_real;
  reg        [15:0]   data_in_61_imag;
  reg        [15:0]   data_in_62_real;
  reg        [15:0]   data_in_62_imag;
  reg        [15:0]   data_in_63_real;
  reg        [15:0]   data_in_63_imag;
  reg        [15:0]   data_in_64_real;
  reg        [15:0]   data_in_64_imag;
  reg        [15:0]   data_in_65_real;
  reg        [15:0]   data_in_65_imag;
  reg        [15:0]   data_in_66_real;
  reg        [15:0]   data_in_66_imag;
  reg        [15:0]   data_in_67_real;
  reg        [15:0]   data_in_67_imag;
  reg        [15:0]   data_in_68_real;
  reg        [15:0]   data_in_68_imag;
  reg        [15:0]   data_in_69_real;
  reg        [15:0]   data_in_69_imag;
  reg        [15:0]   data_in_70_real;
  reg        [15:0]   data_in_70_imag;
  reg        [15:0]   data_in_71_real;
  reg        [15:0]   data_in_71_imag;
  reg        [15:0]   data_in_72_real;
  reg        [15:0]   data_in_72_imag;
  reg        [15:0]   data_in_73_real;
  reg        [15:0]   data_in_73_imag;
  reg        [15:0]   data_in_74_real;
  reg        [15:0]   data_in_74_imag;
  reg        [15:0]   data_in_75_real;
  reg        [15:0]   data_in_75_imag;
  reg        [15:0]   data_in_76_real;
  reg        [15:0]   data_in_76_imag;
  reg        [15:0]   data_in_77_real;
  reg        [15:0]   data_in_77_imag;
  reg        [15:0]   data_in_78_real;
  reg        [15:0]   data_in_78_imag;
  reg        [15:0]   data_in_79_real;
  reg        [15:0]   data_in_79_imag;
  reg        [15:0]   data_in_80_real;
  reg        [15:0]   data_in_80_imag;
  reg        [15:0]   data_in_81_real;
  reg        [15:0]   data_in_81_imag;
  reg        [15:0]   data_in_82_real;
  reg        [15:0]   data_in_82_imag;
  reg        [15:0]   data_in_83_real;
  reg        [15:0]   data_in_83_imag;
  reg        [15:0]   data_in_84_real;
  reg        [15:0]   data_in_84_imag;
  reg        [15:0]   data_in_85_real;
  reg        [15:0]   data_in_85_imag;
  reg        [15:0]   data_in_86_real;
  reg        [15:0]   data_in_86_imag;
  reg        [15:0]   data_in_87_real;
  reg        [15:0]   data_in_87_imag;
  reg        [15:0]   data_in_88_real;
  reg        [15:0]   data_in_88_imag;
  reg        [15:0]   data_in_89_real;
  reg        [15:0]   data_in_89_imag;
  reg        [15:0]   data_in_90_real;
  reg        [15:0]   data_in_90_imag;
  reg        [15:0]   data_in_91_real;
  reg        [15:0]   data_in_91_imag;
  reg        [15:0]   data_in_92_real;
  reg        [15:0]   data_in_92_imag;
  reg        [15:0]   data_in_93_real;
  reg        [15:0]   data_in_93_imag;
  reg        [15:0]   data_in_94_real;
  reg        [15:0]   data_in_94_imag;
  reg        [15:0]   data_in_95_real;
  reg        [15:0]   data_in_95_imag;
  reg        [15:0]   data_in_96_real;
  reg        [15:0]   data_in_96_imag;
  reg        [15:0]   data_in_97_real;
  reg        [15:0]   data_in_97_imag;
  reg        [15:0]   data_in_98_real;
  reg        [15:0]   data_in_98_imag;
  reg        [15:0]   data_in_99_real;
  reg        [15:0]   data_in_99_imag;
  reg        [15:0]   data_in_100_real;
  reg        [15:0]   data_in_100_imag;
  reg        [15:0]   data_in_101_real;
  reg        [15:0]   data_in_101_imag;
  reg        [15:0]   data_in_102_real;
  reg        [15:0]   data_in_102_imag;
  reg        [15:0]   data_in_103_real;
  reg        [15:0]   data_in_103_imag;
  reg        [15:0]   data_in_104_real;
  reg        [15:0]   data_in_104_imag;
  reg        [15:0]   data_in_105_real;
  reg        [15:0]   data_in_105_imag;
  reg        [15:0]   data_in_106_real;
  reg        [15:0]   data_in_106_imag;
  reg        [15:0]   data_in_107_real;
  reg        [15:0]   data_in_107_imag;
  reg        [15:0]   data_in_108_real;
  reg        [15:0]   data_in_108_imag;
  reg        [15:0]   data_in_109_real;
  reg        [15:0]   data_in_109_imag;
  reg        [15:0]   data_in_110_real;
  reg        [15:0]   data_in_110_imag;
  reg        [15:0]   data_in_111_real;
  reg        [15:0]   data_in_111_imag;
  reg        [15:0]   data_in_112_real;
  reg        [15:0]   data_in_112_imag;
  reg        [15:0]   data_in_113_real;
  reg        [15:0]   data_in_113_imag;
  reg        [15:0]   data_in_114_real;
  reg        [15:0]   data_in_114_imag;
  reg        [15:0]   data_in_115_real;
  reg        [15:0]   data_in_115_imag;
  reg        [15:0]   data_in_116_real;
  reg        [15:0]   data_in_116_imag;
  reg        [15:0]   data_in_117_real;
  reg        [15:0]   data_in_117_imag;
  reg        [15:0]   data_in_118_real;
  reg        [15:0]   data_in_118_imag;
  reg        [15:0]   data_in_119_real;
  reg        [15:0]   data_in_119_imag;
  reg        [15:0]   data_in_120_real;
  reg        [15:0]   data_in_120_imag;
  reg        [15:0]   data_in_121_real;
  reg        [15:0]   data_in_121_imag;
  reg        [15:0]   data_in_122_real;
  reg        [15:0]   data_in_122_imag;
  reg        [15:0]   data_in_123_real;
  reg        [15:0]   data_in_123_imag;
  reg        [15:0]   data_in_124_real;
  reg        [15:0]   data_in_124_imag;
  reg        [15:0]   data_in_125_real;
  reg        [15:0]   data_in_125_imag;
  reg        [15:0]   data_in_126_real;
  reg        [15:0]   data_in_126_imag;
  reg        [15:0]   data_in_127_real;
  reg        [15:0]   data_in_127_imag;
  wire       [15:0]   twiddle_factor_table_0_real;
  wire       [15:0]   twiddle_factor_table_0_imag;
  wire       [15:0]   twiddle_factor_table_1_real;
  wire       [15:0]   twiddle_factor_table_1_imag;
  wire       [15:0]   twiddle_factor_table_2_real;
  wire       [15:0]   twiddle_factor_table_2_imag;
  wire       [15:0]   twiddle_factor_table_3_real;
  wire       [15:0]   twiddle_factor_table_3_imag;
  wire       [15:0]   twiddle_factor_table_4_real;
  wire       [15:0]   twiddle_factor_table_4_imag;
  wire       [15:0]   twiddle_factor_table_5_real;
  wire       [15:0]   twiddle_factor_table_5_imag;
  wire       [15:0]   twiddle_factor_table_6_real;
  wire       [15:0]   twiddle_factor_table_6_imag;
  wire       [15:0]   twiddle_factor_table_7_real;
  wire       [15:0]   twiddle_factor_table_7_imag;
  wire       [15:0]   twiddle_factor_table_8_real;
  wire       [15:0]   twiddle_factor_table_8_imag;
  wire       [15:0]   twiddle_factor_table_9_real;
  wire       [15:0]   twiddle_factor_table_9_imag;
  wire       [15:0]   twiddle_factor_table_10_real;
  wire       [15:0]   twiddle_factor_table_10_imag;
  wire       [15:0]   twiddle_factor_table_11_real;
  wire       [15:0]   twiddle_factor_table_11_imag;
  wire       [15:0]   twiddle_factor_table_12_real;
  wire       [15:0]   twiddle_factor_table_12_imag;
  wire       [15:0]   twiddle_factor_table_13_real;
  wire       [15:0]   twiddle_factor_table_13_imag;
  wire       [15:0]   twiddle_factor_table_14_real;
  wire       [15:0]   twiddle_factor_table_14_imag;
  wire       [15:0]   twiddle_factor_table_15_real;
  wire       [15:0]   twiddle_factor_table_15_imag;
  wire       [15:0]   twiddle_factor_table_16_real;
  wire       [15:0]   twiddle_factor_table_16_imag;
  wire       [15:0]   twiddle_factor_table_17_real;
  wire       [15:0]   twiddle_factor_table_17_imag;
  wire       [15:0]   twiddle_factor_table_18_real;
  wire       [15:0]   twiddle_factor_table_18_imag;
  wire       [15:0]   twiddle_factor_table_19_real;
  wire       [15:0]   twiddle_factor_table_19_imag;
  wire       [15:0]   twiddle_factor_table_20_real;
  wire       [15:0]   twiddle_factor_table_20_imag;
  wire       [15:0]   twiddle_factor_table_21_real;
  wire       [15:0]   twiddle_factor_table_21_imag;
  wire       [15:0]   twiddle_factor_table_22_real;
  wire       [15:0]   twiddle_factor_table_22_imag;
  wire       [15:0]   twiddle_factor_table_23_real;
  wire       [15:0]   twiddle_factor_table_23_imag;
  wire       [15:0]   twiddle_factor_table_24_real;
  wire       [15:0]   twiddle_factor_table_24_imag;
  wire       [15:0]   twiddle_factor_table_25_real;
  wire       [15:0]   twiddle_factor_table_25_imag;
  wire       [15:0]   twiddle_factor_table_26_real;
  wire       [15:0]   twiddle_factor_table_26_imag;
  wire       [15:0]   twiddle_factor_table_27_real;
  wire       [15:0]   twiddle_factor_table_27_imag;
  wire       [15:0]   twiddle_factor_table_28_real;
  wire       [15:0]   twiddle_factor_table_28_imag;
  wire       [15:0]   twiddle_factor_table_29_real;
  wire       [15:0]   twiddle_factor_table_29_imag;
  wire       [15:0]   twiddle_factor_table_30_real;
  wire       [15:0]   twiddle_factor_table_30_imag;
  wire       [15:0]   twiddle_factor_table_31_real;
  wire       [15:0]   twiddle_factor_table_31_imag;
  wire       [15:0]   twiddle_factor_table_32_real;
  wire       [15:0]   twiddle_factor_table_32_imag;
  wire       [15:0]   twiddle_factor_table_33_real;
  wire       [15:0]   twiddle_factor_table_33_imag;
  wire       [15:0]   twiddle_factor_table_34_real;
  wire       [15:0]   twiddle_factor_table_34_imag;
  wire       [15:0]   twiddle_factor_table_35_real;
  wire       [15:0]   twiddle_factor_table_35_imag;
  wire       [15:0]   twiddle_factor_table_36_real;
  wire       [15:0]   twiddle_factor_table_36_imag;
  wire       [15:0]   twiddle_factor_table_37_real;
  wire       [15:0]   twiddle_factor_table_37_imag;
  wire       [15:0]   twiddle_factor_table_38_real;
  wire       [15:0]   twiddle_factor_table_38_imag;
  wire       [15:0]   twiddle_factor_table_39_real;
  wire       [15:0]   twiddle_factor_table_39_imag;
  wire       [15:0]   twiddle_factor_table_40_real;
  wire       [15:0]   twiddle_factor_table_40_imag;
  wire       [15:0]   twiddle_factor_table_41_real;
  wire       [15:0]   twiddle_factor_table_41_imag;
  wire       [15:0]   twiddle_factor_table_42_real;
  wire       [15:0]   twiddle_factor_table_42_imag;
  wire       [15:0]   twiddle_factor_table_43_real;
  wire       [15:0]   twiddle_factor_table_43_imag;
  wire       [15:0]   twiddle_factor_table_44_real;
  wire       [15:0]   twiddle_factor_table_44_imag;
  wire       [15:0]   twiddle_factor_table_45_real;
  wire       [15:0]   twiddle_factor_table_45_imag;
  wire       [15:0]   twiddle_factor_table_46_real;
  wire       [15:0]   twiddle_factor_table_46_imag;
  wire       [15:0]   twiddle_factor_table_47_real;
  wire       [15:0]   twiddle_factor_table_47_imag;
  wire       [15:0]   twiddle_factor_table_48_real;
  wire       [15:0]   twiddle_factor_table_48_imag;
  wire       [15:0]   twiddle_factor_table_49_real;
  wire       [15:0]   twiddle_factor_table_49_imag;
  wire       [15:0]   twiddle_factor_table_50_real;
  wire       [15:0]   twiddle_factor_table_50_imag;
  wire       [15:0]   twiddle_factor_table_51_real;
  wire       [15:0]   twiddle_factor_table_51_imag;
  wire       [15:0]   twiddle_factor_table_52_real;
  wire       [15:0]   twiddle_factor_table_52_imag;
  wire       [15:0]   twiddle_factor_table_53_real;
  wire       [15:0]   twiddle_factor_table_53_imag;
  wire       [15:0]   twiddle_factor_table_54_real;
  wire       [15:0]   twiddle_factor_table_54_imag;
  wire       [15:0]   twiddle_factor_table_55_real;
  wire       [15:0]   twiddle_factor_table_55_imag;
  wire       [15:0]   twiddle_factor_table_56_real;
  wire       [15:0]   twiddle_factor_table_56_imag;
  wire       [15:0]   twiddle_factor_table_57_real;
  wire       [15:0]   twiddle_factor_table_57_imag;
  wire       [15:0]   twiddle_factor_table_58_real;
  wire       [15:0]   twiddle_factor_table_58_imag;
  wire       [15:0]   twiddle_factor_table_59_real;
  wire       [15:0]   twiddle_factor_table_59_imag;
  wire       [15:0]   twiddle_factor_table_60_real;
  wire       [15:0]   twiddle_factor_table_60_imag;
  wire       [15:0]   twiddle_factor_table_61_real;
  wire       [15:0]   twiddle_factor_table_61_imag;
  wire       [15:0]   twiddle_factor_table_62_real;
  wire       [15:0]   twiddle_factor_table_62_imag;
  wire       [15:0]   twiddle_factor_table_63_real;
  wire       [15:0]   twiddle_factor_table_63_imag;
  wire       [15:0]   twiddle_factor_table_64_real;
  wire       [15:0]   twiddle_factor_table_64_imag;
  wire       [15:0]   twiddle_factor_table_65_real;
  wire       [15:0]   twiddle_factor_table_65_imag;
  wire       [15:0]   twiddle_factor_table_66_real;
  wire       [15:0]   twiddle_factor_table_66_imag;
  wire       [15:0]   twiddle_factor_table_67_real;
  wire       [15:0]   twiddle_factor_table_67_imag;
  wire       [15:0]   twiddle_factor_table_68_real;
  wire       [15:0]   twiddle_factor_table_68_imag;
  wire       [15:0]   twiddle_factor_table_69_real;
  wire       [15:0]   twiddle_factor_table_69_imag;
  wire       [15:0]   twiddle_factor_table_70_real;
  wire       [15:0]   twiddle_factor_table_70_imag;
  wire       [15:0]   twiddle_factor_table_71_real;
  wire       [15:0]   twiddle_factor_table_71_imag;
  wire       [15:0]   twiddle_factor_table_72_real;
  wire       [15:0]   twiddle_factor_table_72_imag;
  wire       [15:0]   twiddle_factor_table_73_real;
  wire       [15:0]   twiddle_factor_table_73_imag;
  wire       [15:0]   twiddle_factor_table_74_real;
  wire       [15:0]   twiddle_factor_table_74_imag;
  wire       [15:0]   twiddle_factor_table_75_real;
  wire       [15:0]   twiddle_factor_table_75_imag;
  wire       [15:0]   twiddle_factor_table_76_real;
  wire       [15:0]   twiddle_factor_table_76_imag;
  wire       [15:0]   twiddle_factor_table_77_real;
  wire       [15:0]   twiddle_factor_table_77_imag;
  wire       [15:0]   twiddle_factor_table_78_real;
  wire       [15:0]   twiddle_factor_table_78_imag;
  wire       [15:0]   twiddle_factor_table_79_real;
  wire       [15:0]   twiddle_factor_table_79_imag;
  wire       [15:0]   twiddle_factor_table_80_real;
  wire       [15:0]   twiddle_factor_table_80_imag;
  wire       [15:0]   twiddle_factor_table_81_real;
  wire       [15:0]   twiddle_factor_table_81_imag;
  wire       [15:0]   twiddle_factor_table_82_real;
  wire       [15:0]   twiddle_factor_table_82_imag;
  wire       [15:0]   twiddle_factor_table_83_real;
  wire       [15:0]   twiddle_factor_table_83_imag;
  wire       [15:0]   twiddle_factor_table_84_real;
  wire       [15:0]   twiddle_factor_table_84_imag;
  wire       [15:0]   twiddle_factor_table_85_real;
  wire       [15:0]   twiddle_factor_table_85_imag;
  wire       [15:0]   twiddle_factor_table_86_real;
  wire       [15:0]   twiddle_factor_table_86_imag;
  wire       [15:0]   twiddle_factor_table_87_real;
  wire       [15:0]   twiddle_factor_table_87_imag;
  wire       [15:0]   twiddle_factor_table_88_real;
  wire       [15:0]   twiddle_factor_table_88_imag;
  wire       [15:0]   twiddle_factor_table_89_real;
  wire       [15:0]   twiddle_factor_table_89_imag;
  wire       [15:0]   twiddle_factor_table_90_real;
  wire       [15:0]   twiddle_factor_table_90_imag;
  wire       [15:0]   twiddle_factor_table_91_real;
  wire       [15:0]   twiddle_factor_table_91_imag;
  wire       [15:0]   twiddle_factor_table_92_real;
  wire       [15:0]   twiddle_factor_table_92_imag;
  wire       [15:0]   twiddle_factor_table_93_real;
  wire       [15:0]   twiddle_factor_table_93_imag;
  wire       [15:0]   twiddle_factor_table_94_real;
  wire       [15:0]   twiddle_factor_table_94_imag;
  wire       [15:0]   twiddle_factor_table_95_real;
  wire       [15:0]   twiddle_factor_table_95_imag;
  wire       [15:0]   twiddle_factor_table_96_real;
  wire       [15:0]   twiddle_factor_table_96_imag;
  wire       [15:0]   twiddle_factor_table_97_real;
  wire       [15:0]   twiddle_factor_table_97_imag;
  wire       [15:0]   twiddle_factor_table_98_real;
  wire       [15:0]   twiddle_factor_table_98_imag;
  wire       [15:0]   twiddle_factor_table_99_real;
  wire       [15:0]   twiddle_factor_table_99_imag;
  wire       [15:0]   twiddle_factor_table_100_real;
  wire       [15:0]   twiddle_factor_table_100_imag;
  wire       [15:0]   twiddle_factor_table_101_real;
  wire       [15:0]   twiddle_factor_table_101_imag;
  wire       [15:0]   twiddle_factor_table_102_real;
  wire       [15:0]   twiddle_factor_table_102_imag;
  wire       [15:0]   twiddle_factor_table_103_real;
  wire       [15:0]   twiddle_factor_table_103_imag;
  wire       [15:0]   twiddle_factor_table_104_real;
  wire       [15:0]   twiddle_factor_table_104_imag;
  wire       [15:0]   twiddle_factor_table_105_real;
  wire       [15:0]   twiddle_factor_table_105_imag;
  wire       [15:0]   twiddle_factor_table_106_real;
  wire       [15:0]   twiddle_factor_table_106_imag;
  wire       [15:0]   twiddle_factor_table_107_real;
  wire       [15:0]   twiddle_factor_table_107_imag;
  wire       [15:0]   twiddle_factor_table_108_real;
  wire       [15:0]   twiddle_factor_table_108_imag;
  wire       [15:0]   twiddle_factor_table_109_real;
  wire       [15:0]   twiddle_factor_table_109_imag;
  wire       [15:0]   twiddle_factor_table_110_real;
  wire       [15:0]   twiddle_factor_table_110_imag;
  wire       [15:0]   twiddle_factor_table_111_real;
  wire       [15:0]   twiddle_factor_table_111_imag;
  wire       [15:0]   twiddle_factor_table_112_real;
  wire       [15:0]   twiddle_factor_table_112_imag;
  wire       [15:0]   twiddle_factor_table_113_real;
  wire       [15:0]   twiddle_factor_table_113_imag;
  wire       [15:0]   twiddle_factor_table_114_real;
  wire       [15:0]   twiddle_factor_table_114_imag;
  wire       [15:0]   twiddle_factor_table_115_real;
  wire       [15:0]   twiddle_factor_table_115_imag;
  wire       [15:0]   twiddle_factor_table_116_real;
  wire       [15:0]   twiddle_factor_table_116_imag;
  wire       [15:0]   twiddle_factor_table_117_real;
  wire       [15:0]   twiddle_factor_table_117_imag;
  wire       [15:0]   twiddle_factor_table_118_real;
  wire       [15:0]   twiddle_factor_table_118_imag;
  wire       [15:0]   twiddle_factor_table_119_real;
  wire       [15:0]   twiddle_factor_table_119_imag;
  wire       [15:0]   twiddle_factor_table_120_real;
  wire       [15:0]   twiddle_factor_table_120_imag;
  wire       [15:0]   twiddle_factor_table_121_real;
  wire       [15:0]   twiddle_factor_table_121_imag;
  wire       [15:0]   twiddle_factor_table_122_real;
  wire       [15:0]   twiddle_factor_table_122_imag;
  wire       [15:0]   twiddle_factor_table_123_real;
  wire       [15:0]   twiddle_factor_table_123_imag;
  wire       [15:0]   twiddle_factor_table_124_real;
  wire       [15:0]   twiddle_factor_table_124_imag;
  wire       [15:0]   twiddle_factor_table_125_real;
  wire       [15:0]   twiddle_factor_table_125_imag;
  wire       [15:0]   twiddle_factor_table_126_real;
  wire       [15:0]   twiddle_factor_table_126_imag;
  wire       [15:0]   data_reorder_0_real;
  wire       [15:0]   data_reorder_0_imag;
  wire       [15:0]   data_reorder_1_real;
  wire       [15:0]   data_reorder_1_imag;
  wire       [15:0]   data_reorder_2_real;
  wire       [15:0]   data_reorder_2_imag;
  wire       [15:0]   data_reorder_3_real;
  wire       [15:0]   data_reorder_3_imag;
  wire       [15:0]   data_reorder_4_real;
  wire       [15:0]   data_reorder_4_imag;
  wire       [15:0]   data_reorder_5_real;
  wire       [15:0]   data_reorder_5_imag;
  wire       [15:0]   data_reorder_6_real;
  wire       [15:0]   data_reorder_6_imag;
  wire       [15:0]   data_reorder_7_real;
  wire       [15:0]   data_reorder_7_imag;
  wire       [15:0]   data_reorder_8_real;
  wire       [15:0]   data_reorder_8_imag;
  wire       [15:0]   data_reorder_9_real;
  wire       [15:0]   data_reorder_9_imag;
  wire       [15:0]   data_reorder_10_real;
  wire       [15:0]   data_reorder_10_imag;
  wire       [15:0]   data_reorder_11_real;
  wire       [15:0]   data_reorder_11_imag;
  wire       [15:0]   data_reorder_12_real;
  wire       [15:0]   data_reorder_12_imag;
  wire       [15:0]   data_reorder_13_real;
  wire       [15:0]   data_reorder_13_imag;
  wire       [15:0]   data_reorder_14_real;
  wire       [15:0]   data_reorder_14_imag;
  wire       [15:0]   data_reorder_15_real;
  wire       [15:0]   data_reorder_15_imag;
  wire       [15:0]   data_reorder_16_real;
  wire       [15:0]   data_reorder_16_imag;
  wire       [15:0]   data_reorder_17_real;
  wire       [15:0]   data_reorder_17_imag;
  wire       [15:0]   data_reorder_18_real;
  wire       [15:0]   data_reorder_18_imag;
  wire       [15:0]   data_reorder_19_real;
  wire       [15:0]   data_reorder_19_imag;
  wire       [15:0]   data_reorder_20_real;
  wire       [15:0]   data_reorder_20_imag;
  wire       [15:0]   data_reorder_21_real;
  wire       [15:0]   data_reorder_21_imag;
  wire       [15:0]   data_reorder_22_real;
  wire       [15:0]   data_reorder_22_imag;
  wire       [15:0]   data_reorder_23_real;
  wire       [15:0]   data_reorder_23_imag;
  wire       [15:0]   data_reorder_24_real;
  wire       [15:0]   data_reorder_24_imag;
  wire       [15:0]   data_reorder_25_real;
  wire       [15:0]   data_reorder_25_imag;
  wire       [15:0]   data_reorder_26_real;
  wire       [15:0]   data_reorder_26_imag;
  wire       [15:0]   data_reorder_27_real;
  wire       [15:0]   data_reorder_27_imag;
  wire       [15:0]   data_reorder_28_real;
  wire       [15:0]   data_reorder_28_imag;
  wire       [15:0]   data_reorder_29_real;
  wire       [15:0]   data_reorder_29_imag;
  wire       [15:0]   data_reorder_30_real;
  wire       [15:0]   data_reorder_30_imag;
  wire       [15:0]   data_reorder_31_real;
  wire       [15:0]   data_reorder_31_imag;
  wire       [15:0]   data_reorder_32_real;
  wire       [15:0]   data_reorder_32_imag;
  wire       [15:0]   data_reorder_33_real;
  wire       [15:0]   data_reorder_33_imag;
  wire       [15:0]   data_reorder_34_real;
  wire       [15:0]   data_reorder_34_imag;
  wire       [15:0]   data_reorder_35_real;
  wire       [15:0]   data_reorder_35_imag;
  wire       [15:0]   data_reorder_36_real;
  wire       [15:0]   data_reorder_36_imag;
  wire       [15:0]   data_reorder_37_real;
  wire       [15:0]   data_reorder_37_imag;
  wire       [15:0]   data_reorder_38_real;
  wire       [15:0]   data_reorder_38_imag;
  wire       [15:0]   data_reorder_39_real;
  wire       [15:0]   data_reorder_39_imag;
  wire       [15:0]   data_reorder_40_real;
  wire       [15:0]   data_reorder_40_imag;
  wire       [15:0]   data_reorder_41_real;
  wire       [15:0]   data_reorder_41_imag;
  wire       [15:0]   data_reorder_42_real;
  wire       [15:0]   data_reorder_42_imag;
  wire       [15:0]   data_reorder_43_real;
  wire       [15:0]   data_reorder_43_imag;
  wire       [15:0]   data_reorder_44_real;
  wire       [15:0]   data_reorder_44_imag;
  wire       [15:0]   data_reorder_45_real;
  wire       [15:0]   data_reorder_45_imag;
  wire       [15:0]   data_reorder_46_real;
  wire       [15:0]   data_reorder_46_imag;
  wire       [15:0]   data_reorder_47_real;
  wire       [15:0]   data_reorder_47_imag;
  wire       [15:0]   data_reorder_48_real;
  wire       [15:0]   data_reorder_48_imag;
  wire       [15:0]   data_reorder_49_real;
  wire       [15:0]   data_reorder_49_imag;
  wire       [15:0]   data_reorder_50_real;
  wire       [15:0]   data_reorder_50_imag;
  wire       [15:0]   data_reorder_51_real;
  wire       [15:0]   data_reorder_51_imag;
  wire       [15:0]   data_reorder_52_real;
  wire       [15:0]   data_reorder_52_imag;
  wire       [15:0]   data_reorder_53_real;
  wire       [15:0]   data_reorder_53_imag;
  wire       [15:0]   data_reorder_54_real;
  wire       [15:0]   data_reorder_54_imag;
  wire       [15:0]   data_reorder_55_real;
  wire       [15:0]   data_reorder_55_imag;
  wire       [15:0]   data_reorder_56_real;
  wire       [15:0]   data_reorder_56_imag;
  wire       [15:0]   data_reorder_57_real;
  wire       [15:0]   data_reorder_57_imag;
  wire       [15:0]   data_reorder_58_real;
  wire       [15:0]   data_reorder_58_imag;
  wire       [15:0]   data_reorder_59_real;
  wire       [15:0]   data_reorder_59_imag;
  wire       [15:0]   data_reorder_60_real;
  wire       [15:0]   data_reorder_60_imag;
  wire       [15:0]   data_reorder_61_real;
  wire       [15:0]   data_reorder_61_imag;
  wire       [15:0]   data_reorder_62_real;
  wire       [15:0]   data_reorder_62_imag;
  wire       [15:0]   data_reorder_63_real;
  wire       [15:0]   data_reorder_63_imag;
  wire       [15:0]   data_reorder_64_real;
  wire       [15:0]   data_reorder_64_imag;
  wire       [15:0]   data_reorder_65_real;
  wire       [15:0]   data_reorder_65_imag;
  wire       [15:0]   data_reorder_66_real;
  wire       [15:0]   data_reorder_66_imag;
  wire       [15:0]   data_reorder_67_real;
  wire       [15:0]   data_reorder_67_imag;
  wire       [15:0]   data_reorder_68_real;
  wire       [15:0]   data_reorder_68_imag;
  wire       [15:0]   data_reorder_69_real;
  wire       [15:0]   data_reorder_69_imag;
  wire       [15:0]   data_reorder_70_real;
  wire       [15:0]   data_reorder_70_imag;
  wire       [15:0]   data_reorder_71_real;
  wire       [15:0]   data_reorder_71_imag;
  wire       [15:0]   data_reorder_72_real;
  wire       [15:0]   data_reorder_72_imag;
  wire       [15:0]   data_reorder_73_real;
  wire       [15:0]   data_reorder_73_imag;
  wire       [15:0]   data_reorder_74_real;
  wire       [15:0]   data_reorder_74_imag;
  wire       [15:0]   data_reorder_75_real;
  wire       [15:0]   data_reorder_75_imag;
  wire       [15:0]   data_reorder_76_real;
  wire       [15:0]   data_reorder_76_imag;
  wire       [15:0]   data_reorder_77_real;
  wire       [15:0]   data_reorder_77_imag;
  wire       [15:0]   data_reorder_78_real;
  wire       [15:0]   data_reorder_78_imag;
  wire       [15:0]   data_reorder_79_real;
  wire       [15:0]   data_reorder_79_imag;
  wire       [15:0]   data_reorder_80_real;
  wire       [15:0]   data_reorder_80_imag;
  wire       [15:0]   data_reorder_81_real;
  wire       [15:0]   data_reorder_81_imag;
  wire       [15:0]   data_reorder_82_real;
  wire       [15:0]   data_reorder_82_imag;
  wire       [15:0]   data_reorder_83_real;
  wire       [15:0]   data_reorder_83_imag;
  wire       [15:0]   data_reorder_84_real;
  wire       [15:0]   data_reorder_84_imag;
  wire       [15:0]   data_reorder_85_real;
  wire       [15:0]   data_reorder_85_imag;
  wire       [15:0]   data_reorder_86_real;
  wire       [15:0]   data_reorder_86_imag;
  wire       [15:0]   data_reorder_87_real;
  wire       [15:0]   data_reorder_87_imag;
  wire       [15:0]   data_reorder_88_real;
  wire       [15:0]   data_reorder_88_imag;
  wire       [15:0]   data_reorder_89_real;
  wire       [15:0]   data_reorder_89_imag;
  wire       [15:0]   data_reorder_90_real;
  wire       [15:0]   data_reorder_90_imag;
  wire       [15:0]   data_reorder_91_real;
  wire       [15:0]   data_reorder_91_imag;
  wire       [15:0]   data_reorder_92_real;
  wire       [15:0]   data_reorder_92_imag;
  wire       [15:0]   data_reorder_93_real;
  wire       [15:0]   data_reorder_93_imag;
  wire       [15:0]   data_reorder_94_real;
  wire       [15:0]   data_reorder_94_imag;
  wire       [15:0]   data_reorder_95_real;
  wire       [15:0]   data_reorder_95_imag;
  wire       [15:0]   data_reorder_96_real;
  wire       [15:0]   data_reorder_96_imag;
  wire       [15:0]   data_reorder_97_real;
  wire       [15:0]   data_reorder_97_imag;
  wire       [15:0]   data_reorder_98_real;
  wire       [15:0]   data_reorder_98_imag;
  wire       [15:0]   data_reorder_99_real;
  wire       [15:0]   data_reorder_99_imag;
  wire       [15:0]   data_reorder_100_real;
  wire       [15:0]   data_reorder_100_imag;
  wire       [15:0]   data_reorder_101_real;
  wire       [15:0]   data_reorder_101_imag;
  wire       [15:0]   data_reorder_102_real;
  wire       [15:0]   data_reorder_102_imag;
  wire       [15:0]   data_reorder_103_real;
  wire       [15:0]   data_reorder_103_imag;
  wire       [15:0]   data_reorder_104_real;
  wire       [15:0]   data_reorder_104_imag;
  wire       [15:0]   data_reorder_105_real;
  wire       [15:0]   data_reorder_105_imag;
  wire       [15:0]   data_reorder_106_real;
  wire       [15:0]   data_reorder_106_imag;
  wire       [15:0]   data_reorder_107_real;
  wire       [15:0]   data_reorder_107_imag;
  wire       [15:0]   data_reorder_108_real;
  wire       [15:0]   data_reorder_108_imag;
  wire       [15:0]   data_reorder_109_real;
  wire       [15:0]   data_reorder_109_imag;
  wire       [15:0]   data_reorder_110_real;
  wire       [15:0]   data_reorder_110_imag;
  wire       [15:0]   data_reorder_111_real;
  wire       [15:0]   data_reorder_111_imag;
  wire       [15:0]   data_reorder_112_real;
  wire       [15:0]   data_reorder_112_imag;
  wire       [15:0]   data_reorder_113_real;
  wire       [15:0]   data_reorder_113_imag;
  wire       [15:0]   data_reorder_114_real;
  wire       [15:0]   data_reorder_114_imag;
  wire       [15:0]   data_reorder_115_real;
  wire       [15:0]   data_reorder_115_imag;
  wire       [15:0]   data_reorder_116_real;
  wire       [15:0]   data_reorder_116_imag;
  wire       [15:0]   data_reorder_117_real;
  wire       [15:0]   data_reorder_117_imag;
  wire       [15:0]   data_reorder_118_real;
  wire       [15:0]   data_reorder_118_imag;
  wire       [15:0]   data_reorder_119_real;
  wire       [15:0]   data_reorder_119_imag;
  wire       [15:0]   data_reorder_120_real;
  wire       [15:0]   data_reorder_120_imag;
  wire       [15:0]   data_reorder_121_real;
  wire       [15:0]   data_reorder_121_imag;
  wire       [15:0]   data_reorder_122_real;
  wire       [15:0]   data_reorder_122_imag;
  wire       [15:0]   data_reorder_123_real;
  wire       [15:0]   data_reorder_123_imag;
  wire       [15:0]   data_reorder_124_real;
  wire       [15:0]   data_reorder_124_imag;
  wire       [15:0]   data_reorder_125_real;
  wire       [15:0]   data_reorder_125_imag;
  wire       [15:0]   data_reorder_126_real;
  wire       [15:0]   data_reorder_126_imag;
  wire       [15:0]   data_reorder_127_real;
  wire       [15:0]   data_reorder_127_imag;
  reg                 io_data_in_valid_regNext;
  reg                 current_level_willIncrement;
  wire                current_level_willClear;
  reg        [2:0]    current_level_valueNext;
  reg        [2:0]    current_level_value;
  wire                current_level_willOverflowIfInc;
  wire                current_level_willOverflow;
  reg                 null_cond_period_minus_1;
  wire                null_cond_period;
  reg        [15:0]   data_mid_0_real;
  reg        [15:0]   data_mid_0_imag;
  reg        [15:0]   data_mid_1_real;
  reg        [15:0]   data_mid_1_imag;
  reg        [15:0]   data_mid_2_real;
  reg        [15:0]   data_mid_2_imag;
  reg        [15:0]   data_mid_3_real;
  reg        [15:0]   data_mid_3_imag;
  reg        [15:0]   data_mid_4_real;
  reg        [15:0]   data_mid_4_imag;
  reg        [15:0]   data_mid_5_real;
  reg        [15:0]   data_mid_5_imag;
  reg        [15:0]   data_mid_6_real;
  reg        [15:0]   data_mid_6_imag;
  reg        [15:0]   data_mid_7_real;
  reg        [15:0]   data_mid_7_imag;
  reg        [15:0]   data_mid_8_real;
  reg        [15:0]   data_mid_8_imag;
  reg        [15:0]   data_mid_9_real;
  reg        [15:0]   data_mid_9_imag;
  reg        [15:0]   data_mid_10_real;
  reg        [15:0]   data_mid_10_imag;
  reg        [15:0]   data_mid_11_real;
  reg        [15:0]   data_mid_11_imag;
  reg        [15:0]   data_mid_12_real;
  reg        [15:0]   data_mid_12_imag;
  reg        [15:0]   data_mid_13_real;
  reg        [15:0]   data_mid_13_imag;
  reg        [15:0]   data_mid_14_real;
  reg        [15:0]   data_mid_14_imag;
  reg        [15:0]   data_mid_15_real;
  reg        [15:0]   data_mid_15_imag;
  reg        [15:0]   data_mid_16_real;
  reg        [15:0]   data_mid_16_imag;
  reg        [15:0]   data_mid_17_real;
  reg        [15:0]   data_mid_17_imag;
  reg        [15:0]   data_mid_18_real;
  reg        [15:0]   data_mid_18_imag;
  reg        [15:0]   data_mid_19_real;
  reg        [15:0]   data_mid_19_imag;
  reg        [15:0]   data_mid_20_real;
  reg        [15:0]   data_mid_20_imag;
  reg        [15:0]   data_mid_21_real;
  reg        [15:0]   data_mid_21_imag;
  reg        [15:0]   data_mid_22_real;
  reg        [15:0]   data_mid_22_imag;
  reg        [15:0]   data_mid_23_real;
  reg        [15:0]   data_mid_23_imag;
  reg        [15:0]   data_mid_24_real;
  reg        [15:0]   data_mid_24_imag;
  reg        [15:0]   data_mid_25_real;
  reg        [15:0]   data_mid_25_imag;
  reg        [15:0]   data_mid_26_real;
  reg        [15:0]   data_mid_26_imag;
  reg        [15:0]   data_mid_27_real;
  reg        [15:0]   data_mid_27_imag;
  reg        [15:0]   data_mid_28_real;
  reg        [15:0]   data_mid_28_imag;
  reg        [15:0]   data_mid_29_real;
  reg        [15:0]   data_mid_29_imag;
  reg        [15:0]   data_mid_30_real;
  reg        [15:0]   data_mid_30_imag;
  reg        [15:0]   data_mid_31_real;
  reg        [15:0]   data_mid_31_imag;
  reg        [15:0]   data_mid_32_real;
  reg        [15:0]   data_mid_32_imag;
  reg        [15:0]   data_mid_33_real;
  reg        [15:0]   data_mid_33_imag;
  reg        [15:0]   data_mid_34_real;
  reg        [15:0]   data_mid_34_imag;
  reg        [15:0]   data_mid_35_real;
  reg        [15:0]   data_mid_35_imag;
  reg        [15:0]   data_mid_36_real;
  reg        [15:0]   data_mid_36_imag;
  reg        [15:0]   data_mid_37_real;
  reg        [15:0]   data_mid_37_imag;
  reg        [15:0]   data_mid_38_real;
  reg        [15:0]   data_mid_38_imag;
  reg        [15:0]   data_mid_39_real;
  reg        [15:0]   data_mid_39_imag;
  reg        [15:0]   data_mid_40_real;
  reg        [15:0]   data_mid_40_imag;
  reg        [15:0]   data_mid_41_real;
  reg        [15:0]   data_mid_41_imag;
  reg        [15:0]   data_mid_42_real;
  reg        [15:0]   data_mid_42_imag;
  reg        [15:0]   data_mid_43_real;
  reg        [15:0]   data_mid_43_imag;
  reg        [15:0]   data_mid_44_real;
  reg        [15:0]   data_mid_44_imag;
  reg        [15:0]   data_mid_45_real;
  reg        [15:0]   data_mid_45_imag;
  reg        [15:0]   data_mid_46_real;
  reg        [15:0]   data_mid_46_imag;
  reg        [15:0]   data_mid_47_real;
  reg        [15:0]   data_mid_47_imag;
  reg        [15:0]   data_mid_48_real;
  reg        [15:0]   data_mid_48_imag;
  reg        [15:0]   data_mid_49_real;
  reg        [15:0]   data_mid_49_imag;
  reg        [15:0]   data_mid_50_real;
  reg        [15:0]   data_mid_50_imag;
  reg        [15:0]   data_mid_51_real;
  reg        [15:0]   data_mid_51_imag;
  reg        [15:0]   data_mid_52_real;
  reg        [15:0]   data_mid_52_imag;
  reg        [15:0]   data_mid_53_real;
  reg        [15:0]   data_mid_53_imag;
  reg        [15:0]   data_mid_54_real;
  reg        [15:0]   data_mid_54_imag;
  reg        [15:0]   data_mid_55_real;
  reg        [15:0]   data_mid_55_imag;
  reg        [15:0]   data_mid_56_real;
  reg        [15:0]   data_mid_56_imag;
  reg        [15:0]   data_mid_57_real;
  reg        [15:0]   data_mid_57_imag;
  reg        [15:0]   data_mid_58_real;
  reg        [15:0]   data_mid_58_imag;
  reg        [15:0]   data_mid_59_real;
  reg        [15:0]   data_mid_59_imag;
  reg        [15:0]   data_mid_60_real;
  reg        [15:0]   data_mid_60_imag;
  reg        [15:0]   data_mid_61_real;
  reg        [15:0]   data_mid_61_imag;
  reg        [15:0]   data_mid_62_real;
  reg        [15:0]   data_mid_62_imag;
  reg        [15:0]   data_mid_63_real;
  reg        [15:0]   data_mid_63_imag;
  reg        [15:0]   data_mid_64_real;
  reg        [15:0]   data_mid_64_imag;
  reg        [15:0]   data_mid_65_real;
  reg        [15:0]   data_mid_65_imag;
  reg        [15:0]   data_mid_66_real;
  reg        [15:0]   data_mid_66_imag;
  reg        [15:0]   data_mid_67_real;
  reg        [15:0]   data_mid_67_imag;
  reg        [15:0]   data_mid_68_real;
  reg        [15:0]   data_mid_68_imag;
  reg        [15:0]   data_mid_69_real;
  reg        [15:0]   data_mid_69_imag;
  reg        [15:0]   data_mid_70_real;
  reg        [15:0]   data_mid_70_imag;
  reg        [15:0]   data_mid_71_real;
  reg        [15:0]   data_mid_71_imag;
  reg        [15:0]   data_mid_72_real;
  reg        [15:0]   data_mid_72_imag;
  reg        [15:0]   data_mid_73_real;
  reg        [15:0]   data_mid_73_imag;
  reg        [15:0]   data_mid_74_real;
  reg        [15:0]   data_mid_74_imag;
  reg        [15:0]   data_mid_75_real;
  reg        [15:0]   data_mid_75_imag;
  reg        [15:0]   data_mid_76_real;
  reg        [15:0]   data_mid_76_imag;
  reg        [15:0]   data_mid_77_real;
  reg        [15:0]   data_mid_77_imag;
  reg        [15:0]   data_mid_78_real;
  reg        [15:0]   data_mid_78_imag;
  reg        [15:0]   data_mid_79_real;
  reg        [15:0]   data_mid_79_imag;
  reg        [15:0]   data_mid_80_real;
  reg        [15:0]   data_mid_80_imag;
  reg        [15:0]   data_mid_81_real;
  reg        [15:0]   data_mid_81_imag;
  reg        [15:0]   data_mid_82_real;
  reg        [15:0]   data_mid_82_imag;
  reg        [15:0]   data_mid_83_real;
  reg        [15:0]   data_mid_83_imag;
  reg        [15:0]   data_mid_84_real;
  reg        [15:0]   data_mid_84_imag;
  reg        [15:0]   data_mid_85_real;
  reg        [15:0]   data_mid_85_imag;
  reg        [15:0]   data_mid_86_real;
  reg        [15:0]   data_mid_86_imag;
  reg        [15:0]   data_mid_87_real;
  reg        [15:0]   data_mid_87_imag;
  reg        [15:0]   data_mid_88_real;
  reg        [15:0]   data_mid_88_imag;
  reg        [15:0]   data_mid_89_real;
  reg        [15:0]   data_mid_89_imag;
  reg        [15:0]   data_mid_90_real;
  reg        [15:0]   data_mid_90_imag;
  reg        [15:0]   data_mid_91_real;
  reg        [15:0]   data_mid_91_imag;
  reg        [15:0]   data_mid_92_real;
  reg        [15:0]   data_mid_92_imag;
  reg        [15:0]   data_mid_93_real;
  reg        [15:0]   data_mid_93_imag;
  reg        [15:0]   data_mid_94_real;
  reg        [15:0]   data_mid_94_imag;
  reg        [15:0]   data_mid_95_real;
  reg        [15:0]   data_mid_95_imag;
  reg        [15:0]   data_mid_96_real;
  reg        [15:0]   data_mid_96_imag;
  reg        [15:0]   data_mid_97_real;
  reg        [15:0]   data_mid_97_imag;
  reg        [15:0]   data_mid_98_real;
  reg        [15:0]   data_mid_98_imag;
  reg        [15:0]   data_mid_99_real;
  reg        [15:0]   data_mid_99_imag;
  reg        [15:0]   data_mid_100_real;
  reg        [15:0]   data_mid_100_imag;
  reg        [15:0]   data_mid_101_real;
  reg        [15:0]   data_mid_101_imag;
  reg        [15:0]   data_mid_102_real;
  reg        [15:0]   data_mid_102_imag;
  reg        [15:0]   data_mid_103_real;
  reg        [15:0]   data_mid_103_imag;
  reg        [15:0]   data_mid_104_real;
  reg        [15:0]   data_mid_104_imag;
  reg        [15:0]   data_mid_105_real;
  reg        [15:0]   data_mid_105_imag;
  reg        [15:0]   data_mid_106_real;
  reg        [15:0]   data_mid_106_imag;
  reg        [15:0]   data_mid_107_real;
  reg        [15:0]   data_mid_107_imag;
  reg        [15:0]   data_mid_108_real;
  reg        [15:0]   data_mid_108_imag;
  reg        [15:0]   data_mid_109_real;
  reg        [15:0]   data_mid_109_imag;
  reg        [15:0]   data_mid_110_real;
  reg        [15:0]   data_mid_110_imag;
  reg        [15:0]   data_mid_111_real;
  reg        [15:0]   data_mid_111_imag;
  reg        [15:0]   data_mid_112_real;
  reg        [15:0]   data_mid_112_imag;
  reg        [15:0]   data_mid_113_real;
  reg        [15:0]   data_mid_113_imag;
  reg        [15:0]   data_mid_114_real;
  reg        [15:0]   data_mid_114_imag;
  reg        [15:0]   data_mid_115_real;
  reg        [15:0]   data_mid_115_imag;
  reg        [15:0]   data_mid_116_real;
  reg        [15:0]   data_mid_116_imag;
  reg        [15:0]   data_mid_117_real;
  reg        [15:0]   data_mid_117_imag;
  reg        [15:0]   data_mid_118_real;
  reg        [15:0]   data_mid_118_imag;
  reg        [15:0]   data_mid_119_real;
  reg        [15:0]   data_mid_119_imag;
  reg        [15:0]   data_mid_120_real;
  reg        [15:0]   data_mid_120_imag;
  reg        [15:0]   data_mid_121_real;
  reg        [15:0]   data_mid_121_imag;
  reg        [15:0]   data_mid_122_real;
  reg        [15:0]   data_mid_122_imag;
  reg        [15:0]   data_mid_123_real;
  reg        [15:0]   data_mid_123_imag;
  reg        [15:0]   data_mid_124_real;
  reg        [15:0]   data_mid_124_imag;
  reg        [15:0]   data_mid_125_real;
  reg        [15:0]   data_mid_125_imag;
  reg        [15:0]   data_mid_126_real;
  reg        [15:0]   data_mid_126_imag;
  reg        [15:0]   data_mid_127_real;
  reg        [15:0]   data_mid_127_imag;
  wire       [31:0]   _zz_1;
  wire       [31:0]   _zz_2;
  wire       [31:0]   _zz_3;
  wire       [0:0]    _zz_4;
  wire       [0:0]    _zz_5;
  wire       [31:0]   _zz_6;
  wire       [31:0]   _zz_7;
  wire       [31:0]   _zz_8;
  wire       [0:0]    _zz_9;
  wire       [0:0]    _zz_10;
  wire       [31:0]   _zz_11;
  wire       [31:0]   _zz_12;
  wire       [31:0]   _zz_13;
  wire       [0:0]    _zz_14;
  wire       [0:0]    _zz_15;
  wire       [31:0]   _zz_16;
  wire       [31:0]   _zz_17;
  wire       [31:0]   _zz_18;
  wire       [0:0]    _zz_19;
  wire       [0:0]    _zz_20;
  wire       [31:0]   _zz_21;
  wire       [31:0]   _zz_22;
  wire       [31:0]   _zz_23;
  wire       [0:0]    _zz_24;
  wire       [0:0]    _zz_25;
  wire       [31:0]   _zz_26;
  wire       [31:0]   _zz_27;
  wire       [31:0]   _zz_28;
  wire       [0:0]    _zz_29;
  wire       [0:0]    _zz_30;
  wire       [31:0]   _zz_31;
  wire       [31:0]   _zz_32;
  wire       [31:0]   _zz_33;
  wire       [0:0]    _zz_34;
  wire       [0:0]    _zz_35;
  wire       [31:0]   _zz_36;
  wire       [31:0]   _zz_37;
  wire       [31:0]   _zz_38;
  wire       [0:0]    _zz_39;
  wire       [0:0]    _zz_40;
  wire       [31:0]   _zz_41;
  wire       [31:0]   _zz_42;
  wire       [31:0]   _zz_43;
  wire       [0:0]    _zz_44;
  wire       [0:0]    _zz_45;
  wire       [31:0]   _zz_46;
  wire       [31:0]   _zz_47;
  wire       [31:0]   _zz_48;
  wire       [0:0]    _zz_49;
  wire       [0:0]    _zz_50;
  wire       [31:0]   _zz_51;
  wire       [31:0]   _zz_52;
  wire       [31:0]   _zz_53;
  wire       [0:0]    _zz_54;
  wire       [0:0]    _zz_55;
  wire       [31:0]   _zz_56;
  wire       [31:0]   _zz_57;
  wire       [31:0]   _zz_58;
  wire       [0:0]    _zz_59;
  wire       [0:0]    _zz_60;
  wire       [31:0]   _zz_61;
  wire       [31:0]   _zz_62;
  wire       [31:0]   _zz_63;
  wire       [0:0]    _zz_64;
  wire       [0:0]    _zz_65;
  wire       [31:0]   _zz_66;
  wire       [31:0]   _zz_67;
  wire       [31:0]   _zz_68;
  wire       [0:0]    _zz_69;
  wire       [0:0]    _zz_70;
  wire       [31:0]   _zz_71;
  wire       [31:0]   _zz_72;
  wire       [31:0]   _zz_73;
  wire       [0:0]    _zz_74;
  wire       [0:0]    _zz_75;
  wire       [31:0]   _zz_76;
  wire       [31:0]   _zz_77;
  wire       [31:0]   _zz_78;
  wire       [0:0]    _zz_79;
  wire       [0:0]    _zz_80;
  wire       [31:0]   _zz_81;
  wire       [31:0]   _zz_82;
  wire       [31:0]   _zz_83;
  wire       [0:0]    _zz_84;
  wire       [0:0]    _zz_85;
  wire       [31:0]   _zz_86;
  wire       [31:0]   _zz_87;
  wire       [31:0]   _zz_88;
  wire       [0:0]    _zz_89;
  wire       [0:0]    _zz_90;
  wire       [31:0]   _zz_91;
  wire       [31:0]   _zz_92;
  wire       [31:0]   _zz_93;
  wire       [0:0]    _zz_94;
  wire       [0:0]    _zz_95;
  wire       [31:0]   _zz_96;
  wire       [31:0]   _zz_97;
  wire       [31:0]   _zz_98;
  wire       [0:0]    _zz_99;
  wire       [0:0]    _zz_100;
  wire       [31:0]   _zz_101;
  wire       [31:0]   _zz_102;
  wire       [31:0]   _zz_103;
  wire       [0:0]    _zz_104;
  wire       [0:0]    _zz_105;
  wire       [31:0]   _zz_106;
  wire       [31:0]   _zz_107;
  wire       [31:0]   _zz_108;
  wire       [0:0]    _zz_109;
  wire       [0:0]    _zz_110;
  wire       [31:0]   _zz_111;
  wire       [31:0]   _zz_112;
  wire       [31:0]   _zz_113;
  wire       [0:0]    _zz_114;
  wire       [0:0]    _zz_115;
  wire       [31:0]   _zz_116;
  wire       [31:0]   _zz_117;
  wire       [31:0]   _zz_118;
  wire       [0:0]    _zz_119;
  wire       [0:0]    _zz_120;
  wire       [31:0]   _zz_121;
  wire       [31:0]   _zz_122;
  wire       [31:0]   _zz_123;
  wire       [0:0]    _zz_124;
  wire       [0:0]    _zz_125;
  wire       [31:0]   _zz_126;
  wire       [31:0]   _zz_127;
  wire       [31:0]   _zz_128;
  wire       [0:0]    _zz_129;
  wire       [0:0]    _zz_130;
  wire       [31:0]   _zz_131;
  wire       [31:0]   _zz_132;
  wire       [31:0]   _zz_133;
  wire       [0:0]    _zz_134;
  wire       [0:0]    _zz_135;
  wire       [31:0]   _zz_136;
  wire       [31:0]   _zz_137;
  wire       [31:0]   _zz_138;
  wire       [0:0]    _zz_139;
  wire       [0:0]    _zz_140;
  wire       [31:0]   _zz_141;
  wire       [31:0]   _zz_142;
  wire       [31:0]   _zz_143;
  wire       [0:0]    _zz_144;
  wire       [0:0]    _zz_145;
  wire       [31:0]   _zz_146;
  wire       [31:0]   _zz_147;
  wire       [31:0]   _zz_148;
  wire       [0:0]    _zz_149;
  wire       [0:0]    _zz_150;
  wire       [31:0]   _zz_151;
  wire       [31:0]   _zz_152;
  wire       [31:0]   _zz_153;
  wire       [0:0]    _zz_154;
  wire       [0:0]    _zz_155;
  wire       [31:0]   _zz_156;
  wire       [31:0]   _zz_157;
  wire       [31:0]   _zz_158;
  wire       [0:0]    _zz_159;
  wire       [0:0]    _zz_160;
  wire       [31:0]   _zz_161;
  wire       [31:0]   _zz_162;
  wire       [31:0]   _zz_163;
  wire       [0:0]    _zz_164;
  wire       [0:0]    _zz_165;
  wire       [31:0]   _zz_166;
  wire       [31:0]   _zz_167;
  wire       [31:0]   _zz_168;
  wire       [0:0]    _zz_169;
  wire       [0:0]    _zz_170;
  wire       [31:0]   _zz_171;
  wire       [31:0]   _zz_172;
  wire       [31:0]   _zz_173;
  wire       [0:0]    _zz_174;
  wire       [0:0]    _zz_175;
  wire       [31:0]   _zz_176;
  wire       [31:0]   _zz_177;
  wire       [31:0]   _zz_178;
  wire       [0:0]    _zz_179;
  wire       [0:0]    _zz_180;
  wire       [31:0]   _zz_181;
  wire       [31:0]   _zz_182;
  wire       [31:0]   _zz_183;
  wire       [0:0]    _zz_184;
  wire       [0:0]    _zz_185;
  wire       [31:0]   _zz_186;
  wire       [31:0]   _zz_187;
  wire       [31:0]   _zz_188;
  wire       [0:0]    _zz_189;
  wire       [0:0]    _zz_190;
  wire       [31:0]   _zz_191;
  wire       [31:0]   _zz_192;
  wire       [31:0]   _zz_193;
  wire       [0:0]    _zz_194;
  wire       [0:0]    _zz_195;
  wire       [31:0]   _zz_196;
  wire       [31:0]   _zz_197;
  wire       [31:0]   _zz_198;
  wire       [0:0]    _zz_199;
  wire       [0:0]    _zz_200;
  wire       [31:0]   _zz_201;
  wire       [31:0]   _zz_202;
  wire       [31:0]   _zz_203;
  wire       [0:0]    _zz_204;
  wire       [0:0]    _zz_205;
  wire       [31:0]   _zz_206;
  wire       [31:0]   _zz_207;
  wire       [31:0]   _zz_208;
  wire       [0:0]    _zz_209;
  wire       [0:0]    _zz_210;
  wire       [31:0]   _zz_211;
  wire       [31:0]   _zz_212;
  wire       [31:0]   _zz_213;
  wire       [0:0]    _zz_214;
  wire       [0:0]    _zz_215;
  wire       [31:0]   _zz_216;
  wire       [31:0]   _zz_217;
  wire       [31:0]   _zz_218;
  wire       [0:0]    _zz_219;
  wire       [0:0]    _zz_220;
  wire       [31:0]   _zz_221;
  wire       [31:0]   _zz_222;
  wire       [31:0]   _zz_223;
  wire       [0:0]    _zz_224;
  wire       [0:0]    _zz_225;
  wire       [31:0]   _zz_226;
  wire       [31:0]   _zz_227;
  wire       [31:0]   _zz_228;
  wire       [0:0]    _zz_229;
  wire       [0:0]    _zz_230;
  wire       [31:0]   _zz_231;
  wire       [31:0]   _zz_232;
  wire       [31:0]   _zz_233;
  wire       [0:0]    _zz_234;
  wire       [0:0]    _zz_235;
  wire       [31:0]   _zz_236;
  wire       [31:0]   _zz_237;
  wire       [31:0]   _zz_238;
  wire       [0:0]    _zz_239;
  wire       [0:0]    _zz_240;
  wire       [31:0]   _zz_241;
  wire       [31:0]   _zz_242;
  wire       [31:0]   _zz_243;
  wire       [0:0]    _zz_244;
  wire       [0:0]    _zz_245;
  wire       [31:0]   _zz_246;
  wire       [31:0]   _zz_247;
  wire       [31:0]   _zz_248;
  wire       [0:0]    _zz_249;
  wire       [0:0]    _zz_250;
  wire       [31:0]   _zz_251;
  wire       [31:0]   _zz_252;
  wire       [31:0]   _zz_253;
  wire       [0:0]    _zz_254;
  wire       [0:0]    _zz_255;
  wire       [31:0]   _zz_256;
  wire       [31:0]   _zz_257;
  wire       [31:0]   _zz_258;
  wire       [0:0]    _zz_259;
  wire       [0:0]    _zz_260;
  wire       [31:0]   _zz_261;
  wire       [31:0]   _zz_262;
  wire       [31:0]   _zz_263;
  wire       [0:0]    _zz_264;
  wire       [0:0]    _zz_265;
  wire       [31:0]   _zz_266;
  wire       [31:0]   _zz_267;
  wire       [31:0]   _zz_268;
  wire       [0:0]    _zz_269;
  wire       [0:0]    _zz_270;
  wire       [31:0]   _zz_271;
  wire       [31:0]   _zz_272;
  wire       [31:0]   _zz_273;
  wire       [0:0]    _zz_274;
  wire       [0:0]    _zz_275;
  wire       [31:0]   _zz_276;
  wire       [31:0]   _zz_277;
  wire       [31:0]   _zz_278;
  wire       [0:0]    _zz_279;
  wire       [0:0]    _zz_280;
  wire       [31:0]   _zz_281;
  wire       [31:0]   _zz_282;
  wire       [31:0]   _zz_283;
  wire       [0:0]    _zz_284;
  wire       [0:0]    _zz_285;
  wire       [31:0]   _zz_286;
  wire       [31:0]   _zz_287;
  wire       [31:0]   _zz_288;
  wire       [0:0]    _zz_289;
  wire       [0:0]    _zz_290;
  wire       [31:0]   _zz_291;
  wire       [31:0]   _zz_292;
  wire       [31:0]   _zz_293;
  wire       [0:0]    _zz_294;
  wire       [0:0]    _zz_295;
  wire       [31:0]   _zz_296;
  wire       [31:0]   _zz_297;
  wire       [31:0]   _zz_298;
  wire       [0:0]    _zz_299;
  wire       [0:0]    _zz_300;
  wire       [31:0]   _zz_301;
  wire       [31:0]   _zz_302;
  wire       [31:0]   _zz_303;
  wire       [0:0]    _zz_304;
  wire       [0:0]    _zz_305;
  wire       [31:0]   _zz_306;
  wire       [31:0]   _zz_307;
  wire       [31:0]   _zz_308;
  wire       [0:0]    _zz_309;
  wire       [0:0]    _zz_310;
  wire       [31:0]   _zz_311;
  wire       [31:0]   _zz_312;
  wire       [31:0]   _zz_313;
  wire       [0:0]    _zz_314;
  wire       [0:0]    _zz_315;
  wire       [31:0]   _zz_316;
  wire       [31:0]   _zz_317;
  wire       [31:0]   _zz_318;
  wire       [0:0]    _zz_319;
  wire       [0:0]    _zz_320;
  wire       [31:0]   _zz_321;
  wire       [31:0]   _zz_322;
  wire       [31:0]   _zz_323;
  wire       [0:0]    _zz_324;
  wire       [0:0]    _zz_325;
  wire       [31:0]   _zz_326;
  wire       [31:0]   _zz_327;
  wire       [31:0]   _zz_328;
  wire       [0:0]    _zz_329;
  wire       [0:0]    _zz_330;
  wire       [31:0]   _zz_331;
  wire       [31:0]   _zz_332;
  wire       [31:0]   _zz_333;
  wire       [0:0]    _zz_334;
  wire       [0:0]    _zz_335;
  wire       [31:0]   _zz_336;
  wire       [31:0]   _zz_337;
  wire       [31:0]   _zz_338;
  wire       [0:0]    _zz_339;
  wire       [0:0]    _zz_340;
  wire       [31:0]   _zz_341;
  wire       [31:0]   _zz_342;
  wire       [31:0]   _zz_343;
  wire       [0:0]    _zz_344;
  wire       [0:0]    _zz_345;
  wire       [31:0]   _zz_346;
  wire       [31:0]   _zz_347;
  wire       [31:0]   _zz_348;
  wire       [0:0]    _zz_349;
  wire       [0:0]    _zz_350;
  wire       [31:0]   _zz_351;
  wire       [31:0]   _zz_352;
  wire       [31:0]   _zz_353;
  wire       [0:0]    _zz_354;
  wire       [0:0]    _zz_355;
  wire       [31:0]   _zz_356;
  wire       [31:0]   _zz_357;
  wire       [31:0]   _zz_358;
  wire       [0:0]    _zz_359;
  wire       [0:0]    _zz_360;
  wire       [31:0]   _zz_361;
  wire       [31:0]   _zz_362;
  wire       [31:0]   _zz_363;
  wire       [0:0]    _zz_364;
  wire       [0:0]    _zz_365;
  wire       [31:0]   _zz_366;
  wire       [31:0]   _zz_367;
  wire       [31:0]   _zz_368;
  wire       [0:0]    _zz_369;
  wire       [0:0]    _zz_370;
  wire       [31:0]   _zz_371;
  wire       [31:0]   _zz_372;
  wire       [31:0]   _zz_373;
  wire       [0:0]    _zz_374;
  wire       [0:0]    _zz_375;
  wire       [31:0]   _zz_376;
  wire       [31:0]   _zz_377;
  wire       [31:0]   _zz_378;
  wire       [0:0]    _zz_379;
  wire       [0:0]    _zz_380;
  wire       [31:0]   _zz_381;
  wire       [31:0]   _zz_382;
  wire       [31:0]   _zz_383;
  wire       [0:0]    _zz_384;
  wire       [0:0]    _zz_385;
  wire       [31:0]   _zz_386;
  wire       [31:0]   _zz_387;
  wire       [31:0]   _zz_388;
  wire       [0:0]    _zz_389;
  wire       [0:0]    _zz_390;
  wire       [31:0]   _zz_391;
  wire       [31:0]   _zz_392;
  wire       [31:0]   _zz_393;
  wire       [0:0]    _zz_394;
  wire       [0:0]    _zz_395;
  wire       [31:0]   _zz_396;
  wire       [31:0]   _zz_397;
  wire       [31:0]   _zz_398;
  wire       [0:0]    _zz_399;
  wire       [0:0]    _zz_400;
  wire       [31:0]   _zz_401;
  wire       [31:0]   _zz_402;
  wire       [31:0]   _zz_403;
  wire       [0:0]    _zz_404;
  wire       [0:0]    _zz_405;
  wire       [31:0]   _zz_406;
  wire       [31:0]   _zz_407;
  wire       [31:0]   _zz_408;
  wire       [0:0]    _zz_409;
  wire       [0:0]    _zz_410;
  wire       [31:0]   _zz_411;
  wire       [31:0]   _zz_412;
  wire       [31:0]   _zz_413;
  wire       [0:0]    _zz_414;
  wire       [0:0]    _zz_415;
  wire       [31:0]   _zz_416;
  wire       [31:0]   _zz_417;
  wire       [31:0]   _zz_418;
  wire       [0:0]    _zz_419;
  wire       [0:0]    _zz_420;
  wire       [31:0]   _zz_421;
  wire       [31:0]   _zz_422;
  wire       [31:0]   _zz_423;
  wire       [0:0]    _zz_424;
  wire       [0:0]    _zz_425;
  wire       [31:0]   _zz_426;
  wire       [31:0]   _zz_427;
  wire       [31:0]   _zz_428;
  wire       [0:0]    _zz_429;
  wire       [0:0]    _zz_430;
  wire       [31:0]   _zz_431;
  wire       [31:0]   _zz_432;
  wire       [31:0]   _zz_433;
  wire       [0:0]    _zz_434;
  wire       [0:0]    _zz_435;
  wire       [31:0]   _zz_436;
  wire       [31:0]   _zz_437;
  wire       [31:0]   _zz_438;
  wire       [0:0]    _zz_439;
  wire       [0:0]    _zz_440;
  wire       [31:0]   _zz_441;
  wire       [31:0]   _zz_442;
  wire       [31:0]   _zz_443;
  wire       [0:0]    _zz_444;
  wire       [0:0]    _zz_445;
  wire       [31:0]   _zz_446;
  wire       [31:0]   _zz_447;
  wire       [31:0]   _zz_448;
  wire       [0:0]    _zz_449;
  wire       [0:0]    _zz_450;
  wire       [31:0]   _zz_451;
  wire       [31:0]   _zz_452;
  wire       [31:0]   _zz_453;
  wire       [0:0]    _zz_454;
  wire       [0:0]    _zz_455;
  wire       [31:0]   _zz_456;
  wire       [31:0]   _zz_457;
  wire       [31:0]   _zz_458;
  wire       [0:0]    _zz_459;
  wire       [0:0]    _zz_460;
  wire       [31:0]   _zz_461;
  wire       [31:0]   _zz_462;
  wire       [31:0]   _zz_463;
  wire       [0:0]    _zz_464;
  wire       [0:0]    _zz_465;
  wire       [31:0]   _zz_466;
  wire       [31:0]   _zz_467;
  wire       [31:0]   _zz_468;
  wire       [0:0]    _zz_469;
  wire       [0:0]    _zz_470;
  wire       [31:0]   _zz_471;
  wire       [31:0]   _zz_472;
  wire       [31:0]   _zz_473;
  wire       [0:0]    _zz_474;
  wire       [0:0]    _zz_475;
  wire       [31:0]   _zz_476;
  wire       [31:0]   _zz_477;
  wire       [31:0]   _zz_478;
  wire       [0:0]    _zz_479;
  wire       [0:0]    _zz_480;
  wire       [31:0]   _zz_481;
  wire       [31:0]   _zz_482;
  wire       [31:0]   _zz_483;
  wire       [0:0]    _zz_484;
  wire       [0:0]    _zz_485;
  wire       [31:0]   _zz_486;
  wire       [31:0]   _zz_487;
  wire       [31:0]   _zz_488;
  wire       [0:0]    _zz_489;
  wire       [0:0]    _zz_490;
  wire       [31:0]   _zz_491;
  wire       [31:0]   _zz_492;
  wire       [31:0]   _zz_493;
  wire       [0:0]    _zz_494;
  wire       [0:0]    _zz_495;
  wire       [31:0]   _zz_496;
  wire       [31:0]   _zz_497;
  wire       [31:0]   _zz_498;
  wire       [0:0]    _zz_499;
  wire       [0:0]    _zz_500;
  wire       [31:0]   _zz_501;
  wire       [31:0]   _zz_502;
  wire       [31:0]   _zz_503;
  wire       [0:0]    _zz_504;
  wire       [0:0]    _zz_505;
  wire       [31:0]   _zz_506;
  wire       [31:0]   _zz_507;
  wire       [31:0]   _zz_508;
  wire       [0:0]    _zz_509;
  wire       [0:0]    _zz_510;
  wire       [31:0]   _zz_511;
  wire       [31:0]   _zz_512;
  wire       [31:0]   _zz_513;
  wire       [0:0]    _zz_514;
  wire       [0:0]    _zz_515;
  wire       [31:0]   _zz_516;
  wire       [31:0]   _zz_517;
  wire       [31:0]   _zz_518;
  wire       [0:0]    _zz_519;
  wire       [0:0]    _zz_520;
  wire       [31:0]   _zz_521;
  wire       [31:0]   _zz_522;
  wire       [31:0]   _zz_523;
  wire       [0:0]    _zz_524;
  wire       [0:0]    _zz_525;
  wire       [31:0]   _zz_526;
  wire       [31:0]   _zz_527;
  wire       [31:0]   _zz_528;
  wire       [0:0]    _zz_529;
  wire       [0:0]    _zz_530;
  wire       [31:0]   _zz_531;
  wire       [31:0]   _zz_532;
  wire       [31:0]   _zz_533;
  wire       [0:0]    _zz_534;
  wire       [0:0]    _zz_535;
  wire       [31:0]   _zz_536;
  wire       [31:0]   _zz_537;
  wire       [31:0]   _zz_538;
  wire       [0:0]    _zz_539;
  wire       [0:0]    _zz_540;
  wire       [31:0]   _zz_541;
  wire       [31:0]   _zz_542;
  wire       [31:0]   _zz_543;
  wire       [0:0]    _zz_544;
  wire       [0:0]    _zz_545;
  wire       [31:0]   _zz_546;
  wire       [31:0]   _zz_547;
  wire       [31:0]   _zz_548;
  wire       [0:0]    _zz_549;
  wire       [0:0]    _zz_550;
  wire       [31:0]   _zz_551;
  wire       [31:0]   _zz_552;
  wire       [31:0]   _zz_553;
  wire       [0:0]    _zz_554;
  wire       [0:0]    _zz_555;
  wire       [31:0]   _zz_556;
  wire       [31:0]   _zz_557;
  wire       [31:0]   _zz_558;
  wire       [0:0]    _zz_559;
  wire       [0:0]    _zz_560;
  wire       [31:0]   _zz_561;
  wire       [31:0]   _zz_562;
  wire       [31:0]   _zz_563;
  wire       [0:0]    _zz_564;
  wire       [0:0]    _zz_565;
  wire       [31:0]   _zz_566;
  wire       [31:0]   _zz_567;
  wire       [31:0]   _zz_568;
  wire       [0:0]    _zz_569;
  wire       [0:0]    _zz_570;
  wire       [31:0]   _zz_571;
  wire       [31:0]   _zz_572;
  wire       [31:0]   _zz_573;
  wire       [0:0]    _zz_574;
  wire       [0:0]    _zz_575;
  wire       [31:0]   _zz_576;
  wire       [31:0]   _zz_577;
  wire       [31:0]   _zz_578;
  wire       [0:0]    _zz_579;
  wire       [0:0]    _zz_580;
  wire       [31:0]   _zz_581;
  wire       [31:0]   _zz_582;
  wire       [31:0]   _zz_583;
  wire       [0:0]    _zz_584;
  wire       [0:0]    _zz_585;
  wire       [31:0]   _zz_586;
  wire       [31:0]   _zz_587;
  wire       [31:0]   _zz_588;
  wire       [0:0]    _zz_589;
  wire       [0:0]    _zz_590;
  wire       [31:0]   _zz_591;
  wire       [31:0]   _zz_592;
  wire       [31:0]   _zz_593;
  wire       [0:0]    _zz_594;
  wire       [0:0]    _zz_595;
  wire       [31:0]   _zz_596;
  wire       [31:0]   _zz_597;
  wire       [31:0]   _zz_598;
  wire       [0:0]    _zz_599;
  wire       [0:0]    _zz_600;
  wire       [31:0]   _zz_601;
  wire       [31:0]   _zz_602;
  wire       [31:0]   _zz_603;
  wire       [0:0]    _zz_604;
  wire       [0:0]    _zz_605;
  wire       [31:0]   _zz_606;
  wire       [31:0]   _zz_607;
  wire       [31:0]   _zz_608;
  wire       [0:0]    _zz_609;
  wire       [0:0]    _zz_610;
  wire       [31:0]   _zz_611;
  wire       [31:0]   _zz_612;
  wire       [31:0]   _zz_613;
  wire       [0:0]    _zz_614;
  wire       [0:0]    _zz_615;
  wire       [31:0]   _zz_616;
  wire       [31:0]   _zz_617;
  wire       [31:0]   _zz_618;
  wire       [0:0]    _zz_619;
  wire       [0:0]    _zz_620;
  wire       [31:0]   _zz_621;
  wire       [31:0]   _zz_622;
  wire       [31:0]   _zz_623;
  wire       [0:0]    _zz_624;
  wire       [0:0]    _zz_625;
  wire       [31:0]   _zz_626;
  wire       [31:0]   _zz_627;
  wire       [31:0]   _zz_628;
  wire       [0:0]    _zz_629;
  wire       [0:0]    _zz_630;
  wire       [31:0]   _zz_631;
  wire       [31:0]   _zz_632;
  wire       [31:0]   _zz_633;
  wire       [0:0]    _zz_634;
  wire       [0:0]    _zz_635;
  wire       [31:0]   _zz_636;
  wire       [31:0]   _zz_637;
  wire       [31:0]   _zz_638;
  wire       [0:0]    _zz_639;
  wire       [0:0]    _zz_640;
  wire       [31:0]   _zz_641;
  wire       [31:0]   _zz_642;
  wire       [31:0]   _zz_643;
  wire       [0:0]    _zz_644;
  wire       [0:0]    _zz_645;
  wire       [31:0]   _zz_646;
  wire       [31:0]   _zz_647;
  wire       [31:0]   _zz_648;
  wire       [0:0]    _zz_649;
  wire       [0:0]    _zz_650;
  wire       [31:0]   _zz_651;
  wire       [31:0]   _zz_652;
  wire       [31:0]   _zz_653;
  wire       [0:0]    _zz_654;
  wire       [0:0]    _zz_655;
  wire       [31:0]   _zz_656;
  wire       [31:0]   _zz_657;
  wire       [31:0]   _zz_658;
  wire       [0:0]    _zz_659;
  wire       [0:0]    _zz_660;
  wire       [31:0]   _zz_661;
  wire       [31:0]   _zz_662;
  wire       [31:0]   _zz_663;
  wire       [0:0]    _zz_664;
  wire       [0:0]    _zz_665;
  wire       [31:0]   _zz_666;
  wire       [31:0]   _zz_667;
  wire       [31:0]   _zz_668;
  wire       [0:0]    _zz_669;
  wire       [0:0]    _zz_670;
  wire       [31:0]   _zz_671;
  wire       [31:0]   _zz_672;
  wire       [31:0]   _zz_673;
  wire       [0:0]    _zz_674;
  wire       [0:0]    _zz_675;
  wire       [31:0]   _zz_676;
  wire       [31:0]   _zz_677;
  wire       [31:0]   _zz_678;
  wire       [0:0]    _zz_679;
  wire       [0:0]    _zz_680;
  wire       [31:0]   _zz_681;
  wire       [31:0]   _zz_682;
  wire       [31:0]   _zz_683;
  wire       [0:0]    _zz_684;
  wire       [0:0]    _zz_685;
  wire       [31:0]   _zz_686;
  wire       [31:0]   _zz_687;
  wire       [31:0]   _zz_688;
  wire       [0:0]    _zz_689;
  wire       [0:0]    _zz_690;
  wire       [31:0]   _zz_691;
  wire       [31:0]   _zz_692;
  wire       [31:0]   _zz_693;
  wire       [0:0]    _zz_694;
  wire       [0:0]    _zz_695;
  wire       [31:0]   _zz_696;
  wire       [31:0]   _zz_697;
  wire       [31:0]   _zz_698;
  wire       [0:0]    _zz_699;
  wire       [0:0]    _zz_700;
  wire       [31:0]   _zz_701;
  wire       [31:0]   _zz_702;
  wire       [31:0]   _zz_703;
  wire       [0:0]    _zz_704;
  wire       [0:0]    _zz_705;
  wire       [31:0]   _zz_706;
  wire       [31:0]   _zz_707;
  wire       [31:0]   _zz_708;
  wire       [0:0]    _zz_709;
  wire       [0:0]    _zz_710;
  wire       [31:0]   _zz_711;
  wire       [31:0]   _zz_712;
  wire       [31:0]   _zz_713;
  wire       [0:0]    _zz_714;
  wire       [0:0]    _zz_715;
  wire       [31:0]   _zz_716;
  wire       [31:0]   _zz_717;
  wire       [31:0]   _zz_718;
  wire       [0:0]    _zz_719;
  wire       [0:0]    _zz_720;
  wire       [31:0]   _zz_721;
  wire       [31:0]   _zz_722;
  wire       [31:0]   _zz_723;
  wire       [0:0]    _zz_724;
  wire       [0:0]    _zz_725;
  wire       [31:0]   _zz_726;
  wire       [31:0]   _zz_727;
  wire       [31:0]   _zz_728;
  wire       [0:0]    _zz_729;
  wire       [0:0]    _zz_730;
  wire       [31:0]   _zz_731;
  wire       [31:0]   _zz_732;
  wire       [31:0]   _zz_733;
  wire       [0:0]    _zz_734;
  wire       [0:0]    _zz_735;
  wire       [31:0]   _zz_736;
  wire       [31:0]   _zz_737;
  wire       [31:0]   _zz_738;
  wire       [0:0]    _zz_739;
  wire       [0:0]    _zz_740;
  wire       [31:0]   _zz_741;
  wire       [31:0]   _zz_742;
  wire       [31:0]   _zz_743;
  wire       [0:0]    _zz_744;
  wire       [0:0]    _zz_745;
  wire       [31:0]   _zz_746;
  wire       [31:0]   _zz_747;
  wire       [31:0]   _zz_748;
  wire       [0:0]    _zz_749;
  wire       [0:0]    _zz_750;
  wire       [31:0]   _zz_751;
  wire       [31:0]   _zz_752;
  wire       [31:0]   _zz_753;
  wire       [0:0]    _zz_754;
  wire       [0:0]    _zz_755;
  wire       [31:0]   _zz_756;
  wire       [31:0]   _zz_757;
  wire       [31:0]   _zz_758;
  wire       [0:0]    _zz_759;
  wire       [0:0]    _zz_760;
  wire       [31:0]   _zz_761;
  wire       [31:0]   _zz_762;
  wire       [31:0]   _zz_763;
  wire       [0:0]    _zz_764;
  wire       [0:0]    _zz_765;
  wire       [31:0]   _zz_766;
  wire       [31:0]   _zz_767;
  wire       [31:0]   _zz_768;
  wire       [0:0]    _zz_769;
  wire       [0:0]    _zz_770;
  wire       [31:0]   _zz_771;
  wire       [31:0]   _zz_772;
  wire       [31:0]   _zz_773;
  wire       [0:0]    _zz_774;
  wire       [0:0]    _zz_775;
  wire       [31:0]   _zz_776;
  wire       [31:0]   _zz_777;
  wire       [31:0]   _zz_778;
  wire       [0:0]    _zz_779;
  wire       [0:0]    _zz_780;
  wire       [31:0]   _zz_781;
  wire       [31:0]   _zz_782;
  wire       [31:0]   _zz_783;
  wire       [0:0]    _zz_784;
  wire       [0:0]    _zz_785;
  wire       [31:0]   _zz_786;
  wire       [31:0]   _zz_787;
  wire       [31:0]   _zz_788;
  wire       [0:0]    _zz_789;
  wire       [0:0]    _zz_790;
  wire       [31:0]   _zz_791;
  wire       [31:0]   _zz_792;
  wire       [31:0]   _zz_793;
  wire       [0:0]    _zz_794;
  wire       [0:0]    _zz_795;
  wire       [31:0]   _zz_796;
  wire       [31:0]   _zz_797;
  wire       [31:0]   _zz_798;
  wire       [0:0]    _zz_799;
  wire       [0:0]    _zz_800;
  wire       [31:0]   _zz_801;
  wire       [31:0]   _zz_802;
  wire       [31:0]   _zz_803;
  wire       [0:0]    _zz_804;
  wire       [0:0]    _zz_805;
  wire       [31:0]   _zz_806;
  wire       [31:0]   _zz_807;
  wire       [31:0]   _zz_808;
  wire       [0:0]    _zz_809;
  wire       [0:0]    _zz_810;
  wire       [31:0]   _zz_811;
  wire       [31:0]   _zz_812;
  wire       [31:0]   _zz_813;
  wire       [0:0]    _zz_814;
  wire       [0:0]    _zz_815;
  wire       [31:0]   _zz_816;
  wire       [31:0]   _zz_817;
  wire       [31:0]   _zz_818;
  wire       [0:0]    _zz_819;
  wire       [0:0]    _zz_820;
  wire       [31:0]   _zz_821;
  wire       [31:0]   _zz_822;
  wire       [31:0]   _zz_823;
  wire       [0:0]    _zz_824;
  wire       [0:0]    _zz_825;
  wire       [31:0]   _zz_826;
  wire       [31:0]   _zz_827;
  wire       [31:0]   _zz_828;
  wire       [0:0]    _zz_829;
  wire       [0:0]    _zz_830;
  wire       [31:0]   _zz_831;
  wire       [31:0]   _zz_832;
  wire       [31:0]   _zz_833;
  wire       [0:0]    _zz_834;
  wire       [0:0]    _zz_835;
  wire       [31:0]   _zz_836;
  wire       [31:0]   _zz_837;
  wire       [31:0]   _zz_838;
  wire       [0:0]    _zz_839;
  wire       [0:0]    _zz_840;
  wire       [31:0]   _zz_841;
  wire       [31:0]   _zz_842;
  wire       [31:0]   _zz_843;
  wire       [0:0]    _zz_844;
  wire       [0:0]    _zz_845;
  wire       [31:0]   _zz_846;
  wire       [31:0]   _zz_847;
  wire       [31:0]   _zz_848;
  wire       [0:0]    _zz_849;
  wire       [0:0]    _zz_850;
  wire       [31:0]   _zz_851;
  wire       [31:0]   _zz_852;
  wire       [31:0]   _zz_853;
  wire       [0:0]    _zz_854;
  wire       [0:0]    _zz_855;
  wire       [31:0]   _zz_856;
  wire       [31:0]   _zz_857;
  wire       [31:0]   _zz_858;
  wire       [0:0]    _zz_859;
  wire       [0:0]    _zz_860;
  wire       [31:0]   _zz_861;
  wire       [31:0]   _zz_862;
  wire       [31:0]   _zz_863;
  wire       [0:0]    _zz_864;
  wire       [0:0]    _zz_865;
  wire       [31:0]   _zz_866;
  wire       [31:0]   _zz_867;
  wire       [31:0]   _zz_868;
  wire       [0:0]    _zz_869;
  wire       [0:0]    _zz_870;
  wire       [31:0]   _zz_871;
  wire       [31:0]   _zz_872;
  wire       [31:0]   _zz_873;
  wire       [0:0]    _zz_874;
  wire       [0:0]    _zz_875;
  wire       [31:0]   _zz_876;
  wire       [31:0]   _zz_877;
  wire       [31:0]   _zz_878;
  wire       [0:0]    _zz_879;
  wire       [0:0]    _zz_880;
  wire       [31:0]   _zz_881;
  wire       [31:0]   _zz_882;
  wire       [31:0]   _zz_883;
  wire       [0:0]    _zz_884;
  wire       [0:0]    _zz_885;
  wire       [31:0]   _zz_886;
  wire       [31:0]   _zz_887;
  wire       [31:0]   _zz_888;
  wire       [0:0]    _zz_889;
  wire       [0:0]    _zz_890;
  wire       [31:0]   _zz_891;
  wire       [31:0]   _zz_892;
  wire       [31:0]   _zz_893;
  wire       [0:0]    _zz_894;
  wire       [0:0]    _zz_895;
  wire       [31:0]   _zz_896;
  wire       [31:0]   _zz_897;
  wire       [31:0]   _zz_898;
  wire       [0:0]    _zz_899;
  wire       [0:0]    _zz_900;
  wire       [31:0]   _zz_901;
  wire       [31:0]   _zz_902;
  wire       [31:0]   _zz_903;
  wire       [0:0]    _zz_904;
  wire       [0:0]    _zz_905;
  wire       [31:0]   _zz_906;
  wire       [31:0]   _zz_907;
  wire       [31:0]   _zz_908;
  wire       [0:0]    _zz_909;
  wire       [0:0]    _zz_910;
  wire       [31:0]   _zz_911;
  wire       [31:0]   _zz_912;
  wire       [31:0]   _zz_913;
  wire       [0:0]    _zz_914;
  wire       [0:0]    _zz_915;
  wire       [31:0]   _zz_916;
  wire       [31:0]   _zz_917;
  wire       [31:0]   _zz_918;
  wire       [0:0]    _zz_919;
  wire       [0:0]    _zz_920;
  wire       [31:0]   _zz_921;
  wire       [31:0]   _zz_922;
  wire       [31:0]   _zz_923;
  wire       [0:0]    _zz_924;
  wire       [0:0]    _zz_925;
  wire       [31:0]   _zz_926;
  wire       [31:0]   _zz_927;
  wire       [31:0]   _zz_928;
  wire       [0:0]    _zz_929;
  wire       [0:0]    _zz_930;
  wire       [31:0]   _zz_931;
  wire       [31:0]   _zz_932;
  wire       [31:0]   _zz_933;
  wire       [0:0]    _zz_934;
  wire       [0:0]    _zz_935;
  wire       [31:0]   _zz_936;
  wire       [31:0]   _zz_937;
  wire       [31:0]   _zz_938;
  wire       [0:0]    _zz_939;
  wire       [0:0]    _zz_940;
  wire       [31:0]   _zz_941;
  wire       [31:0]   _zz_942;
  wire       [31:0]   _zz_943;
  wire       [0:0]    _zz_944;
  wire       [0:0]    _zz_945;
  wire       [31:0]   _zz_946;
  wire       [31:0]   _zz_947;
  wire       [31:0]   _zz_948;
  wire       [0:0]    _zz_949;
  wire       [0:0]    _zz_950;
  wire       [31:0]   _zz_951;
  wire       [31:0]   _zz_952;
  wire       [31:0]   _zz_953;
  wire       [0:0]    _zz_954;
  wire       [0:0]    _zz_955;
  wire       [31:0]   _zz_956;
  wire       [31:0]   _zz_957;
  wire       [31:0]   _zz_958;
  wire       [0:0]    _zz_959;
  wire       [0:0]    _zz_960;
  wire       [31:0]   _zz_961;
  wire       [31:0]   _zz_962;
  wire       [31:0]   _zz_963;
  wire       [0:0]    _zz_964;
  wire       [0:0]    _zz_965;
  wire       [31:0]   _zz_966;
  wire       [31:0]   _zz_967;
  wire       [31:0]   _zz_968;
  wire       [0:0]    _zz_969;
  wire       [0:0]    _zz_970;
  wire       [31:0]   _zz_971;
  wire       [31:0]   _zz_972;
  wire       [31:0]   _zz_973;
  wire       [0:0]    _zz_974;
  wire       [0:0]    _zz_975;
  wire       [31:0]   _zz_976;
  wire       [31:0]   _zz_977;
  wire       [31:0]   _zz_978;
  wire       [0:0]    _zz_979;
  wire       [0:0]    _zz_980;
  wire       [31:0]   _zz_981;
  wire       [31:0]   _zz_982;
  wire       [31:0]   _zz_983;
  wire       [0:0]    _zz_984;
  wire       [0:0]    _zz_985;
  wire       [31:0]   _zz_986;
  wire       [31:0]   _zz_987;
  wire       [31:0]   _zz_988;
  wire       [0:0]    _zz_989;
  wire       [0:0]    _zz_990;
  wire       [31:0]   _zz_991;
  wire       [31:0]   _zz_992;
  wire       [31:0]   _zz_993;
  wire       [0:0]    _zz_994;
  wire       [0:0]    _zz_995;
  wire       [31:0]   _zz_996;
  wire       [31:0]   _zz_997;
  wire       [31:0]   _zz_998;
  wire       [0:0]    _zz_999;
  wire       [0:0]    _zz_1000;
  wire       [31:0]   _zz_1001;
  wire       [31:0]   _zz_1002;
  wire       [31:0]   _zz_1003;
  wire       [0:0]    _zz_1004;
  wire       [0:0]    _zz_1005;
  wire       [31:0]   _zz_1006;
  wire       [31:0]   _zz_1007;
  wire       [31:0]   _zz_1008;
  wire       [0:0]    _zz_1009;
  wire       [0:0]    _zz_1010;
  wire       [31:0]   _zz_1011;
  wire       [31:0]   _zz_1012;
  wire       [31:0]   _zz_1013;
  wire       [0:0]    _zz_1014;
  wire       [0:0]    _zz_1015;
  wire       [31:0]   _zz_1016;
  wire       [31:0]   _zz_1017;
  wire       [31:0]   _zz_1018;
  wire       [0:0]    _zz_1019;
  wire       [0:0]    _zz_1020;
  wire       [31:0]   _zz_1021;
  wire       [31:0]   _zz_1022;
  wire       [31:0]   _zz_1023;
  wire       [0:0]    _zz_1024;
  wire       [0:0]    _zz_1025;
  wire       [31:0]   _zz_1026;
  wire       [31:0]   _zz_1027;
  wire       [31:0]   _zz_1028;
  wire       [0:0]    _zz_1029;
  wire       [0:0]    _zz_1030;
  wire       [31:0]   _zz_1031;
  wire       [31:0]   _zz_1032;
  wire       [31:0]   _zz_1033;
  wire       [0:0]    _zz_1034;
  wire       [0:0]    _zz_1035;
  wire       [31:0]   _zz_1036;
  wire       [31:0]   _zz_1037;
  wire       [31:0]   _zz_1038;
  wire       [0:0]    _zz_1039;
  wire       [0:0]    _zz_1040;
  wire       [31:0]   _zz_1041;
  wire       [31:0]   _zz_1042;
  wire       [31:0]   _zz_1043;
  wire       [0:0]    _zz_1044;
  wire       [0:0]    _zz_1045;
  wire       [31:0]   _zz_1046;
  wire       [31:0]   _zz_1047;
  wire       [31:0]   _zz_1048;
  wire       [0:0]    _zz_1049;
  wire       [0:0]    _zz_1050;
  wire       [31:0]   _zz_1051;
  wire       [31:0]   _zz_1052;
  wire       [31:0]   _zz_1053;
  wire       [0:0]    _zz_1054;
  wire       [0:0]    _zz_1055;
  wire       [31:0]   _zz_1056;
  wire       [31:0]   _zz_1057;
  wire       [31:0]   _zz_1058;
  wire       [0:0]    _zz_1059;
  wire       [0:0]    _zz_1060;
  wire       [31:0]   _zz_1061;
  wire       [31:0]   _zz_1062;
  wire       [31:0]   _zz_1063;
  wire       [0:0]    _zz_1064;
  wire       [0:0]    _zz_1065;
  wire       [31:0]   _zz_1066;
  wire       [31:0]   _zz_1067;
  wire       [31:0]   _zz_1068;
  wire       [0:0]    _zz_1069;
  wire       [0:0]    _zz_1070;
  wire       [31:0]   _zz_1071;
  wire       [31:0]   _zz_1072;
  wire       [31:0]   _zz_1073;
  wire       [0:0]    _zz_1074;
  wire       [0:0]    _zz_1075;
  wire       [31:0]   _zz_1076;
  wire       [31:0]   _zz_1077;
  wire       [31:0]   _zz_1078;
  wire       [0:0]    _zz_1079;
  wire       [0:0]    _zz_1080;
  wire       [31:0]   _zz_1081;
  wire       [31:0]   _zz_1082;
  wire       [31:0]   _zz_1083;
  wire       [0:0]    _zz_1084;
  wire       [0:0]    _zz_1085;
  wire       [31:0]   _zz_1086;
  wire       [31:0]   _zz_1087;
  wire       [31:0]   _zz_1088;
  wire       [0:0]    _zz_1089;
  wire       [0:0]    _zz_1090;
  wire       [31:0]   _zz_1091;
  wire       [31:0]   _zz_1092;
  wire       [31:0]   _zz_1093;
  wire       [0:0]    _zz_1094;
  wire       [0:0]    _zz_1095;
  wire       [31:0]   _zz_1096;
  wire       [31:0]   _zz_1097;
  wire       [31:0]   _zz_1098;
  wire       [0:0]    _zz_1099;
  wire       [0:0]    _zz_1100;
  wire       [31:0]   _zz_1101;
  wire       [31:0]   _zz_1102;
  wire       [31:0]   _zz_1103;
  wire       [0:0]    _zz_1104;
  wire       [0:0]    _zz_1105;
  wire       [31:0]   _zz_1106;
  wire       [31:0]   _zz_1107;
  wire       [31:0]   _zz_1108;
  wire       [0:0]    _zz_1109;
  wire       [0:0]    _zz_1110;
  wire       [31:0]   _zz_1111;
  wire       [31:0]   _zz_1112;
  wire       [31:0]   _zz_1113;
  wire       [0:0]    _zz_1114;
  wire       [0:0]    _zz_1115;
  wire       [31:0]   _zz_1116;
  wire       [31:0]   _zz_1117;
  wire       [31:0]   _zz_1118;
  wire       [0:0]    _zz_1119;
  wire       [0:0]    _zz_1120;
  wire       [31:0]   _zz_1121;
  wire       [31:0]   _zz_1122;
  wire       [31:0]   _zz_1123;
  wire       [0:0]    _zz_1124;
  wire       [0:0]    _zz_1125;
  wire       [31:0]   _zz_1126;
  wire       [31:0]   _zz_1127;
  wire       [31:0]   _zz_1128;
  wire       [0:0]    _zz_1129;
  wire       [0:0]    _zz_1130;
  wire       [31:0]   _zz_1131;
  wire       [31:0]   _zz_1132;
  wire       [31:0]   _zz_1133;
  wire       [0:0]    _zz_1134;
  wire       [0:0]    _zz_1135;
  wire       [31:0]   _zz_1136;
  wire       [31:0]   _zz_1137;
  wire       [31:0]   _zz_1138;
  wire       [0:0]    _zz_1139;
  wire       [0:0]    _zz_1140;
  wire       [31:0]   _zz_1141;
  wire       [31:0]   _zz_1142;
  wire       [31:0]   _zz_1143;
  wire       [0:0]    _zz_1144;
  wire       [0:0]    _zz_1145;
  wire       [31:0]   _zz_1146;
  wire       [31:0]   _zz_1147;
  wire       [31:0]   _zz_1148;
  wire       [0:0]    _zz_1149;
  wire       [0:0]    _zz_1150;
  wire       [31:0]   _zz_1151;
  wire       [31:0]   _zz_1152;
  wire       [31:0]   _zz_1153;
  wire       [0:0]    _zz_1154;
  wire       [0:0]    _zz_1155;
  wire       [31:0]   _zz_1156;
  wire       [31:0]   _zz_1157;
  wire       [31:0]   _zz_1158;
  wire       [0:0]    _zz_1159;
  wire       [0:0]    _zz_1160;
  wire       [31:0]   _zz_1161;
  wire       [31:0]   _zz_1162;
  wire       [31:0]   _zz_1163;
  wire       [0:0]    _zz_1164;
  wire       [0:0]    _zz_1165;
  wire       [31:0]   _zz_1166;
  wire       [31:0]   _zz_1167;
  wire       [31:0]   _zz_1168;
  wire       [0:0]    _zz_1169;
  wire       [0:0]    _zz_1170;
  wire       [31:0]   _zz_1171;
  wire       [31:0]   _zz_1172;
  wire       [31:0]   _zz_1173;
  wire       [0:0]    _zz_1174;
  wire       [0:0]    _zz_1175;
  wire       [31:0]   _zz_1176;
  wire       [31:0]   _zz_1177;
  wire       [31:0]   _zz_1178;
  wire       [0:0]    _zz_1179;
  wire       [0:0]    _zz_1180;
  wire       [31:0]   _zz_1181;
  wire       [31:0]   _zz_1182;
  wire       [31:0]   _zz_1183;
  wire       [0:0]    _zz_1184;
  wire       [0:0]    _zz_1185;
  wire       [31:0]   _zz_1186;
  wire       [31:0]   _zz_1187;
  wire       [31:0]   _zz_1188;
  wire       [0:0]    _zz_1189;
  wire       [0:0]    _zz_1190;
  wire       [31:0]   _zz_1191;
  wire       [31:0]   _zz_1192;
  wire       [31:0]   _zz_1193;
  wire       [0:0]    _zz_1194;
  wire       [0:0]    _zz_1195;
  wire       [31:0]   _zz_1196;
  wire       [31:0]   _zz_1197;
  wire       [31:0]   _zz_1198;
  wire       [0:0]    _zz_1199;
  wire       [0:0]    _zz_1200;
  wire       [31:0]   _zz_1201;
  wire       [31:0]   _zz_1202;
  wire       [31:0]   _zz_1203;
  wire       [0:0]    _zz_1204;
  wire       [0:0]    _zz_1205;
  wire       [31:0]   _zz_1206;
  wire       [31:0]   _zz_1207;
  wire       [31:0]   _zz_1208;
  wire       [0:0]    _zz_1209;
  wire       [0:0]    _zz_1210;
  wire       [31:0]   _zz_1211;
  wire       [31:0]   _zz_1212;
  wire       [31:0]   _zz_1213;
  wire       [0:0]    _zz_1214;
  wire       [0:0]    _zz_1215;
  wire       [31:0]   _zz_1216;
  wire       [31:0]   _zz_1217;
  wire       [31:0]   _zz_1218;
  wire       [0:0]    _zz_1219;
  wire       [0:0]    _zz_1220;
  wire       [31:0]   _zz_1221;
  wire       [31:0]   _zz_1222;
  wire       [31:0]   _zz_1223;
  wire       [0:0]    _zz_1224;
  wire       [0:0]    _zz_1225;
  wire       [31:0]   _zz_1226;
  wire       [31:0]   _zz_1227;
  wire       [31:0]   _zz_1228;
  wire       [0:0]    _zz_1229;
  wire       [0:0]    _zz_1230;
  wire       [31:0]   _zz_1231;
  wire       [31:0]   _zz_1232;
  wire       [31:0]   _zz_1233;
  wire       [0:0]    _zz_1234;
  wire       [0:0]    _zz_1235;
  wire       [31:0]   _zz_1236;
  wire       [31:0]   _zz_1237;
  wire       [31:0]   _zz_1238;
  wire       [0:0]    _zz_1239;
  wire       [0:0]    _zz_1240;
  wire       [31:0]   _zz_1241;
  wire       [31:0]   _zz_1242;
  wire       [31:0]   _zz_1243;
  wire       [0:0]    _zz_1244;
  wire       [0:0]    _zz_1245;
  wire       [31:0]   _zz_1246;
  wire       [31:0]   _zz_1247;
  wire       [31:0]   _zz_1248;
  wire       [0:0]    _zz_1249;
  wire       [0:0]    _zz_1250;
  wire       [31:0]   _zz_1251;
  wire       [31:0]   _zz_1252;
  wire       [31:0]   _zz_1253;
  wire       [0:0]    _zz_1254;
  wire       [0:0]    _zz_1255;
  wire       [31:0]   _zz_1256;
  wire       [31:0]   _zz_1257;
  wire       [31:0]   _zz_1258;
  wire       [0:0]    _zz_1259;
  wire       [0:0]    _zz_1260;
  wire       [31:0]   _zz_1261;
  wire       [31:0]   _zz_1262;
  wire       [31:0]   _zz_1263;
  wire       [0:0]    _zz_1264;
  wire       [0:0]    _zz_1265;
  wire       [31:0]   _zz_1266;
  wire       [31:0]   _zz_1267;
  wire       [31:0]   _zz_1268;
  wire       [0:0]    _zz_1269;
  wire       [0:0]    _zz_1270;
  wire       [31:0]   _zz_1271;
  wire       [31:0]   _zz_1272;
  wire       [31:0]   _zz_1273;
  wire       [0:0]    _zz_1274;
  wire       [0:0]    _zz_1275;
  wire       [31:0]   _zz_1276;
  wire       [31:0]   _zz_1277;
  wire       [31:0]   _zz_1278;
  wire       [0:0]    _zz_1279;
  wire       [0:0]    _zz_1280;
  wire       [31:0]   _zz_1281;
  wire       [31:0]   _zz_1282;
  wire       [31:0]   _zz_1283;
  wire       [0:0]    _zz_1284;
  wire       [0:0]    _zz_1285;
  wire       [31:0]   _zz_1286;
  wire       [31:0]   _zz_1287;
  wire       [31:0]   _zz_1288;
  wire       [0:0]    _zz_1289;
  wire       [0:0]    _zz_1290;
  wire       [31:0]   _zz_1291;
  wire       [31:0]   _zz_1292;
  wire       [31:0]   _zz_1293;
  wire       [0:0]    _zz_1294;
  wire       [0:0]    _zz_1295;
  wire       [31:0]   _zz_1296;
  wire       [31:0]   _zz_1297;
  wire       [31:0]   _zz_1298;
  wire       [0:0]    _zz_1299;
  wire       [0:0]    _zz_1300;
  wire       [31:0]   _zz_1301;
  wire       [31:0]   _zz_1302;
  wire       [31:0]   _zz_1303;
  wire       [0:0]    _zz_1304;
  wire       [0:0]    _zz_1305;
  wire       [31:0]   _zz_1306;
  wire       [31:0]   _zz_1307;
  wire       [31:0]   _zz_1308;
  wire       [0:0]    _zz_1309;
  wire       [0:0]    _zz_1310;
  wire       [31:0]   _zz_1311;
  wire       [31:0]   _zz_1312;
  wire       [31:0]   _zz_1313;
  wire       [0:0]    _zz_1314;
  wire       [0:0]    _zz_1315;
  wire       [31:0]   _zz_1316;
  wire       [31:0]   _zz_1317;
  wire       [31:0]   _zz_1318;
  wire       [0:0]    _zz_1319;
  wire       [0:0]    _zz_1320;
  wire       [31:0]   _zz_1321;
  wire       [31:0]   _zz_1322;
  wire       [31:0]   _zz_1323;
  wire       [0:0]    _zz_1324;
  wire       [0:0]    _zz_1325;
  wire       [31:0]   _zz_1326;
  wire       [31:0]   _zz_1327;
  wire       [31:0]   _zz_1328;
  wire       [0:0]    _zz_1329;
  wire       [0:0]    _zz_1330;
  wire       [31:0]   _zz_1331;
  wire       [31:0]   _zz_1332;
  wire       [31:0]   _zz_1333;
  wire       [0:0]    _zz_1334;
  wire       [0:0]    _zz_1335;
  wire       [31:0]   _zz_1336;
  wire       [31:0]   _zz_1337;
  wire       [31:0]   _zz_1338;
  wire       [0:0]    _zz_1339;
  wire       [0:0]    _zz_1340;
  wire       [31:0]   _zz_1341;
  wire       [31:0]   _zz_1342;
  wire       [31:0]   _zz_1343;
  wire       [0:0]    _zz_1344;
  wire       [0:0]    _zz_1345;
  wire       [31:0]   _zz_1346;
  wire       [31:0]   _zz_1347;
  wire       [31:0]   _zz_1348;
  wire       [0:0]    _zz_1349;
  wire       [0:0]    _zz_1350;
  wire       [31:0]   _zz_1351;
  wire       [31:0]   _zz_1352;
  wire       [31:0]   _zz_1353;
  wire       [0:0]    _zz_1354;
  wire       [0:0]    _zz_1355;
  wire       [31:0]   _zz_1356;
  wire       [31:0]   _zz_1357;
  wire       [31:0]   _zz_1358;
  wire       [0:0]    _zz_1359;
  wire       [0:0]    _zz_1360;
  wire       [31:0]   _zz_1361;
  wire       [31:0]   _zz_1362;
  wire       [31:0]   _zz_1363;
  wire       [0:0]    _zz_1364;
  wire       [0:0]    _zz_1365;
  wire       [31:0]   _zz_1366;
  wire       [31:0]   _zz_1367;
  wire       [31:0]   _zz_1368;
  wire       [0:0]    _zz_1369;
  wire       [0:0]    _zz_1370;
  wire       [31:0]   _zz_1371;
  wire       [31:0]   _zz_1372;
  wire       [31:0]   _zz_1373;
  wire       [0:0]    _zz_1374;
  wire       [0:0]    _zz_1375;
  wire       [31:0]   _zz_1376;
  wire       [31:0]   _zz_1377;
  wire       [31:0]   _zz_1378;
  wire       [0:0]    _zz_1379;
  wire       [0:0]    _zz_1380;
  wire       [31:0]   _zz_1381;
  wire       [31:0]   _zz_1382;
  wire       [31:0]   _zz_1383;
  wire       [0:0]    _zz_1384;
  wire       [0:0]    _zz_1385;
  wire       [31:0]   _zz_1386;
  wire       [31:0]   _zz_1387;
  wire       [31:0]   _zz_1388;
  wire       [0:0]    _zz_1389;
  wire       [0:0]    _zz_1390;
  wire       [31:0]   _zz_1391;
  wire       [31:0]   _zz_1392;
  wire       [31:0]   _zz_1393;
  wire       [0:0]    _zz_1394;
  wire       [0:0]    _zz_1395;
  wire       [31:0]   _zz_1396;
  wire       [31:0]   _zz_1397;
  wire       [31:0]   _zz_1398;
  wire       [0:0]    _zz_1399;
  wire       [0:0]    _zz_1400;
  wire       [31:0]   _zz_1401;
  wire       [31:0]   _zz_1402;
  wire       [31:0]   _zz_1403;
  wire       [0:0]    _zz_1404;
  wire       [0:0]    _zz_1405;
  wire       [31:0]   _zz_1406;
  wire       [31:0]   _zz_1407;
  wire       [31:0]   _zz_1408;
  wire       [0:0]    _zz_1409;
  wire       [0:0]    _zz_1410;
  wire       [31:0]   _zz_1411;
  wire       [31:0]   _zz_1412;
  wire       [31:0]   _zz_1413;
  wire       [0:0]    _zz_1414;
  wire       [0:0]    _zz_1415;
  wire       [31:0]   _zz_1416;
  wire       [31:0]   _zz_1417;
  wire       [31:0]   _zz_1418;
  wire       [0:0]    _zz_1419;
  wire       [0:0]    _zz_1420;
  wire       [31:0]   _zz_1421;
  wire       [31:0]   _zz_1422;
  wire       [31:0]   _zz_1423;
  wire       [0:0]    _zz_1424;
  wire       [0:0]    _zz_1425;
  wire       [31:0]   _zz_1426;
  wire       [31:0]   _zz_1427;
  wire       [31:0]   _zz_1428;
  wire       [0:0]    _zz_1429;
  wire       [0:0]    _zz_1430;
  wire       [31:0]   _zz_1431;
  wire       [31:0]   _zz_1432;
  wire       [31:0]   _zz_1433;
  wire       [0:0]    _zz_1434;
  wire       [0:0]    _zz_1435;
  wire       [31:0]   _zz_1436;
  wire       [31:0]   _zz_1437;
  wire       [31:0]   _zz_1438;
  wire       [0:0]    _zz_1439;
  wire       [0:0]    _zz_1440;
  wire       [31:0]   _zz_1441;
  wire       [31:0]   _zz_1442;
  wire       [31:0]   _zz_1443;
  wire       [0:0]    _zz_1444;
  wire       [0:0]    _zz_1445;
  wire       [31:0]   _zz_1446;
  wire       [31:0]   _zz_1447;
  wire       [31:0]   _zz_1448;
  wire       [0:0]    _zz_1449;
  wire       [0:0]    _zz_1450;
  wire       [31:0]   _zz_1451;
  wire       [31:0]   _zz_1452;
  wire       [31:0]   _zz_1453;
  wire       [0:0]    _zz_1454;
  wire       [0:0]    _zz_1455;
  wire       [31:0]   _zz_1456;
  wire       [31:0]   _zz_1457;
  wire       [31:0]   _zz_1458;
  wire       [0:0]    _zz_1459;
  wire       [0:0]    _zz_1460;
  wire       [31:0]   _zz_1461;
  wire       [31:0]   _zz_1462;
  wire       [31:0]   _zz_1463;
  wire       [0:0]    _zz_1464;
  wire       [0:0]    _zz_1465;
  wire       [31:0]   _zz_1466;
  wire       [31:0]   _zz_1467;
  wire       [31:0]   _zz_1468;
  wire       [0:0]    _zz_1469;
  wire       [0:0]    _zz_1470;
  wire       [31:0]   _zz_1471;
  wire       [31:0]   _zz_1472;
  wire       [31:0]   _zz_1473;
  wire       [0:0]    _zz_1474;
  wire       [0:0]    _zz_1475;
  wire       [31:0]   _zz_1476;
  wire       [31:0]   _zz_1477;
  wire       [31:0]   _zz_1478;
  wire       [0:0]    _zz_1479;
  wire       [0:0]    _zz_1480;
  wire       [31:0]   _zz_1481;
  wire       [31:0]   _zz_1482;
  wire       [31:0]   _zz_1483;
  wire       [0:0]    _zz_1484;
  wire       [0:0]    _zz_1485;
  wire       [31:0]   _zz_1486;
  wire       [31:0]   _zz_1487;
  wire       [31:0]   _zz_1488;
  wire       [0:0]    _zz_1489;
  wire       [0:0]    _zz_1490;
  wire       [31:0]   _zz_1491;
  wire       [31:0]   _zz_1492;
  wire       [31:0]   _zz_1493;
  wire       [0:0]    _zz_1494;
  wire       [0:0]    _zz_1495;
  wire       [31:0]   _zz_1496;
  wire       [31:0]   _zz_1497;
  wire       [31:0]   _zz_1498;
  wire       [0:0]    _zz_1499;
  wire       [0:0]    _zz_1500;
  wire       [31:0]   _zz_1501;
  wire       [31:0]   _zz_1502;
  wire       [31:0]   _zz_1503;
  wire       [0:0]    _zz_1504;
  wire       [0:0]    _zz_1505;
  wire       [31:0]   _zz_1506;
  wire       [31:0]   _zz_1507;
  wire       [31:0]   _zz_1508;
  wire       [0:0]    _zz_1509;
  wire       [0:0]    _zz_1510;
  wire       [31:0]   _zz_1511;
  wire       [31:0]   _zz_1512;
  wire       [31:0]   _zz_1513;
  wire       [0:0]    _zz_1514;
  wire       [0:0]    _zz_1515;
  wire       [31:0]   _zz_1516;
  wire       [31:0]   _zz_1517;
  wire       [31:0]   _zz_1518;
  wire       [0:0]    _zz_1519;
  wire       [0:0]    _zz_1520;
  wire       [31:0]   _zz_1521;
  wire       [31:0]   _zz_1522;
  wire       [31:0]   _zz_1523;
  wire       [0:0]    _zz_1524;
  wire       [0:0]    _zz_1525;
  wire       [31:0]   _zz_1526;
  wire       [31:0]   _zz_1527;
  wire       [31:0]   _zz_1528;
  wire       [0:0]    _zz_1529;
  wire       [0:0]    _zz_1530;
  wire       [31:0]   _zz_1531;
  wire       [31:0]   _zz_1532;
  wire       [31:0]   _zz_1533;
  wire       [0:0]    _zz_1534;
  wire       [0:0]    _zz_1535;
  wire       [31:0]   _zz_1536;
  wire       [31:0]   _zz_1537;
  wire       [31:0]   _zz_1538;
  wire       [0:0]    _zz_1539;
  wire       [0:0]    _zz_1540;
  wire       [31:0]   _zz_1541;
  wire       [31:0]   _zz_1542;
  wire       [31:0]   _zz_1543;
  wire       [0:0]    _zz_1544;
  wire       [0:0]    _zz_1545;
  wire       [31:0]   _zz_1546;
  wire       [31:0]   _zz_1547;
  wire       [31:0]   _zz_1548;
  wire       [0:0]    _zz_1549;
  wire       [0:0]    _zz_1550;
  wire       [31:0]   _zz_1551;
  wire       [31:0]   _zz_1552;
  wire       [31:0]   _zz_1553;
  wire       [0:0]    _zz_1554;
  wire       [0:0]    _zz_1555;
  wire       [31:0]   _zz_1556;
  wire       [31:0]   _zz_1557;
  wire       [31:0]   _zz_1558;
  wire       [0:0]    _zz_1559;
  wire       [0:0]    _zz_1560;
  wire       [31:0]   _zz_1561;
  wire       [31:0]   _zz_1562;
  wire       [31:0]   _zz_1563;
  wire       [0:0]    _zz_1564;
  wire       [0:0]    _zz_1565;
  wire       [31:0]   _zz_1566;
  wire       [31:0]   _zz_1567;
  wire       [31:0]   _zz_1568;
  wire       [0:0]    _zz_1569;
  wire       [0:0]    _zz_1570;
  wire       [31:0]   _zz_1571;
  wire       [31:0]   _zz_1572;
  wire       [31:0]   _zz_1573;
  wire       [0:0]    _zz_1574;
  wire       [0:0]    _zz_1575;
  wire       [31:0]   _zz_1576;
  wire       [31:0]   _zz_1577;
  wire       [31:0]   _zz_1578;
  wire       [0:0]    _zz_1579;
  wire       [0:0]    _zz_1580;
  wire       [31:0]   _zz_1581;
  wire       [31:0]   _zz_1582;
  wire       [31:0]   _zz_1583;
  wire       [0:0]    _zz_1584;
  wire       [0:0]    _zz_1585;
  wire       [31:0]   _zz_1586;
  wire       [31:0]   _zz_1587;
  wire       [31:0]   _zz_1588;
  wire       [0:0]    _zz_1589;
  wire       [0:0]    _zz_1590;
  wire       [31:0]   _zz_1591;
  wire       [31:0]   _zz_1592;
  wire       [31:0]   _zz_1593;
  wire       [0:0]    _zz_1594;
  wire       [0:0]    _zz_1595;
  wire       [31:0]   _zz_1596;
  wire       [31:0]   _zz_1597;
  wire       [31:0]   _zz_1598;
  wire       [0:0]    _zz_1599;
  wire       [0:0]    _zz_1600;
  wire       [31:0]   _zz_1601;
  wire       [31:0]   _zz_1602;
  wire       [31:0]   _zz_1603;
  wire       [0:0]    _zz_1604;
  wire       [0:0]    _zz_1605;
  wire       [31:0]   _zz_1606;
  wire       [31:0]   _zz_1607;
  wire       [31:0]   _zz_1608;
  wire       [0:0]    _zz_1609;
  wire       [0:0]    _zz_1610;
  wire       [31:0]   _zz_1611;
  wire       [31:0]   _zz_1612;
  wire       [31:0]   _zz_1613;
  wire       [0:0]    _zz_1614;
  wire       [0:0]    _zz_1615;
  wire       [31:0]   _zz_1616;
  wire       [31:0]   _zz_1617;
  wire       [31:0]   _zz_1618;
  wire       [0:0]    _zz_1619;
  wire       [0:0]    _zz_1620;
  wire       [31:0]   _zz_1621;
  wire       [31:0]   _zz_1622;
  wire       [31:0]   _zz_1623;
  wire       [0:0]    _zz_1624;
  wire       [0:0]    _zz_1625;
  wire       [31:0]   _zz_1626;
  wire       [31:0]   _zz_1627;
  wire       [31:0]   _zz_1628;
  wire       [0:0]    _zz_1629;
  wire       [0:0]    _zz_1630;
  wire       [31:0]   _zz_1631;
  wire       [31:0]   _zz_1632;
  wire       [31:0]   _zz_1633;
  wire       [0:0]    _zz_1634;
  wire       [0:0]    _zz_1635;
  wire       [31:0]   _zz_1636;
  wire       [31:0]   _zz_1637;
  wire       [31:0]   _zz_1638;
  wire       [0:0]    _zz_1639;
  wire       [0:0]    _zz_1640;
  wire       [31:0]   _zz_1641;
  wire       [31:0]   _zz_1642;
  wire       [31:0]   _zz_1643;
  wire       [0:0]    _zz_1644;
  wire       [0:0]    _zz_1645;
  wire       [31:0]   _zz_1646;
  wire       [31:0]   _zz_1647;
  wire       [31:0]   _zz_1648;
  wire       [0:0]    _zz_1649;
  wire       [0:0]    _zz_1650;
  wire       [31:0]   _zz_1651;
  wire       [31:0]   _zz_1652;
  wire       [31:0]   _zz_1653;
  wire       [0:0]    _zz_1654;
  wire       [0:0]    _zz_1655;
  wire       [31:0]   _zz_1656;
  wire       [31:0]   _zz_1657;
  wire       [31:0]   _zz_1658;
  wire       [0:0]    _zz_1659;
  wire       [0:0]    _zz_1660;
  wire       [31:0]   _zz_1661;
  wire       [31:0]   _zz_1662;
  wire       [31:0]   _zz_1663;
  wire       [0:0]    _zz_1664;
  wire       [0:0]    _zz_1665;
  wire       [31:0]   _zz_1666;
  wire       [31:0]   _zz_1667;
  wire       [31:0]   _zz_1668;
  wire       [0:0]    _zz_1669;
  wire       [0:0]    _zz_1670;
  wire       [31:0]   _zz_1671;
  wire       [31:0]   _zz_1672;
  wire       [31:0]   _zz_1673;
  wire       [0:0]    _zz_1674;
  wire       [0:0]    _zz_1675;
  wire       [31:0]   _zz_1676;
  wire       [31:0]   _zz_1677;
  wire       [31:0]   _zz_1678;
  wire       [0:0]    _zz_1679;
  wire       [0:0]    _zz_1680;
  wire       [31:0]   _zz_1681;
  wire       [31:0]   _zz_1682;
  wire       [31:0]   _zz_1683;
  wire       [0:0]    _zz_1684;
  wire       [0:0]    _zz_1685;
  wire       [31:0]   _zz_1686;
  wire       [31:0]   _zz_1687;
  wire       [31:0]   _zz_1688;
  wire       [0:0]    _zz_1689;
  wire       [0:0]    _zz_1690;
  wire       [31:0]   _zz_1691;
  wire       [31:0]   _zz_1692;
  wire       [31:0]   _zz_1693;
  wire       [0:0]    _zz_1694;
  wire       [0:0]    _zz_1695;
  wire       [31:0]   _zz_1696;
  wire       [31:0]   _zz_1697;
  wire       [31:0]   _zz_1698;
  wire       [0:0]    _zz_1699;
  wire       [0:0]    _zz_1700;
  wire       [31:0]   _zz_1701;
  wire       [31:0]   _zz_1702;
  wire       [31:0]   _zz_1703;
  wire       [0:0]    _zz_1704;
  wire       [0:0]    _zz_1705;
  wire       [31:0]   _zz_1706;
  wire       [31:0]   _zz_1707;
  wire       [31:0]   _zz_1708;
  wire       [0:0]    _zz_1709;
  wire       [0:0]    _zz_1710;
  wire       [31:0]   _zz_1711;
  wire       [31:0]   _zz_1712;
  wire       [31:0]   _zz_1713;
  wire       [0:0]    _zz_1714;
  wire       [0:0]    _zz_1715;
  wire       [31:0]   _zz_1716;
  wire       [31:0]   _zz_1717;
  wire       [31:0]   _zz_1718;
  wire       [0:0]    _zz_1719;
  wire       [0:0]    _zz_1720;
  wire       [31:0]   _zz_1721;
  wire       [31:0]   _zz_1722;
  wire       [31:0]   _zz_1723;
  wire       [0:0]    _zz_1724;
  wire       [0:0]    _zz_1725;
  wire       [31:0]   _zz_1726;
  wire       [31:0]   _zz_1727;
  wire       [31:0]   _zz_1728;
  wire       [0:0]    _zz_1729;
  wire       [0:0]    _zz_1730;
  wire       [31:0]   _zz_1731;
  wire       [31:0]   _zz_1732;
  wire       [31:0]   _zz_1733;
  wire       [0:0]    _zz_1734;
  wire       [0:0]    _zz_1735;
  wire       [31:0]   _zz_1736;
  wire       [31:0]   _zz_1737;
  wire       [31:0]   _zz_1738;
  wire       [0:0]    _zz_1739;
  wire       [0:0]    _zz_1740;
  wire       [31:0]   _zz_1741;
  wire       [31:0]   _zz_1742;
  wire       [31:0]   _zz_1743;
  wire       [0:0]    _zz_1744;
  wire       [0:0]    _zz_1745;
  wire       [31:0]   _zz_1746;
  wire       [31:0]   _zz_1747;
  wire       [31:0]   _zz_1748;
  wire       [0:0]    _zz_1749;
  wire       [0:0]    _zz_1750;
  wire       [31:0]   _zz_1751;
  wire       [31:0]   _zz_1752;
  wire       [31:0]   _zz_1753;
  wire       [0:0]    _zz_1754;
  wire       [0:0]    _zz_1755;
  wire       [31:0]   _zz_1756;
  wire       [31:0]   _zz_1757;
  wire       [31:0]   _zz_1758;
  wire       [0:0]    _zz_1759;
  wire       [0:0]    _zz_1760;
  wire       [31:0]   _zz_1761;
  wire       [31:0]   _zz_1762;
  wire       [31:0]   _zz_1763;
  wire       [0:0]    _zz_1764;
  wire       [0:0]    _zz_1765;
  wire       [31:0]   _zz_1766;
  wire       [31:0]   _zz_1767;
  wire       [31:0]   _zz_1768;
  wire       [0:0]    _zz_1769;
  wire       [0:0]    _zz_1770;
  wire       [31:0]   _zz_1771;
  wire       [31:0]   _zz_1772;
  wire       [31:0]   _zz_1773;
  wire       [0:0]    _zz_1774;
  wire       [0:0]    _zz_1775;
  wire       [31:0]   _zz_1776;
  wire       [31:0]   _zz_1777;
  wire       [31:0]   _zz_1778;
  wire       [0:0]    _zz_1779;
  wire       [0:0]    _zz_1780;
  wire       [31:0]   _zz_1781;
  wire       [31:0]   _zz_1782;
  wire       [31:0]   _zz_1783;
  wire       [0:0]    _zz_1784;
  wire       [0:0]    _zz_1785;
  wire       [31:0]   _zz_1786;
  wire       [31:0]   _zz_1787;
  wire       [31:0]   _zz_1788;
  wire       [0:0]    _zz_1789;
  wire       [0:0]    _zz_1790;
  wire       [31:0]   _zz_1791;
  wire       [31:0]   _zz_1792;
  wire       [31:0]   _zz_1793;
  wire       [0:0]    _zz_1794;
  wire       [0:0]    _zz_1795;
  wire       [31:0]   _zz_1796;
  wire       [31:0]   _zz_1797;
  wire       [31:0]   _zz_1798;
  wire       [0:0]    _zz_1799;
  wire       [0:0]    _zz_1800;
  wire       [31:0]   _zz_1801;
  wire       [31:0]   _zz_1802;
  wire       [31:0]   _zz_1803;
  wire       [0:0]    _zz_1804;
  wire       [0:0]    _zz_1805;
  wire       [31:0]   _zz_1806;
  wire       [31:0]   _zz_1807;
  wire       [31:0]   _zz_1808;
  wire       [0:0]    _zz_1809;
  wire       [0:0]    _zz_1810;
  wire       [31:0]   _zz_1811;
  wire       [31:0]   _zz_1812;
  wire       [31:0]   _zz_1813;
  wire       [0:0]    _zz_1814;
  wire       [0:0]    _zz_1815;
  wire       [31:0]   _zz_1816;
  wire       [31:0]   _zz_1817;
  wire       [31:0]   _zz_1818;
  wire       [0:0]    _zz_1819;
  wire       [0:0]    _zz_1820;
  wire       [31:0]   _zz_1821;
  wire       [31:0]   _zz_1822;
  wire       [31:0]   _zz_1823;
  wire       [0:0]    _zz_1824;
  wire       [0:0]    _zz_1825;
  wire       [31:0]   _zz_1826;
  wire       [31:0]   _zz_1827;
  wire       [31:0]   _zz_1828;
  wire       [0:0]    _zz_1829;
  wire       [0:0]    _zz_1830;
  wire       [31:0]   _zz_1831;
  wire       [31:0]   _zz_1832;
  wire       [31:0]   _zz_1833;
  wire       [0:0]    _zz_1834;
  wire       [0:0]    _zz_1835;
  wire       [31:0]   _zz_1836;
  wire       [31:0]   _zz_1837;
  wire       [31:0]   _zz_1838;
  wire       [0:0]    _zz_1839;
  wire       [0:0]    _zz_1840;
  wire       [31:0]   _zz_1841;
  wire       [31:0]   _zz_1842;
  wire       [31:0]   _zz_1843;
  wire       [0:0]    _zz_1844;
  wire       [0:0]    _zz_1845;
  wire       [31:0]   _zz_1846;
  wire       [31:0]   _zz_1847;
  wire       [31:0]   _zz_1848;
  wire       [0:0]    _zz_1849;
  wire       [0:0]    _zz_1850;
  wire       [31:0]   _zz_1851;
  wire       [31:0]   _zz_1852;
  wire       [31:0]   _zz_1853;
  wire       [0:0]    _zz_1854;
  wire       [0:0]    _zz_1855;
  wire       [31:0]   _zz_1856;
  wire       [31:0]   _zz_1857;
  wire       [31:0]   _zz_1858;
  wire       [0:0]    _zz_1859;
  wire       [0:0]    _zz_1860;
  wire       [31:0]   _zz_1861;
  wire       [31:0]   _zz_1862;
  wire       [31:0]   _zz_1863;
  wire       [0:0]    _zz_1864;
  wire       [0:0]    _zz_1865;
  wire       [31:0]   _zz_1866;
  wire       [31:0]   _zz_1867;
  wire       [31:0]   _zz_1868;
  wire       [0:0]    _zz_1869;
  wire       [0:0]    _zz_1870;
  wire       [31:0]   _zz_1871;
  wire       [31:0]   _zz_1872;
  wire       [31:0]   _zz_1873;
  wire       [0:0]    _zz_1874;
  wire       [0:0]    _zz_1875;
  wire       [31:0]   _zz_1876;
  wire       [31:0]   _zz_1877;
  wire       [31:0]   _zz_1878;
  wire       [0:0]    _zz_1879;
  wire       [0:0]    _zz_1880;
  wire       [31:0]   _zz_1881;
  wire       [31:0]   _zz_1882;
  wire       [31:0]   _zz_1883;
  wire       [0:0]    _zz_1884;
  wire       [0:0]    _zz_1885;
  wire       [31:0]   _zz_1886;
  wire       [31:0]   _zz_1887;
  wire       [31:0]   _zz_1888;
  wire       [0:0]    _zz_1889;
  wire       [0:0]    _zz_1890;
  wire       [31:0]   _zz_1891;
  wire       [31:0]   _zz_1892;
  wire       [31:0]   _zz_1893;
  wire       [0:0]    _zz_1894;
  wire       [0:0]    _zz_1895;
  wire       [31:0]   _zz_1896;
  wire       [31:0]   _zz_1897;
  wire       [31:0]   _zz_1898;
  wire       [0:0]    _zz_1899;
  wire       [0:0]    _zz_1900;
  wire       [31:0]   _zz_1901;
  wire       [31:0]   _zz_1902;
  wire       [31:0]   _zz_1903;
  wire       [0:0]    _zz_1904;
  wire       [0:0]    _zz_1905;
  wire       [31:0]   _zz_1906;
  wire       [31:0]   _zz_1907;
  wire       [31:0]   _zz_1908;
  wire       [0:0]    _zz_1909;
  wire       [0:0]    _zz_1910;
  wire       [31:0]   _zz_1911;
  wire       [31:0]   _zz_1912;
  wire       [31:0]   _zz_1913;
  wire       [0:0]    _zz_1914;
  wire       [0:0]    _zz_1915;
  wire       [31:0]   _zz_1916;
  wire       [31:0]   _zz_1917;
  wire       [31:0]   _zz_1918;
  wire       [0:0]    _zz_1919;
  wire       [0:0]    _zz_1920;
  wire       [31:0]   _zz_1921;
  wire       [31:0]   _zz_1922;
  wire       [31:0]   _zz_1923;
  wire       [0:0]    _zz_1924;
  wire       [0:0]    _zz_1925;
  wire       [31:0]   _zz_1926;
  wire       [31:0]   _zz_1927;
  wire       [31:0]   _zz_1928;
  wire       [0:0]    _zz_1929;
  wire       [0:0]    _zz_1930;
  wire       [31:0]   _zz_1931;
  wire       [31:0]   _zz_1932;
  wire       [31:0]   _zz_1933;
  wire       [0:0]    _zz_1934;
  wire       [0:0]    _zz_1935;
  wire       [31:0]   _zz_1936;
  wire       [31:0]   _zz_1937;
  wire       [31:0]   _zz_1938;
  wire       [0:0]    _zz_1939;
  wire       [0:0]    _zz_1940;
  wire       [31:0]   _zz_1941;
  wire       [31:0]   _zz_1942;
  wire       [31:0]   _zz_1943;
  wire       [0:0]    _zz_1944;
  wire       [0:0]    _zz_1945;
  wire       [31:0]   _zz_1946;
  wire       [31:0]   _zz_1947;
  wire       [31:0]   _zz_1948;
  wire       [0:0]    _zz_1949;
  wire       [0:0]    _zz_1950;
  wire       [31:0]   _zz_1951;
  wire       [31:0]   _zz_1952;
  wire       [31:0]   _zz_1953;
  wire       [0:0]    _zz_1954;
  wire       [0:0]    _zz_1955;
  wire       [31:0]   _zz_1956;
  wire       [31:0]   _zz_1957;
  wire       [31:0]   _zz_1958;
  wire       [0:0]    _zz_1959;
  wire       [0:0]    _zz_1960;
  wire       [31:0]   _zz_1961;
  wire       [31:0]   _zz_1962;
  wire       [31:0]   _zz_1963;
  wire       [0:0]    _zz_1964;
  wire       [0:0]    _zz_1965;
  wire       [31:0]   _zz_1966;
  wire       [31:0]   _zz_1967;
  wire       [31:0]   _zz_1968;
  wire       [0:0]    _zz_1969;
  wire       [0:0]    _zz_1970;
  wire       [31:0]   _zz_1971;
  wire       [31:0]   _zz_1972;
  wire       [31:0]   _zz_1973;
  wire       [0:0]    _zz_1974;
  wire       [0:0]    _zz_1975;
  wire       [31:0]   _zz_1976;
  wire       [31:0]   _zz_1977;
  wire       [31:0]   _zz_1978;
  wire       [0:0]    _zz_1979;
  wire       [0:0]    _zz_1980;
  wire       [31:0]   _zz_1981;
  wire       [31:0]   _zz_1982;
  wire       [31:0]   _zz_1983;
  wire       [0:0]    _zz_1984;
  wire       [0:0]    _zz_1985;
  wire       [31:0]   _zz_1986;
  wire       [31:0]   _zz_1987;
  wire       [31:0]   _zz_1988;
  wire       [0:0]    _zz_1989;
  wire       [0:0]    _zz_1990;
  wire       [31:0]   _zz_1991;
  wire       [31:0]   _zz_1992;
  wire       [31:0]   _zz_1993;
  wire       [0:0]    _zz_1994;
  wire       [0:0]    _zz_1995;
  wire       [31:0]   _zz_1996;
  wire       [31:0]   _zz_1997;
  wire       [31:0]   _zz_1998;
  wire       [0:0]    _zz_1999;
  wire       [0:0]    _zz_2000;
  wire       [31:0]   _zz_2001;
  wire       [31:0]   _zz_2002;
  wire       [31:0]   _zz_2003;
  wire       [0:0]    _zz_2004;
  wire       [0:0]    _zz_2005;
  wire       [31:0]   _zz_2006;
  wire       [31:0]   _zz_2007;
  wire       [31:0]   _zz_2008;
  wire       [0:0]    _zz_2009;
  wire       [0:0]    _zz_2010;
  wire       [31:0]   _zz_2011;
  wire       [31:0]   _zz_2012;
  wire       [31:0]   _zz_2013;
  wire       [0:0]    _zz_2014;
  wire       [0:0]    _zz_2015;
  wire       [31:0]   _zz_2016;
  wire       [31:0]   _zz_2017;
  wire       [31:0]   _zz_2018;
  wire       [0:0]    _zz_2019;
  wire       [0:0]    _zz_2020;
  wire       [31:0]   _zz_2021;
  wire       [31:0]   _zz_2022;
  wire       [31:0]   _zz_2023;
  wire       [0:0]    _zz_2024;
  wire       [0:0]    _zz_2025;
  wire       [31:0]   _zz_2026;
  wire       [31:0]   _zz_2027;
  wire       [31:0]   _zz_2028;
  wire       [0:0]    _zz_2029;
  wire       [0:0]    _zz_2030;
  wire       [31:0]   _zz_2031;
  wire       [31:0]   _zz_2032;
  wire       [31:0]   _zz_2033;
  wire       [0:0]    _zz_2034;
  wire       [0:0]    _zz_2035;
  wire       [31:0]   _zz_2036;
  wire       [31:0]   _zz_2037;
  wire       [31:0]   _zz_2038;
  wire       [0:0]    _zz_2039;
  wire       [0:0]    _zz_2040;
  wire       [31:0]   _zz_2041;
  wire       [31:0]   _zz_2042;
  wire       [31:0]   _zz_2043;
  wire       [0:0]    _zz_2044;
  wire       [0:0]    _zz_2045;
  wire       [31:0]   _zz_2046;
  wire       [31:0]   _zz_2047;
  wire       [31:0]   _zz_2048;
  wire       [0:0]    _zz_2049;
  wire       [0:0]    _zz_2050;
  wire       [31:0]   _zz_2051;
  wire       [31:0]   _zz_2052;
  wire       [31:0]   _zz_2053;
  wire       [0:0]    _zz_2054;
  wire       [0:0]    _zz_2055;
  wire       [31:0]   _zz_2056;
  wire       [31:0]   _zz_2057;
  wire       [31:0]   _zz_2058;
  wire       [0:0]    _zz_2059;
  wire       [0:0]    _zz_2060;
  wire       [31:0]   _zz_2061;
  wire       [31:0]   _zz_2062;
  wire       [31:0]   _zz_2063;
  wire       [0:0]    _zz_2064;
  wire       [0:0]    _zz_2065;
  wire       [31:0]   _zz_2066;
  wire       [31:0]   _zz_2067;
  wire       [31:0]   _zz_2068;
  wire       [0:0]    _zz_2069;
  wire       [0:0]    _zz_2070;
  wire       [31:0]   _zz_2071;
  wire       [31:0]   _zz_2072;
  wire       [31:0]   _zz_2073;
  wire       [0:0]    _zz_2074;
  wire       [0:0]    _zz_2075;
  wire       [31:0]   _zz_2076;
  wire       [31:0]   _zz_2077;
  wire       [31:0]   _zz_2078;
  wire       [0:0]    _zz_2079;
  wire       [0:0]    _zz_2080;
  wire       [31:0]   _zz_2081;
  wire       [31:0]   _zz_2082;
  wire       [31:0]   _zz_2083;
  wire       [0:0]    _zz_2084;
  wire       [0:0]    _zz_2085;
  wire       [31:0]   _zz_2086;
  wire       [31:0]   _zz_2087;
  wire       [31:0]   _zz_2088;
  wire       [0:0]    _zz_2089;
  wire       [0:0]    _zz_2090;
  wire       [31:0]   _zz_2091;
  wire       [31:0]   _zz_2092;
  wire       [31:0]   _zz_2093;
  wire       [0:0]    _zz_2094;
  wire       [0:0]    _zz_2095;
  wire       [31:0]   _zz_2096;
  wire       [31:0]   _zz_2097;
  wire       [31:0]   _zz_2098;
  wire       [0:0]    _zz_2099;
  wire       [0:0]    _zz_2100;
  wire       [31:0]   _zz_2101;
  wire       [31:0]   _zz_2102;
  wire       [31:0]   _zz_2103;
  wire       [0:0]    _zz_2104;
  wire       [0:0]    _zz_2105;
  wire       [31:0]   _zz_2106;
  wire       [31:0]   _zz_2107;
  wire       [31:0]   _zz_2108;
  wire       [0:0]    _zz_2109;
  wire       [0:0]    _zz_2110;
  wire       [31:0]   _zz_2111;
  wire       [31:0]   _zz_2112;
  wire       [31:0]   _zz_2113;
  wire       [0:0]    _zz_2114;
  wire       [0:0]    _zz_2115;
  wire       [31:0]   _zz_2116;
  wire       [31:0]   _zz_2117;
  wire       [31:0]   _zz_2118;
  wire       [0:0]    _zz_2119;
  wire       [0:0]    _zz_2120;
  wire       [31:0]   _zz_2121;
  wire       [31:0]   _zz_2122;
  wire       [31:0]   _zz_2123;
  wire       [0:0]    _zz_2124;
  wire       [0:0]    _zz_2125;
  wire       [31:0]   _zz_2126;
  wire       [31:0]   _zz_2127;
  wire       [31:0]   _zz_2128;
  wire       [0:0]    _zz_2129;
  wire       [0:0]    _zz_2130;
  wire       [31:0]   _zz_2131;
  wire       [31:0]   _zz_2132;
  wire       [31:0]   _zz_2133;
  wire       [0:0]    _zz_2134;
  wire       [0:0]    _zz_2135;
  wire       [31:0]   _zz_2136;
  wire       [31:0]   _zz_2137;
  wire       [31:0]   _zz_2138;
  wire       [0:0]    _zz_2139;
  wire       [0:0]    _zz_2140;
  wire       [31:0]   _zz_2141;
  wire       [31:0]   _zz_2142;
  wire       [31:0]   _zz_2143;
  wire       [0:0]    _zz_2144;
  wire       [0:0]    _zz_2145;
  wire       [31:0]   _zz_2146;
  wire       [31:0]   _zz_2147;
  wire       [31:0]   _zz_2148;
  wire       [0:0]    _zz_2149;
  wire       [0:0]    _zz_2150;
  wire       [31:0]   _zz_2151;
  wire       [31:0]   _zz_2152;
  wire       [31:0]   _zz_2153;
  wire       [0:0]    _zz_2154;
  wire       [0:0]    _zz_2155;
  wire       [31:0]   _zz_2156;
  wire       [31:0]   _zz_2157;
  wire       [31:0]   _zz_2158;
  wire       [0:0]    _zz_2159;
  wire       [0:0]    _zz_2160;
  wire       [31:0]   _zz_2161;
  wire       [31:0]   _zz_2162;
  wire       [31:0]   _zz_2163;
  wire       [0:0]    _zz_2164;
  wire       [0:0]    _zz_2165;
  wire       [31:0]   _zz_2166;
  wire       [31:0]   _zz_2167;
  wire       [31:0]   _zz_2168;
  wire       [0:0]    _zz_2169;
  wire       [0:0]    _zz_2170;
  wire       [31:0]   _zz_2171;
  wire       [31:0]   _zz_2172;
  wire       [31:0]   _zz_2173;
  wire       [0:0]    _zz_2174;
  wire       [0:0]    _zz_2175;
  wire       [31:0]   _zz_2176;
  wire       [31:0]   _zz_2177;
  wire       [31:0]   _zz_2178;
  wire       [0:0]    _zz_2179;
  wire       [0:0]    _zz_2180;
  wire       [31:0]   _zz_2181;
  wire       [31:0]   _zz_2182;
  wire       [31:0]   _zz_2183;
  wire       [0:0]    _zz_2184;
  wire       [0:0]    _zz_2185;
  wire       [31:0]   _zz_2186;
  wire       [31:0]   _zz_2187;
  wire       [31:0]   _zz_2188;
  wire       [0:0]    _zz_2189;
  wire       [0:0]    _zz_2190;
  wire       [31:0]   _zz_2191;
  wire       [31:0]   _zz_2192;
  wire       [31:0]   _zz_2193;
  wire       [0:0]    _zz_2194;
  wire       [0:0]    _zz_2195;
  wire       [31:0]   _zz_2196;
  wire       [31:0]   _zz_2197;
  wire       [31:0]   _zz_2198;
  wire       [0:0]    _zz_2199;
  wire       [0:0]    _zz_2200;
  wire       [31:0]   _zz_2201;
  wire       [31:0]   _zz_2202;
  wire       [31:0]   _zz_2203;
  wire       [0:0]    _zz_2204;
  wire       [0:0]    _zz_2205;
  wire       [31:0]   _zz_2206;
  wire       [31:0]   _zz_2207;
  wire       [31:0]   _zz_2208;
  wire       [0:0]    _zz_2209;
  wire       [0:0]    _zz_2210;
  wire       [31:0]   _zz_2211;
  wire       [31:0]   _zz_2212;
  wire       [31:0]   _zz_2213;
  wire       [0:0]    _zz_2214;
  wire       [0:0]    _zz_2215;
  wire       [31:0]   _zz_2216;
  wire       [31:0]   _zz_2217;
  wire       [31:0]   _zz_2218;
  wire       [0:0]    _zz_2219;
  wire       [0:0]    _zz_2220;
  wire       [31:0]   _zz_2221;
  wire       [31:0]   _zz_2222;
  wire       [31:0]   _zz_2223;
  wire       [0:0]    _zz_2224;
  wire       [0:0]    _zz_2225;
  wire       [31:0]   _zz_2226;
  wire       [31:0]   _zz_2227;
  wire       [31:0]   _zz_2228;
  wire       [0:0]    _zz_2229;
  wire       [0:0]    _zz_2230;
  wire       [31:0]   _zz_2231;
  wire       [31:0]   _zz_2232;
  wire       [31:0]   _zz_2233;
  wire       [0:0]    _zz_2234;
  wire       [0:0]    _zz_2235;
  wire       [31:0]   _zz_2236;
  wire       [31:0]   _zz_2237;
  wire       [31:0]   _zz_2238;
  wire       [0:0]    _zz_2239;
  wire       [0:0]    _zz_2240;
  reg                 current_level_willOverflow_regNext;

  assign _zz_4929 = current_level_willIncrement;
  assign _zz_4930 = {2'd0, _zz_4929};
  assign _zz_4931 = ($signed(twiddle_factor_table_0_real) + $signed(twiddle_factor_table_0_imag));
  assign _zz_4932 = ($signed(_zz_3) - $signed(_zz_4933));
  assign _zz_4933 = ($signed(_zz_4934) * $signed(twiddle_factor_table_0_imag));
  assign _zz_4934 = ($signed(data_mid_1_real) + $signed(data_mid_1_imag));
  assign _zz_4935 = fixTo_dout;
  assign _zz_4936 = ($signed(_zz_3) + $signed(_zz_4937));
  assign _zz_4937 = ($signed(_zz_4938) * $signed(twiddle_factor_table_0_real));
  assign _zz_4938 = ($signed(data_mid_1_imag) - $signed(data_mid_1_real));
  assign _zz_4939 = fixTo_1_dout;
  assign _zz_4940 = _zz_4941[31 : 0];
  assign _zz_4941 = _zz_4942;
  assign _zz_4942 = ($signed(_zz_4943) >>> _zz_4);
  assign _zz_4943 = _zz_4944;
  assign _zz_4944 = ($signed(_zz_4946) - $signed(_zz_1));
  assign _zz_4945 = ({8'd0,data_mid_0_real} <<< 8);
  assign _zz_4946 = {{8{_zz_4945[23]}}, _zz_4945};
  assign _zz_4947 = fixTo_2_dout;
  assign _zz_4948 = _zz_4949[31 : 0];
  assign _zz_4949 = _zz_4950;
  assign _zz_4950 = ($signed(_zz_4951) >>> _zz_4);
  assign _zz_4951 = _zz_4952;
  assign _zz_4952 = ($signed(_zz_4954) - $signed(_zz_2));
  assign _zz_4953 = ({8'd0,data_mid_0_imag} <<< 8);
  assign _zz_4954 = {{8{_zz_4953[23]}}, _zz_4953};
  assign _zz_4955 = fixTo_3_dout;
  assign _zz_4956 = _zz_4957[31 : 0];
  assign _zz_4957 = _zz_4958;
  assign _zz_4958 = ($signed(_zz_4959) >>> _zz_5);
  assign _zz_4959 = _zz_4960;
  assign _zz_4960 = ($signed(_zz_4962) + $signed(_zz_1));
  assign _zz_4961 = ({8'd0,data_mid_0_real} <<< 8);
  assign _zz_4962 = {{8{_zz_4961[23]}}, _zz_4961};
  assign _zz_4963 = fixTo_4_dout;
  assign _zz_4964 = _zz_4965[31 : 0];
  assign _zz_4965 = _zz_4966;
  assign _zz_4966 = ($signed(_zz_4967) >>> _zz_5);
  assign _zz_4967 = _zz_4968;
  assign _zz_4968 = ($signed(_zz_4970) + $signed(_zz_2));
  assign _zz_4969 = ({8'd0,data_mid_0_imag} <<< 8);
  assign _zz_4970 = {{8{_zz_4969[23]}}, _zz_4969};
  assign _zz_4971 = fixTo_5_dout;
  assign _zz_4972 = ($signed(twiddle_factor_table_0_real) + $signed(twiddle_factor_table_0_imag));
  assign _zz_4973 = ($signed(_zz_8) - $signed(_zz_4974));
  assign _zz_4974 = ($signed(_zz_4975) * $signed(twiddle_factor_table_0_imag));
  assign _zz_4975 = ($signed(data_mid_3_real) + $signed(data_mid_3_imag));
  assign _zz_4976 = fixTo_6_dout;
  assign _zz_4977 = ($signed(_zz_8) + $signed(_zz_4978));
  assign _zz_4978 = ($signed(_zz_4979) * $signed(twiddle_factor_table_0_real));
  assign _zz_4979 = ($signed(data_mid_3_imag) - $signed(data_mid_3_real));
  assign _zz_4980 = fixTo_7_dout;
  assign _zz_4981 = _zz_4982[31 : 0];
  assign _zz_4982 = _zz_4983;
  assign _zz_4983 = ($signed(_zz_4984) >>> _zz_9);
  assign _zz_4984 = _zz_4985;
  assign _zz_4985 = ($signed(_zz_4987) - $signed(_zz_6));
  assign _zz_4986 = ({8'd0,data_mid_2_real} <<< 8);
  assign _zz_4987 = {{8{_zz_4986[23]}}, _zz_4986};
  assign _zz_4988 = fixTo_8_dout;
  assign _zz_4989 = _zz_4990[31 : 0];
  assign _zz_4990 = _zz_4991;
  assign _zz_4991 = ($signed(_zz_4992) >>> _zz_9);
  assign _zz_4992 = _zz_4993;
  assign _zz_4993 = ($signed(_zz_4995) - $signed(_zz_7));
  assign _zz_4994 = ({8'd0,data_mid_2_imag} <<< 8);
  assign _zz_4995 = {{8{_zz_4994[23]}}, _zz_4994};
  assign _zz_4996 = fixTo_9_dout;
  assign _zz_4997 = _zz_4998[31 : 0];
  assign _zz_4998 = _zz_4999;
  assign _zz_4999 = ($signed(_zz_5000) >>> _zz_10);
  assign _zz_5000 = _zz_5001;
  assign _zz_5001 = ($signed(_zz_5003) + $signed(_zz_6));
  assign _zz_5002 = ({8'd0,data_mid_2_real} <<< 8);
  assign _zz_5003 = {{8{_zz_5002[23]}}, _zz_5002};
  assign _zz_5004 = fixTo_10_dout;
  assign _zz_5005 = _zz_5006[31 : 0];
  assign _zz_5006 = _zz_5007;
  assign _zz_5007 = ($signed(_zz_5008) >>> _zz_10);
  assign _zz_5008 = _zz_5009;
  assign _zz_5009 = ($signed(_zz_5011) + $signed(_zz_7));
  assign _zz_5010 = ({8'd0,data_mid_2_imag} <<< 8);
  assign _zz_5011 = {{8{_zz_5010[23]}}, _zz_5010};
  assign _zz_5012 = fixTo_11_dout;
  assign _zz_5013 = ($signed(twiddle_factor_table_0_real) + $signed(twiddle_factor_table_0_imag));
  assign _zz_5014 = ($signed(_zz_13) - $signed(_zz_5015));
  assign _zz_5015 = ($signed(_zz_5016) * $signed(twiddle_factor_table_0_imag));
  assign _zz_5016 = ($signed(data_mid_5_real) + $signed(data_mid_5_imag));
  assign _zz_5017 = fixTo_12_dout;
  assign _zz_5018 = ($signed(_zz_13) + $signed(_zz_5019));
  assign _zz_5019 = ($signed(_zz_5020) * $signed(twiddle_factor_table_0_real));
  assign _zz_5020 = ($signed(data_mid_5_imag) - $signed(data_mid_5_real));
  assign _zz_5021 = fixTo_13_dout;
  assign _zz_5022 = _zz_5023[31 : 0];
  assign _zz_5023 = _zz_5024;
  assign _zz_5024 = ($signed(_zz_5025) >>> _zz_14);
  assign _zz_5025 = _zz_5026;
  assign _zz_5026 = ($signed(_zz_5028) - $signed(_zz_11));
  assign _zz_5027 = ({8'd0,data_mid_4_real} <<< 8);
  assign _zz_5028 = {{8{_zz_5027[23]}}, _zz_5027};
  assign _zz_5029 = fixTo_14_dout;
  assign _zz_5030 = _zz_5031[31 : 0];
  assign _zz_5031 = _zz_5032;
  assign _zz_5032 = ($signed(_zz_5033) >>> _zz_14);
  assign _zz_5033 = _zz_5034;
  assign _zz_5034 = ($signed(_zz_5036) - $signed(_zz_12));
  assign _zz_5035 = ({8'd0,data_mid_4_imag} <<< 8);
  assign _zz_5036 = {{8{_zz_5035[23]}}, _zz_5035};
  assign _zz_5037 = fixTo_15_dout;
  assign _zz_5038 = _zz_5039[31 : 0];
  assign _zz_5039 = _zz_5040;
  assign _zz_5040 = ($signed(_zz_5041) >>> _zz_15);
  assign _zz_5041 = _zz_5042;
  assign _zz_5042 = ($signed(_zz_5044) + $signed(_zz_11));
  assign _zz_5043 = ({8'd0,data_mid_4_real} <<< 8);
  assign _zz_5044 = {{8{_zz_5043[23]}}, _zz_5043};
  assign _zz_5045 = fixTo_16_dout;
  assign _zz_5046 = _zz_5047[31 : 0];
  assign _zz_5047 = _zz_5048;
  assign _zz_5048 = ($signed(_zz_5049) >>> _zz_15);
  assign _zz_5049 = _zz_5050;
  assign _zz_5050 = ($signed(_zz_5052) + $signed(_zz_12));
  assign _zz_5051 = ({8'd0,data_mid_4_imag} <<< 8);
  assign _zz_5052 = {{8{_zz_5051[23]}}, _zz_5051};
  assign _zz_5053 = fixTo_17_dout;
  assign _zz_5054 = ($signed(twiddle_factor_table_0_real) + $signed(twiddle_factor_table_0_imag));
  assign _zz_5055 = ($signed(_zz_18) - $signed(_zz_5056));
  assign _zz_5056 = ($signed(_zz_5057) * $signed(twiddle_factor_table_0_imag));
  assign _zz_5057 = ($signed(data_mid_7_real) + $signed(data_mid_7_imag));
  assign _zz_5058 = fixTo_18_dout;
  assign _zz_5059 = ($signed(_zz_18) + $signed(_zz_5060));
  assign _zz_5060 = ($signed(_zz_5061) * $signed(twiddle_factor_table_0_real));
  assign _zz_5061 = ($signed(data_mid_7_imag) - $signed(data_mid_7_real));
  assign _zz_5062 = fixTo_19_dout;
  assign _zz_5063 = _zz_5064[31 : 0];
  assign _zz_5064 = _zz_5065;
  assign _zz_5065 = ($signed(_zz_5066) >>> _zz_19);
  assign _zz_5066 = _zz_5067;
  assign _zz_5067 = ($signed(_zz_5069) - $signed(_zz_16));
  assign _zz_5068 = ({8'd0,data_mid_6_real} <<< 8);
  assign _zz_5069 = {{8{_zz_5068[23]}}, _zz_5068};
  assign _zz_5070 = fixTo_20_dout;
  assign _zz_5071 = _zz_5072[31 : 0];
  assign _zz_5072 = _zz_5073;
  assign _zz_5073 = ($signed(_zz_5074) >>> _zz_19);
  assign _zz_5074 = _zz_5075;
  assign _zz_5075 = ($signed(_zz_5077) - $signed(_zz_17));
  assign _zz_5076 = ({8'd0,data_mid_6_imag} <<< 8);
  assign _zz_5077 = {{8{_zz_5076[23]}}, _zz_5076};
  assign _zz_5078 = fixTo_21_dout;
  assign _zz_5079 = _zz_5080[31 : 0];
  assign _zz_5080 = _zz_5081;
  assign _zz_5081 = ($signed(_zz_5082) >>> _zz_20);
  assign _zz_5082 = _zz_5083;
  assign _zz_5083 = ($signed(_zz_5085) + $signed(_zz_16));
  assign _zz_5084 = ({8'd0,data_mid_6_real} <<< 8);
  assign _zz_5085 = {{8{_zz_5084[23]}}, _zz_5084};
  assign _zz_5086 = fixTo_22_dout;
  assign _zz_5087 = _zz_5088[31 : 0];
  assign _zz_5088 = _zz_5089;
  assign _zz_5089 = ($signed(_zz_5090) >>> _zz_20);
  assign _zz_5090 = _zz_5091;
  assign _zz_5091 = ($signed(_zz_5093) + $signed(_zz_17));
  assign _zz_5092 = ({8'd0,data_mid_6_imag} <<< 8);
  assign _zz_5093 = {{8{_zz_5092[23]}}, _zz_5092};
  assign _zz_5094 = fixTo_23_dout;
  assign _zz_5095 = ($signed(twiddle_factor_table_0_real) + $signed(twiddle_factor_table_0_imag));
  assign _zz_5096 = ($signed(_zz_23) - $signed(_zz_5097));
  assign _zz_5097 = ($signed(_zz_5098) * $signed(twiddle_factor_table_0_imag));
  assign _zz_5098 = ($signed(data_mid_9_real) + $signed(data_mid_9_imag));
  assign _zz_5099 = fixTo_24_dout;
  assign _zz_5100 = ($signed(_zz_23) + $signed(_zz_5101));
  assign _zz_5101 = ($signed(_zz_5102) * $signed(twiddle_factor_table_0_real));
  assign _zz_5102 = ($signed(data_mid_9_imag) - $signed(data_mid_9_real));
  assign _zz_5103 = fixTo_25_dout;
  assign _zz_5104 = _zz_5105[31 : 0];
  assign _zz_5105 = _zz_5106;
  assign _zz_5106 = ($signed(_zz_5107) >>> _zz_24);
  assign _zz_5107 = _zz_5108;
  assign _zz_5108 = ($signed(_zz_5110) - $signed(_zz_21));
  assign _zz_5109 = ({8'd0,data_mid_8_real} <<< 8);
  assign _zz_5110 = {{8{_zz_5109[23]}}, _zz_5109};
  assign _zz_5111 = fixTo_26_dout;
  assign _zz_5112 = _zz_5113[31 : 0];
  assign _zz_5113 = _zz_5114;
  assign _zz_5114 = ($signed(_zz_5115) >>> _zz_24);
  assign _zz_5115 = _zz_5116;
  assign _zz_5116 = ($signed(_zz_5118) - $signed(_zz_22));
  assign _zz_5117 = ({8'd0,data_mid_8_imag} <<< 8);
  assign _zz_5118 = {{8{_zz_5117[23]}}, _zz_5117};
  assign _zz_5119 = fixTo_27_dout;
  assign _zz_5120 = _zz_5121[31 : 0];
  assign _zz_5121 = _zz_5122;
  assign _zz_5122 = ($signed(_zz_5123) >>> _zz_25);
  assign _zz_5123 = _zz_5124;
  assign _zz_5124 = ($signed(_zz_5126) + $signed(_zz_21));
  assign _zz_5125 = ({8'd0,data_mid_8_real} <<< 8);
  assign _zz_5126 = {{8{_zz_5125[23]}}, _zz_5125};
  assign _zz_5127 = fixTo_28_dout;
  assign _zz_5128 = _zz_5129[31 : 0];
  assign _zz_5129 = _zz_5130;
  assign _zz_5130 = ($signed(_zz_5131) >>> _zz_25);
  assign _zz_5131 = _zz_5132;
  assign _zz_5132 = ($signed(_zz_5134) + $signed(_zz_22));
  assign _zz_5133 = ({8'd0,data_mid_8_imag} <<< 8);
  assign _zz_5134 = {{8{_zz_5133[23]}}, _zz_5133};
  assign _zz_5135 = fixTo_29_dout;
  assign _zz_5136 = ($signed(twiddle_factor_table_0_real) + $signed(twiddle_factor_table_0_imag));
  assign _zz_5137 = ($signed(_zz_28) - $signed(_zz_5138));
  assign _zz_5138 = ($signed(_zz_5139) * $signed(twiddle_factor_table_0_imag));
  assign _zz_5139 = ($signed(data_mid_11_real) + $signed(data_mid_11_imag));
  assign _zz_5140 = fixTo_30_dout;
  assign _zz_5141 = ($signed(_zz_28) + $signed(_zz_5142));
  assign _zz_5142 = ($signed(_zz_5143) * $signed(twiddle_factor_table_0_real));
  assign _zz_5143 = ($signed(data_mid_11_imag) - $signed(data_mid_11_real));
  assign _zz_5144 = fixTo_31_dout;
  assign _zz_5145 = _zz_5146[31 : 0];
  assign _zz_5146 = _zz_5147;
  assign _zz_5147 = ($signed(_zz_5148) >>> _zz_29);
  assign _zz_5148 = _zz_5149;
  assign _zz_5149 = ($signed(_zz_5151) - $signed(_zz_26));
  assign _zz_5150 = ({8'd0,data_mid_10_real} <<< 8);
  assign _zz_5151 = {{8{_zz_5150[23]}}, _zz_5150};
  assign _zz_5152 = fixTo_32_dout;
  assign _zz_5153 = _zz_5154[31 : 0];
  assign _zz_5154 = _zz_5155;
  assign _zz_5155 = ($signed(_zz_5156) >>> _zz_29);
  assign _zz_5156 = _zz_5157;
  assign _zz_5157 = ($signed(_zz_5159) - $signed(_zz_27));
  assign _zz_5158 = ({8'd0,data_mid_10_imag} <<< 8);
  assign _zz_5159 = {{8{_zz_5158[23]}}, _zz_5158};
  assign _zz_5160 = fixTo_33_dout;
  assign _zz_5161 = _zz_5162[31 : 0];
  assign _zz_5162 = _zz_5163;
  assign _zz_5163 = ($signed(_zz_5164) >>> _zz_30);
  assign _zz_5164 = _zz_5165;
  assign _zz_5165 = ($signed(_zz_5167) + $signed(_zz_26));
  assign _zz_5166 = ({8'd0,data_mid_10_real} <<< 8);
  assign _zz_5167 = {{8{_zz_5166[23]}}, _zz_5166};
  assign _zz_5168 = fixTo_34_dout;
  assign _zz_5169 = _zz_5170[31 : 0];
  assign _zz_5170 = _zz_5171;
  assign _zz_5171 = ($signed(_zz_5172) >>> _zz_30);
  assign _zz_5172 = _zz_5173;
  assign _zz_5173 = ($signed(_zz_5175) + $signed(_zz_27));
  assign _zz_5174 = ({8'd0,data_mid_10_imag} <<< 8);
  assign _zz_5175 = {{8{_zz_5174[23]}}, _zz_5174};
  assign _zz_5176 = fixTo_35_dout;
  assign _zz_5177 = ($signed(twiddle_factor_table_0_real) + $signed(twiddle_factor_table_0_imag));
  assign _zz_5178 = ($signed(_zz_33) - $signed(_zz_5179));
  assign _zz_5179 = ($signed(_zz_5180) * $signed(twiddle_factor_table_0_imag));
  assign _zz_5180 = ($signed(data_mid_13_real) + $signed(data_mid_13_imag));
  assign _zz_5181 = fixTo_36_dout;
  assign _zz_5182 = ($signed(_zz_33) + $signed(_zz_5183));
  assign _zz_5183 = ($signed(_zz_5184) * $signed(twiddle_factor_table_0_real));
  assign _zz_5184 = ($signed(data_mid_13_imag) - $signed(data_mid_13_real));
  assign _zz_5185 = fixTo_37_dout;
  assign _zz_5186 = _zz_5187[31 : 0];
  assign _zz_5187 = _zz_5188;
  assign _zz_5188 = ($signed(_zz_5189) >>> _zz_34);
  assign _zz_5189 = _zz_5190;
  assign _zz_5190 = ($signed(_zz_5192) - $signed(_zz_31));
  assign _zz_5191 = ({8'd0,data_mid_12_real} <<< 8);
  assign _zz_5192 = {{8{_zz_5191[23]}}, _zz_5191};
  assign _zz_5193 = fixTo_38_dout;
  assign _zz_5194 = _zz_5195[31 : 0];
  assign _zz_5195 = _zz_5196;
  assign _zz_5196 = ($signed(_zz_5197) >>> _zz_34);
  assign _zz_5197 = _zz_5198;
  assign _zz_5198 = ($signed(_zz_5200) - $signed(_zz_32));
  assign _zz_5199 = ({8'd0,data_mid_12_imag} <<< 8);
  assign _zz_5200 = {{8{_zz_5199[23]}}, _zz_5199};
  assign _zz_5201 = fixTo_39_dout;
  assign _zz_5202 = _zz_5203[31 : 0];
  assign _zz_5203 = _zz_5204;
  assign _zz_5204 = ($signed(_zz_5205) >>> _zz_35);
  assign _zz_5205 = _zz_5206;
  assign _zz_5206 = ($signed(_zz_5208) + $signed(_zz_31));
  assign _zz_5207 = ({8'd0,data_mid_12_real} <<< 8);
  assign _zz_5208 = {{8{_zz_5207[23]}}, _zz_5207};
  assign _zz_5209 = fixTo_40_dout;
  assign _zz_5210 = _zz_5211[31 : 0];
  assign _zz_5211 = _zz_5212;
  assign _zz_5212 = ($signed(_zz_5213) >>> _zz_35);
  assign _zz_5213 = _zz_5214;
  assign _zz_5214 = ($signed(_zz_5216) + $signed(_zz_32));
  assign _zz_5215 = ({8'd0,data_mid_12_imag} <<< 8);
  assign _zz_5216 = {{8{_zz_5215[23]}}, _zz_5215};
  assign _zz_5217 = fixTo_41_dout;
  assign _zz_5218 = ($signed(twiddle_factor_table_0_real) + $signed(twiddle_factor_table_0_imag));
  assign _zz_5219 = ($signed(_zz_38) - $signed(_zz_5220));
  assign _zz_5220 = ($signed(_zz_5221) * $signed(twiddle_factor_table_0_imag));
  assign _zz_5221 = ($signed(data_mid_15_real) + $signed(data_mid_15_imag));
  assign _zz_5222 = fixTo_42_dout;
  assign _zz_5223 = ($signed(_zz_38) + $signed(_zz_5224));
  assign _zz_5224 = ($signed(_zz_5225) * $signed(twiddle_factor_table_0_real));
  assign _zz_5225 = ($signed(data_mid_15_imag) - $signed(data_mid_15_real));
  assign _zz_5226 = fixTo_43_dout;
  assign _zz_5227 = _zz_5228[31 : 0];
  assign _zz_5228 = _zz_5229;
  assign _zz_5229 = ($signed(_zz_5230) >>> _zz_39);
  assign _zz_5230 = _zz_5231;
  assign _zz_5231 = ($signed(_zz_5233) - $signed(_zz_36));
  assign _zz_5232 = ({8'd0,data_mid_14_real} <<< 8);
  assign _zz_5233 = {{8{_zz_5232[23]}}, _zz_5232};
  assign _zz_5234 = fixTo_44_dout;
  assign _zz_5235 = _zz_5236[31 : 0];
  assign _zz_5236 = _zz_5237;
  assign _zz_5237 = ($signed(_zz_5238) >>> _zz_39);
  assign _zz_5238 = _zz_5239;
  assign _zz_5239 = ($signed(_zz_5241) - $signed(_zz_37));
  assign _zz_5240 = ({8'd0,data_mid_14_imag} <<< 8);
  assign _zz_5241 = {{8{_zz_5240[23]}}, _zz_5240};
  assign _zz_5242 = fixTo_45_dout;
  assign _zz_5243 = _zz_5244[31 : 0];
  assign _zz_5244 = _zz_5245;
  assign _zz_5245 = ($signed(_zz_5246) >>> _zz_40);
  assign _zz_5246 = _zz_5247;
  assign _zz_5247 = ($signed(_zz_5249) + $signed(_zz_36));
  assign _zz_5248 = ({8'd0,data_mid_14_real} <<< 8);
  assign _zz_5249 = {{8{_zz_5248[23]}}, _zz_5248};
  assign _zz_5250 = fixTo_46_dout;
  assign _zz_5251 = _zz_5252[31 : 0];
  assign _zz_5252 = _zz_5253;
  assign _zz_5253 = ($signed(_zz_5254) >>> _zz_40);
  assign _zz_5254 = _zz_5255;
  assign _zz_5255 = ($signed(_zz_5257) + $signed(_zz_37));
  assign _zz_5256 = ({8'd0,data_mid_14_imag} <<< 8);
  assign _zz_5257 = {{8{_zz_5256[23]}}, _zz_5256};
  assign _zz_5258 = fixTo_47_dout;
  assign _zz_5259 = ($signed(twiddle_factor_table_0_real) + $signed(twiddle_factor_table_0_imag));
  assign _zz_5260 = ($signed(_zz_43) - $signed(_zz_5261));
  assign _zz_5261 = ($signed(_zz_5262) * $signed(twiddle_factor_table_0_imag));
  assign _zz_5262 = ($signed(data_mid_17_real) + $signed(data_mid_17_imag));
  assign _zz_5263 = fixTo_48_dout;
  assign _zz_5264 = ($signed(_zz_43) + $signed(_zz_5265));
  assign _zz_5265 = ($signed(_zz_5266) * $signed(twiddle_factor_table_0_real));
  assign _zz_5266 = ($signed(data_mid_17_imag) - $signed(data_mid_17_real));
  assign _zz_5267 = fixTo_49_dout;
  assign _zz_5268 = _zz_5269[31 : 0];
  assign _zz_5269 = _zz_5270;
  assign _zz_5270 = ($signed(_zz_5271) >>> _zz_44);
  assign _zz_5271 = _zz_5272;
  assign _zz_5272 = ($signed(_zz_5274) - $signed(_zz_41));
  assign _zz_5273 = ({8'd0,data_mid_16_real} <<< 8);
  assign _zz_5274 = {{8{_zz_5273[23]}}, _zz_5273};
  assign _zz_5275 = fixTo_50_dout;
  assign _zz_5276 = _zz_5277[31 : 0];
  assign _zz_5277 = _zz_5278;
  assign _zz_5278 = ($signed(_zz_5279) >>> _zz_44);
  assign _zz_5279 = _zz_5280;
  assign _zz_5280 = ($signed(_zz_5282) - $signed(_zz_42));
  assign _zz_5281 = ({8'd0,data_mid_16_imag} <<< 8);
  assign _zz_5282 = {{8{_zz_5281[23]}}, _zz_5281};
  assign _zz_5283 = fixTo_51_dout;
  assign _zz_5284 = _zz_5285[31 : 0];
  assign _zz_5285 = _zz_5286;
  assign _zz_5286 = ($signed(_zz_5287) >>> _zz_45);
  assign _zz_5287 = _zz_5288;
  assign _zz_5288 = ($signed(_zz_5290) + $signed(_zz_41));
  assign _zz_5289 = ({8'd0,data_mid_16_real} <<< 8);
  assign _zz_5290 = {{8{_zz_5289[23]}}, _zz_5289};
  assign _zz_5291 = fixTo_52_dout;
  assign _zz_5292 = _zz_5293[31 : 0];
  assign _zz_5293 = _zz_5294;
  assign _zz_5294 = ($signed(_zz_5295) >>> _zz_45);
  assign _zz_5295 = _zz_5296;
  assign _zz_5296 = ($signed(_zz_5298) + $signed(_zz_42));
  assign _zz_5297 = ({8'd0,data_mid_16_imag} <<< 8);
  assign _zz_5298 = {{8{_zz_5297[23]}}, _zz_5297};
  assign _zz_5299 = fixTo_53_dout;
  assign _zz_5300 = ($signed(twiddle_factor_table_0_real) + $signed(twiddle_factor_table_0_imag));
  assign _zz_5301 = ($signed(_zz_48) - $signed(_zz_5302));
  assign _zz_5302 = ($signed(_zz_5303) * $signed(twiddle_factor_table_0_imag));
  assign _zz_5303 = ($signed(data_mid_19_real) + $signed(data_mid_19_imag));
  assign _zz_5304 = fixTo_54_dout;
  assign _zz_5305 = ($signed(_zz_48) + $signed(_zz_5306));
  assign _zz_5306 = ($signed(_zz_5307) * $signed(twiddle_factor_table_0_real));
  assign _zz_5307 = ($signed(data_mid_19_imag) - $signed(data_mid_19_real));
  assign _zz_5308 = fixTo_55_dout;
  assign _zz_5309 = _zz_5310[31 : 0];
  assign _zz_5310 = _zz_5311;
  assign _zz_5311 = ($signed(_zz_5312) >>> _zz_49);
  assign _zz_5312 = _zz_5313;
  assign _zz_5313 = ($signed(_zz_5315) - $signed(_zz_46));
  assign _zz_5314 = ({8'd0,data_mid_18_real} <<< 8);
  assign _zz_5315 = {{8{_zz_5314[23]}}, _zz_5314};
  assign _zz_5316 = fixTo_56_dout;
  assign _zz_5317 = _zz_5318[31 : 0];
  assign _zz_5318 = _zz_5319;
  assign _zz_5319 = ($signed(_zz_5320) >>> _zz_49);
  assign _zz_5320 = _zz_5321;
  assign _zz_5321 = ($signed(_zz_5323) - $signed(_zz_47));
  assign _zz_5322 = ({8'd0,data_mid_18_imag} <<< 8);
  assign _zz_5323 = {{8{_zz_5322[23]}}, _zz_5322};
  assign _zz_5324 = fixTo_57_dout;
  assign _zz_5325 = _zz_5326[31 : 0];
  assign _zz_5326 = _zz_5327;
  assign _zz_5327 = ($signed(_zz_5328) >>> _zz_50);
  assign _zz_5328 = _zz_5329;
  assign _zz_5329 = ($signed(_zz_5331) + $signed(_zz_46));
  assign _zz_5330 = ({8'd0,data_mid_18_real} <<< 8);
  assign _zz_5331 = {{8{_zz_5330[23]}}, _zz_5330};
  assign _zz_5332 = fixTo_58_dout;
  assign _zz_5333 = _zz_5334[31 : 0];
  assign _zz_5334 = _zz_5335;
  assign _zz_5335 = ($signed(_zz_5336) >>> _zz_50);
  assign _zz_5336 = _zz_5337;
  assign _zz_5337 = ($signed(_zz_5339) + $signed(_zz_47));
  assign _zz_5338 = ({8'd0,data_mid_18_imag} <<< 8);
  assign _zz_5339 = {{8{_zz_5338[23]}}, _zz_5338};
  assign _zz_5340 = fixTo_59_dout;
  assign _zz_5341 = ($signed(twiddle_factor_table_0_real) + $signed(twiddle_factor_table_0_imag));
  assign _zz_5342 = ($signed(_zz_53) - $signed(_zz_5343));
  assign _zz_5343 = ($signed(_zz_5344) * $signed(twiddle_factor_table_0_imag));
  assign _zz_5344 = ($signed(data_mid_21_real) + $signed(data_mid_21_imag));
  assign _zz_5345 = fixTo_60_dout;
  assign _zz_5346 = ($signed(_zz_53) + $signed(_zz_5347));
  assign _zz_5347 = ($signed(_zz_5348) * $signed(twiddle_factor_table_0_real));
  assign _zz_5348 = ($signed(data_mid_21_imag) - $signed(data_mid_21_real));
  assign _zz_5349 = fixTo_61_dout;
  assign _zz_5350 = _zz_5351[31 : 0];
  assign _zz_5351 = _zz_5352;
  assign _zz_5352 = ($signed(_zz_5353) >>> _zz_54);
  assign _zz_5353 = _zz_5354;
  assign _zz_5354 = ($signed(_zz_5356) - $signed(_zz_51));
  assign _zz_5355 = ({8'd0,data_mid_20_real} <<< 8);
  assign _zz_5356 = {{8{_zz_5355[23]}}, _zz_5355};
  assign _zz_5357 = fixTo_62_dout;
  assign _zz_5358 = _zz_5359[31 : 0];
  assign _zz_5359 = _zz_5360;
  assign _zz_5360 = ($signed(_zz_5361) >>> _zz_54);
  assign _zz_5361 = _zz_5362;
  assign _zz_5362 = ($signed(_zz_5364) - $signed(_zz_52));
  assign _zz_5363 = ({8'd0,data_mid_20_imag} <<< 8);
  assign _zz_5364 = {{8{_zz_5363[23]}}, _zz_5363};
  assign _zz_5365 = fixTo_63_dout;
  assign _zz_5366 = _zz_5367[31 : 0];
  assign _zz_5367 = _zz_5368;
  assign _zz_5368 = ($signed(_zz_5369) >>> _zz_55);
  assign _zz_5369 = _zz_5370;
  assign _zz_5370 = ($signed(_zz_5372) + $signed(_zz_51));
  assign _zz_5371 = ({8'd0,data_mid_20_real} <<< 8);
  assign _zz_5372 = {{8{_zz_5371[23]}}, _zz_5371};
  assign _zz_5373 = fixTo_64_dout;
  assign _zz_5374 = _zz_5375[31 : 0];
  assign _zz_5375 = _zz_5376;
  assign _zz_5376 = ($signed(_zz_5377) >>> _zz_55);
  assign _zz_5377 = _zz_5378;
  assign _zz_5378 = ($signed(_zz_5380) + $signed(_zz_52));
  assign _zz_5379 = ({8'd0,data_mid_20_imag} <<< 8);
  assign _zz_5380 = {{8{_zz_5379[23]}}, _zz_5379};
  assign _zz_5381 = fixTo_65_dout;
  assign _zz_5382 = ($signed(twiddle_factor_table_0_real) + $signed(twiddle_factor_table_0_imag));
  assign _zz_5383 = ($signed(_zz_58) - $signed(_zz_5384));
  assign _zz_5384 = ($signed(_zz_5385) * $signed(twiddle_factor_table_0_imag));
  assign _zz_5385 = ($signed(data_mid_23_real) + $signed(data_mid_23_imag));
  assign _zz_5386 = fixTo_66_dout;
  assign _zz_5387 = ($signed(_zz_58) + $signed(_zz_5388));
  assign _zz_5388 = ($signed(_zz_5389) * $signed(twiddle_factor_table_0_real));
  assign _zz_5389 = ($signed(data_mid_23_imag) - $signed(data_mid_23_real));
  assign _zz_5390 = fixTo_67_dout;
  assign _zz_5391 = _zz_5392[31 : 0];
  assign _zz_5392 = _zz_5393;
  assign _zz_5393 = ($signed(_zz_5394) >>> _zz_59);
  assign _zz_5394 = _zz_5395;
  assign _zz_5395 = ($signed(_zz_5397) - $signed(_zz_56));
  assign _zz_5396 = ({8'd0,data_mid_22_real} <<< 8);
  assign _zz_5397 = {{8{_zz_5396[23]}}, _zz_5396};
  assign _zz_5398 = fixTo_68_dout;
  assign _zz_5399 = _zz_5400[31 : 0];
  assign _zz_5400 = _zz_5401;
  assign _zz_5401 = ($signed(_zz_5402) >>> _zz_59);
  assign _zz_5402 = _zz_5403;
  assign _zz_5403 = ($signed(_zz_5405) - $signed(_zz_57));
  assign _zz_5404 = ({8'd0,data_mid_22_imag} <<< 8);
  assign _zz_5405 = {{8{_zz_5404[23]}}, _zz_5404};
  assign _zz_5406 = fixTo_69_dout;
  assign _zz_5407 = _zz_5408[31 : 0];
  assign _zz_5408 = _zz_5409;
  assign _zz_5409 = ($signed(_zz_5410) >>> _zz_60);
  assign _zz_5410 = _zz_5411;
  assign _zz_5411 = ($signed(_zz_5413) + $signed(_zz_56));
  assign _zz_5412 = ({8'd0,data_mid_22_real} <<< 8);
  assign _zz_5413 = {{8{_zz_5412[23]}}, _zz_5412};
  assign _zz_5414 = fixTo_70_dout;
  assign _zz_5415 = _zz_5416[31 : 0];
  assign _zz_5416 = _zz_5417;
  assign _zz_5417 = ($signed(_zz_5418) >>> _zz_60);
  assign _zz_5418 = _zz_5419;
  assign _zz_5419 = ($signed(_zz_5421) + $signed(_zz_57));
  assign _zz_5420 = ({8'd0,data_mid_22_imag} <<< 8);
  assign _zz_5421 = {{8{_zz_5420[23]}}, _zz_5420};
  assign _zz_5422 = fixTo_71_dout;
  assign _zz_5423 = ($signed(twiddle_factor_table_0_real) + $signed(twiddle_factor_table_0_imag));
  assign _zz_5424 = ($signed(_zz_63) - $signed(_zz_5425));
  assign _zz_5425 = ($signed(_zz_5426) * $signed(twiddle_factor_table_0_imag));
  assign _zz_5426 = ($signed(data_mid_25_real) + $signed(data_mid_25_imag));
  assign _zz_5427 = fixTo_72_dout;
  assign _zz_5428 = ($signed(_zz_63) + $signed(_zz_5429));
  assign _zz_5429 = ($signed(_zz_5430) * $signed(twiddle_factor_table_0_real));
  assign _zz_5430 = ($signed(data_mid_25_imag) - $signed(data_mid_25_real));
  assign _zz_5431 = fixTo_73_dout;
  assign _zz_5432 = _zz_5433[31 : 0];
  assign _zz_5433 = _zz_5434;
  assign _zz_5434 = ($signed(_zz_5435) >>> _zz_64);
  assign _zz_5435 = _zz_5436;
  assign _zz_5436 = ($signed(_zz_5438) - $signed(_zz_61));
  assign _zz_5437 = ({8'd0,data_mid_24_real} <<< 8);
  assign _zz_5438 = {{8{_zz_5437[23]}}, _zz_5437};
  assign _zz_5439 = fixTo_74_dout;
  assign _zz_5440 = _zz_5441[31 : 0];
  assign _zz_5441 = _zz_5442;
  assign _zz_5442 = ($signed(_zz_5443) >>> _zz_64);
  assign _zz_5443 = _zz_5444;
  assign _zz_5444 = ($signed(_zz_5446) - $signed(_zz_62));
  assign _zz_5445 = ({8'd0,data_mid_24_imag} <<< 8);
  assign _zz_5446 = {{8{_zz_5445[23]}}, _zz_5445};
  assign _zz_5447 = fixTo_75_dout;
  assign _zz_5448 = _zz_5449[31 : 0];
  assign _zz_5449 = _zz_5450;
  assign _zz_5450 = ($signed(_zz_5451) >>> _zz_65);
  assign _zz_5451 = _zz_5452;
  assign _zz_5452 = ($signed(_zz_5454) + $signed(_zz_61));
  assign _zz_5453 = ({8'd0,data_mid_24_real} <<< 8);
  assign _zz_5454 = {{8{_zz_5453[23]}}, _zz_5453};
  assign _zz_5455 = fixTo_76_dout;
  assign _zz_5456 = _zz_5457[31 : 0];
  assign _zz_5457 = _zz_5458;
  assign _zz_5458 = ($signed(_zz_5459) >>> _zz_65);
  assign _zz_5459 = _zz_5460;
  assign _zz_5460 = ($signed(_zz_5462) + $signed(_zz_62));
  assign _zz_5461 = ({8'd0,data_mid_24_imag} <<< 8);
  assign _zz_5462 = {{8{_zz_5461[23]}}, _zz_5461};
  assign _zz_5463 = fixTo_77_dout;
  assign _zz_5464 = ($signed(twiddle_factor_table_0_real) + $signed(twiddle_factor_table_0_imag));
  assign _zz_5465 = ($signed(_zz_68) - $signed(_zz_5466));
  assign _zz_5466 = ($signed(_zz_5467) * $signed(twiddle_factor_table_0_imag));
  assign _zz_5467 = ($signed(data_mid_27_real) + $signed(data_mid_27_imag));
  assign _zz_5468 = fixTo_78_dout;
  assign _zz_5469 = ($signed(_zz_68) + $signed(_zz_5470));
  assign _zz_5470 = ($signed(_zz_5471) * $signed(twiddle_factor_table_0_real));
  assign _zz_5471 = ($signed(data_mid_27_imag) - $signed(data_mid_27_real));
  assign _zz_5472 = fixTo_79_dout;
  assign _zz_5473 = _zz_5474[31 : 0];
  assign _zz_5474 = _zz_5475;
  assign _zz_5475 = ($signed(_zz_5476) >>> _zz_69);
  assign _zz_5476 = _zz_5477;
  assign _zz_5477 = ($signed(_zz_5479) - $signed(_zz_66));
  assign _zz_5478 = ({8'd0,data_mid_26_real} <<< 8);
  assign _zz_5479 = {{8{_zz_5478[23]}}, _zz_5478};
  assign _zz_5480 = fixTo_80_dout;
  assign _zz_5481 = _zz_5482[31 : 0];
  assign _zz_5482 = _zz_5483;
  assign _zz_5483 = ($signed(_zz_5484) >>> _zz_69);
  assign _zz_5484 = _zz_5485;
  assign _zz_5485 = ($signed(_zz_5487) - $signed(_zz_67));
  assign _zz_5486 = ({8'd0,data_mid_26_imag} <<< 8);
  assign _zz_5487 = {{8{_zz_5486[23]}}, _zz_5486};
  assign _zz_5488 = fixTo_81_dout;
  assign _zz_5489 = _zz_5490[31 : 0];
  assign _zz_5490 = _zz_5491;
  assign _zz_5491 = ($signed(_zz_5492) >>> _zz_70);
  assign _zz_5492 = _zz_5493;
  assign _zz_5493 = ($signed(_zz_5495) + $signed(_zz_66));
  assign _zz_5494 = ({8'd0,data_mid_26_real} <<< 8);
  assign _zz_5495 = {{8{_zz_5494[23]}}, _zz_5494};
  assign _zz_5496 = fixTo_82_dout;
  assign _zz_5497 = _zz_5498[31 : 0];
  assign _zz_5498 = _zz_5499;
  assign _zz_5499 = ($signed(_zz_5500) >>> _zz_70);
  assign _zz_5500 = _zz_5501;
  assign _zz_5501 = ($signed(_zz_5503) + $signed(_zz_67));
  assign _zz_5502 = ({8'd0,data_mid_26_imag} <<< 8);
  assign _zz_5503 = {{8{_zz_5502[23]}}, _zz_5502};
  assign _zz_5504 = fixTo_83_dout;
  assign _zz_5505 = ($signed(twiddle_factor_table_0_real) + $signed(twiddle_factor_table_0_imag));
  assign _zz_5506 = ($signed(_zz_73) - $signed(_zz_5507));
  assign _zz_5507 = ($signed(_zz_5508) * $signed(twiddle_factor_table_0_imag));
  assign _zz_5508 = ($signed(data_mid_29_real) + $signed(data_mid_29_imag));
  assign _zz_5509 = fixTo_84_dout;
  assign _zz_5510 = ($signed(_zz_73) + $signed(_zz_5511));
  assign _zz_5511 = ($signed(_zz_5512) * $signed(twiddle_factor_table_0_real));
  assign _zz_5512 = ($signed(data_mid_29_imag) - $signed(data_mid_29_real));
  assign _zz_5513 = fixTo_85_dout;
  assign _zz_5514 = _zz_5515[31 : 0];
  assign _zz_5515 = _zz_5516;
  assign _zz_5516 = ($signed(_zz_5517) >>> _zz_74);
  assign _zz_5517 = _zz_5518;
  assign _zz_5518 = ($signed(_zz_5520) - $signed(_zz_71));
  assign _zz_5519 = ({8'd0,data_mid_28_real} <<< 8);
  assign _zz_5520 = {{8{_zz_5519[23]}}, _zz_5519};
  assign _zz_5521 = fixTo_86_dout;
  assign _zz_5522 = _zz_5523[31 : 0];
  assign _zz_5523 = _zz_5524;
  assign _zz_5524 = ($signed(_zz_5525) >>> _zz_74);
  assign _zz_5525 = _zz_5526;
  assign _zz_5526 = ($signed(_zz_5528) - $signed(_zz_72));
  assign _zz_5527 = ({8'd0,data_mid_28_imag} <<< 8);
  assign _zz_5528 = {{8{_zz_5527[23]}}, _zz_5527};
  assign _zz_5529 = fixTo_87_dout;
  assign _zz_5530 = _zz_5531[31 : 0];
  assign _zz_5531 = _zz_5532;
  assign _zz_5532 = ($signed(_zz_5533) >>> _zz_75);
  assign _zz_5533 = _zz_5534;
  assign _zz_5534 = ($signed(_zz_5536) + $signed(_zz_71));
  assign _zz_5535 = ({8'd0,data_mid_28_real} <<< 8);
  assign _zz_5536 = {{8{_zz_5535[23]}}, _zz_5535};
  assign _zz_5537 = fixTo_88_dout;
  assign _zz_5538 = _zz_5539[31 : 0];
  assign _zz_5539 = _zz_5540;
  assign _zz_5540 = ($signed(_zz_5541) >>> _zz_75);
  assign _zz_5541 = _zz_5542;
  assign _zz_5542 = ($signed(_zz_5544) + $signed(_zz_72));
  assign _zz_5543 = ({8'd0,data_mid_28_imag} <<< 8);
  assign _zz_5544 = {{8{_zz_5543[23]}}, _zz_5543};
  assign _zz_5545 = fixTo_89_dout;
  assign _zz_5546 = ($signed(twiddle_factor_table_0_real) + $signed(twiddle_factor_table_0_imag));
  assign _zz_5547 = ($signed(_zz_78) - $signed(_zz_5548));
  assign _zz_5548 = ($signed(_zz_5549) * $signed(twiddle_factor_table_0_imag));
  assign _zz_5549 = ($signed(data_mid_31_real) + $signed(data_mid_31_imag));
  assign _zz_5550 = fixTo_90_dout;
  assign _zz_5551 = ($signed(_zz_78) + $signed(_zz_5552));
  assign _zz_5552 = ($signed(_zz_5553) * $signed(twiddle_factor_table_0_real));
  assign _zz_5553 = ($signed(data_mid_31_imag) - $signed(data_mid_31_real));
  assign _zz_5554 = fixTo_91_dout;
  assign _zz_5555 = _zz_5556[31 : 0];
  assign _zz_5556 = _zz_5557;
  assign _zz_5557 = ($signed(_zz_5558) >>> _zz_79);
  assign _zz_5558 = _zz_5559;
  assign _zz_5559 = ($signed(_zz_5561) - $signed(_zz_76));
  assign _zz_5560 = ({8'd0,data_mid_30_real} <<< 8);
  assign _zz_5561 = {{8{_zz_5560[23]}}, _zz_5560};
  assign _zz_5562 = fixTo_92_dout;
  assign _zz_5563 = _zz_5564[31 : 0];
  assign _zz_5564 = _zz_5565;
  assign _zz_5565 = ($signed(_zz_5566) >>> _zz_79);
  assign _zz_5566 = _zz_5567;
  assign _zz_5567 = ($signed(_zz_5569) - $signed(_zz_77));
  assign _zz_5568 = ({8'd0,data_mid_30_imag} <<< 8);
  assign _zz_5569 = {{8{_zz_5568[23]}}, _zz_5568};
  assign _zz_5570 = fixTo_93_dout;
  assign _zz_5571 = _zz_5572[31 : 0];
  assign _zz_5572 = _zz_5573;
  assign _zz_5573 = ($signed(_zz_5574) >>> _zz_80);
  assign _zz_5574 = _zz_5575;
  assign _zz_5575 = ($signed(_zz_5577) + $signed(_zz_76));
  assign _zz_5576 = ({8'd0,data_mid_30_real} <<< 8);
  assign _zz_5577 = {{8{_zz_5576[23]}}, _zz_5576};
  assign _zz_5578 = fixTo_94_dout;
  assign _zz_5579 = _zz_5580[31 : 0];
  assign _zz_5580 = _zz_5581;
  assign _zz_5581 = ($signed(_zz_5582) >>> _zz_80);
  assign _zz_5582 = _zz_5583;
  assign _zz_5583 = ($signed(_zz_5585) + $signed(_zz_77));
  assign _zz_5584 = ({8'd0,data_mid_30_imag} <<< 8);
  assign _zz_5585 = {{8{_zz_5584[23]}}, _zz_5584};
  assign _zz_5586 = fixTo_95_dout;
  assign _zz_5587 = ($signed(twiddle_factor_table_0_real) + $signed(twiddle_factor_table_0_imag));
  assign _zz_5588 = ($signed(_zz_83) - $signed(_zz_5589));
  assign _zz_5589 = ($signed(_zz_5590) * $signed(twiddle_factor_table_0_imag));
  assign _zz_5590 = ($signed(data_mid_33_real) + $signed(data_mid_33_imag));
  assign _zz_5591 = fixTo_96_dout;
  assign _zz_5592 = ($signed(_zz_83) + $signed(_zz_5593));
  assign _zz_5593 = ($signed(_zz_5594) * $signed(twiddle_factor_table_0_real));
  assign _zz_5594 = ($signed(data_mid_33_imag) - $signed(data_mid_33_real));
  assign _zz_5595 = fixTo_97_dout;
  assign _zz_5596 = _zz_5597[31 : 0];
  assign _zz_5597 = _zz_5598;
  assign _zz_5598 = ($signed(_zz_5599) >>> _zz_84);
  assign _zz_5599 = _zz_5600;
  assign _zz_5600 = ($signed(_zz_5602) - $signed(_zz_81));
  assign _zz_5601 = ({8'd0,data_mid_32_real} <<< 8);
  assign _zz_5602 = {{8{_zz_5601[23]}}, _zz_5601};
  assign _zz_5603 = fixTo_98_dout;
  assign _zz_5604 = _zz_5605[31 : 0];
  assign _zz_5605 = _zz_5606;
  assign _zz_5606 = ($signed(_zz_5607) >>> _zz_84);
  assign _zz_5607 = _zz_5608;
  assign _zz_5608 = ($signed(_zz_5610) - $signed(_zz_82));
  assign _zz_5609 = ({8'd0,data_mid_32_imag} <<< 8);
  assign _zz_5610 = {{8{_zz_5609[23]}}, _zz_5609};
  assign _zz_5611 = fixTo_99_dout;
  assign _zz_5612 = _zz_5613[31 : 0];
  assign _zz_5613 = _zz_5614;
  assign _zz_5614 = ($signed(_zz_5615) >>> _zz_85);
  assign _zz_5615 = _zz_5616;
  assign _zz_5616 = ($signed(_zz_5618) + $signed(_zz_81));
  assign _zz_5617 = ({8'd0,data_mid_32_real} <<< 8);
  assign _zz_5618 = {{8{_zz_5617[23]}}, _zz_5617};
  assign _zz_5619 = fixTo_100_dout;
  assign _zz_5620 = _zz_5621[31 : 0];
  assign _zz_5621 = _zz_5622;
  assign _zz_5622 = ($signed(_zz_5623) >>> _zz_85);
  assign _zz_5623 = _zz_5624;
  assign _zz_5624 = ($signed(_zz_5626) + $signed(_zz_82));
  assign _zz_5625 = ({8'd0,data_mid_32_imag} <<< 8);
  assign _zz_5626 = {{8{_zz_5625[23]}}, _zz_5625};
  assign _zz_5627 = fixTo_101_dout;
  assign _zz_5628 = ($signed(twiddle_factor_table_0_real) + $signed(twiddle_factor_table_0_imag));
  assign _zz_5629 = ($signed(_zz_88) - $signed(_zz_5630));
  assign _zz_5630 = ($signed(_zz_5631) * $signed(twiddle_factor_table_0_imag));
  assign _zz_5631 = ($signed(data_mid_35_real) + $signed(data_mid_35_imag));
  assign _zz_5632 = fixTo_102_dout;
  assign _zz_5633 = ($signed(_zz_88) + $signed(_zz_5634));
  assign _zz_5634 = ($signed(_zz_5635) * $signed(twiddle_factor_table_0_real));
  assign _zz_5635 = ($signed(data_mid_35_imag) - $signed(data_mid_35_real));
  assign _zz_5636 = fixTo_103_dout;
  assign _zz_5637 = _zz_5638[31 : 0];
  assign _zz_5638 = _zz_5639;
  assign _zz_5639 = ($signed(_zz_5640) >>> _zz_89);
  assign _zz_5640 = _zz_5641;
  assign _zz_5641 = ($signed(_zz_5643) - $signed(_zz_86));
  assign _zz_5642 = ({8'd0,data_mid_34_real} <<< 8);
  assign _zz_5643 = {{8{_zz_5642[23]}}, _zz_5642};
  assign _zz_5644 = fixTo_104_dout;
  assign _zz_5645 = _zz_5646[31 : 0];
  assign _zz_5646 = _zz_5647;
  assign _zz_5647 = ($signed(_zz_5648) >>> _zz_89);
  assign _zz_5648 = _zz_5649;
  assign _zz_5649 = ($signed(_zz_5651) - $signed(_zz_87));
  assign _zz_5650 = ({8'd0,data_mid_34_imag} <<< 8);
  assign _zz_5651 = {{8{_zz_5650[23]}}, _zz_5650};
  assign _zz_5652 = fixTo_105_dout;
  assign _zz_5653 = _zz_5654[31 : 0];
  assign _zz_5654 = _zz_5655;
  assign _zz_5655 = ($signed(_zz_5656) >>> _zz_90);
  assign _zz_5656 = _zz_5657;
  assign _zz_5657 = ($signed(_zz_5659) + $signed(_zz_86));
  assign _zz_5658 = ({8'd0,data_mid_34_real} <<< 8);
  assign _zz_5659 = {{8{_zz_5658[23]}}, _zz_5658};
  assign _zz_5660 = fixTo_106_dout;
  assign _zz_5661 = _zz_5662[31 : 0];
  assign _zz_5662 = _zz_5663;
  assign _zz_5663 = ($signed(_zz_5664) >>> _zz_90);
  assign _zz_5664 = _zz_5665;
  assign _zz_5665 = ($signed(_zz_5667) + $signed(_zz_87));
  assign _zz_5666 = ({8'd0,data_mid_34_imag} <<< 8);
  assign _zz_5667 = {{8{_zz_5666[23]}}, _zz_5666};
  assign _zz_5668 = fixTo_107_dout;
  assign _zz_5669 = ($signed(twiddle_factor_table_0_real) + $signed(twiddle_factor_table_0_imag));
  assign _zz_5670 = ($signed(_zz_93) - $signed(_zz_5671));
  assign _zz_5671 = ($signed(_zz_5672) * $signed(twiddle_factor_table_0_imag));
  assign _zz_5672 = ($signed(data_mid_37_real) + $signed(data_mid_37_imag));
  assign _zz_5673 = fixTo_108_dout;
  assign _zz_5674 = ($signed(_zz_93) + $signed(_zz_5675));
  assign _zz_5675 = ($signed(_zz_5676) * $signed(twiddle_factor_table_0_real));
  assign _zz_5676 = ($signed(data_mid_37_imag) - $signed(data_mid_37_real));
  assign _zz_5677 = fixTo_109_dout;
  assign _zz_5678 = _zz_5679[31 : 0];
  assign _zz_5679 = _zz_5680;
  assign _zz_5680 = ($signed(_zz_5681) >>> _zz_94);
  assign _zz_5681 = _zz_5682;
  assign _zz_5682 = ($signed(_zz_5684) - $signed(_zz_91));
  assign _zz_5683 = ({8'd0,data_mid_36_real} <<< 8);
  assign _zz_5684 = {{8{_zz_5683[23]}}, _zz_5683};
  assign _zz_5685 = fixTo_110_dout;
  assign _zz_5686 = _zz_5687[31 : 0];
  assign _zz_5687 = _zz_5688;
  assign _zz_5688 = ($signed(_zz_5689) >>> _zz_94);
  assign _zz_5689 = _zz_5690;
  assign _zz_5690 = ($signed(_zz_5692) - $signed(_zz_92));
  assign _zz_5691 = ({8'd0,data_mid_36_imag} <<< 8);
  assign _zz_5692 = {{8{_zz_5691[23]}}, _zz_5691};
  assign _zz_5693 = fixTo_111_dout;
  assign _zz_5694 = _zz_5695[31 : 0];
  assign _zz_5695 = _zz_5696;
  assign _zz_5696 = ($signed(_zz_5697) >>> _zz_95);
  assign _zz_5697 = _zz_5698;
  assign _zz_5698 = ($signed(_zz_5700) + $signed(_zz_91));
  assign _zz_5699 = ({8'd0,data_mid_36_real} <<< 8);
  assign _zz_5700 = {{8{_zz_5699[23]}}, _zz_5699};
  assign _zz_5701 = fixTo_112_dout;
  assign _zz_5702 = _zz_5703[31 : 0];
  assign _zz_5703 = _zz_5704;
  assign _zz_5704 = ($signed(_zz_5705) >>> _zz_95);
  assign _zz_5705 = _zz_5706;
  assign _zz_5706 = ($signed(_zz_5708) + $signed(_zz_92));
  assign _zz_5707 = ({8'd0,data_mid_36_imag} <<< 8);
  assign _zz_5708 = {{8{_zz_5707[23]}}, _zz_5707};
  assign _zz_5709 = fixTo_113_dout;
  assign _zz_5710 = ($signed(twiddle_factor_table_0_real) + $signed(twiddle_factor_table_0_imag));
  assign _zz_5711 = ($signed(_zz_98) - $signed(_zz_5712));
  assign _zz_5712 = ($signed(_zz_5713) * $signed(twiddle_factor_table_0_imag));
  assign _zz_5713 = ($signed(data_mid_39_real) + $signed(data_mid_39_imag));
  assign _zz_5714 = fixTo_114_dout;
  assign _zz_5715 = ($signed(_zz_98) + $signed(_zz_5716));
  assign _zz_5716 = ($signed(_zz_5717) * $signed(twiddle_factor_table_0_real));
  assign _zz_5717 = ($signed(data_mid_39_imag) - $signed(data_mid_39_real));
  assign _zz_5718 = fixTo_115_dout;
  assign _zz_5719 = _zz_5720[31 : 0];
  assign _zz_5720 = _zz_5721;
  assign _zz_5721 = ($signed(_zz_5722) >>> _zz_99);
  assign _zz_5722 = _zz_5723;
  assign _zz_5723 = ($signed(_zz_5725) - $signed(_zz_96));
  assign _zz_5724 = ({8'd0,data_mid_38_real} <<< 8);
  assign _zz_5725 = {{8{_zz_5724[23]}}, _zz_5724};
  assign _zz_5726 = fixTo_116_dout;
  assign _zz_5727 = _zz_5728[31 : 0];
  assign _zz_5728 = _zz_5729;
  assign _zz_5729 = ($signed(_zz_5730) >>> _zz_99);
  assign _zz_5730 = _zz_5731;
  assign _zz_5731 = ($signed(_zz_5733) - $signed(_zz_97));
  assign _zz_5732 = ({8'd0,data_mid_38_imag} <<< 8);
  assign _zz_5733 = {{8{_zz_5732[23]}}, _zz_5732};
  assign _zz_5734 = fixTo_117_dout;
  assign _zz_5735 = _zz_5736[31 : 0];
  assign _zz_5736 = _zz_5737;
  assign _zz_5737 = ($signed(_zz_5738) >>> _zz_100);
  assign _zz_5738 = _zz_5739;
  assign _zz_5739 = ($signed(_zz_5741) + $signed(_zz_96));
  assign _zz_5740 = ({8'd0,data_mid_38_real} <<< 8);
  assign _zz_5741 = {{8{_zz_5740[23]}}, _zz_5740};
  assign _zz_5742 = fixTo_118_dout;
  assign _zz_5743 = _zz_5744[31 : 0];
  assign _zz_5744 = _zz_5745;
  assign _zz_5745 = ($signed(_zz_5746) >>> _zz_100);
  assign _zz_5746 = _zz_5747;
  assign _zz_5747 = ($signed(_zz_5749) + $signed(_zz_97));
  assign _zz_5748 = ({8'd0,data_mid_38_imag} <<< 8);
  assign _zz_5749 = {{8{_zz_5748[23]}}, _zz_5748};
  assign _zz_5750 = fixTo_119_dout;
  assign _zz_5751 = ($signed(twiddle_factor_table_0_real) + $signed(twiddle_factor_table_0_imag));
  assign _zz_5752 = ($signed(_zz_103) - $signed(_zz_5753));
  assign _zz_5753 = ($signed(_zz_5754) * $signed(twiddle_factor_table_0_imag));
  assign _zz_5754 = ($signed(data_mid_41_real) + $signed(data_mid_41_imag));
  assign _zz_5755 = fixTo_120_dout;
  assign _zz_5756 = ($signed(_zz_103) + $signed(_zz_5757));
  assign _zz_5757 = ($signed(_zz_5758) * $signed(twiddle_factor_table_0_real));
  assign _zz_5758 = ($signed(data_mid_41_imag) - $signed(data_mid_41_real));
  assign _zz_5759 = fixTo_121_dout;
  assign _zz_5760 = _zz_5761[31 : 0];
  assign _zz_5761 = _zz_5762;
  assign _zz_5762 = ($signed(_zz_5763) >>> _zz_104);
  assign _zz_5763 = _zz_5764;
  assign _zz_5764 = ($signed(_zz_5766) - $signed(_zz_101));
  assign _zz_5765 = ({8'd0,data_mid_40_real} <<< 8);
  assign _zz_5766 = {{8{_zz_5765[23]}}, _zz_5765};
  assign _zz_5767 = fixTo_122_dout;
  assign _zz_5768 = _zz_5769[31 : 0];
  assign _zz_5769 = _zz_5770;
  assign _zz_5770 = ($signed(_zz_5771) >>> _zz_104);
  assign _zz_5771 = _zz_5772;
  assign _zz_5772 = ($signed(_zz_5774) - $signed(_zz_102));
  assign _zz_5773 = ({8'd0,data_mid_40_imag} <<< 8);
  assign _zz_5774 = {{8{_zz_5773[23]}}, _zz_5773};
  assign _zz_5775 = fixTo_123_dout;
  assign _zz_5776 = _zz_5777[31 : 0];
  assign _zz_5777 = _zz_5778;
  assign _zz_5778 = ($signed(_zz_5779) >>> _zz_105);
  assign _zz_5779 = _zz_5780;
  assign _zz_5780 = ($signed(_zz_5782) + $signed(_zz_101));
  assign _zz_5781 = ({8'd0,data_mid_40_real} <<< 8);
  assign _zz_5782 = {{8{_zz_5781[23]}}, _zz_5781};
  assign _zz_5783 = fixTo_124_dout;
  assign _zz_5784 = _zz_5785[31 : 0];
  assign _zz_5785 = _zz_5786;
  assign _zz_5786 = ($signed(_zz_5787) >>> _zz_105);
  assign _zz_5787 = _zz_5788;
  assign _zz_5788 = ($signed(_zz_5790) + $signed(_zz_102));
  assign _zz_5789 = ({8'd0,data_mid_40_imag} <<< 8);
  assign _zz_5790 = {{8{_zz_5789[23]}}, _zz_5789};
  assign _zz_5791 = fixTo_125_dout;
  assign _zz_5792 = ($signed(twiddle_factor_table_0_real) + $signed(twiddle_factor_table_0_imag));
  assign _zz_5793 = ($signed(_zz_108) - $signed(_zz_5794));
  assign _zz_5794 = ($signed(_zz_5795) * $signed(twiddle_factor_table_0_imag));
  assign _zz_5795 = ($signed(data_mid_43_real) + $signed(data_mid_43_imag));
  assign _zz_5796 = fixTo_126_dout;
  assign _zz_5797 = ($signed(_zz_108) + $signed(_zz_5798));
  assign _zz_5798 = ($signed(_zz_5799) * $signed(twiddle_factor_table_0_real));
  assign _zz_5799 = ($signed(data_mid_43_imag) - $signed(data_mid_43_real));
  assign _zz_5800 = fixTo_127_dout;
  assign _zz_5801 = _zz_5802[31 : 0];
  assign _zz_5802 = _zz_5803;
  assign _zz_5803 = ($signed(_zz_5804) >>> _zz_109);
  assign _zz_5804 = _zz_5805;
  assign _zz_5805 = ($signed(_zz_5807) - $signed(_zz_106));
  assign _zz_5806 = ({8'd0,data_mid_42_real} <<< 8);
  assign _zz_5807 = {{8{_zz_5806[23]}}, _zz_5806};
  assign _zz_5808 = fixTo_128_dout;
  assign _zz_5809 = _zz_5810[31 : 0];
  assign _zz_5810 = _zz_5811;
  assign _zz_5811 = ($signed(_zz_5812) >>> _zz_109);
  assign _zz_5812 = _zz_5813;
  assign _zz_5813 = ($signed(_zz_5815) - $signed(_zz_107));
  assign _zz_5814 = ({8'd0,data_mid_42_imag} <<< 8);
  assign _zz_5815 = {{8{_zz_5814[23]}}, _zz_5814};
  assign _zz_5816 = fixTo_129_dout;
  assign _zz_5817 = _zz_5818[31 : 0];
  assign _zz_5818 = _zz_5819;
  assign _zz_5819 = ($signed(_zz_5820) >>> _zz_110);
  assign _zz_5820 = _zz_5821;
  assign _zz_5821 = ($signed(_zz_5823) + $signed(_zz_106));
  assign _zz_5822 = ({8'd0,data_mid_42_real} <<< 8);
  assign _zz_5823 = {{8{_zz_5822[23]}}, _zz_5822};
  assign _zz_5824 = fixTo_130_dout;
  assign _zz_5825 = _zz_5826[31 : 0];
  assign _zz_5826 = _zz_5827;
  assign _zz_5827 = ($signed(_zz_5828) >>> _zz_110);
  assign _zz_5828 = _zz_5829;
  assign _zz_5829 = ($signed(_zz_5831) + $signed(_zz_107));
  assign _zz_5830 = ({8'd0,data_mid_42_imag} <<< 8);
  assign _zz_5831 = {{8{_zz_5830[23]}}, _zz_5830};
  assign _zz_5832 = fixTo_131_dout;
  assign _zz_5833 = ($signed(twiddle_factor_table_0_real) + $signed(twiddle_factor_table_0_imag));
  assign _zz_5834 = ($signed(_zz_113) - $signed(_zz_5835));
  assign _zz_5835 = ($signed(_zz_5836) * $signed(twiddle_factor_table_0_imag));
  assign _zz_5836 = ($signed(data_mid_45_real) + $signed(data_mid_45_imag));
  assign _zz_5837 = fixTo_132_dout;
  assign _zz_5838 = ($signed(_zz_113) + $signed(_zz_5839));
  assign _zz_5839 = ($signed(_zz_5840) * $signed(twiddle_factor_table_0_real));
  assign _zz_5840 = ($signed(data_mid_45_imag) - $signed(data_mid_45_real));
  assign _zz_5841 = fixTo_133_dout;
  assign _zz_5842 = _zz_5843[31 : 0];
  assign _zz_5843 = _zz_5844;
  assign _zz_5844 = ($signed(_zz_5845) >>> _zz_114);
  assign _zz_5845 = _zz_5846;
  assign _zz_5846 = ($signed(_zz_5848) - $signed(_zz_111));
  assign _zz_5847 = ({8'd0,data_mid_44_real} <<< 8);
  assign _zz_5848 = {{8{_zz_5847[23]}}, _zz_5847};
  assign _zz_5849 = fixTo_134_dout;
  assign _zz_5850 = _zz_5851[31 : 0];
  assign _zz_5851 = _zz_5852;
  assign _zz_5852 = ($signed(_zz_5853) >>> _zz_114);
  assign _zz_5853 = _zz_5854;
  assign _zz_5854 = ($signed(_zz_5856) - $signed(_zz_112));
  assign _zz_5855 = ({8'd0,data_mid_44_imag} <<< 8);
  assign _zz_5856 = {{8{_zz_5855[23]}}, _zz_5855};
  assign _zz_5857 = fixTo_135_dout;
  assign _zz_5858 = _zz_5859[31 : 0];
  assign _zz_5859 = _zz_5860;
  assign _zz_5860 = ($signed(_zz_5861) >>> _zz_115);
  assign _zz_5861 = _zz_5862;
  assign _zz_5862 = ($signed(_zz_5864) + $signed(_zz_111));
  assign _zz_5863 = ({8'd0,data_mid_44_real} <<< 8);
  assign _zz_5864 = {{8{_zz_5863[23]}}, _zz_5863};
  assign _zz_5865 = fixTo_136_dout;
  assign _zz_5866 = _zz_5867[31 : 0];
  assign _zz_5867 = _zz_5868;
  assign _zz_5868 = ($signed(_zz_5869) >>> _zz_115);
  assign _zz_5869 = _zz_5870;
  assign _zz_5870 = ($signed(_zz_5872) + $signed(_zz_112));
  assign _zz_5871 = ({8'd0,data_mid_44_imag} <<< 8);
  assign _zz_5872 = {{8{_zz_5871[23]}}, _zz_5871};
  assign _zz_5873 = fixTo_137_dout;
  assign _zz_5874 = ($signed(twiddle_factor_table_0_real) + $signed(twiddle_factor_table_0_imag));
  assign _zz_5875 = ($signed(_zz_118) - $signed(_zz_5876));
  assign _zz_5876 = ($signed(_zz_5877) * $signed(twiddle_factor_table_0_imag));
  assign _zz_5877 = ($signed(data_mid_47_real) + $signed(data_mid_47_imag));
  assign _zz_5878 = fixTo_138_dout;
  assign _zz_5879 = ($signed(_zz_118) + $signed(_zz_5880));
  assign _zz_5880 = ($signed(_zz_5881) * $signed(twiddle_factor_table_0_real));
  assign _zz_5881 = ($signed(data_mid_47_imag) - $signed(data_mid_47_real));
  assign _zz_5882 = fixTo_139_dout;
  assign _zz_5883 = _zz_5884[31 : 0];
  assign _zz_5884 = _zz_5885;
  assign _zz_5885 = ($signed(_zz_5886) >>> _zz_119);
  assign _zz_5886 = _zz_5887;
  assign _zz_5887 = ($signed(_zz_5889) - $signed(_zz_116));
  assign _zz_5888 = ({8'd0,data_mid_46_real} <<< 8);
  assign _zz_5889 = {{8{_zz_5888[23]}}, _zz_5888};
  assign _zz_5890 = fixTo_140_dout;
  assign _zz_5891 = _zz_5892[31 : 0];
  assign _zz_5892 = _zz_5893;
  assign _zz_5893 = ($signed(_zz_5894) >>> _zz_119);
  assign _zz_5894 = _zz_5895;
  assign _zz_5895 = ($signed(_zz_5897) - $signed(_zz_117));
  assign _zz_5896 = ({8'd0,data_mid_46_imag} <<< 8);
  assign _zz_5897 = {{8{_zz_5896[23]}}, _zz_5896};
  assign _zz_5898 = fixTo_141_dout;
  assign _zz_5899 = _zz_5900[31 : 0];
  assign _zz_5900 = _zz_5901;
  assign _zz_5901 = ($signed(_zz_5902) >>> _zz_120);
  assign _zz_5902 = _zz_5903;
  assign _zz_5903 = ($signed(_zz_5905) + $signed(_zz_116));
  assign _zz_5904 = ({8'd0,data_mid_46_real} <<< 8);
  assign _zz_5905 = {{8{_zz_5904[23]}}, _zz_5904};
  assign _zz_5906 = fixTo_142_dout;
  assign _zz_5907 = _zz_5908[31 : 0];
  assign _zz_5908 = _zz_5909;
  assign _zz_5909 = ($signed(_zz_5910) >>> _zz_120);
  assign _zz_5910 = _zz_5911;
  assign _zz_5911 = ($signed(_zz_5913) + $signed(_zz_117));
  assign _zz_5912 = ({8'd0,data_mid_46_imag} <<< 8);
  assign _zz_5913 = {{8{_zz_5912[23]}}, _zz_5912};
  assign _zz_5914 = fixTo_143_dout;
  assign _zz_5915 = ($signed(twiddle_factor_table_0_real) + $signed(twiddle_factor_table_0_imag));
  assign _zz_5916 = ($signed(_zz_123) - $signed(_zz_5917));
  assign _zz_5917 = ($signed(_zz_5918) * $signed(twiddle_factor_table_0_imag));
  assign _zz_5918 = ($signed(data_mid_49_real) + $signed(data_mid_49_imag));
  assign _zz_5919 = fixTo_144_dout;
  assign _zz_5920 = ($signed(_zz_123) + $signed(_zz_5921));
  assign _zz_5921 = ($signed(_zz_5922) * $signed(twiddle_factor_table_0_real));
  assign _zz_5922 = ($signed(data_mid_49_imag) - $signed(data_mid_49_real));
  assign _zz_5923 = fixTo_145_dout;
  assign _zz_5924 = _zz_5925[31 : 0];
  assign _zz_5925 = _zz_5926;
  assign _zz_5926 = ($signed(_zz_5927) >>> _zz_124);
  assign _zz_5927 = _zz_5928;
  assign _zz_5928 = ($signed(_zz_5930) - $signed(_zz_121));
  assign _zz_5929 = ({8'd0,data_mid_48_real} <<< 8);
  assign _zz_5930 = {{8{_zz_5929[23]}}, _zz_5929};
  assign _zz_5931 = fixTo_146_dout;
  assign _zz_5932 = _zz_5933[31 : 0];
  assign _zz_5933 = _zz_5934;
  assign _zz_5934 = ($signed(_zz_5935) >>> _zz_124);
  assign _zz_5935 = _zz_5936;
  assign _zz_5936 = ($signed(_zz_5938) - $signed(_zz_122));
  assign _zz_5937 = ({8'd0,data_mid_48_imag} <<< 8);
  assign _zz_5938 = {{8{_zz_5937[23]}}, _zz_5937};
  assign _zz_5939 = fixTo_147_dout;
  assign _zz_5940 = _zz_5941[31 : 0];
  assign _zz_5941 = _zz_5942;
  assign _zz_5942 = ($signed(_zz_5943) >>> _zz_125);
  assign _zz_5943 = _zz_5944;
  assign _zz_5944 = ($signed(_zz_5946) + $signed(_zz_121));
  assign _zz_5945 = ({8'd0,data_mid_48_real} <<< 8);
  assign _zz_5946 = {{8{_zz_5945[23]}}, _zz_5945};
  assign _zz_5947 = fixTo_148_dout;
  assign _zz_5948 = _zz_5949[31 : 0];
  assign _zz_5949 = _zz_5950;
  assign _zz_5950 = ($signed(_zz_5951) >>> _zz_125);
  assign _zz_5951 = _zz_5952;
  assign _zz_5952 = ($signed(_zz_5954) + $signed(_zz_122));
  assign _zz_5953 = ({8'd0,data_mid_48_imag} <<< 8);
  assign _zz_5954 = {{8{_zz_5953[23]}}, _zz_5953};
  assign _zz_5955 = fixTo_149_dout;
  assign _zz_5956 = ($signed(twiddle_factor_table_0_real) + $signed(twiddle_factor_table_0_imag));
  assign _zz_5957 = ($signed(_zz_128) - $signed(_zz_5958));
  assign _zz_5958 = ($signed(_zz_5959) * $signed(twiddle_factor_table_0_imag));
  assign _zz_5959 = ($signed(data_mid_51_real) + $signed(data_mid_51_imag));
  assign _zz_5960 = fixTo_150_dout;
  assign _zz_5961 = ($signed(_zz_128) + $signed(_zz_5962));
  assign _zz_5962 = ($signed(_zz_5963) * $signed(twiddle_factor_table_0_real));
  assign _zz_5963 = ($signed(data_mid_51_imag) - $signed(data_mid_51_real));
  assign _zz_5964 = fixTo_151_dout;
  assign _zz_5965 = _zz_5966[31 : 0];
  assign _zz_5966 = _zz_5967;
  assign _zz_5967 = ($signed(_zz_5968) >>> _zz_129);
  assign _zz_5968 = _zz_5969;
  assign _zz_5969 = ($signed(_zz_5971) - $signed(_zz_126));
  assign _zz_5970 = ({8'd0,data_mid_50_real} <<< 8);
  assign _zz_5971 = {{8{_zz_5970[23]}}, _zz_5970};
  assign _zz_5972 = fixTo_152_dout;
  assign _zz_5973 = _zz_5974[31 : 0];
  assign _zz_5974 = _zz_5975;
  assign _zz_5975 = ($signed(_zz_5976) >>> _zz_129);
  assign _zz_5976 = _zz_5977;
  assign _zz_5977 = ($signed(_zz_5979) - $signed(_zz_127));
  assign _zz_5978 = ({8'd0,data_mid_50_imag} <<< 8);
  assign _zz_5979 = {{8{_zz_5978[23]}}, _zz_5978};
  assign _zz_5980 = fixTo_153_dout;
  assign _zz_5981 = _zz_5982[31 : 0];
  assign _zz_5982 = _zz_5983;
  assign _zz_5983 = ($signed(_zz_5984) >>> _zz_130);
  assign _zz_5984 = _zz_5985;
  assign _zz_5985 = ($signed(_zz_5987) + $signed(_zz_126));
  assign _zz_5986 = ({8'd0,data_mid_50_real} <<< 8);
  assign _zz_5987 = {{8{_zz_5986[23]}}, _zz_5986};
  assign _zz_5988 = fixTo_154_dout;
  assign _zz_5989 = _zz_5990[31 : 0];
  assign _zz_5990 = _zz_5991;
  assign _zz_5991 = ($signed(_zz_5992) >>> _zz_130);
  assign _zz_5992 = _zz_5993;
  assign _zz_5993 = ($signed(_zz_5995) + $signed(_zz_127));
  assign _zz_5994 = ({8'd0,data_mid_50_imag} <<< 8);
  assign _zz_5995 = {{8{_zz_5994[23]}}, _zz_5994};
  assign _zz_5996 = fixTo_155_dout;
  assign _zz_5997 = ($signed(twiddle_factor_table_0_real) + $signed(twiddle_factor_table_0_imag));
  assign _zz_5998 = ($signed(_zz_133) - $signed(_zz_5999));
  assign _zz_5999 = ($signed(_zz_6000) * $signed(twiddle_factor_table_0_imag));
  assign _zz_6000 = ($signed(data_mid_53_real) + $signed(data_mid_53_imag));
  assign _zz_6001 = fixTo_156_dout;
  assign _zz_6002 = ($signed(_zz_133) + $signed(_zz_6003));
  assign _zz_6003 = ($signed(_zz_6004) * $signed(twiddle_factor_table_0_real));
  assign _zz_6004 = ($signed(data_mid_53_imag) - $signed(data_mid_53_real));
  assign _zz_6005 = fixTo_157_dout;
  assign _zz_6006 = _zz_6007[31 : 0];
  assign _zz_6007 = _zz_6008;
  assign _zz_6008 = ($signed(_zz_6009) >>> _zz_134);
  assign _zz_6009 = _zz_6010;
  assign _zz_6010 = ($signed(_zz_6012) - $signed(_zz_131));
  assign _zz_6011 = ({8'd0,data_mid_52_real} <<< 8);
  assign _zz_6012 = {{8{_zz_6011[23]}}, _zz_6011};
  assign _zz_6013 = fixTo_158_dout;
  assign _zz_6014 = _zz_6015[31 : 0];
  assign _zz_6015 = _zz_6016;
  assign _zz_6016 = ($signed(_zz_6017) >>> _zz_134);
  assign _zz_6017 = _zz_6018;
  assign _zz_6018 = ($signed(_zz_6020) - $signed(_zz_132));
  assign _zz_6019 = ({8'd0,data_mid_52_imag} <<< 8);
  assign _zz_6020 = {{8{_zz_6019[23]}}, _zz_6019};
  assign _zz_6021 = fixTo_159_dout;
  assign _zz_6022 = _zz_6023[31 : 0];
  assign _zz_6023 = _zz_6024;
  assign _zz_6024 = ($signed(_zz_6025) >>> _zz_135);
  assign _zz_6025 = _zz_6026;
  assign _zz_6026 = ($signed(_zz_6028) + $signed(_zz_131));
  assign _zz_6027 = ({8'd0,data_mid_52_real} <<< 8);
  assign _zz_6028 = {{8{_zz_6027[23]}}, _zz_6027};
  assign _zz_6029 = fixTo_160_dout;
  assign _zz_6030 = _zz_6031[31 : 0];
  assign _zz_6031 = _zz_6032;
  assign _zz_6032 = ($signed(_zz_6033) >>> _zz_135);
  assign _zz_6033 = _zz_6034;
  assign _zz_6034 = ($signed(_zz_6036) + $signed(_zz_132));
  assign _zz_6035 = ({8'd0,data_mid_52_imag} <<< 8);
  assign _zz_6036 = {{8{_zz_6035[23]}}, _zz_6035};
  assign _zz_6037 = fixTo_161_dout;
  assign _zz_6038 = ($signed(twiddle_factor_table_0_real) + $signed(twiddle_factor_table_0_imag));
  assign _zz_6039 = ($signed(_zz_138) - $signed(_zz_6040));
  assign _zz_6040 = ($signed(_zz_6041) * $signed(twiddle_factor_table_0_imag));
  assign _zz_6041 = ($signed(data_mid_55_real) + $signed(data_mid_55_imag));
  assign _zz_6042 = fixTo_162_dout;
  assign _zz_6043 = ($signed(_zz_138) + $signed(_zz_6044));
  assign _zz_6044 = ($signed(_zz_6045) * $signed(twiddle_factor_table_0_real));
  assign _zz_6045 = ($signed(data_mid_55_imag) - $signed(data_mid_55_real));
  assign _zz_6046 = fixTo_163_dout;
  assign _zz_6047 = _zz_6048[31 : 0];
  assign _zz_6048 = _zz_6049;
  assign _zz_6049 = ($signed(_zz_6050) >>> _zz_139);
  assign _zz_6050 = _zz_6051;
  assign _zz_6051 = ($signed(_zz_6053) - $signed(_zz_136));
  assign _zz_6052 = ({8'd0,data_mid_54_real} <<< 8);
  assign _zz_6053 = {{8{_zz_6052[23]}}, _zz_6052};
  assign _zz_6054 = fixTo_164_dout;
  assign _zz_6055 = _zz_6056[31 : 0];
  assign _zz_6056 = _zz_6057;
  assign _zz_6057 = ($signed(_zz_6058) >>> _zz_139);
  assign _zz_6058 = _zz_6059;
  assign _zz_6059 = ($signed(_zz_6061) - $signed(_zz_137));
  assign _zz_6060 = ({8'd0,data_mid_54_imag} <<< 8);
  assign _zz_6061 = {{8{_zz_6060[23]}}, _zz_6060};
  assign _zz_6062 = fixTo_165_dout;
  assign _zz_6063 = _zz_6064[31 : 0];
  assign _zz_6064 = _zz_6065;
  assign _zz_6065 = ($signed(_zz_6066) >>> _zz_140);
  assign _zz_6066 = _zz_6067;
  assign _zz_6067 = ($signed(_zz_6069) + $signed(_zz_136));
  assign _zz_6068 = ({8'd0,data_mid_54_real} <<< 8);
  assign _zz_6069 = {{8{_zz_6068[23]}}, _zz_6068};
  assign _zz_6070 = fixTo_166_dout;
  assign _zz_6071 = _zz_6072[31 : 0];
  assign _zz_6072 = _zz_6073;
  assign _zz_6073 = ($signed(_zz_6074) >>> _zz_140);
  assign _zz_6074 = _zz_6075;
  assign _zz_6075 = ($signed(_zz_6077) + $signed(_zz_137));
  assign _zz_6076 = ({8'd0,data_mid_54_imag} <<< 8);
  assign _zz_6077 = {{8{_zz_6076[23]}}, _zz_6076};
  assign _zz_6078 = fixTo_167_dout;
  assign _zz_6079 = ($signed(twiddle_factor_table_0_real) + $signed(twiddle_factor_table_0_imag));
  assign _zz_6080 = ($signed(_zz_143) - $signed(_zz_6081));
  assign _zz_6081 = ($signed(_zz_6082) * $signed(twiddle_factor_table_0_imag));
  assign _zz_6082 = ($signed(data_mid_57_real) + $signed(data_mid_57_imag));
  assign _zz_6083 = fixTo_168_dout;
  assign _zz_6084 = ($signed(_zz_143) + $signed(_zz_6085));
  assign _zz_6085 = ($signed(_zz_6086) * $signed(twiddle_factor_table_0_real));
  assign _zz_6086 = ($signed(data_mid_57_imag) - $signed(data_mid_57_real));
  assign _zz_6087 = fixTo_169_dout;
  assign _zz_6088 = _zz_6089[31 : 0];
  assign _zz_6089 = _zz_6090;
  assign _zz_6090 = ($signed(_zz_6091) >>> _zz_144);
  assign _zz_6091 = _zz_6092;
  assign _zz_6092 = ($signed(_zz_6094) - $signed(_zz_141));
  assign _zz_6093 = ({8'd0,data_mid_56_real} <<< 8);
  assign _zz_6094 = {{8{_zz_6093[23]}}, _zz_6093};
  assign _zz_6095 = fixTo_170_dout;
  assign _zz_6096 = _zz_6097[31 : 0];
  assign _zz_6097 = _zz_6098;
  assign _zz_6098 = ($signed(_zz_6099) >>> _zz_144);
  assign _zz_6099 = _zz_6100;
  assign _zz_6100 = ($signed(_zz_6102) - $signed(_zz_142));
  assign _zz_6101 = ({8'd0,data_mid_56_imag} <<< 8);
  assign _zz_6102 = {{8{_zz_6101[23]}}, _zz_6101};
  assign _zz_6103 = fixTo_171_dout;
  assign _zz_6104 = _zz_6105[31 : 0];
  assign _zz_6105 = _zz_6106;
  assign _zz_6106 = ($signed(_zz_6107) >>> _zz_145);
  assign _zz_6107 = _zz_6108;
  assign _zz_6108 = ($signed(_zz_6110) + $signed(_zz_141));
  assign _zz_6109 = ({8'd0,data_mid_56_real} <<< 8);
  assign _zz_6110 = {{8{_zz_6109[23]}}, _zz_6109};
  assign _zz_6111 = fixTo_172_dout;
  assign _zz_6112 = _zz_6113[31 : 0];
  assign _zz_6113 = _zz_6114;
  assign _zz_6114 = ($signed(_zz_6115) >>> _zz_145);
  assign _zz_6115 = _zz_6116;
  assign _zz_6116 = ($signed(_zz_6118) + $signed(_zz_142));
  assign _zz_6117 = ({8'd0,data_mid_56_imag} <<< 8);
  assign _zz_6118 = {{8{_zz_6117[23]}}, _zz_6117};
  assign _zz_6119 = fixTo_173_dout;
  assign _zz_6120 = ($signed(twiddle_factor_table_0_real) + $signed(twiddle_factor_table_0_imag));
  assign _zz_6121 = ($signed(_zz_148) - $signed(_zz_6122));
  assign _zz_6122 = ($signed(_zz_6123) * $signed(twiddle_factor_table_0_imag));
  assign _zz_6123 = ($signed(data_mid_59_real) + $signed(data_mid_59_imag));
  assign _zz_6124 = fixTo_174_dout;
  assign _zz_6125 = ($signed(_zz_148) + $signed(_zz_6126));
  assign _zz_6126 = ($signed(_zz_6127) * $signed(twiddle_factor_table_0_real));
  assign _zz_6127 = ($signed(data_mid_59_imag) - $signed(data_mid_59_real));
  assign _zz_6128 = fixTo_175_dout;
  assign _zz_6129 = _zz_6130[31 : 0];
  assign _zz_6130 = _zz_6131;
  assign _zz_6131 = ($signed(_zz_6132) >>> _zz_149);
  assign _zz_6132 = _zz_6133;
  assign _zz_6133 = ($signed(_zz_6135) - $signed(_zz_146));
  assign _zz_6134 = ({8'd0,data_mid_58_real} <<< 8);
  assign _zz_6135 = {{8{_zz_6134[23]}}, _zz_6134};
  assign _zz_6136 = fixTo_176_dout;
  assign _zz_6137 = _zz_6138[31 : 0];
  assign _zz_6138 = _zz_6139;
  assign _zz_6139 = ($signed(_zz_6140) >>> _zz_149);
  assign _zz_6140 = _zz_6141;
  assign _zz_6141 = ($signed(_zz_6143) - $signed(_zz_147));
  assign _zz_6142 = ({8'd0,data_mid_58_imag} <<< 8);
  assign _zz_6143 = {{8{_zz_6142[23]}}, _zz_6142};
  assign _zz_6144 = fixTo_177_dout;
  assign _zz_6145 = _zz_6146[31 : 0];
  assign _zz_6146 = _zz_6147;
  assign _zz_6147 = ($signed(_zz_6148) >>> _zz_150);
  assign _zz_6148 = _zz_6149;
  assign _zz_6149 = ($signed(_zz_6151) + $signed(_zz_146));
  assign _zz_6150 = ({8'd0,data_mid_58_real} <<< 8);
  assign _zz_6151 = {{8{_zz_6150[23]}}, _zz_6150};
  assign _zz_6152 = fixTo_178_dout;
  assign _zz_6153 = _zz_6154[31 : 0];
  assign _zz_6154 = _zz_6155;
  assign _zz_6155 = ($signed(_zz_6156) >>> _zz_150);
  assign _zz_6156 = _zz_6157;
  assign _zz_6157 = ($signed(_zz_6159) + $signed(_zz_147));
  assign _zz_6158 = ({8'd0,data_mid_58_imag} <<< 8);
  assign _zz_6159 = {{8{_zz_6158[23]}}, _zz_6158};
  assign _zz_6160 = fixTo_179_dout;
  assign _zz_6161 = ($signed(twiddle_factor_table_0_real) + $signed(twiddle_factor_table_0_imag));
  assign _zz_6162 = ($signed(_zz_153) - $signed(_zz_6163));
  assign _zz_6163 = ($signed(_zz_6164) * $signed(twiddle_factor_table_0_imag));
  assign _zz_6164 = ($signed(data_mid_61_real) + $signed(data_mid_61_imag));
  assign _zz_6165 = fixTo_180_dout;
  assign _zz_6166 = ($signed(_zz_153) + $signed(_zz_6167));
  assign _zz_6167 = ($signed(_zz_6168) * $signed(twiddle_factor_table_0_real));
  assign _zz_6168 = ($signed(data_mid_61_imag) - $signed(data_mid_61_real));
  assign _zz_6169 = fixTo_181_dout;
  assign _zz_6170 = _zz_6171[31 : 0];
  assign _zz_6171 = _zz_6172;
  assign _zz_6172 = ($signed(_zz_6173) >>> _zz_154);
  assign _zz_6173 = _zz_6174;
  assign _zz_6174 = ($signed(_zz_6176) - $signed(_zz_151));
  assign _zz_6175 = ({8'd0,data_mid_60_real} <<< 8);
  assign _zz_6176 = {{8{_zz_6175[23]}}, _zz_6175};
  assign _zz_6177 = fixTo_182_dout;
  assign _zz_6178 = _zz_6179[31 : 0];
  assign _zz_6179 = _zz_6180;
  assign _zz_6180 = ($signed(_zz_6181) >>> _zz_154);
  assign _zz_6181 = _zz_6182;
  assign _zz_6182 = ($signed(_zz_6184) - $signed(_zz_152));
  assign _zz_6183 = ({8'd0,data_mid_60_imag} <<< 8);
  assign _zz_6184 = {{8{_zz_6183[23]}}, _zz_6183};
  assign _zz_6185 = fixTo_183_dout;
  assign _zz_6186 = _zz_6187[31 : 0];
  assign _zz_6187 = _zz_6188;
  assign _zz_6188 = ($signed(_zz_6189) >>> _zz_155);
  assign _zz_6189 = _zz_6190;
  assign _zz_6190 = ($signed(_zz_6192) + $signed(_zz_151));
  assign _zz_6191 = ({8'd0,data_mid_60_real} <<< 8);
  assign _zz_6192 = {{8{_zz_6191[23]}}, _zz_6191};
  assign _zz_6193 = fixTo_184_dout;
  assign _zz_6194 = _zz_6195[31 : 0];
  assign _zz_6195 = _zz_6196;
  assign _zz_6196 = ($signed(_zz_6197) >>> _zz_155);
  assign _zz_6197 = _zz_6198;
  assign _zz_6198 = ($signed(_zz_6200) + $signed(_zz_152));
  assign _zz_6199 = ({8'd0,data_mid_60_imag} <<< 8);
  assign _zz_6200 = {{8{_zz_6199[23]}}, _zz_6199};
  assign _zz_6201 = fixTo_185_dout;
  assign _zz_6202 = ($signed(twiddle_factor_table_0_real) + $signed(twiddle_factor_table_0_imag));
  assign _zz_6203 = ($signed(_zz_158) - $signed(_zz_6204));
  assign _zz_6204 = ($signed(_zz_6205) * $signed(twiddle_factor_table_0_imag));
  assign _zz_6205 = ($signed(data_mid_63_real) + $signed(data_mid_63_imag));
  assign _zz_6206 = fixTo_186_dout;
  assign _zz_6207 = ($signed(_zz_158) + $signed(_zz_6208));
  assign _zz_6208 = ($signed(_zz_6209) * $signed(twiddle_factor_table_0_real));
  assign _zz_6209 = ($signed(data_mid_63_imag) - $signed(data_mid_63_real));
  assign _zz_6210 = fixTo_187_dout;
  assign _zz_6211 = _zz_6212[31 : 0];
  assign _zz_6212 = _zz_6213;
  assign _zz_6213 = ($signed(_zz_6214) >>> _zz_159);
  assign _zz_6214 = _zz_6215;
  assign _zz_6215 = ($signed(_zz_6217) - $signed(_zz_156));
  assign _zz_6216 = ({8'd0,data_mid_62_real} <<< 8);
  assign _zz_6217 = {{8{_zz_6216[23]}}, _zz_6216};
  assign _zz_6218 = fixTo_188_dout;
  assign _zz_6219 = _zz_6220[31 : 0];
  assign _zz_6220 = _zz_6221;
  assign _zz_6221 = ($signed(_zz_6222) >>> _zz_159);
  assign _zz_6222 = _zz_6223;
  assign _zz_6223 = ($signed(_zz_6225) - $signed(_zz_157));
  assign _zz_6224 = ({8'd0,data_mid_62_imag} <<< 8);
  assign _zz_6225 = {{8{_zz_6224[23]}}, _zz_6224};
  assign _zz_6226 = fixTo_189_dout;
  assign _zz_6227 = _zz_6228[31 : 0];
  assign _zz_6228 = _zz_6229;
  assign _zz_6229 = ($signed(_zz_6230) >>> _zz_160);
  assign _zz_6230 = _zz_6231;
  assign _zz_6231 = ($signed(_zz_6233) + $signed(_zz_156));
  assign _zz_6232 = ({8'd0,data_mid_62_real} <<< 8);
  assign _zz_6233 = {{8{_zz_6232[23]}}, _zz_6232};
  assign _zz_6234 = fixTo_190_dout;
  assign _zz_6235 = _zz_6236[31 : 0];
  assign _zz_6236 = _zz_6237;
  assign _zz_6237 = ($signed(_zz_6238) >>> _zz_160);
  assign _zz_6238 = _zz_6239;
  assign _zz_6239 = ($signed(_zz_6241) + $signed(_zz_157));
  assign _zz_6240 = ({8'd0,data_mid_62_imag} <<< 8);
  assign _zz_6241 = {{8{_zz_6240[23]}}, _zz_6240};
  assign _zz_6242 = fixTo_191_dout;
  assign _zz_6243 = ($signed(twiddle_factor_table_0_real) + $signed(twiddle_factor_table_0_imag));
  assign _zz_6244 = ($signed(_zz_163) - $signed(_zz_6245));
  assign _zz_6245 = ($signed(_zz_6246) * $signed(twiddle_factor_table_0_imag));
  assign _zz_6246 = ($signed(data_mid_65_real) + $signed(data_mid_65_imag));
  assign _zz_6247 = fixTo_192_dout;
  assign _zz_6248 = ($signed(_zz_163) + $signed(_zz_6249));
  assign _zz_6249 = ($signed(_zz_6250) * $signed(twiddle_factor_table_0_real));
  assign _zz_6250 = ($signed(data_mid_65_imag) - $signed(data_mid_65_real));
  assign _zz_6251 = fixTo_193_dout;
  assign _zz_6252 = _zz_6253[31 : 0];
  assign _zz_6253 = _zz_6254;
  assign _zz_6254 = ($signed(_zz_6255) >>> _zz_164);
  assign _zz_6255 = _zz_6256;
  assign _zz_6256 = ($signed(_zz_6258) - $signed(_zz_161));
  assign _zz_6257 = ({8'd0,data_mid_64_real} <<< 8);
  assign _zz_6258 = {{8{_zz_6257[23]}}, _zz_6257};
  assign _zz_6259 = fixTo_194_dout;
  assign _zz_6260 = _zz_6261[31 : 0];
  assign _zz_6261 = _zz_6262;
  assign _zz_6262 = ($signed(_zz_6263) >>> _zz_164);
  assign _zz_6263 = _zz_6264;
  assign _zz_6264 = ($signed(_zz_6266) - $signed(_zz_162));
  assign _zz_6265 = ({8'd0,data_mid_64_imag} <<< 8);
  assign _zz_6266 = {{8{_zz_6265[23]}}, _zz_6265};
  assign _zz_6267 = fixTo_195_dout;
  assign _zz_6268 = _zz_6269[31 : 0];
  assign _zz_6269 = _zz_6270;
  assign _zz_6270 = ($signed(_zz_6271) >>> _zz_165);
  assign _zz_6271 = _zz_6272;
  assign _zz_6272 = ($signed(_zz_6274) + $signed(_zz_161));
  assign _zz_6273 = ({8'd0,data_mid_64_real} <<< 8);
  assign _zz_6274 = {{8{_zz_6273[23]}}, _zz_6273};
  assign _zz_6275 = fixTo_196_dout;
  assign _zz_6276 = _zz_6277[31 : 0];
  assign _zz_6277 = _zz_6278;
  assign _zz_6278 = ($signed(_zz_6279) >>> _zz_165);
  assign _zz_6279 = _zz_6280;
  assign _zz_6280 = ($signed(_zz_6282) + $signed(_zz_162));
  assign _zz_6281 = ({8'd0,data_mid_64_imag} <<< 8);
  assign _zz_6282 = {{8{_zz_6281[23]}}, _zz_6281};
  assign _zz_6283 = fixTo_197_dout;
  assign _zz_6284 = ($signed(twiddle_factor_table_0_real) + $signed(twiddle_factor_table_0_imag));
  assign _zz_6285 = ($signed(_zz_168) - $signed(_zz_6286));
  assign _zz_6286 = ($signed(_zz_6287) * $signed(twiddle_factor_table_0_imag));
  assign _zz_6287 = ($signed(data_mid_67_real) + $signed(data_mid_67_imag));
  assign _zz_6288 = fixTo_198_dout;
  assign _zz_6289 = ($signed(_zz_168) + $signed(_zz_6290));
  assign _zz_6290 = ($signed(_zz_6291) * $signed(twiddle_factor_table_0_real));
  assign _zz_6291 = ($signed(data_mid_67_imag) - $signed(data_mid_67_real));
  assign _zz_6292 = fixTo_199_dout;
  assign _zz_6293 = _zz_6294[31 : 0];
  assign _zz_6294 = _zz_6295;
  assign _zz_6295 = ($signed(_zz_6296) >>> _zz_169);
  assign _zz_6296 = _zz_6297;
  assign _zz_6297 = ($signed(_zz_6299) - $signed(_zz_166));
  assign _zz_6298 = ({8'd0,data_mid_66_real} <<< 8);
  assign _zz_6299 = {{8{_zz_6298[23]}}, _zz_6298};
  assign _zz_6300 = fixTo_200_dout;
  assign _zz_6301 = _zz_6302[31 : 0];
  assign _zz_6302 = _zz_6303;
  assign _zz_6303 = ($signed(_zz_6304) >>> _zz_169);
  assign _zz_6304 = _zz_6305;
  assign _zz_6305 = ($signed(_zz_6307) - $signed(_zz_167));
  assign _zz_6306 = ({8'd0,data_mid_66_imag} <<< 8);
  assign _zz_6307 = {{8{_zz_6306[23]}}, _zz_6306};
  assign _zz_6308 = fixTo_201_dout;
  assign _zz_6309 = _zz_6310[31 : 0];
  assign _zz_6310 = _zz_6311;
  assign _zz_6311 = ($signed(_zz_6312) >>> _zz_170);
  assign _zz_6312 = _zz_6313;
  assign _zz_6313 = ($signed(_zz_6315) + $signed(_zz_166));
  assign _zz_6314 = ({8'd0,data_mid_66_real} <<< 8);
  assign _zz_6315 = {{8{_zz_6314[23]}}, _zz_6314};
  assign _zz_6316 = fixTo_202_dout;
  assign _zz_6317 = _zz_6318[31 : 0];
  assign _zz_6318 = _zz_6319;
  assign _zz_6319 = ($signed(_zz_6320) >>> _zz_170);
  assign _zz_6320 = _zz_6321;
  assign _zz_6321 = ($signed(_zz_6323) + $signed(_zz_167));
  assign _zz_6322 = ({8'd0,data_mid_66_imag} <<< 8);
  assign _zz_6323 = {{8{_zz_6322[23]}}, _zz_6322};
  assign _zz_6324 = fixTo_203_dout;
  assign _zz_6325 = ($signed(twiddle_factor_table_0_real) + $signed(twiddle_factor_table_0_imag));
  assign _zz_6326 = ($signed(_zz_173) - $signed(_zz_6327));
  assign _zz_6327 = ($signed(_zz_6328) * $signed(twiddle_factor_table_0_imag));
  assign _zz_6328 = ($signed(data_mid_69_real) + $signed(data_mid_69_imag));
  assign _zz_6329 = fixTo_204_dout;
  assign _zz_6330 = ($signed(_zz_173) + $signed(_zz_6331));
  assign _zz_6331 = ($signed(_zz_6332) * $signed(twiddle_factor_table_0_real));
  assign _zz_6332 = ($signed(data_mid_69_imag) - $signed(data_mid_69_real));
  assign _zz_6333 = fixTo_205_dout;
  assign _zz_6334 = _zz_6335[31 : 0];
  assign _zz_6335 = _zz_6336;
  assign _zz_6336 = ($signed(_zz_6337) >>> _zz_174);
  assign _zz_6337 = _zz_6338;
  assign _zz_6338 = ($signed(_zz_6340) - $signed(_zz_171));
  assign _zz_6339 = ({8'd0,data_mid_68_real} <<< 8);
  assign _zz_6340 = {{8{_zz_6339[23]}}, _zz_6339};
  assign _zz_6341 = fixTo_206_dout;
  assign _zz_6342 = _zz_6343[31 : 0];
  assign _zz_6343 = _zz_6344;
  assign _zz_6344 = ($signed(_zz_6345) >>> _zz_174);
  assign _zz_6345 = _zz_6346;
  assign _zz_6346 = ($signed(_zz_6348) - $signed(_zz_172));
  assign _zz_6347 = ({8'd0,data_mid_68_imag} <<< 8);
  assign _zz_6348 = {{8{_zz_6347[23]}}, _zz_6347};
  assign _zz_6349 = fixTo_207_dout;
  assign _zz_6350 = _zz_6351[31 : 0];
  assign _zz_6351 = _zz_6352;
  assign _zz_6352 = ($signed(_zz_6353) >>> _zz_175);
  assign _zz_6353 = _zz_6354;
  assign _zz_6354 = ($signed(_zz_6356) + $signed(_zz_171));
  assign _zz_6355 = ({8'd0,data_mid_68_real} <<< 8);
  assign _zz_6356 = {{8{_zz_6355[23]}}, _zz_6355};
  assign _zz_6357 = fixTo_208_dout;
  assign _zz_6358 = _zz_6359[31 : 0];
  assign _zz_6359 = _zz_6360;
  assign _zz_6360 = ($signed(_zz_6361) >>> _zz_175);
  assign _zz_6361 = _zz_6362;
  assign _zz_6362 = ($signed(_zz_6364) + $signed(_zz_172));
  assign _zz_6363 = ({8'd0,data_mid_68_imag} <<< 8);
  assign _zz_6364 = {{8{_zz_6363[23]}}, _zz_6363};
  assign _zz_6365 = fixTo_209_dout;
  assign _zz_6366 = ($signed(twiddle_factor_table_0_real) + $signed(twiddle_factor_table_0_imag));
  assign _zz_6367 = ($signed(_zz_178) - $signed(_zz_6368));
  assign _zz_6368 = ($signed(_zz_6369) * $signed(twiddle_factor_table_0_imag));
  assign _zz_6369 = ($signed(data_mid_71_real) + $signed(data_mid_71_imag));
  assign _zz_6370 = fixTo_210_dout;
  assign _zz_6371 = ($signed(_zz_178) + $signed(_zz_6372));
  assign _zz_6372 = ($signed(_zz_6373) * $signed(twiddle_factor_table_0_real));
  assign _zz_6373 = ($signed(data_mid_71_imag) - $signed(data_mid_71_real));
  assign _zz_6374 = fixTo_211_dout;
  assign _zz_6375 = _zz_6376[31 : 0];
  assign _zz_6376 = _zz_6377;
  assign _zz_6377 = ($signed(_zz_6378) >>> _zz_179);
  assign _zz_6378 = _zz_6379;
  assign _zz_6379 = ($signed(_zz_6381) - $signed(_zz_176));
  assign _zz_6380 = ({8'd0,data_mid_70_real} <<< 8);
  assign _zz_6381 = {{8{_zz_6380[23]}}, _zz_6380};
  assign _zz_6382 = fixTo_212_dout;
  assign _zz_6383 = _zz_6384[31 : 0];
  assign _zz_6384 = _zz_6385;
  assign _zz_6385 = ($signed(_zz_6386) >>> _zz_179);
  assign _zz_6386 = _zz_6387;
  assign _zz_6387 = ($signed(_zz_6389) - $signed(_zz_177));
  assign _zz_6388 = ({8'd0,data_mid_70_imag} <<< 8);
  assign _zz_6389 = {{8{_zz_6388[23]}}, _zz_6388};
  assign _zz_6390 = fixTo_213_dout;
  assign _zz_6391 = _zz_6392[31 : 0];
  assign _zz_6392 = _zz_6393;
  assign _zz_6393 = ($signed(_zz_6394) >>> _zz_180);
  assign _zz_6394 = _zz_6395;
  assign _zz_6395 = ($signed(_zz_6397) + $signed(_zz_176));
  assign _zz_6396 = ({8'd0,data_mid_70_real} <<< 8);
  assign _zz_6397 = {{8{_zz_6396[23]}}, _zz_6396};
  assign _zz_6398 = fixTo_214_dout;
  assign _zz_6399 = _zz_6400[31 : 0];
  assign _zz_6400 = _zz_6401;
  assign _zz_6401 = ($signed(_zz_6402) >>> _zz_180);
  assign _zz_6402 = _zz_6403;
  assign _zz_6403 = ($signed(_zz_6405) + $signed(_zz_177));
  assign _zz_6404 = ({8'd0,data_mid_70_imag} <<< 8);
  assign _zz_6405 = {{8{_zz_6404[23]}}, _zz_6404};
  assign _zz_6406 = fixTo_215_dout;
  assign _zz_6407 = ($signed(twiddle_factor_table_0_real) + $signed(twiddle_factor_table_0_imag));
  assign _zz_6408 = ($signed(_zz_183) - $signed(_zz_6409));
  assign _zz_6409 = ($signed(_zz_6410) * $signed(twiddle_factor_table_0_imag));
  assign _zz_6410 = ($signed(data_mid_73_real) + $signed(data_mid_73_imag));
  assign _zz_6411 = fixTo_216_dout;
  assign _zz_6412 = ($signed(_zz_183) + $signed(_zz_6413));
  assign _zz_6413 = ($signed(_zz_6414) * $signed(twiddle_factor_table_0_real));
  assign _zz_6414 = ($signed(data_mid_73_imag) - $signed(data_mid_73_real));
  assign _zz_6415 = fixTo_217_dout;
  assign _zz_6416 = _zz_6417[31 : 0];
  assign _zz_6417 = _zz_6418;
  assign _zz_6418 = ($signed(_zz_6419) >>> _zz_184);
  assign _zz_6419 = _zz_6420;
  assign _zz_6420 = ($signed(_zz_6422) - $signed(_zz_181));
  assign _zz_6421 = ({8'd0,data_mid_72_real} <<< 8);
  assign _zz_6422 = {{8{_zz_6421[23]}}, _zz_6421};
  assign _zz_6423 = fixTo_218_dout;
  assign _zz_6424 = _zz_6425[31 : 0];
  assign _zz_6425 = _zz_6426;
  assign _zz_6426 = ($signed(_zz_6427) >>> _zz_184);
  assign _zz_6427 = _zz_6428;
  assign _zz_6428 = ($signed(_zz_6430) - $signed(_zz_182));
  assign _zz_6429 = ({8'd0,data_mid_72_imag} <<< 8);
  assign _zz_6430 = {{8{_zz_6429[23]}}, _zz_6429};
  assign _zz_6431 = fixTo_219_dout;
  assign _zz_6432 = _zz_6433[31 : 0];
  assign _zz_6433 = _zz_6434;
  assign _zz_6434 = ($signed(_zz_6435) >>> _zz_185);
  assign _zz_6435 = _zz_6436;
  assign _zz_6436 = ($signed(_zz_6438) + $signed(_zz_181));
  assign _zz_6437 = ({8'd0,data_mid_72_real} <<< 8);
  assign _zz_6438 = {{8{_zz_6437[23]}}, _zz_6437};
  assign _zz_6439 = fixTo_220_dout;
  assign _zz_6440 = _zz_6441[31 : 0];
  assign _zz_6441 = _zz_6442;
  assign _zz_6442 = ($signed(_zz_6443) >>> _zz_185);
  assign _zz_6443 = _zz_6444;
  assign _zz_6444 = ($signed(_zz_6446) + $signed(_zz_182));
  assign _zz_6445 = ({8'd0,data_mid_72_imag} <<< 8);
  assign _zz_6446 = {{8{_zz_6445[23]}}, _zz_6445};
  assign _zz_6447 = fixTo_221_dout;
  assign _zz_6448 = ($signed(twiddle_factor_table_0_real) + $signed(twiddle_factor_table_0_imag));
  assign _zz_6449 = ($signed(_zz_188) - $signed(_zz_6450));
  assign _zz_6450 = ($signed(_zz_6451) * $signed(twiddle_factor_table_0_imag));
  assign _zz_6451 = ($signed(data_mid_75_real) + $signed(data_mid_75_imag));
  assign _zz_6452 = fixTo_222_dout;
  assign _zz_6453 = ($signed(_zz_188) + $signed(_zz_6454));
  assign _zz_6454 = ($signed(_zz_6455) * $signed(twiddle_factor_table_0_real));
  assign _zz_6455 = ($signed(data_mid_75_imag) - $signed(data_mid_75_real));
  assign _zz_6456 = fixTo_223_dout;
  assign _zz_6457 = _zz_6458[31 : 0];
  assign _zz_6458 = _zz_6459;
  assign _zz_6459 = ($signed(_zz_6460) >>> _zz_189);
  assign _zz_6460 = _zz_6461;
  assign _zz_6461 = ($signed(_zz_6463) - $signed(_zz_186));
  assign _zz_6462 = ({8'd0,data_mid_74_real} <<< 8);
  assign _zz_6463 = {{8{_zz_6462[23]}}, _zz_6462};
  assign _zz_6464 = fixTo_224_dout;
  assign _zz_6465 = _zz_6466[31 : 0];
  assign _zz_6466 = _zz_6467;
  assign _zz_6467 = ($signed(_zz_6468) >>> _zz_189);
  assign _zz_6468 = _zz_6469;
  assign _zz_6469 = ($signed(_zz_6471) - $signed(_zz_187));
  assign _zz_6470 = ({8'd0,data_mid_74_imag} <<< 8);
  assign _zz_6471 = {{8{_zz_6470[23]}}, _zz_6470};
  assign _zz_6472 = fixTo_225_dout;
  assign _zz_6473 = _zz_6474[31 : 0];
  assign _zz_6474 = _zz_6475;
  assign _zz_6475 = ($signed(_zz_6476) >>> _zz_190);
  assign _zz_6476 = _zz_6477;
  assign _zz_6477 = ($signed(_zz_6479) + $signed(_zz_186));
  assign _zz_6478 = ({8'd0,data_mid_74_real} <<< 8);
  assign _zz_6479 = {{8{_zz_6478[23]}}, _zz_6478};
  assign _zz_6480 = fixTo_226_dout;
  assign _zz_6481 = _zz_6482[31 : 0];
  assign _zz_6482 = _zz_6483;
  assign _zz_6483 = ($signed(_zz_6484) >>> _zz_190);
  assign _zz_6484 = _zz_6485;
  assign _zz_6485 = ($signed(_zz_6487) + $signed(_zz_187));
  assign _zz_6486 = ({8'd0,data_mid_74_imag} <<< 8);
  assign _zz_6487 = {{8{_zz_6486[23]}}, _zz_6486};
  assign _zz_6488 = fixTo_227_dout;
  assign _zz_6489 = ($signed(twiddle_factor_table_0_real) + $signed(twiddle_factor_table_0_imag));
  assign _zz_6490 = ($signed(_zz_193) - $signed(_zz_6491));
  assign _zz_6491 = ($signed(_zz_6492) * $signed(twiddle_factor_table_0_imag));
  assign _zz_6492 = ($signed(data_mid_77_real) + $signed(data_mid_77_imag));
  assign _zz_6493 = fixTo_228_dout;
  assign _zz_6494 = ($signed(_zz_193) + $signed(_zz_6495));
  assign _zz_6495 = ($signed(_zz_6496) * $signed(twiddle_factor_table_0_real));
  assign _zz_6496 = ($signed(data_mid_77_imag) - $signed(data_mid_77_real));
  assign _zz_6497 = fixTo_229_dout;
  assign _zz_6498 = _zz_6499[31 : 0];
  assign _zz_6499 = _zz_6500;
  assign _zz_6500 = ($signed(_zz_6501) >>> _zz_194);
  assign _zz_6501 = _zz_6502;
  assign _zz_6502 = ($signed(_zz_6504) - $signed(_zz_191));
  assign _zz_6503 = ({8'd0,data_mid_76_real} <<< 8);
  assign _zz_6504 = {{8{_zz_6503[23]}}, _zz_6503};
  assign _zz_6505 = fixTo_230_dout;
  assign _zz_6506 = _zz_6507[31 : 0];
  assign _zz_6507 = _zz_6508;
  assign _zz_6508 = ($signed(_zz_6509) >>> _zz_194);
  assign _zz_6509 = _zz_6510;
  assign _zz_6510 = ($signed(_zz_6512) - $signed(_zz_192));
  assign _zz_6511 = ({8'd0,data_mid_76_imag} <<< 8);
  assign _zz_6512 = {{8{_zz_6511[23]}}, _zz_6511};
  assign _zz_6513 = fixTo_231_dout;
  assign _zz_6514 = _zz_6515[31 : 0];
  assign _zz_6515 = _zz_6516;
  assign _zz_6516 = ($signed(_zz_6517) >>> _zz_195);
  assign _zz_6517 = _zz_6518;
  assign _zz_6518 = ($signed(_zz_6520) + $signed(_zz_191));
  assign _zz_6519 = ({8'd0,data_mid_76_real} <<< 8);
  assign _zz_6520 = {{8{_zz_6519[23]}}, _zz_6519};
  assign _zz_6521 = fixTo_232_dout;
  assign _zz_6522 = _zz_6523[31 : 0];
  assign _zz_6523 = _zz_6524;
  assign _zz_6524 = ($signed(_zz_6525) >>> _zz_195);
  assign _zz_6525 = _zz_6526;
  assign _zz_6526 = ($signed(_zz_6528) + $signed(_zz_192));
  assign _zz_6527 = ({8'd0,data_mid_76_imag} <<< 8);
  assign _zz_6528 = {{8{_zz_6527[23]}}, _zz_6527};
  assign _zz_6529 = fixTo_233_dout;
  assign _zz_6530 = ($signed(twiddle_factor_table_0_real) + $signed(twiddle_factor_table_0_imag));
  assign _zz_6531 = ($signed(_zz_198) - $signed(_zz_6532));
  assign _zz_6532 = ($signed(_zz_6533) * $signed(twiddle_factor_table_0_imag));
  assign _zz_6533 = ($signed(data_mid_79_real) + $signed(data_mid_79_imag));
  assign _zz_6534 = fixTo_234_dout;
  assign _zz_6535 = ($signed(_zz_198) + $signed(_zz_6536));
  assign _zz_6536 = ($signed(_zz_6537) * $signed(twiddle_factor_table_0_real));
  assign _zz_6537 = ($signed(data_mid_79_imag) - $signed(data_mid_79_real));
  assign _zz_6538 = fixTo_235_dout;
  assign _zz_6539 = _zz_6540[31 : 0];
  assign _zz_6540 = _zz_6541;
  assign _zz_6541 = ($signed(_zz_6542) >>> _zz_199);
  assign _zz_6542 = _zz_6543;
  assign _zz_6543 = ($signed(_zz_6545) - $signed(_zz_196));
  assign _zz_6544 = ({8'd0,data_mid_78_real} <<< 8);
  assign _zz_6545 = {{8{_zz_6544[23]}}, _zz_6544};
  assign _zz_6546 = fixTo_236_dout;
  assign _zz_6547 = _zz_6548[31 : 0];
  assign _zz_6548 = _zz_6549;
  assign _zz_6549 = ($signed(_zz_6550) >>> _zz_199);
  assign _zz_6550 = _zz_6551;
  assign _zz_6551 = ($signed(_zz_6553) - $signed(_zz_197));
  assign _zz_6552 = ({8'd0,data_mid_78_imag} <<< 8);
  assign _zz_6553 = {{8{_zz_6552[23]}}, _zz_6552};
  assign _zz_6554 = fixTo_237_dout;
  assign _zz_6555 = _zz_6556[31 : 0];
  assign _zz_6556 = _zz_6557;
  assign _zz_6557 = ($signed(_zz_6558) >>> _zz_200);
  assign _zz_6558 = _zz_6559;
  assign _zz_6559 = ($signed(_zz_6561) + $signed(_zz_196));
  assign _zz_6560 = ({8'd0,data_mid_78_real} <<< 8);
  assign _zz_6561 = {{8{_zz_6560[23]}}, _zz_6560};
  assign _zz_6562 = fixTo_238_dout;
  assign _zz_6563 = _zz_6564[31 : 0];
  assign _zz_6564 = _zz_6565;
  assign _zz_6565 = ($signed(_zz_6566) >>> _zz_200);
  assign _zz_6566 = _zz_6567;
  assign _zz_6567 = ($signed(_zz_6569) + $signed(_zz_197));
  assign _zz_6568 = ({8'd0,data_mid_78_imag} <<< 8);
  assign _zz_6569 = {{8{_zz_6568[23]}}, _zz_6568};
  assign _zz_6570 = fixTo_239_dout;
  assign _zz_6571 = ($signed(twiddle_factor_table_0_real) + $signed(twiddle_factor_table_0_imag));
  assign _zz_6572 = ($signed(_zz_203) - $signed(_zz_6573));
  assign _zz_6573 = ($signed(_zz_6574) * $signed(twiddle_factor_table_0_imag));
  assign _zz_6574 = ($signed(data_mid_81_real) + $signed(data_mid_81_imag));
  assign _zz_6575 = fixTo_240_dout;
  assign _zz_6576 = ($signed(_zz_203) + $signed(_zz_6577));
  assign _zz_6577 = ($signed(_zz_6578) * $signed(twiddle_factor_table_0_real));
  assign _zz_6578 = ($signed(data_mid_81_imag) - $signed(data_mid_81_real));
  assign _zz_6579 = fixTo_241_dout;
  assign _zz_6580 = _zz_6581[31 : 0];
  assign _zz_6581 = _zz_6582;
  assign _zz_6582 = ($signed(_zz_6583) >>> _zz_204);
  assign _zz_6583 = _zz_6584;
  assign _zz_6584 = ($signed(_zz_6586) - $signed(_zz_201));
  assign _zz_6585 = ({8'd0,data_mid_80_real} <<< 8);
  assign _zz_6586 = {{8{_zz_6585[23]}}, _zz_6585};
  assign _zz_6587 = fixTo_242_dout;
  assign _zz_6588 = _zz_6589[31 : 0];
  assign _zz_6589 = _zz_6590;
  assign _zz_6590 = ($signed(_zz_6591) >>> _zz_204);
  assign _zz_6591 = _zz_6592;
  assign _zz_6592 = ($signed(_zz_6594) - $signed(_zz_202));
  assign _zz_6593 = ({8'd0,data_mid_80_imag} <<< 8);
  assign _zz_6594 = {{8{_zz_6593[23]}}, _zz_6593};
  assign _zz_6595 = fixTo_243_dout;
  assign _zz_6596 = _zz_6597[31 : 0];
  assign _zz_6597 = _zz_6598;
  assign _zz_6598 = ($signed(_zz_6599) >>> _zz_205);
  assign _zz_6599 = _zz_6600;
  assign _zz_6600 = ($signed(_zz_6602) + $signed(_zz_201));
  assign _zz_6601 = ({8'd0,data_mid_80_real} <<< 8);
  assign _zz_6602 = {{8{_zz_6601[23]}}, _zz_6601};
  assign _zz_6603 = fixTo_244_dout;
  assign _zz_6604 = _zz_6605[31 : 0];
  assign _zz_6605 = _zz_6606;
  assign _zz_6606 = ($signed(_zz_6607) >>> _zz_205);
  assign _zz_6607 = _zz_6608;
  assign _zz_6608 = ($signed(_zz_6610) + $signed(_zz_202));
  assign _zz_6609 = ({8'd0,data_mid_80_imag} <<< 8);
  assign _zz_6610 = {{8{_zz_6609[23]}}, _zz_6609};
  assign _zz_6611 = fixTo_245_dout;
  assign _zz_6612 = ($signed(twiddle_factor_table_0_real) + $signed(twiddle_factor_table_0_imag));
  assign _zz_6613 = ($signed(_zz_208) - $signed(_zz_6614));
  assign _zz_6614 = ($signed(_zz_6615) * $signed(twiddle_factor_table_0_imag));
  assign _zz_6615 = ($signed(data_mid_83_real) + $signed(data_mid_83_imag));
  assign _zz_6616 = fixTo_246_dout;
  assign _zz_6617 = ($signed(_zz_208) + $signed(_zz_6618));
  assign _zz_6618 = ($signed(_zz_6619) * $signed(twiddle_factor_table_0_real));
  assign _zz_6619 = ($signed(data_mid_83_imag) - $signed(data_mid_83_real));
  assign _zz_6620 = fixTo_247_dout;
  assign _zz_6621 = _zz_6622[31 : 0];
  assign _zz_6622 = _zz_6623;
  assign _zz_6623 = ($signed(_zz_6624) >>> _zz_209);
  assign _zz_6624 = _zz_6625;
  assign _zz_6625 = ($signed(_zz_6627) - $signed(_zz_206));
  assign _zz_6626 = ({8'd0,data_mid_82_real} <<< 8);
  assign _zz_6627 = {{8{_zz_6626[23]}}, _zz_6626};
  assign _zz_6628 = fixTo_248_dout;
  assign _zz_6629 = _zz_6630[31 : 0];
  assign _zz_6630 = _zz_6631;
  assign _zz_6631 = ($signed(_zz_6632) >>> _zz_209);
  assign _zz_6632 = _zz_6633;
  assign _zz_6633 = ($signed(_zz_6635) - $signed(_zz_207));
  assign _zz_6634 = ({8'd0,data_mid_82_imag} <<< 8);
  assign _zz_6635 = {{8{_zz_6634[23]}}, _zz_6634};
  assign _zz_6636 = fixTo_249_dout;
  assign _zz_6637 = _zz_6638[31 : 0];
  assign _zz_6638 = _zz_6639;
  assign _zz_6639 = ($signed(_zz_6640) >>> _zz_210);
  assign _zz_6640 = _zz_6641;
  assign _zz_6641 = ($signed(_zz_6643) + $signed(_zz_206));
  assign _zz_6642 = ({8'd0,data_mid_82_real} <<< 8);
  assign _zz_6643 = {{8{_zz_6642[23]}}, _zz_6642};
  assign _zz_6644 = fixTo_250_dout;
  assign _zz_6645 = _zz_6646[31 : 0];
  assign _zz_6646 = _zz_6647;
  assign _zz_6647 = ($signed(_zz_6648) >>> _zz_210);
  assign _zz_6648 = _zz_6649;
  assign _zz_6649 = ($signed(_zz_6651) + $signed(_zz_207));
  assign _zz_6650 = ({8'd0,data_mid_82_imag} <<< 8);
  assign _zz_6651 = {{8{_zz_6650[23]}}, _zz_6650};
  assign _zz_6652 = fixTo_251_dout;
  assign _zz_6653 = ($signed(twiddle_factor_table_0_real) + $signed(twiddle_factor_table_0_imag));
  assign _zz_6654 = ($signed(_zz_213) - $signed(_zz_6655));
  assign _zz_6655 = ($signed(_zz_6656) * $signed(twiddle_factor_table_0_imag));
  assign _zz_6656 = ($signed(data_mid_85_real) + $signed(data_mid_85_imag));
  assign _zz_6657 = fixTo_252_dout;
  assign _zz_6658 = ($signed(_zz_213) + $signed(_zz_6659));
  assign _zz_6659 = ($signed(_zz_6660) * $signed(twiddle_factor_table_0_real));
  assign _zz_6660 = ($signed(data_mid_85_imag) - $signed(data_mid_85_real));
  assign _zz_6661 = fixTo_253_dout;
  assign _zz_6662 = _zz_6663[31 : 0];
  assign _zz_6663 = _zz_6664;
  assign _zz_6664 = ($signed(_zz_6665) >>> _zz_214);
  assign _zz_6665 = _zz_6666;
  assign _zz_6666 = ($signed(_zz_6668) - $signed(_zz_211));
  assign _zz_6667 = ({8'd0,data_mid_84_real} <<< 8);
  assign _zz_6668 = {{8{_zz_6667[23]}}, _zz_6667};
  assign _zz_6669 = fixTo_254_dout;
  assign _zz_6670 = _zz_6671[31 : 0];
  assign _zz_6671 = _zz_6672;
  assign _zz_6672 = ($signed(_zz_6673) >>> _zz_214);
  assign _zz_6673 = _zz_6674;
  assign _zz_6674 = ($signed(_zz_6676) - $signed(_zz_212));
  assign _zz_6675 = ({8'd0,data_mid_84_imag} <<< 8);
  assign _zz_6676 = {{8{_zz_6675[23]}}, _zz_6675};
  assign _zz_6677 = fixTo_255_dout;
  assign _zz_6678 = _zz_6679[31 : 0];
  assign _zz_6679 = _zz_6680;
  assign _zz_6680 = ($signed(_zz_6681) >>> _zz_215);
  assign _zz_6681 = _zz_6682;
  assign _zz_6682 = ($signed(_zz_6684) + $signed(_zz_211));
  assign _zz_6683 = ({8'd0,data_mid_84_real} <<< 8);
  assign _zz_6684 = {{8{_zz_6683[23]}}, _zz_6683};
  assign _zz_6685 = fixTo_256_dout;
  assign _zz_6686 = _zz_6687[31 : 0];
  assign _zz_6687 = _zz_6688;
  assign _zz_6688 = ($signed(_zz_6689) >>> _zz_215);
  assign _zz_6689 = _zz_6690;
  assign _zz_6690 = ($signed(_zz_6692) + $signed(_zz_212));
  assign _zz_6691 = ({8'd0,data_mid_84_imag} <<< 8);
  assign _zz_6692 = {{8{_zz_6691[23]}}, _zz_6691};
  assign _zz_6693 = fixTo_257_dout;
  assign _zz_6694 = ($signed(twiddle_factor_table_0_real) + $signed(twiddle_factor_table_0_imag));
  assign _zz_6695 = ($signed(_zz_218) - $signed(_zz_6696));
  assign _zz_6696 = ($signed(_zz_6697) * $signed(twiddle_factor_table_0_imag));
  assign _zz_6697 = ($signed(data_mid_87_real) + $signed(data_mid_87_imag));
  assign _zz_6698 = fixTo_258_dout;
  assign _zz_6699 = ($signed(_zz_218) + $signed(_zz_6700));
  assign _zz_6700 = ($signed(_zz_6701) * $signed(twiddle_factor_table_0_real));
  assign _zz_6701 = ($signed(data_mid_87_imag) - $signed(data_mid_87_real));
  assign _zz_6702 = fixTo_259_dout;
  assign _zz_6703 = _zz_6704[31 : 0];
  assign _zz_6704 = _zz_6705;
  assign _zz_6705 = ($signed(_zz_6706) >>> _zz_219);
  assign _zz_6706 = _zz_6707;
  assign _zz_6707 = ($signed(_zz_6709) - $signed(_zz_216));
  assign _zz_6708 = ({8'd0,data_mid_86_real} <<< 8);
  assign _zz_6709 = {{8{_zz_6708[23]}}, _zz_6708};
  assign _zz_6710 = fixTo_260_dout;
  assign _zz_6711 = _zz_6712[31 : 0];
  assign _zz_6712 = _zz_6713;
  assign _zz_6713 = ($signed(_zz_6714) >>> _zz_219);
  assign _zz_6714 = _zz_6715;
  assign _zz_6715 = ($signed(_zz_6717) - $signed(_zz_217));
  assign _zz_6716 = ({8'd0,data_mid_86_imag} <<< 8);
  assign _zz_6717 = {{8{_zz_6716[23]}}, _zz_6716};
  assign _zz_6718 = fixTo_261_dout;
  assign _zz_6719 = _zz_6720[31 : 0];
  assign _zz_6720 = _zz_6721;
  assign _zz_6721 = ($signed(_zz_6722) >>> _zz_220);
  assign _zz_6722 = _zz_6723;
  assign _zz_6723 = ($signed(_zz_6725) + $signed(_zz_216));
  assign _zz_6724 = ({8'd0,data_mid_86_real} <<< 8);
  assign _zz_6725 = {{8{_zz_6724[23]}}, _zz_6724};
  assign _zz_6726 = fixTo_262_dout;
  assign _zz_6727 = _zz_6728[31 : 0];
  assign _zz_6728 = _zz_6729;
  assign _zz_6729 = ($signed(_zz_6730) >>> _zz_220);
  assign _zz_6730 = _zz_6731;
  assign _zz_6731 = ($signed(_zz_6733) + $signed(_zz_217));
  assign _zz_6732 = ({8'd0,data_mid_86_imag} <<< 8);
  assign _zz_6733 = {{8{_zz_6732[23]}}, _zz_6732};
  assign _zz_6734 = fixTo_263_dout;
  assign _zz_6735 = ($signed(twiddle_factor_table_0_real) + $signed(twiddle_factor_table_0_imag));
  assign _zz_6736 = ($signed(_zz_223) - $signed(_zz_6737));
  assign _zz_6737 = ($signed(_zz_6738) * $signed(twiddle_factor_table_0_imag));
  assign _zz_6738 = ($signed(data_mid_89_real) + $signed(data_mid_89_imag));
  assign _zz_6739 = fixTo_264_dout;
  assign _zz_6740 = ($signed(_zz_223) + $signed(_zz_6741));
  assign _zz_6741 = ($signed(_zz_6742) * $signed(twiddle_factor_table_0_real));
  assign _zz_6742 = ($signed(data_mid_89_imag) - $signed(data_mid_89_real));
  assign _zz_6743 = fixTo_265_dout;
  assign _zz_6744 = _zz_6745[31 : 0];
  assign _zz_6745 = _zz_6746;
  assign _zz_6746 = ($signed(_zz_6747) >>> _zz_224);
  assign _zz_6747 = _zz_6748;
  assign _zz_6748 = ($signed(_zz_6750) - $signed(_zz_221));
  assign _zz_6749 = ({8'd0,data_mid_88_real} <<< 8);
  assign _zz_6750 = {{8{_zz_6749[23]}}, _zz_6749};
  assign _zz_6751 = fixTo_266_dout;
  assign _zz_6752 = _zz_6753[31 : 0];
  assign _zz_6753 = _zz_6754;
  assign _zz_6754 = ($signed(_zz_6755) >>> _zz_224);
  assign _zz_6755 = _zz_6756;
  assign _zz_6756 = ($signed(_zz_6758) - $signed(_zz_222));
  assign _zz_6757 = ({8'd0,data_mid_88_imag} <<< 8);
  assign _zz_6758 = {{8{_zz_6757[23]}}, _zz_6757};
  assign _zz_6759 = fixTo_267_dout;
  assign _zz_6760 = _zz_6761[31 : 0];
  assign _zz_6761 = _zz_6762;
  assign _zz_6762 = ($signed(_zz_6763) >>> _zz_225);
  assign _zz_6763 = _zz_6764;
  assign _zz_6764 = ($signed(_zz_6766) + $signed(_zz_221));
  assign _zz_6765 = ({8'd0,data_mid_88_real} <<< 8);
  assign _zz_6766 = {{8{_zz_6765[23]}}, _zz_6765};
  assign _zz_6767 = fixTo_268_dout;
  assign _zz_6768 = _zz_6769[31 : 0];
  assign _zz_6769 = _zz_6770;
  assign _zz_6770 = ($signed(_zz_6771) >>> _zz_225);
  assign _zz_6771 = _zz_6772;
  assign _zz_6772 = ($signed(_zz_6774) + $signed(_zz_222));
  assign _zz_6773 = ({8'd0,data_mid_88_imag} <<< 8);
  assign _zz_6774 = {{8{_zz_6773[23]}}, _zz_6773};
  assign _zz_6775 = fixTo_269_dout;
  assign _zz_6776 = ($signed(twiddle_factor_table_0_real) + $signed(twiddle_factor_table_0_imag));
  assign _zz_6777 = ($signed(_zz_228) - $signed(_zz_6778));
  assign _zz_6778 = ($signed(_zz_6779) * $signed(twiddle_factor_table_0_imag));
  assign _zz_6779 = ($signed(data_mid_91_real) + $signed(data_mid_91_imag));
  assign _zz_6780 = fixTo_270_dout;
  assign _zz_6781 = ($signed(_zz_228) + $signed(_zz_6782));
  assign _zz_6782 = ($signed(_zz_6783) * $signed(twiddle_factor_table_0_real));
  assign _zz_6783 = ($signed(data_mid_91_imag) - $signed(data_mid_91_real));
  assign _zz_6784 = fixTo_271_dout;
  assign _zz_6785 = _zz_6786[31 : 0];
  assign _zz_6786 = _zz_6787;
  assign _zz_6787 = ($signed(_zz_6788) >>> _zz_229);
  assign _zz_6788 = _zz_6789;
  assign _zz_6789 = ($signed(_zz_6791) - $signed(_zz_226));
  assign _zz_6790 = ({8'd0,data_mid_90_real} <<< 8);
  assign _zz_6791 = {{8{_zz_6790[23]}}, _zz_6790};
  assign _zz_6792 = fixTo_272_dout;
  assign _zz_6793 = _zz_6794[31 : 0];
  assign _zz_6794 = _zz_6795;
  assign _zz_6795 = ($signed(_zz_6796) >>> _zz_229);
  assign _zz_6796 = _zz_6797;
  assign _zz_6797 = ($signed(_zz_6799) - $signed(_zz_227));
  assign _zz_6798 = ({8'd0,data_mid_90_imag} <<< 8);
  assign _zz_6799 = {{8{_zz_6798[23]}}, _zz_6798};
  assign _zz_6800 = fixTo_273_dout;
  assign _zz_6801 = _zz_6802[31 : 0];
  assign _zz_6802 = _zz_6803;
  assign _zz_6803 = ($signed(_zz_6804) >>> _zz_230);
  assign _zz_6804 = _zz_6805;
  assign _zz_6805 = ($signed(_zz_6807) + $signed(_zz_226));
  assign _zz_6806 = ({8'd0,data_mid_90_real} <<< 8);
  assign _zz_6807 = {{8{_zz_6806[23]}}, _zz_6806};
  assign _zz_6808 = fixTo_274_dout;
  assign _zz_6809 = _zz_6810[31 : 0];
  assign _zz_6810 = _zz_6811;
  assign _zz_6811 = ($signed(_zz_6812) >>> _zz_230);
  assign _zz_6812 = _zz_6813;
  assign _zz_6813 = ($signed(_zz_6815) + $signed(_zz_227));
  assign _zz_6814 = ({8'd0,data_mid_90_imag} <<< 8);
  assign _zz_6815 = {{8{_zz_6814[23]}}, _zz_6814};
  assign _zz_6816 = fixTo_275_dout;
  assign _zz_6817 = ($signed(twiddle_factor_table_0_real) + $signed(twiddle_factor_table_0_imag));
  assign _zz_6818 = ($signed(_zz_233) - $signed(_zz_6819));
  assign _zz_6819 = ($signed(_zz_6820) * $signed(twiddle_factor_table_0_imag));
  assign _zz_6820 = ($signed(data_mid_93_real) + $signed(data_mid_93_imag));
  assign _zz_6821 = fixTo_276_dout;
  assign _zz_6822 = ($signed(_zz_233) + $signed(_zz_6823));
  assign _zz_6823 = ($signed(_zz_6824) * $signed(twiddle_factor_table_0_real));
  assign _zz_6824 = ($signed(data_mid_93_imag) - $signed(data_mid_93_real));
  assign _zz_6825 = fixTo_277_dout;
  assign _zz_6826 = _zz_6827[31 : 0];
  assign _zz_6827 = _zz_6828;
  assign _zz_6828 = ($signed(_zz_6829) >>> _zz_234);
  assign _zz_6829 = _zz_6830;
  assign _zz_6830 = ($signed(_zz_6832) - $signed(_zz_231));
  assign _zz_6831 = ({8'd0,data_mid_92_real} <<< 8);
  assign _zz_6832 = {{8{_zz_6831[23]}}, _zz_6831};
  assign _zz_6833 = fixTo_278_dout;
  assign _zz_6834 = _zz_6835[31 : 0];
  assign _zz_6835 = _zz_6836;
  assign _zz_6836 = ($signed(_zz_6837) >>> _zz_234);
  assign _zz_6837 = _zz_6838;
  assign _zz_6838 = ($signed(_zz_6840) - $signed(_zz_232));
  assign _zz_6839 = ({8'd0,data_mid_92_imag} <<< 8);
  assign _zz_6840 = {{8{_zz_6839[23]}}, _zz_6839};
  assign _zz_6841 = fixTo_279_dout;
  assign _zz_6842 = _zz_6843[31 : 0];
  assign _zz_6843 = _zz_6844;
  assign _zz_6844 = ($signed(_zz_6845) >>> _zz_235);
  assign _zz_6845 = _zz_6846;
  assign _zz_6846 = ($signed(_zz_6848) + $signed(_zz_231));
  assign _zz_6847 = ({8'd0,data_mid_92_real} <<< 8);
  assign _zz_6848 = {{8{_zz_6847[23]}}, _zz_6847};
  assign _zz_6849 = fixTo_280_dout;
  assign _zz_6850 = _zz_6851[31 : 0];
  assign _zz_6851 = _zz_6852;
  assign _zz_6852 = ($signed(_zz_6853) >>> _zz_235);
  assign _zz_6853 = _zz_6854;
  assign _zz_6854 = ($signed(_zz_6856) + $signed(_zz_232));
  assign _zz_6855 = ({8'd0,data_mid_92_imag} <<< 8);
  assign _zz_6856 = {{8{_zz_6855[23]}}, _zz_6855};
  assign _zz_6857 = fixTo_281_dout;
  assign _zz_6858 = ($signed(twiddle_factor_table_0_real) + $signed(twiddle_factor_table_0_imag));
  assign _zz_6859 = ($signed(_zz_238) - $signed(_zz_6860));
  assign _zz_6860 = ($signed(_zz_6861) * $signed(twiddle_factor_table_0_imag));
  assign _zz_6861 = ($signed(data_mid_95_real) + $signed(data_mid_95_imag));
  assign _zz_6862 = fixTo_282_dout;
  assign _zz_6863 = ($signed(_zz_238) + $signed(_zz_6864));
  assign _zz_6864 = ($signed(_zz_6865) * $signed(twiddle_factor_table_0_real));
  assign _zz_6865 = ($signed(data_mid_95_imag) - $signed(data_mid_95_real));
  assign _zz_6866 = fixTo_283_dout;
  assign _zz_6867 = _zz_6868[31 : 0];
  assign _zz_6868 = _zz_6869;
  assign _zz_6869 = ($signed(_zz_6870) >>> _zz_239);
  assign _zz_6870 = _zz_6871;
  assign _zz_6871 = ($signed(_zz_6873) - $signed(_zz_236));
  assign _zz_6872 = ({8'd0,data_mid_94_real} <<< 8);
  assign _zz_6873 = {{8{_zz_6872[23]}}, _zz_6872};
  assign _zz_6874 = fixTo_284_dout;
  assign _zz_6875 = _zz_6876[31 : 0];
  assign _zz_6876 = _zz_6877;
  assign _zz_6877 = ($signed(_zz_6878) >>> _zz_239);
  assign _zz_6878 = _zz_6879;
  assign _zz_6879 = ($signed(_zz_6881) - $signed(_zz_237));
  assign _zz_6880 = ({8'd0,data_mid_94_imag} <<< 8);
  assign _zz_6881 = {{8{_zz_6880[23]}}, _zz_6880};
  assign _zz_6882 = fixTo_285_dout;
  assign _zz_6883 = _zz_6884[31 : 0];
  assign _zz_6884 = _zz_6885;
  assign _zz_6885 = ($signed(_zz_6886) >>> _zz_240);
  assign _zz_6886 = _zz_6887;
  assign _zz_6887 = ($signed(_zz_6889) + $signed(_zz_236));
  assign _zz_6888 = ({8'd0,data_mid_94_real} <<< 8);
  assign _zz_6889 = {{8{_zz_6888[23]}}, _zz_6888};
  assign _zz_6890 = fixTo_286_dout;
  assign _zz_6891 = _zz_6892[31 : 0];
  assign _zz_6892 = _zz_6893;
  assign _zz_6893 = ($signed(_zz_6894) >>> _zz_240);
  assign _zz_6894 = _zz_6895;
  assign _zz_6895 = ($signed(_zz_6897) + $signed(_zz_237));
  assign _zz_6896 = ({8'd0,data_mid_94_imag} <<< 8);
  assign _zz_6897 = {{8{_zz_6896[23]}}, _zz_6896};
  assign _zz_6898 = fixTo_287_dout;
  assign _zz_6899 = ($signed(twiddle_factor_table_0_real) + $signed(twiddle_factor_table_0_imag));
  assign _zz_6900 = ($signed(_zz_243) - $signed(_zz_6901));
  assign _zz_6901 = ($signed(_zz_6902) * $signed(twiddle_factor_table_0_imag));
  assign _zz_6902 = ($signed(data_mid_97_real) + $signed(data_mid_97_imag));
  assign _zz_6903 = fixTo_288_dout;
  assign _zz_6904 = ($signed(_zz_243) + $signed(_zz_6905));
  assign _zz_6905 = ($signed(_zz_6906) * $signed(twiddle_factor_table_0_real));
  assign _zz_6906 = ($signed(data_mid_97_imag) - $signed(data_mid_97_real));
  assign _zz_6907 = fixTo_289_dout;
  assign _zz_6908 = _zz_6909[31 : 0];
  assign _zz_6909 = _zz_6910;
  assign _zz_6910 = ($signed(_zz_6911) >>> _zz_244);
  assign _zz_6911 = _zz_6912;
  assign _zz_6912 = ($signed(_zz_6914) - $signed(_zz_241));
  assign _zz_6913 = ({8'd0,data_mid_96_real} <<< 8);
  assign _zz_6914 = {{8{_zz_6913[23]}}, _zz_6913};
  assign _zz_6915 = fixTo_290_dout;
  assign _zz_6916 = _zz_6917[31 : 0];
  assign _zz_6917 = _zz_6918;
  assign _zz_6918 = ($signed(_zz_6919) >>> _zz_244);
  assign _zz_6919 = _zz_6920;
  assign _zz_6920 = ($signed(_zz_6922) - $signed(_zz_242));
  assign _zz_6921 = ({8'd0,data_mid_96_imag} <<< 8);
  assign _zz_6922 = {{8{_zz_6921[23]}}, _zz_6921};
  assign _zz_6923 = fixTo_291_dout;
  assign _zz_6924 = _zz_6925[31 : 0];
  assign _zz_6925 = _zz_6926;
  assign _zz_6926 = ($signed(_zz_6927) >>> _zz_245);
  assign _zz_6927 = _zz_6928;
  assign _zz_6928 = ($signed(_zz_6930) + $signed(_zz_241));
  assign _zz_6929 = ({8'd0,data_mid_96_real} <<< 8);
  assign _zz_6930 = {{8{_zz_6929[23]}}, _zz_6929};
  assign _zz_6931 = fixTo_292_dout;
  assign _zz_6932 = _zz_6933[31 : 0];
  assign _zz_6933 = _zz_6934;
  assign _zz_6934 = ($signed(_zz_6935) >>> _zz_245);
  assign _zz_6935 = _zz_6936;
  assign _zz_6936 = ($signed(_zz_6938) + $signed(_zz_242));
  assign _zz_6937 = ({8'd0,data_mid_96_imag} <<< 8);
  assign _zz_6938 = {{8{_zz_6937[23]}}, _zz_6937};
  assign _zz_6939 = fixTo_293_dout;
  assign _zz_6940 = ($signed(twiddle_factor_table_0_real) + $signed(twiddle_factor_table_0_imag));
  assign _zz_6941 = ($signed(_zz_248) - $signed(_zz_6942));
  assign _zz_6942 = ($signed(_zz_6943) * $signed(twiddle_factor_table_0_imag));
  assign _zz_6943 = ($signed(data_mid_99_real) + $signed(data_mid_99_imag));
  assign _zz_6944 = fixTo_294_dout;
  assign _zz_6945 = ($signed(_zz_248) + $signed(_zz_6946));
  assign _zz_6946 = ($signed(_zz_6947) * $signed(twiddle_factor_table_0_real));
  assign _zz_6947 = ($signed(data_mid_99_imag) - $signed(data_mid_99_real));
  assign _zz_6948 = fixTo_295_dout;
  assign _zz_6949 = _zz_6950[31 : 0];
  assign _zz_6950 = _zz_6951;
  assign _zz_6951 = ($signed(_zz_6952) >>> _zz_249);
  assign _zz_6952 = _zz_6953;
  assign _zz_6953 = ($signed(_zz_6955) - $signed(_zz_246));
  assign _zz_6954 = ({8'd0,data_mid_98_real} <<< 8);
  assign _zz_6955 = {{8{_zz_6954[23]}}, _zz_6954};
  assign _zz_6956 = fixTo_296_dout;
  assign _zz_6957 = _zz_6958[31 : 0];
  assign _zz_6958 = _zz_6959;
  assign _zz_6959 = ($signed(_zz_6960) >>> _zz_249);
  assign _zz_6960 = _zz_6961;
  assign _zz_6961 = ($signed(_zz_6963) - $signed(_zz_247));
  assign _zz_6962 = ({8'd0,data_mid_98_imag} <<< 8);
  assign _zz_6963 = {{8{_zz_6962[23]}}, _zz_6962};
  assign _zz_6964 = fixTo_297_dout;
  assign _zz_6965 = _zz_6966[31 : 0];
  assign _zz_6966 = _zz_6967;
  assign _zz_6967 = ($signed(_zz_6968) >>> _zz_250);
  assign _zz_6968 = _zz_6969;
  assign _zz_6969 = ($signed(_zz_6971) + $signed(_zz_246));
  assign _zz_6970 = ({8'd0,data_mid_98_real} <<< 8);
  assign _zz_6971 = {{8{_zz_6970[23]}}, _zz_6970};
  assign _zz_6972 = fixTo_298_dout;
  assign _zz_6973 = _zz_6974[31 : 0];
  assign _zz_6974 = _zz_6975;
  assign _zz_6975 = ($signed(_zz_6976) >>> _zz_250);
  assign _zz_6976 = _zz_6977;
  assign _zz_6977 = ($signed(_zz_6979) + $signed(_zz_247));
  assign _zz_6978 = ({8'd0,data_mid_98_imag} <<< 8);
  assign _zz_6979 = {{8{_zz_6978[23]}}, _zz_6978};
  assign _zz_6980 = fixTo_299_dout;
  assign _zz_6981 = ($signed(twiddle_factor_table_0_real) + $signed(twiddle_factor_table_0_imag));
  assign _zz_6982 = ($signed(_zz_253) - $signed(_zz_6983));
  assign _zz_6983 = ($signed(_zz_6984) * $signed(twiddle_factor_table_0_imag));
  assign _zz_6984 = ($signed(data_mid_101_real) + $signed(data_mid_101_imag));
  assign _zz_6985 = fixTo_300_dout;
  assign _zz_6986 = ($signed(_zz_253) + $signed(_zz_6987));
  assign _zz_6987 = ($signed(_zz_6988) * $signed(twiddle_factor_table_0_real));
  assign _zz_6988 = ($signed(data_mid_101_imag) - $signed(data_mid_101_real));
  assign _zz_6989 = fixTo_301_dout;
  assign _zz_6990 = _zz_6991[31 : 0];
  assign _zz_6991 = _zz_6992;
  assign _zz_6992 = ($signed(_zz_6993) >>> _zz_254);
  assign _zz_6993 = _zz_6994;
  assign _zz_6994 = ($signed(_zz_6996) - $signed(_zz_251));
  assign _zz_6995 = ({8'd0,data_mid_100_real} <<< 8);
  assign _zz_6996 = {{8{_zz_6995[23]}}, _zz_6995};
  assign _zz_6997 = fixTo_302_dout;
  assign _zz_6998 = _zz_6999[31 : 0];
  assign _zz_6999 = _zz_7000;
  assign _zz_7000 = ($signed(_zz_7001) >>> _zz_254);
  assign _zz_7001 = _zz_7002;
  assign _zz_7002 = ($signed(_zz_7004) - $signed(_zz_252));
  assign _zz_7003 = ({8'd0,data_mid_100_imag} <<< 8);
  assign _zz_7004 = {{8{_zz_7003[23]}}, _zz_7003};
  assign _zz_7005 = fixTo_303_dout;
  assign _zz_7006 = _zz_7007[31 : 0];
  assign _zz_7007 = _zz_7008;
  assign _zz_7008 = ($signed(_zz_7009) >>> _zz_255);
  assign _zz_7009 = _zz_7010;
  assign _zz_7010 = ($signed(_zz_7012) + $signed(_zz_251));
  assign _zz_7011 = ({8'd0,data_mid_100_real} <<< 8);
  assign _zz_7012 = {{8{_zz_7011[23]}}, _zz_7011};
  assign _zz_7013 = fixTo_304_dout;
  assign _zz_7014 = _zz_7015[31 : 0];
  assign _zz_7015 = _zz_7016;
  assign _zz_7016 = ($signed(_zz_7017) >>> _zz_255);
  assign _zz_7017 = _zz_7018;
  assign _zz_7018 = ($signed(_zz_7020) + $signed(_zz_252));
  assign _zz_7019 = ({8'd0,data_mid_100_imag} <<< 8);
  assign _zz_7020 = {{8{_zz_7019[23]}}, _zz_7019};
  assign _zz_7021 = fixTo_305_dout;
  assign _zz_7022 = ($signed(twiddle_factor_table_0_real) + $signed(twiddle_factor_table_0_imag));
  assign _zz_7023 = ($signed(_zz_258) - $signed(_zz_7024));
  assign _zz_7024 = ($signed(_zz_7025) * $signed(twiddle_factor_table_0_imag));
  assign _zz_7025 = ($signed(data_mid_103_real) + $signed(data_mid_103_imag));
  assign _zz_7026 = fixTo_306_dout;
  assign _zz_7027 = ($signed(_zz_258) + $signed(_zz_7028));
  assign _zz_7028 = ($signed(_zz_7029) * $signed(twiddle_factor_table_0_real));
  assign _zz_7029 = ($signed(data_mid_103_imag) - $signed(data_mid_103_real));
  assign _zz_7030 = fixTo_307_dout;
  assign _zz_7031 = _zz_7032[31 : 0];
  assign _zz_7032 = _zz_7033;
  assign _zz_7033 = ($signed(_zz_7034) >>> _zz_259);
  assign _zz_7034 = _zz_7035;
  assign _zz_7035 = ($signed(_zz_7037) - $signed(_zz_256));
  assign _zz_7036 = ({8'd0,data_mid_102_real} <<< 8);
  assign _zz_7037 = {{8{_zz_7036[23]}}, _zz_7036};
  assign _zz_7038 = fixTo_308_dout;
  assign _zz_7039 = _zz_7040[31 : 0];
  assign _zz_7040 = _zz_7041;
  assign _zz_7041 = ($signed(_zz_7042) >>> _zz_259);
  assign _zz_7042 = _zz_7043;
  assign _zz_7043 = ($signed(_zz_7045) - $signed(_zz_257));
  assign _zz_7044 = ({8'd0,data_mid_102_imag} <<< 8);
  assign _zz_7045 = {{8{_zz_7044[23]}}, _zz_7044};
  assign _zz_7046 = fixTo_309_dout;
  assign _zz_7047 = _zz_7048[31 : 0];
  assign _zz_7048 = _zz_7049;
  assign _zz_7049 = ($signed(_zz_7050) >>> _zz_260);
  assign _zz_7050 = _zz_7051;
  assign _zz_7051 = ($signed(_zz_7053) + $signed(_zz_256));
  assign _zz_7052 = ({8'd0,data_mid_102_real} <<< 8);
  assign _zz_7053 = {{8{_zz_7052[23]}}, _zz_7052};
  assign _zz_7054 = fixTo_310_dout;
  assign _zz_7055 = _zz_7056[31 : 0];
  assign _zz_7056 = _zz_7057;
  assign _zz_7057 = ($signed(_zz_7058) >>> _zz_260);
  assign _zz_7058 = _zz_7059;
  assign _zz_7059 = ($signed(_zz_7061) + $signed(_zz_257));
  assign _zz_7060 = ({8'd0,data_mid_102_imag} <<< 8);
  assign _zz_7061 = {{8{_zz_7060[23]}}, _zz_7060};
  assign _zz_7062 = fixTo_311_dout;
  assign _zz_7063 = ($signed(twiddle_factor_table_0_real) + $signed(twiddle_factor_table_0_imag));
  assign _zz_7064 = ($signed(_zz_263) - $signed(_zz_7065));
  assign _zz_7065 = ($signed(_zz_7066) * $signed(twiddle_factor_table_0_imag));
  assign _zz_7066 = ($signed(data_mid_105_real) + $signed(data_mid_105_imag));
  assign _zz_7067 = fixTo_312_dout;
  assign _zz_7068 = ($signed(_zz_263) + $signed(_zz_7069));
  assign _zz_7069 = ($signed(_zz_7070) * $signed(twiddle_factor_table_0_real));
  assign _zz_7070 = ($signed(data_mid_105_imag) - $signed(data_mid_105_real));
  assign _zz_7071 = fixTo_313_dout;
  assign _zz_7072 = _zz_7073[31 : 0];
  assign _zz_7073 = _zz_7074;
  assign _zz_7074 = ($signed(_zz_7075) >>> _zz_264);
  assign _zz_7075 = _zz_7076;
  assign _zz_7076 = ($signed(_zz_7078) - $signed(_zz_261));
  assign _zz_7077 = ({8'd0,data_mid_104_real} <<< 8);
  assign _zz_7078 = {{8{_zz_7077[23]}}, _zz_7077};
  assign _zz_7079 = fixTo_314_dout;
  assign _zz_7080 = _zz_7081[31 : 0];
  assign _zz_7081 = _zz_7082;
  assign _zz_7082 = ($signed(_zz_7083) >>> _zz_264);
  assign _zz_7083 = _zz_7084;
  assign _zz_7084 = ($signed(_zz_7086) - $signed(_zz_262));
  assign _zz_7085 = ({8'd0,data_mid_104_imag} <<< 8);
  assign _zz_7086 = {{8{_zz_7085[23]}}, _zz_7085};
  assign _zz_7087 = fixTo_315_dout;
  assign _zz_7088 = _zz_7089[31 : 0];
  assign _zz_7089 = _zz_7090;
  assign _zz_7090 = ($signed(_zz_7091) >>> _zz_265);
  assign _zz_7091 = _zz_7092;
  assign _zz_7092 = ($signed(_zz_7094) + $signed(_zz_261));
  assign _zz_7093 = ({8'd0,data_mid_104_real} <<< 8);
  assign _zz_7094 = {{8{_zz_7093[23]}}, _zz_7093};
  assign _zz_7095 = fixTo_316_dout;
  assign _zz_7096 = _zz_7097[31 : 0];
  assign _zz_7097 = _zz_7098;
  assign _zz_7098 = ($signed(_zz_7099) >>> _zz_265);
  assign _zz_7099 = _zz_7100;
  assign _zz_7100 = ($signed(_zz_7102) + $signed(_zz_262));
  assign _zz_7101 = ({8'd0,data_mid_104_imag} <<< 8);
  assign _zz_7102 = {{8{_zz_7101[23]}}, _zz_7101};
  assign _zz_7103 = fixTo_317_dout;
  assign _zz_7104 = ($signed(twiddle_factor_table_0_real) + $signed(twiddle_factor_table_0_imag));
  assign _zz_7105 = ($signed(_zz_268) - $signed(_zz_7106));
  assign _zz_7106 = ($signed(_zz_7107) * $signed(twiddle_factor_table_0_imag));
  assign _zz_7107 = ($signed(data_mid_107_real) + $signed(data_mid_107_imag));
  assign _zz_7108 = fixTo_318_dout;
  assign _zz_7109 = ($signed(_zz_268) + $signed(_zz_7110));
  assign _zz_7110 = ($signed(_zz_7111) * $signed(twiddle_factor_table_0_real));
  assign _zz_7111 = ($signed(data_mid_107_imag) - $signed(data_mid_107_real));
  assign _zz_7112 = fixTo_319_dout;
  assign _zz_7113 = _zz_7114[31 : 0];
  assign _zz_7114 = _zz_7115;
  assign _zz_7115 = ($signed(_zz_7116) >>> _zz_269);
  assign _zz_7116 = _zz_7117;
  assign _zz_7117 = ($signed(_zz_7119) - $signed(_zz_266));
  assign _zz_7118 = ({8'd0,data_mid_106_real} <<< 8);
  assign _zz_7119 = {{8{_zz_7118[23]}}, _zz_7118};
  assign _zz_7120 = fixTo_320_dout;
  assign _zz_7121 = _zz_7122[31 : 0];
  assign _zz_7122 = _zz_7123;
  assign _zz_7123 = ($signed(_zz_7124) >>> _zz_269);
  assign _zz_7124 = _zz_7125;
  assign _zz_7125 = ($signed(_zz_7127) - $signed(_zz_267));
  assign _zz_7126 = ({8'd0,data_mid_106_imag} <<< 8);
  assign _zz_7127 = {{8{_zz_7126[23]}}, _zz_7126};
  assign _zz_7128 = fixTo_321_dout;
  assign _zz_7129 = _zz_7130[31 : 0];
  assign _zz_7130 = _zz_7131;
  assign _zz_7131 = ($signed(_zz_7132) >>> _zz_270);
  assign _zz_7132 = _zz_7133;
  assign _zz_7133 = ($signed(_zz_7135) + $signed(_zz_266));
  assign _zz_7134 = ({8'd0,data_mid_106_real} <<< 8);
  assign _zz_7135 = {{8{_zz_7134[23]}}, _zz_7134};
  assign _zz_7136 = fixTo_322_dout;
  assign _zz_7137 = _zz_7138[31 : 0];
  assign _zz_7138 = _zz_7139;
  assign _zz_7139 = ($signed(_zz_7140) >>> _zz_270);
  assign _zz_7140 = _zz_7141;
  assign _zz_7141 = ($signed(_zz_7143) + $signed(_zz_267));
  assign _zz_7142 = ({8'd0,data_mid_106_imag} <<< 8);
  assign _zz_7143 = {{8{_zz_7142[23]}}, _zz_7142};
  assign _zz_7144 = fixTo_323_dout;
  assign _zz_7145 = ($signed(twiddle_factor_table_0_real) + $signed(twiddle_factor_table_0_imag));
  assign _zz_7146 = ($signed(_zz_273) - $signed(_zz_7147));
  assign _zz_7147 = ($signed(_zz_7148) * $signed(twiddle_factor_table_0_imag));
  assign _zz_7148 = ($signed(data_mid_109_real) + $signed(data_mid_109_imag));
  assign _zz_7149 = fixTo_324_dout;
  assign _zz_7150 = ($signed(_zz_273) + $signed(_zz_7151));
  assign _zz_7151 = ($signed(_zz_7152) * $signed(twiddle_factor_table_0_real));
  assign _zz_7152 = ($signed(data_mid_109_imag) - $signed(data_mid_109_real));
  assign _zz_7153 = fixTo_325_dout;
  assign _zz_7154 = _zz_7155[31 : 0];
  assign _zz_7155 = _zz_7156;
  assign _zz_7156 = ($signed(_zz_7157) >>> _zz_274);
  assign _zz_7157 = _zz_7158;
  assign _zz_7158 = ($signed(_zz_7160) - $signed(_zz_271));
  assign _zz_7159 = ({8'd0,data_mid_108_real} <<< 8);
  assign _zz_7160 = {{8{_zz_7159[23]}}, _zz_7159};
  assign _zz_7161 = fixTo_326_dout;
  assign _zz_7162 = _zz_7163[31 : 0];
  assign _zz_7163 = _zz_7164;
  assign _zz_7164 = ($signed(_zz_7165) >>> _zz_274);
  assign _zz_7165 = _zz_7166;
  assign _zz_7166 = ($signed(_zz_7168) - $signed(_zz_272));
  assign _zz_7167 = ({8'd0,data_mid_108_imag} <<< 8);
  assign _zz_7168 = {{8{_zz_7167[23]}}, _zz_7167};
  assign _zz_7169 = fixTo_327_dout;
  assign _zz_7170 = _zz_7171[31 : 0];
  assign _zz_7171 = _zz_7172;
  assign _zz_7172 = ($signed(_zz_7173) >>> _zz_275);
  assign _zz_7173 = _zz_7174;
  assign _zz_7174 = ($signed(_zz_7176) + $signed(_zz_271));
  assign _zz_7175 = ({8'd0,data_mid_108_real} <<< 8);
  assign _zz_7176 = {{8{_zz_7175[23]}}, _zz_7175};
  assign _zz_7177 = fixTo_328_dout;
  assign _zz_7178 = _zz_7179[31 : 0];
  assign _zz_7179 = _zz_7180;
  assign _zz_7180 = ($signed(_zz_7181) >>> _zz_275);
  assign _zz_7181 = _zz_7182;
  assign _zz_7182 = ($signed(_zz_7184) + $signed(_zz_272));
  assign _zz_7183 = ({8'd0,data_mid_108_imag} <<< 8);
  assign _zz_7184 = {{8{_zz_7183[23]}}, _zz_7183};
  assign _zz_7185 = fixTo_329_dout;
  assign _zz_7186 = ($signed(twiddle_factor_table_0_real) + $signed(twiddle_factor_table_0_imag));
  assign _zz_7187 = ($signed(_zz_278) - $signed(_zz_7188));
  assign _zz_7188 = ($signed(_zz_7189) * $signed(twiddle_factor_table_0_imag));
  assign _zz_7189 = ($signed(data_mid_111_real) + $signed(data_mid_111_imag));
  assign _zz_7190 = fixTo_330_dout;
  assign _zz_7191 = ($signed(_zz_278) + $signed(_zz_7192));
  assign _zz_7192 = ($signed(_zz_7193) * $signed(twiddle_factor_table_0_real));
  assign _zz_7193 = ($signed(data_mid_111_imag) - $signed(data_mid_111_real));
  assign _zz_7194 = fixTo_331_dout;
  assign _zz_7195 = _zz_7196[31 : 0];
  assign _zz_7196 = _zz_7197;
  assign _zz_7197 = ($signed(_zz_7198) >>> _zz_279);
  assign _zz_7198 = _zz_7199;
  assign _zz_7199 = ($signed(_zz_7201) - $signed(_zz_276));
  assign _zz_7200 = ({8'd0,data_mid_110_real} <<< 8);
  assign _zz_7201 = {{8{_zz_7200[23]}}, _zz_7200};
  assign _zz_7202 = fixTo_332_dout;
  assign _zz_7203 = _zz_7204[31 : 0];
  assign _zz_7204 = _zz_7205;
  assign _zz_7205 = ($signed(_zz_7206) >>> _zz_279);
  assign _zz_7206 = _zz_7207;
  assign _zz_7207 = ($signed(_zz_7209) - $signed(_zz_277));
  assign _zz_7208 = ({8'd0,data_mid_110_imag} <<< 8);
  assign _zz_7209 = {{8{_zz_7208[23]}}, _zz_7208};
  assign _zz_7210 = fixTo_333_dout;
  assign _zz_7211 = _zz_7212[31 : 0];
  assign _zz_7212 = _zz_7213;
  assign _zz_7213 = ($signed(_zz_7214) >>> _zz_280);
  assign _zz_7214 = _zz_7215;
  assign _zz_7215 = ($signed(_zz_7217) + $signed(_zz_276));
  assign _zz_7216 = ({8'd0,data_mid_110_real} <<< 8);
  assign _zz_7217 = {{8{_zz_7216[23]}}, _zz_7216};
  assign _zz_7218 = fixTo_334_dout;
  assign _zz_7219 = _zz_7220[31 : 0];
  assign _zz_7220 = _zz_7221;
  assign _zz_7221 = ($signed(_zz_7222) >>> _zz_280);
  assign _zz_7222 = _zz_7223;
  assign _zz_7223 = ($signed(_zz_7225) + $signed(_zz_277));
  assign _zz_7224 = ({8'd0,data_mid_110_imag} <<< 8);
  assign _zz_7225 = {{8{_zz_7224[23]}}, _zz_7224};
  assign _zz_7226 = fixTo_335_dout;
  assign _zz_7227 = ($signed(twiddle_factor_table_0_real) + $signed(twiddle_factor_table_0_imag));
  assign _zz_7228 = ($signed(_zz_283) - $signed(_zz_7229));
  assign _zz_7229 = ($signed(_zz_7230) * $signed(twiddle_factor_table_0_imag));
  assign _zz_7230 = ($signed(data_mid_113_real) + $signed(data_mid_113_imag));
  assign _zz_7231 = fixTo_336_dout;
  assign _zz_7232 = ($signed(_zz_283) + $signed(_zz_7233));
  assign _zz_7233 = ($signed(_zz_7234) * $signed(twiddle_factor_table_0_real));
  assign _zz_7234 = ($signed(data_mid_113_imag) - $signed(data_mid_113_real));
  assign _zz_7235 = fixTo_337_dout;
  assign _zz_7236 = _zz_7237[31 : 0];
  assign _zz_7237 = _zz_7238;
  assign _zz_7238 = ($signed(_zz_7239) >>> _zz_284);
  assign _zz_7239 = _zz_7240;
  assign _zz_7240 = ($signed(_zz_7242) - $signed(_zz_281));
  assign _zz_7241 = ({8'd0,data_mid_112_real} <<< 8);
  assign _zz_7242 = {{8{_zz_7241[23]}}, _zz_7241};
  assign _zz_7243 = fixTo_338_dout;
  assign _zz_7244 = _zz_7245[31 : 0];
  assign _zz_7245 = _zz_7246;
  assign _zz_7246 = ($signed(_zz_7247) >>> _zz_284);
  assign _zz_7247 = _zz_7248;
  assign _zz_7248 = ($signed(_zz_7250) - $signed(_zz_282));
  assign _zz_7249 = ({8'd0,data_mid_112_imag} <<< 8);
  assign _zz_7250 = {{8{_zz_7249[23]}}, _zz_7249};
  assign _zz_7251 = fixTo_339_dout;
  assign _zz_7252 = _zz_7253[31 : 0];
  assign _zz_7253 = _zz_7254;
  assign _zz_7254 = ($signed(_zz_7255) >>> _zz_285);
  assign _zz_7255 = _zz_7256;
  assign _zz_7256 = ($signed(_zz_7258) + $signed(_zz_281));
  assign _zz_7257 = ({8'd0,data_mid_112_real} <<< 8);
  assign _zz_7258 = {{8{_zz_7257[23]}}, _zz_7257};
  assign _zz_7259 = fixTo_340_dout;
  assign _zz_7260 = _zz_7261[31 : 0];
  assign _zz_7261 = _zz_7262;
  assign _zz_7262 = ($signed(_zz_7263) >>> _zz_285);
  assign _zz_7263 = _zz_7264;
  assign _zz_7264 = ($signed(_zz_7266) + $signed(_zz_282));
  assign _zz_7265 = ({8'd0,data_mid_112_imag} <<< 8);
  assign _zz_7266 = {{8{_zz_7265[23]}}, _zz_7265};
  assign _zz_7267 = fixTo_341_dout;
  assign _zz_7268 = ($signed(twiddle_factor_table_0_real) + $signed(twiddle_factor_table_0_imag));
  assign _zz_7269 = ($signed(_zz_288) - $signed(_zz_7270));
  assign _zz_7270 = ($signed(_zz_7271) * $signed(twiddle_factor_table_0_imag));
  assign _zz_7271 = ($signed(data_mid_115_real) + $signed(data_mid_115_imag));
  assign _zz_7272 = fixTo_342_dout;
  assign _zz_7273 = ($signed(_zz_288) + $signed(_zz_7274));
  assign _zz_7274 = ($signed(_zz_7275) * $signed(twiddle_factor_table_0_real));
  assign _zz_7275 = ($signed(data_mid_115_imag) - $signed(data_mid_115_real));
  assign _zz_7276 = fixTo_343_dout;
  assign _zz_7277 = _zz_7278[31 : 0];
  assign _zz_7278 = _zz_7279;
  assign _zz_7279 = ($signed(_zz_7280) >>> _zz_289);
  assign _zz_7280 = _zz_7281;
  assign _zz_7281 = ($signed(_zz_7283) - $signed(_zz_286));
  assign _zz_7282 = ({8'd0,data_mid_114_real} <<< 8);
  assign _zz_7283 = {{8{_zz_7282[23]}}, _zz_7282};
  assign _zz_7284 = fixTo_344_dout;
  assign _zz_7285 = _zz_7286[31 : 0];
  assign _zz_7286 = _zz_7287;
  assign _zz_7287 = ($signed(_zz_7288) >>> _zz_289);
  assign _zz_7288 = _zz_7289;
  assign _zz_7289 = ($signed(_zz_7291) - $signed(_zz_287));
  assign _zz_7290 = ({8'd0,data_mid_114_imag} <<< 8);
  assign _zz_7291 = {{8{_zz_7290[23]}}, _zz_7290};
  assign _zz_7292 = fixTo_345_dout;
  assign _zz_7293 = _zz_7294[31 : 0];
  assign _zz_7294 = _zz_7295;
  assign _zz_7295 = ($signed(_zz_7296) >>> _zz_290);
  assign _zz_7296 = _zz_7297;
  assign _zz_7297 = ($signed(_zz_7299) + $signed(_zz_286));
  assign _zz_7298 = ({8'd0,data_mid_114_real} <<< 8);
  assign _zz_7299 = {{8{_zz_7298[23]}}, _zz_7298};
  assign _zz_7300 = fixTo_346_dout;
  assign _zz_7301 = _zz_7302[31 : 0];
  assign _zz_7302 = _zz_7303;
  assign _zz_7303 = ($signed(_zz_7304) >>> _zz_290);
  assign _zz_7304 = _zz_7305;
  assign _zz_7305 = ($signed(_zz_7307) + $signed(_zz_287));
  assign _zz_7306 = ({8'd0,data_mid_114_imag} <<< 8);
  assign _zz_7307 = {{8{_zz_7306[23]}}, _zz_7306};
  assign _zz_7308 = fixTo_347_dout;
  assign _zz_7309 = ($signed(twiddle_factor_table_0_real) + $signed(twiddle_factor_table_0_imag));
  assign _zz_7310 = ($signed(_zz_293) - $signed(_zz_7311));
  assign _zz_7311 = ($signed(_zz_7312) * $signed(twiddle_factor_table_0_imag));
  assign _zz_7312 = ($signed(data_mid_117_real) + $signed(data_mid_117_imag));
  assign _zz_7313 = fixTo_348_dout;
  assign _zz_7314 = ($signed(_zz_293) + $signed(_zz_7315));
  assign _zz_7315 = ($signed(_zz_7316) * $signed(twiddle_factor_table_0_real));
  assign _zz_7316 = ($signed(data_mid_117_imag) - $signed(data_mid_117_real));
  assign _zz_7317 = fixTo_349_dout;
  assign _zz_7318 = _zz_7319[31 : 0];
  assign _zz_7319 = _zz_7320;
  assign _zz_7320 = ($signed(_zz_7321) >>> _zz_294);
  assign _zz_7321 = _zz_7322;
  assign _zz_7322 = ($signed(_zz_7324) - $signed(_zz_291));
  assign _zz_7323 = ({8'd0,data_mid_116_real} <<< 8);
  assign _zz_7324 = {{8{_zz_7323[23]}}, _zz_7323};
  assign _zz_7325 = fixTo_350_dout;
  assign _zz_7326 = _zz_7327[31 : 0];
  assign _zz_7327 = _zz_7328;
  assign _zz_7328 = ($signed(_zz_7329) >>> _zz_294);
  assign _zz_7329 = _zz_7330;
  assign _zz_7330 = ($signed(_zz_7332) - $signed(_zz_292));
  assign _zz_7331 = ({8'd0,data_mid_116_imag} <<< 8);
  assign _zz_7332 = {{8{_zz_7331[23]}}, _zz_7331};
  assign _zz_7333 = fixTo_351_dout;
  assign _zz_7334 = _zz_7335[31 : 0];
  assign _zz_7335 = _zz_7336;
  assign _zz_7336 = ($signed(_zz_7337) >>> _zz_295);
  assign _zz_7337 = _zz_7338;
  assign _zz_7338 = ($signed(_zz_7340) + $signed(_zz_291));
  assign _zz_7339 = ({8'd0,data_mid_116_real} <<< 8);
  assign _zz_7340 = {{8{_zz_7339[23]}}, _zz_7339};
  assign _zz_7341 = fixTo_352_dout;
  assign _zz_7342 = _zz_7343[31 : 0];
  assign _zz_7343 = _zz_7344;
  assign _zz_7344 = ($signed(_zz_7345) >>> _zz_295);
  assign _zz_7345 = _zz_7346;
  assign _zz_7346 = ($signed(_zz_7348) + $signed(_zz_292));
  assign _zz_7347 = ({8'd0,data_mid_116_imag} <<< 8);
  assign _zz_7348 = {{8{_zz_7347[23]}}, _zz_7347};
  assign _zz_7349 = fixTo_353_dout;
  assign _zz_7350 = ($signed(twiddle_factor_table_0_real) + $signed(twiddle_factor_table_0_imag));
  assign _zz_7351 = ($signed(_zz_298) - $signed(_zz_7352));
  assign _zz_7352 = ($signed(_zz_7353) * $signed(twiddle_factor_table_0_imag));
  assign _zz_7353 = ($signed(data_mid_119_real) + $signed(data_mid_119_imag));
  assign _zz_7354 = fixTo_354_dout;
  assign _zz_7355 = ($signed(_zz_298) + $signed(_zz_7356));
  assign _zz_7356 = ($signed(_zz_7357) * $signed(twiddle_factor_table_0_real));
  assign _zz_7357 = ($signed(data_mid_119_imag) - $signed(data_mid_119_real));
  assign _zz_7358 = fixTo_355_dout;
  assign _zz_7359 = _zz_7360[31 : 0];
  assign _zz_7360 = _zz_7361;
  assign _zz_7361 = ($signed(_zz_7362) >>> _zz_299);
  assign _zz_7362 = _zz_7363;
  assign _zz_7363 = ($signed(_zz_7365) - $signed(_zz_296));
  assign _zz_7364 = ({8'd0,data_mid_118_real} <<< 8);
  assign _zz_7365 = {{8{_zz_7364[23]}}, _zz_7364};
  assign _zz_7366 = fixTo_356_dout;
  assign _zz_7367 = _zz_7368[31 : 0];
  assign _zz_7368 = _zz_7369;
  assign _zz_7369 = ($signed(_zz_7370) >>> _zz_299);
  assign _zz_7370 = _zz_7371;
  assign _zz_7371 = ($signed(_zz_7373) - $signed(_zz_297));
  assign _zz_7372 = ({8'd0,data_mid_118_imag} <<< 8);
  assign _zz_7373 = {{8{_zz_7372[23]}}, _zz_7372};
  assign _zz_7374 = fixTo_357_dout;
  assign _zz_7375 = _zz_7376[31 : 0];
  assign _zz_7376 = _zz_7377;
  assign _zz_7377 = ($signed(_zz_7378) >>> _zz_300);
  assign _zz_7378 = _zz_7379;
  assign _zz_7379 = ($signed(_zz_7381) + $signed(_zz_296));
  assign _zz_7380 = ({8'd0,data_mid_118_real} <<< 8);
  assign _zz_7381 = {{8{_zz_7380[23]}}, _zz_7380};
  assign _zz_7382 = fixTo_358_dout;
  assign _zz_7383 = _zz_7384[31 : 0];
  assign _zz_7384 = _zz_7385;
  assign _zz_7385 = ($signed(_zz_7386) >>> _zz_300);
  assign _zz_7386 = _zz_7387;
  assign _zz_7387 = ($signed(_zz_7389) + $signed(_zz_297));
  assign _zz_7388 = ({8'd0,data_mid_118_imag} <<< 8);
  assign _zz_7389 = {{8{_zz_7388[23]}}, _zz_7388};
  assign _zz_7390 = fixTo_359_dout;
  assign _zz_7391 = ($signed(twiddle_factor_table_0_real) + $signed(twiddle_factor_table_0_imag));
  assign _zz_7392 = ($signed(_zz_303) - $signed(_zz_7393));
  assign _zz_7393 = ($signed(_zz_7394) * $signed(twiddle_factor_table_0_imag));
  assign _zz_7394 = ($signed(data_mid_121_real) + $signed(data_mid_121_imag));
  assign _zz_7395 = fixTo_360_dout;
  assign _zz_7396 = ($signed(_zz_303) + $signed(_zz_7397));
  assign _zz_7397 = ($signed(_zz_7398) * $signed(twiddle_factor_table_0_real));
  assign _zz_7398 = ($signed(data_mid_121_imag) - $signed(data_mid_121_real));
  assign _zz_7399 = fixTo_361_dout;
  assign _zz_7400 = _zz_7401[31 : 0];
  assign _zz_7401 = _zz_7402;
  assign _zz_7402 = ($signed(_zz_7403) >>> _zz_304);
  assign _zz_7403 = _zz_7404;
  assign _zz_7404 = ($signed(_zz_7406) - $signed(_zz_301));
  assign _zz_7405 = ({8'd0,data_mid_120_real} <<< 8);
  assign _zz_7406 = {{8{_zz_7405[23]}}, _zz_7405};
  assign _zz_7407 = fixTo_362_dout;
  assign _zz_7408 = _zz_7409[31 : 0];
  assign _zz_7409 = _zz_7410;
  assign _zz_7410 = ($signed(_zz_7411) >>> _zz_304);
  assign _zz_7411 = _zz_7412;
  assign _zz_7412 = ($signed(_zz_7414) - $signed(_zz_302));
  assign _zz_7413 = ({8'd0,data_mid_120_imag} <<< 8);
  assign _zz_7414 = {{8{_zz_7413[23]}}, _zz_7413};
  assign _zz_7415 = fixTo_363_dout;
  assign _zz_7416 = _zz_7417[31 : 0];
  assign _zz_7417 = _zz_7418;
  assign _zz_7418 = ($signed(_zz_7419) >>> _zz_305);
  assign _zz_7419 = _zz_7420;
  assign _zz_7420 = ($signed(_zz_7422) + $signed(_zz_301));
  assign _zz_7421 = ({8'd0,data_mid_120_real} <<< 8);
  assign _zz_7422 = {{8{_zz_7421[23]}}, _zz_7421};
  assign _zz_7423 = fixTo_364_dout;
  assign _zz_7424 = _zz_7425[31 : 0];
  assign _zz_7425 = _zz_7426;
  assign _zz_7426 = ($signed(_zz_7427) >>> _zz_305);
  assign _zz_7427 = _zz_7428;
  assign _zz_7428 = ($signed(_zz_7430) + $signed(_zz_302));
  assign _zz_7429 = ({8'd0,data_mid_120_imag} <<< 8);
  assign _zz_7430 = {{8{_zz_7429[23]}}, _zz_7429};
  assign _zz_7431 = fixTo_365_dout;
  assign _zz_7432 = ($signed(twiddle_factor_table_0_real) + $signed(twiddle_factor_table_0_imag));
  assign _zz_7433 = ($signed(_zz_308) - $signed(_zz_7434));
  assign _zz_7434 = ($signed(_zz_7435) * $signed(twiddle_factor_table_0_imag));
  assign _zz_7435 = ($signed(data_mid_123_real) + $signed(data_mid_123_imag));
  assign _zz_7436 = fixTo_366_dout;
  assign _zz_7437 = ($signed(_zz_308) + $signed(_zz_7438));
  assign _zz_7438 = ($signed(_zz_7439) * $signed(twiddle_factor_table_0_real));
  assign _zz_7439 = ($signed(data_mid_123_imag) - $signed(data_mid_123_real));
  assign _zz_7440 = fixTo_367_dout;
  assign _zz_7441 = _zz_7442[31 : 0];
  assign _zz_7442 = _zz_7443;
  assign _zz_7443 = ($signed(_zz_7444) >>> _zz_309);
  assign _zz_7444 = _zz_7445;
  assign _zz_7445 = ($signed(_zz_7447) - $signed(_zz_306));
  assign _zz_7446 = ({8'd0,data_mid_122_real} <<< 8);
  assign _zz_7447 = {{8{_zz_7446[23]}}, _zz_7446};
  assign _zz_7448 = fixTo_368_dout;
  assign _zz_7449 = _zz_7450[31 : 0];
  assign _zz_7450 = _zz_7451;
  assign _zz_7451 = ($signed(_zz_7452) >>> _zz_309);
  assign _zz_7452 = _zz_7453;
  assign _zz_7453 = ($signed(_zz_7455) - $signed(_zz_307));
  assign _zz_7454 = ({8'd0,data_mid_122_imag} <<< 8);
  assign _zz_7455 = {{8{_zz_7454[23]}}, _zz_7454};
  assign _zz_7456 = fixTo_369_dout;
  assign _zz_7457 = _zz_7458[31 : 0];
  assign _zz_7458 = _zz_7459;
  assign _zz_7459 = ($signed(_zz_7460) >>> _zz_310);
  assign _zz_7460 = _zz_7461;
  assign _zz_7461 = ($signed(_zz_7463) + $signed(_zz_306));
  assign _zz_7462 = ({8'd0,data_mid_122_real} <<< 8);
  assign _zz_7463 = {{8{_zz_7462[23]}}, _zz_7462};
  assign _zz_7464 = fixTo_370_dout;
  assign _zz_7465 = _zz_7466[31 : 0];
  assign _zz_7466 = _zz_7467;
  assign _zz_7467 = ($signed(_zz_7468) >>> _zz_310);
  assign _zz_7468 = _zz_7469;
  assign _zz_7469 = ($signed(_zz_7471) + $signed(_zz_307));
  assign _zz_7470 = ({8'd0,data_mid_122_imag} <<< 8);
  assign _zz_7471 = {{8{_zz_7470[23]}}, _zz_7470};
  assign _zz_7472 = fixTo_371_dout;
  assign _zz_7473 = ($signed(twiddle_factor_table_0_real) + $signed(twiddle_factor_table_0_imag));
  assign _zz_7474 = ($signed(_zz_313) - $signed(_zz_7475));
  assign _zz_7475 = ($signed(_zz_7476) * $signed(twiddle_factor_table_0_imag));
  assign _zz_7476 = ($signed(data_mid_125_real) + $signed(data_mid_125_imag));
  assign _zz_7477 = fixTo_372_dout;
  assign _zz_7478 = ($signed(_zz_313) + $signed(_zz_7479));
  assign _zz_7479 = ($signed(_zz_7480) * $signed(twiddle_factor_table_0_real));
  assign _zz_7480 = ($signed(data_mid_125_imag) - $signed(data_mid_125_real));
  assign _zz_7481 = fixTo_373_dout;
  assign _zz_7482 = _zz_7483[31 : 0];
  assign _zz_7483 = _zz_7484;
  assign _zz_7484 = ($signed(_zz_7485) >>> _zz_314);
  assign _zz_7485 = _zz_7486;
  assign _zz_7486 = ($signed(_zz_7488) - $signed(_zz_311));
  assign _zz_7487 = ({8'd0,data_mid_124_real} <<< 8);
  assign _zz_7488 = {{8{_zz_7487[23]}}, _zz_7487};
  assign _zz_7489 = fixTo_374_dout;
  assign _zz_7490 = _zz_7491[31 : 0];
  assign _zz_7491 = _zz_7492;
  assign _zz_7492 = ($signed(_zz_7493) >>> _zz_314);
  assign _zz_7493 = _zz_7494;
  assign _zz_7494 = ($signed(_zz_7496) - $signed(_zz_312));
  assign _zz_7495 = ({8'd0,data_mid_124_imag} <<< 8);
  assign _zz_7496 = {{8{_zz_7495[23]}}, _zz_7495};
  assign _zz_7497 = fixTo_375_dout;
  assign _zz_7498 = _zz_7499[31 : 0];
  assign _zz_7499 = _zz_7500;
  assign _zz_7500 = ($signed(_zz_7501) >>> _zz_315);
  assign _zz_7501 = _zz_7502;
  assign _zz_7502 = ($signed(_zz_7504) + $signed(_zz_311));
  assign _zz_7503 = ({8'd0,data_mid_124_real} <<< 8);
  assign _zz_7504 = {{8{_zz_7503[23]}}, _zz_7503};
  assign _zz_7505 = fixTo_376_dout;
  assign _zz_7506 = _zz_7507[31 : 0];
  assign _zz_7507 = _zz_7508;
  assign _zz_7508 = ($signed(_zz_7509) >>> _zz_315);
  assign _zz_7509 = _zz_7510;
  assign _zz_7510 = ($signed(_zz_7512) + $signed(_zz_312));
  assign _zz_7511 = ({8'd0,data_mid_124_imag} <<< 8);
  assign _zz_7512 = {{8{_zz_7511[23]}}, _zz_7511};
  assign _zz_7513 = fixTo_377_dout;
  assign _zz_7514 = ($signed(twiddle_factor_table_0_real) + $signed(twiddle_factor_table_0_imag));
  assign _zz_7515 = ($signed(_zz_318) - $signed(_zz_7516));
  assign _zz_7516 = ($signed(_zz_7517) * $signed(twiddle_factor_table_0_imag));
  assign _zz_7517 = ($signed(data_mid_127_real) + $signed(data_mid_127_imag));
  assign _zz_7518 = fixTo_378_dout;
  assign _zz_7519 = ($signed(_zz_318) + $signed(_zz_7520));
  assign _zz_7520 = ($signed(_zz_7521) * $signed(twiddle_factor_table_0_real));
  assign _zz_7521 = ($signed(data_mid_127_imag) - $signed(data_mid_127_real));
  assign _zz_7522 = fixTo_379_dout;
  assign _zz_7523 = _zz_7524[31 : 0];
  assign _zz_7524 = _zz_7525;
  assign _zz_7525 = ($signed(_zz_7526) >>> _zz_319);
  assign _zz_7526 = _zz_7527;
  assign _zz_7527 = ($signed(_zz_7529) - $signed(_zz_316));
  assign _zz_7528 = ({8'd0,data_mid_126_real} <<< 8);
  assign _zz_7529 = {{8{_zz_7528[23]}}, _zz_7528};
  assign _zz_7530 = fixTo_380_dout;
  assign _zz_7531 = _zz_7532[31 : 0];
  assign _zz_7532 = _zz_7533;
  assign _zz_7533 = ($signed(_zz_7534) >>> _zz_319);
  assign _zz_7534 = _zz_7535;
  assign _zz_7535 = ($signed(_zz_7537) - $signed(_zz_317));
  assign _zz_7536 = ({8'd0,data_mid_126_imag} <<< 8);
  assign _zz_7537 = {{8{_zz_7536[23]}}, _zz_7536};
  assign _zz_7538 = fixTo_381_dout;
  assign _zz_7539 = _zz_7540[31 : 0];
  assign _zz_7540 = _zz_7541;
  assign _zz_7541 = ($signed(_zz_7542) >>> _zz_320);
  assign _zz_7542 = _zz_7543;
  assign _zz_7543 = ($signed(_zz_7545) + $signed(_zz_316));
  assign _zz_7544 = ({8'd0,data_mid_126_real} <<< 8);
  assign _zz_7545 = {{8{_zz_7544[23]}}, _zz_7544};
  assign _zz_7546 = fixTo_382_dout;
  assign _zz_7547 = _zz_7548[31 : 0];
  assign _zz_7548 = _zz_7549;
  assign _zz_7549 = ($signed(_zz_7550) >>> _zz_320);
  assign _zz_7550 = _zz_7551;
  assign _zz_7551 = ($signed(_zz_7553) + $signed(_zz_317));
  assign _zz_7552 = ({8'd0,data_mid_126_imag} <<< 8);
  assign _zz_7553 = {{8{_zz_7552[23]}}, _zz_7552};
  assign _zz_7554 = fixTo_383_dout;
  assign _zz_7555 = ($signed(twiddle_factor_table_1_real) + $signed(twiddle_factor_table_1_imag));
  assign _zz_7556 = ($signed(_zz_323) - $signed(_zz_7557));
  assign _zz_7557 = ($signed(_zz_7558) * $signed(twiddle_factor_table_1_imag));
  assign _zz_7558 = ($signed(data_mid_2_real) + $signed(data_mid_2_imag));
  assign _zz_7559 = fixTo_384_dout;
  assign _zz_7560 = ($signed(_zz_323) + $signed(_zz_7561));
  assign _zz_7561 = ($signed(_zz_7562) * $signed(twiddle_factor_table_1_real));
  assign _zz_7562 = ($signed(data_mid_2_imag) - $signed(data_mid_2_real));
  assign _zz_7563 = fixTo_385_dout;
  assign _zz_7564 = _zz_7565[31 : 0];
  assign _zz_7565 = _zz_7566;
  assign _zz_7566 = ($signed(_zz_7567) >>> _zz_324);
  assign _zz_7567 = _zz_7568;
  assign _zz_7568 = ($signed(_zz_7570) - $signed(_zz_321));
  assign _zz_7569 = ({8'd0,data_mid_0_real} <<< 8);
  assign _zz_7570 = {{8{_zz_7569[23]}}, _zz_7569};
  assign _zz_7571 = fixTo_386_dout;
  assign _zz_7572 = _zz_7573[31 : 0];
  assign _zz_7573 = _zz_7574;
  assign _zz_7574 = ($signed(_zz_7575) >>> _zz_324);
  assign _zz_7575 = _zz_7576;
  assign _zz_7576 = ($signed(_zz_7578) - $signed(_zz_322));
  assign _zz_7577 = ({8'd0,data_mid_0_imag} <<< 8);
  assign _zz_7578 = {{8{_zz_7577[23]}}, _zz_7577};
  assign _zz_7579 = fixTo_387_dout;
  assign _zz_7580 = _zz_7581[31 : 0];
  assign _zz_7581 = _zz_7582;
  assign _zz_7582 = ($signed(_zz_7583) >>> _zz_325);
  assign _zz_7583 = _zz_7584;
  assign _zz_7584 = ($signed(_zz_7586) + $signed(_zz_321));
  assign _zz_7585 = ({8'd0,data_mid_0_real} <<< 8);
  assign _zz_7586 = {{8{_zz_7585[23]}}, _zz_7585};
  assign _zz_7587 = fixTo_388_dout;
  assign _zz_7588 = _zz_7589[31 : 0];
  assign _zz_7589 = _zz_7590;
  assign _zz_7590 = ($signed(_zz_7591) >>> _zz_325);
  assign _zz_7591 = _zz_7592;
  assign _zz_7592 = ($signed(_zz_7594) + $signed(_zz_322));
  assign _zz_7593 = ({8'd0,data_mid_0_imag} <<< 8);
  assign _zz_7594 = {{8{_zz_7593[23]}}, _zz_7593};
  assign _zz_7595 = fixTo_389_dout;
  assign _zz_7596 = ($signed(twiddle_factor_table_2_real) + $signed(twiddle_factor_table_2_imag));
  assign _zz_7597 = ($signed(_zz_328) - $signed(_zz_7598));
  assign _zz_7598 = ($signed(_zz_7599) * $signed(twiddle_factor_table_2_imag));
  assign _zz_7599 = ($signed(data_mid_3_real) + $signed(data_mid_3_imag));
  assign _zz_7600 = fixTo_390_dout;
  assign _zz_7601 = ($signed(_zz_328) + $signed(_zz_7602));
  assign _zz_7602 = ($signed(_zz_7603) * $signed(twiddle_factor_table_2_real));
  assign _zz_7603 = ($signed(data_mid_3_imag) - $signed(data_mid_3_real));
  assign _zz_7604 = fixTo_391_dout;
  assign _zz_7605 = _zz_7606[31 : 0];
  assign _zz_7606 = _zz_7607;
  assign _zz_7607 = ($signed(_zz_7608) >>> _zz_329);
  assign _zz_7608 = _zz_7609;
  assign _zz_7609 = ($signed(_zz_7611) - $signed(_zz_326));
  assign _zz_7610 = ({8'd0,data_mid_1_real} <<< 8);
  assign _zz_7611 = {{8{_zz_7610[23]}}, _zz_7610};
  assign _zz_7612 = fixTo_392_dout;
  assign _zz_7613 = _zz_7614[31 : 0];
  assign _zz_7614 = _zz_7615;
  assign _zz_7615 = ($signed(_zz_7616) >>> _zz_329);
  assign _zz_7616 = _zz_7617;
  assign _zz_7617 = ($signed(_zz_7619) - $signed(_zz_327));
  assign _zz_7618 = ({8'd0,data_mid_1_imag} <<< 8);
  assign _zz_7619 = {{8{_zz_7618[23]}}, _zz_7618};
  assign _zz_7620 = fixTo_393_dout;
  assign _zz_7621 = _zz_7622[31 : 0];
  assign _zz_7622 = _zz_7623;
  assign _zz_7623 = ($signed(_zz_7624) >>> _zz_330);
  assign _zz_7624 = _zz_7625;
  assign _zz_7625 = ($signed(_zz_7627) + $signed(_zz_326));
  assign _zz_7626 = ({8'd0,data_mid_1_real} <<< 8);
  assign _zz_7627 = {{8{_zz_7626[23]}}, _zz_7626};
  assign _zz_7628 = fixTo_394_dout;
  assign _zz_7629 = _zz_7630[31 : 0];
  assign _zz_7630 = _zz_7631;
  assign _zz_7631 = ($signed(_zz_7632) >>> _zz_330);
  assign _zz_7632 = _zz_7633;
  assign _zz_7633 = ($signed(_zz_7635) + $signed(_zz_327));
  assign _zz_7634 = ({8'd0,data_mid_1_imag} <<< 8);
  assign _zz_7635 = {{8{_zz_7634[23]}}, _zz_7634};
  assign _zz_7636 = fixTo_395_dout;
  assign _zz_7637 = ($signed(twiddle_factor_table_1_real) + $signed(twiddle_factor_table_1_imag));
  assign _zz_7638 = ($signed(_zz_333) - $signed(_zz_7639));
  assign _zz_7639 = ($signed(_zz_7640) * $signed(twiddle_factor_table_1_imag));
  assign _zz_7640 = ($signed(data_mid_6_real) + $signed(data_mid_6_imag));
  assign _zz_7641 = fixTo_396_dout;
  assign _zz_7642 = ($signed(_zz_333) + $signed(_zz_7643));
  assign _zz_7643 = ($signed(_zz_7644) * $signed(twiddle_factor_table_1_real));
  assign _zz_7644 = ($signed(data_mid_6_imag) - $signed(data_mid_6_real));
  assign _zz_7645 = fixTo_397_dout;
  assign _zz_7646 = _zz_7647[31 : 0];
  assign _zz_7647 = _zz_7648;
  assign _zz_7648 = ($signed(_zz_7649) >>> _zz_334);
  assign _zz_7649 = _zz_7650;
  assign _zz_7650 = ($signed(_zz_7652) - $signed(_zz_331));
  assign _zz_7651 = ({8'd0,data_mid_4_real} <<< 8);
  assign _zz_7652 = {{8{_zz_7651[23]}}, _zz_7651};
  assign _zz_7653 = fixTo_398_dout;
  assign _zz_7654 = _zz_7655[31 : 0];
  assign _zz_7655 = _zz_7656;
  assign _zz_7656 = ($signed(_zz_7657) >>> _zz_334);
  assign _zz_7657 = _zz_7658;
  assign _zz_7658 = ($signed(_zz_7660) - $signed(_zz_332));
  assign _zz_7659 = ({8'd0,data_mid_4_imag} <<< 8);
  assign _zz_7660 = {{8{_zz_7659[23]}}, _zz_7659};
  assign _zz_7661 = fixTo_399_dout;
  assign _zz_7662 = _zz_7663[31 : 0];
  assign _zz_7663 = _zz_7664;
  assign _zz_7664 = ($signed(_zz_7665) >>> _zz_335);
  assign _zz_7665 = _zz_7666;
  assign _zz_7666 = ($signed(_zz_7668) + $signed(_zz_331));
  assign _zz_7667 = ({8'd0,data_mid_4_real} <<< 8);
  assign _zz_7668 = {{8{_zz_7667[23]}}, _zz_7667};
  assign _zz_7669 = fixTo_400_dout;
  assign _zz_7670 = _zz_7671[31 : 0];
  assign _zz_7671 = _zz_7672;
  assign _zz_7672 = ($signed(_zz_7673) >>> _zz_335);
  assign _zz_7673 = _zz_7674;
  assign _zz_7674 = ($signed(_zz_7676) + $signed(_zz_332));
  assign _zz_7675 = ({8'd0,data_mid_4_imag} <<< 8);
  assign _zz_7676 = {{8{_zz_7675[23]}}, _zz_7675};
  assign _zz_7677 = fixTo_401_dout;
  assign _zz_7678 = ($signed(twiddle_factor_table_2_real) + $signed(twiddle_factor_table_2_imag));
  assign _zz_7679 = ($signed(_zz_338) - $signed(_zz_7680));
  assign _zz_7680 = ($signed(_zz_7681) * $signed(twiddle_factor_table_2_imag));
  assign _zz_7681 = ($signed(data_mid_7_real) + $signed(data_mid_7_imag));
  assign _zz_7682 = fixTo_402_dout;
  assign _zz_7683 = ($signed(_zz_338) + $signed(_zz_7684));
  assign _zz_7684 = ($signed(_zz_7685) * $signed(twiddle_factor_table_2_real));
  assign _zz_7685 = ($signed(data_mid_7_imag) - $signed(data_mid_7_real));
  assign _zz_7686 = fixTo_403_dout;
  assign _zz_7687 = _zz_7688[31 : 0];
  assign _zz_7688 = _zz_7689;
  assign _zz_7689 = ($signed(_zz_7690) >>> _zz_339);
  assign _zz_7690 = _zz_7691;
  assign _zz_7691 = ($signed(_zz_7693) - $signed(_zz_336));
  assign _zz_7692 = ({8'd0,data_mid_5_real} <<< 8);
  assign _zz_7693 = {{8{_zz_7692[23]}}, _zz_7692};
  assign _zz_7694 = fixTo_404_dout;
  assign _zz_7695 = _zz_7696[31 : 0];
  assign _zz_7696 = _zz_7697;
  assign _zz_7697 = ($signed(_zz_7698) >>> _zz_339);
  assign _zz_7698 = _zz_7699;
  assign _zz_7699 = ($signed(_zz_7701) - $signed(_zz_337));
  assign _zz_7700 = ({8'd0,data_mid_5_imag} <<< 8);
  assign _zz_7701 = {{8{_zz_7700[23]}}, _zz_7700};
  assign _zz_7702 = fixTo_405_dout;
  assign _zz_7703 = _zz_7704[31 : 0];
  assign _zz_7704 = _zz_7705;
  assign _zz_7705 = ($signed(_zz_7706) >>> _zz_340);
  assign _zz_7706 = _zz_7707;
  assign _zz_7707 = ($signed(_zz_7709) + $signed(_zz_336));
  assign _zz_7708 = ({8'd0,data_mid_5_real} <<< 8);
  assign _zz_7709 = {{8{_zz_7708[23]}}, _zz_7708};
  assign _zz_7710 = fixTo_406_dout;
  assign _zz_7711 = _zz_7712[31 : 0];
  assign _zz_7712 = _zz_7713;
  assign _zz_7713 = ($signed(_zz_7714) >>> _zz_340);
  assign _zz_7714 = _zz_7715;
  assign _zz_7715 = ($signed(_zz_7717) + $signed(_zz_337));
  assign _zz_7716 = ({8'd0,data_mid_5_imag} <<< 8);
  assign _zz_7717 = {{8{_zz_7716[23]}}, _zz_7716};
  assign _zz_7718 = fixTo_407_dout;
  assign _zz_7719 = ($signed(twiddle_factor_table_1_real) + $signed(twiddle_factor_table_1_imag));
  assign _zz_7720 = ($signed(_zz_343) - $signed(_zz_7721));
  assign _zz_7721 = ($signed(_zz_7722) * $signed(twiddle_factor_table_1_imag));
  assign _zz_7722 = ($signed(data_mid_10_real) + $signed(data_mid_10_imag));
  assign _zz_7723 = fixTo_408_dout;
  assign _zz_7724 = ($signed(_zz_343) + $signed(_zz_7725));
  assign _zz_7725 = ($signed(_zz_7726) * $signed(twiddle_factor_table_1_real));
  assign _zz_7726 = ($signed(data_mid_10_imag) - $signed(data_mid_10_real));
  assign _zz_7727 = fixTo_409_dout;
  assign _zz_7728 = _zz_7729[31 : 0];
  assign _zz_7729 = _zz_7730;
  assign _zz_7730 = ($signed(_zz_7731) >>> _zz_344);
  assign _zz_7731 = _zz_7732;
  assign _zz_7732 = ($signed(_zz_7734) - $signed(_zz_341));
  assign _zz_7733 = ({8'd0,data_mid_8_real} <<< 8);
  assign _zz_7734 = {{8{_zz_7733[23]}}, _zz_7733};
  assign _zz_7735 = fixTo_410_dout;
  assign _zz_7736 = _zz_7737[31 : 0];
  assign _zz_7737 = _zz_7738;
  assign _zz_7738 = ($signed(_zz_7739) >>> _zz_344);
  assign _zz_7739 = _zz_7740;
  assign _zz_7740 = ($signed(_zz_7742) - $signed(_zz_342));
  assign _zz_7741 = ({8'd0,data_mid_8_imag} <<< 8);
  assign _zz_7742 = {{8{_zz_7741[23]}}, _zz_7741};
  assign _zz_7743 = fixTo_411_dout;
  assign _zz_7744 = _zz_7745[31 : 0];
  assign _zz_7745 = _zz_7746;
  assign _zz_7746 = ($signed(_zz_7747) >>> _zz_345);
  assign _zz_7747 = _zz_7748;
  assign _zz_7748 = ($signed(_zz_7750) + $signed(_zz_341));
  assign _zz_7749 = ({8'd0,data_mid_8_real} <<< 8);
  assign _zz_7750 = {{8{_zz_7749[23]}}, _zz_7749};
  assign _zz_7751 = fixTo_412_dout;
  assign _zz_7752 = _zz_7753[31 : 0];
  assign _zz_7753 = _zz_7754;
  assign _zz_7754 = ($signed(_zz_7755) >>> _zz_345);
  assign _zz_7755 = _zz_7756;
  assign _zz_7756 = ($signed(_zz_7758) + $signed(_zz_342));
  assign _zz_7757 = ({8'd0,data_mid_8_imag} <<< 8);
  assign _zz_7758 = {{8{_zz_7757[23]}}, _zz_7757};
  assign _zz_7759 = fixTo_413_dout;
  assign _zz_7760 = ($signed(twiddle_factor_table_2_real) + $signed(twiddle_factor_table_2_imag));
  assign _zz_7761 = ($signed(_zz_348) - $signed(_zz_7762));
  assign _zz_7762 = ($signed(_zz_7763) * $signed(twiddle_factor_table_2_imag));
  assign _zz_7763 = ($signed(data_mid_11_real) + $signed(data_mid_11_imag));
  assign _zz_7764 = fixTo_414_dout;
  assign _zz_7765 = ($signed(_zz_348) + $signed(_zz_7766));
  assign _zz_7766 = ($signed(_zz_7767) * $signed(twiddle_factor_table_2_real));
  assign _zz_7767 = ($signed(data_mid_11_imag) - $signed(data_mid_11_real));
  assign _zz_7768 = fixTo_415_dout;
  assign _zz_7769 = _zz_7770[31 : 0];
  assign _zz_7770 = _zz_7771;
  assign _zz_7771 = ($signed(_zz_7772) >>> _zz_349);
  assign _zz_7772 = _zz_7773;
  assign _zz_7773 = ($signed(_zz_7775) - $signed(_zz_346));
  assign _zz_7774 = ({8'd0,data_mid_9_real} <<< 8);
  assign _zz_7775 = {{8{_zz_7774[23]}}, _zz_7774};
  assign _zz_7776 = fixTo_416_dout;
  assign _zz_7777 = _zz_7778[31 : 0];
  assign _zz_7778 = _zz_7779;
  assign _zz_7779 = ($signed(_zz_7780) >>> _zz_349);
  assign _zz_7780 = _zz_7781;
  assign _zz_7781 = ($signed(_zz_7783) - $signed(_zz_347));
  assign _zz_7782 = ({8'd0,data_mid_9_imag} <<< 8);
  assign _zz_7783 = {{8{_zz_7782[23]}}, _zz_7782};
  assign _zz_7784 = fixTo_417_dout;
  assign _zz_7785 = _zz_7786[31 : 0];
  assign _zz_7786 = _zz_7787;
  assign _zz_7787 = ($signed(_zz_7788) >>> _zz_350);
  assign _zz_7788 = _zz_7789;
  assign _zz_7789 = ($signed(_zz_7791) + $signed(_zz_346));
  assign _zz_7790 = ({8'd0,data_mid_9_real} <<< 8);
  assign _zz_7791 = {{8{_zz_7790[23]}}, _zz_7790};
  assign _zz_7792 = fixTo_418_dout;
  assign _zz_7793 = _zz_7794[31 : 0];
  assign _zz_7794 = _zz_7795;
  assign _zz_7795 = ($signed(_zz_7796) >>> _zz_350);
  assign _zz_7796 = _zz_7797;
  assign _zz_7797 = ($signed(_zz_7799) + $signed(_zz_347));
  assign _zz_7798 = ({8'd0,data_mid_9_imag} <<< 8);
  assign _zz_7799 = {{8{_zz_7798[23]}}, _zz_7798};
  assign _zz_7800 = fixTo_419_dout;
  assign _zz_7801 = ($signed(twiddle_factor_table_1_real) + $signed(twiddle_factor_table_1_imag));
  assign _zz_7802 = ($signed(_zz_353) - $signed(_zz_7803));
  assign _zz_7803 = ($signed(_zz_7804) * $signed(twiddle_factor_table_1_imag));
  assign _zz_7804 = ($signed(data_mid_14_real) + $signed(data_mid_14_imag));
  assign _zz_7805 = fixTo_420_dout;
  assign _zz_7806 = ($signed(_zz_353) + $signed(_zz_7807));
  assign _zz_7807 = ($signed(_zz_7808) * $signed(twiddle_factor_table_1_real));
  assign _zz_7808 = ($signed(data_mid_14_imag) - $signed(data_mid_14_real));
  assign _zz_7809 = fixTo_421_dout;
  assign _zz_7810 = _zz_7811[31 : 0];
  assign _zz_7811 = _zz_7812;
  assign _zz_7812 = ($signed(_zz_7813) >>> _zz_354);
  assign _zz_7813 = _zz_7814;
  assign _zz_7814 = ($signed(_zz_7816) - $signed(_zz_351));
  assign _zz_7815 = ({8'd0,data_mid_12_real} <<< 8);
  assign _zz_7816 = {{8{_zz_7815[23]}}, _zz_7815};
  assign _zz_7817 = fixTo_422_dout;
  assign _zz_7818 = _zz_7819[31 : 0];
  assign _zz_7819 = _zz_7820;
  assign _zz_7820 = ($signed(_zz_7821) >>> _zz_354);
  assign _zz_7821 = _zz_7822;
  assign _zz_7822 = ($signed(_zz_7824) - $signed(_zz_352));
  assign _zz_7823 = ({8'd0,data_mid_12_imag} <<< 8);
  assign _zz_7824 = {{8{_zz_7823[23]}}, _zz_7823};
  assign _zz_7825 = fixTo_423_dout;
  assign _zz_7826 = _zz_7827[31 : 0];
  assign _zz_7827 = _zz_7828;
  assign _zz_7828 = ($signed(_zz_7829) >>> _zz_355);
  assign _zz_7829 = _zz_7830;
  assign _zz_7830 = ($signed(_zz_7832) + $signed(_zz_351));
  assign _zz_7831 = ({8'd0,data_mid_12_real} <<< 8);
  assign _zz_7832 = {{8{_zz_7831[23]}}, _zz_7831};
  assign _zz_7833 = fixTo_424_dout;
  assign _zz_7834 = _zz_7835[31 : 0];
  assign _zz_7835 = _zz_7836;
  assign _zz_7836 = ($signed(_zz_7837) >>> _zz_355);
  assign _zz_7837 = _zz_7838;
  assign _zz_7838 = ($signed(_zz_7840) + $signed(_zz_352));
  assign _zz_7839 = ({8'd0,data_mid_12_imag} <<< 8);
  assign _zz_7840 = {{8{_zz_7839[23]}}, _zz_7839};
  assign _zz_7841 = fixTo_425_dout;
  assign _zz_7842 = ($signed(twiddle_factor_table_2_real) + $signed(twiddle_factor_table_2_imag));
  assign _zz_7843 = ($signed(_zz_358) - $signed(_zz_7844));
  assign _zz_7844 = ($signed(_zz_7845) * $signed(twiddle_factor_table_2_imag));
  assign _zz_7845 = ($signed(data_mid_15_real) + $signed(data_mid_15_imag));
  assign _zz_7846 = fixTo_426_dout;
  assign _zz_7847 = ($signed(_zz_358) + $signed(_zz_7848));
  assign _zz_7848 = ($signed(_zz_7849) * $signed(twiddle_factor_table_2_real));
  assign _zz_7849 = ($signed(data_mid_15_imag) - $signed(data_mid_15_real));
  assign _zz_7850 = fixTo_427_dout;
  assign _zz_7851 = _zz_7852[31 : 0];
  assign _zz_7852 = _zz_7853;
  assign _zz_7853 = ($signed(_zz_7854) >>> _zz_359);
  assign _zz_7854 = _zz_7855;
  assign _zz_7855 = ($signed(_zz_7857) - $signed(_zz_356));
  assign _zz_7856 = ({8'd0,data_mid_13_real} <<< 8);
  assign _zz_7857 = {{8{_zz_7856[23]}}, _zz_7856};
  assign _zz_7858 = fixTo_428_dout;
  assign _zz_7859 = _zz_7860[31 : 0];
  assign _zz_7860 = _zz_7861;
  assign _zz_7861 = ($signed(_zz_7862) >>> _zz_359);
  assign _zz_7862 = _zz_7863;
  assign _zz_7863 = ($signed(_zz_7865) - $signed(_zz_357));
  assign _zz_7864 = ({8'd0,data_mid_13_imag} <<< 8);
  assign _zz_7865 = {{8{_zz_7864[23]}}, _zz_7864};
  assign _zz_7866 = fixTo_429_dout;
  assign _zz_7867 = _zz_7868[31 : 0];
  assign _zz_7868 = _zz_7869;
  assign _zz_7869 = ($signed(_zz_7870) >>> _zz_360);
  assign _zz_7870 = _zz_7871;
  assign _zz_7871 = ($signed(_zz_7873) + $signed(_zz_356));
  assign _zz_7872 = ({8'd0,data_mid_13_real} <<< 8);
  assign _zz_7873 = {{8{_zz_7872[23]}}, _zz_7872};
  assign _zz_7874 = fixTo_430_dout;
  assign _zz_7875 = _zz_7876[31 : 0];
  assign _zz_7876 = _zz_7877;
  assign _zz_7877 = ($signed(_zz_7878) >>> _zz_360);
  assign _zz_7878 = _zz_7879;
  assign _zz_7879 = ($signed(_zz_7881) + $signed(_zz_357));
  assign _zz_7880 = ({8'd0,data_mid_13_imag} <<< 8);
  assign _zz_7881 = {{8{_zz_7880[23]}}, _zz_7880};
  assign _zz_7882 = fixTo_431_dout;
  assign _zz_7883 = ($signed(twiddle_factor_table_1_real) + $signed(twiddle_factor_table_1_imag));
  assign _zz_7884 = ($signed(_zz_363) - $signed(_zz_7885));
  assign _zz_7885 = ($signed(_zz_7886) * $signed(twiddle_factor_table_1_imag));
  assign _zz_7886 = ($signed(data_mid_18_real) + $signed(data_mid_18_imag));
  assign _zz_7887 = fixTo_432_dout;
  assign _zz_7888 = ($signed(_zz_363) + $signed(_zz_7889));
  assign _zz_7889 = ($signed(_zz_7890) * $signed(twiddle_factor_table_1_real));
  assign _zz_7890 = ($signed(data_mid_18_imag) - $signed(data_mid_18_real));
  assign _zz_7891 = fixTo_433_dout;
  assign _zz_7892 = _zz_7893[31 : 0];
  assign _zz_7893 = _zz_7894;
  assign _zz_7894 = ($signed(_zz_7895) >>> _zz_364);
  assign _zz_7895 = _zz_7896;
  assign _zz_7896 = ($signed(_zz_7898) - $signed(_zz_361));
  assign _zz_7897 = ({8'd0,data_mid_16_real} <<< 8);
  assign _zz_7898 = {{8{_zz_7897[23]}}, _zz_7897};
  assign _zz_7899 = fixTo_434_dout;
  assign _zz_7900 = _zz_7901[31 : 0];
  assign _zz_7901 = _zz_7902;
  assign _zz_7902 = ($signed(_zz_7903) >>> _zz_364);
  assign _zz_7903 = _zz_7904;
  assign _zz_7904 = ($signed(_zz_7906) - $signed(_zz_362));
  assign _zz_7905 = ({8'd0,data_mid_16_imag} <<< 8);
  assign _zz_7906 = {{8{_zz_7905[23]}}, _zz_7905};
  assign _zz_7907 = fixTo_435_dout;
  assign _zz_7908 = _zz_7909[31 : 0];
  assign _zz_7909 = _zz_7910;
  assign _zz_7910 = ($signed(_zz_7911) >>> _zz_365);
  assign _zz_7911 = _zz_7912;
  assign _zz_7912 = ($signed(_zz_7914) + $signed(_zz_361));
  assign _zz_7913 = ({8'd0,data_mid_16_real} <<< 8);
  assign _zz_7914 = {{8{_zz_7913[23]}}, _zz_7913};
  assign _zz_7915 = fixTo_436_dout;
  assign _zz_7916 = _zz_7917[31 : 0];
  assign _zz_7917 = _zz_7918;
  assign _zz_7918 = ($signed(_zz_7919) >>> _zz_365);
  assign _zz_7919 = _zz_7920;
  assign _zz_7920 = ($signed(_zz_7922) + $signed(_zz_362));
  assign _zz_7921 = ({8'd0,data_mid_16_imag} <<< 8);
  assign _zz_7922 = {{8{_zz_7921[23]}}, _zz_7921};
  assign _zz_7923 = fixTo_437_dout;
  assign _zz_7924 = ($signed(twiddle_factor_table_2_real) + $signed(twiddle_factor_table_2_imag));
  assign _zz_7925 = ($signed(_zz_368) - $signed(_zz_7926));
  assign _zz_7926 = ($signed(_zz_7927) * $signed(twiddle_factor_table_2_imag));
  assign _zz_7927 = ($signed(data_mid_19_real) + $signed(data_mid_19_imag));
  assign _zz_7928 = fixTo_438_dout;
  assign _zz_7929 = ($signed(_zz_368) + $signed(_zz_7930));
  assign _zz_7930 = ($signed(_zz_7931) * $signed(twiddle_factor_table_2_real));
  assign _zz_7931 = ($signed(data_mid_19_imag) - $signed(data_mid_19_real));
  assign _zz_7932 = fixTo_439_dout;
  assign _zz_7933 = _zz_7934[31 : 0];
  assign _zz_7934 = _zz_7935;
  assign _zz_7935 = ($signed(_zz_7936) >>> _zz_369);
  assign _zz_7936 = _zz_7937;
  assign _zz_7937 = ($signed(_zz_7939) - $signed(_zz_366));
  assign _zz_7938 = ({8'd0,data_mid_17_real} <<< 8);
  assign _zz_7939 = {{8{_zz_7938[23]}}, _zz_7938};
  assign _zz_7940 = fixTo_440_dout;
  assign _zz_7941 = _zz_7942[31 : 0];
  assign _zz_7942 = _zz_7943;
  assign _zz_7943 = ($signed(_zz_7944) >>> _zz_369);
  assign _zz_7944 = _zz_7945;
  assign _zz_7945 = ($signed(_zz_7947) - $signed(_zz_367));
  assign _zz_7946 = ({8'd0,data_mid_17_imag} <<< 8);
  assign _zz_7947 = {{8{_zz_7946[23]}}, _zz_7946};
  assign _zz_7948 = fixTo_441_dout;
  assign _zz_7949 = _zz_7950[31 : 0];
  assign _zz_7950 = _zz_7951;
  assign _zz_7951 = ($signed(_zz_7952) >>> _zz_370);
  assign _zz_7952 = _zz_7953;
  assign _zz_7953 = ($signed(_zz_7955) + $signed(_zz_366));
  assign _zz_7954 = ({8'd0,data_mid_17_real} <<< 8);
  assign _zz_7955 = {{8{_zz_7954[23]}}, _zz_7954};
  assign _zz_7956 = fixTo_442_dout;
  assign _zz_7957 = _zz_7958[31 : 0];
  assign _zz_7958 = _zz_7959;
  assign _zz_7959 = ($signed(_zz_7960) >>> _zz_370);
  assign _zz_7960 = _zz_7961;
  assign _zz_7961 = ($signed(_zz_7963) + $signed(_zz_367));
  assign _zz_7962 = ({8'd0,data_mid_17_imag} <<< 8);
  assign _zz_7963 = {{8{_zz_7962[23]}}, _zz_7962};
  assign _zz_7964 = fixTo_443_dout;
  assign _zz_7965 = ($signed(twiddle_factor_table_1_real) + $signed(twiddle_factor_table_1_imag));
  assign _zz_7966 = ($signed(_zz_373) - $signed(_zz_7967));
  assign _zz_7967 = ($signed(_zz_7968) * $signed(twiddle_factor_table_1_imag));
  assign _zz_7968 = ($signed(data_mid_22_real) + $signed(data_mid_22_imag));
  assign _zz_7969 = fixTo_444_dout;
  assign _zz_7970 = ($signed(_zz_373) + $signed(_zz_7971));
  assign _zz_7971 = ($signed(_zz_7972) * $signed(twiddle_factor_table_1_real));
  assign _zz_7972 = ($signed(data_mid_22_imag) - $signed(data_mid_22_real));
  assign _zz_7973 = fixTo_445_dout;
  assign _zz_7974 = _zz_7975[31 : 0];
  assign _zz_7975 = _zz_7976;
  assign _zz_7976 = ($signed(_zz_7977) >>> _zz_374);
  assign _zz_7977 = _zz_7978;
  assign _zz_7978 = ($signed(_zz_7980) - $signed(_zz_371));
  assign _zz_7979 = ({8'd0,data_mid_20_real} <<< 8);
  assign _zz_7980 = {{8{_zz_7979[23]}}, _zz_7979};
  assign _zz_7981 = fixTo_446_dout;
  assign _zz_7982 = _zz_7983[31 : 0];
  assign _zz_7983 = _zz_7984;
  assign _zz_7984 = ($signed(_zz_7985) >>> _zz_374);
  assign _zz_7985 = _zz_7986;
  assign _zz_7986 = ($signed(_zz_7988) - $signed(_zz_372));
  assign _zz_7987 = ({8'd0,data_mid_20_imag} <<< 8);
  assign _zz_7988 = {{8{_zz_7987[23]}}, _zz_7987};
  assign _zz_7989 = fixTo_447_dout;
  assign _zz_7990 = _zz_7991[31 : 0];
  assign _zz_7991 = _zz_7992;
  assign _zz_7992 = ($signed(_zz_7993) >>> _zz_375);
  assign _zz_7993 = _zz_7994;
  assign _zz_7994 = ($signed(_zz_7996) + $signed(_zz_371));
  assign _zz_7995 = ({8'd0,data_mid_20_real} <<< 8);
  assign _zz_7996 = {{8{_zz_7995[23]}}, _zz_7995};
  assign _zz_7997 = fixTo_448_dout;
  assign _zz_7998 = _zz_7999[31 : 0];
  assign _zz_7999 = _zz_8000;
  assign _zz_8000 = ($signed(_zz_8001) >>> _zz_375);
  assign _zz_8001 = _zz_8002;
  assign _zz_8002 = ($signed(_zz_8004) + $signed(_zz_372));
  assign _zz_8003 = ({8'd0,data_mid_20_imag} <<< 8);
  assign _zz_8004 = {{8{_zz_8003[23]}}, _zz_8003};
  assign _zz_8005 = fixTo_449_dout;
  assign _zz_8006 = ($signed(twiddle_factor_table_2_real) + $signed(twiddle_factor_table_2_imag));
  assign _zz_8007 = ($signed(_zz_378) - $signed(_zz_8008));
  assign _zz_8008 = ($signed(_zz_8009) * $signed(twiddle_factor_table_2_imag));
  assign _zz_8009 = ($signed(data_mid_23_real) + $signed(data_mid_23_imag));
  assign _zz_8010 = fixTo_450_dout;
  assign _zz_8011 = ($signed(_zz_378) + $signed(_zz_8012));
  assign _zz_8012 = ($signed(_zz_8013) * $signed(twiddle_factor_table_2_real));
  assign _zz_8013 = ($signed(data_mid_23_imag) - $signed(data_mid_23_real));
  assign _zz_8014 = fixTo_451_dout;
  assign _zz_8015 = _zz_8016[31 : 0];
  assign _zz_8016 = _zz_8017;
  assign _zz_8017 = ($signed(_zz_8018) >>> _zz_379);
  assign _zz_8018 = _zz_8019;
  assign _zz_8019 = ($signed(_zz_8021) - $signed(_zz_376));
  assign _zz_8020 = ({8'd0,data_mid_21_real} <<< 8);
  assign _zz_8021 = {{8{_zz_8020[23]}}, _zz_8020};
  assign _zz_8022 = fixTo_452_dout;
  assign _zz_8023 = _zz_8024[31 : 0];
  assign _zz_8024 = _zz_8025;
  assign _zz_8025 = ($signed(_zz_8026) >>> _zz_379);
  assign _zz_8026 = _zz_8027;
  assign _zz_8027 = ($signed(_zz_8029) - $signed(_zz_377));
  assign _zz_8028 = ({8'd0,data_mid_21_imag} <<< 8);
  assign _zz_8029 = {{8{_zz_8028[23]}}, _zz_8028};
  assign _zz_8030 = fixTo_453_dout;
  assign _zz_8031 = _zz_8032[31 : 0];
  assign _zz_8032 = _zz_8033;
  assign _zz_8033 = ($signed(_zz_8034) >>> _zz_380);
  assign _zz_8034 = _zz_8035;
  assign _zz_8035 = ($signed(_zz_8037) + $signed(_zz_376));
  assign _zz_8036 = ({8'd0,data_mid_21_real} <<< 8);
  assign _zz_8037 = {{8{_zz_8036[23]}}, _zz_8036};
  assign _zz_8038 = fixTo_454_dout;
  assign _zz_8039 = _zz_8040[31 : 0];
  assign _zz_8040 = _zz_8041;
  assign _zz_8041 = ($signed(_zz_8042) >>> _zz_380);
  assign _zz_8042 = _zz_8043;
  assign _zz_8043 = ($signed(_zz_8045) + $signed(_zz_377));
  assign _zz_8044 = ({8'd0,data_mid_21_imag} <<< 8);
  assign _zz_8045 = {{8{_zz_8044[23]}}, _zz_8044};
  assign _zz_8046 = fixTo_455_dout;
  assign _zz_8047 = ($signed(twiddle_factor_table_1_real) + $signed(twiddle_factor_table_1_imag));
  assign _zz_8048 = ($signed(_zz_383) - $signed(_zz_8049));
  assign _zz_8049 = ($signed(_zz_8050) * $signed(twiddle_factor_table_1_imag));
  assign _zz_8050 = ($signed(data_mid_26_real) + $signed(data_mid_26_imag));
  assign _zz_8051 = fixTo_456_dout;
  assign _zz_8052 = ($signed(_zz_383) + $signed(_zz_8053));
  assign _zz_8053 = ($signed(_zz_8054) * $signed(twiddle_factor_table_1_real));
  assign _zz_8054 = ($signed(data_mid_26_imag) - $signed(data_mid_26_real));
  assign _zz_8055 = fixTo_457_dout;
  assign _zz_8056 = _zz_8057[31 : 0];
  assign _zz_8057 = _zz_8058;
  assign _zz_8058 = ($signed(_zz_8059) >>> _zz_384);
  assign _zz_8059 = _zz_8060;
  assign _zz_8060 = ($signed(_zz_8062) - $signed(_zz_381));
  assign _zz_8061 = ({8'd0,data_mid_24_real} <<< 8);
  assign _zz_8062 = {{8{_zz_8061[23]}}, _zz_8061};
  assign _zz_8063 = fixTo_458_dout;
  assign _zz_8064 = _zz_8065[31 : 0];
  assign _zz_8065 = _zz_8066;
  assign _zz_8066 = ($signed(_zz_8067) >>> _zz_384);
  assign _zz_8067 = _zz_8068;
  assign _zz_8068 = ($signed(_zz_8070) - $signed(_zz_382));
  assign _zz_8069 = ({8'd0,data_mid_24_imag} <<< 8);
  assign _zz_8070 = {{8{_zz_8069[23]}}, _zz_8069};
  assign _zz_8071 = fixTo_459_dout;
  assign _zz_8072 = _zz_8073[31 : 0];
  assign _zz_8073 = _zz_8074;
  assign _zz_8074 = ($signed(_zz_8075) >>> _zz_385);
  assign _zz_8075 = _zz_8076;
  assign _zz_8076 = ($signed(_zz_8078) + $signed(_zz_381));
  assign _zz_8077 = ({8'd0,data_mid_24_real} <<< 8);
  assign _zz_8078 = {{8{_zz_8077[23]}}, _zz_8077};
  assign _zz_8079 = fixTo_460_dout;
  assign _zz_8080 = _zz_8081[31 : 0];
  assign _zz_8081 = _zz_8082;
  assign _zz_8082 = ($signed(_zz_8083) >>> _zz_385);
  assign _zz_8083 = _zz_8084;
  assign _zz_8084 = ($signed(_zz_8086) + $signed(_zz_382));
  assign _zz_8085 = ({8'd0,data_mid_24_imag} <<< 8);
  assign _zz_8086 = {{8{_zz_8085[23]}}, _zz_8085};
  assign _zz_8087 = fixTo_461_dout;
  assign _zz_8088 = ($signed(twiddle_factor_table_2_real) + $signed(twiddle_factor_table_2_imag));
  assign _zz_8089 = ($signed(_zz_388) - $signed(_zz_8090));
  assign _zz_8090 = ($signed(_zz_8091) * $signed(twiddle_factor_table_2_imag));
  assign _zz_8091 = ($signed(data_mid_27_real) + $signed(data_mid_27_imag));
  assign _zz_8092 = fixTo_462_dout;
  assign _zz_8093 = ($signed(_zz_388) + $signed(_zz_8094));
  assign _zz_8094 = ($signed(_zz_8095) * $signed(twiddle_factor_table_2_real));
  assign _zz_8095 = ($signed(data_mid_27_imag) - $signed(data_mid_27_real));
  assign _zz_8096 = fixTo_463_dout;
  assign _zz_8097 = _zz_8098[31 : 0];
  assign _zz_8098 = _zz_8099;
  assign _zz_8099 = ($signed(_zz_8100) >>> _zz_389);
  assign _zz_8100 = _zz_8101;
  assign _zz_8101 = ($signed(_zz_8103) - $signed(_zz_386));
  assign _zz_8102 = ({8'd0,data_mid_25_real} <<< 8);
  assign _zz_8103 = {{8{_zz_8102[23]}}, _zz_8102};
  assign _zz_8104 = fixTo_464_dout;
  assign _zz_8105 = _zz_8106[31 : 0];
  assign _zz_8106 = _zz_8107;
  assign _zz_8107 = ($signed(_zz_8108) >>> _zz_389);
  assign _zz_8108 = _zz_8109;
  assign _zz_8109 = ($signed(_zz_8111) - $signed(_zz_387));
  assign _zz_8110 = ({8'd0,data_mid_25_imag} <<< 8);
  assign _zz_8111 = {{8{_zz_8110[23]}}, _zz_8110};
  assign _zz_8112 = fixTo_465_dout;
  assign _zz_8113 = _zz_8114[31 : 0];
  assign _zz_8114 = _zz_8115;
  assign _zz_8115 = ($signed(_zz_8116) >>> _zz_390);
  assign _zz_8116 = _zz_8117;
  assign _zz_8117 = ($signed(_zz_8119) + $signed(_zz_386));
  assign _zz_8118 = ({8'd0,data_mid_25_real} <<< 8);
  assign _zz_8119 = {{8{_zz_8118[23]}}, _zz_8118};
  assign _zz_8120 = fixTo_466_dout;
  assign _zz_8121 = _zz_8122[31 : 0];
  assign _zz_8122 = _zz_8123;
  assign _zz_8123 = ($signed(_zz_8124) >>> _zz_390);
  assign _zz_8124 = _zz_8125;
  assign _zz_8125 = ($signed(_zz_8127) + $signed(_zz_387));
  assign _zz_8126 = ({8'd0,data_mid_25_imag} <<< 8);
  assign _zz_8127 = {{8{_zz_8126[23]}}, _zz_8126};
  assign _zz_8128 = fixTo_467_dout;
  assign _zz_8129 = ($signed(twiddle_factor_table_1_real) + $signed(twiddle_factor_table_1_imag));
  assign _zz_8130 = ($signed(_zz_393) - $signed(_zz_8131));
  assign _zz_8131 = ($signed(_zz_8132) * $signed(twiddle_factor_table_1_imag));
  assign _zz_8132 = ($signed(data_mid_30_real) + $signed(data_mid_30_imag));
  assign _zz_8133 = fixTo_468_dout;
  assign _zz_8134 = ($signed(_zz_393) + $signed(_zz_8135));
  assign _zz_8135 = ($signed(_zz_8136) * $signed(twiddle_factor_table_1_real));
  assign _zz_8136 = ($signed(data_mid_30_imag) - $signed(data_mid_30_real));
  assign _zz_8137 = fixTo_469_dout;
  assign _zz_8138 = _zz_8139[31 : 0];
  assign _zz_8139 = _zz_8140;
  assign _zz_8140 = ($signed(_zz_8141) >>> _zz_394);
  assign _zz_8141 = _zz_8142;
  assign _zz_8142 = ($signed(_zz_8144) - $signed(_zz_391));
  assign _zz_8143 = ({8'd0,data_mid_28_real} <<< 8);
  assign _zz_8144 = {{8{_zz_8143[23]}}, _zz_8143};
  assign _zz_8145 = fixTo_470_dout;
  assign _zz_8146 = _zz_8147[31 : 0];
  assign _zz_8147 = _zz_8148;
  assign _zz_8148 = ($signed(_zz_8149) >>> _zz_394);
  assign _zz_8149 = _zz_8150;
  assign _zz_8150 = ($signed(_zz_8152) - $signed(_zz_392));
  assign _zz_8151 = ({8'd0,data_mid_28_imag} <<< 8);
  assign _zz_8152 = {{8{_zz_8151[23]}}, _zz_8151};
  assign _zz_8153 = fixTo_471_dout;
  assign _zz_8154 = _zz_8155[31 : 0];
  assign _zz_8155 = _zz_8156;
  assign _zz_8156 = ($signed(_zz_8157) >>> _zz_395);
  assign _zz_8157 = _zz_8158;
  assign _zz_8158 = ($signed(_zz_8160) + $signed(_zz_391));
  assign _zz_8159 = ({8'd0,data_mid_28_real} <<< 8);
  assign _zz_8160 = {{8{_zz_8159[23]}}, _zz_8159};
  assign _zz_8161 = fixTo_472_dout;
  assign _zz_8162 = _zz_8163[31 : 0];
  assign _zz_8163 = _zz_8164;
  assign _zz_8164 = ($signed(_zz_8165) >>> _zz_395);
  assign _zz_8165 = _zz_8166;
  assign _zz_8166 = ($signed(_zz_8168) + $signed(_zz_392));
  assign _zz_8167 = ({8'd0,data_mid_28_imag} <<< 8);
  assign _zz_8168 = {{8{_zz_8167[23]}}, _zz_8167};
  assign _zz_8169 = fixTo_473_dout;
  assign _zz_8170 = ($signed(twiddle_factor_table_2_real) + $signed(twiddle_factor_table_2_imag));
  assign _zz_8171 = ($signed(_zz_398) - $signed(_zz_8172));
  assign _zz_8172 = ($signed(_zz_8173) * $signed(twiddle_factor_table_2_imag));
  assign _zz_8173 = ($signed(data_mid_31_real) + $signed(data_mid_31_imag));
  assign _zz_8174 = fixTo_474_dout;
  assign _zz_8175 = ($signed(_zz_398) + $signed(_zz_8176));
  assign _zz_8176 = ($signed(_zz_8177) * $signed(twiddle_factor_table_2_real));
  assign _zz_8177 = ($signed(data_mid_31_imag) - $signed(data_mid_31_real));
  assign _zz_8178 = fixTo_475_dout;
  assign _zz_8179 = _zz_8180[31 : 0];
  assign _zz_8180 = _zz_8181;
  assign _zz_8181 = ($signed(_zz_8182) >>> _zz_399);
  assign _zz_8182 = _zz_8183;
  assign _zz_8183 = ($signed(_zz_8185) - $signed(_zz_396));
  assign _zz_8184 = ({8'd0,data_mid_29_real} <<< 8);
  assign _zz_8185 = {{8{_zz_8184[23]}}, _zz_8184};
  assign _zz_8186 = fixTo_476_dout;
  assign _zz_8187 = _zz_8188[31 : 0];
  assign _zz_8188 = _zz_8189;
  assign _zz_8189 = ($signed(_zz_8190) >>> _zz_399);
  assign _zz_8190 = _zz_8191;
  assign _zz_8191 = ($signed(_zz_8193) - $signed(_zz_397));
  assign _zz_8192 = ({8'd0,data_mid_29_imag} <<< 8);
  assign _zz_8193 = {{8{_zz_8192[23]}}, _zz_8192};
  assign _zz_8194 = fixTo_477_dout;
  assign _zz_8195 = _zz_8196[31 : 0];
  assign _zz_8196 = _zz_8197;
  assign _zz_8197 = ($signed(_zz_8198) >>> _zz_400);
  assign _zz_8198 = _zz_8199;
  assign _zz_8199 = ($signed(_zz_8201) + $signed(_zz_396));
  assign _zz_8200 = ({8'd0,data_mid_29_real} <<< 8);
  assign _zz_8201 = {{8{_zz_8200[23]}}, _zz_8200};
  assign _zz_8202 = fixTo_478_dout;
  assign _zz_8203 = _zz_8204[31 : 0];
  assign _zz_8204 = _zz_8205;
  assign _zz_8205 = ($signed(_zz_8206) >>> _zz_400);
  assign _zz_8206 = _zz_8207;
  assign _zz_8207 = ($signed(_zz_8209) + $signed(_zz_397));
  assign _zz_8208 = ({8'd0,data_mid_29_imag} <<< 8);
  assign _zz_8209 = {{8{_zz_8208[23]}}, _zz_8208};
  assign _zz_8210 = fixTo_479_dout;
  assign _zz_8211 = ($signed(twiddle_factor_table_1_real) + $signed(twiddle_factor_table_1_imag));
  assign _zz_8212 = ($signed(_zz_403) - $signed(_zz_8213));
  assign _zz_8213 = ($signed(_zz_8214) * $signed(twiddle_factor_table_1_imag));
  assign _zz_8214 = ($signed(data_mid_34_real) + $signed(data_mid_34_imag));
  assign _zz_8215 = fixTo_480_dout;
  assign _zz_8216 = ($signed(_zz_403) + $signed(_zz_8217));
  assign _zz_8217 = ($signed(_zz_8218) * $signed(twiddle_factor_table_1_real));
  assign _zz_8218 = ($signed(data_mid_34_imag) - $signed(data_mid_34_real));
  assign _zz_8219 = fixTo_481_dout;
  assign _zz_8220 = _zz_8221[31 : 0];
  assign _zz_8221 = _zz_8222;
  assign _zz_8222 = ($signed(_zz_8223) >>> _zz_404);
  assign _zz_8223 = _zz_8224;
  assign _zz_8224 = ($signed(_zz_8226) - $signed(_zz_401));
  assign _zz_8225 = ({8'd0,data_mid_32_real} <<< 8);
  assign _zz_8226 = {{8{_zz_8225[23]}}, _zz_8225};
  assign _zz_8227 = fixTo_482_dout;
  assign _zz_8228 = _zz_8229[31 : 0];
  assign _zz_8229 = _zz_8230;
  assign _zz_8230 = ($signed(_zz_8231) >>> _zz_404);
  assign _zz_8231 = _zz_8232;
  assign _zz_8232 = ($signed(_zz_8234) - $signed(_zz_402));
  assign _zz_8233 = ({8'd0,data_mid_32_imag} <<< 8);
  assign _zz_8234 = {{8{_zz_8233[23]}}, _zz_8233};
  assign _zz_8235 = fixTo_483_dout;
  assign _zz_8236 = _zz_8237[31 : 0];
  assign _zz_8237 = _zz_8238;
  assign _zz_8238 = ($signed(_zz_8239) >>> _zz_405);
  assign _zz_8239 = _zz_8240;
  assign _zz_8240 = ($signed(_zz_8242) + $signed(_zz_401));
  assign _zz_8241 = ({8'd0,data_mid_32_real} <<< 8);
  assign _zz_8242 = {{8{_zz_8241[23]}}, _zz_8241};
  assign _zz_8243 = fixTo_484_dout;
  assign _zz_8244 = _zz_8245[31 : 0];
  assign _zz_8245 = _zz_8246;
  assign _zz_8246 = ($signed(_zz_8247) >>> _zz_405);
  assign _zz_8247 = _zz_8248;
  assign _zz_8248 = ($signed(_zz_8250) + $signed(_zz_402));
  assign _zz_8249 = ({8'd0,data_mid_32_imag} <<< 8);
  assign _zz_8250 = {{8{_zz_8249[23]}}, _zz_8249};
  assign _zz_8251 = fixTo_485_dout;
  assign _zz_8252 = ($signed(twiddle_factor_table_2_real) + $signed(twiddle_factor_table_2_imag));
  assign _zz_8253 = ($signed(_zz_408) - $signed(_zz_8254));
  assign _zz_8254 = ($signed(_zz_8255) * $signed(twiddle_factor_table_2_imag));
  assign _zz_8255 = ($signed(data_mid_35_real) + $signed(data_mid_35_imag));
  assign _zz_8256 = fixTo_486_dout;
  assign _zz_8257 = ($signed(_zz_408) + $signed(_zz_8258));
  assign _zz_8258 = ($signed(_zz_8259) * $signed(twiddle_factor_table_2_real));
  assign _zz_8259 = ($signed(data_mid_35_imag) - $signed(data_mid_35_real));
  assign _zz_8260 = fixTo_487_dout;
  assign _zz_8261 = _zz_8262[31 : 0];
  assign _zz_8262 = _zz_8263;
  assign _zz_8263 = ($signed(_zz_8264) >>> _zz_409);
  assign _zz_8264 = _zz_8265;
  assign _zz_8265 = ($signed(_zz_8267) - $signed(_zz_406));
  assign _zz_8266 = ({8'd0,data_mid_33_real} <<< 8);
  assign _zz_8267 = {{8{_zz_8266[23]}}, _zz_8266};
  assign _zz_8268 = fixTo_488_dout;
  assign _zz_8269 = _zz_8270[31 : 0];
  assign _zz_8270 = _zz_8271;
  assign _zz_8271 = ($signed(_zz_8272) >>> _zz_409);
  assign _zz_8272 = _zz_8273;
  assign _zz_8273 = ($signed(_zz_8275) - $signed(_zz_407));
  assign _zz_8274 = ({8'd0,data_mid_33_imag} <<< 8);
  assign _zz_8275 = {{8{_zz_8274[23]}}, _zz_8274};
  assign _zz_8276 = fixTo_489_dout;
  assign _zz_8277 = _zz_8278[31 : 0];
  assign _zz_8278 = _zz_8279;
  assign _zz_8279 = ($signed(_zz_8280) >>> _zz_410);
  assign _zz_8280 = _zz_8281;
  assign _zz_8281 = ($signed(_zz_8283) + $signed(_zz_406));
  assign _zz_8282 = ({8'd0,data_mid_33_real} <<< 8);
  assign _zz_8283 = {{8{_zz_8282[23]}}, _zz_8282};
  assign _zz_8284 = fixTo_490_dout;
  assign _zz_8285 = _zz_8286[31 : 0];
  assign _zz_8286 = _zz_8287;
  assign _zz_8287 = ($signed(_zz_8288) >>> _zz_410);
  assign _zz_8288 = _zz_8289;
  assign _zz_8289 = ($signed(_zz_8291) + $signed(_zz_407));
  assign _zz_8290 = ({8'd0,data_mid_33_imag} <<< 8);
  assign _zz_8291 = {{8{_zz_8290[23]}}, _zz_8290};
  assign _zz_8292 = fixTo_491_dout;
  assign _zz_8293 = ($signed(twiddle_factor_table_1_real) + $signed(twiddle_factor_table_1_imag));
  assign _zz_8294 = ($signed(_zz_413) - $signed(_zz_8295));
  assign _zz_8295 = ($signed(_zz_8296) * $signed(twiddle_factor_table_1_imag));
  assign _zz_8296 = ($signed(data_mid_38_real) + $signed(data_mid_38_imag));
  assign _zz_8297 = fixTo_492_dout;
  assign _zz_8298 = ($signed(_zz_413) + $signed(_zz_8299));
  assign _zz_8299 = ($signed(_zz_8300) * $signed(twiddle_factor_table_1_real));
  assign _zz_8300 = ($signed(data_mid_38_imag) - $signed(data_mid_38_real));
  assign _zz_8301 = fixTo_493_dout;
  assign _zz_8302 = _zz_8303[31 : 0];
  assign _zz_8303 = _zz_8304;
  assign _zz_8304 = ($signed(_zz_8305) >>> _zz_414);
  assign _zz_8305 = _zz_8306;
  assign _zz_8306 = ($signed(_zz_8308) - $signed(_zz_411));
  assign _zz_8307 = ({8'd0,data_mid_36_real} <<< 8);
  assign _zz_8308 = {{8{_zz_8307[23]}}, _zz_8307};
  assign _zz_8309 = fixTo_494_dout;
  assign _zz_8310 = _zz_8311[31 : 0];
  assign _zz_8311 = _zz_8312;
  assign _zz_8312 = ($signed(_zz_8313) >>> _zz_414);
  assign _zz_8313 = _zz_8314;
  assign _zz_8314 = ($signed(_zz_8316) - $signed(_zz_412));
  assign _zz_8315 = ({8'd0,data_mid_36_imag} <<< 8);
  assign _zz_8316 = {{8{_zz_8315[23]}}, _zz_8315};
  assign _zz_8317 = fixTo_495_dout;
  assign _zz_8318 = _zz_8319[31 : 0];
  assign _zz_8319 = _zz_8320;
  assign _zz_8320 = ($signed(_zz_8321) >>> _zz_415);
  assign _zz_8321 = _zz_8322;
  assign _zz_8322 = ($signed(_zz_8324) + $signed(_zz_411));
  assign _zz_8323 = ({8'd0,data_mid_36_real} <<< 8);
  assign _zz_8324 = {{8{_zz_8323[23]}}, _zz_8323};
  assign _zz_8325 = fixTo_496_dout;
  assign _zz_8326 = _zz_8327[31 : 0];
  assign _zz_8327 = _zz_8328;
  assign _zz_8328 = ($signed(_zz_8329) >>> _zz_415);
  assign _zz_8329 = _zz_8330;
  assign _zz_8330 = ($signed(_zz_8332) + $signed(_zz_412));
  assign _zz_8331 = ({8'd0,data_mid_36_imag} <<< 8);
  assign _zz_8332 = {{8{_zz_8331[23]}}, _zz_8331};
  assign _zz_8333 = fixTo_497_dout;
  assign _zz_8334 = ($signed(twiddle_factor_table_2_real) + $signed(twiddle_factor_table_2_imag));
  assign _zz_8335 = ($signed(_zz_418) - $signed(_zz_8336));
  assign _zz_8336 = ($signed(_zz_8337) * $signed(twiddle_factor_table_2_imag));
  assign _zz_8337 = ($signed(data_mid_39_real) + $signed(data_mid_39_imag));
  assign _zz_8338 = fixTo_498_dout;
  assign _zz_8339 = ($signed(_zz_418) + $signed(_zz_8340));
  assign _zz_8340 = ($signed(_zz_8341) * $signed(twiddle_factor_table_2_real));
  assign _zz_8341 = ($signed(data_mid_39_imag) - $signed(data_mid_39_real));
  assign _zz_8342 = fixTo_499_dout;
  assign _zz_8343 = _zz_8344[31 : 0];
  assign _zz_8344 = _zz_8345;
  assign _zz_8345 = ($signed(_zz_8346) >>> _zz_419);
  assign _zz_8346 = _zz_8347;
  assign _zz_8347 = ($signed(_zz_8349) - $signed(_zz_416));
  assign _zz_8348 = ({8'd0,data_mid_37_real} <<< 8);
  assign _zz_8349 = {{8{_zz_8348[23]}}, _zz_8348};
  assign _zz_8350 = fixTo_500_dout;
  assign _zz_8351 = _zz_8352[31 : 0];
  assign _zz_8352 = _zz_8353;
  assign _zz_8353 = ($signed(_zz_8354) >>> _zz_419);
  assign _zz_8354 = _zz_8355;
  assign _zz_8355 = ($signed(_zz_8357) - $signed(_zz_417));
  assign _zz_8356 = ({8'd0,data_mid_37_imag} <<< 8);
  assign _zz_8357 = {{8{_zz_8356[23]}}, _zz_8356};
  assign _zz_8358 = fixTo_501_dout;
  assign _zz_8359 = _zz_8360[31 : 0];
  assign _zz_8360 = _zz_8361;
  assign _zz_8361 = ($signed(_zz_8362) >>> _zz_420);
  assign _zz_8362 = _zz_8363;
  assign _zz_8363 = ($signed(_zz_8365) + $signed(_zz_416));
  assign _zz_8364 = ({8'd0,data_mid_37_real} <<< 8);
  assign _zz_8365 = {{8{_zz_8364[23]}}, _zz_8364};
  assign _zz_8366 = fixTo_502_dout;
  assign _zz_8367 = _zz_8368[31 : 0];
  assign _zz_8368 = _zz_8369;
  assign _zz_8369 = ($signed(_zz_8370) >>> _zz_420);
  assign _zz_8370 = _zz_8371;
  assign _zz_8371 = ($signed(_zz_8373) + $signed(_zz_417));
  assign _zz_8372 = ({8'd0,data_mid_37_imag} <<< 8);
  assign _zz_8373 = {{8{_zz_8372[23]}}, _zz_8372};
  assign _zz_8374 = fixTo_503_dout;
  assign _zz_8375 = ($signed(twiddle_factor_table_1_real) + $signed(twiddle_factor_table_1_imag));
  assign _zz_8376 = ($signed(_zz_423) - $signed(_zz_8377));
  assign _zz_8377 = ($signed(_zz_8378) * $signed(twiddle_factor_table_1_imag));
  assign _zz_8378 = ($signed(data_mid_42_real) + $signed(data_mid_42_imag));
  assign _zz_8379 = fixTo_504_dout;
  assign _zz_8380 = ($signed(_zz_423) + $signed(_zz_8381));
  assign _zz_8381 = ($signed(_zz_8382) * $signed(twiddle_factor_table_1_real));
  assign _zz_8382 = ($signed(data_mid_42_imag) - $signed(data_mid_42_real));
  assign _zz_8383 = fixTo_505_dout;
  assign _zz_8384 = _zz_8385[31 : 0];
  assign _zz_8385 = _zz_8386;
  assign _zz_8386 = ($signed(_zz_8387) >>> _zz_424);
  assign _zz_8387 = _zz_8388;
  assign _zz_8388 = ($signed(_zz_8390) - $signed(_zz_421));
  assign _zz_8389 = ({8'd0,data_mid_40_real} <<< 8);
  assign _zz_8390 = {{8{_zz_8389[23]}}, _zz_8389};
  assign _zz_8391 = fixTo_506_dout;
  assign _zz_8392 = _zz_8393[31 : 0];
  assign _zz_8393 = _zz_8394;
  assign _zz_8394 = ($signed(_zz_8395) >>> _zz_424);
  assign _zz_8395 = _zz_8396;
  assign _zz_8396 = ($signed(_zz_8398) - $signed(_zz_422));
  assign _zz_8397 = ({8'd0,data_mid_40_imag} <<< 8);
  assign _zz_8398 = {{8{_zz_8397[23]}}, _zz_8397};
  assign _zz_8399 = fixTo_507_dout;
  assign _zz_8400 = _zz_8401[31 : 0];
  assign _zz_8401 = _zz_8402;
  assign _zz_8402 = ($signed(_zz_8403) >>> _zz_425);
  assign _zz_8403 = _zz_8404;
  assign _zz_8404 = ($signed(_zz_8406) + $signed(_zz_421));
  assign _zz_8405 = ({8'd0,data_mid_40_real} <<< 8);
  assign _zz_8406 = {{8{_zz_8405[23]}}, _zz_8405};
  assign _zz_8407 = fixTo_508_dout;
  assign _zz_8408 = _zz_8409[31 : 0];
  assign _zz_8409 = _zz_8410;
  assign _zz_8410 = ($signed(_zz_8411) >>> _zz_425);
  assign _zz_8411 = _zz_8412;
  assign _zz_8412 = ($signed(_zz_8414) + $signed(_zz_422));
  assign _zz_8413 = ({8'd0,data_mid_40_imag} <<< 8);
  assign _zz_8414 = {{8{_zz_8413[23]}}, _zz_8413};
  assign _zz_8415 = fixTo_509_dout;
  assign _zz_8416 = ($signed(twiddle_factor_table_2_real) + $signed(twiddle_factor_table_2_imag));
  assign _zz_8417 = ($signed(_zz_428) - $signed(_zz_8418));
  assign _zz_8418 = ($signed(_zz_8419) * $signed(twiddle_factor_table_2_imag));
  assign _zz_8419 = ($signed(data_mid_43_real) + $signed(data_mid_43_imag));
  assign _zz_8420 = fixTo_510_dout;
  assign _zz_8421 = ($signed(_zz_428) + $signed(_zz_8422));
  assign _zz_8422 = ($signed(_zz_8423) * $signed(twiddle_factor_table_2_real));
  assign _zz_8423 = ($signed(data_mid_43_imag) - $signed(data_mid_43_real));
  assign _zz_8424 = fixTo_511_dout;
  assign _zz_8425 = _zz_8426[31 : 0];
  assign _zz_8426 = _zz_8427;
  assign _zz_8427 = ($signed(_zz_8428) >>> _zz_429);
  assign _zz_8428 = _zz_8429;
  assign _zz_8429 = ($signed(_zz_8431) - $signed(_zz_426));
  assign _zz_8430 = ({8'd0,data_mid_41_real} <<< 8);
  assign _zz_8431 = {{8{_zz_8430[23]}}, _zz_8430};
  assign _zz_8432 = fixTo_512_dout;
  assign _zz_8433 = _zz_8434[31 : 0];
  assign _zz_8434 = _zz_8435;
  assign _zz_8435 = ($signed(_zz_8436) >>> _zz_429);
  assign _zz_8436 = _zz_8437;
  assign _zz_8437 = ($signed(_zz_8439) - $signed(_zz_427));
  assign _zz_8438 = ({8'd0,data_mid_41_imag} <<< 8);
  assign _zz_8439 = {{8{_zz_8438[23]}}, _zz_8438};
  assign _zz_8440 = fixTo_513_dout;
  assign _zz_8441 = _zz_8442[31 : 0];
  assign _zz_8442 = _zz_8443;
  assign _zz_8443 = ($signed(_zz_8444) >>> _zz_430);
  assign _zz_8444 = _zz_8445;
  assign _zz_8445 = ($signed(_zz_8447) + $signed(_zz_426));
  assign _zz_8446 = ({8'd0,data_mid_41_real} <<< 8);
  assign _zz_8447 = {{8{_zz_8446[23]}}, _zz_8446};
  assign _zz_8448 = fixTo_514_dout;
  assign _zz_8449 = _zz_8450[31 : 0];
  assign _zz_8450 = _zz_8451;
  assign _zz_8451 = ($signed(_zz_8452) >>> _zz_430);
  assign _zz_8452 = _zz_8453;
  assign _zz_8453 = ($signed(_zz_8455) + $signed(_zz_427));
  assign _zz_8454 = ({8'd0,data_mid_41_imag} <<< 8);
  assign _zz_8455 = {{8{_zz_8454[23]}}, _zz_8454};
  assign _zz_8456 = fixTo_515_dout;
  assign _zz_8457 = ($signed(twiddle_factor_table_1_real) + $signed(twiddle_factor_table_1_imag));
  assign _zz_8458 = ($signed(_zz_433) - $signed(_zz_8459));
  assign _zz_8459 = ($signed(_zz_8460) * $signed(twiddle_factor_table_1_imag));
  assign _zz_8460 = ($signed(data_mid_46_real) + $signed(data_mid_46_imag));
  assign _zz_8461 = fixTo_516_dout;
  assign _zz_8462 = ($signed(_zz_433) + $signed(_zz_8463));
  assign _zz_8463 = ($signed(_zz_8464) * $signed(twiddle_factor_table_1_real));
  assign _zz_8464 = ($signed(data_mid_46_imag) - $signed(data_mid_46_real));
  assign _zz_8465 = fixTo_517_dout;
  assign _zz_8466 = _zz_8467[31 : 0];
  assign _zz_8467 = _zz_8468;
  assign _zz_8468 = ($signed(_zz_8469) >>> _zz_434);
  assign _zz_8469 = _zz_8470;
  assign _zz_8470 = ($signed(_zz_8472) - $signed(_zz_431));
  assign _zz_8471 = ({8'd0,data_mid_44_real} <<< 8);
  assign _zz_8472 = {{8{_zz_8471[23]}}, _zz_8471};
  assign _zz_8473 = fixTo_518_dout;
  assign _zz_8474 = _zz_8475[31 : 0];
  assign _zz_8475 = _zz_8476;
  assign _zz_8476 = ($signed(_zz_8477) >>> _zz_434);
  assign _zz_8477 = _zz_8478;
  assign _zz_8478 = ($signed(_zz_8480) - $signed(_zz_432));
  assign _zz_8479 = ({8'd0,data_mid_44_imag} <<< 8);
  assign _zz_8480 = {{8{_zz_8479[23]}}, _zz_8479};
  assign _zz_8481 = fixTo_519_dout;
  assign _zz_8482 = _zz_8483[31 : 0];
  assign _zz_8483 = _zz_8484;
  assign _zz_8484 = ($signed(_zz_8485) >>> _zz_435);
  assign _zz_8485 = _zz_8486;
  assign _zz_8486 = ($signed(_zz_8488) + $signed(_zz_431));
  assign _zz_8487 = ({8'd0,data_mid_44_real} <<< 8);
  assign _zz_8488 = {{8{_zz_8487[23]}}, _zz_8487};
  assign _zz_8489 = fixTo_520_dout;
  assign _zz_8490 = _zz_8491[31 : 0];
  assign _zz_8491 = _zz_8492;
  assign _zz_8492 = ($signed(_zz_8493) >>> _zz_435);
  assign _zz_8493 = _zz_8494;
  assign _zz_8494 = ($signed(_zz_8496) + $signed(_zz_432));
  assign _zz_8495 = ({8'd0,data_mid_44_imag} <<< 8);
  assign _zz_8496 = {{8{_zz_8495[23]}}, _zz_8495};
  assign _zz_8497 = fixTo_521_dout;
  assign _zz_8498 = ($signed(twiddle_factor_table_2_real) + $signed(twiddle_factor_table_2_imag));
  assign _zz_8499 = ($signed(_zz_438) - $signed(_zz_8500));
  assign _zz_8500 = ($signed(_zz_8501) * $signed(twiddle_factor_table_2_imag));
  assign _zz_8501 = ($signed(data_mid_47_real) + $signed(data_mid_47_imag));
  assign _zz_8502 = fixTo_522_dout;
  assign _zz_8503 = ($signed(_zz_438) + $signed(_zz_8504));
  assign _zz_8504 = ($signed(_zz_8505) * $signed(twiddle_factor_table_2_real));
  assign _zz_8505 = ($signed(data_mid_47_imag) - $signed(data_mid_47_real));
  assign _zz_8506 = fixTo_523_dout;
  assign _zz_8507 = _zz_8508[31 : 0];
  assign _zz_8508 = _zz_8509;
  assign _zz_8509 = ($signed(_zz_8510) >>> _zz_439);
  assign _zz_8510 = _zz_8511;
  assign _zz_8511 = ($signed(_zz_8513) - $signed(_zz_436));
  assign _zz_8512 = ({8'd0,data_mid_45_real} <<< 8);
  assign _zz_8513 = {{8{_zz_8512[23]}}, _zz_8512};
  assign _zz_8514 = fixTo_524_dout;
  assign _zz_8515 = _zz_8516[31 : 0];
  assign _zz_8516 = _zz_8517;
  assign _zz_8517 = ($signed(_zz_8518) >>> _zz_439);
  assign _zz_8518 = _zz_8519;
  assign _zz_8519 = ($signed(_zz_8521) - $signed(_zz_437));
  assign _zz_8520 = ({8'd0,data_mid_45_imag} <<< 8);
  assign _zz_8521 = {{8{_zz_8520[23]}}, _zz_8520};
  assign _zz_8522 = fixTo_525_dout;
  assign _zz_8523 = _zz_8524[31 : 0];
  assign _zz_8524 = _zz_8525;
  assign _zz_8525 = ($signed(_zz_8526) >>> _zz_440);
  assign _zz_8526 = _zz_8527;
  assign _zz_8527 = ($signed(_zz_8529) + $signed(_zz_436));
  assign _zz_8528 = ({8'd0,data_mid_45_real} <<< 8);
  assign _zz_8529 = {{8{_zz_8528[23]}}, _zz_8528};
  assign _zz_8530 = fixTo_526_dout;
  assign _zz_8531 = _zz_8532[31 : 0];
  assign _zz_8532 = _zz_8533;
  assign _zz_8533 = ($signed(_zz_8534) >>> _zz_440);
  assign _zz_8534 = _zz_8535;
  assign _zz_8535 = ($signed(_zz_8537) + $signed(_zz_437));
  assign _zz_8536 = ({8'd0,data_mid_45_imag} <<< 8);
  assign _zz_8537 = {{8{_zz_8536[23]}}, _zz_8536};
  assign _zz_8538 = fixTo_527_dout;
  assign _zz_8539 = ($signed(twiddle_factor_table_1_real) + $signed(twiddle_factor_table_1_imag));
  assign _zz_8540 = ($signed(_zz_443) - $signed(_zz_8541));
  assign _zz_8541 = ($signed(_zz_8542) * $signed(twiddle_factor_table_1_imag));
  assign _zz_8542 = ($signed(data_mid_50_real) + $signed(data_mid_50_imag));
  assign _zz_8543 = fixTo_528_dout;
  assign _zz_8544 = ($signed(_zz_443) + $signed(_zz_8545));
  assign _zz_8545 = ($signed(_zz_8546) * $signed(twiddle_factor_table_1_real));
  assign _zz_8546 = ($signed(data_mid_50_imag) - $signed(data_mid_50_real));
  assign _zz_8547 = fixTo_529_dout;
  assign _zz_8548 = _zz_8549[31 : 0];
  assign _zz_8549 = _zz_8550;
  assign _zz_8550 = ($signed(_zz_8551) >>> _zz_444);
  assign _zz_8551 = _zz_8552;
  assign _zz_8552 = ($signed(_zz_8554) - $signed(_zz_441));
  assign _zz_8553 = ({8'd0,data_mid_48_real} <<< 8);
  assign _zz_8554 = {{8{_zz_8553[23]}}, _zz_8553};
  assign _zz_8555 = fixTo_530_dout;
  assign _zz_8556 = _zz_8557[31 : 0];
  assign _zz_8557 = _zz_8558;
  assign _zz_8558 = ($signed(_zz_8559) >>> _zz_444);
  assign _zz_8559 = _zz_8560;
  assign _zz_8560 = ($signed(_zz_8562) - $signed(_zz_442));
  assign _zz_8561 = ({8'd0,data_mid_48_imag} <<< 8);
  assign _zz_8562 = {{8{_zz_8561[23]}}, _zz_8561};
  assign _zz_8563 = fixTo_531_dout;
  assign _zz_8564 = _zz_8565[31 : 0];
  assign _zz_8565 = _zz_8566;
  assign _zz_8566 = ($signed(_zz_8567) >>> _zz_445);
  assign _zz_8567 = _zz_8568;
  assign _zz_8568 = ($signed(_zz_8570) + $signed(_zz_441));
  assign _zz_8569 = ({8'd0,data_mid_48_real} <<< 8);
  assign _zz_8570 = {{8{_zz_8569[23]}}, _zz_8569};
  assign _zz_8571 = fixTo_532_dout;
  assign _zz_8572 = _zz_8573[31 : 0];
  assign _zz_8573 = _zz_8574;
  assign _zz_8574 = ($signed(_zz_8575) >>> _zz_445);
  assign _zz_8575 = _zz_8576;
  assign _zz_8576 = ($signed(_zz_8578) + $signed(_zz_442));
  assign _zz_8577 = ({8'd0,data_mid_48_imag} <<< 8);
  assign _zz_8578 = {{8{_zz_8577[23]}}, _zz_8577};
  assign _zz_8579 = fixTo_533_dout;
  assign _zz_8580 = ($signed(twiddle_factor_table_2_real) + $signed(twiddle_factor_table_2_imag));
  assign _zz_8581 = ($signed(_zz_448) - $signed(_zz_8582));
  assign _zz_8582 = ($signed(_zz_8583) * $signed(twiddle_factor_table_2_imag));
  assign _zz_8583 = ($signed(data_mid_51_real) + $signed(data_mid_51_imag));
  assign _zz_8584 = fixTo_534_dout;
  assign _zz_8585 = ($signed(_zz_448) + $signed(_zz_8586));
  assign _zz_8586 = ($signed(_zz_8587) * $signed(twiddle_factor_table_2_real));
  assign _zz_8587 = ($signed(data_mid_51_imag) - $signed(data_mid_51_real));
  assign _zz_8588 = fixTo_535_dout;
  assign _zz_8589 = _zz_8590[31 : 0];
  assign _zz_8590 = _zz_8591;
  assign _zz_8591 = ($signed(_zz_8592) >>> _zz_449);
  assign _zz_8592 = _zz_8593;
  assign _zz_8593 = ($signed(_zz_8595) - $signed(_zz_446));
  assign _zz_8594 = ({8'd0,data_mid_49_real} <<< 8);
  assign _zz_8595 = {{8{_zz_8594[23]}}, _zz_8594};
  assign _zz_8596 = fixTo_536_dout;
  assign _zz_8597 = _zz_8598[31 : 0];
  assign _zz_8598 = _zz_8599;
  assign _zz_8599 = ($signed(_zz_8600) >>> _zz_449);
  assign _zz_8600 = _zz_8601;
  assign _zz_8601 = ($signed(_zz_8603) - $signed(_zz_447));
  assign _zz_8602 = ({8'd0,data_mid_49_imag} <<< 8);
  assign _zz_8603 = {{8{_zz_8602[23]}}, _zz_8602};
  assign _zz_8604 = fixTo_537_dout;
  assign _zz_8605 = _zz_8606[31 : 0];
  assign _zz_8606 = _zz_8607;
  assign _zz_8607 = ($signed(_zz_8608) >>> _zz_450);
  assign _zz_8608 = _zz_8609;
  assign _zz_8609 = ($signed(_zz_8611) + $signed(_zz_446));
  assign _zz_8610 = ({8'd0,data_mid_49_real} <<< 8);
  assign _zz_8611 = {{8{_zz_8610[23]}}, _zz_8610};
  assign _zz_8612 = fixTo_538_dout;
  assign _zz_8613 = _zz_8614[31 : 0];
  assign _zz_8614 = _zz_8615;
  assign _zz_8615 = ($signed(_zz_8616) >>> _zz_450);
  assign _zz_8616 = _zz_8617;
  assign _zz_8617 = ($signed(_zz_8619) + $signed(_zz_447));
  assign _zz_8618 = ({8'd0,data_mid_49_imag} <<< 8);
  assign _zz_8619 = {{8{_zz_8618[23]}}, _zz_8618};
  assign _zz_8620 = fixTo_539_dout;
  assign _zz_8621 = ($signed(twiddle_factor_table_1_real) + $signed(twiddle_factor_table_1_imag));
  assign _zz_8622 = ($signed(_zz_453) - $signed(_zz_8623));
  assign _zz_8623 = ($signed(_zz_8624) * $signed(twiddle_factor_table_1_imag));
  assign _zz_8624 = ($signed(data_mid_54_real) + $signed(data_mid_54_imag));
  assign _zz_8625 = fixTo_540_dout;
  assign _zz_8626 = ($signed(_zz_453) + $signed(_zz_8627));
  assign _zz_8627 = ($signed(_zz_8628) * $signed(twiddle_factor_table_1_real));
  assign _zz_8628 = ($signed(data_mid_54_imag) - $signed(data_mid_54_real));
  assign _zz_8629 = fixTo_541_dout;
  assign _zz_8630 = _zz_8631[31 : 0];
  assign _zz_8631 = _zz_8632;
  assign _zz_8632 = ($signed(_zz_8633) >>> _zz_454);
  assign _zz_8633 = _zz_8634;
  assign _zz_8634 = ($signed(_zz_8636) - $signed(_zz_451));
  assign _zz_8635 = ({8'd0,data_mid_52_real} <<< 8);
  assign _zz_8636 = {{8{_zz_8635[23]}}, _zz_8635};
  assign _zz_8637 = fixTo_542_dout;
  assign _zz_8638 = _zz_8639[31 : 0];
  assign _zz_8639 = _zz_8640;
  assign _zz_8640 = ($signed(_zz_8641) >>> _zz_454);
  assign _zz_8641 = _zz_8642;
  assign _zz_8642 = ($signed(_zz_8644) - $signed(_zz_452));
  assign _zz_8643 = ({8'd0,data_mid_52_imag} <<< 8);
  assign _zz_8644 = {{8{_zz_8643[23]}}, _zz_8643};
  assign _zz_8645 = fixTo_543_dout;
  assign _zz_8646 = _zz_8647[31 : 0];
  assign _zz_8647 = _zz_8648;
  assign _zz_8648 = ($signed(_zz_8649) >>> _zz_455);
  assign _zz_8649 = _zz_8650;
  assign _zz_8650 = ($signed(_zz_8652) + $signed(_zz_451));
  assign _zz_8651 = ({8'd0,data_mid_52_real} <<< 8);
  assign _zz_8652 = {{8{_zz_8651[23]}}, _zz_8651};
  assign _zz_8653 = fixTo_544_dout;
  assign _zz_8654 = _zz_8655[31 : 0];
  assign _zz_8655 = _zz_8656;
  assign _zz_8656 = ($signed(_zz_8657) >>> _zz_455);
  assign _zz_8657 = _zz_8658;
  assign _zz_8658 = ($signed(_zz_8660) + $signed(_zz_452));
  assign _zz_8659 = ({8'd0,data_mid_52_imag} <<< 8);
  assign _zz_8660 = {{8{_zz_8659[23]}}, _zz_8659};
  assign _zz_8661 = fixTo_545_dout;
  assign _zz_8662 = ($signed(twiddle_factor_table_2_real) + $signed(twiddle_factor_table_2_imag));
  assign _zz_8663 = ($signed(_zz_458) - $signed(_zz_8664));
  assign _zz_8664 = ($signed(_zz_8665) * $signed(twiddle_factor_table_2_imag));
  assign _zz_8665 = ($signed(data_mid_55_real) + $signed(data_mid_55_imag));
  assign _zz_8666 = fixTo_546_dout;
  assign _zz_8667 = ($signed(_zz_458) + $signed(_zz_8668));
  assign _zz_8668 = ($signed(_zz_8669) * $signed(twiddle_factor_table_2_real));
  assign _zz_8669 = ($signed(data_mid_55_imag) - $signed(data_mid_55_real));
  assign _zz_8670 = fixTo_547_dout;
  assign _zz_8671 = _zz_8672[31 : 0];
  assign _zz_8672 = _zz_8673;
  assign _zz_8673 = ($signed(_zz_8674) >>> _zz_459);
  assign _zz_8674 = _zz_8675;
  assign _zz_8675 = ($signed(_zz_8677) - $signed(_zz_456));
  assign _zz_8676 = ({8'd0,data_mid_53_real} <<< 8);
  assign _zz_8677 = {{8{_zz_8676[23]}}, _zz_8676};
  assign _zz_8678 = fixTo_548_dout;
  assign _zz_8679 = _zz_8680[31 : 0];
  assign _zz_8680 = _zz_8681;
  assign _zz_8681 = ($signed(_zz_8682) >>> _zz_459);
  assign _zz_8682 = _zz_8683;
  assign _zz_8683 = ($signed(_zz_8685) - $signed(_zz_457));
  assign _zz_8684 = ({8'd0,data_mid_53_imag} <<< 8);
  assign _zz_8685 = {{8{_zz_8684[23]}}, _zz_8684};
  assign _zz_8686 = fixTo_549_dout;
  assign _zz_8687 = _zz_8688[31 : 0];
  assign _zz_8688 = _zz_8689;
  assign _zz_8689 = ($signed(_zz_8690) >>> _zz_460);
  assign _zz_8690 = _zz_8691;
  assign _zz_8691 = ($signed(_zz_8693) + $signed(_zz_456));
  assign _zz_8692 = ({8'd0,data_mid_53_real} <<< 8);
  assign _zz_8693 = {{8{_zz_8692[23]}}, _zz_8692};
  assign _zz_8694 = fixTo_550_dout;
  assign _zz_8695 = _zz_8696[31 : 0];
  assign _zz_8696 = _zz_8697;
  assign _zz_8697 = ($signed(_zz_8698) >>> _zz_460);
  assign _zz_8698 = _zz_8699;
  assign _zz_8699 = ($signed(_zz_8701) + $signed(_zz_457));
  assign _zz_8700 = ({8'd0,data_mid_53_imag} <<< 8);
  assign _zz_8701 = {{8{_zz_8700[23]}}, _zz_8700};
  assign _zz_8702 = fixTo_551_dout;
  assign _zz_8703 = ($signed(twiddle_factor_table_1_real) + $signed(twiddle_factor_table_1_imag));
  assign _zz_8704 = ($signed(_zz_463) - $signed(_zz_8705));
  assign _zz_8705 = ($signed(_zz_8706) * $signed(twiddle_factor_table_1_imag));
  assign _zz_8706 = ($signed(data_mid_58_real) + $signed(data_mid_58_imag));
  assign _zz_8707 = fixTo_552_dout;
  assign _zz_8708 = ($signed(_zz_463) + $signed(_zz_8709));
  assign _zz_8709 = ($signed(_zz_8710) * $signed(twiddle_factor_table_1_real));
  assign _zz_8710 = ($signed(data_mid_58_imag) - $signed(data_mid_58_real));
  assign _zz_8711 = fixTo_553_dout;
  assign _zz_8712 = _zz_8713[31 : 0];
  assign _zz_8713 = _zz_8714;
  assign _zz_8714 = ($signed(_zz_8715) >>> _zz_464);
  assign _zz_8715 = _zz_8716;
  assign _zz_8716 = ($signed(_zz_8718) - $signed(_zz_461));
  assign _zz_8717 = ({8'd0,data_mid_56_real} <<< 8);
  assign _zz_8718 = {{8{_zz_8717[23]}}, _zz_8717};
  assign _zz_8719 = fixTo_554_dout;
  assign _zz_8720 = _zz_8721[31 : 0];
  assign _zz_8721 = _zz_8722;
  assign _zz_8722 = ($signed(_zz_8723) >>> _zz_464);
  assign _zz_8723 = _zz_8724;
  assign _zz_8724 = ($signed(_zz_8726) - $signed(_zz_462));
  assign _zz_8725 = ({8'd0,data_mid_56_imag} <<< 8);
  assign _zz_8726 = {{8{_zz_8725[23]}}, _zz_8725};
  assign _zz_8727 = fixTo_555_dout;
  assign _zz_8728 = _zz_8729[31 : 0];
  assign _zz_8729 = _zz_8730;
  assign _zz_8730 = ($signed(_zz_8731) >>> _zz_465);
  assign _zz_8731 = _zz_8732;
  assign _zz_8732 = ($signed(_zz_8734) + $signed(_zz_461));
  assign _zz_8733 = ({8'd0,data_mid_56_real} <<< 8);
  assign _zz_8734 = {{8{_zz_8733[23]}}, _zz_8733};
  assign _zz_8735 = fixTo_556_dout;
  assign _zz_8736 = _zz_8737[31 : 0];
  assign _zz_8737 = _zz_8738;
  assign _zz_8738 = ($signed(_zz_8739) >>> _zz_465);
  assign _zz_8739 = _zz_8740;
  assign _zz_8740 = ($signed(_zz_8742) + $signed(_zz_462));
  assign _zz_8741 = ({8'd0,data_mid_56_imag} <<< 8);
  assign _zz_8742 = {{8{_zz_8741[23]}}, _zz_8741};
  assign _zz_8743 = fixTo_557_dout;
  assign _zz_8744 = ($signed(twiddle_factor_table_2_real) + $signed(twiddle_factor_table_2_imag));
  assign _zz_8745 = ($signed(_zz_468) - $signed(_zz_8746));
  assign _zz_8746 = ($signed(_zz_8747) * $signed(twiddle_factor_table_2_imag));
  assign _zz_8747 = ($signed(data_mid_59_real) + $signed(data_mid_59_imag));
  assign _zz_8748 = fixTo_558_dout;
  assign _zz_8749 = ($signed(_zz_468) + $signed(_zz_8750));
  assign _zz_8750 = ($signed(_zz_8751) * $signed(twiddle_factor_table_2_real));
  assign _zz_8751 = ($signed(data_mid_59_imag) - $signed(data_mid_59_real));
  assign _zz_8752 = fixTo_559_dout;
  assign _zz_8753 = _zz_8754[31 : 0];
  assign _zz_8754 = _zz_8755;
  assign _zz_8755 = ($signed(_zz_8756) >>> _zz_469);
  assign _zz_8756 = _zz_8757;
  assign _zz_8757 = ($signed(_zz_8759) - $signed(_zz_466));
  assign _zz_8758 = ({8'd0,data_mid_57_real} <<< 8);
  assign _zz_8759 = {{8{_zz_8758[23]}}, _zz_8758};
  assign _zz_8760 = fixTo_560_dout;
  assign _zz_8761 = _zz_8762[31 : 0];
  assign _zz_8762 = _zz_8763;
  assign _zz_8763 = ($signed(_zz_8764) >>> _zz_469);
  assign _zz_8764 = _zz_8765;
  assign _zz_8765 = ($signed(_zz_8767) - $signed(_zz_467));
  assign _zz_8766 = ({8'd0,data_mid_57_imag} <<< 8);
  assign _zz_8767 = {{8{_zz_8766[23]}}, _zz_8766};
  assign _zz_8768 = fixTo_561_dout;
  assign _zz_8769 = _zz_8770[31 : 0];
  assign _zz_8770 = _zz_8771;
  assign _zz_8771 = ($signed(_zz_8772) >>> _zz_470);
  assign _zz_8772 = _zz_8773;
  assign _zz_8773 = ($signed(_zz_8775) + $signed(_zz_466));
  assign _zz_8774 = ({8'd0,data_mid_57_real} <<< 8);
  assign _zz_8775 = {{8{_zz_8774[23]}}, _zz_8774};
  assign _zz_8776 = fixTo_562_dout;
  assign _zz_8777 = _zz_8778[31 : 0];
  assign _zz_8778 = _zz_8779;
  assign _zz_8779 = ($signed(_zz_8780) >>> _zz_470);
  assign _zz_8780 = _zz_8781;
  assign _zz_8781 = ($signed(_zz_8783) + $signed(_zz_467));
  assign _zz_8782 = ({8'd0,data_mid_57_imag} <<< 8);
  assign _zz_8783 = {{8{_zz_8782[23]}}, _zz_8782};
  assign _zz_8784 = fixTo_563_dout;
  assign _zz_8785 = ($signed(twiddle_factor_table_1_real) + $signed(twiddle_factor_table_1_imag));
  assign _zz_8786 = ($signed(_zz_473) - $signed(_zz_8787));
  assign _zz_8787 = ($signed(_zz_8788) * $signed(twiddle_factor_table_1_imag));
  assign _zz_8788 = ($signed(data_mid_62_real) + $signed(data_mid_62_imag));
  assign _zz_8789 = fixTo_564_dout;
  assign _zz_8790 = ($signed(_zz_473) + $signed(_zz_8791));
  assign _zz_8791 = ($signed(_zz_8792) * $signed(twiddle_factor_table_1_real));
  assign _zz_8792 = ($signed(data_mid_62_imag) - $signed(data_mid_62_real));
  assign _zz_8793 = fixTo_565_dout;
  assign _zz_8794 = _zz_8795[31 : 0];
  assign _zz_8795 = _zz_8796;
  assign _zz_8796 = ($signed(_zz_8797) >>> _zz_474);
  assign _zz_8797 = _zz_8798;
  assign _zz_8798 = ($signed(_zz_8800) - $signed(_zz_471));
  assign _zz_8799 = ({8'd0,data_mid_60_real} <<< 8);
  assign _zz_8800 = {{8{_zz_8799[23]}}, _zz_8799};
  assign _zz_8801 = fixTo_566_dout;
  assign _zz_8802 = _zz_8803[31 : 0];
  assign _zz_8803 = _zz_8804;
  assign _zz_8804 = ($signed(_zz_8805) >>> _zz_474);
  assign _zz_8805 = _zz_8806;
  assign _zz_8806 = ($signed(_zz_8808) - $signed(_zz_472));
  assign _zz_8807 = ({8'd0,data_mid_60_imag} <<< 8);
  assign _zz_8808 = {{8{_zz_8807[23]}}, _zz_8807};
  assign _zz_8809 = fixTo_567_dout;
  assign _zz_8810 = _zz_8811[31 : 0];
  assign _zz_8811 = _zz_8812;
  assign _zz_8812 = ($signed(_zz_8813) >>> _zz_475);
  assign _zz_8813 = _zz_8814;
  assign _zz_8814 = ($signed(_zz_8816) + $signed(_zz_471));
  assign _zz_8815 = ({8'd0,data_mid_60_real} <<< 8);
  assign _zz_8816 = {{8{_zz_8815[23]}}, _zz_8815};
  assign _zz_8817 = fixTo_568_dout;
  assign _zz_8818 = _zz_8819[31 : 0];
  assign _zz_8819 = _zz_8820;
  assign _zz_8820 = ($signed(_zz_8821) >>> _zz_475);
  assign _zz_8821 = _zz_8822;
  assign _zz_8822 = ($signed(_zz_8824) + $signed(_zz_472));
  assign _zz_8823 = ({8'd0,data_mid_60_imag} <<< 8);
  assign _zz_8824 = {{8{_zz_8823[23]}}, _zz_8823};
  assign _zz_8825 = fixTo_569_dout;
  assign _zz_8826 = ($signed(twiddle_factor_table_2_real) + $signed(twiddle_factor_table_2_imag));
  assign _zz_8827 = ($signed(_zz_478) - $signed(_zz_8828));
  assign _zz_8828 = ($signed(_zz_8829) * $signed(twiddle_factor_table_2_imag));
  assign _zz_8829 = ($signed(data_mid_63_real) + $signed(data_mid_63_imag));
  assign _zz_8830 = fixTo_570_dout;
  assign _zz_8831 = ($signed(_zz_478) + $signed(_zz_8832));
  assign _zz_8832 = ($signed(_zz_8833) * $signed(twiddle_factor_table_2_real));
  assign _zz_8833 = ($signed(data_mid_63_imag) - $signed(data_mid_63_real));
  assign _zz_8834 = fixTo_571_dout;
  assign _zz_8835 = _zz_8836[31 : 0];
  assign _zz_8836 = _zz_8837;
  assign _zz_8837 = ($signed(_zz_8838) >>> _zz_479);
  assign _zz_8838 = _zz_8839;
  assign _zz_8839 = ($signed(_zz_8841) - $signed(_zz_476));
  assign _zz_8840 = ({8'd0,data_mid_61_real} <<< 8);
  assign _zz_8841 = {{8{_zz_8840[23]}}, _zz_8840};
  assign _zz_8842 = fixTo_572_dout;
  assign _zz_8843 = _zz_8844[31 : 0];
  assign _zz_8844 = _zz_8845;
  assign _zz_8845 = ($signed(_zz_8846) >>> _zz_479);
  assign _zz_8846 = _zz_8847;
  assign _zz_8847 = ($signed(_zz_8849) - $signed(_zz_477));
  assign _zz_8848 = ({8'd0,data_mid_61_imag} <<< 8);
  assign _zz_8849 = {{8{_zz_8848[23]}}, _zz_8848};
  assign _zz_8850 = fixTo_573_dout;
  assign _zz_8851 = _zz_8852[31 : 0];
  assign _zz_8852 = _zz_8853;
  assign _zz_8853 = ($signed(_zz_8854) >>> _zz_480);
  assign _zz_8854 = _zz_8855;
  assign _zz_8855 = ($signed(_zz_8857) + $signed(_zz_476));
  assign _zz_8856 = ({8'd0,data_mid_61_real} <<< 8);
  assign _zz_8857 = {{8{_zz_8856[23]}}, _zz_8856};
  assign _zz_8858 = fixTo_574_dout;
  assign _zz_8859 = _zz_8860[31 : 0];
  assign _zz_8860 = _zz_8861;
  assign _zz_8861 = ($signed(_zz_8862) >>> _zz_480);
  assign _zz_8862 = _zz_8863;
  assign _zz_8863 = ($signed(_zz_8865) + $signed(_zz_477));
  assign _zz_8864 = ({8'd0,data_mid_61_imag} <<< 8);
  assign _zz_8865 = {{8{_zz_8864[23]}}, _zz_8864};
  assign _zz_8866 = fixTo_575_dout;
  assign _zz_8867 = ($signed(twiddle_factor_table_1_real) + $signed(twiddle_factor_table_1_imag));
  assign _zz_8868 = ($signed(_zz_483) - $signed(_zz_8869));
  assign _zz_8869 = ($signed(_zz_8870) * $signed(twiddle_factor_table_1_imag));
  assign _zz_8870 = ($signed(data_mid_66_real) + $signed(data_mid_66_imag));
  assign _zz_8871 = fixTo_576_dout;
  assign _zz_8872 = ($signed(_zz_483) + $signed(_zz_8873));
  assign _zz_8873 = ($signed(_zz_8874) * $signed(twiddle_factor_table_1_real));
  assign _zz_8874 = ($signed(data_mid_66_imag) - $signed(data_mid_66_real));
  assign _zz_8875 = fixTo_577_dout;
  assign _zz_8876 = _zz_8877[31 : 0];
  assign _zz_8877 = _zz_8878;
  assign _zz_8878 = ($signed(_zz_8879) >>> _zz_484);
  assign _zz_8879 = _zz_8880;
  assign _zz_8880 = ($signed(_zz_8882) - $signed(_zz_481));
  assign _zz_8881 = ({8'd0,data_mid_64_real} <<< 8);
  assign _zz_8882 = {{8{_zz_8881[23]}}, _zz_8881};
  assign _zz_8883 = fixTo_578_dout;
  assign _zz_8884 = _zz_8885[31 : 0];
  assign _zz_8885 = _zz_8886;
  assign _zz_8886 = ($signed(_zz_8887) >>> _zz_484);
  assign _zz_8887 = _zz_8888;
  assign _zz_8888 = ($signed(_zz_8890) - $signed(_zz_482));
  assign _zz_8889 = ({8'd0,data_mid_64_imag} <<< 8);
  assign _zz_8890 = {{8{_zz_8889[23]}}, _zz_8889};
  assign _zz_8891 = fixTo_579_dout;
  assign _zz_8892 = _zz_8893[31 : 0];
  assign _zz_8893 = _zz_8894;
  assign _zz_8894 = ($signed(_zz_8895) >>> _zz_485);
  assign _zz_8895 = _zz_8896;
  assign _zz_8896 = ($signed(_zz_8898) + $signed(_zz_481));
  assign _zz_8897 = ({8'd0,data_mid_64_real} <<< 8);
  assign _zz_8898 = {{8{_zz_8897[23]}}, _zz_8897};
  assign _zz_8899 = fixTo_580_dout;
  assign _zz_8900 = _zz_8901[31 : 0];
  assign _zz_8901 = _zz_8902;
  assign _zz_8902 = ($signed(_zz_8903) >>> _zz_485);
  assign _zz_8903 = _zz_8904;
  assign _zz_8904 = ($signed(_zz_8906) + $signed(_zz_482));
  assign _zz_8905 = ({8'd0,data_mid_64_imag} <<< 8);
  assign _zz_8906 = {{8{_zz_8905[23]}}, _zz_8905};
  assign _zz_8907 = fixTo_581_dout;
  assign _zz_8908 = ($signed(twiddle_factor_table_2_real) + $signed(twiddle_factor_table_2_imag));
  assign _zz_8909 = ($signed(_zz_488) - $signed(_zz_8910));
  assign _zz_8910 = ($signed(_zz_8911) * $signed(twiddle_factor_table_2_imag));
  assign _zz_8911 = ($signed(data_mid_67_real) + $signed(data_mid_67_imag));
  assign _zz_8912 = fixTo_582_dout;
  assign _zz_8913 = ($signed(_zz_488) + $signed(_zz_8914));
  assign _zz_8914 = ($signed(_zz_8915) * $signed(twiddle_factor_table_2_real));
  assign _zz_8915 = ($signed(data_mid_67_imag) - $signed(data_mid_67_real));
  assign _zz_8916 = fixTo_583_dout;
  assign _zz_8917 = _zz_8918[31 : 0];
  assign _zz_8918 = _zz_8919;
  assign _zz_8919 = ($signed(_zz_8920) >>> _zz_489);
  assign _zz_8920 = _zz_8921;
  assign _zz_8921 = ($signed(_zz_8923) - $signed(_zz_486));
  assign _zz_8922 = ({8'd0,data_mid_65_real} <<< 8);
  assign _zz_8923 = {{8{_zz_8922[23]}}, _zz_8922};
  assign _zz_8924 = fixTo_584_dout;
  assign _zz_8925 = _zz_8926[31 : 0];
  assign _zz_8926 = _zz_8927;
  assign _zz_8927 = ($signed(_zz_8928) >>> _zz_489);
  assign _zz_8928 = _zz_8929;
  assign _zz_8929 = ($signed(_zz_8931) - $signed(_zz_487));
  assign _zz_8930 = ({8'd0,data_mid_65_imag} <<< 8);
  assign _zz_8931 = {{8{_zz_8930[23]}}, _zz_8930};
  assign _zz_8932 = fixTo_585_dout;
  assign _zz_8933 = _zz_8934[31 : 0];
  assign _zz_8934 = _zz_8935;
  assign _zz_8935 = ($signed(_zz_8936) >>> _zz_490);
  assign _zz_8936 = _zz_8937;
  assign _zz_8937 = ($signed(_zz_8939) + $signed(_zz_486));
  assign _zz_8938 = ({8'd0,data_mid_65_real} <<< 8);
  assign _zz_8939 = {{8{_zz_8938[23]}}, _zz_8938};
  assign _zz_8940 = fixTo_586_dout;
  assign _zz_8941 = _zz_8942[31 : 0];
  assign _zz_8942 = _zz_8943;
  assign _zz_8943 = ($signed(_zz_8944) >>> _zz_490);
  assign _zz_8944 = _zz_8945;
  assign _zz_8945 = ($signed(_zz_8947) + $signed(_zz_487));
  assign _zz_8946 = ({8'd0,data_mid_65_imag} <<< 8);
  assign _zz_8947 = {{8{_zz_8946[23]}}, _zz_8946};
  assign _zz_8948 = fixTo_587_dout;
  assign _zz_8949 = ($signed(twiddle_factor_table_1_real) + $signed(twiddle_factor_table_1_imag));
  assign _zz_8950 = ($signed(_zz_493) - $signed(_zz_8951));
  assign _zz_8951 = ($signed(_zz_8952) * $signed(twiddle_factor_table_1_imag));
  assign _zz_8952 = ($signed(data_mid_70_real) + $signed(data_mid_70_imag));
  assign _zz_8953 = fixTo_588_dout;
  assign _zz_8954 = ($signed(_zz_493) + $signed(_zz_8955));
  assign _zz_8955 = ($signed(_zz_8956) * $signed(twiddle_factor_table_1_real));
  assign _zz_8956 = ($signed(data_mid_70_imag) - $signed(data_mid_70_real));
  assign _zz_8957 = fixTo_589_dout;
  assign _zz_8958 = _zz_8959[31 : 0];
  assign _zz_8959 = _zz_8960;
  assign _zz_8960 = ($signed(_zz_8961) >>> _zz_494);
  assign _zz_8961 = _zz_8962;
  assign _zz_8962 = ($signed(_zz_8964) - $signed(_zz_491));
  assign _zz_8963 = ({8'd0,data_mid_68_real} <<< 8);
  assign _zz_8964 = {{8{_zz_8963[23]}}, _zz_8963};
  assign _zz_8965 = fixTo_590_dout;
  assign _zz_8966 = _zz_8967[31 : 0];
  assign _zz_8967 = _zz_8968;
  assign _zz_8968 = ($signed(_zz_8969) >>> _zz_494);
  assign _zz_8969 = _zz_8970;
  assign _zz_8970 = ($signed(_zz_8972) - $signed(_zz_492));
  assign _zz_8971 = ({8'd0,data_mid_68_imag} <<< 8);
  assign _zz_8972 = {{8{_zz_8971[23]}}, _zz_8971};
  assign _zz_8973 = fixTo_591_dout;
  assign _zz_8974 = _zz_8975[31 : 0];
  assign _zz_8975 = _zz_8976;
  assign _zz_8976 = ($signed(_zz_8977) >>> _zz_495);
  assign _zz_8977 = _zz_8978;
  assign _zz_8978 = ($signed(_zz_8980) + $signed(_zz_491));
  assign _zz_8979 = ({8'd0,data_mid_68_real} <<< 8);
  assign _zz_8980 = {{8{_zz_8979[23]}}, _zz_8979};
  assign _zz_8981 = fixTo_592_dout;
  assign _zz_8982 = _zz_8983[31 : 0];
  assign _zz_8983 = _zz_8984;
  assign _zz_8984 = ($signed(_zz_8985) >>> _zz_495);
  assign _zz_8985 = _zz_8986;
  assign _zz_8986 = ($signed(_zz_8988) + $signed(_zz_492));
  assign _zz_8987 = ({8'd0,data_mid_68_imag} <<< 8);
  assign _zz_8988 = {{8{_zz_8987[23]}}, _zz_8987};
  assign _zz_8989 = fixTo_593_dout;
  assign _zz_8990 = ($signed(twiddle_factor_table_2_real) + $signed(twiddle_factor_table_2_imag));
  assign _zz_8991 = ($signed(_zz_498) - $signed(_zz_8992));
  assign _zz_8992 = ($signed(_zz_8993) * $signed(twiddle_factor_table_2_imag));
  assign _zz_8993 = ($signed(data_mid_71_real) + $signed(data_mid_71_imag));
  assign _zz_8994 = fixTo_594_dout;
  assign _zz_8995 = ($signed(_zz_498) + $signed(_zz_8996));
  assign _zz_8996 = ($signed(_zz_8997) * $signed(twiddle_factor_table_2_real));
  assign _zz_8997 = ($signed(data_mid_71_imag) - $signed(data_mid_71_real));
  assign _zz_8998 = fixTo_595_dout;
  assign _zz_8999 = _zz_9000[31 : 0];
  assign _zz_9000 = _zz_9001;
  assign _zz_9001 = ($signed(_zz_9002) >>> _zz_499);
  assign _zz_9002 = _zz_9003;
  assign _zz_9003 = ($signed(_zz_9005) - $signed(_zz_496));
  assign _zz_9004 = ({8'd0,data_mid_69_real} <<< 8);
  assign _zz_9005 = {{8{_zz_9004[23]}}, _zz_9004};
  assign _zz_9006 = fixTo_596_dout;
  assign _zz_9007 = _zz_9008[31 : 0];
  assign _zz_9008 = _zz_9009;
  assign _zz_9009 = ($signed(_zz_9010) >>> _zz_499);
  assign _zz_9010 = _zz_9011;
  assign _zz_9011 = ($signed(_zz_9013) - $signed(_zz_497));
  assign _zz_9012 = ({8'd0,data_mid_69_imag} <<< 8);
  assign _zz_9013 = {{8{_zz_9012[23]}}, _zz_9012};
  assign _zz_9014 = fixTo_597_dout;
  assign _zz_9015 = _zz_9016[31 : 0];
  assign _zz_9016 = _zz_9017;
  assign _zz_9017 = ($signed(_zz_9018) >>> _zz_500);
  assign _zz_9018 = _zz_9019;
  assign _zz_9019 = ($signed(_zz_9021) + $signed(_zz_496));
  assign _zz_9020 = ({8'd0,data_mid_69_real} <<< 8);
  assign _zz_9021 = {{8{_zz_9020[23]}}, _zz_9020};
  assign _zz_9022 = fixTo_598_dout;
  assign _zz_9023 = _zz_9024[31 : 0];
  assign _zz_9024 = _zz_9025;
  assign _zz_9025 = ($signed(_zz_9026) >>> _zz_500);
  assign _zz_9026 = _zz_9027;
  assign _zz_9027 = ($signed(_zz_9029) + $signed(_zz_497));
  assign _zz_9028 = ({8'd0,data_mid_69_imag} <<< 8);
  assign _zz_9029 = {{8{_zz_9028[23]}}, _zz_9028};
  assign _zz_9030 = fixTo_599_dout;
  assign _zz_9031 = ($signed(twiddle_factor_table_1_real) + $signed(twiddle_factor_table_1_imag));
  assign _zz_9032 = ($signed(_zz_503) - $signed(_zz_9033));
  assign _zz_9033 = ($signed(_zz_9034) * $signed(twiddle_factor_table_1_imag));
  assign _zz_9034 = ($signed(data_mid_74_real) + $signed(data_mid_74_imag));
  assign _zz_9035 = fixTo_600_dout;
  assign _zz_9036 = ($signed(_zz_503) + $signed(_zz_9037));
  assign _zz_9037 = ($signed(_zz_9038) * $signed(twiddle_factor_table_1_real));
  assign _zz_9038 = ($signed(data_mid_74_imag) - $signed(data_mid_74_real));
  assign _zz_9039 = fixTo_601_dout;
  assign _zz_9040 = _zz_9041[31 : 0];
  assign _zz_9041 = _zz_9042;
  assign _zz_9042 = ($signed(_zz_9043) >>> _zz_504);
  assign _zz_9043 = _zz_9044;
  assign _zz_9044 = ($signed(_zz_9046) - $signed(_zz_501));
  assign _zz_9045 = ({8'd0,data_mid_72_real} <<< 8);
  assign _zz_9046 = {{8{_zz_9045[23]}}, _zz_9045};
  assign _zz_9047 = fixTo_602_dout;
  assign _zz_9048 = _zz_9049[31 : 0];
  assign _zz_9049 = _zz_9050;
  assign _zz_9050 = ($signed(_zz_9051) >>> _zz_504);
  assign _zz_9051 = _zz_9052;
  assign _zz_9052 = ($signed(_zz_9054) - $signed(_zz_502));
  assign _zz_9053 = ({8'd0,data_mid_72_imag} <<< 8);
  assign _zz_9054 = {{8{_zz_9053[23]}}, _zz_9053};
  assign _zz_9055 = fixTo_603_dout;
  assign _zz_9056 = _zz_9057[31 : 0];
  assign _zz_9057 = _zz_9058;
  assign _zz_9058 = ($signed(_zz_9059) >>> _zz_505);
  assign _zz_9059 = _zz_9060;
  assign _zz_9060 = ($signed(_zz_9062) + $signed(_zz_501));
  assign _zz_9061 = ({8'd0,data_mid_72_real} <<< 8);
  assign _zz_9062 = {{8{_zz_9061[23]}}, _zz_9061};
  assign _zz_9063 = fixTo_604_dout;
  assign _zz_9064 = _zz_9065[31 : 0];
  assign _zz_9065 = _zz_9066;
  assign _zz_9066 = ($signed(_zz_9067) >>> _zz_505);
  assign _zz_9067 = _zz_9068;
  assign _zz_9068 = ($signed(_zz_9070) + $signed(_zz_502));
  assign _zz_9069 = ({8'd0,data_mid_72_imag} <<< 8);
  assign _zz_9070 = {{8{_zz_9069[23]}}, _zz_9069};
  assign _zz_9071 = fixTo_605_dout;
  assign _zz_9072 = ($signed(twiddle_factor_table_2_real) + $signed(twiddle_factor_table_2_imag));
  assign _zz_9073 = ($signed(_zz_508) - $signed(_zz_9074));
  assign _zz_9074 = ($signed(_zz_9075) * $signed(twiddle_factor_table_2_imag));
  assign _zz_9075 = ($signed(data_mid_75_real) + $signed(data_mid_75_imag));
  assign _zz_9076 = fixTo_606_dout;
  assign _zz_9077 = ($signed(_zz_508) + $signed(_zz_9078));
  assign _zz_9078 = ($signed(_zz_9079) * $signed(twiddle_factor_table_2_real));
  assign _zz_9079 = ($signed(data_mid_75_imag) - $signed(data_mid_75_real));
  assign _zz_9080 = fixTo_607_dout;
  assign _zz_9081 = _zz_9082[31 : 0];
  assign _zz_9082 = _zz_9083;
  assign _zz_9083 = ($signed(_zz_9084) >>> _zz_509);
  assign _zz_9084 = _zz_9085;
  assign _zz_9085 = ($signed(_zz_9087) - $signed(_zz_506));
  assign _zz_9086 = ({8'd0,data_mid_73_real} <<< 8);
  assign _zz_9087 = {{8{_zz_9086[23]}}, _zz_9086};
  assign _zz_9088 = fixTo_608_dout;
  assign _zz_9089 = _zz_9090[31 : 0];
  assign _zz_9090 = _zz_9091;
  assign _zz_9091 = ($signed(_zz_9092) >>> _zz_509);
  assign _zz_9092 = _zz_9093;
  assign _zz_9093 = ($signed(_zz_9095) - $signed(_zz_507));
  assign _zz_9094 = ({8'd0,data_mid_73_imag} <<< 8);
  assign _zz_9095 = {{8{_zz_9094[23]}}, _zz_9094};
  assign _zz_9096 = fixTo_609_dout;
  assign _zz_9097 = _zz_9098[31 : 0];
  assign _zz_9098 = _zz_9099;
  assign _zz_9099 = ($signed(_zz_9100) >>> _zz_510);
  assign _zz_9100 = _zz_9101;
  assign _zz_9101 = ($signed(_zz_9103) + $signed(_zz_506));
  assign _zz_9102 = ({8'd0,data_mid_73_real} <<< 8);
  assign _zz_9103 = {{8{_zz_9102[23]}}, _zz_9102};
  assign _zz_9104 = fixTo_610_dout;
  assign _zz_9105 = _zz_9106[31 : 0];
  assign _zz_9106 = _zz_9107;
  assign _zz_9107 = ($signed(_zz_9108) >>> _zz_510);
  assign _zz_9108 = _zz_9109;
  assign _zz_9109 = ($signed(_zz_9111) + $signed(_zz_507));
  assign _zz_9110 = ({8'd0,data_mid_73_imag} <<< 8);
  assign _zz_9111 = {{8{_zz_9110[23]}}, _zz_9110};
  assign _zz_9112 = fixTo_611_dout;
  assign _zz_9113 = ($signed(twiddle_factor_table_1_real) + $signed(twiddle_factor_table_1_imag));
  assign _zz_9114 = ($signed(_zz_513) - $signed(_zz_9115));
  assign _zz_9115 = ($signed(_zz_9116) * $signed(twiddle_factor_table_1_imag));
  assign _zz_9116 = ($signed(data_mid_78_real) + $signed(data_mid_78_imag));
  assign _zz_9117 = fixTo_612_dout;
  assign _zz_9118 = ($signed(_zz_513) + $signed(_zz_9119));
  assign _zz_9119 = ($signed(_zz_9120) * $signed(twiddle_factor_table_1_real));
  assign _zz_9120 = ($signed(data_mid_78_imag) - $signed(data_mid_78_real));
  assign _zz_9121 = fixTo_613_dout;
  assign _zz_9122 = _zz_9123[31 : 0];
  assign _zz_9123 = _zz_9124;
  assign _zz_9124 = ($signed(_zz_9125) >>> _zz_514);
  assign _zz_9125 = _zz_9126;
  assign _zz_9126 = ($signed(_zz_9128) - $signed(_zz_511));
  assign _zz_9127 = ({8'd0,data_mid_76_real} <<< 8);
  assign _zz_9128 = {{8{_zz_9127[23]}}, _zz_9127};
  assign _zz_9129 = fixTo_614_dout;
  assign _zz_9130 = _zz_9131[31 : 0];
  assign _zz_9131 = _zz_9132;
  assign _zz_9132 = ($signed(_zz_9133) >>> _zz_514);
  assign _zz_9133 = _zz_9134;
  assign _zz_9134 = ($signed(_zz_9136) - $signed(_zz_512));
  assign _zz_9135 = ({8'd0,data_mid_76_imag} <<< 8);
  assign _zz_9136 = {{8{_zz_9135[23]}}, _zz_9135};
  assign _zz_9137 = fixTo_615_dout;
  assign _zz_9138 = _zz_9139[31 : 0];
  assign _zz_9139 = _zz_9140;
  assign _zz_9140 = ($signed(_zz_9141) >>> _zz_515);
  assign _zz_9141 = _zz_9142;
  assign _zz_9142 = ($signed(_zz_9144) + $signed(_zz_511));
  assign _zz_9143 = ({8'd0,data_mid_76_real} <<< 8);
  assign _zz_9144 = {{8{_zz_9143[23]}}, _zz_9143};
  assign _zz_9145 = fixTo_616_dout;
  assign _zz_9146 = _zz_9147[31 : 0];
  assign _zz_9147 = _zz_9148;
  assign _zz_9148 = ($signed(_zz_9149) >>> _zz_515);
  assign _zz_9149 = _zz_9150;
  assign _zz_9150 = ($signed(_zz_9152) + $signed(_zz_512));
  assign _zz_9151 = ({8'd0,data_mid_76_imag} <<< 8);
  assign _zz_9152 = {{8{_zz_9151[23]}}, _zz_9151};
  assign _zz_9153 = fixTo_617_dout;
  assign _zz_9154 = ($signed(twiddle_factor_table_2_real) + $signed(twiddle_factor_table_2_imag));
  assign _zz_9155 = ($signed(_zz_518) - $signed(_zz_9156));
  assign _zz_9156 = ($signed(_zz_9157) * $signed(twiddle_factor_table_2_imag));
  assign _zz_9157 = ($signed(data_mid_79_real) + $signed(data_mid_79_imag));
  assign _zz_9158 = fixTo_618_dout;
  assign _zz_9159 = ($signed(_zz_518) + $signed(_zz_9160));
  assign _zz_9160 = ($signed(_zz_9161) * $signed(twiddle_factor_table_2_real));
  assign _zz_9161 = ($signed(data_mid_79_imag) - $signed(data_mid_79_real));
  assign _zz_9162 = fixTo_619_dout;
  assign _zz_9163 = _zz_9164[31 : 0];
  assign _zz_9164 = _zz_9165;
  assign _zz_9165 = ($signed(_zz_9166) >>> _zz_519);
  assign _zz_9166 = _zz_9167;
  assign _zz_9167 = ($signed(_zz_9169) - $signed(_zz_516));
  assign _zz_9168 = ({8'd0,data_mid_77_real} <<< 8);
  assign _zz_9169 = {{8{_zz_9168[23]}}, _zz_9168};
  assign _zz_9170 = fixTo_620_dout;
  assign _zz_9171 = _zz_9172[31 : 0];
  assign _zz_9172 = _zz_9173;
  assign _zz_9173 = ($signed(_zz_9174) >>> _zz_519);
  assign _zz_9174 = _zz_9175;
  assign _zz_9175 = ($signed(_zz_9177) - $signed(_zz_517));
  assign _zz_9176 = ({8'd0,data_mid_77_imag} <<< 8);
  assign _zz_9177 = {{8{_zz_9176[23]}}, _zz_9176};
  assign _zz_9178 = fixTo_621_dout;
  assign _zz_9179 = _zz_9180[31 : 0];
  assign _zz_9180 = _zz_9181;
  assign _zz_9181 = ($signed(_zz_9182) >>> _zz_520);
  assign _zz_9182 = _zz_9183;
  assign _zz_9183 = ($signed(_zz_9185) + $signed(_zz_516));
  assign _zz_9184 = ({8'd0,data_mid_77_real} <<< 8);
  assign _zz_9185 = {{8{_zz_9184[23]}}, _zz_9184};
  assign _zz_9186 = fixTo_622_dout;
  assign _zz_9187 = _zz_9188[31 : 0];
  assign _zz_9188 = _zz_9189;
  assign _zz_9189 = ($signed(_zz_9190) >>> _zz_520);
  assign _zz_9190 = _zz_9191;
  assign _zz_9191 = ($signed(_zz_9193) + $signed(_zz_517));
  assign _zz_9192 = ({8'd0,data_mid_77_imag} <<< 8);
  assign _zz_9193 = {{8{_zz_9192[23]}}, _zz_9192};
  assign _zz_9194 = fixTo_623_dout;
  assign _zz_9195 = ($signed(twiddle_factor_table_1_real) + $signed(twiddle_factor_table_1_imag));
  assign _zz_9196 = ($signed(_zz_523) - $signed(_zz_9197));
  assign _zz_9197 = ($signed(_zz_9198) * $signed(twiddle_factor_table_1_imag));
  assign _zz_9198 = ($signed(data_mid_82_real) + $signed(data_mid_82_imag));
  assign _zz_9199 = fixTo_624_dout;
  assign _zz_9200 = ($signed(_zz_523) + $signed(_zz_9201));
  assign _zz_9201 = ($signed(_zz_9202) * $signed(twiddle_factor_table_1_real));
  assign _zz_9202 = ($signed(data_mid_82_imag) - $signed(data_mid_82_real));
  assign _zz_9203 = fixTo_625_dout;
  assign _zz_9204 = _zz_9205[31 : 0];
  assign _zz_9205 = _zz_9206;
  assign _zz_9206 = ($signed(_zz_9207) >>> _zz_524);
  assign _zz_9207 = _zz_9208;
  assign _zz_9208 = ($signed(_zz_9210) - $signed(_zz_521));
  assign _zz_9209 = ({8'd0,data_mid_80_real} <<< 8);
  assign _zz_9210 = {{8{_zz_9209[23]}}, _zz_9209};
  assign _zz_9211 = fixTo_626_dout;
  assign _zz_9212 = _zz_9213[31 : 0];
  assign _zz_9213 = _zz_9214;
  assign _zz_9214 = ($signed(_zz_9215) >>> _zz_524);
  assign _zz_9215 = _zz_9216;
  assign _zz_9216 = ($signed(_zz_9218) - $signed(_zz_522));
  assign _zz_9217 = ({8'd0,data_mid_80_imag} <<< 8);
  assign _zz_9218 = {{8{_zz_9217[23]}}, _zz_9217};
  assign _zz_9219 = fixTo_627_dout;
  assign _zz_9220 = _zz_9221[31 : 0];
  assign _zz_9221 = _zz_9222;
  assign _zz_9222 = ($signed(_zz_9223) >>> _zz_525);
  assign _zz_9223 = _zz_9224;
  assign _zz_9224 = ($signed(_zz_9226) + $signed(_zz_521));
  assign _zz_9225 = ({8'd0,data_mid_80_real} <<< 8);
  assign _zz_9226 = {{8{_zz_9225[23]}}, _zz_9225};
  assign _zz_9227 = fixTo_628_dout;
  assign _zz_9228 = _zz_9229[31 : 0];
  assign _zz_9229 = _zz_9230;
  assign _zz_9230 = ($signed(_zz_9231) >>> _zz_525);
  assign _zz_9231 = _zz_9232;
  assign _zz_9232 = ($signed(_zz_9234) + $signed(_zz_522));
  assign _zz_9233 = ({8'd0,data_mid_80_imag} <<< 8);
  assign _zz_9234 = {{8{_zz_9233[23]}}, _zz_9233};
  assign _zz_9235 = fixTo_629_dout;
  assign _zz_9236 = ($signed(twiddle_factor_table_2_real) + $signed(twiddle_factor_table_2_imag));
  assign _zz_9237 = ($signed(_zz_528) - $signed(_zz_9238));
  assign _zz_9238 = ($signed(_zz_9239) * $signed(twiddle_factor_table_2_imag));
  assign _zz_9239 = ($signed(data_mid_83_real) + $signed(data_mid_83_imag));
  assign _zz_9240 = fixTo_630_dout;
  assign _zz_9241 = ($signed(_zz_528) + $signed(_zz_9242));
  assign _zz_9242 = ($signed(_zz_9243) * $signed(twiddle_factor_table_2_real));
  assign _zz_9243 = ($signed(data_mid_83_imag) - $signed(data_mid_83_real));
  assign _zz_9244 = fixTo_631_dout;
  assign _zz_9245 = _zz_9246[31 : 0];
  assign _zz_9246 = _zz_9247;
  assign _zz_9247 = ($signed(_zz_9248) >>> _zz_529);
  assign _zz_9248 = _zz_9249;
  assign _zz_9249 = ($signed(_zz_9251) - $signed(_zz_526));
  assign _zz_9250 = ({8'd0,data_mid_81_real} <<< 8);
  assign _zz_9251 = {{8{_zz_9250[23]}}, _zz_9250};
  assign _zz_9252 = fixTo_632_dout;
  assign _zz_9253 = _zz_9254[31 : 0];
  assign _zz_9254 = _zz_9255;
  assign _zz_9255 = ($signed(_zz_9256) >>> _zz_529);
  assign _zz_9256 = _zz_9257;
  assign _zz_9257 = ($signed(_zz_9259) - $signed(_zz_527));
  assign _zz_9258 = ({8'd0,data_mid_81_imag} <<< 8);
  assign _zz_9259 = {{8{_zz_9258[23]}}, _zz_9258};
  assign _zz_9260 = fixTo_633_dout;
  assign _zz_9261 = _zz_9262[31 : 0];
  assign _zz_9262 = _zz_9263;
  assign _zz_9263 = ($signed(_zz_9264) >>> _zz_530);
  assign _zz_9264 = _zz_9265;
  assign _zz_9265 = ($signed(_zz_9267) + $signed(_zz_526));
  assign _zz_9266 = ({8'd0,data_mid_81_real} <<< 8);
  assign _zz_9267 = {{8{_zz_9266[23]}}, _zz_9266};
  assign _zz_9268 = fixTo_634_dout;
  assign _zz_9269 = _zz_9270[31 : 0];
  assign _zz_9270 = _zz_9271;
  assign _zz_9271 = ($signed(_zz_9272) >>> _zz_530);
  assign _zz_9272 = _zz_9273;
  assign _zz_9273 = ($signed(_zz_9275) + $signed(_zz_527));
  assign _zz_9274 = ({8'd0,data_mid_81_imag} <<< 8);
  assign _zz_9275 = {{8{_zz_9274[23]}}, _zz_9274};
  assign _zz_9276 = fixTo_635_dout;
  assign _zz_9277 = ($signed(twiddle_factor_table_1_real) + $signed(twiddle_factor_table_1_imag));
  assign _zz_9278 = ($signed(_zz_533) - $signed(_zz_9279));
  assign _zz_9279 = ($signed(_zz_9280) * $signed(twiddle_factor_table_1_imag));
  assign _zz_9280 = ($signed(data_mid_86_real) + $signed(data_mid_86_imag));
  assign _zz_9281 = fixTo_636_dout;
  assign _zz_9282 = ($signed(_zz_533) + $signed(_zz_9283));
  assign _zz_9283 = ($signed(_zz_9284) * $signed(twiddle_factor_table_1_real));
  assign _zz_9284 = ($signed(data_mid_86_imag) - $signed(data_mid_86_real));
  assign _zz_9285 = fixTo_637_dout;
  assign _zz_9286 = _zz_9287[31 : 0];
  assign _zz_9287 = _zz_9288;
  assign _zz_9288 = ($signed(_zz_9289) >>> _zz_534);
  assign _zz_9289 = _zz_9290;
  assign _zz_9290 = ($signed(_zz_9292) - $signed(_zz_531));
  assign _zz_9291 = ({8'd0,data_mid_84_real} <<< 8);
  assign _zz_9292 = {{8{_zz_9291[23]}}, _zz_9291};
  assign _zz_9293 = fixTo_638_dout;
  assign _zz_9294 = _zz_9295[31 : 0];
  assign _zz_9295 = _zz_9296;
  assign _zz_9296 = ($signed(_zz_9297) >>> _zz_534);
  assign _zz_9297 = _zz_9298;
  assign _zz_9298 = ($signed(_zz_9300) - $signed(_zz_532));
  assign _zz_9299 = ({8'd0,data_mid_84_imag} <<< 8);
  assign _zz_9300 = {{8{_zz_9299[23]}}, _zz_9299};
  assign _zz_9301 = fixTo_639_dout;
  assign _zz_9302 = _zz_9303[31 : 0];
  assign _zz_9303 = _zz_9304;
  assign _zz_9304 = ($signed(_zz_9305) >>> _zz_535);
  assign _zz_9305 = _zz_9306;
  assign _zz_9306 = ($signed(_zz_9308) + $signed(_zz_531));
  assign _zz_9307 = ({8'd0,data_mid_84_real} <<< 8);
  assign _zz_9308 = {{8{_zz_9307[23]}}, _zz_9307};
  assign _zz_9309 = fixTo_640_dout;
  assign _zz_9310 = _zz_9311[31 : 0];
  assign _zz_9311 = _zz_9312;
  assign _zz_9312 = ($signed(_zz_9313) >>> _zz_535);
  assign _zz_9313 = _zz_9314;
  assign _zz_9314 = ($signed(_zz_9316) + $signed(_zz_532));
  assign _zz_9315 = ({8'd0,data_mid_84_imag} <<< 8);
  assign _zz_9316 = {{8{_zz_9315[23]}}, _zz_9315};
  assign _zz_9317 = fixTo_641_dout;
  assign _zz_9318 = ($signed(twiddle_factor_table_2_real) + $signed(twiddle_factor_table_2_imag));
  assign _zz_9319 = ($signed(_zz_538) - $signed(_zz_9320));
  assign _zz_9320 = ($signed(_zz_9321) * $signed(twiddle_factor_table_2_imag));
  assign _zz_9321 = ($signed(data_mid_87_real) + $signed(data_mid_87_imag));
  assign _zz_9322 = fixTo_642_dout;
  assign _zz_9323 = ($signed(_zz_538) + $signed(_zz_9324));
  assign _zz_9324 = ($signed(_zz_9325) * $signed(twiddle_factor_table_2_real));
  assign _zz_9325 = ($signed(data_mid_87_imag) - $signed(data_mid_87_real));
  assign _zz_9326 = fixTo_643_dout;
  assign _zz_9327 = _zz_9328[31 : 0];
  assign _zz_9328 = _zz_9329;
  assign _zz_9329 = ($signed(_zz_9330) >>> _zz_539);
  assign _zz_9330 = _zz_9331;
  assign _zz_9331 = ($signed(_zz_9333) - $signed(_zz_536));
  assign _zz_9332 = ({8'd0,data_mid_85_real} <<< 8);
  assign _zz_9333 = {{8{_zz_9332[23]}}, _zz_9332};
  assign _zz_9334 = fixTo_644_dout;
  assign _zz_9335 = _zz_9336[31 : 0];
  assign _zz_9336 = _zz_9337;
  assign _zz_9337 = ($signed(_zz_9338) >>> _zz_539);
  assign _zz_9338 = _zz_9339;
  assign _zz_9339 = ($signed(_zz_9341) - $signed(_zz_537));
  assign _zz_9340 = ({8'd0,data_mid_85_imag} <<< 8);
  assign _zz_9341 = {{8{_zz_9340[23]}}, _zz_9340};
  assign _zz_9342 = fixTo_645_dout;
  assign _zz_9343 = _zz_9344[31 : 0];
  assign _zz_9344 = _zz_9345;
  assign _zz_9345 = ($signed(_zz_9346) >>> _zz_540);
  assign _zz_9346 = _zz_9347;
  assign _zz_9347 = ($signed(_zz_9349) + $signed(_zz_536));
  assign _zz_9348 = ({8'd0,data_mid_85_real} <<< 8);
  assign _zz_9349 = {{8{_zz_9348[23]}}, _zz_9348};
  assign _zz_9350 = fixTo_646_dout;
  assign _zz_9351 = _zz_9352[31 : 0];
  assign _zz_9352 = _zz_9353;
  assign _zz_9353 = ($signed(_zz_9354) >>> _zz_540);
  assign _zz_9354 = _zz_9355;
  assign _zz_9355 = ($signed(_zz_9357) + $signed(_zz_537));
  assign _zz_9356 = ({8'd0,data_mid_85_imag} <<< 8);
  assign _zz_9357 = {{8{_zz_9356[23]}}, _zz_9356};
  assign _zz_9358 = fixTo_647_dout;
  assign _zz_9359 = ($signed(twiddle_factor_table_1_real) + $signed(twiddle_factor_table_1_imag));
  assign _zz_9360 = ($signed(_zz_543) - $signed(_zz_9361));
  assign _zz_9361 = ($signed(_zz_9362) * $signed(twiddle_factor_table_1_imag));
  assign _zz_9362 = ($signed(data_mid_90_real) + $signed(data_mid_90_imag));
  assign _zz_9363 = fixTo_648_dout;
  assign _zz_9364 = ($signed(_zz_543) + $signed(_zz_9365));
  assign _zz_9365 = ($signed(_zz_9366) * $signed(twiddle_factor_table_1_real));
  assign _zz_9366 = ($signed(data_mid_90_imag) - $signed(data_mid_90_real));
  assign _zz_9367 = fixTo_649_dout;
  assign _zz_9368 = _zz_9369[31 : 0];
  assign _zz_9369 = _zz_9370;
  assign _zz_9370 = ($signed(_zz_9371) >>> _zz_544);
  assign _zz_9371 = _zz_9372;
  assign _zz_9372 = ($signed(_zz_9374) - $signed(_zz_541));
  assign _zz_9373 = ({8'd0,data_mid_88_real} <<< 8);
  assign _zz_9374 = {{8{_zz_9373[23]}}, _zz_9373};
  assign _zz_9375 = fixTo_650_dout;
  assign _zz_9376 = _zz_9377[31 : 0];
  assign _zz_9377 = _zz_9378;
  assign _zz_9378 = ($signed(_zz_9379) >>> _zz_544);
  assign _zz_9379 = _zz_9380;
  assign _zz_9380 = ($signed(_zz_9382) - $signed(_zz_542));
  assign _zz_9381 = ({8'd0,data_mid_88_imag} <<< 8);
  assign _zz_9382 = {{8{_zz_9381[23]}}, _zz_9381};
  assign _zz_9383 = fixTo_651_dout;
  assign _zz_9384 = _zz_9385[31 : 0];
  assign _zz_9385 = _zz_9386;
  assign _zz_9386 = ($signed(_zz_9387) >>> _zz_545);
  assign _zz_9387 = _zz_9388;
  assign _zz_9388 = ($signed(_zz_9390) + $signed(_zz_541));
  assign _zz_9389 = ({8'd0,data_mid_88_real} <<< 8);
  assign _zz_9390 = {{8{_zz_9389[23]}}, _zz_9389};
  assign _zz_9391 = fixTo_652_dout;
  assign _zz_9392 = _zz_9393[31 : 0];
  assign _zz_9393 = _zz_9394;
  assign _zz_9394 = ($signed(_zz_9395) >>> _zz_545);
  assign _zz_9395 = _zz_9396;
  assign _zz_9396 = ($signed(_zz_9398) + $signed(_zz_542));
  assign _zz_9397 = ({8'd0,data_mid_88_imag} <<< 8);
  assign _zz_9398 = {{8{_zz_9397[23]}}, _zz_9397};
  assign _zz_9399 = fixTo_653_dout;
  assign _zz_9400 = ($signed(twiddle_factor_table_2_real) + $signed(twiddle_factor_table_2_imag));
  assign _zz_9401 = ($signed(_zz_548) - $signed(_zz_9402));
  assign _zz_9402 = ($signed(_zz_9403) * $signed(twiddle_factor_table_2_imag));
  assign _zz_9403 = ($signed(data_mid_91_real) + $signed(data_mid_91_imag));
  assign _zz_9404 = fixTo_654_dout;
  assign _zz_9405 = ($signed(_zz_548) + $signed(_zz_9406));
  assign _zz_9406 = ($signed(_zz_9407) * $signed(twiddle_factor_table_2_real));
  assign _zz_9407 = ($signed(data_mid_91_imag) - $signed(data_mid_91_real));
  assign _zz_9408 = fixTo_655_dout;
  assign _zz_9409 = _zz_9410[31 : 0];
  assign _zz_9410 = _zz_9411;
  assign _zz_9411 = ($signed(_zz_9412) >>> _zz_549);
  assign _zz_9412 = _zz_9413;
  assign _zz_9413 = ($signed(_zz_9415) - $signed(_zz_546));
  assign _zz_9414 = ({8'd0,data_mid_89_real} <<< 8);
  assign _zz_9415 = {{8{_zz_9414[23]}}, _zz_9414};
  assign _zz_9416 = fixTo_656_dout;
  assign _zz_9417 = _zz_9418[31 : 0];
  assign _zz_9418 = _zz_9419;
  assign _zz_9419 = ($signed(_zz_9420) >>> _zz_549);
  assign _zz_9420 = _zz_9421;
  assign _zz_9421 = ($signed(_zz_9423) - $signed(_zz_547));
  assign _zz_9422 = ({8'd0,data_mid_89_imag} <<< 8);
  assign _zz_9423 = {{8{_zz_9422[23]}}, _zz_9422};
  assign _zz_9424 = fixTo_657_dout;
  assign _zz_9425 = _zz_9426[31 : 0];
  assign _zz_9426 = _zz_9427;
  assign _zz_9427 = ($signed(_zz_9428) >>> _zz_550);
  assign _zz_9428 = _zz_9429;
  assign _zz_9429 = ($signed(_zz_9431) + $signed(_zz_546));
  assign _zz_9430 = ({8'd0,data_mid_89_real} <<< 8);
  assign _zz_9431 = {{8{_zz_9430[23]}}, _zz_9430};
  assign _zz_9432 = fixTo_658_dout;
  assign _zz_9433 = _zz_9434[31 : 0];
  assign _zz_9434 = _zz_9435;
  assign _zz_9435 = ($signed(_zz_9436) >>> _zz_550);
  assign _zz_9436 = _zz_9437;
  assign _zz_9437 = ($signed(_zz_9439) + $signed(_zz_547));
  assign _zz_9438 = ({8'd0,data_mid_89_imag} <<< 8);
  assign _zz_9439 = {{8{_zz_9438[23]}}, _zz_9438};
  assign _zz_9440 = fixTo_659_dout;
  assign _zz_9441 = ($signed(twiddle_factor_table_1_real) + $signed(twiddle_factor_table_1_imag));
  assign _zz_9442 = ($signed(_zz_553) - $signed(_zz_9443));
  assign _zz_9443 = ($signed(_zz_9444) * $signed(twiddle_factor_table_1_imag));
  assign _zz_9444 = ($signed(data_mid_94_real) + $signed(data_mid_94_imag));
  assign _zz_9445 = fixTo_660_dout;
  assign _zz_9446 = ($signed(_zz_553) + $signed(_zz_9447));
  assign _zz_9447 = ($signed(_zz_9448) * $signed(twiddle_factor_table_1_real));
  assign _zz_9448 = ($signed(data_mid_94_imag) - $signed(data_mid_94_real));
  assign _zz_9449 = fixTo_661_dout;
  assign _zz_9450 = _zz_9451[31 : 0];
  assign _zz_9451 = _zz_9452;
  assign _zz_9452 = ($signed(_zz_9453) >>> _zz_554);
  assign _zz_9453 = _zz_9454;
  assign _zz_9454 = ($signed(_zz_9456) - $signed(_zz_551));
  assign _zz_9455 = ({8'd0,data_mid_92_real} <<< 8);
  assign _zz_9456 = {{8{_zz_9455[23]}}, _zz_9455};
  assign _zz_9457 = fixTo_662_dout;
  assign _zz_9458 = _zz_9459[31 : 0];
  assign _zz_9459 = _zz_9460;
  assign _zz_9460 = ($signed(_zz_9461) >>> _zz_554);
  assign _zz_9461 = _zz_9462;
  assign _zz_9462 = ($signed(_zz_9464) - $signed(_zz_552));
  assign _zz_9463 = ({8'd0,data_mid_92_imag} <<< 8);
  assign _zz_9464 = {{8{_zz_9463[23]}}, _zz_9463};
  assign _zz_9465 = fixTo_663_dout;
  assign _zz_9466 = _zz_9467[31 : 0];
  assign _zz_9467 = _zz_9468;
  assign _zz_9468 = ($signed(_zz_9469) >>> _zz_555);
  assign _zz_9469 = _zz_9470;
  assign _zz_9470 = ($signed(_zz_9472) + $signed(_zz_551));
  assign _zz_9471 = ({8'd0,data_mid_92_real} <<< 8);
  assign _zz_9472 = {{8{_zz_9471[23]}}, _zz_9471};
  assign _zz_9473 = fixTo_664_dout;
  assign _zz_9474 = _zz_9475[31 : 0];
  assign _zz_9475 = _zz_9476;
  assign _zz_9476 = ($signed(_zz_9477) >>> _zz_555);
  assign _zz_9477 = _zz_9478;
  assign _zz_9478 = ($signed(_zz_9480) + $signed(_zz_552));
  assign _zz_9479 = ({8'd0,data_mid_92_imag} <<< 8);
  assign _zz_9480 = {{8{_zz_9479[23]}}, _zz_9479};
  assign _zz_9481 = fixTo_665_dout;
  assign _zz_9482 = ($signed(twiddle_factor_table_2_real) + $signed(twiddle_factor_table_2_imag));
  assign _zz_9483 = ($signed(_zz_558) - $signed(_zz_9484));
  assign _zz_9484 = ($signed(_zz_9485) * $signed(twiddle_factor_table_2_imag));
  assign _zz_9485 = ($signed(data_mid_95_real) + $signed(data_mid_95_imag));
  assign _zz_9486 = fixTo_666_dout;
  assign _zz_9487 = ($signed(_zz_558) + $signed(_zz_9488));
  assign _zz_9488 = ($signed(_zz_9489) * $signed(twiddle_factor_table_2_real));
  assign _zz_9489 = ($signed(data_mid_95_imag) - $signed(data_mid_95_real));
  assign _zz_9490 = fixTo_667_dout;
  assign _zz_9491 = _zz_9492[31 : 0];
  assign _zz_9492 = _zz_9493;
  assign _zz_9493 = ($signed(_zz_9494) >>> _zz_559);
  assign _zz_9494 = _zz_9495;
  assign _zz_9495 = ($signed(_zz_9497) - $signed(_zz_556));
  assign _zz_9496 = ({8'd0,data_mid_93_real} <<< 8);
  assign _zz_9497 = {{8{_zz_9496[23]}}, _zz_9496};
  assign _zz_9498 = fixTo_668_dout;
  assign _zz_9499 = _zz_9500[31 : 0];
  assign _zz_9500 = _zz_9501;
  assign _zz_9501 = ($signed(_zz_9502) >>> _zz_559);
  assign _zz_9502 = _zz_9503;
  assign _zz_9503 = ($signed(_zz_9505) - $signed(_zz_557));
  assign _zz_9504 = ({8'd0,data_mid_93_imag} <<< 8);
  assign _zz_9505 = {{8{_zz_9504[23]}}, _zz_9504};
  assign _zz_9506 = fixTo_669_dout;
  assign _zz_9507 = _zz_9508[31 : 0];
  assign _zz_9508 = _zz_9509;
  assign _zz_9509 = ($signed(_zz_9510) >>> _zz_560);
  assign _zz_9510 = _zz_9511;
  assign _zz_9511 = ($signed(_zz_9513) + $signed(_zz_556));
  assign _zz_9512 = ({8'd0,data_mid_93_real} <<< 8);
  assign _zz_9513 = {{8{_zz_9512[23]}}, _zz_9512};
  assign _zz_9514 = fixTo_670_dout;
  assign _zz_9515 = _zz_9516[31 : 0];
  assign _zz_9516 = _zz_9517;
  assign _zz_9517 = ($signed(_zz_9518) >>> _zz_560);
  assign _zz_9518 = _zz_9519;
  assign _zz_9519 = ($signed(_zz_9521) + $signed(_zz_557));
  assign _zz_9520 = ({8'd0,data_mid_93_imag} <<< 8);
  assign _zz_9521 = {{8{_zz_9520[23]}}, _zz_9520};
  assign _zz_9522 = fixTo_671_dout;
  assign _zz_9523 = ($signed(twiddle_factor_table_1_real) + $signed(twiddle_factor_table_1_imag));
  assign _zz_9524 = ($signed(_zz_563) - $signed(_zz_9525));
  assign _zz_9525 = ($signed(_zz_9526) * $signed(twiddle_factor_table_1_imag));
  assign _zz_9526 = ($signed(data_mid_98_real) + $signed(data_mid_98_imag));
  assign _zz_9527 = fixTo_672_dout;
  assign _zz_9528 = ($signed(_zz_563) + $signed(_zz_9529));
  assign _zz_9529 = ($signed(_zz_9530) * $signed(twiddle_factor_table_1_real));
  assign _zz_9530 = ($signed(data_mid_98_imag) - $signed(data_mid_98_real));
  assign _zz_9531 = fixTo_673_dout;
  assign _zz_9532 = _zz_9533[31 : 0];
  assign _zz_9533 = _zz_9534;
  assign _zz_9534 = ($signed(_zz_9535) >>> _zz_564);
  assign _zz_9535 = _zz_9536;
  assign _zz_9536 = ($signed(_zz_9538) - $signed(_zz_561));
  assign _zz_9537 = ({8'd0,data_mid_96_real} <<< 8);
  assign _zz_9538 = {{8{_zz_9537[23]}}, _zz_9537};
  assign _zz_9539 = fixTo_674_dout;
  assign _zz_9540 = _zz_9541[31 : 0];
  assign _zz_9541 = _zz_9542;
  assign _zz_9542 = ($signed(_zz_9543) >>> _zz_564);
  assign _zz_9543 = _zz_9544;
  assign _zz_9544 = ($signed(_zz_9546) - $signed(_zz_562));
  assign _zz_9545 = ({8'd0,data_mid_96_imag} <<< 8);
  assign _zz_9546 = {{8{_zz_9545[23]}}, _zz_9545};
  assign _zz_9547 = fixTo_675_dout;
  assign _zz_9548 = _zz_9549[31 : 0];
  assign _zz_9549 = _zz_9550;
  assign _zz_9550 = ($signed(_zz_9551) >>> _zz_565);
  assign _zz_9551 = _zz_9552;
  assign _zz_9552 = ($signed(_zz_9554) + $signed(_zz_561));
  assign _zz_9553 = ({8'd0,data_mid_96_real} <<< 8);
  assign _zz_9554 = {{8{_zz_9553[23]}}, _zz_9553};
  assign _zz_9555 = fixTo_676_dout;
  assign _zz_9556 = _zz_9557[31 : 0];
  assign _zz_9557 = _zz_9558;
  assign _zz_9558 = ($signed(_zz_9559) >>> _zz_565);
  assign _zz_9559 = _zz_9560;
  assign _zz_9560 = ($signed(_zz_9562) + $signed(_zz_562));
  assign _zz_9561 = ({8'd0,data_mid_96_imag} <<< 8);
  assign _zz_9562 = {{8{_zz_9561[23]}}, _zz_9561};
  assign _zz_9563 = fixTo_677_dout;
  assign _zz_9564 = ($signed(twiddle_factor_table_2_real) + $signed(twiddle_factor_table_2_imag));
  assign _zz_9565 = ($signed(_zz_568) - $signed(_zz_9566));
  assign _zz_9566 = ($signed(_zz_9567) * $signed(twiddle_factor_table_2_imag));
  assign _zz_9567 = ($signed(data_mid_99_real) + $signed(data_mid_99_imag));
  assign _zz_9568 = fixTo_678_dout;
  assign _zz_9569 = ($signed(_zz_568) + $signed(_zz_9570));
  assign _zz_9570 = ($signed(_zz_9571) * $signed(twiddle_factor_table_2_real));
  assign _zz_9571 = ($signed(data_mid_99_imag) - $signed(data_mid_99_real));
  assign _zz_9572 = fixTo_679_dout;
  assign _zz_9573 = _zz_9574[31 : 0];
  assign _zz_9574 = _zz_9575;
  assign _zz_9575 = ($signed(_zz_9576) >>> _zz_569);
  assign _zz_9576 = _zz_9577;
  assign _zz_9577 = ($signed(_zz_9579) - $signed(_zz_566));
  assign _zz_9578 = ({8'd0,data_mid_97_real} <<< 8);
  assign _zz_9579 = {{8{_zz_9578[23]}}, _zz_9578};
  assign _zz_9580 = fixTo_680_dout;
  assign _zz_9581 = _zz_9582[31 : 0];
  assign _zz_9582 = _zz_9583;
  assign _zz_9583 = ($signed(_zz_9584) >>> _zz_569);
  assign _zz_9584 = _zz_9585;
  assign _zz_9585 = ($signed(_zz_9587) - $signed(_zz_567));
  assign _zz_9586 = ({8'd0,data_mid_97_imag} <<< 8);
  assign _zz_9587 = {{8{_zz_9586[23]}}, _zz_9586};
  assign _zz_9588 = fixTo_681_dout;
  assign _zz_9589 = _zz_9590[31 : 0];
  assign _zz_9590 = _zz_9591;
  assign _zz_9591 = ($signed(_zz_9592) >>> _zz_570);
  assign _zz_9592 = _zz_9593;
  assign _zz_9593 = ($signed(_zz_9595) + $signed(_zz_566));
  assign _zz_9594 = ({8'd0,data_mid_97_real} <<< 8);
  assign _zz_9595 = {{8{_zz_9594[23]}}, _zz_9594};
  assign _zz_9596 = fixTo_682_dout;
  assign _zz_9597 = _zz_9598[31 : 0];
  assign _zz_9598 = _zz_9599;
  assign _zz_9599 = ($signed(_zz_9600) >>> _zz_570);
  assign _zz_9600 = _zz_9601;
  assign _zz_9601 = ($signed(_zz_9603) + $signed(_zz_567));
  assign _zz_9602 = ({8'd0,data_mid_97_imag} <<< 8);
  assign _zz_9603 = {{8{_zz_9602[23]}}, _zz_9602};
  assign _zz_9604 = fixTo_683_dout;
  assign _zz_9605 = ($signed(twiddle_factor_table_1_real) + $signed(twiddle_factor_table_1_imag));
  assign _zz_9606 = ($signed(_zz_573) - $signed(_zz_9607));
  assign _zz_9607 = ($signed(_zz_9608) * $signed(twiddle_factor_table_1_imag));
  assign _zz_9608 = ($signed(data_mid_102_real) + $signed(data_mid_102_imag));
  assign _zz_9609 = fixTo_684_dout;
  assign _zz_9610 = ($signed(_zz_573) + $signed(_zz_9611));
  assign _zz_9611 = ($signed(_zz_9612) * $signed(twiddle_factor_table_1_real));
  assign _zz_9612 = ($signed(data_mid_102_imag) - $signed(data_mid_102_real));
  assign _zz_9613 = fixTo_685_dout;
  assign _zz_9614 = _zz_9615[31 : 0];
  assign _zz_9615 = _zz_9616;
  assign _zz_9616 = ($signed(_zz_9617) >>> _zz_574);
  assign _zz_9617 = _zz_9618;
  assign _zz_9618 = ($signed(_zz_9620) - $signed(_zz_571));
  assign _zz_9619 = ({8'd0,data_mid_100_real} <<< 8);
  assign _zz_9620 = {{8{_zz_9619[23]}}, _zz_9619};
  assign _zz_9621 = fixTo_686_dout;
  assign _zz_9622 = _zz_9623[31 : 0];
  assign _zz_9623 = _zz_9624;
  assign _zz_9624 = ($signed(_zz_9625) >>> _zz_574);
  assign _zz_9625 = _zz_9626;
  assign _zz_9626 = ($signed(_zz_9628) - $signed(_zz_572));
  assign _zz_9627 = ({8'd0,data_mid_100_imag} <<< 8);
  assign _zz_9628 = {{8{_zz_9627[23]}}, _zz_9627};
  assign _zz_9629 = fixTo_687_dout;
  assign _zz_9630 = _zz_9631[31 : 0];
  assign _zz_9631 = _zz_9632;
  assign _zz_9632 = ($signed(_zz_9633) >>> _zz_575);
  assign _zz_9633 = _zz_9634;
  assign _zz_9634 = ($signed(_zz_9636) + $signed(_zz_571));
  assign _zz_9635 = ({8'd0,data_mid_100_real} <<< 8);
  assign _zz_9636 = {{8{_zz_9635[23]}}, _zz_9635};
  assign _zz_9637 = fixTo_688_dout;
  assign _zz_9638 = _zz_9639[31 : 0];
  assign _zz_9639 = _zz_9640;
  assign _zz_9640 = ($signed(_zz_9641) >>> _zz_575);
  assign _zz_9641 = _zz_9642;
  assign _zz_9642 = ($signed(_zz_9644) + $signed(_zz_572));
  assign _zz_9643 = ({8'd0,data_mid_100_imag} <<< 8);
  assign _zz_9644 = {{8{_zz_9643[23]}}, _zz_9643};
  assign _zz_9645 = fixTo_689_dout;
  assign _zz_9646 = ($signed(twiddle_factor_table_2_real) + $signed(twiddle_factor_table_2_imag));
  assign _zz_9647 = ($signed(_zz_578) - $signed(_zz_9648));
  assign _zz_9648 = ($signed(_zz_9649) * $signed(twiddle_factor_table_2_imag));
  assign _zz_9649 = ($signed(data_mid_103_real) + $signed(data_mid_103_imag));
  assign _zz_9650 = fixTo_690_dout;
  assign _zz_9651 = ($signed(_zz_578) + $signed(_zz_9652));
  assign _zz_9652 = ($signed(_zz_9653) * $signed(twiddle_factor_table_2_real));
  assign _zz_9653 = ($signed(data_mid_103_imag) - $signed(data_mid_103_real));
  assign _zz_9654 = fixTo_691_dout;
  assign _zz_9655 = _zz_9656[31 : 0];
  assign _zz_9656 = _zz_9657;
  assign _zz_9657 = ($signed(_zz_9658) >>> _zz_579);
  assign _zz_9658 = _zz_9659;
  assign _zz_9659 = ($signed(_zz_9661) - $signed(_zz_576));
  assign _zz_9660 = ({8'd0,data_mid_101_real} <<< 8);
  assign _zz_9661 = {{8{_zz_9660[23]}}, _zz_9660};
  assign _zz_9662 = fixTo_692_dout;
  assign _zz_9663 = _zz_9664[31 : 0];
  assign _zz_9664 = _zz_9665;
  assign _zz_9665 = ($signed(_zz_9666) >>> _zz_579);
  assign _zz_9666 = _zz_9667;
  assign _zz_9667 = ($signed(_zz_9669) - $signed(_zz_577));
  assign _zz_9668 = ({8'd0,data_mid_101_imag} <<< 8);
  assign _zz_9669 = {{8{_zz_9668[23]}}, _zz_9668};
  assign _zz_9670 = fixTo_693_dout;
  assign _zz_9671 = _zz_9672[31 : 0];
  assign _zz_9672 = _zz_9673;
  assign _zz_9673 = ($signed(_zz_9674) >>> _zz_580);
  assign _zz_9674 = _zz_9675;
  assign _zz_9675 = ($signed(_zz_9677) + $signed(_zz_576));
  assign _zz_9676 = ({8'd0,data_mid_101_real} <<< 8);
  assign _zz_9677 = {{8{_zz_9676[23]}}, _zz_9676};
  assign _zz_9678 = fixTo_694_dout;
  assign _zz_9679 = _zz_9680[31 : 0];
  assign _zz_9680 = _zz_9681;
  assign _zz_9681 = ($signed(_zz_9682) >>> _zz_580);
  assign _zz_9682 = _zz_9683;
  assign _zz_9683 = ($signed(_zz_9685) + $signed(_zz_577));
  assign _zz_9684 = ({8'd0,data_mid_101_imag} <<< 8);
  assign _zz_9685 = {{8{_zz_9684[23]}}, _zz_9684};
  assign _zz_9686 = fixTo_695_dout;
  assign _zz_9687 = ($signed(twiddle_factor_table_1_real) + $signed(twiddle_factor_table_1_imag));
  assign _zz_9688 = ($signed(_zz_583) - $signed(_zz_9689));
  assign _zz_9689 = ($signed(_zz_9690) * $signed(twiddle_factor_table_1_imag));
  assign _zz_9690 = ($signed(data_mid_106_real) + $signed(data_mid_106_imag));
  assign _zz_9691 = fixTo_696_dout;
  assign _zz_9692 = ($signed(_zz_583) + $signed(_zz_9693));
  assign _zz_9693 = ($signed(_zz_9694) * $signed(twiddle_factor_table_1_real));
  assign _zz_9694 = ($signed(data_mid_106_imag) - $signed(data_mid_106_real));
  assign _zz_9695 = fixTo_697_dout;
  assign _zz_9696 = _zz_9697[31 : 0];
  assign _zz_9697 = _zz_9698;
  assign _zz_9698 = ($signed(_zz_9699) >>> _zz_584);
  assign _zz_9699 = _zz_9700;
  assign _zz_9700 = ($signed(_zz_9702) - $signed(_zz_581));
  assign _zz_9701 = ({8'd0,data_mid_104_real} <<< 8);
  assign _zz_9702 = {{8{_zz_9701[23]}}, _zz_9701};
  assign _zz_9703 = fixTo_698_dout;
  assign _zz_9704 = _zz_9705[31 : 0];
  assign _zz_9705 = _zz_9706;
  assign _zz_9706 = ($signed(_zz_9707) >>> _zz_584);
  assign _zz_9707 = _zz_9708;
  assign _zz_9708 = ($signed(_zz_9710) - $signed(_zz_582));
  assign _zz_9709 = ({8'd0,data_mid_104_imag} <<< 8);
  assign _zz_9710 = {{8{_zz_9709[23]}}, _zz_9709};
  assign _zz_9711 = fixTo_699_dout;
  assign _zz_9712 = _zz_9713[31 : 0];
  assign _zz_9713 = _zz_9714;
  assign _zz_9714 = ($signed(_zz_9715) >>> _zz_585);
  assign _zz_9715 = _zz_9716;
  assign _zz_9716 = ($signed(_zz_9718) + $signed(_zz_581));
  assign _zz_9717 = ({8'd0,data_mid_104_real} <<< 8);
  assign _zz_9718 = {{8{_zz_9717[23]}}, _zz_9717};
  assign _zz_9719 = fixTo_700_dout;
  assign _zz_9720 = _zz_9721[31 : 0];
  assign _zz_9721 = _zz_9722;
  assign _zz_9722 = ($signed(_zz_9723) >>> _zz_585);
  assign _zz_9723 = _zz_9724;
  assign _zz_9724 = ($signed(_zz_9726) + $signed(_zz_582));
  assign _zz_9725 = ({8'd0,data_mid_104_imag} <<< 8);
  assign _zz_9726 = {{8{_zz_9725[23]}}, _zz_9725};
  assign _zz_9727 = fixTo_701_dout;
  assign _zz_9728 = ($signed(twiddle_factor_table_2_real) + $signed(twiddle_factor_table_2_imag));
  assign _zz_9729 = ($signed(_zz_588) - $signed(_zz_9730));
  assign _zz_9730 = ($signed(_zz_9731) * $signed(twiddle_factor_table_2_imag));
  assign _zz_9731 = ($signed(data_mid_107_real) + $signed(data_mid_107_imag));
  assign _zz_9732 = fixTo_702_dout;
  assign _zz_9733 = ($signed(_zz_588) + $signed(_zz_9734));
  assign _zz_9734 = ($signed(_zz_9735) * $signed(twiddle_factor_table_2_real));
  assign _zz_9735 = ($signed(data_mid_107_imag) - $signed(data_mid_107_real));
  assign _zz_9736 = fixTo_703_dout;
  assign _zz_9737 = _zz_9738[31 : 0];
  assign _zz_9738 = _zz_9739;
  assign _zz_9739 = ($signed(_zz_9740) >>> _zz_589);
  assign _zz_9740 = _zz_9741;
  assign _zz_9741 = ($signed(_zz_9743) - $signed(_zz_586));
  assign _zz_9742 = ({8'd0,data_mid_105_real} <<< 8);
  assign _zz_9743 = {{8{_zz_9742[23]}}, _zz_9742};
  assign _zz_9744 = fixTo_704_dout;
  assign _zz_9745 = _zz_9746[31 : 0];
  assign _zz_9746 = _zz_9747;
  assign _zz_9747 = ($signed(_zz_9748) >>> _zz_589);
  assign _zz_9748 = _zz_9749;
  assign _zz_9749 = ($signed(_zz_9751) - $signed(_zz_587));
  assign _zz_9750 = ({8'd0,data_mid_105_imag} <<< 8);
  assign _zz_9751 = {{8{_zz_9750[23]}}, _zz_9750};
  assign _zz_9752 = fixTo_705_dout;
  assign _zz_9753 = _zz_9754[31 : 0];
  assign _zz_9754 = _zz_9755;
  assign _zz_9755 = ($signed(_zz_9756) >>> _zz_590);
  assign _zz_9756 = _zz_9757;
  assign _zz_9757 = ($signed(_zz_9759) + $signed(_zz_586));
  assign _zz_9758 = ({8'd0,data_mid_105_real} <<< 8);
  assign _zz_9759 = {{8{_zz_9758[23]}}, _zz_9758};
  assign _zz_9760 = fixTo_706_dout;
  assign _zz_9761 = _zz_9762[31 : 0];
  assign _zz_9762 = _zz_9763;
  assign _zz_9763 = ($signed(_zz_9764) >>> _zz_590);
  assign _zz_9764 = _zz_9765;
  assign _zz_9765 = ($signed(_zz_9767) + $signed(_zz_587));
  assign _zz_9766 = ({8'd0,data_mid_105_imag} <<< 8);
  assign _zz_9767 = {{8{_zz_9766[23]}}, _zz_9766};
  assign _zz_9768 = fixTo_707_dout;
  assign _zz_9769 = ($signed(twiddle_factor_table_1_real) + $signed(twiddle_factor_table_1_imag));
  assign _zz_9770 = ($signed(_zz_593) - $signed(_zz_9771));
  assign _zz_9771 = ($signed(_zz_9772) * $signed(twiddle_factor_table_1_imag));
  assign _zz_9772 = ($signed(data_mid_110_real) + $signed(data_mid_110_imag));
  assign _zz_9773 = fixTo_708_dout;
  assign _zz_9774 = ($signed(_zz_593) + $signed(_zz_9775));
  assign _zz_9775 = ($signed(_zz_9776) * $signed(twiddle_factor_table_1_real));
  assign _zz_9776 = ($signed(data_mid_110_imag) - $signed(data_mid_110_real));
  assign _zz_9777 = fixTo_709_dout;
  assign _zz_9778 = _zz_9779[31 : 0];
  assign _zz_9779 = _zz_9780;
  assign _zz_9780 = ($signed(_zz_9781) >>> _zz_594);
  assign _zz_9781 = _zz_9782;
  assign _zz_9782 = ($signed(_zz_9784) - $signed(_zz_591));
  assign _zz_9783 = ({8'd0,data_mid_108_real} <<< 8);
  assign _zz_9784 = {{8{_zz_9783[23]}}, _zz_9783};
  assign _zz_9785 = fixTo_710_dout;
  assign _zz_9786 = _zz_9787[31 : 0];
  assign _zz_9787 = _zz_9788;
  assign _zz_9788 = ($signed(_zz_9789) >>> _zz_594);
  assign _zz_9789 = _zz_9790;
  assign _zz_9790 = ($signed(_zz_9792) - $signed(_zz_592));
  assign _zz_9791 = ({8'd0,data_mid_108_imag} <<< 8);
  assign _zz_9792 = {{8{_zz_9791[23]}}, _zz_9791};
  assign _zz_9793 = fixTo_711_dout;
  assign _zz_9794 = _zz_9795[31 : 0];
  assign _zz_9795 = _zz_9796;
  assign _zz_9796 = ($signed(_zz_9797) >>> _zz_595);
  assign _zz_9797 = _zz_9798;
  assign _zz_9798 = ($signed(_zz_9800) + $signed(_zz_591));
  assign _zz_9799 = ({8'd0,data_mid_108_real} <<< 8);
  assign _zz_9800 = {{8{_zz_9799[23]}}, _zz_9799};
  assign _zz_9801 = fixTo_712_dout;
  assign _zz_9802 = _zz_9803[31 : 0];
  assign _zz_9803 = _zz_9804;
  assign _zz_9804 = ($signed(_zz_9805) >>> _zz_595);
  assign _zz_9805 = _zz_9806;
  assign _zz_9806 = ($signed(_zz_9808) + $signed(_zz_592));
  assign _zz_9807 = ({8'd0,data_mid_108_imag} <<< 8);
  assign _zz_9808 = {{8{_zz_9807[23]}}, _zz_9807};
  assign _zz_9809 = fixTo_713_dout;
  assign _zz_9810 = ($signed(twiddle_factor_table_2_real) + $signed(twiddle_factor_table_2_imag));
  assign _zz_9811 = ($signed(_zz_598) - $signed(_zz_9812));
  assign _zz_9812 = ($signed(_zz_9813) * $signed(twiddle_factor_table_2_imag));
  assign _zz_9813 = ($signed(data_mid_111_real) + $signed(data_mid_111_imag));
  assign _zz_9814 = fixTo_714_dout;
  assign _zz_9815 = ($signed(_zz_598) + $signed(_zz_9816));
  assign _zz_9816 = ($signed(_zz_9817) * $signed(twiddle_factor_table_2_real));
  assign _zz_9817 = ($signed(data_mid_111_imag) - $signed(data_mid_111_real));
  assign _zz_9818 = fixTo_715_dout;
  assign _zz_9819 = _zz_9820[31 : 0];
  assign _zz_9820 = _zz_9821;
  assign _zz_9821 = ($signed(_zz_9822) >>> _zz_599);
  assign _zz_9822 = _zz_9823;
  assign _zz_9823 = ($signed(_zz_9825) - $signed(_zz_596));
  assign _zz_9824 = ({8'd0,data_mid_109_real} <<< 8);
  assign _zz_9825 = {{8{_zz_9824[23]}}, _zz_9824};
  assign _zz_9826 = fixTo_716_dout;
  assign _zz_9827 = _zz_9828[31 : 0];
  assign _zz_9828 = _zz_9829;
  assign _zz_9829 = ($signed(_zz_9830) >>> _zz_599);
  assign _zz_9830 = _zz_9831;
  assign _zz_9831 = ($signed(_zz_9833) - $signed(_zz_597));
  assign _zz_9832 = ({8'd0,data_mid_109_imag} <<< 8);
  assign _zz_9833 = {{8{_zz_9832[23]}}, _zz_9832};
  assign _zz_9834 = fixTo_717_dout;
  assign _zz_9835 = _zz_9836[31 : 0];
  assign _zz_9836 = _zz_9837;
  assign _zz_9837 = ($signed(_zz_9838) >>> _zz_600);
  assign _zz_9838 = _zz_9839;
  assign _zz_9839 = ($signed(_zz_9841) + $signed(_zz_596));
  assign _zz_9840 = ({8'd0,data_mid_109_real} <<< 8);
  assign _zz_9841 = {{8{_zz_9840[23]}}, _zz_9840};
  assign _zz_9842 = fixTo_718_dout;
  assign _zz_9843 = _zz_9844[31 : 0];
  assign _zz_9844 = _zz_9845;
  assign _zz_9845 = ($signed(_zz_9846) >>> _zz_600);
  assign _zz_9846 = _zz_9847;
  assign _zz_9847 = ($signed(_zz_9849) + $signed(_zz_597));
  assign _zz_9848 = ({8'd0,data_mid_109_imag} <<< 8);
  assign _zz_9849 = {{8{_zz_9848[23]}}, _zz_9848};
  assign _zz_9850 = fixTo_719_dout;
  assign _zz_9851 = ($signed(twiddle_factor_table_1_real) + $signed(twiddle_factor_table_1_imag));
  assign _zz_9852 = ($signed(_zz_603) - $signed(_zz_9853));
  assign _zz_9853 = ($signed(_zz_9854) * $signed(twiddle_factor_table_1_imag));
  assign _zz_9854 = ($signed(data_mid_114_real) + $signed(data_mid_114_imag));
  assign _zz_9855 = fixTo_720_dout;
  assign _zz_9856 = ($signed(_zz_603) + $signed(_zz_9857));
  assign _zz_9857 = ($signed(_zz_9858) * $signed(twiddle_factor_table_1_real));
  assign _zz_9858 = ($signed(data_mid_114_imag) - $signed(data_mid_114_real));
  assign _zz_9859 = fixTo_721_dout;
  assign _zz_9860 = _zz_9861[31 : 0];
  assign _zz_9861 = _zz_9862;
  assign _zz_9862 = ($signed(_zz_9863) >>> _zz_604);
  assign _zz_9863 = _zz_9864;
  assign _zz_9864 = ($signed(_zz_9866) - $signed(_zz_601));
  assign _zz_9865 = ({8'd0,data_mid_112_real} <<< 8);
  assign _zz_9866 = {{8{_zz_9865[23]}}, _zz_9865};
  assign _zz_9867 = fixTo_722_dout;
  assign _zz_9868 = _zz_9869[31 : 0];
  assign _zz_9869 = _zz_9870;
  assign _zz_9870 = ($signed(_zz_9871) >>> _zz_604);
  assign _zz_9871 = _zz_9872;
  assign _zz_9872 = ($signed(_zz_9874) - $signed(_zz_602));
  assign _zz_9873 = ({8'd0,data_mid_112_imag} <<< 8);
  assign _zz_9874 = {{8{_zz_9873[23]}}, _zz_9873};
  assign _zz_9875 = fixTo_723_dout;
  assign _zz_9876 = _zz_9877[31 : 0];
  assign _zz_9877 = _zz_9878;
  assign _zz_9878 = ($signed(_zz_9879) >>> _zz_605);
  assign _zz_9879 = _zz_9880;
  assign _zz_9880 = ($signed(_zz_9882) + $signed(_zz_601));
  assign _zz_9881 = ({8'd0,data_mid_112_real} <<< 8);
  assign _zz_9882 = {{8{_zz_9881[23]}}, _zz_9881};
  assign _zz_9883 = fixTo_724_dout;
  assign _zz_9884 = _zz_9885[31 : 0];
  assign _zz_9885 = _zz_9886;
  assign _zz_9886 = ($signed(_zz_9887) >>> _zz_605);
  assign _zz_9887 = _zz_9888;
  assign _zz_9888 = ($signed(_zz_9890) + $signed(_zz_602));
  assign _zz_9889 = ({8'd0,data_mid_112_imag} <<< 8);
  assign _zz_9890 = {{8{_zz_9889[23]}}, _zz_9889};
  assign _zz_9891 = fixTo_725_dout;
  assign _zz_9892 = ($signed(twiddle_factor_table_2_real) + $signed(twiddle_factor_table_2_imag));
  assign _zz_9893 = ($signed(_zz_608) - $signed(_zz_9894));
  assign _zz_9894 = ($signed(_zz_9895) * $signed(twiddle_factor_table_2_imag));
  assign _zz_9895 = ($signed(data_mid_115_real) + $signed(data_mid_115_imag));
  assign _zz_9896 = fixTo_726_dout;
  assign _zz_9897 = ($signed(_zz_608) + $signed(_zz_9898));
  assign _zz_9898 = ($signed(_zz_9899) * $signed(twiddle_factor_table_2_real));
  assign _zz_9899 = ($signed(data_mid_115_imag) - $signed(data_mid_115_real));
  assign _zz_9900 = fixTo_727_dout;
  assign _zz_9901 = _zz_9902[31 : 0];
  assign _zz_9902 = _zz_9903;
  assign _zz_9903 = ($signed(_zz_9904) >>> _zz_609);
  assign _zz_9904 = _zz_9905;
  assign _zz_9905 = ($signed(_zz_9907) - $signed(_zz_606));
  assign _zz_9906 = ({8'd0,data_mid_113_real} <<< 8);
  assign _zz_9907 = {{8{_zz_9906[23]}}, _zz_9906};
  assign _zz_9908 = fixTo_728_dout;
  assign _zz_9909 = _zz_9910[31 : 0];
  assign _zz_9910 = _zz_9911;
  assign _zz_9911 = ($signed(_zz_9912) >>> _zz_609);
  assign _zz_9912 = _zz_9913;
  assign _zz_9913 = ($signed(_zz_9915) - $signed(_zz_607));
  assign _zz_9914 = ({8'd0,data_mid_113_imag} <<< 8);
  assign _zz_9915 = {{8{_zz_9914[23]}}, _zz_9914};
  assign _zz_9916 = fixTo_729_dout;
  assign _zz_9917 = _zz_9918[31 : 0];
  assign _zz_9918 = _zz_9919;
  assign _zz_9919 = ($signed(_zz_9920) >>> _zz_610);
  assign _zz_9920 = _zz_9921;
  assign _zz_9921 = ($signed(_zz_9923) + $signed(_zz_606));
  assign _zz_9922 = ({8'd0,data_mid_113_real} <<< 8);
  assign _zz_9923 = {{8{_zz_9922[23]}}, _zz_9922};
  assign _zz_9924 = fixTo_730_dout;
  assign _zz_9925 = _zz_9926[31 : 0];
  assign _zz_9926 = _zz_9927;
  assign _zz_9927 = ($signed(_zz_9928) >>> _zz_610);
  assign _zz_9928 = _zz_9929;
  assign _zz_9929 = ($signed(_zz_9931) + $signed(_zz_607));
  assign _zz_9930 = ({8'd0,data_mid_113_imag} <<< 8);
  assign _zz_9931 = {{8{_zz_9930[23]}}, _zz_9930};
  assign _zz_9932 = fixTo_731_dout;
  assign _zz_9933 = ($signed(twiddle_factor_table_1_real) + $signed(twiddle_factor_table_1_imag));
  assign _zz_9934 = ($signed(_zz_613) - $signed(_zz_9935));
  assign _zz_9935 = ($signed(_zz_9936) * $signed(twiddle_factor_table_1_imag));
  assign _zz_9936 = ($signed(data_mid_118_real) + $signed(data_mid_118_imag));
  assign _zz_9937 = fixTo_732_dout;
  assign _zz_9938 = ($signed(_zz_613) + $signed(_zz_9939));
  assign _zz_9939 = ($signed(_zz_9940) * $signed(twiddle_factor_table_1_real));
  assign _zz_9940 = ($signed(data_mid_118_imag) - $signed(data_mid_118_real));
  assign _zz_9941 = fixTo_733_dout;
  assign _zz_9942 = _zz_9943[31 : 0];
  assign _zz_9943 = _zz_9944;
  assign _zz_9944 = ($signed(_zz_9945) >>> _zz_614);
  assign _zz_9945 = _zz_9946;
  assign _zz_9946 = ($signed(_zz_9948) - $signed(_zz_611));
  assign _zz_9947 = ({8'd0,data_mid_116_real} <<< 8);
  assign _zz_9948 = {{8{_zz_9947[23]}}, _zz_9947};
  assign _zz_9949 = fixTo_734_dout;
  assign _zz_9950 = _zz_9951[31 : 0];
  assign _zz_9951 = _zz_9952;
  assign _zz_9952 = ($signed(_zz_9953) >>> _zz_614);
  assign _zz_9953 = _zz_9954;
  assign _zz_9954 = ($signed(_zz_9956) - $signed(_zz_612));
  assign _zz_9955 = ({8'd0,data_mid_116_imag} <<< 8);
  assign _zz_9956 = {{8{_zz_9955[23]}}, _zz_9955};
  assign _zz_9957 = fixTo_735_dout;
  assign _zz_9958 = _zz_9959[31 : 0];
  assign _zz_9959 = _zz_9960;
  assign _zz_9960 = ($signed(_zz_9961) >>> _zz_615);
  assign _zz_9961 = _zz_9962;
  assign _zz_9962 = ($signed(_zz_9964) + $signed(_zz_611));
  assign _zz_9963 = ({8'd0,data_mid_116_real} <<< 8);
  assign _zz_9964 = {{8{_zz_9963[23]}}, _zz_9963};
  assign _zz_9965 = fixTo_736_dout;
  assign _zz_9966 = _zz_9967[31 : 0];
  assign _zz_9967 = _zz_9968;
  assign _zz_9968 = ($signed(_zz_9969) >>> _zz_615);
  assign _zz_9969 = _zz_9970;
  assign _zz_9970 = ($signed(_zz_9972) + $signed(_zz_612));
  assign _zz_9971 = ({8'd0,data_mid_116_imag} <<< 8);
  assign _zz_9972 = {{8{_zz_9971[23]}}, _zz_9971};
  assign _zz_9973 = fixTo_737_dout;
  assign _zz_9974 = ($signed(twiddle_factor_table_2_real) + $signed(twiddle_factor_table_2_imag));
  assign _zz_9975 = ($signed(_zz_618) - $signed(_zz_9976));
  assign _zz_9976 = ($signed(_zz_9977) * $signed(twiddle_factor_table_2_imag));
  assign _zz_9977 = ($signed(data_mid_119_real) + $signed(data_mid_119_imag));
  assign _zz_9978 = fixTo_738_dout;
  assign _zz_9979 = ($signed(_zz_618) + $signed(_zz_9980));
  assign _zz_9980 = ($signed(_zz_9981) * $signed(twiddle_factor_table_2_real));
  assign _zz_9981 = ($signed(data_mid_119_imag) - $signed(data_mid_119_real));
  assign _zz_9982 = fixTo_739_dout;
  assign _zz_9983 = _zz_9984[31 : 0];
  assign _zz_9984 = _zz_9985;
  assign _zz_9985 = ($signed(_zz_9986) >>> _zz_619);
  assign _zz_9986 = _zz_9987;
  assign _zz_9987 = ($signed(_zz_9989) - $signed(_zz_616));
  assign _zz_9988 = ({8'd0,data_mid_117_real} <<< 8);
  assign _zz_9989 = {{8{_zz_9988[23]}}, _zz_9988};
  assign _zz_9990 = fixTo_740_dout;
  assign _zz_9991 = _zz_9992[31 : 0];
  assign _zz_9992 = _zz_9993;
  assign _zz_9993 = ($signed(_zz_9994) >>> _zz_619);
  assign _zz_9994 = _zz_9995;
  assign _zz_9995 = ($signed(_zz_9997) - $signed(_zz_617));
  assign _zz_9996 = ({8'd0,data_mid_117_imag} <<< 8);
  assign _zz_9997 = {{8{_zz_9996[23]}}, _zz_9996};
  assign _zz_9998 = fixTo_741_dout;
  assign _zz_9999 = _zz_10000[31 : 0];
  assign _zz_10000 = _zz_10001;
  assign _zz_10001 = ($signed(_zz_10002) >>> _zz_620);
  assign _zz_10002 = _zz_10003;
  assign _zz_10003 = ($signed(_zz_10005) + $signed(_zz_616));
  assign _zz_10004 = ({8'd0,data_mid_117_real} <<< 8);
  assign _zz_10005 = {{8{_zz_10004[23]}}, _zz_10004};
  assign _zz_10006 = fixTo_742_dout;
  assign _zz_10007 = _zz_10008[31 : 0];
  assign _zz_10008 = _zz_10009;
  assign _zz_10009 = ($signed(_zz_10010) >>> _zz_620);
  assign _zz_10010 = _zz_10011;
  assign _zz_10011 = ($signed(_zz_10013) + $signed(_zz_617));
  assign _zz_10012 = ({8'd0,data_mid_117_imag} <<< 8);
  assign _zz_10013 = {{8{_zz_10012[23]}}, _zz_10012};
  assign _zz_10014 = fixTo_743_dout;
  assign _zz_10015 = ($signed(twiddle_factor_table_1_real) + $signed(twiddle_factor_table_1_imag));
  assign _zz_10016 = ($signed(_zz_623) - $signed(_zz_10017));
  assign _zz_10017 = ($signed(_zz_10018) * $signed(twiddle_factor_table_1_imag));
  assign _zz_10018 = ($signed(data_mid_122_real) + $signed(data_mid_122_imag));
  assign _zz_10019 = fixTo_744_dout;
  assign _zz_10020 = ($signed(_zz_623) + $signed(_zz_10021));
  assign _zz_10021 = ($signed(_zz_10022) * $signed(twiddle_factor_table_1_real));
  assign _zz_10022 = ($signed(data_mid_122_imag) - $signed(data_mid_122_real));
  assign _zz_10023 = fixTo_745_dout;
  assign _zz_10024 = _zz_10025[31 : 0];
  assign _zz_10025 = _zz_10026;
  assign _zz_10026 = ($signed(_zz_10027) >>> _zz_624);
  assign _zz_10027 = _zz_10028;
  assign _zz_10028 = ($signed(_zz_10030) - $signed(_zz_621));
  assign _zz_10029 = ({8'd0,data_mid_120_real} <<< 8);
  assign _zz_10030 = {{8{_zz_10029[23]}}, _zz_10029};
  assign _zz_10031 = fixTo_746_dout;
  assign _zz_10032 = _zz_10033[31 : 0];
  assign _zz_10033 = _zz_10034;
  assign _zz_10034 = ($signed(_zz_10035) >>> _zz_624);
  assign _zz_10035 = _zz_10036;
  assign _zz_10036 = ($signed(_zz_10038) - $signed(_zz_622));
  assign _zz_10037 = ({8'd0,data_mid_120_imag} <<< 8);
  assign _zz_10038 = {{8{_zz_10037[23]}}, _zz_10037};
  assign _zz_10039 = fixTo_747_dout;
  assign _zz_10040 = _zz_10041[31 : 0];
  assign _zz_10041 = _zz_10042;
  assign _zz_10042 = ($signed(_zz_10043) >>> _zz_625);
  assign _zz_10043 = _zz_10044;
  assign _zz_10044 = ($signed(_zz_10046) + $signed(_zz_621));
  assign _zz_10045 = ({8'd0,data_mid_120_real} <<< 8);
  assign _zz_10046 = {{8{_zz_10045[23]}}, _zz_10045};
  assign _zz_10047 = fixTo_748_dout;
  assign _zz_10048 = _zz_10049[31 : 0];
  assign _zz_10049 = _zz_10050;
  assign _zz_10050 = ($signed(_zz_10051) >>> _zz_625);
  assign _zz_10051 = _zz_10052;
  assign _zz_10052 = ($signed(_zz_10054) + $signed(_zz_622));
  assign _zz_10053 = ({8'd0,data_mid_120_imag} <<< 8);
  assign _zz_10054 = {{8{_zz_10053[23]}}, _zz_10053};
  assign _zz_10055 = fixTo_749_dout;
  assign _zz_10056 = ($signed(twiddle_factor_table_2_real) + $signed(twiddle_factor_table_2_imag));
  assign _zz_10057 = ($signed(_zz_628) - $signed(_zz_10058));
  assign _zz_10058 = ($signed(_zz_10059) * $signed(twiddle_factor_table_2_imag));
  assign _zz_10059 = ($signed(data_mid_123_real) + $signed(data_mid_123_imag));
  assign _zz_10060 = fixTo_750_dout;
  assign _zz_10061 = ($signed(_zz_628) + $signed(_zz_10062));
  assign _zz_10062 = ($signed(_zz_10063) * $signed(twiddle_factor_table_2_real));
  assign _zz_10063 = ($signed(data_mid_123_imag) - $signed(data_mid_123_real));
  assign _zz_10064 = fixTo_751_dout;
  assign _zz_10065 = _zz_10066[31 : 0];
  assign _zz_10066 = _zz_10067;
  assign _zz_10067 = ($signed(_zz_10068) >>> _zz_629);
  assign _zz_10068 = _zz_10069;
  assign _zz_10069 = ($signed(_zz_10071) - $signed(_zz_626));
  assign _zz_10070 = ({8'd0,data_mid_121_real} <<< 8);
  assign _zz_10071 = {{8{_zz_10070[23]}}, _zz_10070};
  assign _zz_10072 = fixTo_752_dout;
  assign _zz_10073 = _zz_10074[31 : 0];
  assign _zz_10074 = _zz_10075;
  assign _zz_10075 = ($signed(_zz_10076) >>> _zz_629);
  assign _zz_10076 = _zz_10077;
  assign _zz_10077 = ($signed(_zz_10079) - $signed(_zz_627));
  assign _zz_10078 = ({8'd0,data_mid_121_imag} <<< 8);
  assign _zz_10079 = {{8{_zz_10078[23]}}, _zz_10078};
  assign _zz_10080 = fixTo_753_dout;
  assign _zz_10081 = _zz_10082[31 : 0];
  assign _zz_10082 = _zz_10083;
  assign _zz_10083 = ($signed(_zz_10084) >>> _zz_630);
  assign _zz_10084 = _zz_10085;
  assign _zz_10085 = ($signed(_zz_10087) + $signed(_zz_626));
  assign _zz_10086 = ({8'd0,data_mid_121_real} <<< 8);
  assign _zz_10087 = {{8{_zz_10086[23]}}, _zz_10086};
  assign _zz_10088 = fixTo_754_dout;
  assign _zz_10089 = _zz_10090[31 : 0];
  assign _zz_10090 = _zz_10091;
  assign _zz_10091 = ($signed(_zz_10092) >>> _zz_630);
  assign _zz_10092 = _zz_10093;
  assign _zz_10093 = ($signed(_zz_10095) + $signed(_zz_627));
  assign _zz_10094 = ({8'd0,data_mid_121_imag} <<< 8);
  assign _zz_10095 = {{8{_zz_10094[23]}}, _zz_10094};
  assign _zz_10096 = fixTo_755_dout;
  assign _zz_10097 = ($signed(twiddle_factor_table_1_real) + $signed(twiddle_factor_table_1_imag));
  assign _zz_10098 = ($signed(_zz_633) - $signed(_zz_10099));
  assign _zz_10099 = ($signed(_zz_10100) * $signed(twiddle_factor_table_1_imag));
  assign _zz_10100 = ($signed(data_mid_126_real) + $signed(data_mid_126_imag));
  assign _zz_10101 = fixTo_756_dout;
  assign _zz_10102 = ($signed(_zz_633) + $signed(_zz_10103));
  assign _zz_10103 = ($signed(_zz_10104) * $signed(twiddle_factor_table_1_real));
  assign _zz_10104 = ($signed(data_mid_126_imag) - $signed(data_mid_126_real));
  assign _zz_10105 = fixTo_757_dout;
  assign _zz_10106 = _zz_10107[31 : 0];
  assign _zz_10107 = _zz_10108;
  assign _zz_10108 = ($signed(_zz_10109) >>> _zz_634);
  assign _zz_10109 = _zz_10110;
  assign _zz_10110 = ($signed(_zz_10112) - $signed(_zz_631));
  assign _zz_10111 = ({8'd0,data_mid_124_real} <<< 8);
  assign _zz_10112 = {{8{_zz_10111[23]}}, _zz_10111};
  assign _zz_10113 = fixTo_758_dout;
  assign _zz_10114 = _zz_10115[31 : 0];
  assign _zz_10115 = _zz_10116;
  assign _zz_10116 = ($signed(_zz_10117) >>> _zz_634);
  assign _zz_10117 = _zz_10118;
  assign _zz_10118 = ($signed(_zz_10120) - $signed(_zz_632));
  assign _zz_10119 = ({8'd0,data_mid_124_imag} <<< 8);
  assign _zz_10120 = {{8{_zz_10119[23]}}, _zz_10119};
  assign _zz_10121 = fixTo_759_dout;
  assign _zz_10122 = _zz_10123[31 : 0];
  assign _zz_10123 = _zz_10124;
  assign _zz_10124 = ($signed(_zz_10125) >>> _zz_635);
  assign _zz_10125 = _zz_10126;
  assign _zz_10126 = ($signed(_zz_10128) + $signed(_zz_631));
  assign _zz_10127 = ({8'd0,data_mid_124_real} <<< 8);
  assign _zz_10128 = {{8{_zz_10127[23]}}, _zz_10127};
  assign _zz_10129 = fixTo_760_dout;
  assign _zz_10130 = _zz_10131[31 : 0];
  assign _zz_10131 = _zz_10132;
  assign _zz_10132 = ($signed(_zz_10133) >>> _zz_635);
  assign _zz_10133 = _zz_10134;
  assign _zz_10134 = ($signed(_zz_10136) + $signed(_zz_632));
  assign _zz_10135 = ({8'd0,data_mid_124_imag} <<< 8);
  assign _zz_10136 = {{8{_zz_10135[23]}}, _zz_10135};
  assign _zz_10137 = fixTo_761_dout;
  assign _zz_10138 = ($signed(twiddle_factor_table_2_real) + $signed(twiddle_factor_table_2_imag));
  assign _zz_10139 = ($signed(_zz_638) - $signed(_zz_10140));
  assign _zz_10140 = ($signed(_zz_10141) * $signed(twiddle_factor_table_2_imag));
  assign _zz_10141 = ($signed(data_mid_127_real) + $signed(data_mid_127_imag));
  assign _zz_10142 = fixTo_762_dout;
  assign _zz_10143 = ($signed(_zz_638) + $signed(_zz_10144));
  assign _zz_10144 = ($signed(_zz_10145) * $signed(twiddle_factor_table_2_real));
  assign _zz_10145 = ($signed(data_mid_127_imag) - $signed(data_mid_127_real));
  assign _zz_10146 = fixTo_763_dout;
  assign _zz_10147 = _zz_10148[31 : 0];
  assign _zz_10148 = _zz_10149;
  assign _zz_10149 = ($signed(_zz_10150) >>> _zz_639);
  assign _zz_10150 = _zz_10151;
  assign _zz_10151 = ($signed(_zz_10153) - $signed(_zz_636));
  assign _zz_10152 = ({8'd0,data_mid_125_real} <<< 8);
  assign _zz_10153 = {{8{_zz_10152[23]}}, _zz_10152};
  assign _zz_10154 = fixTo_764_dout;
  assign _zz_10155 = _zz_10156[31 : 0];
  assign _zz_10156 = _zz_10157;
  assign _zz_10157 = ($signed(_zz_10158) >>> _zz_639);
  assign _zz_10158 = _zz_10159;
  assign _zz_10159 = ($signed(_zz_10161) - $signed(_zz_637));
  assign _zz_10160 = ({8'd0,data_mid_125_imag} <<< 8);
  assign _zz_10161 = {{8{_zz_10160[23]}}, _zz_10160};
  assign _zz_10162 = fixTo_765_dout;
  assign _zz_10163 = _zz_10164[31 : 0];
  assign _zz_10164 = _zz_10165;
  assign _zz_10165 = ($signed(_zz_10166) >>> _zz_640);
  assign _zz_10166 = _zz_10167;
  assign _zz_10167 = ($signed(_zz_10169) + $signed(_zz_636));
  assign _zz_10168 = ({8'd0,data_mid_125_real} <<< 8);
  assign _zz_10169 = {{8{_zz_10168[23]}}, _zz_10168};
  assign _zz_10170 = fixTo_766_dout;
  assign _zz_10171 = _zz_10172[31 : 0];
  assign _zz_10172 = _zz_10173;
  assign _zz_10173 = ($signed(_zz_10174) >>> _zz_640);
  assign _zz_10174 = _zz_10175;
  assign _zz_10175 = ($signed(_zz_10177) + $signed(_zz_637));
  assign _zz_10176 = ({8'd0,data_mid_125_imag} <<< 8);
  assign _zz_10177 = {{8{_zz_10176[23]}}, _zz_10176};
  assign _zz_10178 = fixTo_767_dout;
  assign _zz_10179 = ($signed(twiddle_factor_table_3_real) + $signed(twiddle_factor_table_3_imag));
  assign _zz_10180 = ($signed(_zz_643) - $signed(_zz_10181));
  assign _zz_10181 = ($signed(_zz_10182) * $signed(twiddle_factor_table_3_imag));
  assign _zz_10182 = ($signed(data_mid_4_real) + $signed(data_mid_4_imag));
  assign _zz_10183 = fixTo_768_dout;
  assign _zz_10184 = ($signed(_zz_643) + $signed(_zz_10185));
  assign _zz_10185 = ($signed(_zz_10186) * $signed(twiddle_factor_table_3_real));
  assign _zz_10186 = ($signed(data_mid_4_imag) - $signed(data_mid_4_real));
  assign _zz_10187 = fixTo_769_dout;
  assign _zz_10188 = _zz_10189[31 : 0];
  assign _zz_10189 = _zz_10190;
  assign _zz_10190 = ($signed(_zz_10191) >>> _zz_644);
  assign _zz_10191 = _zz_10192;
  assign _zz_10192 = ($signed(_zz_10194) - $signed(_zz_641));
  assign _zz_10193 = ({8'd0,data_mid_0_real} <<< 8);
  assign _zz_10194 = {{8{_zz_10193[23]}}, _zz_10193};
  assign _zz_10195 = fixTo_770_dout;
  assign _zz_10196 = _zz_10197[31 : 0];
  assign _zz_10197 = _zz_10198;
  assign _zz_10198 = ($signed(_zz_10199) >>> _zz_644);
  assign _zz_10199 = _zz_10200;
  assign _zz_10200 = ($signed(_zz_10202) - $signed(_zz_642));
  assign _zz_10201 = ({8'd0,data_mid_0_imag} <<< 8);
  assign _zz_10202 = {{8{_zz_10201[23]}}, _zz_10201};
  assign _zz_10203 = fixTo_771_dout;
  assign _zz_10204 = _zz_10205[31 : 0];
  assign _zz_10205 = _zz_10206;
  assign _zz_10206 = ($signed(_zz_10207) >>> _zz_645);
  assign _zz_10207 = _zz_10208;
  assign _zz_10208 = ($signed(_zz_10210) + $signed(_zz_641));
  assign _zz_10209 = ({8'd0,data_mid_0_real} <<< 8);
  assign _zz_10210 = {{8{_zz_10209[23]}}, _zz_10209};
  assign _zz_10211 = fixTo_772_dout;
  assign _zz_10212 = _zz_10213[31 : 0];
  assign _zz_10213 = _zz_10214;
  assign _zz_10214 = ($signed(_zz_10215) >>> _zz_645);
  assign _zz_10215 = _zz_10216;
  assign _zz_10216 = ($signed(_zz_10218) + $signed(_zz_642));
  assign _zz_10217 = ({8'd0,data_mid_0_imag} <<< 8);
  assign _zz_10218 = {{8{_zz_10217[23]}}, _zz_10217};
  assign _zz_10219 = fixTo_773_dout;
  assign _zz_10220 = ($signed(twiddle_factor_table_4_real) + $signed(twiddle_factor_table_4_imag));
  assign _zz_10221 = ($signed(_zz_648) - $signed(_zz_10222));
  assign _zz_10222 = ($signed(_zz_10223) * $signed(twiddle_factor_table_4_imag));
  assign _zz_10223 = ($signed(data_mid_5_real) + $signed(data_mid_5_imag));
  assign _zz_10224 = fixTo_774_dout;
  assign _zz_10225 = ($signed(_zz_648) + $signed(_zz_10226));
  assign _zz_10226 = ($signed(_zz_10227) * $signed(twiddle_factor_table_4_real));
  assign _zz_10227 = ($signed(data_mid_5_imag) - $signed(data_mid_5_real));
  assign _zz_10228 = fixTo_775_dout;
  assign _zz_10229 = _zz_10230[31 : 0];
  assign _zz_10230 = _zz_10231;
  assign _zz_10231 = ($signed(_zz_10232) >>> _zz_649);
  assign _zz_10232 = _zz_10233;
  assign _zz_10233 = ($signed(_zz_10235) - $signed(_zz_646));
  assign _zz_10234 = ({8'd0,data_mid_1_real} <<< 8);
  assign _zz_10235 = {{8{_zz_10234[23]}}, _zz_10234};
  assign _zz_10236 = fixTo_776_dout;
  assign _zz_10237 = _zz_10238[31 : 0];
  assign _zz_10238 = _zz_10239;
  assign _zz_10239 = ($signed(_zz_10240) >>> _zz_649);
  assign _zz_10240 = _zz_10241;
  assign _zz_10241 = ($signed(_zz_10243) - $signed(_zz_647));
  assign _zz_10242 = ({8'd0,data_mid_1_imag} <<< 8);
  assign _zz_10243 = {{8{_zz_10242[23]}}, _zz_10242};
  assign _zz_10244 = fixTo_777_dout;
  assign _zz_10245 = _zz_10246[31 : 0];
  assign _zz_10246 = _zz_10247;
  assign _zz_10247 = ($signed(_zz_10248) >>> _zz_650);
  assign _zz_10248 = _zz_10249;
  assign _zz_10249 = ($signed(_zz_10251) + $signed(_zz_646));
  assign _zz_10250 = ({8'd0,data_mid_1_real} <<< 8);
  assign _zz_10251 = {{8{_zz_10250[23]}}, _zz_10250};
  assign _zz_10252 = fixTo_778_dout;
  assign _zz_10253 = _zz_10254[31 : 0];
  assign _zz_10254 = _zz_10255;
  assign _zz_10255 = ($signed(_zz_10256) >>> _zz_650);
  assign _zz_10256 = _zz_10257;
  assign _zz_10257 = ($signed(_zz_10259) + $signed(_zz_647));
  assign _zz_10258 = ({8'd0,data_mid_1_imag} <<< 8);
  assign _zz_10259 = {{8{_zz_10258[23]}}, _zz_10258};
  assign _zz_10260 = fixTo_779_dout;
  assign _zz_10261 = ($signed(twiddle_factor_table_5_real) + $signed(twiddle_factor_table_5_imag));
  assign _zz_10262 = ($signed(_zz_653) - $signed(_zz_10263));
  assign _zz_10263 = ($signed(_zz_10264) * $signed(twiddle_factor_table_5_imag));
  assign _zz_10264 = ($signed(data_mid_6_real) + $signed(data_mid_6_imag));
  assign _zz_10265 = fixTo_780_dout;
  assign _zz_10266 = ($signed(_zz_653) + $signed(_zz_10267));
  assign _zz_10267 = ($signed(_zz_10268) * $signed(twiddle_factor_table_5_real));
  assign _zz_10268 = ($signed(data_mid_6_imag) - $signed(data_mid_6_real));
  assign _zz_10269 = fixTo_781_dout;
  assign _zz_10270 = _zz_10271[31 : 0];
  assign _zz_10271 = _zz_10272;
  assign _zz_10272 = ($signed(_zz_10273) >>> _zz_654);
  assign _zz_10273 = _zz_10274;
  assign _zz_10274 = ($signed(_zz_10276) - $signed(_zz_651));
  assign _zz_10275 = ({8'd0,data_mid_2_real} <<< 8);
  assign _zz_10276 = {{8{_zz_10275[23]}}, _zz_10275};
  assign _zz_10277 = fixTo_782_dout;
  assign _zz_10278 = _zz_10279[31 : 0];
  assign _zz_10279 = _zz_10280;
  assign _zz_10280 = ($signed(_zz_10281) >>> _zz_654);
  assign _zz_10281 = _zz_10282;
  assign _zz_10282 = ($signed(_zz_10284) - $signed(_zz_652));
  assign _zz_10283 = ({8'd0,data_mid_2_imag} <<< 8);
  assign _zz_10284 = {{8{_zz_10283[23]}}, _zz_10283};
  assign _zz_10285 = fixTo_783_dout;
  assign _zz_10286 = _zz_10287[31 : 0];
  assign _zz_10287 = _zz_10288;
  assign _zz_10288 = ($signed(_zz_10289) >>> _zz_655);
  assign _zz_10289 = _zz_10290;
  assign _zz_10290 = ($signed(_zz_10292) + $signed(_zz_651));
  assign _zz_10291 = ({8'd0,data_mid_2_real} <<< 8);
  assign _zz_10292 = {{8{_zz_10291[23]}}, _zz_10291};
  assign _zz_10293 = fixTo_784_dout;
  assign _zz_10294 = _zz_10295[31 : 0];
  assign _zz_10295 = _zz_10296;
  assign _zz_10296 = ($signed(_zz_10297) >>> _zz_655);
  assign _zz_10297 = _zz_10298;
  assign _zz_10298 = ($signed(_zz_10300) + $signed(_zz_652));
  assign _zz_10299 = ({8'd0,data_mid_2_imag} <<< 8);
  assign _zz_10300 = {{8{_zz_10299[23]}}, _zz_10299};
  assign _zz_10301 = fixTo_785_dout;
  assign _zz_10302 = ($signed(twiddle_factor_table_6_real) + $signed(twiddle_factor_table_6_imag));
  assign _zz_10303 = ($signed(_zz_658) - $signed(_zz_10304));
  assign _zz_10304 = ($signed(_zz_10305) * $signed(twiddle_factor_table_6_imag));
  assign _zz_10305 = ($signed(data_mid_7_real) + $signed(data_mid_7_imag));
  assign _zz_10306 = fixTo_786_dout;
  assign _zz_10307 = ($signed(_zz_658) + $signed(_zz_10308));
  assign _zz_10308 = ($signed(_zz_10309) * $signed(twiddle_factor_table_6_real));
  assign _zz_10309 = ($signed(data_mid_7_imag) - $signed(data_mid_7_real));
  assign _zz_10310 = fixTo_787_dout;
  assign _zz_10311 = _zz_10312[31 : 0];
  assign _zz_10312 = _zz_10313;
  assign _zz_10313 = ($signed(_zz_10314) >>> _zz_659);
  assign _zz_10314 = _zz_10315;
  assign _zz_10315 = ($signed(_zz_10317) - $signed(_zz_656));
  assign _zz_10316 = ({8'd0,data_mid_3_real} <<< 8);
  assign _zz_10317 = {{8{_zz_10316[23]}}, _zz_10316};
  assign _zz_10318 = fixTo_788_dout;
  assign _zz_10319 = _zz_10320[31 : 0];
  assign _zz_10320 = _zz_10321;
  assign _zz_10321 = ($signed(_zz_10322) >>> _zz_659);
  assign _zz_10322 = _zz_10323;
  assign _zz_10323 = ($signed(_zz_10325) - $signed(_zz_657));
  assign _zz_10324 = ({8'd0,data_mid_3_imag} <<< 8);
  assign _zz_10325 = {{8{_zz_10324[23]}}, _zz_10324};
  assign _zz_10326 = fixTo_789_dout;
  assign _zz_10327 = _zz_10328[31 : 0];
  assign _zz_10328 = _zz_10329;
  assign _zz_10329 = ($signed(_zz_10330) >>> _zz_660);
  assign _zz_10330 = _zz_10331;
  assign _zz_10331 = ($signed(_zz_10333) + $signed(_zz_656));
  assign _zz_10332 = ({8'd0,data_mid_3_real} <<< 8);
  assign _zz_10333 = {{8{_zz_10332[23]}}, _zz_10332};
  assign _zz_10334 = fixTo_790_dout;
  assign _zz_10335 = _zz_10336[31 : 0];
  assign _zz_10336 = _zz_10337;
  assign _zz_10337 = ($signed(_zz_10338) >>> _zz_660);
  assign _zz_10338 = _zz_10339;
  assign _zz_10339 = ($signed(_zz_10341) + $signed(_zz_657));
  assign _zz_10340 = ({8'd0,data_mid_3_imag} <<< 8);
  assign _zz_10341 = {{8{_zz_10340[23]}}, _zz_10340};
  assign _zz_10342 = fixTo_791_dout;
  assign _zz_10343 = ($signed(twiddle_factor_table_3_real) + $signed(twiddle_factor_table_3_imag));
  assign _zz_10344 = ($signed(_zz_663) - $signed(_zz_10345));
  assign _zz_10345 = ($signed(_zz_10346) * $signed(twiddle_factor_table_3_imag));
  assign _zz_10346 = ($signed(data_mid_12_real) + $signed(data_mid_12_imag));
  assign _zz_10347 = fixTo_792_dout;
  assign _zz_10348 = ($signed(_zz_663) + $signed(_zz_10349));
  assign _zz_10349 = ($signed(_zz_10350) * $signed(twiddle_factor_table_3_real));
  assign _zz_10350 = ($signed(data_mid_12_imag) - $signed(data_mid_12_real));
  assign _zz_10351 = fixTo_793_dout;
  assign _zz_10352 = _zz_10353[31 : 0];
  assign _zz_10353 = _zz_10354;
  assign _zz_10354 = ($signed(_zz_10355) >>> _zz_664);
  assign _zz_10355 = _zz_10356;
  assign _zz_10356 = ($signed(_zz_10358) - $signed(_zz_661));
  assign _zz_10357 = ({8'd0,data_mid_8_real} <<< 8);
  assign _zz_10358 = {{8{_zz_10357[23]}}, _zz_10357};
  assign _zz_10359 = fixTo_794_dout;
  assign _zz_10360 = _zz_10361[31 : 0];
  assign _zz_10361 = _zz_10362;
  assign _zz_10362 = ($signed(_zz_10363) >>> _zz_664);
  assign _zz_10363 = _zz_10364;
  assign _zz_10364 = ($signed(_zz_10366) - $signed(_zz_662));
  assign _zz_10365 = ({8'd0,data_mid_8_imag} <<< 8);
  assign _zz_10366 = {{8{_zz_10365[23]}}, _zz_10365};
  assign _zz_10367 = fixTo_795_dout;
  assign _zz_10368 = _zz_10369[31 : 0];
  assign _zz_10369 = _zz_10370;
  assign _zz_10370 = ($signed(_zz_10371) >>> _zz_665);
  assign _zz_10371 = _zz_10372;
  assign _zz_10372 = ($signed(_zz_10374) + $signed(_zz_661));
  assign _zz_10373 = ({8'd0,data_mid_8_real} <<< 8);
  assign _zz_10374 = {{8{_zz_10373[23]}}, _zz_10373};
  assign _zz_10375 = fixTo_796_dout;
  assign _zz_10376 = _zz_10377[31 : 0];
  assign _zz_10377 = _zz_10378;
  assign _zz_10378 = ($signed(_zz_10379) >>> _zz_665);
  assign _zz_10379 = _zz_10380;
  assign _zz_10380 = ($signed(_zz_10382) + $signed(_zz_662));
  assign _zz_10381 = ({8'd0,data_mid_8_imag} <<< 8);
  assign _zz_10382 = {{8{_zz_10381[23]}}, _zz_10381};
  assign _zz_10383 = fixTo_797_dout;
  assign _zz_10384 = ($signed(twiddle_factor_table_4_real) + $signed(twiddle_factor_table_4_imag));
  assign _zz_10385 = ($signed(_zz_668) - $signed(_zz_10386));
  assign _zz_10386 = ($signed(_zz_10387) * $signed(twiddle_factor_table_4_imag));
  assign _zz_10387 = ($signed(data_mid_13_real) + $signed(data_mid_13_imag));
  assign _zz_10388 = fixTo_798_dout;
  assign _zz_10389 = ($signed(_zz_668) + $signed(_zz_10390));
  assign _zz_10390 = ($signed(_zz_10391) * $signed(twiddle_factor_table_4_real));
  assign _zz_10391 = ($signed(data_mid_13_imag) - $signed(data_mid_13_real));
  assign _zz_10392 = fixTo_799_dout;
  assign _zz_10393 = _zz_10394[31 : 0];
  assign _zz_10394 = _zz_10395;
  assign _zz_10395 = ($signed(_zz_10396) >>> _zz_669);
  assign _zz_10396 = _zz_10397;
  assign _zz_10397 = ($signed(_zz_10399) - $signed(_zz_666));
  assign _zz_10398 = ({8'd0,data_mid_9_real} <<< 8);
  assign _zz_10399 = {{8{_zz_10398[23]}}, _zz_10398};
  assign _zz_10400 = fixTo_800_dout;
  assign _zz_10401 = _zz_10402[31 : 0];
  assign _zz_10402 = _zz_10403;
  assign _zz_10403 = ($signed(_zz_10404) >>> _zz_669);
  assign _zz_10404 = _zz_10405;
  assign _zz_10405 = ($signed(_zz_10407) - $signed(_zz_667));
  assign _zz_10406 = ({8'd0,data_mid_9_imag} <<< 8);
  assign _zz_10407 = {{8{_zz_10406[23]}}, _zz_10406};
  assign _zz_10408 = fixTo_801_dout;
  assign _zz_10409 = _zz_10410[31 : 0];
  assign _zz_10410 = _zz_10411;
  assign _zz_10411 = ($signed(_zz_10412) >>> _zz_670);
  assign _zz_10412 = _zz_10413;
  assign _zz_10413 = ($signed(_zz_10415) + $signed(_zz_666));
  assign _zz_10414 = ({8'd0,data_mid_9_real} <<< 8);
  assign _zz_10415 = {{8{_zz_10414[23]}}, _zz_10414};
  assign _zz_10416 = fixTo_802_dout;
  assign _zz_10417 = _zz_10418[31 : 0];
  assign _zz_10418 = _zz_10419;
  assign _zz_10419 = ($signed(_zz_10420) >>> _zz_670);
  assign _zz_10420 = _zz_10421;
  assign _zz_10421 = ($signed(_zz_10423) + $signed(_zz_667));
  assign _zz_10422 = ({8'd0,data_mid_9_imag} <<< 8);
  assign _zz_10423 = {{8{_zz_10422[23]}}, _zz_10422};
  assign _zz_10424 = fixTo_803_dout;
  assign _zz_10425 = ($signed(twiddle_factor_table_5_real) + $signed(twiddle_factor_table_5_imag));
  assign _zz_10426 = ($signed(_zz_673) - $signed(_zz_10427));
  assign _zz_10427 = ($signed(_zz_10428) * $signed(twiddle_factor_table_5_imag));
  assign _zz_10428 = ($signed(data_mid_14_real) + $signed(data_mid_14_imag));
  assign _zz_10429 = fixTo_804_dout;
  assign _zz_10430 = ($signed(_zz_673) + $signed(_zz_10431));
  assign _zz_10431 = ($signed(_zz_10432) * $signed(twiddle_factor_table_5_real));
  assign _zz_10432 = ($signed(data_mid_14_imag) - $signed(data_mid_14_real));
  assign _zz_10433 = fixTo_805_dout;
  assign _zz_10434 = _zz_10435[31 : 0];
  assign _zz_10435 = _zz_10436;
  assign _zz_10436 = ($signed(_zz_10437) >>> _zz_674);
  assign _zz_10437 = _zz_10438;
  assign _zz_10438 = ($signed(_zz_10440) - $signed(_zz_671));
  assign _zz_10439 = ({8'd0,data_mid_10_real} <<< 8);
  assign _zz_10440 = {{8{_zz_10439[23]}}, _zz_10439};
  assign _zz_10441 = fixTo_806_dout;
  assign _zz_10442 = _zz_10443[31 : 0];
  assign _zz_10443 = _zz_10444;
  assign _zz_10444 = ($signed(_zz_10445) >>> _zz_674);
  assign _zz_10445 = _zz_10446;
  assign _zz_10446 = ($signed(_zz_10448) - $signed(_zz_672));
  assign _zz_10447 = ({8'd0,data_mid_10_imag} <<< 8);
  assign _zz_10448 = {{8{_zz_10447[23]}}, _zz_10447};
  assign _zz_10449 = fixTo_807_dout;
  assign _zz_10450 = _zz_10451[31 : 0];
  assign _zz_10451 = _zz_10452;
  assign _zz_10452 = ($signed(_zz_10453) >>> _zz_675);
  assign _zz_10453 = _zz_10454;
  assign _zz_10454 = ($signed(_zz_10456) + $signed(_zz_671));
  assign _zz_10455 = ({8'd0,data_mid_10_real} <<< 8);
  assign _zz_10456 = {{8{_zz_10455[23]}}, _zz_10455};
  assign _zz_10457 = fixTo_808_dout;
  assign _zz_10458 = _zz_10459[31 : 0];
  assign _zz_10459 = _zz_10460;
  assign _zz_10460 = ($signed(_zz_10461) >>> _zz_675);
  assign _zz_10461 = _zz_10462;
  assign _zz_10462 = ($signed(_zz_10464) + $signed(_zz_672));
  assign _zz_10463 = ({8'd0,data_mid_10_imag} <<< 8);
  assign _zz_10464 = {{8{_zz_10463[23]}}, _zz_10463};
  assign _zz_10465 = fixTo_809_dout;
  assign _zz_10466 = ($signed(twiddle_factor_table_6_real) + $signed(twiddle_factor_table_6_imag));
  assign _zz_10467 = ($signed(_zz_678) - $signed(_zz_10468));
  assign _zz_10468 = ($signed(_zz_10469) * $signed(twiddle_factor_table_6_imag));
  assign _zz_10469 = ($signed(data_mid_15_real) + $signed(data_mid_15_imag));
  assign _zz_10470 = fixTo_810_dout;
  assign _zz_10471 = ($signed(_zz_678) + $signed(_zz_10472));
  assign _zz_10472 = ($signed(_zz_10473) * $signed(twiddle_factor_table_6_real));
  assign _zz_10473 = ($signed(data_mid_15_imag) - $signed(data_mid_15_real));
  assign _zz_10474 = fixTo_811_dout;
  assign _zz_10475 = _zz_10476[31 : 0];
  assign _zz_10476 = _zz_10477;
  assign _zz_10477 = ($signed(_zz_10478) >>> _zz_679);
  assign _zz_10478 = _zz_10479;
  assign _zz_10479 = ($signed(_zz_10481) - $signed(_zz_676));
  assign _zz_10480 = ({8'd0,data_mid_11_real} <<< 8);
  assign _zz_10481 = {{8{_zz_10480[23]}}, _zz_10480};
  assign _zz_10482 = fixTo_812_dout;
  assign _zz_10483 = _zz_10484[31 : 0];
  assign _zz_10484 = _zz_10485;
  assign _zz_10485 = ($signed(_zz_10486) >>> _zz_679);
  assign _zz_10486 = _zz_10487;
  assign _zz_10487 = ($signed(_zz_10489) - $signed(_zz_677));
  assign _zz_10488 = ({8'd0,data_mid_11_imag} <<< 8);
  assign _zz_10489 = {{8{_zz_10488[23]}}, _zz_10488};
  assign _zz_10490 = fixTo_813_dout;
  assign _zz_10491 = _zz_10492[31 : 0];
  assign _zz_10492 = _zz_10493;
  assign _zz_10493 = ($signed(_zz_10494) >>> _zz_680);
  assign _zz_10494 = _zz_10495;
  assign _zz_10495 = ($signed(_zz_10497) + $signed(_zz_676));
  assign _zz_10496 = ({8'd0,data_mid_11_real} <<< 8);
  assign _zz_10497 = {{8{_zz_10496[23]}}, _zz_10496};
  assign _zz_10498 = fixTo_814_dout;
  assign _zz_10499 = _zz_10500[31 : 0];
  assign _zz_10500 = _zz_10501;
  assign _zz_10501 = ($signed(_zz_10502) >>> _zz_680);
  assign _zz_10502 = _zz_10503;
  assign _zz_10503 = ($signed(_zz_10505) + $signed(_zz_677));
  assign _zz_10504 = ({8'd0,data_mid_11_imag} <<< 8);
  assign _zz_10505 = {{8{_zz_10504[23]}}, _zz_10504};
  assign _zz_10506 = fixTo_815_dout;
  assign _zz_10507 = ($signed(twiddle_factor_table_3_real) + $signed(twiddle_factor_table_3_imag));
  assign _zz_10508 = ($signed(_zz_683) - $signed(_zz_10509));
  assign _zz_10509 = ($signed(_zz_10510) * $signed(twiddle_factor_table_3_imag));
  assign _zz_10510 = ($signed(data_mid_20_real) + $signed(data_mid_20_imag));
  assign _zz_10511 = fixTo_816_dout;
  assign _zz_10512 = ($signed(_zz_683) + $signed(_zz_10513));
  assign _zz_10513 = ($signed(_zz_10514) * $signed(twiddle_factor_table_3_real));
  assign _zz_10514 = ($signed(data_mid_20_imag) - $signed(data_mid_20_real));
  assign _zz_10515 = fixTo_817_dout;
  assign _zz_10516 = _zz_10517[31 : 0];
  assign _zz_10517 = _zz_10518;
  assign _zz_10518 = ($signed(_zz_10519) >>> _zz_684);
  assign _zz_10519 = _zz_10520;
  assign _zz_10520 = ($signed(_zz_10522) - $signed(_zz_681));
  assign _zz_10521 = ({8'd0,data_mid_16_real} <<< 8);
  assign _zz_10522 = {{8{_zz_10521[23]}}, _zz_10521};
  assign _zz_10523 = fixTo_818_dout;
  assign _zz_10524 = _zz_10525[31 : 0];
  assign _zz_10525 = _zz_10526;
  assign _zz_10526 = ($signed(_zz_10527) >>> _zz_684);
  assign _zz_10527 = _zz_10528;
  assign _zz_10528 = ($signed(_zz_10530) - $signed(_zz_682));
  assign _zz_10529 = ({8'd0,data_mid_16_imag} <<< 8);
  assign _zz_10530 = {{8{_zz_10529[23]}}, _zz_10529};
  assign _zz_10531 = fixTo_819_dout;
  assign _zz_10532 = _zz_10533[31 : 0];
  assign _zz_10533 = _zz_10534;
  assign _zz_10534 = ($signed(_zz_10535) >>> _zz_685);
  assign _zz_10535 = _zz_10536;
  assign _zz_10536 = ($signed(_zz_10538) + $signed(_zz_681));
  assign _zz_10537 = ({8'd0,data_mid_16_real} <<< 8);
  assign _zz_10538 = {{8{_zz_10537[23]}}, _zz_10537};
  assign _zz_10539 = fixTo_820_dout;
  assign _zz_10540 = _zz_10541[31 : 0];
  assign _zz_10541 = _zz_10542;
  assign _zz_10542 = ($signed(_zz_10543) >>> _zz_685);
  assign _zz_10543 = _zz_10544;
  assign _zz_10544 = ($signed(_zz_10546) + $signed(_zz_682));
  assign _zz_10545 = ({8'd0,data_mid_16_imag} <<< 8);
  assign _zz_10546 = {{8{_zz_10545[23]}}, _zz_10545};
  assign _zz_10547 = fixTo_821_dout;
  assign _zz_10548 = ($signed(twiddle_factor_table_4_real) + $signed(twiddle_factor_table_4_imag));
  assign _zz_10549 = ($signed(_zz_688) - $signed(_zz_10550));
  assign _zz_10550 = ($signed(_zz_10551) * $signed(twiddle_factor_table_4_imag));
  assign _zz_10551 = ($signed(data_mid_21_real) + $signed(data_mid_21_imag));
  assign _zz_10552 = fixTo_822_dout;
  assign _zz_10553 = ($signed(_zz_688) + $signed(_zz_10554));
  assign _zz_10554 = ($signed(_zz_10555) * $signed(twiddle_factor_table_4_real));
  assign _zz_10555 = ($signed(data_mid_21_imag) - $signed(data_mid_21_real));
  assign _zz_10556 = fixTo_823_dout;
  assign _zz_10557 = _zz_10558[31 : 0];
  assign _zz_10558 = _zz_10559;
  assign _zz_10559 = ($signed(_zz_10560) >>> _zz_689);
  assign _zz_10560 = _zz_10561;
  assign _zz_10561 = ($signed(_zz_10563) - $signed(_zz_686));
  assign _zz_10562 = ({8'd0,data_mid_17_real} <<< 8);
  assign _zz_10563 = {{8{_zz_10562[23]}}, _zz_10562};
  assign _zz_10564 = fixTo_824_dout;
  assign _zz_10565 = _zz_10566[31 : 0];
  assign _zz_10566 = _zz_10567;
  assign _zz_10567 = ($signed(_zz_10568) >>> _zz_689);
  assign _zz_10568 = _zz_10569;
  assign _zz_10569 = ($signed(_zz_10571) - $signed(_zz_687));
  assign _zz_10570 = ({8'd0,data_mid_17_imag} <<< 8);
  assign _zz_10571 = {{8{_zz_10570[23]}}, _zz_10570};
  assign _zz_10572 = fixTo_825_dout;
  assign _zz_10573 = _zz_10574[31 : 0];
  assign _zz_10574 = _zz_10575;
  assign _zz_10575 = ($signed(_zz_10576) >>> _zz_690);
  assign _zz_10576 = _zz_10577;
  assign _zz_10577 = ($signed(_zz_10579) + $signed(_zz_686));
  assign _zz_10578 = ({8'd0,data_mid_17_real} <<< 8);
  assign _zz_10579 = {{8{_zz_10578[23]}}, _zz_10578};
  assign _zz_10580 = fixTo_826_dout;
  assign _zz_10581 = _zz_10582[31 : 0];
  assign _zz_10582 = _zz_10583;
  assign _zz_10583 = ($signed(_zz_10584) >>> _zz_690);
  assign _zz_10584 = _zz_10585;
  assign _zz_10585 = ($signed(_zz_10587) + $signed(_zz_687));
  assign _zz_10586 = ({8'd0,data_mid_17_imag} <<< 8);
  assign _zz_10587 = {{8{_zz_10586[23]}}, _zz_10586};
  assign _zz_10588 = fixTo_827_dout;
  assign _zz_10589 = ($signed(twiddle_factor_table_5_real) + $signed(twiddle_factor_table_5_imag));
  assign _zz_10590 = ($signed(_zz_693) - $signed(_zz_10591));
  assign _zz_10591 = ($signed(_zz_10592) * $signed(twiddle_factor_table_5_imag));
  assign _zz_10592 = ($signed(data_mid_22_real) + $signed(data_mid_22_imag));
  assign _zz_10593 = fixTo_828_dout;
  assign _zz_10594 = ($signed(_zz_693) + $signed(_zz_10595));
  assign _zz_10595 = ($signed(_zz_10596) * $signed(twiddle_factor_table_5_real));
  assign _zz_10596 = ($signed(data_mid_22_imag) - $signed(data_mid_22_real));
  assign _zz_10597 = fixTo_829_dout;
  assign _zz_10598 = _zz_10599[31 : 0];
  assign _zz_10599 = _zz_10600;
  assign _zz_10600 = ($signed(_zz_10601) >>> _zz_694);
  assign _zz_10601 = _zz_10602;
  assign _zz_10602 = ($signed(_zz_10604) - $signed(_zz_691));
  assign _zz_10603 = ({8'd0,data_mid_18_real} <<< 8);
  assign _zz_10604 = {{8{_zz_10603[23]}}, _zz_10603};
  assign _zz_10605 = fixTo_830_dout;
  assign _zz_10606 = _zz_10607[31 : 0];
  assign _zz_10607 = _zz_10608;
  assign _zz_10608 = ($signed(_zz_10609) >>> _zz_694);
  assign _zz_10609 = _zz_10610;
  assign _zz_10610 = ($signed(_zz_10612) - $signed(_zz_692));
  assign _zz_10611 = ({8'd0,data_mid_18_imag} <<< 8);
  assign _zz_10612 = {{8{_zz_10611[23]}}, _zz_10611};
  assign _zz_10613 = fixTo_831_dout;
  assign _zz_10614 = _zz_10615[31 : 0];
  assign _zz_10615 = _zz_10616;
  assign _zz_10616 = ($signed(_zz_10617) >>> _zz_695);
  assign _zz_10617 = _zz_10618;
  assign _zz_10618 = ($signed(_zz_10620) + $signed(_zz_691));
  assign _zz_10619 = ({8'd0,data_mid_18_real} <<< 8);
  assign _zz_10620 = {{8{_zz_10619[23]}}, _zz_10619};
  assign _zz_10621 = fixTo_832_dout;
  assign _zz_10622 = _zz_10623[31 : 0];
  assign _zz_10623 = _zz_10624;
  assign _zz_10624 = ($signed(_zz_10625) >>> _zz_695);
  assign _zz_10625 = _zz_10626;
  assign _zz_10626 = ($signed(_zz_10628) + $signed(_zz_692));
  assign _zz_10627 = ({8'd0,data_mid_18_imag} <<< 8);
  assign _zz_10628 = {{8{_zz_10627[23]}}, _zz_10627};
  assign _zz_10629 = fixTo_833_dout;
  assign _zz_10630 = ($signed(twiddle_factor_table_6_real) + $signed(twiddle_factor_table_6_imag));
  assign _zz_10631 = ($signed(_zz_698) - $signed(_zz_10632));
  assign _zz_10632 = ($signed(_zz_10633) * $signed(twiddle_factor_table_6_imag));
  assign _zz_10633 = ($signed(data_mid_23_real) + $signed(data_mid_23_imag));
  assign _zz_10634 = fixTo_834_dout;
  assign _zz_10635 = ($signed(_zz_698) + $signed(_zz_10636));
  assign _zz_10636 = ($signed(_zz_10637) * $signed(twiddle_factor_table_6_real));
  assign _zz_10637 = ($signed(data_mid_23_imag) - $signed(data_mid_23_real));
  assign _zz_10638 = fixTo_835_dout;
  assign _zz_10639 = _zz_10640[31 : 0];
  assign _zz_10640 = _zz_10641;
  assign _zz_10641 = ($signed(_zz_10642) >>> _zz_699);
  assign _zz_10642 = _zz_10643;
  assign _zz_10643 = ($signed(_zz_10645) - $signed(_zz_696));
  assign _zz_10644 = ({8'd0,data_mid_19_real} <<< 8);
  assign _zz_10645 = {{8{_zz_10644[23]}}, _zz_10644};
  assign _zz_10646 = fixTo_836_dout;
  assign _zz_10647 = _zz_10648[31 : 0];
  assign _zz_10648 = _zz_10649;
  assign _zz_10649 = ($signed(_zz_10650) >>> _zz_699);
  assign _zz_10650 = _zz_10651;
  assign _zz_10651 = ($signed(_zz_10653) - $signed(_zz_697));
  assign _zz_10652 = ({8'd0,data_mid_19_imag} <<< 8);
  assign _zz_10653 = {{8{_zz_10652[23]}}, _zz_10652};
  assign _zz_10654 = fixTo_837_dout;
  assign _zz_10655 = _zz_10656[31 : 0];
  assign _zz_10656 = _zz_10657;
  assign _zz_10657 = ($signed(_zz_10658) >>> _zz_700);
  assign _zz_10658 = _zz_10659;
  assign _zz_10659 = ($signed(_zz_10661) + $signed(_zz_696));
  assign _zz_10660 = ({8'd0,data_mid_19_real} <<< 8);
  assign _zz_10661 = {{8{_zz_10660[23]}}, _zz_10660};
  assign _zz_10662 = fixTo_838_dout;
  assign _zz_10663 = _zz_10664[31 : 0];
  assign _zz_10664 = _zz_10665;
  assign _zz_10665 = ($signed(_zz_10666) >>> _zz_700);
  assign _zz_10666 = _zz_10667;
  assign _zz_10667 = ($signed(_zz_10669) + $signed(_zz_697));
  assign _zz_10668 = ({8'd0,data_mid_19_imag} <<< 8);
  assign _zz_10669 = {{8{_zz_10668[23]}}, _zz_10668};
  assign _zz_10670 = fixTo_839_dout;
  assign _zz_10671 = ($signed(twiddle_factor_table_3_real) + $signed(twiddle_factor_table_3_imag));
  assign _zz_10672 = ($signed(_zz_703) - $signed(_zz_10673));
  assign _zz_10673 = ($signed(_zz_10674) * $signed(twiddle_factor_table_3_imag));
  assign _zz_10674 = ($signed(data_mid_28_real) + $signed(data_mid_28_imag));
  assign _zz_10675 = fixTo_840_dout;
  assign _zz_10676 = ($signed(_zz_703) + $signed(_zz_10677));
  assign _zz_10677 = ($signed(_zz_10678) * $signed(twiddle_factor_table_3_real));
  assign _zz_10678 = ($signed(data_mid_28_imag) - $signed(data_mid_28_real));
  assign _zz_10679 = fixTo_841_dout;
  assign _zz_10680 = _zz_10681[31 : 0];
  assign _zz_10681 = _zz_10682;
  assign _zz_10682 = ($signed(_zz_10683) >>> _zz_704);
  assign _zz_10683 = _zz_10684;
  assign _zz_10684 = ($signed(_zz_10686) - $signed(_zz_701));
  assign _zz_10685 = ({8'd0,data_mid_24_real} <<< 8);
  assign _zz_10686 = {{8{_zz_10685[23]}}, _zz_10685};
  assign _zz_10687 = fixTo_842_dout;
  assign _zz_10688 = _zz_10689[31 : 0];
  assign _zz_10689 = _zz_10690;
  assign _zz_10690 = ($signed(_zz_10691) >>> _zz_704);
  assign _zz_10691 = _zz_10692;
  assign _zz_10692 = ($signed(_zz_10694) - $signed(_zz_702));
  assign _zz_10693 = ({8'd0,data_mid_24_imag} <<< 8);
  assign _zz_10694 = {{8{_zz_10693[23]}}, _zz_10693};
  assign _zz_10695 = fixTo_843_dout;
  assign _zz_10696 = _zz_10697[31 : 0];
  assign _zz_10697 = _zz_10698;
  assign _zz_10698 = ($signed(_zz_10699) >>> _zz_705);
  assign _zz_10699 = _zz_10700;
  assign _zz_10700 = ($signed(_zz_10702) + $signed(_zz_701));
  assign _zz_10701 = ({8'd0,data_mid_24_real} <<< 8);
  assign _zz_10702 = {{8{_zz_10701[23]}}, _zz_10701};
  assign _zz_10703 = fixTo_844_dout;
  assign _zz_10704 = _zz_10705[31 : 0];
  assign _zz_10705 = _zz_10706;
  assign _zz_10706 = ($signed(_zz_10707) >>> _zz_705);
  assign _zz_10707 = _zz_10708;
  assign _zz_10708 = ($signed(_zz_10710) + $signed(_zz_702));
  assign _zz_10709 = ({8'd0,data_mid_24_imag} <<< 8);
  assign _zz_10710 = {{8{_zz_10709[23]}}, _zz_10709};
  assign _zz_10711 = fixTo_845_dout;
  assign _zz_10712 = ($signed(twiddle_factor_table_4_real) + $signed(twiddle_factor_table_4_imag));
  assign _zz_10713 = ($signed(_zz_708) - $signed(_zz_10714));
  assign _zz_10714 = ($signed(_zz_10715) * $signed(twiddle_factor_table_4_imag));
  assign _zz_10715 = ($signed(data_mid_29_real) + $signed(data_mid_29_imag));
  assign _zz_10716 = fixTo_846_dout;
  assign _zz_10717 = ($signed(_zz_708) + $signed(_zz_10718));
  assign _zz_10718 = ($signed(_zz_10719) * $signed(twiddle_factor_table_4_real));
  assign _zz_10719 = ($signed(data_mid_29_imag) - $signed(data_mid_29_real));
  assign _zz_10720 = fixTo_847_dout;
  assign _zz_10721 = _zz_10722[31 : 0];
  assign _zz_10722 = _zz_10723;
  assign _zz_10723 = ($signed(_zz_10724) >>> _zz_709);
  assign _zz_10724 = _zz_10725;
  assign _zz_10725 = ($signed(_zz_10727) - $signed(_zz_706));
  assign _zz_10726 = ({8'd0,data_mid_25_real} <<< 8);
  assign _zz_10727 = {{8{_zz_10726[23]}}, _zz_10726};
  assign _zz_10728 = fixTo_848_dout;
  assign _zz_10729 = _zz_10730[31 : 0];
  assign _zz_10730 = _zz_10731;
  assign _zz_10731 = ($signed(_zz_10732) >>> _zz_709);
  assign _zz_10732 = _zz_10733;
  assign _zz_10733 = ($signed(_zz_10735) - $signed(_zz_707));
  assign _zz_10734 = ({8'd0,data_mid_25_imag} <<< 8);
  assign _zz_10735 = {{8{_zz_10734[23]}}, _zz_10734};
  assign _zz_10736 = fixTo_849_dout;
  assign _zz_10737 = _zz_10738[31 : 0];
  assign _zz_10738 = _zz_10739;
  assign _zz_10739 = ($signed(_zz_10740) >>> _zz_710);
  assign _zz_10740 = _zz_10741;
  assign _zz_10741 = ($signed(_zz_10743) + $signed(_zz_706));
  assign _zz_10742 = ({8'd0,data_mid_25_real} <<< 8);
  assign _zz_10743 = {{8{_zz_10742[23]}}, _zz_10742};
  assign _zz_10744 = fixTo_850_dout;
  assign _zz_10745 = _zz_10746[31 : 0];
  assign _zz_10746 = _zz_10747;
  assign _zz_10747 = ($signed(_zz_10748) >>> _zz_710);
  assign _zz_10748 = _zz_10749;
  assign _zz_10749 = ($signed(_zz_10751) + $signed(_zz_707));
  assign _zz_10750 = ({8'd0,data_mid_25_imag} <<< 8);
  assign _zz_10751 = {{8{_zz_10750[23]}}, _zz_10750};
  assign _zz_10752 = fixTo_851_dout;
  assign _zz_10753 = ($signed(twiddle_factor_table_5_real) + $signed(twiddle_factor_table_5_imag));
  assign _zz_10754 = ($signed(_zz_713) - $signed(_zz_10755));
  assign _zz_10755 = ($signed(_zz_10756) * $signed(twiddle_factor_table_5_imag));
  assign _zz_10756 = ($signed(data_mid_30_real) + $signed(data_mid_30_imag));
  assign _zz_10757 = fixTo_852_dout;
  assign _zz_10758 = ($signed(_zz_713) + $signed(_zz_10759));
  assign _zz_10759 = ($signed(_zz_10760) * $signed(twiddle_factor_table_5_real));
  assign _zz_10760 = ($signed(data_mid_30_imag) - $signed(data_mid_30_real));
  assign _zz_10761 = fixTo_853_dout;
  assign _zz_10762 = _zz_10763[31 : 0];
  assign _zz_10763 = _zz_10764;
  assign _zz_10764 = ($signed(_zz_10765) >>> _zz_714);
  assign _zz_10765 = _zz_10766;
  assign _zz_10766 = ($signed(_zz_10768) - $signed(_zz_711));
  assign _zz_10767 = ({8'd0,data_mid_26_real} <<< 8);
  assign _zz_10768 = {{8{_zz_10767[23]}}, _zz_10767};
  assign _zz_10769 = fixTo_854_dout;
  assign _zz_10770 = _zz_10771[31 : 0];
  assign _zz_10771 = _zz_10772;
  assign _zz_10772 = ($signed(_zz_10773) >>> _zz_714);
  assign _zz_10773 = _zz_10774;
  assign _zz_10774 = ($signed(_zz_10776) - $signed(_zz_712));
  assign _zz_10775 = ({8'd0,data_mid_26_imag} <<< 8);
  assign _zz_10776 = {{8{_zz_10775[23]}}, _zz_10775};
  assign _zz_10777 = fixTo_855_dout;
  assign _zz_10778 = _zz_10779[31 : 0];
  assign _zz_10779 = _zz_10780;
  assign _zz_10780 = ($signed(_zz_10781) >>> _zz_715);
  assign _zz_10781 = _zz_10782;
  assign _zz_10782 = ($signed(_zz_10784) + $signed(_zz_711));
  assign _zz_10783 = ({8'd0,data_mid_26_real} <<< 8);
  assign _zz_10784 = {{8{_zz_10783[23]}}, _zz_10783};
  assign _zz_10785 = fixTo_856_dout;
  assign _zz_10786 = _zz_10787[31 : 0];
  assign _zz_10787 = _zz_10788;
  assign _zz_10788 = ($signed(_zz_10789) >>> _zz_715);
  assign _zz_10789 = _zz_10790;
  assign _zz_10790 = ($signed(_zz_10792) + $signed(_zz_712));
  assign _zz_10791 = ({8'd0,data_mid_26_imag} <<< 8);
  assign _zz_10792 = {{8{_zz_10791[23]}}, _zz_10791};
  assign _zz_10793 = fixTo_857_dout;
  assign _zz_10794 = ($signed(twiddle_factor_table_6_real) + $signed(twiddle_factor_table_6_imag));
  assign _zz_10795 = ($signed(_zz_718) - $signed(_zz_10796));
  assign _zz_10796 = ($signed(_zz_10797) * $signed(twiddle_factor_table_6_imag));
  assign _zz_10797 = ($signed(data_mid_31_real) + $signed(data_mid_31_imag));
  assign _zz_10798 = fixTo_858_dout;
  assign _zz_10799 = ($signed(_zz_718) + $signed(_zz_10800));
  assign _zz_10800 = ($signed(_zz_10801) * $signed(twiddle_factor_table_6_real));
  assign _zz_10801 = ($signed(data_mid_31_imag) - $signed(data_mid_31_real));
  assign _zz_10802 = fixTo_859_dout;
  assign _zz_10803 = _zz_10804[31 : 0];
  assign _zz_10804 = _zz_10805;
  assign _zz_10805 = ($signed(_zz_10806) >>> _zz_719);
  assign _zz_10806 = _zz_10807;
  assign _zz_10807 = ($signed(_zz_10809) - $signed(_zz_716));
  assign _zz_10808 = ({8'd0,data_mid_27_real} <<< 8);
  assign _zz_10809 = {{8{_zz_10808[23]}}, _zz_10808};
  assign _zz_10810 = fixTo_860_dout;
  assign _zz_10811 = _zz_10812[31 : 0];
  assign _zz_10812 = _zz_10813;
  assign _zz_10813 = ($signed(_zz_10814) >>> _zz_719);
  assign _zz_10814 = _zz_10815;
  assign _zz_10815 = ($signed(_zz_10817) - $signed(_zz_717));
  assign _zz_10816 = ({8'd0,data_mid_27_imag} <<< 8);
  assign _zz_10817 = {{8{_zz_10816[23]}}, _zz_10816};
  assign _zz_10818 = fixTo_861_dout;
  assign _zz_10819 = _zz_10820[31 : 0];
  assign _zz_10820 = _zz_10821;
  assign _zz_10821 = ($signed(_zz_10822) >>> _zz_720);
  assign _zz_10822 = _zz_10823;
  assign _zz_10823 = ($signed(_zz_10825) + $signed(_zz_716));
  assign _zz_10824 = ({8'd0,data_mid_27_real} <<< 8);
  assign _zz_10825 = {{8{_zz_10824[23]}}, _zz_10824};
  assign _zz_10826 = fixTo_862_dout;
  assign _zz_10827 = _zz_10828[31 : 0];
  assign _zz_10828 = _zz_10829;
  assign _zz_10829 = ($signed(_zz_10830) >>> _zz_720);
  assign _zz_10830 = _zz_10831;
  assign _zz_10831 = ($signed(_zz_10833) + $signed(_zz_717));
  assign _zz_10832 = ({8'd0,data_mid_27_imag} <<< 8);
  assign _zz_10833 = {{8{_zz_10832[23]}}, _zz_10832};
  assign _zz_10834 = fixTo_863_dout;
  assign _zz_10835 = ($signed(twiddle_factor_table_3_real) + $signed(twiddle_factor_table_3_imag));
  assign _zz_10836 = ($signed(_zz_723) - $signed(_zz_10837));
  assign _zz_10837 = ($signed(_zz_10838) * $signed(twiddle_factor_table_3_imag));
  assign _zz_10838 = ($signed(data_mid_36_real) + $signed(data_mid_36_imag));
  assign _zz_10839 = fixTo_864_dout;
  assign _zz_10840 = ($signed(_zz_723) + $signed(_zz_10841));
  assign _zz_10841 = ($signed(_zz_10842) * $signed(twiddle_factor_table_3_real));
  assign _zz_10842 = ($signed(data_mid_36_imag) - $signed(data_mid_36_real));
  assign _zz_10843 = fixTo_865_dout;
  assign _zz_10844 = _zz_10845[31 : 0];
  assign _zz_10845 = _zz_10846;
  assign _zz_10846 = ($signed(_zz_10847) >>> _zz_724);
  assign _zz_10847 = _zz_10848;
  assign _zz_10848 = ($signed(_zz_10850) - $signed(_zz_721));
  assign _zz_10849 = ({8'd0,data_mid_32_real} <<< 8);
  assign _zz_10850 = {{8{_zz_10849[23]}}, _zz_10849};
  assign _zz_10851 = fixTo_866_dout;
  assign _zz_10852 = _zz_10853[31 : 0];
  assign _zz_10853 = _zz_10854;
  assign _zz_10854 = ($signed(_zz_10855) >>> _zz_724);
  assign _zz_10855 = _zz_10856;
  assign _zz_10856 = ($signed(_zz_10858) - $signed(_zz_722));
  assign _zz_10857 = ({8'd0,data_mid_32_imag} <<< 8);
  assign _zz_10858 = {{8{_zz_10857[23]}}, _zz_10857};
  assign _zz_10859 = fixTo_867_dout;
  assign _zz_10860 = _zz_10861[31 : 0];
  assign _zz_10861 = _zz_10862;
  assign _zz_10862 = ($signed(_zz_10863) >>> _zz_725);
  assign _zz_10863 = _zz_10864;
  assign _zz_10864 = ($signed(_zz_10866) + $signed(_zz_721));
  assign _zz_10865 = ({8'd0,data_mid_32_real} <<< 8);
  assign _zz_10866 = {{8{_zz_10865[23]}}, _zz_10865};
  assign _zz_10867 = fixTo_868_dout;
  assign _zz_10868 = _zz_10869[31 : 0];
  assign _zz_10869 = _zz_10870;
  assign _zz_10870 = ($signed(_zz_10871) >>> _zz_725);
  assign _zz_10871 = _zz_10872;
  assign _zz_10872 = ($signed(_zz_10874) + $signed(_zz_722));
  assign _zz_10873 = ({8'd0,data_mid_32_imag} <<< 8);
  assign _zz_10874 = {{8{_zz_10873[23]}}, _zz_10873};
  assign _zz_10875 = fixTo_869_dout;
  assign _zz_10876 = ($signed(twiddle_factor_table_4_real) + $signed(twiddle_factor_table_4_imag));
  assign _zz_10877 = ($signed(_zz_728) - $signed(_zz_10878));
  assign _zz_10878 = ($signed(_zz_10879) * $signed(twiddle_factor_table_4_imag));
  assign _zz_10879 = ($signed(data_mid_37_real) + $signed(data_mid_37_imag));
  assign _zz_10880 = fixTo_870_dout;
  assign _zz_10881 = ($signed(_zz_728) + $signed(_zz_10882));
  assign _zz_10882 = ($signed(_zz_10883) * $signed(twiddle_factor_table_4_real));
  assign _zz_10883 = ($signed(data_mid_37_imag) - $signed(data_mid_37_real));
  assign _zz_10884 = fixTo_871_dout;
  assign _zz_10885 = _zz_10886[31 : 0];
  assign _zz_10886 = _zz_10887;
  assign _zz_10887 = ($signed(_zz_10888) >>> _zz_729);
  assign _zz_10888 = _zz_10889;
  assign _zz_10889 = ($signed(_zz_10891) - $signed(_zz_726));
  assign _zz_10890 = ({8'd0,data_mid_33_real} <<< 8);
  assign _zz_10891 = {{8{_zz_10890[23]}}, _zz_10890};
  assign _zz_10892 = fixTo_872_dout;
  assign _zz_10893 = _zz_10894[31 : 0];
  assign _zz_10894 = _zz_10895;
  assign _zz_10895 = ($signed(_zz_10896) >>> _zz_729);
  assign _zz_10896 = _zz_10897;
  assign _zz_10897 = ($signed(_zz_10899) - $signed(_zz_727));
  assign _zz_10898 = ({8'd0,data_mid_33_imag} <<< 8);
  assign _zz_10899 = {{8{_zz_10898[23]}}, _zz_10898};
  assign _zz_10900 = fixTo_873_dout;
  assign _zz_10901 = _zz_10902[31 : 0];
  assign _zz_10902 = _zz_10903;
  assign _zz_10903 = ($signed(_zz_10904) >>> _zz_730);
  assign _zz_10904 = _zz_10905;
  assign _zz_10905 = ($signed(_zz_10907) + $signed(_zz_726));
  assign _zz_10906 = ({8'd0,data_mid_33_real} <<< 8);
  assign _zz_10907 = {{8{_zz_10906[23]}}, _zz_10906};
  assign _zz_10908 = fixTo_874_dout;
  assign _zz_10909 = _zz_10910[31 : 0];
  assign _zz_10910 = _zz_10911;
  assign _zz_10911 = ($signed(_zz_10912) >>> _zz_730);
  assign _zz_10912 = _zz_10913;
  assign _zz_10913 = ($signed(_zz_10915) + $signed(_zz_727));
  assign _zz_10914 = ({8'd0,data_mid_33_imag} <<< 8);
  assign _zz_10915 = {{8{_zz_10914[23]}}, _zz_10914};
  assign _zz_10916 = fixTo_875_dout;
  assign _zz_10917 = ($signed(twiddle_factor_table_5_real) + $signed(twiddle_factor_table_5_imag));
  assign _zz_10918 = ($signed(_zz_733) - $signed(_zz_10919));
  assign _zz_10919 = ($signed(_zz_10920) * $signed(twiddle_factor_table_5_imag));
  assign _zz_10920 = ($signed(data_mid_38_real) + $signed(data_mid_38_imag));
  assign _zz_10921 = fixTo_876_dout;
  assign _zz_10922 = ($signed(_zz_733) + $signed(_zz_10923));
  assign _zz_10923 = ($signed(_zz_10924) * $signed(twiddle_factor_table_5_real));
  assign _zz_10924 = ($signed(data_mid_38_imag) - $signed(data_mid_38_real));
  assign _zz_10925 = fixTo_877_dout;
  assign _zz_10926 = _zz_10927[31 : 0];
  assign _zz_10927 = _zz_10928;
  assign _zz_10928 = ($signed(_zz_10929) >>> _zz_734);
  assign _zz_10929 = _zz_10930;
  assign _zz_10930 = ($signed(_zz_10932) - $signed(_zz_731));
  assign _zz_10931 = ({8'd0,data_mid_34_real} <<< 8);
  assign _zz_10932 = {{8{_zz_10931[23]}}, _zz_10931};
  assign _zz_10933 = fixTo_878_dout;
  assign _zz_10934 = _zz_10935[31 : 0];
  assign _zz_10935 = _zz_10936;
  assign _zz_10936 = ($signed(_zz_10937) >>> _zz_734);
  assign _zz_10937 = _zz_10938;
  assign _zz_10938 = ($signed(_zz_10940) - $signed(_zz_732));
  assign _zz_10939 = ({8'd0,data_mid_34_imag} <<< 8);
  assign _zz_10940 = {{8{_zz_10939[23]}}, _zz_10939};
  assign _zz_10941 = fixTo_879_dout;
  assign _zz_10942 = _zz_10943[31 : 0];
  assign _zz_10943 = _zz_10944;
  assign _zz_10944 = ($signed(_zz_10945) >>> _zz_735);
  assign _zz_10945 = _zz_10946;
  assign _zz_10946 = ($signed(_zz_10948) + $signed(_zz_731));
  assign _zz_10947 = ({8'd0,data_mid_34_real} <<< 8);
  assign _zz_10948 = {{8{_zz_10947[23]}}, _zz_10947};
  assign _zz_10949 = fixTo_880_dout;
  assign _zz_10950 = _zz_10951[31 : 0];
  assign _zz_10951 = _zz_10952;
  assign _zz_10952 = ($signed(_zz_10953) >>> _zz_735);
  assign _zz_10953 = _zz_10954;
  assign _zz_10954 = ($signed(_zz_10956) + $signed(_zz_732));
  assign _zz_10955 = ({8'd0,data_mid_34_imag} <<< 8);
  assign _zz_10956 = {{8{_zz_10955[23]}}, _zz_10955};
  assign _zz_10957 = fixTo_881_dout;
  assign _zz_10958 = ($signed(twiddle_factor_table_6_real) + $signed(twiddle_factor_table_6_imag));
  assign _zz_10959 = ($signed(_zz_738) - $signed(_zz_10960));
  assign _zz_10960 = ($signed(_zz_10961) * $signed(twiddle_factor_table_6_imag));
  assign _zz_10961 = ($signed(data_mid_39_real) + $signed(data_mid_39_imag));
  assign _zz_10962 = fixTo_882_dout;
  assign _zz_10963 = ($signed(_zz_738) + $signed(_zz_10964));
  assign _zz_10964 = ($signed(_zz_10965) * $signed(twiddle_factor_table_6_real));
  assign _zz_10965 = ($signed(data_mid_39_imag) - $signed(data_mid_39_real));
  assign _zz_10966 = fixTo_883_dout;
  assign _zz_10967 = _zz_10968[31 : 0];
  assign _zz_10968 = _zz_10969;
  assign _zz_10969 = ($signed(_zz_10970) >>> _zz_739);
  assign _zz_10970 = _zz_10971;
  assign _zz_10971 = ($signed(_zz_10973) - $signed(_zz_736));
  assign _zz_10972 = ({8'd0,data_mid_35_real} <<< 8);
  assign _zz_10973 = {{8{_zz_10972[23]}}, _zz_10972};
  assign _zz_10974 = fixTo_884_dout;
  assign _zz_10975 = _zz_10976[31 : 0];
  assign _zz_10976 = _zz_10977;
  assign _zz_10977 = ($signed(_zz_10978) >>> _zz_739);
  assign _zz_10978 = _zz_10979;
  assign _zz_10979 = ($signed(_zz_10981) - $signed(_zz_737));
  assign _zz_10980 = ({8'd0,data_mid_35_imag} <<< 8);
  assign _zz_10981 = {{8{_zz_10980[23]}}, _zz_10980};
  assign _zz_10982 = fixTo_885_dout;
  assign _zz_10983 = _zz_10984[31 : 0];
  assign _zz_10984 = _zz_10985;
  assign _zz_10985 = ($signed(_zz_10986) >>> _zz_740);
  assign _zz_10986 = _zz_10987;
  assign _zz_10987 = ($signed(_zz_10989) + $signed(_zz_736));
  assign _zz_10988 = ({8'd0,data_mid_35_real} <<< 8);
  assign _zz_10989 = {{8{_zz_10988[23]}}, _zz_10988};
  assign _zz_10990 = fixTo_886_dout;
  assign _zz_10991 = _zz_10992[31 : 0];
  assign _zz_10992 = _zz_10993;
  assign _zz_10993 = ($signed(_zz_10994) >>> _zz_740);
  assign _zz_10994 = _zz_10995;
  assign _zz_10995 = ($signed(_zz_10997) + $signed(_zz_737));
  assign _zz_10996 = ({8'd0,data_mid_35_imag} <<< 8);
  assign _zz_10997 = {{8{_zz_10996[23]}}, _zz_10996};
  assign _zz_10998 = fixTo_887_dout;
  assign _zz_10999 = ($signed(twiddle_factor_table_3_real) + $signed(twiddle_factor_table_3_imag));
  assign _zz_11000 = ($signed(_zz_743) - $signed(_zz_11001));
  assign _zz_11001 = ($signed(_zz_11002) * $signed(twiddle_factor_table_3_imag));
  assign _zz_11002 = ($signed(data_mid_44_real) + $signed(data_mid_44_imag));
  assign _zz_11003 = fixTo_888_dout;
  assign _zz_11004 = ($signed(_zz_743) + $signed(_zz_11005));
  assign _zz_11005 = ($signed(_zz_11006) * $signed(twiddle_factor_table_3_real));
  assign _zz_11006 = ($signed(data_mid_44_imag) - $signed(data_mid_44_real));
  assign _zz_11007 = fixTo_889_dout;
  assign _zz_11008 = _zz_11009[31 : 0];
  assign _zz_11009 = _zz_11010;
  assign _zz_11010 = ($signed(_zz_11011) >>> _zz_744);
  assign _zz_11011 = _zz_11012;
  assign _zz_11012 = ($signed(_zz_11014) - $signed(_zz_741));
  assign _zz_11013 = ({8'd0,data_mid_40_real} <<< 8);
  assign _zz_11014 = {{8{_zz_11013[23]}}, _zz_11013};
  assign _zz_11015 = fixTo_890_dout;
  assign _zz_11016 = _zz_11017[31 : 0];
  assign _zz_11017 = _zz_11018;
  assign _zz_11018 = ($signed(_zz_11019) >>> _zz_744);
  assign _zz_11019 = _zz_11020;
  assign _zz_11020 = ($signed(_zz_11022) - $signed(_zz_742));
  assign _zz_11021 = ({8'd0,data_mid_40_imag} <<< 8);
  assign _zz_11022 = {{8{_zz_11021[23]}}, _zz_11021};
  assign _zz_11023 = fixTo_891_dout;
  assign _zz_11024 = _zz_11025[31 : 0];
  assign _zz_11025 = _zz_11026;
  assign _zz_11026 = ($signed(_zz_11027) >>> _zz_745);
  assign _zz_11027 = _zz_11028;
  assign _zz_11028 = ($signed(_zz_11030) + $signed(_zz_741));
  assign _zz_11029 = ({8'd0,data_mid_40_real} <<< 8);
  assign _zz_11030 = {{8{_zz_11029[23]}}, _zz_11029};
  assign _zz_11031 = fixTo_892_dout;
  assign _zz_11032 = _zz_11033[31 : 0];
  assign _zz_11033 = _zz_11034;
  assign _zz_11034 = ($signed(_zz_11035) >>> _zz_745);
  assign _zz_11035 = _zz_11036;
  assign _zz_11036 = ($signed(_zz_11038) + $signed(_zz_742));
  assign _zz_11037 = ({8'd0,data_mid_40_imag} <<< 8);
  assign _zz_11038 = {{8{_zz_11037[23]}}, _zz_11037};
  assign _zz_11039 = fixTo_893_dout;
  assign _zz_11040 = ($signed(twiddle_factor_table_4_real) + $signed(twiddle_factor_table_4_imag));
  assign _zz_11041 = ($signed(_zz_748) - $signed(_zz_11042));
  assign _zz_11042 = ($signed(_zz_11043) * $signed(twiddle_factor_table_4_imag));
  assign _zz_11043 = ($signed(data_mid_45_real) + $signed(data_mid_45_imag));
  assign _zz_11044 = fixTo_894_dout;
  assign _zz_11045 = ($signed(_zz_748) + $signed(_zz_11046));
  assign _zz_11046 = ($signed(_zz_11047) * $signed(twiddle_factor_table_4_real));
  assign _zz_11047 = ($signed(data_mid_45_imag) - $signed(data_mid_45_real));
  assign _zz_11048 = fixTo_895_dout;
  assign _zz_11049 = _zz_11050[31 : 0];
  assign _zz_11050 = _zz_11051;
  assign _zz_11051 = ($signed(_zz_11052) >>> _zz_749);
  assign _zz_11052 = _zz_11053;
  assign _zz_11053 = ($signed(_zz_11055) - $signed(_zz_746));
  assign _zz_11054 = ({8'd0,data_mid_41_real} <<< 8);
  assign _zz_11055 = {{8{_zz_11054[23]}}, _zz_11054};
  assign _zz_11056 = fixTo_896_dout;
  assign _zz_11057 = _zz_11058[31 : 0];
  assign _zz_11058 = _zz_11059;
  assign _zz_11059 = ($signed(_zz_11060) >>> _zz_749);
  assign _zz_11060 = _zz_11061;
  assign _zz_11061 = ($signed(_zz_11063) - $signed(_zz_747));
  assign _zz_11062 = ({8'd0,data_mid_41_imag} <<< 8);
  assign _zz_11063 = {{8{_zz_11062[23]}}, _zz_11062};
  assign _zz_11064 = fixTo_897_dout;
  assign _zz_11065 = _zz_11066[31 : 0];
  assign _zz_11066 = _zz_11067;
  assign _zz_11067 = ($signed(_zz_11068) >>> _zz_750);
  assign _zz_11068 = _zz_11069;
  assign _zz_11069 = ($signed(_zz_11071) + $signed(_zz_746));
  assign _zz_11070 = ({8'd0,data_mid_41_real} <<< 8);
  assign _zz_11071 = {{8{_zz_11070[23]}}, _zz_11070};
  assign _zz_11072 = fixTo_898_dout;
  assign _zz_11073 = _zz_11074[31 : 0];
  assign _zz_11074 = _zz_11075;
  assign _zz_11075 = ($signed(_zz_11076) >>> _zz_750);
  assign _zz_11076 = _zz_11077;
  assign _zz_11077 = ($signed(_zz_11079) + $signed(_zz_747));
  assign _zz_11078 = ({8'd0,data_mid_41_imag} <<< 8);
  assign _zz_11079 = {{8{_zz_11078[23]}}, _zz_11078};
  assign _zz_11080 = fixTo_899_dout;
  assign _zz_11081 = ($signed(twiddle_factor_table_5_real) + $signed(twiddle_factor_table_5_imag));
  assign _zz_11082 = ($signed(_zz_753) - $signed(_zz_11083));
  assign _zz_11083 = ($signed(_zz_11084) * $signed(twiddle_factor_table_5_imag));
  assign _zz_11084 = ($signed(data_mid_46_real) + $signed(data_mid_46_imag));
  assign _zz_11085 = fixTo_900_dout;
  assign _zz_11086 = ($signed(_zz_753) + $signed(_zz_11087));
  assign _zz_11087 = ($signed(_zz_11088) * $signed(twiddle_factor_table_5_real));
  assign _zz_11088 = ($signed(data_mid_46_imag) - $signed(data_mid_46_real));
  assign _zz_11089 = fixTo_901_dout;
  assign _zz_11090 = _zz_11091[31 : 0];
  assign _zz_11091 = _zz_11092;
  assign _zz_11092 = ($signed(_zz_11093) >>> _zz_754);
  assign _zz_11093 = _zz_11094;
  assign _zz_11094 = ($signed(_zz_11096) - $signed(_zz_751));
  assign _zz_11095 = ({8'd0,data_mid_42_real} <<< 8);
  assign _zz_11096 = {{8{_zz_11095[23]}}, _zz_11095};
  assign _zz_11097 = fixTo_902_dout;
  assign _zz_11098 = _zz_11099[31 : 0];
  assign _zz_11099 = _zz_11100;
  assign _zz_11100 = ($signed(_zz_11101) >>> _zz_754);
  assign _zz_11101 = _zz_11102;
  assign _zz_11102 = ($signed(_zz_11104) - $signed(_zz_752));
  assign _zz_11103 = ({8'd0,data_mid_42_imag} <<< 8);
  assign _zz_11104 = {{8{_zz_11103[23]}}, _zz_11103};
  assign _zz_11105 = fixTo_903_dout;
  assign _zz_11106 = _zz_11107[31 : 0];
  assign _zz_11107 = _zz_11108;
  assign _zz_11108 = ($signed(_zz_11109) >>> _zz_755);
  assign _zz_11109 = _zz_11110;
  assign _zz_11110 = ($signed(_zz_11112) + $signed(_zz_751));
  assign _zz_11111 = ({8'd0,data_mid_42_real} <<< 8);
  assign _zz_11112 = {{8{_zz_11111[23]}}, _zz_11111};
  assign _zz_11113 = fixTo_904_dout;
  assign _zz_11114 = _zz_11115[31 : 0];
  assign _zz_11115 = _zz_11116;
  assign _zz_11116 = ($signed(_zz_11117) >>> _zz_755);
  assign _zz_11117 = _zz_11118;
  assign _zz_11118 = ($signed(_zz_11120) + $signed(_zz_752));
  assign _zz_11119 = ({8'd0,data_mid_42_imag} <<< 8);
  assign _zz_11120 = {{8{_zz_11119[23]}}, _zz_11119};
  assign _zz_11121 = fixTo_905_dout;
  assign _zz_11122 = ($signed(twiddle_factor_table_6_real) + $signed(twiddle_factor_table_6_imag));
  assign _zz_11123 = ($signed(_zz_758) - $signed(_zz_11124));
  assign _zz_11124 = ($signed(_zz_11125) * $signed(twiddle_factor_table_6_imag));
  assign _zz_11125 = ($signed(data_mid_47_real) + $signed(data_mid_47_imag));
  assign _zz_11126 = fixTo_906_dout;
  assign _zz_11127 = ($signed(_zz_758) + $signed(_zz_11128));
  assign _zz_11128 = ($signed(_zz_11129) * $signed(twiddle_factor_table_6_real));
  assign _zz_11129 = ($signed(data_mid_47_imag) - $signed(data_mid_47_real));
  assign _zz_11130 = fixTo_907_dout;
  assign _zz_11131 = _zz_11132[31 : 0];
  assign _zz_11132 = _zz_11133;
  assign _zz_11133 = ($signed(_zz_11134) >>> _zz_759);
  assign _zz_11134 = _zz_11135;
  assign _zz_11135 = ($signed(_zz_11137) - $signed(_zz_756));
  assign _zz_11136 = ({8'd0,data_mid_43_real} <<< 8);
  assign _zz_11137 = {{8{_zz_11136[23]}}, _zz_11136};
  assign _zz_11138 = fixTo_908_dout;
  assign _zz_11139 = _zz_11140[31 : 0];
  assign _zz_11140 = _zz_11141;
  assign _zz_11141 = ($signed(_zz_11142) >>> _zz_759);
  assign _zz_11142 = _zz_11143;
  assign _zz_11143 = ($signed(_zz_11145) - $signed(_zz_757));
  assign _zz_11144 = ({8'd0,data_mid_43_imag} <<< 8);
  assign _zz_11145 = {{8{_zz_11144[23]}}, _zz_11144};
  assign _zz_11146 = fixTo_909_dout;
  assign _zz_11147 = _zz_11148[31 : 0];
  assign _zz_11148 = _zz_11149;
  assign _zz_11149 = ($signed(_zz_11150) >>> _zz_760);
  assign _zz_11150 = _zz_11151;
  assign _zz_11151 = ($signed(_zz_11153) + $signed(_zz_756));
  assign _zz_11152 = ({8'd0,data_mid_43_real} <<< 8);
  assign _zz_11153 = {{8{_zz_11152[23]}}, _zz_11152};
  assign _zz_11154 = fixTo_910_dout;
  assign _zz_11155 = _zz_11156[31 : 0];
  assign _zz_11156 = _zz_11157;
  assign _zz_11157 = ($signed(_zz_11158) >>> _zz_760);
  assign _zz_11158 = _zz_11159;
  assign _zz_11159 = ($signed(_zz_11161) + $signed(_zz_757));
  assign _zz_11160 = ({8'd0,data_mid_43_imag} <<< 8);
  assign _zz_11161 = {{8{_zz_11160[23]}}, _zz_11160};
  assign _zz_11162 = fixTo_911_dout;
  assign _zz_11163 = ($signed(twiddle_factor_table_3_real) + $signed(twiddle_factor_table_3_imag));
  assign _zz_11164 = ($signed(_zz_763) - $signed(_zz_11165));
  assign _zz_11165 = ($signed(_zz_11166) * $signed(twiddle_factor_table_3_imag));
  assign _zz_11166 = ($signed(data_mid_52_real) + $signed(data_mid_52_imag));
  assign _zz_11167 = fixTo_912_dout;
  assign _zz_11168 = ($signed(_zz_763) + $signed(_zz_11169));
  assign _zz_11169 = ($signed(_zz_11170) * $signed(twiddle_factor_table_3_real));
  assign _zz_11170 = ($signed(data_mid_52_imag) - $signed(data_mid_52_real));
  assign _zz_11171 = fixTo_913_dout;
  assign _zz_11172 = _zz_11173[31 : 0];
  assign _zz_11173 = _zz_11174;
  assign _zz_11174 = ($signed(_zz_11175) >>> _zz_764);
  assign _zz_11175 = _zz_11176;
  assign _zz_11176 = ($signed(_zz_11178) - $signed(_zz_761));
  assign _zz_11177 = ({8'd0,data_mid_48_real} <<< 8);
  assign _zz_11178 = {{8{_zz_11177[23]}}, _zz_11177};
  assign _zz_11179 = fixTo_914_dout;
  assign _zz_11180 = _zz_11181[31 : 0];
  assign _zz_11181 = _zz_11182;
  assign _zz_11182 = ($signed(_zz_11183) >>> _zz_764);
  assign _zz_11183 = _zz_11184;
  assign _zz_11184 = ($signed(_zz_11186) - $signed(_zz_762));
  assign _zz_11185 = ({8'd0,data_mid_48_imag} <<< 8);
  assign _zz_11186 = {{8{_zz_11185[23]}}, _zz_11185};
  assign _zz_11187 = fixTo_915_dout;
  assign _zz_11188 = _zz_11189[31 : 0];
  assign _zz_11189 = _zz_11190;
  assign _zz_11190 = ($signed(_zz_11191) >>> _zz_765);
  assign _zz_11191 = _zz_11192;
  assign _zz_11192 = ($signed(_zz_11194) + $signed(_zz_761));
  assign _zz_11193 = ({8'd0,data_mid_48_real} <<< 8);
  assign _zz_11194 = {{8{_zz_11193[23]}}, _zz_11193};
  assign _zz_11195 = fixTo_916_dout;
  assign _zz_11196 = _zz_11197[31 : 0];
  assign _zz_11197 = _zz_11198;
  assign _zz_11198 = ($signed(_zz_11199) >>> _zz_765);
  assign _zz_11199 = _zz_11200;
  assign _zz_11200 = ($signed(_zz_11202) + $signed(_zz_762));
  assign _zz_11201 = ({8'd0,data_mid_48_imag} <<< 8);
  assign _zz_11202 = {{8{_zz_11201[23]}}, _zz_11201};
  assign _zz_11203 = fixTo_917_dout;
  assign _zz_11204 = ($signed(twiddle_factor_table_4_real) + $signed(twiddle_factor_table_4_imag));
  assign _zz_11205 = ($signed(_zz_768) - $signed(_zz_11206));
  assign _zz_11206 = ($signed(_zz_11207) * $signed(twiddle_factor_table_4_imag));
  assign _zz_11207 = ($signed(data_mid_53_real) + $signed(data_mid_53_imag));
  assign _zz_11208 = fixTo_918_dout;
  assign _zz_11209 = ($signed(_zz_768) + $signed(_zz_11210));
  assign _zz_11210 = ($signed(_zz_11211) * $signed(twiddle_factor_table_4_real));
  assign _zz_11211 = ($signed(data_mid_53_imag) - $signed(data_mid_53_real));
  assign _zz_11212 = fixTo_919_dout;
  assign _zz_11213 = _zz_11214[31 : 0];
  assign _zz_11214 = _zz_11215;
  assign _zz_11215 = ($signed(_zz_11216) >>> _zz_769);
  assign _zz_11216 = _zz_11217;
  assign _zz_11217 = ($signed(_zz_11219) - $signed(_zz_766));
  assign _zz_11218 = ({8'd0,data_mid_49_real} <<< 8);
  assign _zz_11219 = {{8{_zz_11218[23]}}, _zz_11218};
  assign _zz_11220 = fixTo_920_dout;
  assign _zz_11221 = _zz_11222[31 : 0];
  assign _zz_11222 = _zz_11223;
  assign _zz_11223 = ($signed(_zz_11224) >>> _zz_769);
  assign _zz_11224 = _zz_11225;
  assign _zz_11225 = ($signed(_zz_11227) - $signed(_zz_767));
  assign _zz_11226 = ({8'd0,data_mid_49_imag} <<< 8);
  assign _zz_11227 = {{8{_zz_11226[23]}}, _zz_11226};
  assign _zz_11228 = fixTo_921_dout;
  assign _zz_11229 = _zz_11230[31 : 0];
  assign _zz_11230 = _zz_11231;
  assign _zz_11231 = ($signed(_zz_11232) >>> _zz_770);
  assign _zz_11232 = _zz_11233;
  assign _zz_11233 = ($signed(_zz_11235) + $signed(_zz_766));
  assign _zz_11234 = ({8'd0,data_mid_49_real} <<< 8);
  assign _zz_11235 = {{8{_zz_11234[23]}}, _zz_11234};
  assign _zz_11236 = fixTo_922_dout;
  assign _zz_11237 = _zz_11238[31 : 0];
  assign _zz_11238 = _zz_11239;
  assign _zz_11239 = ($signed(_zz_11240) >>> _zz_770);
  assign _zz_11240 = _zz_11241;
  assign _zz_11241 = ($signed(_zz_11243) + $signed(_zz_767));
  assign _zz_11242 = ({8'd0,data_mid_49_imag} <<< 8);
  assign _zz_11243 = {{8{_zz_11242[23]}}, _zz_11242};
  assign _zz_11244 = fixTo_923_dout;
  assign _zz_11245 = ($signed(twiddle_factor_table_5_real) + $signed(twiddle_factor_table_5_imag));
  assign _zz_11246 = ($signed(_zz_773) - $signed(_zz_11247));
  assign _zz_11247 = ($signed(_zz_11248) * $signed(twiddle_factor_table_5_imag));
  assign _zz_11248 = ($signed(data_mid_54_real) + $signed(data_mid_54_imag));
  assign _zz_11249 = fixTo_924_dout;
  assign _zz_11250 = ($signed(_zz_773) + $signed(_zz_11251));
  assign _zz_11251 = ($signed(_zz_11252) * $signed(twiddle_factor_table_5_real));
  assign _zz_11252 = ($signed(data_mid_54_imag) - $signed(data_mid_54_real));
  assign _zz_11253 = fixTo_925_dout;
  assign _zz_11254 = _zz_11255[31 : 0];
  assign _zz_11255 = _zz_11256;
  assign _zz_11256 = ($signed(_zz_11257) >>> _zz_774);
  assign _zz_11257 = _zz_11258;
  assign _zz_11258 = ($signed(_zz_11260) - $signed(_zz_771));
  assign _zz_11259 = ({8'd0,data_mid_50_real} <<< 8);
  assign _zz_11260 = {{8{_zz_11259[23]}}, _zz_11259};
  assign _zz_11261 = fixTo_926_dout;
  assign _zz_11262 = _zz_11263[31 : 0];
  assign _zz_11263 = _zz_11264;
  assign _zz_11264 = ($signed(_zz_11265) >>> _zz_774);
  assign _zz_11265 = _zz_11266;
  assign _zz_11266 = ($signed(_zz_11268) - $signed(_zz_772));
  assign _zz_11267 = ({8'd0,data_mid_50_imag} <<< 8);
  assign _zz_11268 = {{8{_zz_11267[23]}}, _zz_11267};
  assign _zz_11269 = fixTo_927_dout;
  assign _zz_11270 = _zz_11271[31 : 0];
  assign _zz_11271 = _zz_11272;
  assign _zz_11272 = ($signed(_zz_11273) >>> _zz_775);
  assign _zz_11273 = _zz_11274;
  assign _zz_11274 = ($signed(_zz_11276) + $signed(_zz_771));
  assign _zz_11275 = ({8'd0,data_mid_50_real} <<< 8);
  assign _zz_11276 = {{8{_zz_11275[23]}}, _zz_11275};
  assign _zz_11277 = fixTo_928_dout;
  assign _zz_11278 = _zz_11279[31 : 0];
  assign _zz_11279 = _zz_11280;
  assign _zz_11280 = ($signed(_zz_11281) >>> _zz_775);
  assign _zz_11281 = _zz_11282;
  assign _zz_11282 = ($signed(_zz_11284) + $signed(_zz_772));
  assign _zz_11283 = ({8'd0,data_mid_50_imag} <<< 8);
  assign _zz_11284 = {{8{_zz_11283[23]}}, _zz_11283};
  assign _zz_11285 = fixTo_929_dout;
  assign _zz_11286 = ($signed(twiddle_factor_table_6_real) + $signed(twiddle_factor_table_6_imag));
  assign _zz_11287 = ($signed(_zz_778) - $signed(_zz_11288));
  assign _zz_11288 = ($signed(_zz_11289) * $signed(twiddle_factor_table_6_imag));
  assign _zz_11289 = ($signed(data_mid_55_real) + $signed(data_mid_55_imag));
  assign _zz_11290 = fixTo_930_dout;
  assign _zz_11291 = ($signed(_zz_778) + $signed(_zz_11292));
  assign _zz_11292 = ($signed(_zz_11293) * $signed(twiddle_factor_table_6_real));
  assign _zz_11293 = ($signed(data_mid_55_imag) - $signed(data_mid_55_real));
  assign _zz_11294 = fixTo_931_dout;
  assign _zz_11295 = _zz_11296[31 : 0];
  assign _zz_11296 = _zz_11297;
  assign _zz_11297 = ($signed(_zz_11298) >>> _zz_779);
  assign _zz_11298 = _zz_11299;
  assign _zz_11299 = ($signed(_zz_11301) - $signed(_zz_776));
  assign _zz_11300 = ({8'd0,data_mid_51_real} <<< 8);
  assign _zz_11301 = {{8{_zz_11300[23]}}, _zz_11300};
  assign _zz_11302 = fixTo_932_dout;
  assign _zz_11303 = _zz_11304[31 : 0];
  assign _zz_11304 = _zz_11305;
  assign _zz_11305 = ($signed(_zz_11306) >>> _zz_779);
  assign _zz_11306 = _zz_11307;
  assign _zz_11307 = ($signed(_zz_11309) - $signed(_zz_777));
  assign _zz_11308 = ({8'd0,data_mid_51_imag} <<< 8);
  assign _zz_11309 = {{8{_zz_11308[23]}}, _zz_11308};
  assign _zz_11310 = fixTo_933_dout;
  assign _zz_11311 = _zz_11312[31 : 0];
  assign _zz_11312 = _zz_11313;
  assign _zz_11313 = ($signed(_zz_11314) >>> _zz_780);
  assign _zz_11314 = _zz_11315;
  assign _zz_11315 = ($signed(_zz_11317) + $signed(_zz_776));
  assign _zz_11316 = ({8'd0,data_mid_51_real} <<< 8);
  assign _zz_11317 = {{8{_zz_11316[23]}}, _zz_11316};
  assign _zz_11318 = fixTo_934_dout;
  assign _zz_11319 = _zz_11320[31 : 0];
  assign _zz_11320 = _zz_11321;
  assign _zz_11321 = ($signed(_zz_11322) >>> _zz_780);
  assign _zz_11322 = _zz_11323;
  assign _zz_11323 = ($signed(_zz_11325) + $signed(_zz_777));
  assign _zz_11324 = ({8'd0,data_mid_51_imag} <<< 8);
  assign _zz_11325 = {{8{_zz_11324[23]}}, _zz_11324};
  assign _zz_11326 = fixTo_935_dout;
  assign _zz_11327 = ($signed(twiddle_factor_table_3_real) + $signed(twiddle_factor_table_3_imag));
  assign _zz_11328 = ($signed(_zz_783) - $signed(_zz_11329));
  assign _zz_11329 = ($signed(_zz_11330) * $signed(twiddle_factor_table_3_imag));
  assign _zz_11330 = ($signed(data_mid_60_real) + $signed(data_mid_60_imag));
  assign _zz_11331 = fixTo_936_dout;
  assign _zz_11332 = ($signed(_zz_783) + $signed(_zz_11333));
  assign _zz_11333 = ($signed(_zz_11334) * $signed(twiddle_factor_table_3_real));
  assign _zz_11334 = ($signed(data_mid_60_imag) - $signed(data_mid_60_real));
  assign _zz_11335 = fixTo_937_dout;
  assign _zz_11336 = _zz_11337[31 : 0];
  assign _zz_11337 = _zz_11338;
  assign _zz_11338 = ($signed(_zz_11339) >>> _zz_784);
  assign _zz_11339 = _zz_11340;
  assign _zz_11340 = ($signed(_zz_11342) - $signed(_zz_781));
  assign _zz_11341 = ({8'd0,data_mid_56_real} <<< 8);
  assign _zz_11342 = {{8{_zz_11341[23]}}, _zz_11341};
  assign _zz_11343 = fixTo_938_dout;
  assign _zz_11344 = _zz_11345[31 : 0];
  assign _zz_11345 = _zz_11346;
  assign _zz_11346 = ($signed(_zz_11347) >>> _zz_784);
  assign _zz_11347 = _zz_11348;
  assign _zz_11348 = ($signed(_zz_11350) - $signed(_zz_782));
  assign _zz_11349 = ({8'd0,data_mid_56_imag} <<< 8);
  assign _zz_11350 = {{8{_zz_11349[23]}}, _zz_11349};
  assign _zz_11351 = fixTo_939_dout;
  assign _zz_11352 = _zz_11353[31 : 0];
  assign _zz_11353 = _zz_11354;
  assign _zz_11354 = ($signed(_zz_11355) >>> _zz_785);
  assign _zz_11355 = _zz_11356;
  assign _zz_11356 = ($signed(_zz_11358) + $signed(_zz_781));
  assign _zz_11357 = ({8'd0,data_mid_56_real} <<< 8);
  assign _zz_11358 = {{8{_zz_11357[23]}}, _zz_11357};
  assign _zz_11359 = fixTo_940_dout;
  assign _zz_11360 = _zz_11361[31 : 0];
  assign _zz_11361 = _zz_11362;
  assign _zz_11362 = ($signed(_zz_11363) >>> _zz_785);
  assign _zz_11363 = _zz_11364;
  assign _zz_11364 = ($signed(_zz_11366) + $signed(_zz_782));
  assign _zz_11365 = ({8'd0,data_mid_56_imag} <<< 8);
  assign _zz_11366 = {{8{_zz_11365[23]}}, _zz_11365};
  assign _zz_11367 = fixTo_941_dout;
  assign _zz_11368 = ($signed(twiddle_factor_table_4_real) + $signed(twiddle_factor_table_4_imag));
  assign _zz_11369 = ($signed(_zz_788) - $signed(_zz_11370));
  assign _zz_11370 = ($signed(_zz_11371) * $signed(twiddle_factor_table_4_imag));
  assign _zz_11371 = ($signed(data_mid_61_real) + $signed(data_mid_61_imag));
  assign _zz_11372 = fixTo_942_dout;
  assign _zz_11373 = ($signed(_zz_788) + $signed(_zz_11374));
  assign _zz_11374 = ($signed(_zz_11375) * $signed(twiddle_factor_table_4_real));
  assign _zz_11375 = ($signed(data_mid_61_imag) - $signed(data_mid_61_real));
  assign _zz_11376 = fixTo_943_dout;
  assign _zz_11377 = _zz_11378[31 : 0];
  assign _zz_11378 = _zz_11379;
  assign _zz_11379 = ($signed(_zz_11380) >>> _zz_789);
  assign _zz_11380 = _zz_11381;
  assign _zz_11381 = ($signed(_zz_11383) - $signed(_zz_786));
  assign _zz_11382 = ({8'd0,data_mid_57_real} <<< 8);
  assign _zz_11383 = {{8{_zz_11382[23]}}, _zz_11382};
  assign _zz_11384 = fixTo_944_dout;
  assign _zz_11385 = _zz_11386[31 : 0];
  assign _zz_11386 = _zz_11387;
  assign _zz_11387 = ($signed(_zz_11388) >>> _zz_789);
  assign _zz_11388 = _zz_11389;
  assign _zz_11389 = ($signed(_zz_11391) - $signed(_zz_787));
  assign _zz_11390 = ({8'd0,data_mid_57_imag} <<< 8);
  assign _zz_11391 = {{8{_zz_11390[23]}}, _zz_11390};
  assign _zz_11392 = fixTo_945_dout;
  assign _zz_11393 = _zz_11394[31 : 0];
  assign _zz_11394 = _zz_11395;
  assign _zz_11395 = ($signed(_zz_11396) >>> _zz_790);
  assign _zz_11396 = _zz_11397;
  assign _zz_11397 = ($signed(_zz_11399) + $signed(_zz_786));
  assign _zz_11398 = ({8'd0,data_mid_57_real} <<< 8);
  assign _zz_11399 = {{8{_zz_11398[23]}}, _zz_11398};
  assign _zz_11400 = fixTo_946_dout;
  assign _zz_11401 = _zz_11402[31 : 0];
  assign _zz_11402 = _zz_11403;
  assign _zz_11403 = ($signed(_zz_11404) >>> _zz_790);
  assign _zz_11404 = _zz_11405;
  assign _zz_11405 = ($signed(_zz_11407) + $signed(_zz_787));
  assign _zz_11406 = ({8'd0,data_mid_57_imag} <<< 8);
  assign _zz_11407 = {{8{_zz_11406[23]}}, _zz_11406};
  assign _zz_11408 = fixTo_947_dout;
  assign _zz_11409 = ($signed(twiddle_factor_table_5_real) + $signed(twiddle_factor_table_5_imag));
  assign _zz_11410 = ($signed(_zz_793) - $signed(_zz_11411));
  assign _zz_11411 = ($signed(_zz_11412) * $signed(twiddle_factor_table_5_imag));
  assign _zz_11412 = ($signed(data_mid_62_real) + $signed(data_mid_62_imag));
  assign _zz_11413 = fixTo_948_dout;
  assign _zz_11414 = ($signed(_zz_793) + $signed(_zz_11415));
  assign _zz_11415 = ($signed(_zz_11416) * $signed(twiddle_factor_table_5_real));
  assign _zz_11416 = ($signed(data_mid_62_imag) - $signed(data_mid_62_real));
  assign _zz_11417 = fixTo_949_dout;
  assign _zz_11418 = _zz_11419[31 : 0];
  assign _zz_11419 = _zz_11420;
  assign _zz_11420 = ($signed(_zz_11421) >>> _zz_794);
  assign _zz_11421 = _zz_11422;
  assign _zz_11422 = ($signed(_zz_11424) - $signed(_zz_791));
  assign _zz_11423 = ({8'd0,data_mid_58_real} <<< 8);
  assign _zz_11424 = {{8{_zz_11423[23]}}, _zz_11423};
  assign _zz_11425 = fixTo_950_dout;
  assign _zz_11426 = _zz_11427[31 : 0];
  assign _zz_11427 = _zz_11428;
  assign _zz_11428 = ($signed(_zz_11429) >>> _zz_794);
  assign _zz_11429 = _zz_11430;
  assign _zz_11430 = ($signed(_zz_11432) - $signed(_zz_792));
  assign _zz_11431 = ({8'd0,data_mid_58_imag} <<< 8);
  assign _zz_11432 = {{8{_zz_11431[23]}}, _zz_11431};
  assign _zz_11433 = fixTo_951_dout;
  assign _zz_11434 = _zz_11435[31 : 0];
  assign _zz_11435 = _zz_11436;
  assign _zz_11436 = ($signed(_zz_11437) >>> _zz_795);
  assign _zz_11437 = _zz_11438;
  assign _zz_11438 = ($signed(_zz_11440) + $signed(_zz_791));
  assign _zz_11439 = ({8'd0,data_mid_58_real} <<< 8);
  assign _zz_11440 = {{8{_zz_11439[23]}}, _zz_11439};
  assign _zz_11441 = fixTo_952_dout;
  assign _zz_11442 = _zz_11443[31 : 0];
  assign _zz_11443 = _zz_11444;
  assign _zz_11444 = ($signed(_zz_11445) >>> _zz_795);
  assign _zz_11445 = _zz_11446;
  assign _zz_11446 = ($signed(_zz_11448) + $signed(_zz_792));
  assign _zz_11447 = ({8'd0,data_mid_58_imag} <<< 8);
  assign _zz_11448 = {{8{_zz_11447[23]}}, _zz_11447};
  assign _zz_11449 = fixTo_953_dout;
  assign _zz_11450 = ($signed(twiddle_factor_table_6_real) + $signed(twiddle_factor_table_6_imag));
  assign _zz_11451 = ($signed(_zz_798) - $signed(_zz_11452));
  assign _zz_11452 = ($signed(_zz_11453) * $signed(twiddle_factor_table_6_imag));
  assign _zz_11453 = ($signed(data_mid_63_real) + $signed(data_mid_63_imag));
  assign _zz_11454 = fixTo_954_dout;
  assign _zz_11455 = ($signed(_zz_798) + $signed(_zz_11456));
  assign _zz_11456 = ($signed(_zz_11457) * $signed(twiddle_factor_table_6_real));
  assign _zz_11457 = ($signed(data_mid_63_imag) - $signed(data_mid_63_real));
  assign _zz_11458 = fixTo_955_dout;
  assign _zz_11459 = _zz_11460[31 : 0];
  assign _zz_11460 = _zz_11461;
  assign _zz_11461 = ($signed(_zz_11462) >>> _zz_799);
  assign _zz_11462 = _zz_11463;
  assign _zz_11463 = ($signed(_zz_11465) - $signed(_zz_796));
  assign _zz_11464 = ({8'd0,data_mid_59_real} <<< 8);
  assign _zz_11465 = {{8{_zz_11464[23]}}, _zz_11464};
  assign _zz_11466 = fixTo_956_dout;
  assign _zz_11467 = _zz_11468[31 : 0];
  assign _zz_11468 = _zz_11469;
  assign _zz_11469 = ($signed(_zz_11470) >>> _zz_799);
  assign _zz_11470 = _zz_11471;
  assign _zz_11471 = ($signed(_zz_11473) - $signed(_zz_797));
  assign _zz_11472 = ({8'd0,data_mid_59_imag} <<< 8);
  assign _zz_11473 = {{8{_zz_11472[23]}}, _zz_11472};
  assign _zz_11474 = fixTo_957_dout;
  assign _zz_11475 = _zz_11476[31 : 0];
  assign _zz_11476 = _zz_11477;
  assign _zz_11477 = ($signed(_zz_11478) >>> _zz_800);
  assign _zz_11478 = _zz_11479;
  assign _zz_11479 = ($signed(_zz_11481) + $signed(_zz_796));
  assign _zz_11480 = ({8'd0,data_mid_59_real} <<< 8);
  assign _zz_11481 = {{8{_zz_11480[23]}}, _zz_11480};
  assign _zz_11482 = fixTo_958_dout;
  assign _zz_11483 = _zz_11484[31 : 0];
  assign _zz_11484 = _zz_11485;
  assign _zz_11485 = ($signed(_zz_11486) >>> _zz_800);
  assign _zz_11486 = _zz_11487;
  assign _zz_11487 = ($signed(_zz_11489) + $signed(_zz_797));
  assign _zz_11488 = ({8'd0,data_mid_59_imag} <<< 8);
  assign _zz_11489 = {{8{_zz_11488[23]}}, _zz_11488};
  assign _zz_11490 = fixTo_959_dout;
  assign _zz_11491 = ($signed(twiddle_factor_table_3_real) + $signed(twiddle_factor_table_3_imag));
  assign _zz_11492 = ($signed(_zz_803) - $signed(_zz_11493));
  assign _zz_11493 = ($signed(_zz_11494) * $signed(twiddle_factor_table_3_imag));
  assign _zz_11494 = ($signed(data_mid_68_real) + $signed(data_mid_68_imag));
  assign _zz_11495 = fixTo_960_dout;
  assign _zz_11496 = ($signed(_zz_803) + $signed(_zz_11497));
  assign _zz_11497 = ($signed(_zz_11498) * $signed(twiddle_factor_table_3_real));
  assign _zz_11498 = ($signed(data_mid_68_imag) - $signed(data_mid_68_real));
  assign _zz_11499 = fixTo_961_dout;
  assign _zz_11500 = _zz_11501[31 : 0];
  assign _zz_11501 = _zz_11502;
  assign _zz_11502 = ($signed(_zz_11503) >>> _zz_804);
  assign _zz_11503 = _zz_11504;
  assign _zz_11504 = ($signed(_zz_11506) - $signed(_zz_801));
  assign _zz_11505 = ({8'd0,data_mid_64_real} <<< 8);
  assign _zz_11506 = {{8{_zz_11505[23]}}, _zz_11505};
  assign _zz_11507 = fixTo_962_dout;
  assign _zz_11508 = _zz_11509[31 : 0];
  assign _zz_11509 = _zz_11510;
  assign _zz_11510 = ($signed(_zz_11511) >>> _zz_804);
  assign _zz_11511 = _zz_11512;
  assign _zz_11512 = ($signed(_zz_11514) - $signed(_zz_802));
  assign _zz_11513 = ({8'd0,data_mid_64_imag} <<< 8);
  assign _zz_11514 = {{8{_zz_11513[23]}}, _zz_11513};
  assign _zz_11515 = fixTo_963_dout;
  assign _zz_11516 = _zz_11517[31 : 0];
  assign _zz_11517 = _zz_11518;
  assign _zz_11518 = ($signed(_zz_11519) >>> _zz_805);
  assign _zz_11519 = _zz_11520;
  assign _zz_11520 = ($signed(_zz_11522) + $signed(_zz_801));
  assign _zz_11521 = ({8'd0,data_mid_64_real} <<< 8);
  assign _zz_11522 = {{8{_zz_11521[23]}}, _zz_11521};
  assign _zz_11523 = fixTo_964_dout;
  assign _zz_11524 = _zz_11525[31 : 0];
  assign _zz_11525 = _zz_11526;
  assign _zz_11526 = ($signed(_zz_11527) >>> _zz_805);
  assign _zz_11527 = _zz_11528;
  assign _zz_11528 = ($signed(_zz_11530) + $signed(_zz_802));
  assign _zz_11529 = ({8'd0,data_mid_64_imag} <<< 8);
  assign _zz_11530 = {{8{_zz_11529[23]}}, _zz_11529};
  assign _zz_11531 = fixTo_965_dout;
  assign _zz_11532 = ($signed(twiddle_factor_table_4_real) + $signed(twiddle_factor_table_4_imag));
  assign _zz_11533 = ($signed(_zz_808) - $signed(_zz_11534));
  assign _zz_11534 = ($signed(_zz_11535) * $signed(twiddle_factor_table_4_imag));
  assign _zz_11535 = ($signed(data_mid_69_real) + $signed(data_mid_69_imag));
  assign _zz_11536 = fixTo_966_dout;
  assign _zz_11537 = ($signed(_zz_808) + $signed(_zz_11538));
  assign _zz_11538 = ($signed(_zz_11539) * $signed(twiddle_factor_table_4_real));
  assign _zz_11539 = ($signed(data_mid_69_imag) - $signed(data_mid_69_real));
  assign _zz_11540 = fixTo_967_dout;
  assign _zz_11541 = _zz_11542[31 : 0];
  assign _zz_11542 = _zz_11543;
  assign _zz_11543 = ($signed(_zz_11544) >>> _zz_809);
  assign _zz_11544 = _zz_11545;
  assign _zz_11545 = ($signed(_zz_11547) - $signed(_zz_806));
  assign _zz_11546 = ({8'd0,data_mid_65_real} <<< 8);
  assign _zz_11547 = {{8{_zz_11546[23]}}, _zz_11546};
  assign _zz_11548 = fixTo_968_dout;
  assign _zz_11549 = _zz_11550[31 : 0];
  assign _zz_11550 = _zz_11551;
  assign _zz_11551 = ($signed(_zz_11552) >>> _zz_809);
  assign _zz_11552 = _zz_11553;
  assign _zz_11553 = ($signed(_zz_11555) - $signed(_zz_807));
  assign _zz_11554 = ({8'd0,data_mid_65_imag} <<< 8);
  assign _zz_11555 = {{8{_zz_11554[23]}}, _zz_11554};
  assign _zz_11556 = fixTo_969_dout;
  assign _zz_11557 = _zz_11558[31 : 0];
  assign _zz_11558 = _zz_11559;
  assign _zz_11559 = ($signed(_zz_11560) >>> _zz_810);
  assign _zz_11560 = _zz_11561;
  assign _zz_11561 = ($signed(_zz_11563) + $signed(_zz_806));
  assign _zz_11562 = ({8'd0,data_mid_65_real} <<< 8);
  assign _zz_11563 = {{8{_zz_11562[23]}}, _zz_11562};
  assign _zz_11564 = fixTo_970_dout;
  assign _zz_11565 = _zz_11566[31 : 0];
  assign _zz_11566 = _zz_11567;
  assign _zz_11567 = ($signed(_zz_11568) >>> _zz_810);
  assign _zz_11568 = _zz_11569;
  assign _zz_11569 = ($signed(_zz_11571) + $signed(_zz_807));
  assign _zz_11570 = ({8'd0,data_mid_65_imag} <<< 8);
  assign _zz_11571 = {{8{_zz_11570[23]}}, _zz_11570};
  assign _zz_11572 = fixTo_971_dout;
  assign _zz_11573 = ($signed(twiddle_factor_table_5_real) + $signed(twiddle_factor_table_5_imag));
  assign _zz_11574 = ($signed(_zz_813) - $signed(_zz_11575));
  assign _zz_11575 = ($signed(_zz_11576) * $signed(twiddle_factor_table_5_imag));
  assign _zz_11576 = ($signed(data_mid_70_real) + $signed(data_mid_70_imag));
  assign _zz_11577 = fixTo_972_dout;
  assign _zz_11578 = ($signed(_zz_813) + $signed(_zz_11579));
  assign _zz_11579 = ($signed(_zz_11580) * $signed(twiddle_factor_table_5_real));
  assign _zz_11580 = ($signed(data_mid_70_imag) - $signed(data_mid_70_real));
  assign _zz_11581 = fixTo_973_dout;
  assign _zz_11582 = _zz_11583[31 : 0];
  assign _zz_11583 = _zz_11584;
  assign _zz_11584 = ($signed(_zz_11585) >>> _zz_814);
  assign _zz_11585 = _zz_11586;
  assign _zz_11586 = ($signed(_zz_11588) - $signed(_zz_811));
  assign _zz_11587 = ({8'd0,data_mid_66_real} <<< 8);
  assign _zz_11588 = {{8{_zz_11587[23]}}, _zz_11587};
  assign _zz_11589 = fixTo_974_dout;
  assign _zz_11590 = _zz_11591[31 : 0];
  assign _zz_11591 = _zz_11592;
  assign _zz_11592 = ($signed(_zz_11593) >>> _zz_814);
  assign _zz_11593 = _zz_11594;
  assign _zz_11594 = ($signed(_zz_11596) - $signed(_zz_812));
  assign _zz_11595 = ({8'd0,data_mid_66_imag} <<< 8);
  assign _zz_11596 = {{8{_zz_11595[23]}}, _zz_11595};
  assign _zz_11597 = fixTo_975_dout;
  assign _zz_11598 = _zz_11599[31 : 0];
  assign _zz_11599 = _zz_11600;
  assign _zz_11600 = ($signed(_zz_11601) >>> _zz_815);
  assign _zz_11601 = _zz_11602;
  assign _zz_11602 = ($signed(_zz_11604) + $signed(_zz_811));
  assign _zz_11603 = ({8'd0,data_mid_66_real} <<< 8);
  assign _zz_11604 = {{8{_zz_11603[23]}}, _zz_11603};
  assign _zz_11605 = fixTo_976_dout;
  assign _zz_11606 = _zz_11607[31 : 0];
  assign _zz_11607 = _zz_11608;
  assign _zz_11608 = ($signed(_zz_11609) >>> _zz_815);
  assign _zz_11609 = _zz_11610;
  assign _zz_11610 = ($signed(_zz_11612) + $signed(_zz_812));
  assign _zz_11611 = ({8'd0,data_mid_66_imag} <<< 8);
  assign _zz_11612 = {{8{_zz_11611[23]}}, _zz_11611};
  assign _zz_11613 = fixTo_977_dout;
  assign _zz_11614 = ($signed(twiddle_factor_table_6_real) + $signed(twiddle_factor_table_6_imag));
  assign _zz_11615 = ($signed(_zz_818) - $signed(_zz_11616));
  assign _zz_11616 = ($signed(_zz_11617) * $signed(twiddle_factor_table_6_imag));
  assign _zz_11617 = ($signed(data_mid_71_real) + $signed(data_mid_71_imag));
  assign _zz_11618 = fixTo_978_dout;
  assign _zz_11619 = ($signed(_zz_818) + $signed(_zz_11620));
  assign _zz_11620 = ($signed(_zz_11621) * $signed(twiddle_factor_table_6_real));
  assign _zz_11621 = ($signed(data_mid_71_imag) - $signed(data_mid_71_real));
  assign _zz_11622 = fixTo_979_dout;
  assign _zz_11623 = _zz_11624[31 : 0];
  assign _zz_11624 = _zz_11625;
  assign _zz_11625 = ($signed(_zz_11626) >>> _zz_819);
  assign _zz_11626 = _zz_11627;
  assign _zz_11627 = ($signed(_zz_11629) - $signed(_zz_816));
  assign _zz_11628 = ({8'd0,data_mid_67_real} <<< 8);
  assign _zz_11629 = {{8{_zz_11628[23]}}, _zz_11628};
  assign _zz_11630 = fixTo_980_dout;
  assign _zz_11631 = _zz_11632[31 : 0];
  assign _zz_11632 = _zz_11633;
  assign _zz_11633 = ($signed(_zz_11634) >>> _zz_819);
  assign _zz_11634 = _zz_11635;
  assign _zz_11635 = ($signed(_zz_11637) - $signed(_zz_817));
  assign _zz_11636 = ({8'd0,data_mid_67_imag} <<< 8);
  assign _zz_11637 = {{8{_zz_11636[23]}}, _zz_11636};
  assign _zz_11638 = fixTo_981_dout;
  assign _zz_11639 = _zz_11640[31 : 0];
  assign _zz_11640 = _zz_11641;
  assign _zz_11641 = ($signed(_zz_11642) >>> _zz_820);
  assign _zz_11642 = _zz_11643;
  assign _zz_11643 = ($signed(_zz_11645) + $signed(_zz_816));
  assign _zz_11644 = ({8'd0,data_mid_67_real} <<< 8);
  assign _zz_11645 = {{8{_zz_11644[23]}}, _zz_11644};
  assign _zz_11646 = fixTo_982_dout;
  assign _zz_11647 = _zz_11648[31 : 0];
  assign _zz_11648 = _zz_11649;
  assign _zz_11649 = ($signed(_zz_11650) >>> _zz_820);
  assign _zz_11650 = _zz_11651;
  assign _zz_11651 = ($signed(_zz_11653) + $signed(_zz_817));
  assign _zz_11652 = ({8'd0,data_mid_67_imag} <<< 8);
  assign _zz_11653 = {{8{_zz_11652[23]}}, _zz_11652};
  assign _zz_11654 = fixTo_983_dout;
  assign _zz_11655 = ($signed(twiddle_factor_table_3_real) + $signed(twiddle_factor_table_3_imag));
  assign _zz_11656 = ($signed(_zz_823) - $signed(_zz_11657));
  assign _zz_11657 = ($signed(_zz_11658) * $signed(twiddle_factor_table_3_imag));
  assign _zz_11658 = ($signed(data_mid_76_real) + $signed(data_mid_76_imag));
  assign _zz_11659 = fixTo_984_dout;
  assign _zz_11660 = ($signed(_zz_823) + $signed(_zz_11661));
  assign _zz_11661 = ($signed(_zz_11662) * $signed(twiddle_factor_table_3_real));
  assign _zz_11662 = ($signed(data_mid_76_imag) - $signed(data_mid_76_real));
  assign _zz_11663 = fixTo_985_dout;
  assign _zz_11664 = _zz_11665[31 : 0];
  assign _zz_11665 = _zz_11666;
  assign _zz_11666 = ($signed(_zz_11667) >>> _zz_824);
  assign _zz_11667 = _zz_11668;
  assign _zz_11668 = ($signed(_zz_11670) - $signed(_zz_821));
  assign _zz_11669 = ({8'd0,data_mid_72_real} <<< 8);
  assign _zz_11670 = {{8{_zz_11669[23]}}, _zz_11669};
  assign _zz_11671 = fixTo_986_dout;
  assign _zz_11672 = _zz_11673[31 : 0];
  assign _zz_11673 = _zz_11674;
  assign _zz_11674 = ($signed(_zz_11675) >>> _zz_824);
  assign _zz_11675 = _zz_11676;
  assign _zz_11676 = ($signed(_zz_11678) - $signed(_zz_822));
  assign _zz_11677 = ({8'd0,data_mid_72_imag} <<< 8);
  assign _zz_11678 = {{8{_zz_11677[23]}}, _zz_11677};
  assign _zz_11679 = fixTo_987_dout;
  assign _zz_11680 = _zz_11681[31 : 0];
  assign _zz_11681 = _zz_11682;
  assign _zz_11682 = ($signed(_zz_11683) >>> _zz_825);
  assign _zz_11683 = _zz_11684;
  assign _zz_11684 = ($signed(_zz_11686) + $signed(_zz_821));
  assign _zz_11685 = ({8'd0,data_mid_72_real} <<< 8);
  assign _zz_11686 = {{8{_zz_11685[23]}}, _zz_11685};
  assign _zz_11687 = fixTo_988_dout;
  assign _zz_11688 = _zz_11689[31 : 0];
  assign _zz_11689 = _zz_11690;
  assign _zz_11690 = ($signed(_zz_11691) >>> _zz_825);
  assign _zz_11691 = _zz_11692;
  assign _zz_11692 = ($signed(_zz_11694) + $signed(_zz_822));
  assign _zz_11693 = ({8'd0,data_mid_72_imag} <<< 8);
  assign _zz_11694 = {{8{_zz_11693[23]}}, _zz_11693};
  assign _zz_11695 = fixTo_989_dout;
  assign _zz_11696 = ($signed(twiddle_factor_table_4_real) + $signed(twiddle_factor_table_4_imag));
  assign _zz_11697 = ($signed(_zz_828) - $signed(_zz_11698));
  assign _zz_11698 = ($signed(_zz_11699) * $signed(twiddle_factor_table_4_imag));
  assign _zz_11699 = ($signed(data_mid_77_real) + $signed(data_mid_77_imag));
  assign _zz_11700 = fixTo_990_dout;
  assign _zz_11701 = ($signed(_zz_828) + $signed(_zz_11702));
  assign _zz_11702 = ($signed(_zz_11703) * $signed(twiddle_factor_table_4_real));
  assign _zz_11703 = ($signed(data_mid_77_imag) - $signed(data_mid_77_real));
  assign _zz_11704 = fixTo_991_dout;
  assign _zz_11705 = _zz_11706[31 : 0];
  assign _zz_11706 = _zz_11707;
  assign _zz_11707 = ($signed(_zz_11708) >>> _zz_829);
  assign _zz_11708 = _zz_11709;
  assign _zz_11709 = ($signed(_zz_11711) - $signed(_zz_826));
  assign _zz_11710 = ({8'd0,data_mid_73_real} <<< 8);
  assign _zz_11711 = {{8{_zz_11710[23]}}, _zz_11710};
  assign _zz_11712 = fixTo_992_dout;
  assign _zz_11713 = _zz_11714[31 : 0];
  assign _zz_11714 = _zz_11715;
  assign _zz_11715 = ($signed(_zz_11716) >>> _zz_829);
  assign _zz_11716 = _zz_11717;
  assign _zz_11717 = ($signed(_zz_11719) - $signed(_zz_827));
  assign _zz_11718 = ({8'd0,data_mid_73_imag} <<< 8);
  assign _zz_11719 = {{8{_zz_11718[23]}}, _zz_11718};
  assign _zz_11720 = fixTo_993_dout;
  assign _zz_11721 = _zz_11722[31 : 0];
  assign _zz_11722 = _zz_11723;
  assign _zz_11723 = ($signed(_zz_11724) >>> _zz_830);
  assign _zz_11724 = _zz_11725;
  assign _zz_11725 = ($signed(_zz_11727) + $signed(_zz_826));
  assign _zz_11726 = ({8'd0,data_mid_73_real} <<< 8);
  assign _zz_11727 = {{8{_zz_11726[23]}}, _zz_11726};
  assign _zz_11728 = fixTo_994_dout;
  assign _zz_11729 = _zz_11730[31 : 0];
  assign _zz_11730 = _zz_11731;
  assign _zz_11731 = ($signed(_zz_11732) >>> _zz_830);
  assign _zz_11732 = _zz_11733;
  assign _zz_11733 = ($signed(_zz_11735) + $signed(_zz_827));
  assign _zz_11734 = ({8'd0,data_mid_73_imag} <<< 8);
  assign _zz_11735 = {{8{_zz_11734[23]}}, _zz_11734};
  assign _zz_11736 = fixTo_995_dout;
  assign _zz_11737 = ($signed(twiddle_factor_table_5_real) + $signed(twiddle_factor_table_5_imag));
  assign _zz_11738 = ($signed(_zz_833) - $signed(_zz_11739));
  assign _zz_11739 = ($signed(_zz_11740) * $signed(twiddle_factor_table_5_imag));
  assign _zz_11740 = ($signed(data_mid_78_real) + $signed(data_mid_78_imag));
  assign _zz_11741 = fixTo_996_dout;
  assign _zz_11742 = ($signed(_zz_833) + $signed(_zz_11743));
  assign _zz_11743 = ($signed(_zz_11744) * $signed(twiddle_factor_table_5_real));
  assign _zz_11744 = ($signed(data_mid_78_imag) - $signed(data_mid_78_real));
  assign _zz_11745 = fixTo_997_dout;
  assign _zz_11746 = _zz_11747[31 : 0];
  assign _zz_11747 = _zz_11748;
  assign _zz_11748 = ($signed(_zz_11749) >>> _zz_834);
  assign _zz_11749 = _zz_11750;
  assign _zz_11750 = ($signed(_zz_11752) - $signed(_zz_831));
  assign _zz_11751 = ({8'd0,data_mid_74_real} <<< 8);
  assign _zz_11752 = {{8{_zz_11751[23]}}, _zz_11751};
  assign _zz_11753 = fixTo_998_dout;
  assign _zz_11754 = _zz_11755[31 : 0];
  assign _zz_11755 = _zz_11756;
  assign _zz_11756 = ($signed(_zz_11757) >>> _zz_834);
  assign _zz_11757 = _zz_11758;
  assign _zz_11758 = ($signed(_zz_11760) - $signed(_zz_832));
  assign _zz_11759 = ({8'd0,data_mid_74_imag} <<< 8);
  assign _zz_11760 = {{8{_zz_11759[23]}}, _zz_11759};
  assign _zz_11761 = fixTo_999_dout;
  assign _zz_11762 = _zz_11763[31 : 0];
  assign _zz_11763 = _zz_11764;
  assign _zz_11764 = ($signed(_zz_11765) >>> _zz_835);
  assign _zz_11765 = _zz_11766;
  assign _zz_11766 = ($signed(_zz_11768) + $signed(_zz_831));
  assign _zz_11767 = ({8'd0,data_mid_74_real} <<< 8);
  assign _zz_11768 = {{8{_zz_11767[23]}}, _zz_11767};
  assign _zz_11769 = fixTo_1000_dout;
  assign _zz_11770 = _zz_11771[31 : 0];
  assign _zz_11771 = _zz_11772;
  assign _zz_11772 = ($signed(_zz_11773) >>> _zz_835);
  assign _zz_11773 = _zz_11774;
  assign _zz_11774 = ($signed(_zz_11776) + $signed(_zz_832));
  assign _zz_11775 = ({8'd0,data_mid_74_imag} <<< 8);
  assign _zz_11776 = {{8{_zz_11775[23]}}, _zz_11775};
  assign _zz_11777 = fixTo_1001_dout;
  assign _zz_11778 = ($signed(twiddle_factor_table_6_real) + $signed(twiddle_factor_table_6_imag));
  assign _zz_11779 = ($signed(_zz_838) - $signed(_zz_11780));
  assign _zz_11780 = ($signed(_zz_11781) * $signed(twiddle_factor_table_6_imag));
  assign _zz_11781 = ($signed(data_mid_79_real) + $signed(data_mid_79_imag));
  assign _zz_11782 = fixTo_1002_dout;
  assign _zz_11783 = ($signed(_zz_838) + $signed(_zz_11784));
  assign _zz_11784 = ($signed(_zz_11785) * $signed(twiddle_factor_table_6_real));
  assign _zz_11785 = ($signed(data_mid_79_imag) - $signed(data_mid_79_real));
  assign _zz_11786 = fixTo_1003_dout;
  assign _zz_11787 = _zz_11788[31 : 0];
  assign _zz_11788 = _zz_11789;
  assign _zz_11789 = ($signed(_zz_11790) >>> _zz_839);
  assign _zz_11790 = _zz_11791;
  assign _zz_11791 = ($signed(_zz_11793) - $signed(_zz_836));
  assign _zz_11792 = ({8'd0,data_mid_75_real} <<< 8);
  assign _zz_11793 = {{8{_zz_11792[23]}}, _zz_11792};
  assign _zz_11794 = fixTo_1004_dout;
  assign _zz_11795 = _zz_11796[31 : 0];
  assign _zz_11796 = _zz_11797;
  assign _zz_11797 = ($signed(_zz_11798) >>> _zz_839);
  assign _zz_11798 = _zz_11799;
  assign _zz_11799 = ($signed(_zz_11801) - $signed(_zz_837));
  assign _zz_11800 = ({8'd0,data_mid_75_imag} <<< 8);
  assign _zz_11801 = {{8{_zz_11800[23]}}, _zz_11800};
  assign _zz_11802 = fixTo_1005_dout;
  assign _zz_11803 = _zz_11804[31 : 0];
  assign _zz_11804 = _zz_11805;
  assign _zz_11805 = ($signed(_zz_11806) >>> _zz_840);
  assign _zz_11806 = _zz_11807;
  assign _zz_11807 = ($signed(_zz_11809) + $signed(_zz_836));
  assign _zz_11808 = ({8'd0,data_mid_75_real} <<< 8);
  assign _zz_11809 = {{8{_zz_11808[23]}}, _zz_11808};
  assign _zz_11810 = fixTo_1006_dout;
  assign _zz_11811 = _zz_11812[31 : 0];
  assign _zz_11812 = _zz_11813;
  assign _zz_11813 = ($signed(_zz_11814) >>> _zz_840);
  assign _zz_11814 = _zz_11815;
  assign _zz_11815 = ($signed(_zz_11817) + $signed(_zz_837));
  assign _zz_11816 = ({8'd0,data_mid_75_imag} <<< 8);
  assign _zz_11817 = {{8{_zz_11816[23]}}, _zz_11816};
  assign _zz_11818 = fixTo_1007_dout;
  assign _zz_11819 = ($signed(twiddle_factor_table_3_real) + $signed(twiddle_factor_table_3_imag));
  assign _zz_11820 = ($signed(_zz_843) - $signed(_zz_11821));
  assign _zz_11821 = ($signed(_zz_11822) * $signed(twiddle_factor_table_3_imag));
  assign _zz_11822 = ($signed(data_mid_84_real) + $signed(data_mid_84_imag));
  assign _zz_11823 = fixTo_1008_dout;
  assign _zz_11824 = ($signed(_zz_843) + $signed(_zz_11825));
  assign _zz_11825 = ($signed(_zz_11826) * $signed(twiddle_factor_table_3_real));
  assign _zz_11826 = ($signed(data_mid_84_imag) - $signed(data_mid_84_real));
  assign _zz_11827 = fixTo_1009_dout;
  assign _zz_11828 = _zz_11829[31 : 0];
  assign _zz_11829 = _zz_11830;
  assign _zz_11830 = ($signed(_zz_11831) >>> _zz_844);
  assign _zz_11831 = _zz_11832;
  assign _zz_11832 = ($signed(_zz_11834) - $signed(_zz_841));
  assign _zz_11833 = ({8'd0,data_mid_80_real} <<< 8);
  assign _zz_11834 = {{8{_zz_11833[23]}}, _zz_11833};
  assign _zz_11835 = fixTo_1010_dout;
  assign _zz_11836 = _zz_11837[31 : 0];
  assign _zz_11837 = _zz_11838;
  assign _zz_11838 = ($signed(_zz_11839) >>> _zz_844);
  assign _zz_11839 = _zz_11840;
  assign _zz_11840 = ($signed(_zz_11842) - $signed(_zz_842));
  assign _zz_11841 = ({8'd0,data_mid_80_imag} <<< 8);
  assign _zz_11842 = {{8{_zz_11841[23]}}, _zz_11841};
  assign _zz_11843 = fixTo_1011_dout;
  assign _zz_11844 = _zz_11845[31 : 0];
  assign _zz_11845 = _zz_11846;
  assign _zz_11846 = ($signed(_zz_11847) >>> _zz_845);
  assign _zz_11847 = _zz_11848;
  assign _zz_11848 = ($signed(_zz_11850) + $signed(_zz_841));
  assign _zz_11849 = ({8'd0,data_mid_80_real} <<< 8);
  assign _zz_11850 = {{8{_zz_11849[23]}}, _zz_11849};
  assign _zz_11851 = fixTo_1012_dout;
  assign _zz_11852 = _zz_11853[31 : 0];
  assign _zz_11853 = _zz_11854;
  assign _zz_11854 = ($signed(_zz_11855) >>> _zz_845);
  assign _zz_11855 = _zz_11856;
  assign _zz_11856 = ($signed(_zz_11858) + $signed(_zz_842));
  assign _zz_11857 = ({8'd0,data_mid_80_imag} <<< 8);
  assign _zz_11858 = {{8{_zz_11857[23]}}, _zz_11857};
  assign _zz_11859 = fixTo_1013_dout;
  assign _zz_11860 = ($signed(twiddle_factor_table_4_real) + $signed(twiddle_factor_table_4_imag));
  assign _zz_11861 = ($signed(_zz_848) - $signed(_zz_11862));
  assign _zz_11862 = ($signed(_zz_11863) * $signed(twiddle_factor_table_4_imag));
  assign _zz_11863 = ($signed(data_mid_85_real) + $signed(data_mid_85_imag));
  assign _zz_11864 = fixTo_1014_dout;
  assign _zz_11865 = ($signed(_zz_848) + $signed(_zz_11866));
  assign _zz_11866 = ($signed(_zz_11867) * $signed(twiddle_factor_table_4_real));
  assign _zz_11867 = ($signed(data_mid_85_imag) - $signed(data_mid_85_real));
  assign _zz_11868 = fixTo_1015_dout;
  assign _zz_11869 = _zz_11870[31 : 0];
  assign _zz_11870 = _zz_11871;
  assign _zz_11871 = ($signed(_zz_11872) >>> _zz_849);
  assign _zz_11872 = _zz_11873;
  assign _zz_11873 = ($signed(_zz_11875) - $signed(_zz_846));
  assign _zz_11874 = ({8'd0,data_mid_81_real} <<< 8);
  assign _zz_11875 = {{8{_zz_11874[23]}}, _zz_11874};
  assign _zz_11876 = fixTo_1016_dout;
  assign _zz_11877 = _zz_11878[31 : 0];
  assign _zz_11878 = _zz_11879;
  assign _zz_11879 = ($signed(_zz_11880) >>> _zz_849);
  assign _zz_11880 = _zz_11881;
  assign _zz_11881 = ($signed(_zz_11883) - $signed(_zz_847));
  assign _zz_11882 = ({8'd0,data_mid_81_imag} <<< 8);
  assign _zz_11883 = {{8{_zz_11882[23]}}, _zz_11882};
  assign _zz_11884 = fixTo_1017_dout;
  assign _zz_11885 = _zz_11886[31 : 0];
  assign _zz_11886 = _zz_11887;
  assign _zz_11887 = ($signed(_zz_11888) >>> _zz_850);
  assign _zz_11888 = _zz_11889;
  assign _zz_11889 = ($signed(_zz_11891) + $signed(_zz_846));
  assign _zz_11890 = ({8'd0,data_mid_81_real} <<< 8);
  assign _zz_11891 = {{8{_zz_11890[23]}}, _zz_11890};
  assign _zz_11892 = fixTo_1018_dout;
  assign _zz_11893 = _zz_11894[31 : 0];
  assign _zz_11894 = _zz_11895;
  assign _zz_11895 = ($signed(_zz_11896) >>> _zz_850);
  assign _zz_11896 = _zz_11897;
  assign _zz_11897 = ($signed(_zz_11899) + $signed(_zz_847));
  assign _zz_11898 = ({8'd0,data_mid_81_imag} <<< 8);
  assign _zz_11899 = {{8{_zz_11898[23]}}, _zz_11898};
  assign _zz_11900 = fixTo_1019_dout;
  assign _zz_11901 = ($signed(twiddle_factor_table_5_real) + $signed(twiddle_factor_table_5_imag));
  assign _zz_11902 = ($signed(_zz_853) - $signed(_zz_11903));
  assign _zz_11903 = ($signed(_zz_11904) * $signed(twiddle_factor_table_5_imag));
  assign _zz_11904 = ($signed(data_mid_86_real) + $signed(data_mid_86_imag));
  assign _zz_11905 = fixTo_1020_dout;
  assign _zz_11906 = ($signed(_zz_853) + $signed(_zz_11907));
  assign _zz_11907 = ($signed(_zz_11908) * $signed(twiddle_factor_table_5_real));
  assign _zz_11908 = ($signed(data_mid_86_imag) - $signed(data_mid_86_real));
  assign _zz_11909 = fixTo_1021_dout;
  assign _zz_11910 = _zz_11911[31 : 0];
  assign _zz_11911 = _zz_11912;
  assign _zz_11912 = ($signed(_zz_11913) >>> _zz_854);
  assign _zz_11913 = _zz_11914;
  assign _zz_11914 = ($signed(_zz_11916) - $signed(_zz_851));
  assign _zz_11915 = ({8'd0,data_mid_82_real} <<< 8);
  assign _zz_11916 = {{8{_zz_11915[23]}}, _zz_11915};
  assign _zz_11917 = fixTo_1022_dout;
  assign _zz_11918 = _zz_11919[31 : 0];
  assign _zz_11919 = _zz_11920;
  assign _zz_11920 = ($signed(_zz_11921) >>> _zz_854);
  assign _zz_11921 = _zz_11922;
  assign _zz_11922 = ($signed(_zz_11924) - $signed(_zz_852));
  assign _zz_11923 = ({8'd0,data_mid_82_imag} <<< 8);
  assign _zz_11924 = {{8{_zz_11923[23]}}, _zz_11923};
  assign _zz_11925 = fixTo_1023_dout;
  assign _zz_11926 = _zz_11927[31 : 0];
  assign _zz_11927 = _zz_11928;
  assign _zz_11928 = ($signed(_zz_11929) >>> _zz_855);
  assign _zz_11929 = _zz_11930;
  assign _zz_11930 = ($signed(_zz_11932) + $signed(_zz_851));
  assign _zz_11931 = ({8'd0,data_mid_82_real} <<< 8);
  assign _zz_11932 = {{8{_zz_11931[23]}}, _zz_11931};
  assign _zz_11933 = fixTo_1024_dout;
  assign _zz_11934 = _zz_11935[31 : 0];
  assign _zz_11935 = _zz_11936;
  assign _zz_11936 = ($signed(_zz_11937) >>> _zz_855);
  assign _zz_11937 = _zz_11938;
  assign _zz_11938 = ($signed(_zz_11940) + $signed(_zz_852));
  assign _zz_11939 = ({8'd0,data_mid_82_imag} <<< 8);
  assign _zz_11940 = {{8{_zz_11939[23]}}, _zz_11939};
  assign _zz_11941 = fixTo_1025_dout;
  assign _zz_11942 = ($signed(twiddle_factor_table_6_real) + $signed(twiddle_factor_table_6_imag));
  assign _zz_11943 = ($signed(_zz_858) - $signed(_zz_11944));
  assign _zz_11944 = ($signed(_zz_11945) * $signed(twiddle_factor_table_6_imag));
  assign _zz_11945 = ($signed(data_mid_87_real) + $signed(data_mid_87_imag));
  assign _zz_11946 = fixTo_1026_dout;
  assign _zz_11947 = ($signed(_zz_858) + $signed(_zz_11948));
  assign _zz_11948 = ($signed(_zz_11949) * $signed(twiddle_factor_table_6_real));
  assign _zz_11949 = ($signed(data_mid_87_imag) - $signed(data_mid_87_real));
  assign _zz_11950 = fixTo_1027_dout;
  assign _zz_11951 = _zz_11952[31 : 0];
  assign _zz_11952 = _zz_11953;
  assign _zz_11953 = ($signed(_zz_11954) >>> _zz_859);
  assign _zz_11954 = _zz_11955;
  assign _zz_11955 = ($signed(_zz_11957) - $signed(_zz_856));
  assign _zz_11956 = ({8'd0,data_mid_83_real} <<< 8);
  assign _zz_11957 = {{8{_zz_11956[23]}}, _zz_11956};
  assign _zz_11958 = fixTo_1028_dout;
  assign _zz_11959 = _zz_11960[31 : 0];
  assign _zz_11960 = _zz_11961;
  assign _zz_11961 = ($signed(_zz_11962) >>> _zz_859);
  assign _zz_11962 = _zz_11963;
  assign _zz_11963 = ($signed(_zz_11965) - $signed(_zz_857));
  assign _zz_11964 = ({8'd0,data_mid_83_imag} <<< 8);
  assign _zz_11965 = {{8{_zz_11964[23]}}, _zz_11964};
  assign _zz_11966 = fixTo_1029_dout;
  assign _zz_11967 = _zz_11968[31 : 0];
  assign _zz_11968 = _zz_11969;
  assign _zz_11969 = ($signed(_zz_11970) >>> _zz_860);
  assign _zz_11970 = _zz_11971;
  assign _zz_11971 = ($signed(_zz_11973) + $signed(_zz_856));
  assign _zz_11972 = ({8'd0,data_mid_83_real} <<< 8);
  assign _zz_11973 = {{8{_zz_11972[23]}}, _zz_11972};
  assign _zz_11974 = fixTo_1030_dout;
  assign _zz_11975 = _zz_11976[31 : 0];
  assign _zz_11976 = _zz_11977;
  assign _zz_11977 = ($signed(_zz_11978) >>> _zz_860);
  assign _zz_11978 = _zz_11979;
  assign _zz_11979 = ($signed(_zz_11981) + $signed(_zz_857));
  assign _zz_11980 = ({8'd0,data_mid_83_imag} <<< 8);
  assign _zz_11981 = {{8{_zz_11980[23]}}, _zz_11980};
  assign _zz_11982 = fixTo_1031_dout;
  assign _zz_11983 = ($signed(twiddle_factor_table_3_real) + $signed(twiddle_factor_table_3_imag));
  assign _zz_11984 = ($signed(_zz_863) - $signed(_zz_11985));
  assign _zz_11985 = ($signed(_zz_11986) * $signed(twiddle_factor_table_3_imag));
  assign _zz_11986 = ($signed(data_mid_92_real) + $signed(data_mid_92_imag));
  assign _zz_11987 = fixTo_1032_dout;
  assign _zz_11988 = ($signed(_zz_863) + $signed(_zz_11989));
  assign _zz_11989 = ($signed(_zz_11990) * $signed(twiddle_factor_table_3_real));
  assign _zz_11990 = ($signed(data_mid_92_imag) - $signed(data_mid_92_real));
  assign _zz_11991 = fixTo_1033_dout;
  assign _zz_11992 = _zz_11993[31 : 0];
  assign _zz_11993 = _zz_11994;
  assign _zz_11994 = ($signed(_zz_11995) >>> _zz_864);
  assign _zz_11995 = _zz_11996;
  assign _zz_11996 = ($signed(_zz_11998) - $signed(_zz_861));
  assign _zz_11997 = ({8'd0,data_mid_88_real} <<< 8);
  assign _zz_11998 = {{8{_zz_11997[23]}}, _zz_11997};
  assign _zz_11999 = fixTo_1034_dout;
  assign _zz_12000 = _zz_12001[31 : 0];
  assign _zz_12001 = _zz_12002;
  assign _zz_12002 = ($signed(_zz_12003) >>> _zz_864);
  assign _zz_12003 = _zz_12004;
  assign _zz_12004 = ($signed(_zz_12006) - $signed(_zz_862));
  assign _zz_12005 = ({8'd0,data_mid_88_imag} <<< 8);
  assign _zz_12006 = {{8{_zz_12005[23]}}, _zz_12005};
  assign _zz_12007 = fixTo_1035_dout;
  assign _zz_12008 = _zz_12009[31 : 0];
  assign _zz_12009 = _zz_12010;
  assign _zz_12010 = ($signed(_zz_12011) >>> _zz_865);
  assign _zz_12011 = _zz_12012;
  assign _zz_12012 = ($signed(_zz_12014) + $signed(_zz_861));
  assign _zz_12013 = ({8'd0,data_mid_88_real} <<< 8);
  assign _zz_12014 = {{8{_zz_12013[23]}}, _zz_12013};
  assign _zz_12015 = fixTo_1036_dout;
  assign _zz_12016 = _zz_12017[31 : 0];
  assign _zz_12017 = _zz_12018;
  assign _zz_12018 = ($signed(_zz_12019) >>> _zz_865);
  assign _zz_12019 = _zz_12020;
  assign _zz_12020 = ($signed(_zz_12022) + $signed(_zz_862));
  assign _zz_12021 = ({8'd0,data_mid_88_imag} <<< 8);
  assign _zz_12022 = {{8{_zz_12021[23]}}, _zz_12021};
  assign _zz_12023 = fixTo_1037_dout;
  assign _zz_12024 = ($signed(twiddle_factor_table_4_real) + $signed(twiddle_factor_table_4_imag));
  assign _zz_12025 = ($signed(_zz_868) - $signed(_zz_12026));
  assign _zz_12026 = ($signed(_zz_12027) * $signed(twiddle_factor_table_4_imag));
  assign _zz_12027 = ($signed(data_mid_93_real) + $signed(data_mid_93_imag));
  assign _zz_12028 = fixTo_1038_dout;
  assign _zz_12029 = ($signed(_zz_868) + $signed(_zz_12030));
  assign _zz_12030 = ($signed(_zz_12031) * $signed(twiddle_factor_table_4_real));
  assign _zz_12031 = ($signed(data_mid_93_imag) - $signed(data_mid_93_real));
  assign _zz_12032 = fixTo_1039_dout;
  assign _zz_12033 = _zz_12034[31 : 0];
  assign _zz_12034 = _zz_12035;
  assign _zz_12035 = ($signed(_zz_12036) >>> _zz_869);
  assign _zz_12036 = _zz_12037;
  assign _zz_12037 = ($signed(_zz_12039) - $signed(_zz_866));
  assign _zz_12038 = ({8'd0,data_mid_89_real} <<< 8);
  assign _zz_12039 = {{8{_zz_12038[23]}}, _zz_12038};
  assign _zz_12040 = fixTo_1040_dout;
  assign _zz_12041 = _zz_12042[31 : 0];
  assign _zz_12042 = _zz_12043;
  assign _zz_12043 = ($signed(_zz_12044) >>> _zz_869);
  assign _zz_12044 = _zz_12045;
  assign _zz_12045 = ($signed(_zz_12047) - $signed(_zz_867));
  assign _zz_12046 = ({8'd0,data_mid_89_imag} <<< 8);
  assign _zz_12047 = {{8{_zz_12046[23]}}, _zz_12046};
  assign _zz_12048 = fixTo_1041_dout;
  assign _zz_12049 = _zz_12050[31 : 0];
  assign _zz_12050 = _zz_12051;
  assign _zz_12051 = ($signed(_zz_12052) >>> _zz_870);
  assign _zz_12052 = _zz_12053;
  assign _zz_12053 = ($signed(_zz_12055) + $signed(_zz_866));
  assign _zz_12054 = ({8'd0,data_mid_89_real} <<< 8);
  assign _zz_12055 = {{8{_zz_12054[23]}}, _zz_12054};
  assign _zz_12056 = fixTo_1042_dout;
  assign _zz_12057 = _zz_12058[31 : 0];
  assign _zz_12058 = _zz_12059;
  assign _zz_12059 = ($signed(_zz_12060) >>> _zz_870);
  assign _zz_12060 = _zz_12061;
  assign _zz_12061 = ($signed(_zz_12063) + $signed(_zz_867));
  assign _zz_12062 = ({8'd0,data_mid_89_imag} <<< 8);
  assign _zz_12063 = {{8{_zz_12062[23]}}, _zz_12062};
  assign _zz_12064 = fixTo_1043_dout;
  assign _zz_12065 = ($signed(twiddle_factor_table_5_real) + $signed(twiddle_factor_table_5_imag));
  assign _zz_12066 = ($signed(_zz_873) - $signed(_zz_12067));
  assign _zz_12067 = ($signed(_zz_12068) * $signed(twiddle_factor_table_5_imag));
  assign _zz_12068 = ($signed(data_mid_94_real) + $signed(data_mid_94_imag));
  assign _zz_12069 = fixTo_1044_dout;
  assign _zz_12070 = ($signed(_zz_873) + $signed(_zz_12071));
  assign _zz_12071 = ($signed(_zz_12072) * $signed(twiddle_factor_table_5_real));
  assign _zz_12072 = ($signed(data_mid_94_imag) - $signed(data_mid_94_real));
  assign _zz_12073 = fixTo_1045_dout;
  assign _zz_12074 = _zz_12075[31 : 0];
  assign _zz_12075 = _zz_12076;
  assign _zz_12076 = ($signed(_zz_12077) >>> _zz_874);
  assign _zz_12077 = _zz_12078;
  assign _zz_12078 = ($signed(_zz_12080) - $signed(_zz_871));
  assign _zz_12079 = ({8'd0,data_mid_90_real} <<< 8);
  assign _zz_12080 = {{8{_zz_12079[23]}}, _zz_12079};
  assign _zz_12081 = fixTo_1046_dout;
  assign _zz_12082 = _zz_12083[31 : 0];
  assign _zz_12083 = _zz_12084;
  assign _zz_12084 = ($signed(_zz_12085) >>> _zz_874);
  assign _zz_12085 = _zz_12086;
  assign _zz_12086 = ($signed(_zz_12088) - $signed(_zz_872));
  assign _zz_12087 = ({8'd0,data_mid_90_imag} <<< 8);
  assign _zz_12088 = {{8{_zz_12087[23]}}, _zz_12087};
  assign _zz_12089 = fixTo_1047_dout;
  assign _zz_12090 = _zz_12091[31 : 0];
  assign _zz_12091 = _zz_12092;
  assign _zz_12092 = ($signed(_zz_12093) >>> _zz_875);
  assign _zz_12093 = _zz_12094;
  assign _zz_12094 = ($signed(_zz_12096) + $signed(_zz_871));
  assign _zz_12095 = ({8'd0,data_mid_90_real} <<< 8);
  assign _zz_12096 = {{8{_zz_12095[23]}}, _zz_12095};
  assign _zz_12097 = fixTo_1048_dout;
  assign _zz_12098 = _zz_12099[31 : 0];
  assign _zz_12099 = _zz_12100;
  assign _zz_12100 = ($signed(_zz_12101) >>> _zz_875);
  assign _zz_12101 = _zz_12102;
  assign _zz_12102 = ($signed(_zz_12104) + $signed(_zz_872));
  assign _zz_12103 = ({8'd0,data_mid_90_imag} <<< 8);
  assign _zz_12104 = {{8{_zz_12103[23]}}, _zz_12103};
  assign _zz_12105 = fixTo_1049_dout;
  assign _zz_12106 = ($signed(twiddle_factor_table_6_real) + $signed(twiddle_factor_table_6_imag));
  assign _zz_12107 = ($signed(_zz_878) - $signed(_zz_12108));
  assign _zz_12108 = ($signed(_zz_12109) * $signed(twiddle_factor_table_6_imag));
  assign _zz_12109 = ($signed(data_mid_95_real) + $signed(data_mid_95_imag));
  assign _zz_12110 = fixTo_1050_dout;
  assign _zz_12111 = ($signed(_zz_878) + $signed(_zz_12112));
  assign _zz_12112 = ($signed(_zz_12113) * $signed(twiddle_factor_table_6_real));
  assign _zz_12113 = ($signed(data_mid_95_imag) - $signed(data_mid_95_real));
  assign _zz_12114 = fixTo_1051_dout;
  assign _zz_12115 = _zz_12116[31 : 0];
  assign _zz_12116 = _zz_12117;
  assign _zz_12117 = ($signed(_zz_12118) >>> _zz_879);
  assign _zz_12118 = _zz_12119;
  assign _zz_12119 = ($signed(_zz_12121) - $signed(_zz_876));
  assign _zz_12120 = ({8'd0,data_mid_91_real} <<< 8);
  assign _zz_12121 = {{8{_zz_12120[23]}}, _zz_12120};
  assign _zz_12122 = fixTo_1052_dout;
  assign _zz_12123 = _zz_12124[31 : 0];
  assign _zz_12124 = _zz_12125;
  assign _zz_12125 = ($signed(_zz_12126) >>> _zz_879);
  assign _zz_12126 = _zz_12127;
  assign _zz_12127 = ($signed(_zz_12129) - $signed(_zz_877));
  assign _zz_12128 = ({8'd0,data_mid_91_imag} <<< 8);
  assign _zz_12129 = {{8{_zz_12128[23]}}, _zz_12128};
  assign _zz_12130 = fixTo_1053_dout;
  assign _zz_12131 = _zz_12132[31 : 0];
  assign _zz_12132 = _zz_12133;
  assign _zz_12133 = ($signed(_zz_12134) >>> _zz_880);
  assign _zz_12134 = _zz_12135;
  assign _zz_12135 = ($signed(_zz_12137) + $signed(_zz_876));
  assign _zz_12136 = ({8'd0,data_mid_91_real} <<< 8);
  assign _zz_12137 = {{8{_zz_12136[23]}}, _zz_12136};
  assign _zz_12138 = fixTo_1054_dout;
  assign _zz_12139 = _zz_12140[31 : 0];
  assign _zz_12140 = _zz_12141;
  assign _zz_12141 = ($signed(_zz_12142) >>> _zz_880);
  assign _zz_12142 = _zz_12143;
  assign _zz_12143 = ($signed(_zz_12145) + $signed(_zz_877));
  assign _zz_12144 = ({8'd0,data_mid_91_imag} <<< 8);
  assign _zz_12145 = {{8{_zz_12144[23]}}, _zz_12144};
  assign _zz_12146 = fixTo_1055_dout;
  assign _zz_12147 = ($signed(twiddle_factor_table_3_real) + $signed(twiddle_factor_table_3_imag));
  assign _zz_12148 = ($signed(_zz_883) - $signed(_zz_12149));
  assign _zz_12149 = ($signed(_zz_12150) * $signed(twiddle_factor_table_3_imag));
  assign _zz_12150 = ($signed(data_mid_100_real) + $signed(data_mid_100_imag));
  assign _zz_12151 = fixTo_1056_dout;
  assign _zz_12152 = ($signed(_zz_883) + $signed(_zz_12153));
  assign _zz_12153 = ($signed(_zz_12154) * $signed(twiddle_factor_table_3_real));
  assign _zz_12154 = ($signed(data_mid_100_imag) - $signed(data_mid_100_real));
  assign _zz_12155 = fixTo_1057_dout;
  assign _zz_12156 = _zz_12157[31 : 0];
  assign _zz_12157 = _zz_12158;
  assign _zz_12158 = ($signed(_zz_12159) >>> _zz_884);
  assign _zz_12159 = _zz_12160;
  assign _zz_12160 = ($signed(_zz_12162) - $signed(_zz_881));
  assign _zz_12161 = ({8'd0,data_mid_96_real} <<< 8);
  assign _zz_12162 = {{8{_zz_12161[23]}}, _zz_12161};
  assign _zz_12163 = fixTo_1058_dout;
  assign _zz_12164 = _zz_12165[31 : 0];
  assign _zz_12165 = _zz_12166;
  assign _zz_12166 = ($signed(_zz_12167) >>> _zz_884);
  assign _zz_12167 = _zz_12168;
  assign _zz_12168 = ($signed(_zz_12170) - $signed(_zz_882));
  assign _zz_12169 = ({8'd0,data_mid_96_imag} <<< 8);
  assign _zz_12170 = {{8{_zz_12169[23]}}, _zz_12169};
  assign _zz_12171 = fixTo_1059_dout;
  assign _zz_12172 = _zz_12173[31 : 0];
  assign _zz_12173 = _zz_12174;
  assign _zz_12174 = ($signed(_zz_12175) >>> _zz_885);
  assign _zz_12175 = _zz_12176;
  assign _zz_12176 = ($signed(_zz_12178) + $signed(_zz_881));
  assign _zz_12177 = ({8'd0,data_mid_96_real} <<< 8);
  assign _zz_12178 = {{8{_zz_12177[23]}}, _zz_12177};
  assign _zz_12179 = fixTo_1060_dout;
  assign _zz_12180 = _zz_12181[31 : 0];
  assign _zz_12181 = _zz_12182;
  assign _zz_12182 = ($signed(_zz_12183) >>> _zz_885);
  assign _zz_12183 = _zz_12184;
  assign _zz_12184 = ($signed(_zz_12186) + $signed(_zz_882));
  assign _zz_12185 = ({8'd0,data_mid_96_imag} <<< 8);
  assign _zz_12186 = {{8{_zz_12185[23]}}, _zz_12185};
  assign _zz_12187 = fixTo_1061_dout;
  assign _zz_12188 = ($signed(twiddle_factor_table_4_real) + $signed(twiddle_factor_table_4_imag));
  assign _zz_12189 = ($signed(_zz_888) - $signed(_zz_12190));
  assign _zz_12190 = ($signed(_zz_12191) * $signed(twiddle_factor_table_4_imag));
  assign _zz_12191 = ($signed(data_mid_101_real) + $signed(data_mid_101_imag));
  assign _zz_12192 = fixTo_1062_dout;
  assign _zz_12193 = ($signed(_zz_888) + $signed(_zz_12194));
  assign _zz_12194 = ($signed(_zz_12195) * $signed(twiddle_factor_table_4_real));
  assign _zz_12195 = ($signed(data_mid_101_imag) - $signed(data_mid_101_real));
  assign _zz_12196 = fixTo_1063_dout;
  assign _zz_12197 = _zz_12198[31 : 0];
  assign _zz_12198 = _zz_12199;
  assign _zz_12199 = ($signed(_zz_12200) >>> _zz_889);
  assign _zz_12200 = _zz_12201;
  assign _zz_12201 = ($signed(_zz_12203) - $signed(_zz_886));
  assign _zz_12202 = ({8'd0,data_mid_97_real} <<< 8);
  assign _zz_12203 = {{8{_zz_12202[23]}}, _zz_12202};
  assign _zz_12204 = fixTo_1064_dout;
  assign _zz_12205 = _zz_12206[31 : 0];
  assign _zz_12206 = _zz_12207;
  assign _zz_12207 = ($signed(_zz_12208) >>> _zz_889);
  assign _zz_12208 = _zz_12209;
  assign _zz_12209 = ($signed(_zz_12211) - $signed(_zz_887));
  assign _zz_12210 = ({8'd0,data_mid_97_imag} <<< 8);
  assign _zz_12211 = {{8{_zz_12210[23]}}, _zz_12210};
  assign _zz_12212 = fixTo_1065_dout;
  assign _zz_12213 = _zz_12214[31 : 0];
  assign _zz_12214 = _zz_12215;
  assign _zz_12215 = ($signed(_zz_12216) >>> _zz_890);
  assign _zz_12216 = _zz_12217;
  assign _zz_12217 = ($signed(_zz_12219) + $signed(_zz_886));
  assign _zz_12218 = ({8'd0,data_mid_97_real} <<< 8);
  assign _zz_12219 = {{8{_zz_12218[23]}}, _zz_12218};
  assign _zz_12220 = fixTo_1066_dout;
  assign _zz_12221 = _zz_12222[31 : 0];
  assign _zz_12222 = _zz_12223;
  assign _zz_12223 = ($signed(_zz_12224) >>> _zz_890);
  assign _zz_12224 = _zz_12225;
  assign _zz_12225 = ($signed(_zz_12227) + $signed(_zz_887));
  assign _zz_12226 = ({8'd0,data_mid_97_imag} <<< 8);
  assign _zz_12227 = {{8{_zz_12226[23]}}, _zz_12226};
  assign _zz_12228 = fixTo_1067_dout;
  assign _zz_12229 = ($signed(twiddle_factor_table_5_real) + $signed(twiddle_factor_table_5_imag));
  assign _zz_12230 = ($signed(_zz_893) - $signed(_zz_12231));
  assign _zz_12231 = ($signed(_zz_12232) * $signed(twiddle_factor_table_5_imag));
  assign _zz_12232 = ($signed(data_mid_102_real) + $signed(data_mid_102_imag));
  assign _zz_12233 = fixTo_1068_dout;
  assign _zz_12234 = ($signed(_zz_893) + $signed(_zz_12235));
  assign _zz_12235 = ($signed(_zz_12236) * $signed(twiddle_factor_table_5_real));
  assign _zz_12236 = ($signed(data_mid_102_imag) - $signed(data_mid_102_real));
  assign _zz_12237 = fixTo_1069_dout;
  assign _zz_12238 = _zz_12239[31 : 0];
  assign _zz_12239 = _zz_12240;
  assign _zz_12240 = ($signed(_zz_12241) >>> _zz_894);
  assign _zz_12241 = _zz_12242;
  assign _zz_12242 = ($signed(_zz_12244) - $signed(_zz_891));
  assign _zz_12243 = ({8'd0,data_mid_98_real} <<< 8);
  assign _zz_12244 = {{8{_zz_12243[23]}}, _zz_12243};
  assign _zz_12245 = fixTo_1070_dout;
  assign _zz_12246 = _zz_12247[31 : 0];
  assign _zz_12247 = _zz_12248;
  assign _zz_12248 = ($signed(_zz_12249) >>> _zz_894);
  assign _zz_12249 = _zz_12250;
  assign _zz_12250 = ($signed(_zz_12252) - $signed(_zz_892));
  assign _zz_12251 = ({8'd0,data_mid_98_imag} <<< 8);
  assign _zz_12252 = {{8{_zz_12251[23]}}, _zz_12251};
  assign _zz_12253 = fixTo_1071_dout;
  assign _zz_12254 = _zz_12255[31 : 0];
  assign _zz_12255 = _zz_12256;
  assign _zz_12256 = ($signed(_zz_12257) >>> _zz_895);
  assign _zz_12257 = _zz_12258;
  assign _zz_12258 = ($signed(_zz_12260) + $signed(_zz_891));
  assign _zz_12259 = ({8'd0,data_mid_98_real} <<< 8);
  assign _zz_12260 = {{8{_zz_12259[23]}}, _zz_12259};
  assign _zz_12261 = fixTo_1072_dout;
  assign _zz_12262 = _zz_12263[31 : 0];
  assign _zz_12263 = _zz_12264;
  assign _zz_12264 = ($signed(_zz_12265) >>> _zz_895);
  assign _zz_12265 = _zz_12266;
  assign _zz_12266 = ($signed(_zz_12268) + $signed(_zz_892));
  assign _zz_12267 = ({8'd0,data_mid_98_imag} <<< 8);
  assign _zz_12268 = {{8{_zz_12267[23]}}, _zz_12267};
  assign _zz_12269 = fixTo_1073_dout;
  assign _zz_12270 = ($signed(twiddle_factor_table_6_real) + $signed(twiddle_factor_table_6_imag));
  assign _zz_12271 = ($signed(_zz_898) - $signed(_zz_12272));
  assign _zz_12272 = ($signed(_zz_12273) * $signed(twiddle_factor_table_6_imag));
  assign _zz_12273 = ($signed(data_mid_103_real) + $signed(data_mid_103_imag));
  assign _zz_12274 = fixTo_1074_dout;
  assign _zz_12275 = ($signed(_zz_898) + $signed(_zz_12276));
  assign _zz_12276 = ($signed(_zz_12277) * $signed(twiddle_factor_table_6_real));
  assign _zz_12277 = ($signed(data_mid_103_imag) - $signed(data_mid_103_real));
  assign _zz_12278 = fixTo_1075_dout;
  assign _zz_12279 = _zz_12280[31 : 0];
  assign _zz_12280 = _zz_12281;
  assign _zz_12281 = ($signed(_zz_12282) >>> _zz_899);
  assign _zz_12282 = _zz_12283;
  assign _zz_12283 = ($signed(_zz_12285) - $signed(_zz_896));
  assign _zz_12284 = ({8'd0,data_mid_99_real} <<< 8);
  assign _zz_12285 = {{8{_zz_12284[23]}}, _zz_12284};
  assign _zz_12286 = fixTo_1076_dout;
  assign _zz_12287 = _zz_12288[31 : 0];
  assign _zz_12288 = _zz_12289;
  assign _zz_12289 = ($signed(_zz_12290) >>> _zz_899);
  assign _zz_12290 = _zz_12291;
  assign _zz_12291 = ($signed(_zz_12293) - $signed(_zz_897));
  assign _zz_12292 = ({8'd0,data_mid_99_imag} <<< 8);
  assign _zz_12293 = {{8{_zz_12292[23]}}, _zz_12292};
  assign _zz_12294 = fixTo_1077_dout;
  assign _zz_12295 = _zz_12296[31 : 0];
  assign _zz_12296 = _zz_12297;
  assign _zz_12297 = ($signed(_zz_12298) >>> _zz_900);
  assign _zz_12298 = _zz_12299;
  assign _zz_12299 = ($signed(_zz_12301) + $signed(_zz_896));
  assign _zz_12300 = ({8'd0,data_mid_99_real} <<< 8);
  assign _zz_12301 = {{8{_zz_12300[23]}}, _zz_12300};
  assign _zz_12302 = fixTo_1078_dout;
  assign _zz_12303 = _zz_12304[31 : 0];
  assign _zz_12304 = _zz_12305;
  assign _zz_12305 = ($signed(_zz_12306) >>> _zz_900);
  assign _zz_12306 = _zz_12307;
  assign _zz_12307 = ($signed(_zz_12309) + $signed(_zz_897));
  assign _zz_12308 = ({8'd0,data_mid_99_imag} <<< 8);
  assign _zz_12309 = {{8{_zz_12308[23]}}, _zz_12308};
  assign _zz_12310 = fixTo_1079_dout;
  assign _zz_12311 = ($signed(twiddle_factor_table_3_real) + $signed(twiddle_factor_table_3_imag));
  assign _zz_12312 = ($signed(_zz_903) - $signed(_zz_12313));
  assign _zz_12313 = ($signed(_zz_12314) * $signed(twiddle_factor_table_3_imag));
  assign _zz_12314 = ($signed(data_mid_108_real) + $signed(data_mid_108_imag));
  assign _zz_12315 = fixTo_1080_dout;
  assign _zz_12316 = ($signed(_zz_903) + $signed(_zz_12317));
  assign _zz_12317 = ($signed(_zz_12318) * $signed(twiddle_factor_table_3_real));
  assign _zz_12318 = ($signed(data_mid_108_imag) - $signed(data_mid_108_real));
  assign _zz_12319 = fixTo_1081_dout;
  assign _zz_12320 = _zz_12321[31 : 0];
  assign _zz_12321 = _zz_12322;
  assign _zz_12322 = ($signed(_zz_12323) >>> _zz_904);
  assign _zz_12323 = _zz_12324;
  assign _zz_12324 = ($signed(_zz_12326) - $signed(_zz_901));
  assign _zz_12325 = ({8'd0,data_mid_104_real} <<< 8);
  assign _zz_12326 = {{8{_zz_12325[23]}}, _zz_12325};
  assign _zz_12327 = fixTo_1082_dout;
  assign _zz_12328 = _zz_12329[31 : 0];
  assign _zz_12329 = _zz_12330;
  assign _zz_12330 = ($signed(_zz_12331) >>> _zz_904);
  assign _zz_12331 = _zz_12332;
  assign _zz_12332 = ($signed(_zz_12334) - $signed(_zz_902));
  assign _zz_12333 = ({8'd0,data_mid_104_imag} <<< 8);
  assign _zz_12334 = {{8{_zz_12333[23]}}, _zz_12333};
  assign _zz_12335 = fixTo_1083_dout;
  assign _zz_12336 = _zz_12337[31 : 0];
  assign _zz_12337 = _zz_12338;
  assign _zz_12338 = ($signed(_zz_12339) >>> _zz_905);
  assign _zz_12339 = _zz_12340;
  assign _zz_12340 = ($signed(_zz_12342) + $signed(_zz_901));
  assign _zz_12341 = ({8'd0,data_mid_104_real} <<< 8);
  assign _zz_12342 = {{8{_zz_12341[23]}}, _zz_12341};
  assign _zz_12343 = fixTo_1084_dout;
  assign _zz_12344 = _zz_12345[31 : 0];
  assign _zz_12345 = _zz_12346;
  assign _zz_12346 = ($signed(_zz_12347) >>> _zz_905);
  assign _zz_12347 = _zz_12348;
  assign _zz_12348 = ($signed(_zz_12350) + $signed(_zz_902));
  assign _zz_12349 = ({8'd0,data_mid_104_imag} <<< 8);
  assign _zz_12350 = {{8{_zz_12349[23]}}, _zz_12349};
  assign _zz_12351 = fixTo_1085_dout;
  assign _zz_12352 = ($signed(twiddle_factor_table_4_real) + $signed(twiddle_factor_table_4_imag));
  assign _zz_12353 = ($signed(_zz_908) - $signed(_zz_12354));
  assign _zz_12354 = ($signed(_zz_12355) * $signed(twiddle_factor_table_4_imag));
  assign _zz_12355 = ($signed(data_mid_109_real) + $signed(data_mid_109_imag));
  assign _zz_12356 = fixTo_1086_dout;
  assign _zz_12357 = ($signed(_zz_908) + $signed(_zz_12358));
  assign _zz_12358 = ($signed(_zz_12359) * $signed(twiddle_factor_table_4_real));
  assign _zz_12359 = ($signed(data_mid_109_imag) - $signed(data_mid_109_real));
  assign _zz_12360 = fixTo_1087_dout;
  assign _zz_12361 = _zz_12362[31 : 0];
  assign _zz_12362 = _zz_12363;
  assign _zz_12363 = ($signed(_zz_12364) >>> _zz_909);
  assign _zz_12364 = _zz_12365;
  assign _zz_12365 = ($signed(_zz_12367) - $signed(_zz_906));
  assign _zz_12366 = ({8'd0,data_mid_105_real} <<< 8);
  assign _zz_12367 = {{8{_zz_12366[23]}}, _zz_12366};
  assign _zz_12368 = fixTo_1088_dout;
  assign _zz_12369 = _zz_12370[31 : 0];
  assign _zz_12370 = _zz_12371;
  assign _zz_12371 = ($signed(_zz_12372) >>> _zz_909);
  assign _zz_12372 = _zz_12373;
  assign _zz_12373 = ($signed(_zz_12375) - $signed(_zz_907));
  assign _zz_12374 = ({8'd0,data_mid_105_imag} <<< 8);
  assign _zz_12375 = {{8{_zz_12374[23]}}, _zz_12374};
  assign _zz_12376 = fixTo_1089_dout;
  assign _zz_12377 = _zz_12378[31 : 0];
  assign _zz_12378 = _zz_12379;
  assign _zz_12379 = ($signed(_zz_12380) >>> _zz_910);
  assign _zz_12380 = _zz_12381;
  assign _zz_12381 = ($signed(_zz_12383) + $signed(_zz_906));
  assign _zz_12382 = ({8'd0,data_mid_105_real} <<< 8);
  assign _zz_12383 = {{8{_zz_12382[23]}}, _zz_12382};
  assign _zz_12384 = fixTo_1090_dout;
  assign _zz_12385 = _zz_12386[31 : 0];
  assign _zz_12386 = _zz_12387;
  assign _zz_12387 = ($signed(_zz_12388) >>> _zz_910);
  assign _zz_12388 = _zz_12389;
  assign _zz_12389 = ($signed(_zz_12391) + $signed(_zz_907));
  assign _zz_12390 = ({8'd0,data_mid_105_imag} <<< 8);
  assign _zz_12391 = {{8{_zz_12390[23]}}, _zz_12390};
  assign _zz_12392 = fixTo_1091_dout;
  assign _zz_12393 = ($signed(twiddle_factor_table_5_real) + $signed(twiddle_factor_table_5_imag));
  assign _zz_12394 = ($signed(_zz_913) - $signed(_zz_12395));
  assign _zz_12395 = ($signed(_zz_12396) * $signed(twiddle_factor_table_5_imag));
  assign _zz_12396 = ($signed(data_mid_110_real) + $signed(data_mid_110_imag));
  assign _zz_12397 = fixTo_1092_dout;
  assign _zz_12398 = ($signed(_zz_913) + $signed(_zz_12399));
  assign _zz_12399 = ($signed(_zz_12400) * $signed(twiddle_factor_table_5_real));
  assign _zz_12400 = ($signed(data_mid_110_imag) - $signed(data_mid_110_real));
  assign _zz_12401 = fixTo_1093_dout;
  assign _zz_12402 = _zz_12403[31 : 0];
  assign _zz_12403 = _zz_12404;
  assign _zz_12404 = ($signed(_zz_12405) >>> _zz_914);
  assign _zz_12405 = _zz_12406;
  assign _zz_12406 = ($signed(_zz_12408) - $signed(_zz_911));
  assign _zz_12407 = ({8'd0,data_mid_106_real} <<< 8);
  assign _zz_12408 = {{8{_zz_12407[23]}}, _zz_12407};
  assign _zz_12409 = fixTo_1094_dout;
  assign _zz_12410 = _zz_12411[31 : 0];
  assign _zz_12411 = _zz_12412;
  assign _zz_12412 = ($signed(_zz_12413) >>> _zz_914);
  assign _zz_12413 = _zz_12414;
  assign _zz_12414 = ($signed(_zz_12416) - $signed(_zz_912));
  assign _zz_12415 = ({8'd0,data_mid_106_imag} <<< 8);
  assign _zz_12416 = {{8{_zz_12415[23]}}, _zz_12415};
  assign _zz_12417 = fixTo_1095_dout;
  assign _zz_12418 = _zz_12419[31 : 0];
  assign _zz_12419 = _zz_12420;
  assign _zz_12420 = ($signed(_zz_12421) >>> _zz_915);
  assign _zz_12421 = _zz_12422;
  assign _zz_12422 = ($signed(_zz_12424) + $signed(_zz_911));
  assign _zz_12423 = ({8'd0,data_mid_106_real} <<< 8);
  assign _zz_12424 = {{8{_zz_12423[23]}}, _zz_12423};
  assign _zz_12425 = fixTo_1096_dout;
  assign _zz_12426 = _zz_12427[31 : 0];
  assign _zz_12427 = _zz_12428;
  assign _zz_12428 = ($signed(_zz_12429) >>> _zz_915);
  assign _zz_12429 = _zz_12430;
  assign _zz_12430 = ($signed(_zz_12432) + $signed(_zz_912));
  assign _zz_12431 = ({8'd0,data_mid_106_imag} <<< 8);
  assign _zz_12432 = {{8{_zz_12431[23]}}, _zz_12431};
  assign _zz_12433 = fixTo_1097_dout;
  assign _zz_12434 = ($signed(twiddle_factor_table_6_real) + $signed(twiddle_factor_table_6_imag));
  assign _zz_12435 = ($signed(_zz_918) - $signed(_zz_12436));
  assign _zz_12436 = ($signed(_zz_12437) * $signed(twiddle_factor_table_6_imag));
  assign _zz_12437 = ($signed(data_mid_111_real) + $signed(data_mid_111_imag));
  assign _zz_12438 = fixTo_1098_dout;
  assign _zz_12439 = ($signed(_zz_918) + $signed(_zz_12440));
  assign _zz_12440 = ($signed(_zz_12441) * $signed(twiddle_factor_table_6_real));
  assign _zz_12441 = ($signed(data_mid_111_imag) - $signed(data_mid_111_real));
  assign _zz_12442 = fixTo_1099_dout;
  assign _zz_12443 = _zz_12444[31 : 0];
  assign _zz_12444 = _zz_12445;
  assign _zz_12445 = ($signed(_zz_12446) >>> _zz_919);
  assign _zz_12446 = _zz_12447;
  assign _zz_12447 = ($signed(_zz_12449) - $signed(_zz_916));
  assign _zz_12448 = ({8'd0,data_mid_107_real} <<< 8);
  assign _zz_12449 = {{8{_zz_12448[23]}}, _zz_12448};
  assign _zz_12450 = fixTo_1100_dout;
  assign _zz_12451 = _zz_12452[31 : 0];
  assign _zz_12452 = _zz_12453;
  assign _zz_12453 = ($signed(_zz_12454) >>> _zz_919);
  assign _zz_12454 = _zz_12455;
  assign _zz_12455 = ($signed(_zz_12457) - $signed(_zz_917));
  assign _zz_12456 = ({8'd0,data_mid_107_imag} <<< 8);
  assign _zz_12457 = {{8{_zz_12456[23]}}, _zz_12456};
  assign _zz_12458 = fixTo_1101_dout;
  assign _zz_12459 = _zz_12460[31 : 0];
  assign _zz_12460 = _zz_12461;
  assign _zz_12461 = ($signed(_zz_12462) >>> _zz_920);
  assign _zz_12462 = _zz_12463;
  assign _zz_12463 = ($signed(_zz_12465) + $signed(_zz_916));
  assign _zz_12464 = ({8'd0,data_mid_107_real} <<< 8);
  assign _zz_12465 = {{8{_zz_12464[23]}}, _zz_12464};
  assign _zz_12466 = fixTo_1102_dout;
  assign _zz_12467 = _zz_12468[31 : 0];
  assign _zz_12468 = _zz_12469;
  assign _zz_12469 = ($signed(_zz_12470) >>> _zz_920);
  assign _zz_12470 = _zz_12471;
  assign _zz_12471 = ($signed(_zz_12473) + $signed(_zz_917));
  assign _zz_12472 = ({8'd0,data_mid_107_imag} <<< 8);
  assign _zz_12473 = {{8{_zz_12472[23]}}, _zz_12472};
  assign _zz_12474 = fixTo_1103_dout;
  assign _zz_12475 = ($signed(twiddle_factor_table_3_real) + $signed(twiddle_factor_table_3_imag));
  assign _zz_12476 = ($signed(_zz_923) - $signed(_zz_12477));
  assign _zz_12477 = ($signed(_zz_12478) * $signed(twiddle_factor_table_3_imag));
  assign _zz_12478 = ($signed(data_mid_116_real) + $signed(data_mid_116_imag));
  assign _zz_12479 = fixTo_1104_dout;
  assign _zz_12480 = ($signed(_zz_923) + $signed(_zz_12481));
  assign _zz_12481 = ($signed(_zz_12482) * $signed(twiddle_factor_table_3_real));
  assign _zz_12482 = ($signed(data_mid_116_imag) - $signed(data_mid_116_real));
  assign _zz_12483 = fixTo_1105_dout;
  assign _zz_12484 = _zz_12485[31 : 0];
  assign _zz_12485 = _zz_12486;
  assign _zz_12486 = ($signed(_zz_12487) >>> _zz_924);
  assign _zz_12487 = _zz_12488;
  assign _zz_12488 = ($signed(_zz_12490) - $signed(_zz_921));
  assign _zz_12489 = ({8'd0,data_mid_112_real} <<< 8);
  assign _zz_12490 = {{8{_zz_12489[23]}}, _zz_12489};
  assign _zz_12491 = fixTo_1106_dout;
  assign _zz_12492 = _zz_12493[31 : 0];
  assign _zz_12493 = _zz_12494;
  assign _zz_12494 = ($signed(_zz_12495) >>> _zz_924);
  assign _zz_12495 = _zz_12496;
  assign _zz_12496 = ($signed(_zz_12498) - $signed(_zz_922));
  assign _zz_12497 = ({8'd0,data_mid_112_imag} <<< 8);
  assign _zz_12498 = {{8{_zz_12497[23]}}, _zz_12497};
  assign _zz_12499 = fixTo_1107_dout;
  assign _zz_12500 = _zz_12501[31 : 0];
  assign _zz_12501 = _zz_12502;
  assign _zz_12502 = ($signed(_zz_12503) >>> _zz_925);
  assign _zz_12503 = _zz_12504;
  assign _zz_12504 = ($signed(_zz_12506) + $signed(_zz_921));
  assign _zz_12505 = ({8'd0,data_mid_112_real} <<< 8);
  assign _zz_12506 = {{8{_zz_12505[23]}}, _zz_12505};
  assign _zz_12507 = fixTo_1108_dout;
  assign _zz_12508 = _zz_12509[31 : 0];
  assign _zz_12509 = _zz_12510;
  assign _zz_12510 = ($signed(_zz_12511) >>> _zz_925);
  assign _zz_12511 = _zz_12512;
  assign _zz_12512 = ($signed(_zz_12514) + $signed(_zz_922));
  assign _zz_12513 = ({8'd0,data_mid_112_imag} <<< 8);
  assign _zz_12514 = {{8{_zz_12513[23]}}, _zz_12513};
  assign _zz_12515 = fixTo_1109_dout;
  assign _zz_12516 = ($signed(twiddle_factor_table_4_real) + $signed(twiddle_factor_table_4_imag));
  assign _zz_12517 = ($signed(_zz_928) - $signed(_zz_12518));
  assign _zz_12518 = ($signed(_zz_12519) * $signed(twiddle_factor_table_4_imag));
  assign _zz_12519 = ($signed(data_mid_117_real) + $signed(data_mid_117_imag));
  assign _zz_12520 = fixTo_1110_dout;
  assign _zz_12521 = ($signed(_zz_928) + $signed(_zz_12522));
  assign _zz_12522 = ($signed(_zz_12523) * $signed(twiddle_factor_table_4_real));
  assign _zz_12523 = ($signed(data_mid_117_imag) - $signed(data_mid_117_real));
  assign _zz_12524 = fixTo_1111_dout;
  assign _zz_12525 = _zz_12526[31 : 0];
  assign _zz_12526 = _zz_12527;
  assign _zz_12527 = ($signed(_zz_12528) >>> _zz_929);
  assign _zz_12528 = _zz_12529;
  assign _zz_12529 = ($signed(_zz_12531) - $signed(_zz_926));
  assign _zz_12530 = ({8'd0,data_mid_113_real} <<< 8);
  assign _zz_12531 = {{8{_zz_12530[23]}}, _zz_12530};
  assign _zz_12532 = fixTo_1112_dout;
  assign _zz_12533 = _zz_12534[31 : 0];
  assign _zz_12534 = _zz_12535;
  assign _zz_12535 = ($signed(_zz_12536) >>> _zz_929);
  assign _zz_12536 = _zz_12537;
  assign _zz_12537 = ($signed(_zz_12539) - $signed(_zz_927));
  assign _zz_12538 = ({8'd0,data_mid_113_imag} <<< 8);
  assign _zz_12539 = {{8{_zz_12538[23]}}, _zz_12538};
  assign _zz_12540 = fixTo_1113_dout;
  assign _zz_12541 = _zz_12542[31 : 0];
  assign _zz_12542 = _zz_12543;
  assign _zz_12543 = ($signed(_zz_12544) >>> _zz_930);
  assign _zz_12544 = _zz_12545;
  assign _zz_12545 = ($signed(_zz_12547) + $signed(_zz_926));
  assign _zz_12546 = ({8'd0,data_mid_113_real} <<< 8);
  assign _zz_12547 = {{8{_zz_12546[23]}}, _zz_12546};
  assign _zz_12548 = fixTo_1114_dout;
  assign _zz_12549 = _zz_12550[31 : 0];
  assign _zz_12550 = _zz_12551;
  assign _zz_12551 = ($signed(_zz_12552) >>> _zz_930);
  assign _zz_12552 = _zz_12553;
  assign _zz_12553 = ($signed(_zz_12555) + $signed(_zz_927));
  assign _zz_12554 = ({8'd0,data_mid_113_imag} <<< 8);
  assign _zz_12555 = {{8{_zz_12554[23]}}, _zz_12554};
  assign _zz_12556 = fixTo_1115_dout;
  assign _zz_12557 = ($signed(twiddle_factor_table_5_real) + $signed(twiddle_factor_table_5_imag));
  assign _zz_12558 = ($signed(_zz_933) - $signed(_zz_12559));
  assign _zz_12559 = ($signed(_zz_12560) * $signed(twiddle_factor_table_5_imag));
  assign _zz_12560 = ($signed(data_mid_118_real) + $signed(data_mid_118_imag));
  assign _zz_12561 = fixTo_1116_dout;
  assign _zz_12562 = ($signed(_zz_933) + $signed(_zz_12563));
  assign _zz_12563 = ($signed(_zz_12564) * $signed(twiddle_factor_table_5_real));
  assign _zz_12564 = ($signed(data_mid_118_imag) - $signed(data_mid_118_real));
  assign _zz_12565 = fixTo_1117_dout;
  assign _zz_12566 = _zz_12567[31 : 0];
  assign _zz_12567 = _zz_12568;
  assign _zz_12568 = ($signed(_zz_12569) >>> _zz_934);
  assign _zz_12569 = _zz_12570;
  assign _zz_12570 = ($signed(_zz_12572) - $signed(_zz_931));
  assign _zz_12571 = ({8'd0,data_mid_114_real} <<< 8);
  assign _zz_12572 = {{8{_zz_12571[23]}}, _zz_12571};
  assign _zz_12573 = fixTo_1118_dout;
  assign _zz_12574 = _zz_12575[31 : 0];
  assign _zz_12575 = _zz_12576;
  assign _zz_12576 = ($signed(_zz_12577) >>> _zz_934);
  assign _zz_12577 = _zz_12578;
  assign _zz_12578 = ($signed(_zz_12580) - $signed(_zz_932));
  assign _zz_12579 = ({8'd0,data_mid_114_imag} <<< 8);
  assign _zz_12580 = {{8{_zz_12579[23]}}, _zz_12579};
  assign _zz_12581 = fixTo_1119_dout;
  assign _zz_12582 = _zz_12583[31 : 0];
  assign _zz_12583 = _zz_12584;
  assign _zz_12584 = ($signed(_zz_12585) >>> _zz_935);
  assign _zz_12585 = _zz_12586;
  assign _zz_12586 = ($signed(_zz_12588) + $signed(_zz_931));
  assign _zz_12587 = ({8'd0,data_mid_114_real} <<< 8);
  assign _zz_12588 = {{8{_zz_12587[23]}}, _zz_12587};
  assign _zz_12589 = fixTo_1120_dout;
  assign _zz_12590 = _zz_12591[31 : 0];
  assign _zz_12591 = _zz_12592;
  assign _zz_12592 = ($signed(_zz_12593) >>> _zz_935);
  assign _zz_12593 = _zz_12594;
  assign _zz_12594 = ($signed(_zz_12596) + $signed(_zz_932));
  assign _zz_12595 = ({8'd0,data_mid_114_imag} <<< 8);
  assign _zz_12596 = {{8{_zz_12595[23]}}, _zz_12595};
  assign _zz_12597 = fixTo_1121_dout;
  assign _zz_12598 = ($signed(twiddle_factor_table_6_real) + $signed(twiddle_factor_table_6_imag));
  assign _zz_12599 = ($signed(_zz_938) - $signed(_zz_12600));
  assign _zz_12600 = ($signed(_zz_12601) * $signed(twiddle_factor_table_6_imag));
  assign _zz_12601 = ($signed(data_mid_119_real) + $signed(data_mid_119_imag));
  assign _zz_12602 = fixTo_1122_dout;
  assign _zz_12603 = ($signed(_zz_938) + $signed(_zz_12604));
  assign _zz_12604 = ($signed(_zz_12605) * $signed(twiddle_factor_table_6_real));
  assign _zz_12605 = ($signed(data_mid_119_imag) - $signed(data_mid_119_real));
  assign _zz_12606 = fixTo_1123_dout;
  assign _zz_12607 = _zz_12608[31 : 0];
  assign _zz_12608 = _zz_12609;
  assign _zz_12609 = ($signed(_zz_12610) >>> _zz_939);
  assign _zz_12610 = _zz_12611;
  assign _zz_12611 = ($signed(_zz_12613) - $signed(_zz_936));
  assign _zz_12612 = ({8'd0,data_mid_115_real} <<< 8);
  assign _zz_12613 = {{8{_zz_12612[23]}}, _zz_12612};
  assign _zz_12614 = fixTo_1124_dout;
  assign _zz_12615 = _zz_12616[31 : 0];
  assign _zz_12616 = _zz_12617;
  assign _zz_12617 = ($signed(_zz_12618) >>> _zz_939);
  assign _zz_12618 = _zz_12619;
  assign _zz_12619 = ($signed(_zz_12621) - $signed(_zz_937));
  assign _zz_12620 = ({8'd0,data_mid_115_imag} <<< 8);
  assign _zz_12621 = {{8{_zz_12620[23]}}, _zz_12620};
  assign _zz_12622 = fixTo_1125_dout;
  assign _zz_12623 = _zz_12624[31 : 0];
  assign _zz_12624 = _zz_12625;
  assign _zz_12625 = ($signed(_zz_12626) >>> _zz_940);
  assign _zz_12626 = _zz_12627;
  assign _zz_12627 = ($signed(_zz_12629) + $signed(_zz_936));
  assign _zz_12628 = ({8'd0,data_mid_115_real} <<< 8);
  assign _zz_12629 = {{8{_zz_12628[23]}}, _zz_12628};
  assign _zz_12630 = fixTo_1126_dout;
  assign _zz_12631 = _zz_12632[31 : 0];
  assign _zz_12632 = _zz_12633;
  assign _zz_12633 = ($signed(_zz_12634) >>> _zz_940);
  assign _zz_12634 = _zz_12635;
  assign _zz_12635 = ($signed(_zz_12637) + $signed(_zz_937));
  assign _zz_12636 = ({8'd0,data_mid_115_imag} <<< 8);
  assign _zz_12637 = {{8{_zz_12636[23]}}, _zz_12636};
  assign _zz_12638 = fixTo_1127_dout;
  assign _zz_12639 = ($signed(twiddle_factor_table_3_real) + $signed(twiddle_factor_table_3_imag));
  assign _zz_12640 = ($signed(_zz_943) - $signed(_zz_12641));
  assign _zz_12641 = ($signed(_zz_12642) * $signed(twiddle_factor_table_3_imag));
  assign _zz_12642 = ($signed(data_mid_124_real) + $signed(data_mid_124_imag));
  assign _zz_12643 = fixTo_1128_dout;
  assign _zz_12644 = ($signed(_zz_943) + $signed(_zz_12645));
  assign _zz_12645 = ($signed(_zz_12646) * $signed(twiddle_factor_table_3_real));
  assign _zz_12646 = ($signed(data_mid_124_imag) - $signed(data_mid_124_real));
  assign _zz_12647 = fixTo_1129_dout;
  assign _zz_12648 = _zz_12649[31 : 0];
  assign _zz_12649 = _zz_12650;
  assign _zz_12650 = ($signed(_zz_12651) >>> _zz_944);
  assign _zz_12651 = _zz_12652;
  assign _zz_12652 = ($signed(_zz_12654) - $signed(_zz_941));
  assign _zz_12653 = ({8'd0,data_mid_120_real} <<< 8);
  assign _zz_12654 = {{8{_zz_12653[23]}}, _zz_12653};
  assign _zz_12655 = fixTo_1130_dout;
  assign _zz_12656 = _zz_12657[31 : 0];
  assign _zz_12657 = _zz_12658;
  assign _zz_12658 = ($signed(_zz_12659) >>> _zz_944);
  assign _zz_12659 = _zz_12660;
  assign _zz_12660 = ($signed(_zz_12662) - $signed(_zz_942));
  assign _zz_12661 = ({8'd0,data_mid_120_imag} <<< 8);
  assign _zz_12662 = {{8{_zz_12661[23]}}, _zz_12661};
  assign _zz_12663 = fixTo_1131_dout;
  assign _zz_12664 = _zz_12665[31 : 0];
  assign _zz_12665 = _zz_12666;
  assign _zz_12666 = ($signed(_zz_12667) >>> _zz_945);
  assign _zz_12667 = _zz_12668;
  assign _zz_12668 = ($signed(_zz_12670) + $signed(_zz_941));
  assign _zz_12669 = ({8'd0,data_mid_120_real} <<< 8);
  assign _zz_12670 = {{8{_zz_12669[23]}}, _zz_12669};
  assign _zz_12671 = fixTo_1132_dout;
  assign _zz_12672 = _zz_12673[31 : 0];
  assign _zz_12673 = _zz_12674;
  assign _zz_12674 = ($signed(_zz_12675) >>> _zz_945);
  assign _zz_12675 = _zz_12676;
  assign _zz_12676 = ($signed(_zz_12678) + $signed(_zz_942));
  assign _zz_12677 = ({8'd0,data_mid_120_imag} <<< 8);
  assign _zz_12678 = {{8{_zz_12677[23]}}, _zz_12677};
  assign _zz_12679 = fixTo_1133_dout;
  assign _zz_12680 = ($signed(twiddle_factor_table_4_real) + $signed(twiddle_factor_table_4_imag));
  assign _zz_12681 = ($signed(_zz_948) - $signed(_zz_12682));
  assign _zz_12682 = ($signed(_zz_12683) * $signed(twiddle_factor_table_4_imag));
  assign _zz_12683 = ($signed(data_mid_125_real) + $signed(data_mid_125_imag));
  assign _zz_12684 = fixTo_1134_dout;
  assign _zz_12685 = ($signed(_zz_948) + $signed(_zz_12686));
  assign _zz_12686 = ($signed(_zz_12687) * $signed(twiddle_factor_table_4_real));
  assign _zz_12687 = ($signed(data_mid_125_imag) - $signed(data_mid_125_real));
  assign _zz_12688 = fixTo_1135_dout;
  assign _zz_12689 = _zz_12690[31 : 0];
  assign _zz_12690 = _zz_12691;
  assign _zz_12691 = ($signed(_zz_12692) >>> _zz_949);
  assign _zz_12692 = _zz_12693;
  assign _zz_12693 = ($signed(_zz_12695) - $signed(_zz_946));
  assign _zz_12694 = ({8'd0,data_mid_121_real} <<< 8);
  assign _zz_12695 = {{8{_zz_12694[23]}}, _zz_12694};
  assign _zz_12696 = fixTo_1136_dout;
  assign _zz_12697 = _zz_12698[31 : 0];
  assign _zz_12698 = _zz_12699;
  assign _zz_12699 = ($signed(_zz_12700) >>> _zz_949);
  assign _zz_12700 = _zz_12701;
  assign _zz_12701 = ($signed(_zz_12703) - $signed(_zz_947));
  assign _zz_12702 = ({8'd0,data_mid_121_imag} <<< 8);
  assign _zz_12703 = {{8{_zz_12702[23]}}, _zz_12702};
  assign _zz_12704 = fixTo_1137_dout;
  assign _zz_12705 = _zz_12706[31 : 0];
  assign _zz_12706 = _zz_12707;
  assign _zz_12707 = ($signed(_zz_12708) >>> _zz_950);
  assign _zz_12708 = _zz_12709;
  assign _zz_12709 = ($signed(_zz_12711) + $signed(_zz_946));
  assign _zz_12710 = ({8'd0,data_mid_121_real} <<< 8);
  assign _zz_12711 = {{8{_zz_12710[23]}}, _zz_12710};
  assign _zz_12712 = fixTo_1138_dout;
  assign _zz_12713 = _zz_12714[31 : 0];
  assign _zz_12714 = _zz_12715;
  assign _zz_12715 = ($signed(_zz_12716) >>> _zz_950);
  assign _zz_12716 = _zz_12717;
  assign _zz_12717 = ($signed(_zz_12719) + $signed(_zz_947));
  assign _zz_12718 = ({8'd0,data_mid_121_imag} <<< 8);
  assign _zz_12719 = {{8{_zz_12718[23]}}, _zz_12718};
  assign _zz_12720 = fixTo_1139_dout;
  assign _zz_12721 = ($signed(twiddle_factor_table_5_real) + $signed(twiddle_factor_table_5_imag));
  assign _zz_12722 = ($signed(_zz_953) - $signed(_zz_12723));
  assign _zz_12723 = ($signed(_zz_12724) * $signed(twiddle_factor_table_5_imag));
  assign _zz_12724 = ($signed(data_mid_126_real) + $signed(data_mid_126_imag));
  assign _zz_12725 = fixTo_1140_dout;
  assign _zz_12726 = ($signed(_zz_953) + $signed(_zz_12727));
  assign _zz_12727 = ($signed(_zz_12728) * $signed(twiddle_factor_table_5_real));
  assign _zz_12728 = ($signed(data_mid_126_imag) - $signed(data_mid_126_real));
  assign _zz_12729 = fixTo_1141_dout;
  assign _zz_12730 = _zz_12731[31 : 0];
  assign _zz_12731 = _zz_12732;
  assign _zz_12732 = ($signed(_zz_12733) >>> _zz_954);
  assign _zz_12733 = _zz_12734;
  assign _zz_12734 = ($signed(_zz_12736) - $signed(_zz_951));
  assign _zz_12735 = ({8'd0,data_mid_122_real} <<< 8);
  assign _zz_12736 = {{8{_zz_12735[23]}}, _zz_12735};
  assign _zz_12737 = fixTo_1142_dout;
  assign _zz_12738 = _zz_12739[31 : 0];
  assign _zz_12739 = _zz_12740;
  assign _zz_12740 = ($signed(_zz_12741) >>> _zz_954);
  assign _zz_12741 = _zz_12742;
  assign _zz_12742 = ($signed(_zz_12744) - $signed(_zz_952));
  assign _zz_12743 = ({8'd0,data_mid_122_imag} <<< 8);
  assign _zz_12744 = {{8{_zz_12743[23]}}, _zz_12743};
  assign _zz_12745 = fixTo_1143_dout;
  assign _zz_12746 = _zz_12747[31 : 0];
  assign _zz_12747 = _zz_12748;
  assign _zz_12748 = ($signed(_zz_12749) >>> _zz_955);
  assign _zz_12749 = _zz_12750;
  assign _zz_12750 = ($signed(_zz_12752) + $signed(_zz_951));
  assign _zz_12751 = ({8'd0,data_mid_122_real} <<< 8);
  assign _zz_12752 = {{8{_zz_12751[23]}}, _zz_12751};
  assign _zz_12753 = fixTo_1144_dout;
  assign _zz_12754 = _zz_12755[31 : 0];
  assign _zz_12755 = _zz_12756;
  assign _zz_12756 = ($signed(_zz_12757) >>> _zz_955);
  assign _zz_12757 = _zz_12758;
  assign _zz_12758 = ($signed(_zz_12760) + $signed(_zz_952));
  assign _zz_12759 = ({8'd0,data_mid_122_imag} <<< 8);
  assign _zz_12760 = {{8{_zz_12759[23]}}, _zz_12759};
  assign _zz_12761 = fixTo_1145_dout;
  assign _zz_12762 = ($signed(twiddle_factor_table_6_real) + $signed(twiddle_factor_table_6_imag));
  assign _zz_12763 = ($signed(_zz_958) - $signed(_zz_12764));
  assign _zz_12764 = ($signed(_zz_12765) * $signed(twiddle_factor_table_6_imag));
  assign _zz_12765 = ($signed(data_mid_127_real) + $signed(data_mid_127_imag));
  assign _zz_12766 = fixTo_1146_dout;
  assign _zz_12767 = ($signed(_zz_958) + $signed(_zz_12768));
  assign _zz_12768 = ($signed(_zz_12769) * $signed(twiddle_factor_table_6_real));
  assign _zz_12769 = ($signed(data_mid_127_imag) - $signed(data_mid_127_real));
  assign _zz_12770 = fixTo_1147_dout;
  assign _zz_12771 = _zz_12772[31 : 0];
  assign _zz_12772 = _zz_12773;
  assign _zz_12773 = ($signed(_zz_12774) >>> _zz_959);
  assign _zz_12774 = _zz_12775;
  assign _zz_12775 = ($signed(_zz_12777) - $signed(_zz_956));
  assign _zz_12776 = ({8'd0,data_mid_123_real} <<< 8);
  assign _zz_12777 = {{8{_zz_12776[23]}}, _zz_12776};
  assign _zz_12778 = fixTo_1148_dout;
  assign _zz_12779 = _zz_12780[31 : 0];
  assign _zz_12780 = _zz_12781;
  assign _zz_12781 = ($signed(_zz_12782) >>> _zz_959);
  assign _zz_12782 = _zz_12783;
  assign _zz_12783 = ($signed(_zz_12785) - $signed(_zz_957));
  assign _zz_12784 = ({8'd0,data_mid_123_imag} <<< 8);
  assign _zz_12785 = {{8{_zz_12784[23]}}, _zz_12784};
  assign _zz_12786 = fixTo_1149_dout;
  assign _zz_12787 = _zz_12788[31 : 0];
  assign _zz_12788 = _zz_12789;
  assign _zz_12789 = ($signed(_zz_12790) >>> _zz_960);
  assign _zz_12790 = _zz_12791;
  assign _zz_12791 = ($signed(_zz_12793) + $signed(_zz_956));
  assign _zz_12792 = ({8'd0,data_mid_123_real} <<< 8);
  assign _zz_12793 = {{8{_zz_12792[23]}}, _zz_12792};
  assign _zz_12794 = fixTo_1150_dout;
  assign _zz_12795 = _zz_12796[31 : 0];
  assign _zz_12796 = _zz_12797;
  assign _zz_12797 = ($signed(_zz_12798) >>> _zz_960);
  assign _zz_12798 = _zz_12799;
  assign _zz_12799 = ($signed(_zz_12801) + $signed(_zz_957));
  assign _zz_12800 = ({8'd0,data_mid_123_imag} <<< 8);
  assign _zz_12801 = {{8{_zz_12800[23]}}, _zz_12800};
  assign _zz_12802 = fixTo_1151_dout;
  assign _zz_12803 = ($signed(twiddle_factor_table_7_real) + $signed(twiddle_factor_table_7_imag));
  assign _zz_12804 = ($signed(_zz_963) - $signed(_zz_12805));
  assign _zz_12805 = ($signed(_zz_12806) * $signed(twiddle_factor_table_7_imag));
  assign _zz_12806 = ($signed(data_mid_8_real) + $signed(data_mid_8_imag));
  assign _zz_12807 = fixTo_1152_dout;
  assign _zz_12808 = ($signed(_zz_963) + $signed(_zz_12809));
  assign _zz_12809 = ($signed(_zz_12810) * $signed(twiddle_factor_table_7_real));
  assign _zz_12810 = ($signed(data_mid_8_imag) - $signed(data_mid_8_real));
  assign _zz_12811 = fixTo_1153_dout;
  assign _zz_12812 = _zz_12813[31 : 0];
  assign _zz_12813 = _zz_12814;
  assign _zz_12814 = ($signed(_zz_12815) >>> _zz_964);
  assign _zz_12815 = _zz_12816;
  assign _zz_12816 = ($signed(_zz_12818) - $signed(_zz_961));
  assign _zz_12817 = ({8'd0,data_mid_0_real} <<< 8);
  assign _zz_12818 = {{8{_zz_12817[23]}}, _zz_12817};
  assign _zz_12819 = fixTo_1154_dout;
  assign _zz_12820 = _zz_12821[31 : 0];
  assign _zz_12821 = _zz_12822;
  assign _zz_12822 = ($signed(_zz_12823) >>> _zz_964);
  assign _zz_12823 = _zz_12824;
  assign _zz_12824 = ($signed(_zz_12826) - $signed(_zz_962));
  assign _zz_12825 = ({8'd0,data_mid_0_imag} <<< 8);
  assign _zz_12826 = {{8{_zz_12825[23]}}, _zz_12825};
  assign _zz_12827 = fixTo_1155_dout;
  assign _zz_12828 = _zz_12829[31 : 0];
  assign _zz_12829 = _zz_12830;
  assign _zz_12830 = ($signed(_zz_12831) >>> _zz_965);
  assign _zz_12831 = _zz_12832;
  assign _zz_12832 = ($signed(_zz_12834) + $signed(_zz_961));
  assign _zz_12833 = ({8'd0,data_mid_0_real} <<< 8);
  assign _zz_12834 = {{8{_zz_12833[23]}}, _zz_12833};
  assign _zz_12835 = fixTo_1156_dout;
  assign _zz_12836 = _zz_12837[31 : 0];
  assign _zz_12837 = _zz_12838;
  assign _zz_12838 = ($signed(_zz_12839) >>> _zz_965);
  assign _zz_12839 = _zz_12840;
  assign _zz_12840 = ($signed(_zz_12842) + $signed(_zz_962));
  assign _zz_12841 = ({8'd0,data_mid_0_imag} <<< 8);
  assign _zz_12842 = {{8{_zz_12841[23]}}, _zz_12841};
  assign _zz_12843 = fixTo_1157_dout;
  assign _zz_12844 = ($signed(twiddle_factor_table_8_real) + $signed(twiddle_factor_table_8_imag));
  assign _zz_12845 = ($signed(_zz_968) - $signed(_zz_12846));
  assign _zz_12846 = ($signed(_zz_12847) * $signed(twiddle_factor_table_8_imag));
  assign _zz_12847 = ($signed(data_mid_9_real) + $signed(data_mid_9_imag));
  assign _zz_12848 = fixTo_1158_dout;
  assign _zz_12849 = ($signed(_zz_968) + $signed(_zz_12850));
  assign _zz_12850 = ($signed(_zz_12851) * $signed(twiddle_factor_table_8_real));
  assign _zz_12851 = ($signed(data_mid_9_imag) - $signed(data_mid_9_real));
  assign _zz_12852 = fixTo_1159_dout;
  assign _zz_12853 = _zz_12854[31 : 0];
  assign _zz_12854 = _zz_12855;
  assign _zz_12855 = ($signed(_zz_12856) >>> _zz_969);
  assign _zz_12856 = _zz_12857;
  assign _zz_12857 = ($signed(_zz_12859) - $signed(_zz_966));
  assign _zz_12858 = ({8'd0,data_mid_1_real} <<< 8);
  assign _zz_12859 = {{8{_zz_12858[23]}}, _zz_12858};
  assign _zz_12860 = fixTo_1160_dout;
  assign _zz_12861 = _zz_12862[31 : 0];
  assign _zz_12862 = _zz_12863;
  assign _zz_12863 = ($signed(_zz_12864) >>> _zz_969);
  assign _zz_12864 = _zz_12865;
  assign _zz_12865 = ($signed(_zz_12867) - $signed(_zz_967));
  assign _zz_12866 = ({8'd0,data_mid_1_imag} <<< 8);
  assign _zz_12867 = {{8{_zz_12866[23]}}, _zz_12866};
  assign _zz_12868 = fixTo_1161_dout;
  assign _zz_12869 = _zz_12870[31 : 0];
  assign _zz_12870 = _zz_12871;
  assign _zz_12871 = ($signed(_zz_12872) >>> _zz_970);
  assign _zz_12872 = _zz_12873;
  assign _zz_12873 = ($signed(_zz_12875) + $signed(_zz_966));
  assign _zz_12874 = ({8'd0,data_mid_1_real} <<< 8);
  assign _zz_12875 = {{8{_zz_12874[23]}}, _zz_12874};
  assign _zz_12876 = fixTo_1162_dout;
  assign _zz_12877 = _zz_12878[31 : 0];
  assign _zz_12878 = _zz_12879;
  assign _zz_12879 = ($signed(_zz_12880) >>> _zz_970);
  assign _zz_12880 = _zz_12881;
  assign _zz_12881 = ($signed(_zz_12883) + $signed(_zz_967));
  assign _zz_12882 = ({8'd0,data_mid_1_imag} <<< 8);
  assign _zz_12883 = {{8{_zz_12882[23]}}, _zz_12882};
  assign _zz_12884 = fixTo_1163_dout;
  assign _zz_12885 = ($signed(twiddle_factor_table_9_real) + $signed(twiddle_factor_table_9_imag));
  assign _zz_12886 = ($signed(_zz_973) - $signed(_zz_12887));
  assign _zz_12887 = ($signed(_zz_12888) * $signed(twiddle_factor_table_9_imag));
  assign _zz_12888 = ($signed(data_mid_10_real) + $signed(data_mid_10_imag));
  assign _zz_12889 = fixTo_1164_dout;
  assign _zz_12890 = ($signed(_zz_973) + $signed(_zz_12891));
  assign _zz_12891 = ($signed(_zz_12892) * $signed(twiddle_factor_table_9_real));
  assign _zz_12892 = ($signed(data_mid_10_imag) - $signed(data_mid_10_real));
  assign _zz_12893 = fixTo_1165_dout;
  assign _zz_12894 = _zz_12895[31 : 0];
  assign _zz_12895 = _zz_12896;
  assign _zz_12896 = ($signed(_zz_12897) >>> _zz_974);
  assign _zz_12897 = _zz_12898;
  assign _zz_12898 = ($signed(_zz_12900) - $signed(_zz_971));
  assign _zz_12899 = ({8'd0,data_mid_2_real} <<< 8);
  assign _zz_12900 = {{8{_zz_12899[23]}}, _zz_12899};
  assign _zz_12901 = fixTo_1166_dout;
  assign _zz_12902 = _zz_12903[31 : 0];
  assign _zz_12903 = _zz_12904;
  assign _zz_12904 = ($signed(_zz_12905) >>> _zz_974);
  assign _zz_12905 = _zz_12906;
  assign _zz_12906 = ($signed(_zz_12908) - $signed(_zz_972));
  assign _zz_12907 = ({8'd0,data_mid_2_imag} <<< 8);
  assign _zz_12908 = {{8{_zz_12907[23]}}, _zz_12907};
  assign _zz_12909 = fixTo_1167_dout;
  assign _zz_12910 = _zz_12911[31 : 0];
  assign _zz_12911 = _zz_12912;
  assign _zz_12912 = ($signed(_zz_12913) >>> _zz_975);
  assign _zz_12913 = _zz_12914;
  assign _zz_12914 = ($signed(_zz_12916) + $signed(_zz_971));
  assign _zz_12915 = ({8'd0,data_mid_2_real} <<< 8);
  assign _zz_12916 = {{8{_zz_12915[23]}}, _zz_12915};
  assign _zz_12917 = fixTo_1168_dout;
  assign _zz_12918 = _zz_12919[31 : 0];
  assign _zz_12919 = _zz_12920;
  assign _zz_12920 = ($signed(_zz_12921) >>> _zz_975);
  assign _zz_12921 = _zz_12922;
  assign _zz_12922 = ($signed(_zz_12924) + $signed(_zz_972));
  assign _zz_12923 = ({8'd0,data_mid_2_imag} <<< 8);
  assign _zz_12924 = {{8{_zz_12923[23]}}, _zz_12923};
  assign _zz_12925 = fixTo_1169_dout;
  assign _zz_12926 = ($signed(twiddle_factor_table_10_real) + $signed(twiddle_factor_table_10_imag));
  assign _zz_12927 = ($signed(_zz_978) - $signed(_zz_12928));
  assign _zz_12928 = ($signed(_zz_12929) * $signed(twiddle_factor_table_10_imag));
  assign _zz_12929 = ($signed(data_mid_11_real) + $signed(data_mid_11_imag));
  assign _zz_12930 = fixTo_1170_dout;
  assign _zz_12931 = ($signed(_zz_978) + $signed(_zz_12932));
  assign _zz_12932 = ($signed(_zz_12933) * $signed(twiddle_factor_table_10_real));
  assign _zz_12933 = ($signed(data_mid_11_imag) - $signed(data_mid_11_real));
  assign _zz_12934 = fixTo_1171_dout;
  assign _zz_12935 = _zz_12936[31 : 0];
  assign _zz_12936 = _zz_12937;
  assign _zz_12937 = ($signed(_zz_12938) >>> _zz_979);
  assign _zz_12938 = _zz_12939;
  assign _zz_12939 = ($signed(_zz_12941) - $signed(_zz_976));
  assign _zz_12940 = ({8'd0,data_mid_3_real} <<< 8);
  assign _zz_12941 = {{8{_zz_12940[23]}}, _zz_12940};
  assign _zz_12942 = fixTo_1172_dout;
  assign _zz_12943 = _zz_12944[31 : 0];
  assign _zz_12944 = _zz_12945;
  assign _zz_12945 = ($signed(_zz_12946) >>> _zz_979);
  assign _zz_12946 = _zz_12947;
  assign _zz_12947 = ($signed(_zz_12949) - $signed(_zz_977));
  assign _zz_12948 = ({8'd0,data_mid_3_imag} <<< 8);
  assign _zz_12949 = {{8{_zz_12948[23]}}, _zz_12948};
  assign _zz_12950 = fixTo_1173_dout;
  assign _zz_12951 = _zz_12952[31 : 0];
  assign _zz_12952 = _zz_12953;
  assign _zz_12953 = ($signed(_zz_12954) >>> _zz_980);
  assign _zz_12954 = _zz_12955;
  assign _zz_12955 = ($signed(_zz_12957) + $signed(_zz_976));
  assign _zz_12956 = ({8'd0,data_mid_3_real} <<< 8);
  assign _zz_12957 = {{8{_zz_12956[23]}}, _zz_12956};
  assign _zz_12958 = fixTo_1174_dout;
  assign _zz_12959 = _zz_12960[31 : 0];
  assign _zz_12960 = _zz_12961;
  assign _zz_12961 = ($signed(_zz_12962) >>> _zz_980);
  assign _zz_12962 = _zz_12963;
  assign _zz_12963 = ($signed(_zz_12965) + $signed(_zz_977));
  assign _zz_12964 = ({8'd0,data_mid_3_imag} <<< 8);
  assign _zz_12965 = {{8{_zz_12964[23]}}, _zz_12964};
  assign _zz_12966 = fixTo_1175_dout;
  assign _zz_12967 = ($signed(twiddle_factor_table_11_real) + $signed(twiddle_factor_table_11_imag));
  assign _zz_12968 = ($signed(_zz_983) - $signed(_zz_12969));
  assign _zz_12969 = ($signed(_zz_12970) * $signed(twiddle_factor_table_11_imag));
  assign _zz_12970 = ($signed(data_mid_12_real) + $signed(data_mid_12_imag));
  assign _zz_12971 = fixTo_1176_dout;
  assign _zz_12972 = ($signed(_zz_983) + $signed(_zz_12973));
  assign _zz_12973 = ($signed(_zz_12974) * $signed(twiddle_factor_table_11_real));
  assign _zz_12974 = ($signed(data_mid_12_imag) - $signed(data_mid_12_real));
  assign _zz_12975 = fixTo_1177_dout;
  assign _zz_12976 = _zz_12977[31 : 0];
  assign _zz_12977 = _zz_12978;
  assign _zz_12978 = ($signed(_zz_12979) >>> _zz_984);
  assign _zz_12979 = _zz_12980;
  assign _zz_12980 = ($signed(_zz_12982) - $signed(_zz_981));
  assign _zz_12981 = ({8'd0,data_mid_4_real} <<< 8);
  assign _zz_12982 = {{8{_zz_12981[23]}}, _zz_12981};
  assign _zz_12983 = fixTo_1178_dout;
  assign _zz_12984 = _zz_12985[31 : 0];
  assign _zz_12985 = _zz_12986;
  assign _zz_12986 = ($signed(_zz_12987) >>> _zz_984);
  assign _zz_12987 = _zz_12988;
  assign _zz_12988 = ($signed(_zz_12990) - $signed(_zz_982));
  assign _zz_12989 = ({8'd0,data_mid_4_imag} <<< 8);
  assign _zz_12990 = {{8{_zz_12989[23]}}, _zz_12989};
  assign _zz_12991 = fixTo_1179_dout;
  assign _zz_12992 = _zz_12993[31 : 0];
  assign _zz_12993 = _zz_12994;
  assign _zz_12994 = ($signed(_zz_12995) >>> _zz_985);
  assign _zz_12995 = _zz_12996;
  assign _zz_12996 = ($signed(_zz_12998) + $signed(_zz_981));
  assign _zz_12997 = ({8'd0,data_mid_4_real} <<< 8);
  assign _zz_12998 = {{8{_zz_12997[23]}}, _zz_12997};
  assign _zz_12999 = fixTo_1180_dout;
  assign _zz_13000 = _zz_13001[31 : 0];
  assign _zz_13001 = _zz_13002;
  assign _zz_13002 = ($signed(_zz_13003) >>> _zz_985);
  assign _zz_13003 = _zz_13004;
  assign _zz_13004 = ($signed(_zz_13006) + $signed(_zz_982));
  assign _zz_13005 = ({8'd0,data_mid_4_imag} <<< 8);
  assign _zz_13006 = {{8{_zz_13005[23]}}, _zz_13005};
  assign _zz_13007 = fixTo_1181_dout;
  assign _zz_13008 = ($signed(twiddle_factor_table_12_real) + $signed(twiddle_factor_table_12_imag));
  assign _zz_13009 = ($signed(_zz_988) - $signed(_zz_13010));
  assign _zz_13010 = ($signed(_zz_13011) * $signed(twiddle_factor_table_12_imag));
  assign _zz_13011 = ($signed(data_mid_13_real) + $signed(data_mid_13_imag));
  assign _zz_13012 = fixTo_1182_dout;
  assign _zz_13013 = ($signed(_zz_988) + $signed(_zz_13014));
  assign _zz_13014 = ($signed(_zz_13015) * $signed(twiddle_factor_table_12_real));
  assign _zz_13015 = ($signed(data_mid_13_imag) - $signed(data_mid_13_real));
  assign _zz_13016 = fixTo_1183_dout;
  assign _zz_13017 = _zz_13018[31 : 0];
  assign _zz_13018 = _zz_13019;
  assign _zz_13019 = ($signed(_zz_13020) >>> _zz_989);
  assign _zz_13020 = _zz_13021;
  assign _zz_13021 = ($signed(_zz_13023) - $signed(_zz_986));
  assign _zz_13022 = ({8'd0,data_mid_5_real} <<< 8);
  assign _zz_13023 = {{8{_zz_13022[23]}}, _zz_13022};
  assign _zz_13024 = fixTo_1184_dout;
  assign _zz_13025 = _zz_13026[31 : 0];
  assign _zz_13026 = _zz_13027;
  assign _zz_13027 = ($signed(_zz_13028) >>> _zz_989);
  assign _zz_13028 = _zz_13029;
  assign _zz_13029 = ($signed(_zz_13031) - $signed(_zz_987));
  assign _zz_13030 = ({8'd0,data_mid_5_imag} <<< 8);
  assign _zz_13031 = {{8{_zz_13030[23]}}, _zz_13030};
  assign _zz_13032 = fixTo_1185_dout;
  assign _zz_13033 = _zz_13034[31 : 0];
  assign _zz_13034 = _zz_13035;
  assign _zz_13035 = ($signed(_zz_13036) >>> _zz_990);
  assign _zz_13036 = _zz_13037;
  assign _zz_13037 = ($signed(_zz_13039) + $signed(_zz_986));
  assign _zz_13038 = ({8'd0,data_mid_5_real} <<< 8);
  assign _zz_13039 = {{8{_zz_13038[23]}}, _zz_13038};
  assign _zz_13040 = fixTo_1186_dout;
  assign _zz_13041 = _zz_13042[31 : 0];
  assign _zz_13042 = _zz_13043;
  assign _zz_13043 = ($signed(_zz_13044) >>> _zz_990);
  assign _zz_13044 = _zz_13045;
  assign _zz_13045 = ($signed(_zz_13047) + $signed(_zz_987));
  assign _zz_13046 = ({8'd0,data_mid_5_imag} <<< 8);
  assign _zz_13047 = {{8{_zz_13046[23]}}, _zz_13046};
  assign _zz_13048 = fixTo_1187_dout;
  assign _zz_13049 = ($signed(twiddle_factor_table_13_real) + $signed(twiddle_factor_table_13_imag));
  assign _zz_13050 = ($signed(_zz_993) - $signed(_zz_13051));
  assign _zz_13051 = ($signed(_zz_13052) * $signed(twiddle_factor_table_13_imag));
  assign _zz_13052 = ($signed(data_mid_14_real) + $signed(data_mid_14_imag));
  assign _zz_13053 = fixTo_1188_dout;
  assign _zz_13054 = ($signed(_zz_993) + $signed(_zz_13055));
  assign _zz_13055 = ($signed(_zz_13056) * $signed(twiddle_factor_table_13_real));
  assign _zz_13056 = ($signed(data_mid_14_imag) - $signed(data_mid_14_real));
  assign _zz_13057 = fixTo_1189_dout;
  assign _zz_13058 = _zz_13059[31 : 0];
  assign _zz_13059 = _zz_13060;
  assign _zz_13060 = ($signed(_zz_13061) >>> _zz_994);
  assign _zz_13061 = _zz_13062;
  assign _zz_13062 = ($signed(_zz_13064) - $signed(_zz_991));
  assign _zz_13063 = ({8'd0,data_mid_6_real} <<< 8);
  assign _zz_13064 = {{8{_zz_13063[23]}}, _zz_13063};
  assign _zz_13065 = fixTo_1190_dout;
  assign _zz_13066 = _zz_13067[31 : 0];
  assign _zz_13067 = _zz_13068;
  assign _zz_13068 = ($signed(_zz_13069) >>> _zz_994);
  assign _zz_13069 = _zz_13070;
  assign _zz_13070 = ($signed(_zz_13072) - $signed(_zz_992));
  assign _zz_13071 = ({8'd0,data_mid_6_imag} <<< 8);
  assign _zz_13072 = {{8{_zz_13071[23]}}, _zz_13071};
  assign _zz_13073 = fixTo_1191_dout;
  assign _zz_13074 = _zz_13075[31 : 0];
  assign _zz_13075 = _zz_13076;
  assign _zz_13076 = ($signed(_zz_13077) >>> _zz_995);
  assign _zz_13077 = _zz_13078;
  assign _zz_13078 = ($signed(_zz_13080) + $signed(_zz_991));
  assign _zz_13079 = ({8'd0,data_mid_6_real} <<< 8);
  assign _zz_13080 = {{8{_zz_13079[23]}}, _zz_13079};
  assign _zz_13081 = fixTo_1192_dout;
  assign _zz_13082 = _zz_13083[31 : 0];
  assign _zz_13083 = _zz_13084;
  assign _zz_13084 = ($signed(_zz_13085) >>> _zz_995);
  assign _zz_13085 = _zz_13086;
  assign _zz_13086 = ($signed(_zz_13088) + $signed(_zz_992));
  assign _zz_13087 = ({8'd0,data_mid_6_imag} <<< 8);
  assign _zz_13088 = {{8{_zz_13087[23]}}, _zz_13087};
  assign _zz_13089 = fixTo_1193_dout;
  assign _zz_13090 = ($signed(twiddle_factor_table_14_real) + $signed(twiddle_factor_table_14_imag));
  assign _zz_13091 = ($signed(_zz_998) - $signed(_zz_13092));
  assign _zz_13092 = ($signed(_zz_13093) * $signed(twiddle_factor_table_14_imag));
  assign _zz_13093 = ($signed(data_mid_15_real) + $signed(data_mid_15_imag));
  assign _zz_13094 = fixTo_1194_dout;
  assign _zz_13095 = ($signed(_zz_998) + $signed(_zz_13096));
  assign _zz_13096 = ($signed(_zz_13097) * $signed(twiddle_factor_table_14_real));
  assign _zz_13097 = ($signed(data_mid_15_imag) - $signed(data_mid_15_real));
  assign _zz_13098 = fixTo_1195_dout;
  assign _zz_13099 = _zz_13100[31 : 0];
  assign _zz_13100 = _zz_13101;
  assign _zz_13101 = ($signed(_zz_13102) >>> _zz_999);
  assign _zz_13102 = _zz_13103;
  assign _zz_13103 = ($signed(_zz_13105) - $signed(_zz_996));
  assign _zz_13104 = ({8'd0,data_mid_7_real} <<< 8);
  assign _zz_13105 = {{8{_zz_13104[23]}}, _zz_13104};
  assign _zz_13106 = fixTo_1196_dout;
  assign _zz_13107 = _zz_13108[31 : 0];
  assign _zz_13108 = _zz_13109;
  assign _zz_13109 = ($signed(_zz_13110) >>> _zz_999);
  assign _zz_13110 = _zz_13111;
  assign _zz_13111 = ($signed(_zz_13113) - $signed(_zz_997));
  assign _zz_13112 = ({8'd0,data_mid_7_imag} <<< 8);
  assign _zz_13113 = {{8{_zz_13112[23]}}, _zz_13112};
  assign _zz_13114 = fixTo_1197_dout;
  assign _zz_13115 = _zz_13116[31 : 0];
  assign _zz_13116 = _zz_13117;
  assign _zz_13117 = ($signed(_zz_13118) >>> _zz_1000);
  assign _zz_13118 = _zz_13119;
  assign _zz_13119 = ($signed(_zz_13121) + $signed(_zz_996));
  assign _zz_13120 = ({8'd0,data_mid_7_real} <<< 8);
  assign _zz_13121 = {{8{_zz_13120[23]}}, _zz_13120};
  assign _zz_13122 = fixTo_1198_dout;
  assign _zz_13123 = _zz_13124[31 : 0];
  assign _zz_13124 = _zz_13125;
  assign _zz_13125 = ($signed(_zz_13126) >>> _zz_1000);
  assign _zz_13126 = _zz_13127;
  assign _zz_13127 = ($signed(_zz_13129) + $signed(_zz_997));
  assign _zz_13128 = ({8'd0,data_mid_7_imag} <<< 8);
  assign _zz_13129 = {{8{_zz_13128[23]}}, _zz_13128};
  assign _zz_13130 = fixTo_1199_dout;
  assign _zz_13131 = ($signed(twiddle_factor_table_7_real) + $signed(twiddle_factor_table_7_imag));
  assign _zz_13132 = ($signed(_zz_1003) - $signed(_zz_13133));
  assign _zz_13133 = ($signed(_zz_13134) * $signed(twiddle_factor_table_7_imag));
  assign _zz_13134 = ($signed(data_mid_24_real) + $signed(data_mid_24_imag));
  assign _zz_13135 = fixTo_1200_dout;
  assign _zz_13136 = ($signed(_zz_1003) + $signed(_zz_13137));
  assign _zz_13137 = ($signed(_zz_13138) * $signed(twiddle_factor_table_7_real));
  assign _zz_13138 = ($signed(data_mid_24_imag) - $signed(data_mid_24_real));
  assign _zz_13139 = fixTo_1201_dout;
  assign _zz_13140 = _zz_13141[31 : 0];
  assign _zz_13141 = _zz_13142;
  assign _zz_13142 = ($signed(_zz_13143) >>> _zz_1004);
  assign _zz_13143 = _zz_13144;
  assign _zz_13144 = ($signed(_zz_13146) - $signed(_zz_1001));
  assign _zz_13145 = ({8'd0,data_mid_16_real} <<< 8);
  assign _zz_13146 = {{8{_zz_13145[23]}}, _zz_13145};
  assign _zz_13147 = fixTo_1202_dout;
  assign _zz_13148 = _zz_13149[31 : 0];
  assign _zz_13149 = _zz_13150;
  assign _zz_13150 = ($signed(_zz_13151) >>> _zz_1004);
  assign _zz_13151 = _zz_13152;
  assign _zz_13152 = ($signed(_zz_13154) - $signed(_zz_1002));
  assign _zz_13153 = ({8'd0,data_mid_16_imag} <<< 8);
  assign _zz_13154 = {{8{_zz_13153[23]}}, _zz_13153};
  assign _zz_13155 = fixTo_1203_dout;
  assign _zz_13156 = _zz_13157[31 : 0];
  assign _zz_13157 = _zz_13158;
  assign _zz_13158 = ($signed(_zz_13159) >>> _zz_1005);
  assign _zz_13159 = _zz_13160;
  assign _zz_13160 = ($signed(_zz_13162) + $signed(_zz_1001));
  assign _zz_13161 = ({8'd0,data_mid_16_real} <<< 8);
  assign _zz_13162 = {{8{_zz_13161[23]}}, _zz_13161};
  assign _zz_13163 = fixTo_1204_dout;
  assign _zz_13164 = _zz_13165[31 : 0];
  assign _zz_13165 = _zz_13166;
  assign _zz_13166 = ($signed(_zz_13167) >>> _zz_1005);
  assign _zz_13167 = _zz_13168;
  assign _zz_13168 = ($signed(_zz_13170) + $signed(_zz_1002));
  assign _zz_13169 = ({8'd0,data_mid_16_imag} <<< 8);
  assign _zz_13170 = {{8{_zz_13169[23]}}, _zz_13169};
  assign _zz_13171 = fixTo_1205_dout;
  assign _zz_13172 = ($signed(twiddle_factor_table_8_real) + $signed(twiddle_factor_table_8_imag));
  assign _zz_13173 = ($signed(_zz_1008) - $signed(_zz_13174));
  assign _zz_13174 = ($signed(_zz_13175) * $signed(twiddle_factor_table_8_imag));
  assign _zz_13175 = ($signed(data_mid_25_real) + $signed(data_mid_25_imag));
  assign _zz_13176 = fixTo_1206_dout;
  assign _zz_13177 = ($signed(_zz_1008) + $signed(_zz_13178));
  assign _zz_13178 = ($signed(_zz_13179) * $signed(twiddle_factor_table_8_real));
  assign _zz_13179 = ($signed(data_mid_25_imag) - $signed(data_mid_25_real));
  assign _zz_13180 = fixTo_1207_dout;
  assign _zz_13181 = _zz_13182[31 : 0];
  assign _zz_13182 = _zz_13183;
  assign _zz_13183 = ($signed(_zz_13184) >>> _zz_1009);
  assign _zz_13184 = _zz_13185;
  assign _zz_13185 = ($signed(_zz_13187) - $signed(_zz_1006));
  assign _zz_13186 = ({8'd0,data_mid_17_real} <<< 8);
  assign _zz_13187 = {{8{_zz_13186[23]}}, _zz_13186};
  assign _zz_13188 = fixTo_1208_dout;
  assign _zz_13189 = _zz_13190[31 : 0];
  assign _zz_13190 = _zz_13191;
  assign _zz_13191 = ($signed(_zz_13192) >>> _zz_1009);
  assign _zz_13192 = _zz_13193;
  assign _zz_13193 = ($signed(_zz_13195) - $signed(_zz_1007));
  assign _zz_13194 = ({8'd0,data_mid_17_imag} <<< 8);
  assign _zz_13195 = {{8{_zz_13194[23]}}, _zz_13194};
  assign _zz_13196 = fixTo_1209_dout;
  assign _zz_13197 = _zz_13198[31 : 0];
  assign _zz_13198 = _zz_13199;
  assign _zz_13199 = ($signed(_zz_13200) >>> _zz_1010);
  assign _zz_13200 = _zz_13201;
  assign _zz_13201 = ($signed(_zz_13203) + $signed(_zz_1006));
  assign _zz_13202 = ({8'd0,data_mid_17_real} <<< 8);
  assign _zz_13203 = {{8{_zz_13202[23]}}, _zz_13202};
  assign _zz_13204 = fixTo_1210_dout;
  assign _zz_13205 = _zz_13206[31 : 0];
  assign _zz_13206 = _zz_13207;
  assign _zz_13207 = ($signed(_zz_13208) >>> _zz_1010);
  assign _zz_13208 = _zz_13209;
  assign _zz_13209 = ($signed(_zz_13211) + $signed(_zz_1007));
  assign _zz_13210 = ({8'd0,data_mid_17_imag} <<< 8);
  assign _zz_13211 = {{8{_zz_13210[23]}}, _zz_13210};
  assign _zz_13212 = fixTo_1211_dout;
  assign _zz_13213 = ($signed(twiddle_factor_table_9_real) + $signed(twiddle_factor_table_9_imag));
  assign _zz_13214 = ($signed(_zz_1013) - $signed(_zz_13215));
  assign _zz_13215 = ($signed(_zz_13216) * $signed(twiddle_factor_table_9_imag));
  assign _zz_13216 = ($signed(data_mid_26_real) + $signed(data_mid_26_imag));
  assign _zz_13217 = fixTo_1212_dout;
  assign _zz_13218 = ($signed(_zz_1013) + $signed(_zz_13219));
  assign _zz_13219 = ($signed(_zz_13220) * $signed(twiddle_factor_table_9_real));
  assign _zz_13220 = ($signed(data_mid_26_imag) - $signed(data_mid_26_real));
  assign _zz_13221 = fixTo_1213_dout;
  assign _zz_13222 = _zz_13223[31 : 0];
  assign _zz_13223 = _zz_13224;
  assign _zz_13224 = ($signed(_zz_13225) >>> _zz_1014);
  assign _zz_13225 = _zz_13226;
  assign _zz_13226 = ($signed(_zz_13228) - $signed(_zz_1011));
  assign _zz_13227 = ({8'd0,data_mid_18_real} <<< 8);
  assign _zz_13228 = {{8{_zz_13227[23]}}, _zz_13227};
  assign _zz_13229 = fixTo_1214_dout;
  assign _zz_13230 = _zz_13231[31 : 0];
  assign _zz_13231 = _zz_13232;
  assign _zz_13232 = ($signed(_zz_13233) >>> _zz_1014);
  assign _zz_13233 = _zz_13234;
  assign _zz_13234 = ($signed(_zz_13236) - $signed(_zz_1012));
  assign _zz_13235 = ({8'd0,data_mid_18_imag} <<< 8);
  assign _zz_13236 = {{8{_zz_13235[23]}}, _zz_13235};
  assign _zz_13237 = fixTo_1215_dout;
  assign _zz_13238 = _zz_13239[31 : 0];
  assign _zz_13239 = _zz_13240;
  assign _zz_13240 = ($signed(_zz_13241) >>> _zz_1015);
  assign _zz_13241 = _zz_13242;
  assign _zz_13242 = ($signed(_zz_13244) + $signed(_zz_1011));
  assign _zz_13243 = ({8'd0,data_mid_18_real} <<< 8);
  assign _zz_13244 = {{8{_zz_13243[23]}}, _zz_13243};
  assign _zz_13245 = fixTo_1216_dout;
  assign _zz_13246 = _zz_13247[31 : 0];
  assign _zz_13247 = _zz_13248;
  assign _zz_13248 = ($signed(_zz_13249) >>> _zz_1015);
  assign _zz_13249 = _zz_13250;
  assign _zz_13250 = ($signed(_zz_13252) + $signed(_zz_1012));
  assign _zz_13251 = ({8'd0,data_mid_18_imag} <<< 8);
  assign _zz_13252 = {{8{_zz_13251[23]}}, _zz_13251};
  assign _zz_13253 = fixTo_1217_dout;
  assign _zz_13254 = ($signed(twiddle_factor_table_10_real) + $signed(twiddle_factor_table_10_imag));
  assign _zz_13255 = ($signed(_zz_1018) - $signed(_zz_13256));
  assign _zz_13256 = ($signed(_zz_13257) * $signed(twiddle_factor_table_10_imag));
  assign _zz_13257 = ($signed(data_mid_27_real) + $signed(data_mid_27_imag));
  assign _zz_13258 = fixTo_1218_dout;
  assign _zz_13259 = ($signed(_zz_1018) + $signed(_zz_13260));
  assign _zz_13260 = ($signed(_zz_13261) * $signed(twiddle_factor_table_10_real));
  assign _zz_13261 = ($signed(data_mid_27_imag) - $signed(data_mid_27_real));
  assign _zz_13262 = fixTo_1219_dout;
  assign _zz_13263 = _zz_13264[31 : 0];
  assign _zz_13264 = _zz_13265;
  assign _zz_13265 = ($signed(_zz_13266) >>> _zz_1019);
  assign _zz_13266 = _zz_13267;
  assign _zz_13267 = ($signed(_zz_13269) - $signed(_zz_1016));
  assign _zz_13268 = ({8'd0,data_mid_19_real} <<< 8);
  assign _zz_13269 = {{8{_zz_13268[23]}}, _zz_13268};
  assign _zz_13270 = fixTo_1220_dout;
  assign _zz_13271 = _zz_13272[31 : 0];
  assign _zz_13272 = _zz_13273;
  assign _zz_13273 = ($signed(_zz_13274) >>> _zz_1019);
  assign _zz_13274 = _zz_13275;
  assign _zz_13275 = ($signed(_zz_13277) - $signed(_zz_1017));
  assign _zz_13276 = ({8'd0,data_mid_19_imag} <<< 8);
  assign _zz_13277 = {{8{_zz_13276[23]}}, _zz_13276};
  assign _zz_13278 = fixTo_1221_dout;
  assign _zz_13279 = _zz_13280[31 : 0];
  assign _zz_13280 = _zz_13281;
  assign _zz_13281 = ($signed(_zz_13282) >>> _zz_1020);
  assign _zz_13282 = _zz_13283;
  assign _zz_13283 = ($signed(_zz_13285) + $signed(_zz_1016));
  assign _zz_13284 = ({8'd0,data_mid_19_real} <<< 8);
  assign _zz_13285 = {{8{_zz_13284[23]}}, _zz_13284};
  assign _zz_13286 = fixTo_1222_dout;
  assign _zz_13287 = _zz_13288[31 : 0];
  assign _zz_13288 = _zz_13289;
  assign _zz_13289 = ($signed(_zz_13290) >>> _zz_1020);
  assign _zz_13290 = _zz_13291;
  assign _zz_13291 = ($signed(_zz_13293) + $signed(_zz_1017));
  assign _zz_13292 = ({8'd0,data_mid_19_imag} <<< 8);
  assign _zz_13293 = {{8{_zz_13292[23]}}, _zz_13292};
  assign _zz_13294 = fixTo_1223_dout;
  assign _zz_13295 = ($signed(twiddle_factor_table_11_real) + $signed(twiddle_factor_table_11_imag));
  assign _zz_13296 = ($signed(_zz_1023) - $signed(_zz_13297));
  assign _zz_13297 = ($signed(_zz_13298) * $signed(twiddle_factor_table_11_imag));
  assign _zz_13298 = ($signed(data_mid_28_real) + $signed(data_mid_28_imag));
  assign _zz_13299 = fixTo_1224_dout;
  assign _zz_13300 = ($signed(_zz_1023) + $signed(_zz_13301));
  assign _zz_13301 = ($signed(_zz_13302) * $signed(twiddle_factor_table_11_real));
  assign _zz_13302 = ($signed(data_mid_28_imag) - $signed(data_mid_28_real));
  assign _zz_13303 = fixTo_1225_dout;
  assign _zz_13304 = _zz_13305[31 : 0];
  assign _zz_13305 = _zz_13306;
  assign _zz_13306 = ($signed(_zz_13307) >>> _zz_1024);
  assign _zz_13307 = _zz_13308;
  assign _zz_13308 = ($signed(_zz_13310) - $signed(_zz_1021));
  assign _zz_13309 = ({8'd0,data_mid_20_real} <<< 8);
  assign _zz_13310 = {{8{_zz_13309[23]}}, _zz_13309};
  assign _zz_13311 = fixTo_1226_dout;
  assign _zz_13312 = _zz_13313[31 : 0];
  assign _zz_13313 = _zz_13314;
  assign _zz_13314 = ($signed(_zz_13315) >>> _zz_1024);
  assign _zz_13315 = _zz_13316;
  assign _zz_13316 = ($signed(_zz_13318) - $signed(_zz_1022));
  assign _zz_13317 = ({8'd0,data_mid_20_imag} <<< 8);
  assign _zz_13318 = {{8{_zz_13317[23]}}, _zz_13317};
  assign _zz_13319 = fixTo_1227_dout;
  assign _zz_13320 = _zz_13321[31 : 0];
  assign _zz_13321 = _zz_13322;
  assign _zz_13322 = ($signed(_zz_13323) >>> _zz_1025);
  assign _zz_13323 = _zz_13324;
  assign _zz_13324 = ($signed(_zz_13326) + $signed(_zz_1021));
  assign _zz_13325 = ({8'd0,data_mid_20_real} <<< 8);
  assign _zz_13326 = {{8{_zz_13325[23]}}, _zz_13325};
  assign _zz_13327 = fixTo_1228_dout;
  assign _zz_13328 = _zz_13329[31 : 0];
  assign _zz_13329 = _zz_13330;
  assign _zz_13330 = ($signed(_zz_13331) >>> _zz_1025);
  assign _zz_13331 = _zz_13332;
  assign _zz_13332 = ($signed(_zz_13334) + $signed(_zz_1022));
  assign _zz_13333 = ({8'd0,data_mid_20_imag} <<< 8);
  assign _zz_13334 = {{8{_zz_13333[23]}}, _zz_13333};
  assign _zz_13335 = fixTo_1229_dout;
  assign _zz_13336 = ($signed(twiddle_factor_table_12_real) + $signed(twiddle_factor_table_12_imag));
  assign _zz_13337 = ($signed(_zz_1028) - $signed(_zz_13338));
  assign _zz_13338 = ($signed(_zz_13339) * $signed(twiddle_factor_table_12_imag));
  assign _zz_13339 = ($signed(data_mid_29_real) + $signed(data_mid_29_imag));
  assign _zz_13340 = fixTo_1230_dout;
  assign _zz_13341 = ($signed(_zz_1028) + $signed(_zz_13342));
  assign _zz_13342 = ($signed(_zz_13343) * $signed(twiddle_factor_table_12_real));
  assign _zz_13343 = ($signed(data_mid_29_imag) - $signed(data_mid_29_real));
  assign _zz_13344 = fixTo_1231_dout;
  assign _zz_13345 = _zz_13346[31 : 0];
  assign _zz_13346 = _zz_13347;
  assign _zz_13347 = ($signed(_zz_13348) >>> _zz_1029);
  assign _zz_13348 = _zz_13349;
  assign _zz_13349 = ($signed(_zz_13351) - $signed(_zz_1026));
  assign _zz_13350 = ({8'd0,data_mid_21_real} <<< 8);
  assign _zz_13351 = {{8{_zz_13350[23]}}, _zz_13350};
  assign _zz_13352 = fixTo_1232_dout;
  assign _zz_13353 = _zz_13354[31 : 0];
  assign _zz_13354 = _zz_13355;
  assign _zz_13355 = ($signed(_zz_13356) >>> _zz_1029);
  assign _zz_13356 = _zz_13357;
  assign _zz_13357 = ($signed(_zz_13359) - $signed(_zz_1027));
  assign _zz_13358 = ({8'd0,data_mid_21_imag} <<< 8);
  assign _zz_13359 = {{8{_zz_13358[23]}}, _zz_13358};
  assign _zz_13360 = fixTo_1233_dout;
  assign _zz_13361 = _zz_13362[31 : 0];
  assign _zz_13362 = _zz_13363;
  assign _zz_13363 = ($signed(_zz_13364) >>> _zz_1030);
  assign _zz_13364 = _zz_13365;
  assign _zz_13365 = ($signed(_zz_13367) + $signed(_zz_1026));
  assign _zz_13366 = ({8'd0,data_mid_21_real} <<< 8);
  assign _zz_13367 = {{8{_zz_13366[23]}}, _zz_13366};
  assign _zz_13368 = fixTo_1234_dout;
  assign _zz_13369 = _zz_13370[31 : 0];
  assign _zz_13370 = _zz_13371;
  assign _zz_13371 = ($signed(_zz_13372) >>> _zz_1030);
  assign _zz_13372 = _zz_13373;
  assign _zz_13373 = ($signed(_zz_13375) + $signed(_zz_1027));
  assign _zz_13374 = ({8'd0,data_mid_21_imag} <<< 8);
  assign _zz_13375 = {{8{_zz_13374[23]}}, _zz_13374};
  assign _zz_13376 = fixTo_1235_dout;
  assign _zz_13377 = ($signed(twiddle_factor_table_13_real) + $signed(twiddle_factor_table_13_imag));
  assign _zz_13378 = ($signed(_zz_1033) - $signed(_zz_13379));
  assign _zz_13379 = ($signed(_zz_13380) * $signed(twiddle_factor_table_13_imag));
  assign _zz_13380 = ($signed(data_mid_30_real) + $signed(data_mid_30_imag));
  assign _zz_13381 = fixTo_1236_dout;
  assign _zz_13382 = ($signed(_zz_1033) + $signed(_zz_13383));
  assign _zz_13383 = ($signed(_zz_13384) * $signed(twiddle_factor_table_13_real));
  assign _zz_13384 = ($signed(data_mid_30_imag) - $signed(data_mid_30_real));
  assign _zz_13385 = fixTo_1237_dout;
  assign _zz_13386 = _zz_13387[31 : 0];
  assign _zz_13387 = _zz_13388;
  assign _zz_13388 = ($signed(_zz_13389) >>> _zz_1034);
  assign _zz_13389 = _zz_13390;
  assign _zz_13390 = ($signed(_zz_13392) - $signed(_zz_1031));
  assign _zz_13391 = ({8'd0,data_mid_22_real} <<< 8);
  assign _zz_13392 = {{8{_zz_13391[23]}}, _zz_13391};
  assign _zz_13393 = fixTo_1238_dout;
  assign _zz_13394 = _zz_13395[31 : 0];
  assign _zz_13395 = _zz_13396;
  assign _zz_13396 = ($signed(_zz_13397) >>> _zz_1034);
  assign _zz_13397 = _zz_13398;
  assign _zz_13398 = ($signed(_zz_13400) - $signed(_zz_1032));
  assign _zz_13399 = ({8'd0,data_mid_22_imag} <<< 8);
  assign _zz_13400 = {{8{_zz_13399[23]}}, _zz_13399};
  assign _zz_13401 = fixTo_1239_dout;
  assign _zz_13402 = _zz_13403[31 : 0];
  assign _zz_13403 = _zz_13404;
  assign _zz_13404 = ($signed(_zz_13405) >>> _zz_1035);
  assign _zz_13405 = _zz_13406;
  assign _zz_13406 = ($signed(_zz_13408) + $signed(_zz_1031));
  assign _zz_13407 = ({8'd0,data_mid_22_real} <<< 8);
  assign _zz_13408 = {{8{_zz_13407[23]}}, _zz_13407};
  assign _zz_13409 = fixTo_1240_dout;
  assign _zz_13410 = _zz_13411[31 : 0];
  assign _zz_13411 = _zz_13412;
  assign _zz_13412 = ($signed(_zz_13413) >>> _zz_1035);
  assign _zz_13413 = _zz_13414;
  assign _zz_13414 = ($signed(_zz_13416) + $signed(_zz_1032));
  assign _zz_13415 = ({8'd0,data_mid_22_imag} <<< 8);
  assign _zz_13416 = {{8{_zz_13415[23]}}, _zz_13415};
  assign _zz_13417 = fixTo_1241_dout;
  assign _zz_13418 = ($signed(twiddle_factor_table_14_real) + $signed(twiddle_factor_table_14_imag));
  assign _zz_13419 = ($signed(_zz_1038) - $signed(_zz_13420));
  assign _zz_13420 = ($signed(_zz_13421) * $signed(twiddle_factor_table_14_imag));
  assign _zz_13421 = ($signed(data_mid_31_real) + $signed(data_mid_31_imag));
  assign _zz_13422 = fixTo_1242_dout;
  assign _zz_13423 = ($signed(_zz_1038) + $signed(_zz_13424));
  assign _zz_13424 = ($signed(_zz_13425) * $signed(twiddle_factor_table_14_real));
  assign _zz_13425 = ($signed(data_mid_31_imag) - $signed(data_mid_31_real));
  assign _zz_13426 = fixTo_1243_dout;
  assign _zz_13427 = _zz_13428[31 : 0];
  assign _zz_13428 = _zz_13429;
  assign _zz_13429 = ($signed(_zz_13430) >>> _zz_1039);
  assign _zz_13430 = _zz_13431;
  assign _zz_13431 = ($signed(_zz_13433) - $signed(_zz_1036));
  assign _zz_13432 = ({8'd0,data_mid_23_real} <<< 8);
  assign _zz_13433 = {{8{_zz_13432[23]}}, _zz_13432};
  assign _zz_13434 = fixTo_1244_dout;
  assign _zz_13435 = _zz_13436[31 : 0];
  assign _zz_13436 = _zz_13437;
  assign _zz_13437 = ($signed(_zz_13438) >>> _zz_1039);
  assign _zz_13438 = _zz_13439;
  assign _zz_13439 = ($signed(_zz_13441) - $signed(_zz_1037));
  assign _zz_13440 = ({8'd0,data_mid_23_imag} <<< 8);
  assign _zz_13441 = {{8{_zz_13440[23]}}, _zz_13440};
  assign _zz_13442 = fixTo_1245_dout;
  assign _zz_13443 = _zz_13444[31 : 0];
  assign _zz_13444 = _zz_13445;
  assign _zz_13445 = ($signed(_zz_13446) >>> _zz_1040);
  assign _zz_13446 = _zz_13447;
  assign _zz_13447 = ($signed(_zz_13449) + $signed(_zz_1036));
  assign _zz_13448 = ({8'd0,data_mid_23_real} <<< 8);
  assign _zz_13449 = {{8{_zz_13448[23]}}, _zz_13448};
  assign _zz_13450 = fixTo_1246_dout;
  assign _zz_13451 = _zz_13452[31 : 0];
  assign _zz_13452 = _zz_13453;
  assign _zz_13453 = ($signed(_zz_13454) >>> _zz_1040);
  assign _zz_13454 = _zz_13455;
  assign _zz_13455 = ($signed(_zz_13457) + $signed(_zz_1037));
  assign _zz_13456 = ({8'd0,data_mid_23_imag} <<< 8);
  assign _zz_13457 = {{8{_zz_13456[23]}}, _zz_13456};
  assign _zz_13458 = fixTo_1247_dout;
  assign _zz_13459 = ($signed(twiddle_factor_table_7_real) + $signed(twiddle_factor_table_7_imag));
  assign _zz_13460 = ($signed(_zz_1043) - $signed(_zz_13461));
  assign _zz_13461 = ($signed(_zz_13462) * $signed(twiddle_factor_table_7_imag));
  assign _zz_13462 = ($signed(data_mid_40_real) + $signed(data_mid_40_imag));
  assign _zz_13463 = fixTo_1248_dout;
  assign _zz_13464 = ($signed(_zz_1043) + $signed(_zz_13465));
  assign _zz_13465 = ($signed(_zz_13466) * $signed(twiddle_factor_table_7_real));
  assign _zz_13466 = ($signed(data_mid_40_imag) - $signed(data_mid_40_real));
  assign _zz_13467 = fixTo_1249_dout;
  assign _zz_13468 = _zz_13469[31 : 0];
  assign _zz_13469 = _zz_13470;
  assign _zz_13470 = ($signed(_zz_13471) >>> _zz_1044);
  assign _zz_13471 = _zz_13472;
  assign _zz_13472 = ($signed(_zz_13474) - $signed(_zz_1041));
  assign _zz_13473 = ({8'd0,data_mid_32_real} <<< 8);
  assign _zz_13474 = {{8{_zz_13473[23]}}, _zz_13473};
  assign _zz_13475 = fixTo_1250_dout;
  assign _zz_13476 = _zz_13477[31 : 0];
  assign _zz_13477 = _zz_13478;
  assign _zz_13478 = ($signed(_zz_13479) >>> _zz_1044);
  assign _zz_13479 = _zz_13480;
  assign _zz_13480 = ($signed(_zz_13482) - $signed(_zz_1042));
  assign _zz_13481 = ({8'd0,data_mid_32_imag} <<< 8);
  assign _zz_13482 = {{8{_zz_13481[23]}}, _zz_13481};
  assign _zz_13483 = fixTo_1251_dout;
  assign _zz_13484 = _zz_13485[31 : 0];
  assign _zz_13485 = _zz_13486;
  assign _zz_13486 = ($signed(_zz_13487) >>> _zz_1045);
  assign _zz_13487 = _zz_13488;
  assign _zz_13488 = ($signed(_zz_13490) + $signed(_zz_1041));
  assign _zz_13489 = ({8'd0,data_mid_32_real} <<< 8);
  assign _zz_13490 = {{8{_zz_13489[23]}}, _zz_13489};
  assign _zz_13491 = fixTo_1252_dout;
  assign _zz_13492 = _zz_13493[31 : 0];
  assign _zz_13493 = _zz_13494;
  assign _zz_13494 = ($signed(_zz_13495) >>> _zz_1045);
  assign _zz_13495 = _zz_13496;
  assign _zz_13496 = ($signed(_zz_13498) + $signed(_zz_1042));
  assign _zz_13497 = ({8'd0,data_mid_32_imag} <<< 8);
  assign _zz_13498 = {{8{_zz_13497[23]}}, _zz_13497};
  assign _zz_13499 = fixTo_1253_dout;
  assign _zz_13500 = ($signed(twiddle_factor_table_8_real) + $signed(twiddle_factor_table_8_imag));
  assign _zz_13501 = ($signed(_zz_1048) - $signed(_zz_13502));
  assign _zz_13502 = ($signed(_zz_13503) * $signed(twiddle_factor_table_8_imag));
  assign _zz_13503 = ($signed(data_mid_41_real) + $signed(data_mid_41_imag));
  assign _zz_13504 = fixTo_1254_dout;
  assign _zz_13505 = ($signed(_zz_1048) + $signed(_zz_13506));
  assign _zz_13506 = ($signed(_zz_13507) * $signed(twiddle_factor_table_8_real));
  assign _zz_13507 = ($signed(data_mid_41_imag) - $signed(data_mid_41_real));
  assign _zz_13508 = fixTo_1255_dout;
  assign _zz_13509 = _zz_13510[31 : 0];
  assign _zz_13510 = _zz_13511;
  assign _zz_13511 = ($signed(_zz_13512) >>> _zz_1049);
  assign _zz_13512 = _zz_13513;
  assign _zz_13513 = ($signed(_zz_13515) - $signed(_zz_1046));
  assign _zz_13514 = ({8'd0,data_mid_33_real} <<< 8);
  assign _zz_13515 = {{8{_zz_13514[23]}}, _zz_13514};
  assign _zz_13516 = fixTo_1256_dout;
  assign _zz_13517 = _zz_13518[31 : 0];
  assign _zz_13518 = _zz_13519;
  assign _zz_13519 = ($signed(_zz_13520) >>> _zz_1049);
  assign _zz_13520 = _zz_13521;
  assign _zz_13521 = ($signed(_zz_13523) - $signed(_zz_1047));
  assign _zz_13522 = ({8'd0,data_mid_33_imag} <<< 8);
  assign _zz_13523 = {{8{_zz_13522[23]}}, _zz_13522};
  assign _zz_13524 = fixTo_1257_dout;
  assign _zz_13525 = _zz_13526[31 : 0];
  assign _zz_13526 = _zz_13527;
  assign _zz_13527 = ($signed(_zz_13528) >>> _zz_1050);
  assign _zz_13528 = _zz_13529;
  assign _zz_13529 = ($signed(_zz_13531) + $signed(_zz_1046));
  assign _zz_13530 = ({8'd0,data_mid_33_real} <<< 8);
  assign _zz_13531 = {{8{_zz_13530[23]}}, _zz_13530};
  assign _zz_13532 = fixTo_1258_dout;
  assign _zz_13533 = _zz_13534[31 : 0];
  assign _zz_13534 = _zz_13535;
  assign _zz_13535 = ($signed(_zz_13536) >>> _zz_1050);
  assign _zz_13536 = _zz_13537;
  assign _zz_13537 = ($signed(_zz_13539) + $signed(_zz_1047));
  assign _zz_13538 = ({8'd0,data_mid_33_imag} <<< 8);
  assign _zz_13539 = {{8{_zz_13538[23]}}, _zz_13538};
  assign _zz_13540 = fixTo_1259_dout;
  assign _zz_13541 = ($signed(twiddle_factor_table_9_real) + $signed(twiddle_factor_table_9_imag));
  assign _zz_13542 = ($signed(_zz_1053) - $signed(_zz_13543));
  assign _zz_13543 = ($signed(_zz_13544) * $signed(twiddle_factor_table_9_imag));
  assign _zz_13544 = ($signed(data_mid_42_real) + $signed(data_mid_42_imag));
  assign _zz_13545 = fixTo_1260_dout;
  assign _zz_13546 = ($signed(_zz_1053) + $signed(_zz_13547));
  assign _zz_13547 = ($signed(_zz_13548) * $signed(twiddle_factor_table_9_real));
  assign _zz_13548 = ($signed(data_mid_42_imag) - $signed(data_mid_42_real));
  assign _zz_13549 = fixTo_1261_dout;
  assign _zz_13550 = _zz_13551[31 : 0];
  assign _zz_13551 = _zz_13552;
  assign _zz_13552 = ($signed(_zz_13553) >>> _zz_1054);
  assign _zz_13553 = _zz_13554;
  assign _zz_13554 = ($signed(_zz_13556) - $signed(_zz_1051));
  assign _zz_13555 = ({8'd0,data_mid_34_real} <<< 8);
  assign _zz_13556 = {{8{_zz_13555[23]}}, _zz_13555};
  assign _zz_13557 = fixTo_1262_dout;
  assign _zz_13558 = _zz_13559[31 : 0];
  assign _zz_13559 = _zz_13560;
  assign _zz_13560 = ($signed(_zz_13561) >>> _zz_1054);
  assign _zz_13561 = _zz_13562;
  assign _zz_13562 = ($signed(_zz_13564) - $signed(_zz_1052));
  assign _zz_13563 = ({8'd0,data_mid_34_imag} <<< 8);
  assign _zz_13564 = {{8{_zz_13563[23]}}, _zz_13563};
  assign _zz_13565 = fixTo_1263_dout;
  assign _zz_13566 = _zz_13567[31 : 0];
  assign _zz_13567 = _zz_13568;
  assign _zz_13568 = ($signed(_zz_13569) >>> _zz_1055);
  assign _zz_13569 = _zz_13570;
  assign _zz_13570 = ($signed(_zz_13572) + $signed(_zz_1051));
  assign _zz_13571 = ({8'd0,data_mid_34_real} <<< 8);
  assign _zz_13572 = {{8{_zz_13571[23]}}, _zz_13571};
  assign _zz_13573 = fixTo_1264_dout;
  assign _zz_13574 = _zz_13575[31 : 0];
  assign _zz_13575 = _zz_13576;
  assign _zz_13576 = ($signed(_zz_13577) >>> _zz_1055);
  assign _zz_13577 = _zz_13578;
  assign _zz_13578 = ($signed(_zz_13580) + $signed(_zz_1052));
  assign _zz_13579 = ({8'd0,data_mid_34_imag} <<< 8);
  assign _zz_13580 = {{8{_zz_13579[23]}}, _zz_13579};
  assign _zz_13581 = fixTo_1265_dout;
  assign _zz_13582 = ($signed(twiddle_factor_table_10_real) + $signed(twiddle_factor_table_10_imag));
  assign _zz_13583 = ($signed(_zz_1058) - $signed(_zz_13584));
  assign _zz_13584 = ($signed(_zz_13585) * $signed(twiddle_factor_table_10_imag));
  assign _zz_13585 = ($signed(data_mid_43_real) + $signed(data_mid_43_imag));
  assign _zz_13586 = fixTo_1266_dout;
  assign _zz_13587 = ($signed(_zz_1058) + $signed(_zz_13588));
  assign _zz_13588 = ($signed(_zz_13589) * $signed(twiddle_factor_table_10_real));
  assign _zz_13589 = ($signed(data_mid_43_imag) - $signed(data_mid_43_real));
  assign _zz_13590 = fixTo_1267_dout;
  assign _zz_13591 = _zz_13592[31 : 0];
  assign _zz_13592 = _zz_13593;
  assign _zz_13593 = ($signed(_zz_13594) >>> _zz_1059);
  assign _zz_13594 = _zz_13595;
  assign _zz_13595 = ($signed(_zz_13597) - $signed(_zz_1056));
  assign _zz_13596 = ({8'd0,data_mid_35_real} <<< 8);
  assign _zz_13597 = {{8{_zz_13596[23]}}, _zz_13596};
  assign _zz_13598 = fixTo_1268_dout;
  assign _zz_13599 = _zz_13600[31 : 0];
  assign _zz_13600 = _zz_13601;
  assign _zz_13601 = ($signed(_zz_13602) >>> _zz_1059);
  assign _zz_13602 = _zz_13603;
  assign _zz_13603 = ($signed(_zz_13605) - $signed(_zz_1057));
  assign _zz_13604 = ({8'd0,data_mid_35_imag} <<< 8);
  assign _zz_13605 = {{8{_zz_13604[23]}}, _zz_13604};
  assign _zz_13606 = fixTo_1269_dout;
  assign _zz_13607 = _zz_13608[31 : 0];
  assign _zz_13608 = _zz_13609;
  assign _zz_13609 = ($signed(_zz_13610) >>> _zz_1060);
  assign _zz_13610 = _zz_13611;
  assign _zz_13611 = ($signed(_zz_13613) + $signed(_zz_1056));
  assign _zz_13612 = ({8'd0,data_mid_35_real} <<< 8);
  assign _zz_13613 = {{8{_zz_13612[23]}}, _zz_13612};
  assign _zz_13614 = fixTo_1270_dout;
  assign _zz_13615 = _zz_13616[31 : 0];
  assign _zz_13616 = _zz_13617;
  assign _zz_13617 = ($signed(_zz_13618) >>> _zz_1060);
  assign _zz_13618 = _zz_13619;
  assign _zz_13619 = ($signed(_zz_13621) + $signed(_zz_1057));
  assign _zz_13620 = ({8'd0,data_mid_35_imag} <<< 8);
  assign _zz_13621 = {{8{_zz_13620[23]}}, _zz_13620};
  assign _zz_13622 = fixTo_1271_dout;
  assign _zz_13623 = ($signed(twiddle_factor_table_11_real) + $signed(twiddle_factor_table_11_imag));
  assign _zz_13624 = ($signed(_zz_1063) - $signed(_zz_13625));
  assign _zz_13625 = ($signed(_zz_13626) * $signed(twiddle_factor_table_11_imag));
  assign _zz_13626 = ($signed(data_mid_44_real) + $signed(data_mid_44_imag));
  assign _zz_13627 = fixTo_1272_dout;
  assign _zz_13628 = ($signed(_zz_1063) + $signed(_zz_13629));
  assign _zz_13629 = ($signed(_zz_13630) * $signed(twiddle_factor_table_11_real));
  assign _zz_13630 = ($signed(data_mid_44_imag) - $signed(data_mid_44_real));
  assign _zz_13631 = fixTo_1273_dout;
  assign _zz_13632 = _zz_13633[31 : 0];
  assign _zz_13633 = _zz_13634;
  assign _zz_13634 = ($signed(_zz_13635) >>> _zz_1064);
  assign _zz_13635 = _zz_13636;
  assign _zz_13636 = ($signed(_zz_13638) - $signed(_zz_1061));
  assign _zz_13637 = ({8'd0,data_mid_36_real} <<< 8);
  assign _zz_13638 = {{8{_zz_13637[23]}}, _zz_13637};
  assign _zz_13639 = fixTo_1274_dout;
  assign _zz_13640 = _zz_13641[31 : 0];
  assign _zz_13641 = _zz_13642;
  assign _zz_13642 = ($signed(_zz_13643) >>> _zz_1064);
  assign _zz_13643 = _zz_13644;
  assign _zz_13644 = ($signed(_zz_13646) - $signed(_zz_1062));
  assign _zz_13645 = ({8'd0,data_mid_36_imag} <<< 8);
  assign _zz_13646 = {{8{_zz_13645[23]}}, _zz_13645};
  assign _zz_13647 = fixTo_1275_dout;
  assign _zz_13648 = _zz_13649[31 : 0];
  assign _zz_13649 = _zz_13650;
  assign _zz_13650 = ($signed(_zz_13651) >>> _zz_1065);
  assign _zz_13651 = _zz_13652;
  assign _zz_13652 = ($signed(_zz_13654) + $signed(_zz_1061));
  assign _zz_13653 = ({8'd0,data_mid_36_real} <<< 8);
  assign _zz_13654 = {{8{_zz_13653[23]}}, _zz_13653};
  assign _zz_13655 = fixTo_1276_dout;
  assign _zz_13656 = _zz_13657[31 : 0];
  assign _zz_13657 = _zz_13658;
  assign _zz_13658 = ($signed(_zz_13659) >>> _zz_1065);
  assign _zz_13659 = _zz_13660;
  assign _zz_13660 = ($signed(_zz_13662) + $signed(_zz_1062));
  assign _zz_13661 = ({8'd0,data_mid_36_imag} <<< 8);
  assign _zz_13662 = {{8{_zz_13661[23]}}, _zz_13661};
  assign _zz_13663 = fixTo_1277_dout;
  assign _zz_13664 = ($signed(twiddle_factor_table_12_real) + $signed(twiddle_factor_table_12_imag));
  assign _zz_13665 = ($signed(_zz_1068) - $signed(_zz_13666));
  assign _zz_13666 = ($signed(_zz_13667) * $signed(twiddle_factor_table_12_imag));
  assign _zz_13667 = ($signed(data_mid_45_real) + $signed(data_mid_45_imag));
  assign _zz_13668 = fixTo_1278_dout;
  assign _zz_13669 = ($signed(_zz_1068) + $signed(_zz_13670));
  assign _zz_13670 = ($signed(_zz_13671) * $signed(twiddle_factor_table_12_real));
  assign _zz_13671 = ($signed(data_mid_45_imag) - $signed(data_mid_45_real));
  assign _zz_13672 = fixTo_1279_dout;
  assign _zz_13673 = _zz_13674[31 : 0];
  assign _zz_13674 = _zz_13675;
  assign _zz_13675 = ($signed(_zz_13676) >>> _zz_1069);
  assign _zz_13676 = _zz_13677;
  assign _zz_13677 = ($signed(_zz_13679) - $signed(_zz_1066));
  assign _zz_13678 = ({8'd0,data_mid_37_real} <<< 8);
  assign _zz_13679 = {{8{_zz_13678[23]}}, _zz_13678};
  assign _zz_13680 = fixTo_1280_dout;
  assign _zz_13681 = _zz_13682[31 : 0];
  assign _zz_13682 = _zz_13683;
  assign _zz_13683 = ($signed(_zz_13684) >>> _zz_1069);
  assign _zz_13684 = _zz_13685;
  assign _zz_13685 = ($signed(_zz_13687) - $signed(_zz_1067));
  assign _zz_13686 = ({8'd0,data_mid_37_imag} <<< 8);
  assign _zz_13687 = {{8{_zz_13686[23]}}, _zz_13686};
  assign _zz_13688 = fixTo_1281_dout;
  assign _zz_13689 = _zz_13690[31 : 0];
  assign _zz_13690 = _zz_13691;
  assign _zz_13691 = ($signed(_zz_13692) >>> _zz_1070);
  assign _zz_13692 = _zz_13693;
  assign _zz_13693 = ($signed(_zz_13695) + $signed(_zz_1066));
  assign _zz_13694 = ({8'd0,data_mid_37_real} <<< 8);
  assign _zz_13695 = {{8{_zz_13694[23]}}, _zz_13694};
  assign _zz_13696 = fixTo_1282_dout;
  assign _zz_13697 = _zz_13698[31 : 0];
  assign _zz_13698 = _zz_13699;
  assign _zz_13699 = ($signed(_zz_13700) >>> _zz_1070);
  assign _zz_13700 = _zz_13701;
  assign _zz_13701 = ($signed(_zz_13703) + $signed(_zz_1067));
  assign _zz_13702 = ({8'd0,data_mid_37_imag} <<< 8);
  assign _zz_13703 = {{8{_zz_13702[23]}}, _zz_13702};
  assign _zz_13704 = fixTo_1283_dout;
  assign _zz_13705 = ($signed(twiddle_factor_table_13_real) + $signed(twiddle_factor_table_13_imag));
  assign _zz_13706 = ($signed(_zz_1073) - $signed(_zz_13707));
  assign _zz_13707 = ($signed(_zz_13708) * $signed(twiddle_factor_table_13_imag));
  assign _zz_13708 = ($signed(data_mid_46_real) + $signed(data_mid_46_imag));
  assign _zz_13709 = fixTo_1284_dout;
  assign _zz_13710 = ($signed(_zz_1073) + $signed(_zz_13711));
  assign _zz_13711 = ($signed(_zz_13712) * $signed(twiddle_factor_table_13_real));
  assign _zz_13712 = ($signed(data_mid_46_imag) - $signed(data_mid_46_real));
  assign _zz_13713 = fixTo_1285_dout;
  assign _zz_13714 = _zz_13715[31 : 0];
  assign _zz_13715 = _zz_13716;
  assign _zz_13716 = ($signed(_zz_13717) >>> _zz_1074);
  assign _zz_13717 = _zz_13718;
  assign _zz_13718 = ($signed(_zz_13720) - $signed(_zz_1071));
  assign _zz_13719 = ({8'd0,data_mid_38_real} <<< 8);
  assign _zz_13720 = {{8{_zz_13719[23]}}, _zz_13719};
  assign _zz_13721 = fixTo_1286_dout;
  assign _zz_13722 = _zz_13723[31 : 0];
  assign _zz_13723 = _zz_13724;
  assign _zz_13724 = ($signed(_zz_13725) >>> _zz_1074);
  assign _zz_13725 = _zz_13726;
  assign _zz_13726 = ($signed(_zz_13728) - $signed(_zz_1072));
  assign _zz_13727 = ({8'd0,data_mid_38_imag} <<< 8);
  assign _zz_13728 = {{8{_zz_13727[23]}}, _zz_13727};
  assign _zz_13729 = fixTo_1287_dout;
  assign _zz_13730 = _zz_13731[31 : 0];
  assign _zz_13731 = _zz_13732;
  assign _zz_13732 = ($signed(_zz_13733) >>> _zz_1075);
  assign _zz_13733 = _zz_13734;
  assign _zz_13734 = ($signed(_zz_13736) + $signed(_zz_1071));
  assign _zz_13735 = ({8'd0,data_mid_38_real} <<< 8);
  assign _zz_13736 = {{8{_zz_13735[23]}}, _zz_13735};
  assign _zz_13737 = fixTo_1288_dout;
  assign _zz_13738 = _zz_13739[31 : 0];
  assign _zz_13739 = _zz_13740;
  assign _zz_13740 = ($signed(_zz_13741) >>> _zz_1075);
  assign _zz_13741 = _zz_13742;
  assign _zz_13742 = ($signed(_zz_13744) + $signed(_zz_1072));
  assign _zz_13743 = ({8'd0,data_mid_38_imag} <<< 8);
  assign _zz_13744 = {{8{_zz_13743[23]}}, _zz_13743};
  assign _zz_13745 = fixTo_1289_dout;
  assign _zz_13746 = ($signed(twiddle_factor_table_14_real) + $signed(twiddle_factor_table_14_imag));
  assign _zz_13747 = ($signed(_zz_1078) - $signed(_zz_13748));
  assign _zz_13748 = ($signed(_zz_13749) * $signed(twiddle_factor_table_14_imag));
  assign _zz_13749 = ($signed(data_mid_47_real) + $signed(data_mid_47_imag));
  assign _zz_13750 = fixTo_1290_dout;
  assign _zz_13751 = ($signed(_zz_1078) + $signed(_zz_13752));
  assign _zz_13752 = ($signed(_zz_13753) * $signed(twiddle_factor_table_14_real));
  assign _zz_13753 = ($signed(data_mid_47_imag) - $signed(data_mid_47_real));
  assign _zz_13754 = fixTo_1291_dout;
  assign _zz_13755 = _zz_13756[31 : 0];
  assign _zz_13756 = _zz_13757;
  assign _zz_13757 = ($signed(_zz_13758) >>> _zz_1079);
  assign _zz_13758 = _zz_13759;
  assign _zz_13759 = ($signed(_zz_13761) - $signed(_zz_1076));
  assign _zz_13760 = ({8'd0,data_mid_39_real} <<< 8);
  assign _zz_13761 = {{8{_zz_13760[23]}}, _zz_13760};
  assign _zz_13762 = fixTo_1292_dout;
  assign _zz_13763 = _zz_13764[31 : 0];
  assign _zz_13764 = _zz_13765;
  assign _zz_13765 = ($signed(_zz_13766) >>> _zz_1079);
  assign _zz_13766 = _zz_13767;
  assign _zz_13767 = ($signed(_zz_13769) - $signed(_zz_1077));
  assign _zz_13768 = ({8'd0,data_mid_39_imag} <<< 8);
  assign _zz_13769 = {{8{_zz_13768[23]}}, _zz_13768};
  assign _zz_13770 = fixTo_1293_dout;
  assign _zz_13771 = _zz_13772[31 : 0];
  assign _zz_13772 = _zz_13773;
  assign _zz_13773 = ($signed(_zz_13774) >>> _zz_1080);
  assign _zz_13774 = _zz_13775;
  assign _zz_13775 = ($signed(_zz_13777) + $signed(_zz_1076));
  assign _zz_13776 = ({8'd0,data_mid_39_real} <<< 8);
  assign _zz_13777 = {{8{_zz_13776[23]}}, _zz_13776};
  assign _zz_13778 = fixTo_1294_dout;
  assign _zz_13779 = _zz_13780[31 : 0];
  assign _zz_13780 = _zz_13781;
  assign _zz_13781 = ($signed(_zz_13782) >>> _zz_1080);
  assign _zz_13782 = _zz_13783;
  assign _zz_13783 = ($signed(_zz_13785) + $signed(_zz_1077));
  assign _zz_13784 = ({8'd0,data_mid_39_imag} <<< 8);
  assign _zz_13785 = {{8{_zz_13784[23]}}, _zz_13784};
  assign _zz_13786 = fixTo_1295_dout;
  assign _zz_13787 = ($signed(twiddle_factor_table_7_real) + $signed(twiddle_factor_table_7_imag));
  assign _zz_13788 = ($signed(_zz_1083) - $signed(_zz_13789));
  assign _zz_13789 = ($signed(_zz_13790) * $signed(twiddle_factor_table_7_imag));
  assign _zz_13790 = ($signed(data_mid_56_real) + $signed(data_mid_56_imag));
  assign _zz_13791 = fixTo_1296_dout;
  assign _zz_13792 = ($signed(_zz_1083) + $signed(_zz_13793));
  assign _zz_13793 = ($signed(_zz_13794) * $signed(twiddle_factor_table_7_real));
  assign _zz_13794 = ($signed(data_mid_56_imag) - $signed(data_mid_56_real));
  assign _zz_13795 = fixTo_1297_dout;
  assign _zz_13796 = _zz_13797[31 : 0];
  assign _zz_13797 = _zz_13798;
  assign _zz_13798 = ($signed(_zz_13799) >>> _zz_1084);
  assign _zz_13799 = _zz_13800;
  assign _zz_13800 = ($signed(_zz_13802) - $signed(_zz_1081));
  assign _zz_13801 = ({8'd0,data_mid_48_real} <<< 8);
  assign _zz_13802 = {{8{_zz_13801[23]}}, _zz_13801};
  assign _zz_13803 = fixTo_1298_dout;
  assign _zz_13804 = _zz_13805[31 : 0];
  assign _zz_13805 = _zz_13806;
  assign _zz_13806 = ($signed(_zz_13807) >>> _zz_1084);
  assign _zz_13807 = _zz_13808;
  assign _zz_13808 = ($signed(_zz_13810) - $signed(_zz_1082));
  assign _zz_13809 = ({8'd0,data_mid_48_imag} <<< 8);
  assign _zz_13810 = {{8{_zz_13809[23]}}, _zz_13809};
  assign _zz_13811 = fixTo_1299_dout;
  assign _zz_13812 = _zz_13813[31 : 0];
  assign _zz_13813 = _zz_13814;
  assign _zz_13814 = ($signed(_zz_13815) >>> _zz_1085);
  assign _zz_13815 = _zz_13816;
  assign _zz_13816 = ($signed(_zz_13818) + $signed(_zz_1081));
  assign _zz_13817 = ({8'd0,data_mid_48_real} <<< 8);
  assign _zz_13818 = {{8{_zz_13817[23]}}, _zz_13817};
  assign _zz_13819 = fixTo_1300_dout;
  assign _zz_13820 = _zz_13821[31 : 0];
  assign _zz_13821 = _zz_13822;
  assign _zz_13822 = ($signed(_zz_13823) >>> _zz_1085);
  assign _zz_13823 = _zz_13824;
  assign _zz_13824 = ($signed(_zz_13826) + $signed(_zz_1082));
  assign _zz_13825 = ({8'd0,data_mid_48_imag} <<< 8);
  assign _zz_13826 = {{8{_zz_13825[23]}}, _zz_13825};
  assign _zz_13827 = fixTo_1301_dout;
  assign _zz_13828 = ($signed(twiddle_factor_table_8_real) + $signed(twiddle_factor_table_8_imag));
  assign _zz_13829 = ($signed(_zz_1088) - $signed(_zz_13830));
  assign _zz_13830 = ($signed(_zz_13831) * $signed(twiddle_factor_table_8_imag));
  assign _zz_13831 = ($signed(data_mid_57_real) + $signed(data_mid_57_imag));
  assign _zz_13832 = fixTo_1302_dout;
  assign _zz_13833 = ($signed(_zz_1088) + $signed(_zz_13834));
  assign _zz_13834 = ($signed(_zz_13835) * $signed(twiddle_factor_table_8_real));
  assign _zz_13835 = ($signed(data_mid_57_imag) - $signed(data_mid_57_real));
  assign _zz_13836 = fixTo_1303_dout;
  assign _zz_13837 = _zz_13838[31 : 0];
  assign _zz_13838 = _zz_13839;
  assign _zz_13839 = ($signed(_zz_13840) >>> _zz_1089);
  assign _zz_13840 = _zz_13841;
  assign _zz_13841 = ($signed(_zz_13843) - $signed(_zz_1086));
  assign _zz_13842 = ({8'd0,data_mid_49_real} <<< 8);
  assign _zz_13843 = {{8{_zz_13842[23]}}, _zz_13842};
  assign _zz_13844 = fixTo_1304_dout;
  assign _zz_13845 = _zz_13846[31 : 0];
  assign _zz_13846 = _zz_13847;
  assign _zz_13847 = ($signed(_zz_13848) >>> _zz_1089);
  assign _zz_13848 = _zz_13849;
  assign _zz_13849 = ($signed(_zz_13851) - $signed(_zz_1087));
  assign _zz_13850 = ({8'd0,data_mid_49_imag} <<< 8);
  assign _zz_13851 = {{8{_zz_13850[23]}}, _zz_13850};
  assign _zz_13852 = fixTo_1305_dout;
  assign _zz_13853 = _zz_13854[31 : 0];
  assign _zz_13854 = _zz_13855;
  assign _zz_13855 = ($signed(_zz_13856) >>> _zz_1090);
  assign _zz_13856 = _zz_13857;
  assign _zz_13857 = ($signed(_zz_13859) + $signed(_zz_1086));
  assign _zz_13858 = ({8'd0,data_mid_49_real} <<< 8);
  assign _zz_13859 = {{8{_zz_13858[23]}}, _zz_13858};
  assign _zz_13860 = fixTo_1306_dout;
  assign _zz_13861 = _zz_13862[31 : 0];
  assign _zz_13862 = _zz_13863;
  assign _zz_13863 = ($signed(_zz_13864) >>> _zz_1090);
  assign _zz_13864 = _zz_13865;
  assign _zz_13865 = ($signed(_zz_13867) + $signed(_zz_1087));
  assign _zz_13866 = ({8'd0,data_mid_49_imag} <<< 8);
  assign _zz_13867 = {{8{_zz_13866[23]}}, _zz_13866};
  assign _zz_13868 = fixTo_1307_dout;
  assign _zz_13869 = ($signed(twiddle_factor_table_9_real) + $signed(twiddle_factor_table_9_imag));
  assign _zz_13870 = ($signed(_zz_1093) - $signed(_zz_13871));
  assign _zz_13871 = ($signed(_zz_13872) * $signed(twiddle_factor_table_9_imag));
  assign _zz_13872 = ($signed(data_mid_58_real) + $signed(data_mid_58_imag));
  assign _zz_13873 = fixTo_1308_dout;
  assign _zz_13874 = ($signed(_zz_1093) + $signed(_zz_13875));
  assign _zz_13875 = ($signed(_zz_13876) * $signed(twiddle_factor_table_9_real));
  assign _zz_13876 = ($signed(data_mid_58_imag) - $signed(data_mid_58_real));
  assign _zz_13877 = fixTo_1309_dout;
  assign _zz_13878 = _zz_13879[31 : 0];
  assign _zz_13879 = _zz_13880;
  assign _zz_13880 = ($signed(_zz_13881) >>> _zz_1094);
  assign _zz_13881 = _zz_13882;
  assign _zz_13882 = ($signed(_zz_13884) - $signed(_zz_1091));
  assign _zz_13883 = ({8'd0,data_mid_50_real} <<< 8);
  assign _zz_13884 = {{8{_zz_13883[23]}}, _zz_13883};
  assign _zz_13885 = fixTo_1310_dout;
  assign _zz_13886 = _zz_13887[31 : 0];
  assign _zz_13887 = _zz_13888;
  assign _zz_13888 = ($signed(_zz_13889) >>> _zz_1094);
  assign _zz_13889 = _zz_13890;
  assign _zz_13890 = ($signed(_zz_13892) - $signed(_zz_1092));
  assign _zz_13891 = ({8'd0,data_mid_50_imag} <<< 8);
  assign _zz_13892 = {{8{_zz_13891[23]}}, _zz_13891};
  assign _zz_13893 = fixTo_1311_dout;
  assign _zz_13894 = _zz_13895[31 : 0];
  assign _zz_13895 = _zz_13896;
  assign _zz_13896 = ($signed(_zz_13897) >>> _zz_1095);
  assign _zz_13897 = _zz_13898;
  assign _zz_13898 = ($signed(_zz_13900) + $signed(_zz_1091));
  assign _zz_13899 = ({8'd0,data_mid_50_real} <<< 8);
  assign _zz_13900 = {{8{_zz_13899[23]}}, _zz_13899};
  assign _zz_13901 = fixTo_1312_dout;
  assign _zz_13902 = _zz_13903[31 : 0];
  assign _zz_13903 = _zz_13904;
  assign _zz_13904 = ($signed(_zz_13905) >>> _zz_1095);
  assign _zz_13905 = _zz_13906;
  assign _zz_13906 = ($signed(_zz_13908) + $signed(_zz_1092));
  assign _zz_13907 = ({8'd0,data_mid_50_imag} <<< 8);
  assign _zz_13908 = {{8{_zz_13907[23]}}, _zz_13907};
  assign _zz_13909 = fixTo_1313_dout;
  assign _zz_13910 = ($signed(twiddle_factor_table_10_real) + $signed(twiddle_factor_table_10_imag));
  assign _zz_13911 = ($signed(_zz_1098) - $signed(_zz_13912));
  assign _zz_13912 = ($signed(_zz_13913) * $signed(twiddle_factor_table_10_imag));
  assign _zz_13913 = ($signed(data_mid_59_real) + $signed(data_mid_59_imag));
  assign _zz_13914 = fixTo_1314_dout;
  assign _zz_13915 = ($signed(_zz_1098) + $signed(_zz_13916));
  assign _zz_13916 = ($signed(_zz_13917) * $signed(twiddle_factor_table_10_real));
  assign _zz_13917 = ($signed(data_mid_59_imag) - $signed(data_mid_59_real));
  assign _zz_13918 = fixTo_1315_dout;
  assign _zz_13919 = _zz_13920[31 : 0];
  assign _zz_13920 = _zz_13921;
  assign _zz_13921 = ($signed(_zz_13922) >>> _zz_1099);
  assign _zz_13922 = _zz_13923;
  assign _zz_13923 = ($signed(_zz_13925) - $signed(_zz_1096));
  assign _zz_13924 = ({8'd0,data_mid_51_real} <<< 8);
  assign _zz_13925 = {{8{_zz_13924[23]}}, _zz_13924};
  assign _zz_13926 = fixTo_1316_dout;
  assign _zz_13927 = _zz_13928[31 : 0];
  assign _zz_13928 = _zz_13929;
  assign _zz_13929 = ($signed(_zz_13930) >>> _zz_1099);
  assign _zz_13930 = _zz_13931;
  assign _zz_13931 = ($signed(_zz_13933) - $signed(_zz_1097));
  assign _zz_13932 = ({8'd0,data_mid_51_imag} <<< 8);
  assign _zz_13933 = {{8{_zz_13932[23]}}, _zz_13932};
  assign _zz_13934 = fixTo_1317_dout;
  assign _zz_13935 = _zz_13936[31 : 0];
  assign _zz_13936 = _zz_13937;
  assign _zz_13937 = ($signed(_zz_13938) >>> _zz_1100);
  assign _zz_13938 = _zz_13939;
  assign _zz_13939 = ($signed(_zz_13941) + $signed(_zz_1096));
  assign _zz_13940 = ({8'd0,data_mid_51_real} <<< 8);
  assign _zz_13941 = {{8{_zz_13940[23]}}, _zz_13940};
  assign _zz_13942 = fixTo_1318_dout;
  assign _zz_13943 = _zz_13944[31 : 0];
  assign _zz_13944 = _zz_13945;
  assign _zz_13945 = ($signed(_zz_13946) >>> _zz_1100);
  assign _zz_13946 = _zz_13947;
  assign _zz_13947 = ($signed(_zz_13949) + $signed(_zz_1097));
  assign _zz_13948 = ({8'd0,data_mid_51_imag} <<< 8);
  assign _zz_13949 = {{8{_zz_13948[23]}}, _zz_13948};
  assign _zz_13950 = fixTo_1319_dout;
  assign _zz_13951 = ($signed(twiddle_factor_table_11_real) + $signed(twiddle_factor_table_11_imag));
  assign _zz_13952 = ($signed(_zz_1103) - $signed(_zz_13953));
  assign _zz_13953 = ($signed(_zz_13954) * $signed(twiddle_factor_table_11_imag));
  assign _zz_13954 = ($signed(data_mid_60_real) + $signed(data_mid_60_imag));
  assign _zz_13955 = fixTo_1320_dout;
  assign _zz_13956 = ($signed(_zz_1103) + $signed(_zz_13957));
  assign _zz_13957 = ($signed(_zz_13958) * $signed(twiddle_factor_table_11_real));
  assign _zz_13958 = ($signed(data_mid_60_imag) - $signed(data_mid_60_real));
  assign _zz_13959 = fixTo_1321_dout;
  assign _zz_13960 = _zz_13961[31 : 0];
  assign _zz_13961 = _zz_13962;
  assign _zz_13962 = ($signed(_zz_13963) >>> _zz_1104);
  assign _zz_13963 = _zz_13964;
  assign _zz_13964 = ($signed(_zz_13966) - $signed(_zz_1101));
  assign _zz_13965 = ({8'd0,data_mid_52_real} <<< 8);
  assign _zz_13966 = {{8{_zz_13965[23]}}, _zz_13965};
  assign _zz_13967 = fixTo_1322_dout;
  assign _zz_13968 = _zz_13969[31 : 0];
  assign _zz_13969 = _zz_13970;
  assign _zz_13970 = ($signed(_zz_13971) >>> _zz_1104);
  assign _zz_13971 = _zz_13972;
  assign _zz_13972 = ($signed(_zz_13974) - $signed(_zz_1102));
  assign _zz_13973 = ({8'd0,data_mid_52_imag} <<< 8);
  assign _zz_13974 = {{8{_zz_13973[23]}}, _zz_13973};
  assign _zz_13975 = fixTo_1323_dout;
  assign _zz_13976 = _zz_13977[31 : 0];
  assign _zz_13977 = _zz_13978;
  assign _zz_13978 = ($signed(_zz_13979) >>> _zz_1105);
  assign _zz_13979 = _zz_13980;
  assign _zz_13980 = ($signed(_zz_13982) + $signed(_zz_1101));
  assign _zz_13981 = ({8'd0,data_mid_52_real} <<< 8);
  assign _zz_13982 = {{8{_zz_13981[23]}}, _zz_13981};
  assign _zz_13983 = fixTo_1324_dout;
  assign _zz_13984 = _zz_13985[31 : 0];
  assign _zz_13985 = _zz_13986;
  assign _zz_13986 = ($signed(_zz_13987) >>> _zz_1105);
  assign _zz_13987 = _zz_13988;
  assign _zz_13988 = ($signed(_zz_13990) + $signed(_zz_1102));
  assign _zz_13989 = ({8'd0,data_mid_52_imag} <<< 8);
  assign _zz_13990 = {{8{_zz_13989[23]}}, _zz_13989};
  assign _zz_13991 = fixTo_1325_dout;
  assign _zz_13992 = ($signed(twiddle_factor_table_12_real) + $signed(twiddle_factor_table_12_imag));
  assign _zz_13993 = ($signed(_zz_1108) - $signed(_zz_13994));
  assign _zz_13994 = ($signed(_zz_13995) * $signed(twiddle_factor_table_12_imag));
  assign _zz_13995 = ($signed(data_mid_61_real) + $signed(data_mid_61_imag));
  assign _zz_13996 = fixTo_1326_dout;
  assign _zz_13997 = ($signed(_zz_1108) + $signed(_zz_13998));
  assign _zz_13998 = ($signed(_zz_13999) * $signed(twiddle_factor_table_12_real));
  assign _zz_13999 = ($signed(data_mid_61_imag) - $signed(data_mid_61_real));
  assign _zz_14000 = fixTo_1327_dout;
  assign _zz_14001 = _zz_14002[31 : 0];
  assign _zz_14002 = _zz_14003;
  assign _zz_14003 = ($signed(_zz_14004) >>> _zz_1109);
  assign _zz_14004 = _zz_14005;
  assign _zz_14005 = ($signed(_zz_14007) - $signed(_zz_1106));
  assign _zz_14006 = ({8'd0,data_mid_53_real} <<< 8);
  assign _zz_14007 = {{8{_zz_14006[23]}}, _zz_14006};
  assign _zz_14008 = fixTo_1328_dout;
  assign _zz_14009 = _zz_14010[31 : 0];
  assign _zz_14010 = _zz_14011;
  assign _zz_14011 = ($signed(_zz_14012) >>> _zz_1109);
  assign _zz_14012 = _zz_14013;
  assign _zz_14013 = ($signed(_zz_14015) - $signed(_zz_1107));
  assign _zz_14014 = ({8'd0,data_mid_53_imag} <<< 8);
  assign _zz_14015 = {{8{_zz_14014[23]}}, _zz_14014};
  assign _zz_14016 = fixTo_1329_dout;
  assign _zz_14017 = _zz_14018[31 : 0];
  assign _zz_14018 = _zz_14019;
  assign _zz_14019 = ($signed(_zz_14020) >>> _zz_1110);
  assign _zz_14020 = _zz_14021;
  assign _zz_14021 = ($signed(_zz_14023) + $signed(_zz_1106));
  assign _zz_14022 = ({8'd0,data_mid_53_real} <<< 8);
  assign _zz_14023 = {{8{_zz_14022[23]}}, _zz_14022};
  assign _zz_14024 = fixTo_1330_dout;
  assign _zz_14025 = _zz_14026[31 : 0];
  assign _zz_14026 = _zz_14027;
  assign _zz_14027 = ($signed(_zz_14028) >>> _zz_1110);
  assign _zz_14028 = _zz_14029;
  assign _zz_14029 = ($signed(_zz_14031) + $signed(_zz_1107));
  assign _zz_14030 = ({8'd0,data_mid_53_imag} <<< 8);
  assign _zz_14031 = {{8{_zz_14030[23]}}, _zz_14030};
  assign _zz_14032 = fixTo_1331_dout;
  assign _zz_14033 = ($signed(twiddle_factor_table_13_real) + $signed(twiddle_factor_table_13_imag));
  assign _zz_14034 = ($signed(_zz_1113) - $signed(_zz_14035));
  assign _zz_14035 = ($signed(_zz_14036) * $signed(twiddle_factor_table_13_imag));
  assign _zz_14036 = ($signed(data_mid_62_real) + $signed(data_mid_62_imag));
  assign _zz_14037 = fixTo_1332_dout;
  assign _zz_14038 = ($signed(_zz_1113) + $signed(_zz_14039));
  assign _zz_14039 = ($signed(_zz_14040) * $signed(twiddle_factor_table_13_real));
  assign _zz_14040 = ($signed(data_mid_62_imag) - $signed(data_mid_62_real));
  assign _zz_14041 = fixTo_1333_dout;
  assign _zz_14042 = _zz_14043[31 : 0];
  assign _zz_14043 = _zz_14044;
  assign _zz_14044 = ($signed(_zz_14045) >>> _zz_1114);
  assign _zz_14045 = _zz_14046;
  assign _zz_14046 = ($signed(_zz_14048) - $signed(_zz_1111));
  assign _zz_14047 = ({8'd0,data_mid_54_real} <<< 8);
  assign _zz_14048 = {{8{_zz_14047[23]}}, _zz_14047};
  assign _zz_14049 = fixTo_1334_dout;
  assign _zz_14050 = _zz_14051[31 : 0];
  assign _zz_14051 = _zz_14052;
  assign _zz_14052 = ($signed(_zz_14053) >>> _zz_1114);
  assign _zz_14053 = _zz_14054;
  assign _zz_14054 = ($signed(_zz_14056) - $signed(_zz_1112));
  assign _zz_14055 = ({8'd0,data_mid_54_imag} <<< 8);
  assign _zz_14056 = {{8{_zz_14055[23]}}, _zz_14055};
  assign _zz_14057 = fixTo_1335_dout;
  assign _zz_14058 = _zz_14059[31 : 0];
  assign _zz_14059 = _zz_14060;
  assign _zz_14060 = ($signed(_zz_14061) >>> _zz_1115);
  assign _zz_14061 = _zz_14062;
  assign _zz_14062 = ($signed(_zz_14064) + $signed(_zz_1111));
  assign _zz_14063 = ({8'd0,data_mid_54_real} <<< 8);
  assign _zz_14064 = {{8{_zz_14063[23]}}, _zz_14063};
  assign _zz_14065 = fixTo_1336_dout;
  assign _zz_14066 = _zz_14067[31 : 0];
  assign _zz_14067 = _zz_14068;
  assign _zz_14068 = ($signed(_zz_14069) >>> _zz_1115);
  assign _zz_14069 = _zz_14070;
  assign _zz_14070 = ($signed(_zz_14072) + $signed(_zz_1112));
  assign _zz_14071 = ({8'd0,data_mid_54_imag} <<< 8);
  assign _zz_14072 = {{8{_zz_14071[23]}}, _zz_14071};
  assign _zz_14073 = fixTo_1337_dout;
  assign _zz_14074 = ($signed(twiddle_factor_table_14_real) + $signed(twiddle_factor_table_14_imag));
  assign _zz_14075 = ($signed(_zz_1118) - $signed(_zz_14076));
  assign _zz_14076 = ($signed(_zz_14077) * $signed(twiddle_factor_table_14_imag));
  assign _zz_14077 = ($signed(data_mid_63_real) + $signed(data_mid_63_imag));
  assign _zz_14078 = fixTo_1338_dout;
  assign _zz_14079 = ($signed(_zz_1118) + $signed(_zz_14080));
  assign _zz_14080 = ($signed(_zz_14081) * $signed(twiddle_factor_table_14_real));
  assign _zz_14081 = ($signed(data_mid_63_imag) - $signed(data_mid_63_real));
  assign _zz_14082 = fixTo_1339_dout;
  assign _zz_14083 = _zz_14084[31 : 0];
  assign _zz_14084 = _zz_14085;
  assign _zz_14085 = ($signed(_zz_14086) >>> _zz_1119);
  assign _zz_14086 = _zz_14087;
  assign _zz_14087 = ($signed(_zz_14089) - $signed(_zz_1116));
  assign _zz_14088 = ({8'd0,data_mid_55_real} <<< 8);
  assign _zz_14089 = {{8{_zz_14088[23]}}, _zz_14088};
  assign _zz_14090 = fixTo_1340_dout;
  assign _zz_14091 = _zz_14092[31 : 0];
  assign _zz_14092 = _zz_14093;
  assign _zz_14093 = ($signed(_zz_14094) >>> _zz_1119);
  assign _zz_14094 = _zz_14095;
  assign _zz_14095 = ($signed(_zz_14097) - $signed(_zz_1117));
  assign _zz_14096 = ({8'd0,data_mid_55_imag} <<< 8);
  assign _zz_14097 = {{8{_zz_14096[23]}}, _zz_14096};
  assign _zz_14098 = fixTo_1341_dout;
  assign _zz_14099 = _zz_14100[31 : 0];
  assign _zz_14100 = _zz_14101;
  assign _zz_14101 = ($signed(_zz_14102) >>> _zz_1120);
  assign _zz_14102 = _zz_14103;
  assign _zz_14103 = ($signed(_zz_14105) + $signed(_zz_1116));
  assign _zz_14104 = ({8'd0,data_mid_55_real} <<< 8);
  assign _zz_14105 = {{8{_zz_14104[23]}}, _zz_14104};
  assign _zz_14106 = fixTo_1342_dout;
  assign _zz_14107 = _zz_14108[31 : 0];
  assign _zz_14108 = _zz_14109;
  assign _zz_14109 = ($signed(_zz_14110) >>> _zz_1120);
  assign _zz_14110 = _zz_14111;
  assign _zz_14111 = ($signed(_zz_14113) + $signed(_zz_1117));
  assign _zz_14112 = ({8'd0,data_mid_55_imag} <<< 8);
  assign _zz_14113 = {{8{_zz_14112[23]}}, _zz_14112};
  assign _zz_14114 = fixTo_1343_dout;
  assign _zz_14115 = ($signed(twiddle_factor_table_7_real) + $signed(twiddle_factor_table_7_imag));
  assign _zz_14116 = ($signed(_zz_1123) - $signed(_zz_14117));
  assign _zz_14117 = ($signed(_zz_14118) * $signed(twiddle_factor_table_7_imag));
  assign _zz_14118 = ($signed(data_mid_72_real) + $signed(data_mid_72_imag));
  assign _zz_14119 = fixTo_1344_dout;
  assign _zz_14120 = ($signed(_zz_1123) + $signed(_zz_14121));
  assign _zz_14121 = ($signed(_zz_14122) * $signed(twiddle_factor_table_7_real));
  assign _zz_14122 = ($signed(data_mid_72_imag) - $signed(data_mid_72_real));
  assign _zz_14123 = fixTo_1345_dout;
  assign _zz_14124 = _zz_14125[31 : 0];
  assign _zz_14125 = _zz_14126;
  assign _zz_14126 = ($signed(_zz_14127) >>> _zz_1124);
  assign _zz_14127 = _zz_14128;
  assign _zz_14128 = ($signed(_zz_14130) - $signed(_zz_1121));
  assign _zz_14129 = ({8'd0,data_mid_64_real} <<< 8);
  assign _zz_14130 = {{8{_zz_14129[23]}}, _zz_14129};
  assign _zz_14131 = fixTo_1346_dout;
  assign _zz_14132 = _zz_14133[31 : 0];
  assign _zz_14133 = _zz_14134;
  assign _zz_14134 = ($signed(_zz_14135) >>> _zz_1124);
  assign _zz_14135 = _zz_14136;
  assign _zz_14136 = ($signed(_zz_14138) - $signed(_zz_1122));
  assign _zz_14137 = ({8'd0,data_mid_64_imag} <<< 8);
  assign _zz_14138 = {{8{_zz_14137[23]}}, _zz_14137};
  assign _zz_14139 = fixTo_1347_dout;
  assign _zz_14140 = _zz_14141[31 : 0];
  assign _zz_14141 = _zz_14142;
  assign _zz_14142 = ($signed(_zz_14143) >>> _zz_1125);
  assign _zz_14143 = _zz_14144;
  assign _zz_14144 = ($signed(_zz_14146) + $signed(_zz_1121));
  assign _zz_14145 = ({8'd0,data_mid_64_real} <<< 8);
  assign _zz_14146 = {{8{_zz_14145[23]}}, _zz_14145};
  assign _zz_14147 = fixTo_1348_dout;
  assign _zz_14148 = _zz_14149[31 : 0];
  assign _zz_14149 = _zz_14150;
  assign _zz_14150 = ($signed(_zz_14151) >>> _zz_1125);
  assign _zz_14151 = _zz_14152;
  assign _zz_14152 = ($signed(_zz_14154) + $signed(_zz_1122));
  assign _zz_14153 = ({8'd0,data_mid_64_imag} <<< 8);
  assign _zz_14154 = {{8{_zz_14153[23]}}, _zz_14153};
  assign _zz_14155 = fixTo_1349_dout;
  assign _zz_14156 = ($signed(twiddle_factor_table_8_real) + $signed(twiddle_factor_table_8_imag));
  assign _zz_14157 = ($signed(_zz_1128) - $signed(_zz_14158));
  assign _zz_14158 = ($signed(_zz_14159) * $signed(twiddle_factor_table_8_imag));
  assign _zz_14159 = ($signed(data_mid_73_real) + $signed(data_mid_73_imag));
  assign _zz_14160 = fixTo_1350_dout;
  assign _zz_14161 = ($signed(_zz_1128) + $signed(_zz_14162));
  assign _zz_14162 = ($signed(_zz_14163) * $signed(twiddle_factor_table_8_real));
  assign _zz_14163 = ($signed(data_mid_73_imag) - $signed(data_mid_73_real));
  assign _zz_14164 = fixTo_1351_dout;
  assign _zz_14165 = _zz_14166[31 : 0];
  assign _zz_14166 = _zz_14167;
  assign _zz_14167 = ($signed(_zz_14168) >>> _zz_1129);
  assign _zz_14168 = _zz_14169;
  assign _zz_14169 = ($signed(_zz_14171) - $signed(_zz_1126));
  assign _zz_14170 = ({8'd0,data_mid_65_real} <<< 8);
  assign _zz_14171 = {{8{_zz_14170[23]}}, _zz_14170};
  assign _zz_14172 = fixTo_1352_dout;
  assign _zz_14173 = _zz_14174[31 : 0];
  assign _zz_14174 = _zz_14175;
  assign _zz_14175 = ($signed(_zz_14176) >>> _zz_1129);
  assign _zz_14176 = _zz_14177;
  assign _zz_14177 = ($signed(_zz_14179) - $signed(_zz_1127));
  assign _zz_14178 = ({8'd0,data_mid_65_imag} <<< 8);
  assign _zz_14179 = {{8{_zz_14178[23]}}, _zz_14178};
  assign _zz_14180 = fixTo_1353_dout;
  assign _zz_14181 = _zz_14182[31 : 0];
  assign _zz_14182 = _zz_14183;
  assign _zz_14183 = ($signed(_zz_14184) >>> _zz_1130);
  assign _zz_14184 = _zz_14185;
  assign _zz_14185 = ($signed(_zz_14187) + $signed(_zz_1126));
  assign _zz_14186 = ({8'd0,data_mid_65_real} <<< 8);
  assign _zz_14187 = {{8{_zz_14186[23]}}, _zz_14186};
  assign _zz_14188 = fixTo_1354_dout;
  assign _zz_14189 = _zz_14190[31 : 0];
  assign _zz_14190 = _zz_14191;
  assign _zz_14191 = ($signed(_zz_14192) >>> _zz_1130);
  assign _zz_14192 = _zz_14193;
  assign _zz_14193 = ($signed(_zz_14195) + $signed(_zz_1127));
  assign _zz_14194 = ({8'd0,data_mid_65_imag} <<< 8);
  assign _zz_14195 = {{8{_zz_14194[23]}}, _zz_14194};
  assign _zz_14196 = fixTo_1355_dout;
  assign _zz_14197 = ($signed(twiddle_factor_table_9_real) + $signed(twiddle_factor_table_9_imag));
  assign _zz_14198 = ($signed(_zz_1133) - $signed(_zz_14199));
  assign _zz_14199 = ($signed(_zz_14200) * $signed(twiddle_factor_table_9_imag));
  assign _zz_14200 = ($signed(data_mid_74_real) + $signed(data_mid_74_imag));
  assign _zz_14201 = fixTo_1356_dout;
  assign _zz_14202 = ($signed(_zz_1133) + $signed(_zz_14203));
  assign _zz_14203 = ($signed(_zz_14204) * $signed(twiddle_factor_table_9_real));
  assign _zz_14204 = ($signed(data_mid_74_imag) - $signed(data_mid_74_real));
  assign _zz_14205 = fixTo_1357_dout;
  assign _zz_14206 = _zz_14207[31 : 0];
  assign _zz_14207 = _zz_14208;
  assign _zz_14208 = ($signed(_zz_14209) >>> _zz_1134);
  assign _zz_14209 = _zz_14210;
  assign _zz_14210 = ($signed(_zz_14212) - $signed(_zz_1131));
  assign _zz_14211 = ({8'd0,data_mid_66_real} <<< 8);
  assign _zz_14212 = {{8{_zz_14211[23]}}, _zz_14211};
  assign _zz_14213 = fixTo_1358_dout;
  assign _zz_14214 = _zz_14215[31 : 0];
  assign _zz_14215 = _zz_14216;
  assign _zz_14216 = ($signed(_zz_14217) >>> _zz_1134);
  assign _zz_14217 = _zz_14218;
  assign _zz_14218 = ($signed(_zz_14220) - $signed(_zz_1132));
  assign _zz_14219 = ({8'd0,data_mid_66_imag} <<< 8);
  assign _zz_14220 = {{8{_zz_14219[23]}}, _zz_14219};
  assign _zz_14221 = fixTo_1359_dout;
  assign _zz_14222 = _zz_14223[31 : 0];
  assign _zz_14223 = _zz_14224;
  assign _zz_14224 = ($signed(_zz_14225) >>> _zz_1135);
  assign _zz_14225 = _zz_14226;
  assign _zz_14226 = ($signed(_zz_14228) + $signed(_zz_1131));
  assign _zz_14227 = ({8'd0,data_mid_66_real} <<< 8);
  assign _zz_14228 = {{8{_zz_14227[23]}}, _zz_14227};
  assign _zz_14229 = fixTo_1360_dout;
  assign _zz_14230 = _zz_14231[31 : 0];
  assign _zz_14231 = _zz_14232;
  assign _zz_14232 = ($signed(_zz_14233) >>> _zz_1135);
  assign _zz_14233 = _zz_14234;
  assign _zz_14234 = ($signed(_zz_14236) + $signed(_zz_1132));
  assign _zz_14235 = ({8'd0,data_mid_66_imag} <<< 8);
  assign _zz_14236 = {{8{_zz_14235[23]}}, _zz_14235};
  assign _zz_14237 = fixTo_1361_dout;
  assign _zz_14238 = ($signed(twiddle_factor_table_10_real) + $signed(twiddle_factor_table_10_imag));
  assign _zz_14239 = ($signed(_zz_1138) - $signed(_zz_14240));
  assign _zz_14240 = ($signed(_zz_14241) * $signed(twiddle_factor_table_10_imag));
  assign _zz_14241 = ($signed(data_mid_75_real) + $signed(data_mid_75_imag));
  assign _zz_14242 = fixTo_1362_dout;
  assign _zz_14243 = ($signed(_zz_1138) + $signed(_zz_14244));
  assign _zz_14244 = ($signed(_zz_14245) * $signed(twiddle_factor_table_10_real));
  assign _zz_14245 = ($signed(data_mid_75_imag) - $signed(data_mid_75_real));
  assign _zz_14246 = fixTo_1363_dout;
  assign _zz_14247 = _zz_14248[31 : 0];
  assign _zz_14248 = _zz_14249;
  assign _zz_14249 = ($signed(_zz_14250) >>> _zz_1139);
  assign _zz_14250 = _zz_14251;
  assign _zz_14251 = ($signed(_zz_14253) - $signed(_zz_1136));
  assign _zz_14252 = ({8'd0,data_mid_67_real} <<< 8);
  assign _zz_14253 = {{8{_zz_14252[23]}}, _zz_14252};
  assign _zz_14254 = fixTo_1364_dout;
  assign _zz_14255 = _zz_14256[31 : 0];
  assign _zz_14256 = _zz_14257;
  assign _zz_14257 = ($signed(_zz_14258) >>> _zz_1139);
  assign _zz_14258 = _zz_14259;
  assign _zz_14259 = ($signed(_zz_14261) - $signed(_zz_1137));
  assign _zz_14260 = ({8'd0,data_mid_67_imag} <<< 8);
  assign _zz_14261 = {{8{_zz_14260[23]}}, _zz_14260};
  assign _zz_14262 = fixTo_1365_dout;
  assign _zz_14263 = _zz_14264[31 : 0];
  assign _zz_14264 = _zz_14265;
  assign _zz_14265 = ($signed(_zz_14266) >>> _zz_1140);
  assign _zz_14266 = _zz_14267;
  assign _zz_14267 = ($signed(_zz_14269) + $signed(_zz_1136));
  assign _zz_14268 = ({8'd0,data_mid_67_real} <<< 8);
  assign _zz_14269 = {{8{_zz_14268[23]}}, _zz_14268};
  assign _zz_14270 = fixTo_1366_dout;
  assign _zz_14271 = _zz_14272[31 : 0];
  assign _zz_14272 = _zz_14273;
  assign _zz_14273 = ($signed(_zz_14274) >>> _zz_1140);
  assign _zz_14274 = _zz_14275;
  assign _zz_14275 = ($signed(_zz_14277) + $signed(_zz_1137));
  assign _zz_14276 = ({8'd0,data_mid_67_imag} <<< 8);
  assign _zz_14277 = {{8{_zz_14276[23]}}, _zz_14276};
  assign _zz_14278 = fixTo_1367_dout;
  assign _zz_14279 = ($signed(twiddle_factor_table_11_real) + $signed(twiddle_factor_table_11_imag));
  assign _zz_14280 = ($signed(_zz_1143) - $signed(_zz_14281));
  assign _zz_14281 = ($signed(_zz_14282) * $signed(twiddle_factor_table_11_imag));
  assign _zz_14282 = ($signed(data_mid_76_real) + $signed(data_mid_76_imag));
  assign _zz_14283 = fixTo_1368_dout;
  assign _zz_14284 = ($signed(_zz_1143) + $signed(_zz_14285));
  assign _zz_14285 = ($signed(_zz_14286) * $signed(twiddle_factor_table_11_real));
  assign _zz_14286 = ($signed(data_mid_76_imag) - $signed(data_mid_76_real));
  assign _zz_14287 = fixTo_1369_dout;
  assign _zz_14288 = _zz_14289[31 : 0];
  assign _zz_14289 = _zz_14290;
  assign _zz_14290 = ($signed(_zz_14291) >>> _zz_1144);
  assign _zz_14291 = _zz_14292;
  assign _zz_14292 = ($signed(_zz_14294) - $signed(_zz_1141));
  assign _zz_14293 = ({8'd0,data_mid_68_real} <<< 8);
  assign _zz_14294 = {{8{_zz_14293[23]}}, _zz_14293};
  assign _zz_14295 = fixTo_1370_dout;
  assign _zz_14296 = _zz_14297[31 : 0];
  assign _zz_14297 = _zz_14298;
  assign _zz_14298 = ($signed(_zz_14299) >>> _zz_1144);
  assign _zz_14299 = _zz_14300;
  assign _zz_14300 = ($signed(_zz_14302) - $signed(_zz_1142));
  assign _zz_14301 = ({8'd0,data_mid_68_imag} <<< 8);
  assign _zz_14302 = {{8{_zz_14301[23]}}, _zz_14301};
  assign _zz_14303 = fixTo_1371_dout;
  assign _zz_14304 = _zz_14305[31 : 0];
  assign _zz_14305 = _zz_14306;
  assign _zz_14306 = ($signed(_zz_14307) >>> _zz_1145);
  assign _zz_14307 = _zz_14308;
  assign _zz_14308 = ($signed(_zz_14310) + $signed(_zz_1141));
  assign _zz_14309 = ({8'd0,data_mid_68_real} <<< 8);
  assign _zz_14310 = {{8{_zz_14309[23]}}, _zz_14309};
  assign _zz_14311 = fixTo_1372_dout;
  assign _zz_14312 = _zz_14313[31 : 0];
  assign _zz_14313 = _zz_14314;
  assign _zz_14314 = ($signed(_zz_14315) >>> _zz_1145);
  assign _zz_14315 = _zz_14316;
  assign _zz_14316 = ($signed(_zz_14318) + $signed(_zz_1142));
  assign _zz_14317 = ({8'd0,data_mid_68_imag} <<< 8);
  assign _zz_14318 = {{8{_zz_14317[23]}}, _zz_14317};
  assign _zz_14319 = fixTo_1373_dout;
  assign _zz_14320 = ($signed(twiddle_factor_table_12_real) + $signed(twiddle_factor_table_12_imag));
  assign _zz_14321 = ($signed(_zz_1148) - $signed(_zz_14322));
  assign _zz_14322 = ($signed(_zz_14323) * $signed(twiddle_factor_table_12_imag));
  assign _zz_14323 = ($signed(data_mid_77_real) + $signed(data_mid_77_imag));
  assign _zz_14324 = fixTo_1374_dout;
  assign _zz_14325 = ($signed(_zz_1148) + $signed(_zz_14326));
  assign _zz_14326 = ($signed(_zz_14327) * $signed(twiddle_factor_table_12_real));
  assign _zz_14327 = ($signed(data_mid_77_imag) - $signed(data_mid_77_real));
  assign _zz_14328 = fixTo_1375_dout;
  assign _zz_14329 = _zz_14330[31 : 0];
  assign _zz_14330 = _zz_14331;
  assign _zz_14331 = ($signed(_zz_14332) >>> _zz_1149);
  assign _zz_14332 = _zz_14333;
  assign _zz_14333 = ($signed(_zz_14335) - $signed(_zz_1146));
  assign _zz_14334 = ({8'd0,data_mid_69_real} <<< 8);
  assign _zz_14335 = {{8{_zz_14334[23]}}, _zz_14334};
  assign _zz_14336 = fixTo_1376_dout;
  assign _zz_14337 = _zz_14338[31 : 0];
  assign _zz_14338 = _zz_14339;
  assign _zz_14339 = ($signed(_zz_14340) >>> _zz_1149);
  assign _zz_14340 = _zz_14341;
  assign _zz_14341 = ($signed(_zz_14343) - $signed(_zz_1147));
  assign _zz_14342 = ({8'd0,data_mid_69_imag} <<< 8);
  assign _zz_14343 = {{8{_zz_14342[23]}}, _zz_14342};
  assign _zz_14344 = fixTo_1377_dout;
  assign _zz_14345 = _zz_14346[31 : 0];
  assign _zz_14346 = _zz_14347;
  assign _zz_14347 = ($signed(_zz_14348) >>> _zz_1150);
  assign _zz_14348 = _zz_14349;
  assign _zz_14349 = ($signed(_zz_14351) + $signed(_zz_1146));
  assign _zz_14350 = ({8'd0,data_mid_69_real} <<< 8);
  assign _zz_14351 = {{8{_zz_14350[23]}}, _zz_14350};
  assign _zz_14352 = fixTo_1378_dout;
  assign _zz_14353 = _zz_14354[31 : 0];
  assign _zz_14354 = _zz_14355;
  assign _zz_14355 = ($signed(_zz_14356) >>> _zz_1150);
  assign _zz_14356 = _zz_14357;
  assign _zz_14357 = ($signed(_zz_14359) + $signed(_zz_1147));
  assign _zz_14358 = ({8'd0,data_mid_69_imag} <<< 8);
  assign _zz_14359 = {{8{_zz_14358[23]}}, _zz_14358};
  assign _zz_14360 = fixTo_1379_dout;
  assign _zz_14361 = ($signed(twiddle_factor_table_13_real) + $signed(twiddle_factor_table_13_imag));
  assign _zz_14362 = ($signed(_zz_1153) - $signed(_zz_14363));
  assign _zz_14363 = ($signed(_zz_14364) * $signed(twiddle_factor_table_13_imag));
  assign _zz_14364 = ($signed(data_mid_78_real) + $signed(data_mid_78_imag));
  assign _zz_14365 = fixTo_1380_dout;
  assign _zz_14366 = ($signed(_zz_1153) + $signed(_zz_14367));
  assign _zz_14367 = ($signed(_zz_14368) * $signed(twiddle_factor_table_13_real));
  assign _zz_14368 = ($signed(data_mid_78_imag) - $signed(data_mid_78_real));
  assign _zz_14369 = fixTo_1381_dout;
  assign _zz_14370 = _zz_14371[31 : 0];
  assign _zz_14371 = _zz_14372;
  assign _zz_14372 = ($signed(_zz_14373) >>> _zz_1154);
  assign _zz_14373 = _zz_14374;
  assign _zz_14374 = ($signed(_zz_14376) - $signed(_zz_1151));
  assign _zz_14375 = ({8'd0,data_mid_70_real} <<< 8);
  assign _zz_14376 = {{8{_zz_14375[23]}}, _zz_14375};
  assign _zz_14377 = fixTo_1382_dout;
  assign _zz_14378 = _zz_14379[31 : 0];
  assign _zz_14379 = _zz_14380;
  assign _zz_14380 = ($signed(_zz_14381) >>> _zz_1154);
  assign _zz_14381 = _zz_14382;
  assign _zz_14382 = ($signed(_zz_14384) - $signed(_zz_1152));
  assign _zz_14383 = ({8'd0,data_mid_70_imag} <<< 8);
  assign _zz_14384 = {{8{_zz_14383[23]}}, _zz_14383};
  assign _zz_14385 = fixTo_1383_dout;
  assign _zz_14386 = _zz_14387[31 : 0];
  assign _zz_14387 = _zz_14388;
  assign _zz_14388 = ($signed(_zz_14389) >>> _zz_1155);
  assign _zz_14389 = _zz_14390;
  assign _zz_14390 = ($signed(_zz_14392) + $signed(_zz_1151));
  assign _zz_14391 = ({8'd0,data_mid_70_real} <<< 8);
  assign _zz_14392 = {{8{_zz_14391[23]}}, _zz_14391};
  assign _zz_14393 = fixTo_1384_dout;
  assign _zz_14394 = _zz_14395[31 : 0];
  assign _zz_14395 = _zz_14396;
  assign _zz_14396 = ($signed(_zz_14397) >>> _zz_1155);
  assign _zz_14397 = _zz_14398;
  assign _zz_14398 = ($signed(_zz_14400) + $signed(_zz_1152));
  assign _zz_14399 = ({8'd0,data_mid_70_imag} <<< 8);
  assign _zz_14400 = {{8{_zz_14399[23]}}, _zz_14399};
  assign _zz_14401 = fixTo_1385_dout;
  assign _zz_14402 = ($signed(twiddle_factor_table_14_real) + $signed(twiddle_factor_table_14_imag));
  assign _zz_14403 = ($signed(_zz_1158) - $signed(_zz_14404));
  assign _zz_14404 = ($signed(_zz_14405) * $signed(twiddle_factor_table_14_imag));
  assign _zz_14405 = ($signed(data_mid_79_real) + $signed(data_mid_79_imag));
  assign _zz_14406 = fixTo_1386_dout;
  assign _zz_14407 = ($signed(_zz_1158) + $signed(_zz_14408));
  assign _zz_14408 = ($signed(_zz_14409) * $signed(twiddle_factor_table_14_real));
  assign _zz_14409 = ($signed(data_mid_79_imag) - $signed(data_mid_79_real));
  assign _zz_14410 = fixTo_1387_dout;
  assign _zz_14411 = _zz_14412[31 : 0];
  assign _zz_14412 = _zz_14413;
  assign _zz_14413 = ($signed(_zz_14414) >>> _zz_1159);
  assign _zz_14414 = _zz_14415;
  assign _zz_14415 = ($signed(_zz_14417) - $signed(_zz_1156));
  assign _zz_14416 = ({8'd0,data_mid_71_real} <<< 8);
  assign _zz_14417 = {{8{_zz_14416[23]}}, _zz_14416};
  assign _zz_14418 = fixTo_1388_dout;
  assign _zz_14419 = _zz_14420[31 : 0];
  assign _zz_14420 = _zz_14421;
  assign _zz_14421 = ($signed(_zz_14422) >>> _zz_1159);
  assign _zz_14422 = _zz_14423;
  assign _zz_14423 = ($signed(_zz_14425) - $signed(_zz_1157));
  assign _zz_14424 = ({8'd0,data_mid_71_imag} <<< 8);
  assign _zz_14425 = {{8{_zz_14424[23]}}, _zz_14424};
  assign _zz_14426 = fixTo_1389_dout;
  assign _zz_14427 = _zz_14428[31 : 0];
  assign _zz_14428 = _zz_14429;
  assign _zz_14429 = ($signed(_zz_14430) >>> _zz_1160);
  assign _zz_14430 = _zz_14431;
  assign _zz_14431 = ($signed(_zz_14433) + $signed(_zz_1156));
  assign _zz_14432 = ({8'd0,data_mid_71_real} <<< 8);
  assign _zz_14433 = {{8{_zz_14432[23]}}, _zz_14432};
  assign _zz_14434 = fixTo_1390_dout;
  assign _zz_14435 = _zz_14436[31 : 0];
  assign _zz_14436 = _zz_14437;
  assign _zz_14437 = ($signed(_zz_14438) >>> _zz_1160);
  assign _zz_14438 = _zz_14439;
  assign _zz_14439 = ($signed(_zz_14441) + $signed(_zz_1157));
  assign _zz_14440 = ({8'd0,data_mid_71_imag} <<< 8);
  assign _zz_14441 = {{8{_zz_14440[23]}}, _zz_14440};
  assign _zz_14442 = fixTo_1391_dout;
  assign _zz_14443 = ($signed(twiddle_factor_table_7_real) + $signed(twiddle_factor_table_7_imag));
  assign _zz_14444 = ($signed(_zz_1163) - $signed(_zz_14445));
  assign _zz_14445 = ($signed(_zz_14446) * $signed(twiddle_factor_table_7_imag));
  assign _zz_14446 = ($signed(data_mid_88_real) + $signed(data_mid_88_imag));
  assign _zz_14447 = fixTo_1392_dout;
  assign _zz_14448 = ($signed(_zz_1163) + $signed(_zz_14449));
  assign _zz_14449 = ($signed(_zz_14450) * $signed(twiddle_factor_table_7_real));
  assign _zz_14450 = ($signed(data_mid_88_imag) - $signed(data_mid_88_real));
  assign _zz_14451 = fixTo_1393_dout;
  assign _zz_14452 = _zz_14453[31 : 0];
  assign _zz_14453 = _zz_14454;
  assign _zz_14454 = ($signed(_zz_14455) >>> _zz_1164);
  assign _zz_14455 = _zz_14456;
  assign _zz_14456 = ($signed(_zz_14458) - $signed(_zz_1161));
  assign _zz_14457 = ({8'd0,data_mid_80_real} <<< 8);
  assign _zz_14458 = {{8{_zz_14457[23]}}, _zz_14457};
  assign _zz_14459 = fixTo_1394_dout;
  assign _zz_14460 = _zz_14461[31 : 0];
  assign _zz_14461 = _zz_14462;
  assign _zz_14462 = ($signed(_zz_14463) >>> _zz_1164);
  assign _zz_14463 = _zz_14464;
  assign _zz_14464 = ($signed(_zz_14466) - $signed(_zz_1162));
  assign _zz_14465 = ({8'd0,data_mid_80_imag} <<< 8);
  assign _zz_14466 = {{8{_zz_14465[23]}}, _zz_14465};
  assign _zz_14467 = fixTo_1395_dout;
  assign _zz_14468 = _zz_14469[31 : 0];
  assign _zz_14469 = _zz_14470;
  assign _zz_14470 = ($signed(_zz_14471) >>> _zz_1165);
  assign _zz_14471 = _zz_14472;
  assign _zz_14472 = ($signed(_zz_14474) + $signed(_zz_1161));
  assign _zz_14473 = ({8'd0,data_mid_80_real} <<< 8);
  assign _zz_14474 = {{8{_zz_14473[23]}}, _zz_14473};
  assign _zz_14475 = fixTo_1396_dout;
  assign _zz_14476 = _zz_14477[31 : 0];
  assign _zz_14477 = _zz_14478;
  assign _zz_14478 = ($signed(_zz_14479) >>> _zz_1165);
  assign _zz_14479 = _zz_14480;
  assign _zz_14480 = ($signed(_zz_14482) + $signed(_zz_1162));
  assign _zz_14481 = ({8'd0,data_mid_80_imag} <<< 8);
  assign _zz_14482 = {{8{_zz_14481[23]}}, _zz_14481};
  assign _zz_14483 = fixTo_1397_dout;
  assign _zz_14484 = ($signed(twiddle_factor_table_8_real) + $signed(twiddle_factor_table_8_imag));
  assign _zz_14485 = ($signed(_zz_1168) - $signed(_zz_14486));
  assign _zz_14486 = ($signed(_zz_14487) * $signed(twiddle_factor_table_8_imag));
  assign _zz_14487 = ($signed(data_mid_89_real) + $signed(data_mid_89_imag));
  assign _zz_14488 = fixTo_1398_dout;
  assign _zz_14489 = ($signed(_zz_1168) + $signed(_zz_14490));
  assign _zz_14490 = ($signed(_zz_14491) * $signed(twiddle_factor_table_8_real));
  assign _zz_14491 = ($signed(data_mid_89_imag) - $signed(data_mid_89_real));
  assign _zz_14492 = fixTo_1399_dout;
  assign _zz_14493 = _zz_14494[31 : 0];
  assign _zz_14494 = _zz_14495;
  assign _zz_14495 = ($signed(_zz_14496) >>> _zz_1169);
  assign _zz_14496 = _zz_14497;
  assign _zz_14497 = ($signed(_zz_14499) - $signed(_zz_1166));
  assign _zz_14498 = ({8'd0,data_mid_81_real} <<< 8);
  assign _zz_14499 = {{8{_zz_14498[23]}}, _zz_14498};
  assign _zz_14500 = fixTo_1400_dout;
  assign _zz_14501 = _zz_14502[31 : 0];
  assign _zz_14502 = _zz_14503;
  assign _zz_14503 = ($signed(_zz_14504) >>> _zz_1169);
  assign _zz_14504 = _zz_14505;
  assign _zz_14505 = ($signed(_zz_14507) - $signed(_zz_1167));
  assign _zz_14506 = ({8'd0,data_mid_81_imag} <<< 8);
  assign _zz_14507 = {{8{_zz_14506[23]}}, _zz_14506};
  assign _zz_14508 = fixTo_1401_dout;
  assign _zz_14509 = _zz_14510[31 : 0];
  assign _zz_14510 = _zz_14511;
  assign _zz_14511 = ($signed(_zz_14512) >>> _zz_1170);
  assign _zz_14512 = _zz_14513;
  assign _zz_14513 = ($signed(_zz_14515) + $signed(_zz_1166));
  assign _zz_14514 = ({8'd0,data_mid_81_real} <<< 8);
  assign _zz_14515 = {{8{_zz_14514[23]}}, _zz_14514};
  assign _zz_14516 = fixTo_1402_dout;
  assign _zz_14517 = _zz_14518[31 : 0];
  assign _zz_14518 = _zz_14519;
  assign _zz_14519 = ($signed(_zz_14520) >>> _zz_1170);
  assign _zz_14520 = _zz_14521;
  assign _zz_14521 = ($signed(_zz_14523) + $signed(_zz_1167));
  assign _zz_14522 = ({8'd0,data_mid_81_imag} <<< 8);
  assign _zz_14523 = {{8{_zz_14522[23]}}, _zz_14522};
  assign _zz_14524 = fixTo_1403_dout;
  assign _zz_14525 = ($signed(twiddle_factor_table_9_real) + $signed(twiddle_factor_table_9_imag));
  assign _zz_14526 = ($signed(_zz_1173) - $signed(_zz_14527));
  assign _zz_14527 = ($signed(_zz_14528) * $signed(twiddle_factor_table_9_imag));
  assign _zz_14528 = ($signed(data_mid_90_real) + $signed(data_mid_90_imag));
  assign _zz_14529 = fixTo_1404_dout;
  assign _zz_14530 = ($signed(_zz_1173) + $signed(_zz_14531));
  assign _zz_14531 = ($signed(_zz_14532) * $signed(twiddle_factor_table_9_real));
  assign _zz_14532 = ($signed(data_mid_90_imag) - $signed(data_mid_90_real));
  assign _zz_14533 = fixTo_1405_dout;
  assign _zz_14534 = _zz_14535[31 : 0];
  assign _zz_14535 = _zz_14536;
  assign _zz_14536 = ($signed(_zz_14537) >>> _zz_1174);
  assign _zz_14537 = _zz_14538;
  assign _zz_14538 = ($signed(_zz_14540) - $signed(_zz_1171));
  assign _zz_14539 = ({8'd0,data_mid_82_real} <<< 8);
  assign _zz_14540 = {{8{_zz_14539[23]}}, _zz_14539};
  assign _zz_14541 = fixTo_1406_dout;
  assign _zz_14542 = _zz_14543[31 : 0];
  assign _zz_14543 = _zz_14544;
  assign _zz_14544 = ($signed(_zz_14545) >>> _zz_1174);
  assign _zz_14545 = _zz_14546;
  assign _zz_14546 = ($signed(_zz_14548) - $signed(_zz_1172));
  assign _zz_14547 = ({8'd0,data_mid_82_imag} <<< 8);
  assign _zz_14548 = {{8{_zz_14547[23]}}, _zz_14547};
  assign _zz_14549 = fixTo_1407_dout;
  assign _zz_14550 = _zz_14551[31 : 0];
  assign _zz_14551 = _zz_14552;
  assign _zz_14552 = ($signed(_zz_14553) >>> _zz_1175);
  assign _zz_14553 = _zz_14554;
  assign _zz_14554 = ($signed(_zz_14556) + $signed(_zz_1171));
  assign _zz_14555 = ({8'd0,data_mid_82_real} <<< 8);
  assign _zz_14556 = {{8{_zz_14555[23]}}, _zz_14555};
  assign _zz_14557 = fixTo_1408_dout;
  assign _zz_14558 = _zz_14559[31 : 0];
  assign _zz_14559 = _zz_14560;
  assign _zz_14560 = ($signed(_zz_14561) >>> _zz_1175);
  assign _zz_14561 = _zz_14562;
  assign _zz_14562 = ($signed(_zz_14564) + $signed(_zz_1172));
  assign _zz_14563 = ({8'd0,data_mid_82_imag} <<< 8);
  assign _zz_14564 = {{8{_zz_14563[23]}}, _zz_14563};
  assign _zz_14565 = fixTo_1409_dout;
  assign _zz_14566 = ($signed(twiddle_factor_table_10_real) + $signed(twiddle_factor_table_10_imag));
  assign _zz_14567 = ($signed(_zz_1178) - $signed(_zz_14568));
  assign _zz_14568 = ($signed(_zz_14569) * $signed(twiddle_factor_table_10_imag));
  assign _zz_14569 = ($signed(data_mid_91_real) + $signed(data_mid_91_imag));
  assign _zz_14570 = fixTo_1410_dout;
  assign _zz_14571 = ($signed(_zz_1178) + $signed(_zz_14572));
  assign _zz_14572 = ($signed(_zz_14573) * $signed(twiddle_factor_table_10_real));
  assign _zz_14573 = ($signed(data_mid_91_imag) - $signed(data_mid_91_real));
  assign _zz_14574 = fixTo_1411_dout;
  assign _zz_14575 = _zz_14576[31 : 0];
  assign _zz_14576 = _zz_14577;
  assign _zz_14577 = ($signed(_zz_14578) >>> _zz_1179);
  assign _zz_14578 = _zz_14579;
  assign _zz_14579 = ($signed(_zz_14581) - $signed(_zz_1176));
  assign _zz_14580 = ({8'd0,data_mid_83_real} <<< 8);
  assign _zz_14581 = {{8{_zz_14580[23]}}, _zz_14580};
  assign _zz_14582 = fixTo_1412_dout;
  assign _zz_14583 = _zz_14584[31 : 0];
  assign _zz_14584 = _zz_14585;
  assign _zz_14585 = ($signed(_zz_14586) >>> _zz_1179);
  assign _zz_14586 = _zz_14587;
  assign _zz_14587 = ($signed(_zz_14589) - $signed(_zz_1177));
  assign _zz_14588 = ({8'd0,data_mid_83_imag} <<< 8);
  assign _zz_14589 = {{8{_zz_14588[23]}}, _zz_14588};
  assign _zz_14590 = fixTo_1413_dout;
  assign _zz_14591 = _zz_14592[31 : 0];
  assign _zz_14592 = _zz_14593;
  assign _zz_14593 = ($signed(_zz_14594) >>> _zz_1180);
  assign _zz_14594 = _zz_14595;
  assign _zz_14595 = ($signed(_zz_14597) + $signed(_zz_1176));
  assign _zz_14596 = ({8'd0,data_mid_83_real} <<< 8);
  assign _zz_14597 = {{8{_zz_14596[23]}}, _zz_14596};
  assign _zz_14598 = fixTo_1414_dout;
  assign _zz_14599 = _zz_14600[31 : 0];
  assign _zz_14600 = _zz_14601;
  assign _zz_14601 = ($signed(_zz_14602) >>> _zz_1180);
  assign _zz_14602 = _zz_14603;
  assign _zz_14603 = ($signed(_zz_14605) + $signed(_zz_1177));
  assign _zz_14604 = ({8'd0,data_mid_83_imag} <<< 8);
  assign _zz_14605 = {{8{_zz_14604[23]}}, _zz_14604};
  assign _zz_14606 = fixTo_1415_dout;
  assign _zz_14607 = ($signed(twiddle_factor_table_11_real) + $signed(twiddle_factor_table_11_imag));
  assign _zz_14608 = ($signed(_zz_1183) - $signed(_zz_14609));
  assign _zz_14609 = ($signed(_zz_14610) * $signed(twiddle_factor_table_11_imag));
  assign _zz_14610 = ($signed(data_mid_92_real) + $signed(data_mid_92_imag));
  assign _zz_14611 = fixTo_1416_dout;
  assign _zz_14612 = ($signed(_zz_1183) + $signed(_zz_14613));
  assign _zz_14613 = ($signed(_zz_14614) * $signed(twiddle_factor_table_11_real));
  assign _zz_14614 = ($signed(data_mid_92_imag) - $signed(data_mid_92_real));
  assign _zz_14615 = fixTo_1417_dout;
  assign _zz_14616 = _zz_14617[31 : 0];
  assign _zz_14617 = _zz_14618;
  assign _zz_14618 = ($signed(_zz_14619) >>> _zz_1184);
  assign _zz_14619 = _zz_14620;
  assign _zz_14620 = ($signed(_zz_14622) - $signed(_zz_1181));
  assign _zz_14621 = ({8'd0,data_mid_84_real} <<< 8);
  assign _zz_14622 = {{8{_zz_14621[23]}}, _zz_14621};
  assign _zz_14623 = fixTo_1418_dout;
  assign _zz_14624 = _zz_14625[31 : 0];
  assign _zz_14625 = _zz_14626;
  assign _zz_14626 = ($signed(_zz_14627) >>> _zz_1184);
  assign _zz_14627 = _zz_14628;
  assign _zz_14628 = ($signed(_zz_14630) - $signed(_zz_1182));
  assign _zz_14629 = ({8'd0,data_mid_84_imag} <<< 8);
  assign _zz_14630 = {{8{_zz_14629[23]}}, _zz_14629};
  assign _zz_14631 = fixTo_1419_dout;
  assign _zz_14632 = _zz_14633[31 : 0];
  assign _zz_14633 = _zz_14634;
  assign _zz_14634 = ($signed(_zz_14635) >>> _zz_1185);
  assign _zz_14635 = _zz_14636;
  assign _zz_14636 = ($signed(_zz_14638) + $signed(_zz_1181));
  assign _zz_14637 = ({8'd0,data_mid_84_real} <<< 8);
  assign _zz_14638 = {{8{_zz_14637[23]}}, _zz_14637};
  assign _zz_14639 = fixTo_1420_dout;
  assign _zz_14640 = _zz_14641[31 : 0];
  assign _zz_14641 = _zz_14642;
  assign _zz_14642 = ($signed(_zz_14643) >>> _zz_1185);
  assign _zz_14643 = _zz_14644;
  assign _zz_14644 = ($signed(_zz_14646) + $signed(_zz_1182));
  assign _zz_14645 = ({8'd0,data_mid_84_imag} <<< 8);
  assign _zz_14646 = {{8{_zz_14645[23]}}, _zz_14645};
  assign _zz_14647 = fixTo_1421_dout;
  assign _zz_14648 = ($signed(twiddle_factor_table_12_real) + $signed(twiddle_factor_table_12_imag));
  assign _zz_14649 = ($signed(_zz_1188) - $signed(_zz_14650));
  assign _zz_14650 = ($signed(_zz_14651) * $signed(twiddle_factor_table_12_imag));
  assign _zz_14651 = ($signed(data_mid_93_real) + $signed(data_mid_93_imag));
  assign _zz_14652 = fixTo_1422_dout;
  assign _zz_14653 = ($signed(_zz_1188) + $signed(_zz_14654));
  assign _zz_14654 = ($signed(_zz_14655) * $signed(twiddle_factor_table_12_real));
  assign _zz_14655 = ($signed(data_mid_93_imag) - $signed(data_mid_93_real));
  assign _zz_14656 = fixTo_1423_dout;
  assign _zz_14657 = _zz_14658[31 : 0];
  assign _zz_14658 = _zz_14659;
  assign _zz_14659 = ($signed(_zz_14660) >>> _zz_1189);
  assign _zz_14660 = _zz_14661;
  assign _zz_14661 = ($signed(_zz_14663) - $signed(_zz_1186));
  assign _zz_14662 = ({8'd0,data_mid_85_real} <<< 8);
  assign _zz_14663 = {{8{_zz_14662[23]}}, _zz_14662};
  assign _zz_14664 = fixTo_1424_dout;
  assign _zz_14665 = _zz_14666[31 : 0];
  assign _zz_14666 = _zz_14667;
  assign _zz_14667 = ($signed(_zz_14668) >>> _zz_1189);
  assign _zz_14668 = _zz_14669;
  assign _zz_14669 = ($signed(_zz_14671) - $signed(_zz_1187));
  assign _zz_14670 = ({8'd0,data_mid_85_imag} <<< 8);
  assign _zz_14671 = {{8{_zz_14670[23]}}, _zz_14670};
  assign _zz_14672 = fixTo_1425_dout;
  assign _zz_14673 = _zz_14674[31 : 0];
  assign _zz_14674 = _zz_14675;
  assign _zz_14675 = ($signed(_zz_14676) >>> _zz_1190);
  assign _zz_14676 = _zz_14677;
  assign _zz_14677 = ($signed(_zz_14679) + $signed(_zz_1186));
  assign _zz_14678 = ({8'd0,data_mid_85_real} <<< 8);
  assign _zz_14679 = {{8{_zz_14678[23]}}, _zz_14678};
  assign _zz_14680 = fixTo_1426_dout;
  assign _zz_14681 = _zz_14682[31 : 0];
  assign _zz_14682 = _zz_14683;
  assign _zz_14683 = ($signed(_zz_14684) >>> _zz_1190);
  assign _zz_14684 = _zz_14685;
  assign _zz_14685 = ($signed(_zz_14687) + $signed(_zz_1187));
  assign _zz_14686 = ({8'd0,data_mid_85_imag} <<< 8);
  assign _zz_14687 = {{8{_zz_14686[23]}}, _zz_14686};
  assign _zz_14688 = fixTo_1427_dout;
  assign _zz_14689 = ($signed(twiddle_factor_table_13_real) + $signed(twiddle_factor_table_13_imag));
  assign _zz_14690 = ($signed(_zz_1193) - $signed(_zz_14691));
  assign _zz_14691 = ($signed(_zz_14692) * $signed(twiddle_factor_table_13_imag));
  assign _zz_14692 = ($signed(data_mid_94_real) + $signed(data_mid_94_imag));
  assign _zz_14693 = fixTo_1428_dout;
  assign _zz_14694 = ($signed(_zz_1193) + $signed(_zz_14695));
  assign _zz_14695 = ($signed(_zz_14696) * $signed(twiddle_factor_table_13_real));
  assign _zz_14696 = ($signed(data_mid_94_imag) - $signed(data_mid_94_real));
  assign _zz_14697 = fixTo_1429_dout;
  assign _zz_14698 = _zz_14699[31 : 0];
  assign _zz_14699 = _zz_14700;
  assign _zz_14700 = ($signed(_zz_14701) >>> _zz_1194);
  assign _zz_14701 = _zz_14702;
  assign _zz_14702 = ($signed(_zz_14704) - $signed(_zz_1191));
  assign _zz_14703 = ({8'd0,data_mid_86_real} <<< 8);
  assign _zz_14704 = {{8{_zz_14703[23]}}, _zz_14703};
  assign _zz_14705 = fixTo_1430_dout;
  assign _zz_14706 = _zz_14707[31 : 0];
  assign _zz_14707 = _zz_14708;
  assign _zz_14708 = ($signed(_zz_14709) >>> _zz_1194);
  assign _zz_14709 = _zz_14710;
  assign _zz_14710 = ($signed(_zz_14712) - $signed(_zz_1192));
  assign _zz_14711 = ({8'd0,data_mid_86_imag} <<< 8);
  assign _zz_14712 = {{8{_zz_14711[23]}}, _zz_14711};
  assign _zz_14713 = fixTo_1431_dout;
  assign _zz_14714 = _zz_14715[31 : 0];
  assign _zz_14715 = _zz_14716;
  assign _zz_14716 = ($signed(_zz_14717) >>> _zz_1195);
  assign _zz_14717 = _zz_14718;
  assign _zz_14718 = ($signed(_zz_14720) + $signed(_zz_1191));
  assign _zz_14719 = ({8'd0,data_mid_86_real} <<< 8);
  assign _zz_14720 = {{8{_zz_14719[23]}}, _zz_14719};
  assign _zz_14721 = fixTo_1432_dout;
  assign _zz_14722 = _zz_14723[31 : 0];
  assign _zz_14723 = _zz_14724;
  assign _zz_14724 = ($signed(_zz_14725) >>> _zz_1195);
  assign _zz_14725 = _zz_14726;
  assign _zz_14726 = ($signed(_zz_14728) + $signed(_zz_1192));
  assign _zz_14727 = ({8'd0,data_mid_86_imag} <<< 8);
  assign _zz_14728 = {{8{_zz_14727[23]}}, _zz_14727};
  assign _zz_14729 = fixTo_1433_dout;
  assign _zz_14730 = ($signed(twiddle_factor_table_14_real) + $signed(twiddle_factor_table_14_imag));
  assign _zz_14731 = ($signed(_zz_1198) - $signed(_zz_14732));
  assign _zz_14732 = ($signed(_zz_14733) * $signed(twiddle_factor_table_14_imag));
  assign _zz_14733 = ($signed(data_mid_95_real) + $signed(data_mid_95_imag));
  assign _zz_14734 = fixTo_1434_dout;
  assign _zz_14735 = ($signed(_zz_1198) + $signed(_zz_14736));
  assign _zz_14736 = ($signed(_zz_14737) * $signed(twiddle_factor_table_14_real));
  assign _zz_14737 = ($signed(data_mid_95_imag) - $signed(data_mid_95_real));
  assign _zz_14738 = fixTo_1435_dout;
  assign _zz_14739 = _zz_14740[31 : 0];
  assign _zz_14740 = _zz_14741;
  assign _zz_14741 = ($signed(_zz_14742) >>> _zz_1199);
  assign _zz_14742 = _zz_14743;
  assign _zz_14743 = ($signed(_zz_14745) - $signed(_zz_1196));
  assign _zz_14744 = ({8'd0,data_mid_87_real} <<< 8);
  assign _zz_14745 = {{8{_zz_14744[23]}}, _zz_14744};
  assign _zz_14746 = fixTo_1436_dout;
  assign _zz_14747 = _zz_14748[31 : 0];
  assign _zz_14748 = _zz_14749;
  assign _zz_14749 = ($signed(_zz_14750) >>> _zz_1199);
  assign _zz_14750 = _zz_14751;
  assign _zz_14751 = ($signed(_zz_14753) - $signed(_zz_1197));
  assign _zz_14752 = ({8'd0,data_mid_87_imag} <<< 8);
  assign _zz_14753 = {{8{_zz_14752[23]}}, _zz_14752};
  assign _zz_14754 = fixTo_1437_dout;
  assign _zz_14755 = _zz_14756[31 : 0];
  assign _zz_14756 = _zz_14757;
  assign _zz_14757 = ($signed(_zz_14758) >>> _zz_1200);
  assign _zz_14758 = _zz_14759;
  assign _zz_14759 = ($signed(_zz_14761) + $signed(_zz_1196));
  assign _zz_14760 = ({8'd0,data_mid_87_real} <<< 8);
  assign _zz_14761 = {{8{_zz_14760[23]}}, _zz_14760};
  assign _zz_14762 = fixTo_1438_dout;
  assign _zz_14763 = _zz_14764[31 : 0];
  assign _zz_14764 = _zz_14765;
  assign _zz_14765 = ($signed(_zz_14766) >>> _zz_1200);
  assign _zz_14766 = _zz_14767;
  assign _zz_14767 = ($signed(_zz_14769) + $signed(_zz_1197));
  assign _zz_14768 = ({8'd0,data_mid_87_imag} <<< 8);
  assign _zz_14769 = {{8{_zz_14768[23]}}, _zz_14768};
  assign _zz_14770 = fixTo_1439_dout;
  assign _zz_14771 = ($signed(twiddle_factor_table_7_real) + $signed(twiddle_factor_table_7_imag));
  assign _zz_14772 = ($signed(_zz_1203) - $signed(_zz_14773));
  assign _zz_14773 = ($signed(_zz_14774) * $signed(twiddle_factor_table_7_imag));
  assign _zz_14774 = ($signed(data_mid_104_real) + $signed(data_mid_104_imag));
  assign _zz_14775 = fixTo_1440_dout;
  assign _zz_14776 = ($signed(_zz_1203) + $signed(_zz_14777));
  assign _zz_14777 = ($signed(_zz_14778) * $signed(twiddle_factor_table_7_real));
  assign _zz_14778 = ($signed(data_mid_104_imag) - $signed(data_mid_104_real));
  assign _zz_14779 = fixTo_1441_dout;
  assign _zz_14780 = _zz_14781[31 : 0];
  assign _zz_14781 = _zz_14782;
  assign _zz_14782 = ($signed(_zz_14783) >>> _zz_1204);
  assign _zz_14783 = _zz_14784;
  assign _zz_14784 = ($signed(_zz_14786) - $signed(_zz_1201));
  assign _zz_14785 = ({8'd0,data_mid_96_real} <<< 8);
  assign _zz_14786 = {{8{_zz_14785[23]}}, _zz_14785};
  assign _zz_14787 = fixTo_1442_dout;
  assign _zz_14788 = _zz_14789[31 : 0];
  assign _zz_14789 = _zz_14790;
  assign _zz_14790 = ($signed(_zz_14791) >>> _zz_1204);
  assign _zz_14791 = _zz_14792;
  assign _zz_14792 = ($signed(_zz_14794) - $signed(_zz_1202));
  assign _zz_14793 = ({8'd0,data_mid_96_imag} <<< 8);
  assign _zz_14794 = {{8{_zz_14793[23]}}, _zz_14793};
  assign _zz_14795 = fixTo_1443_dout;
  assign _zz_14796 = _zz_14797[31 : 0];
  assign _zz_14797 = _zz_14798;
  assign _zz_14798 = ($signed(_zz_14799) >>> _zz_1205);
  assign _zz_14799 = _zz_14800;
  assign _zz_14800 = ($signed(_zz_14802) + $signed(_zz_1201));
  assign _zz_14801 = ({8'd0,data_mid_96_real} <<< 8);
  assign _zz_14802 = {{8{_zz_14801[23]}}, _zz_14801};
  assign _zz_14803 = fixTo_1444_dout;
  assign _zz_14804 = _zz_14805[31 : 0];
  assign _zz_14805 = _zz_14806;
  assign _zz_14806 = ($signed(_zz_14807) >>> _zz_1205);
  assign _zz_14807 = _zz_14808;
  assign _zz_14808 = ($signed(_zz_14810) + $signed(_zz_1202));
  assign _zz_14809 = ({8'd0,data_mid_96_imag} <<< 8);
  assign _zz_14810 = {{8{_zz_14809[23]}}, _zz_14809};
  assign _zz_14811 = fixTo_1445_dout;
  assign _zz_14812 = ($signed(twiddle_factor_table_8_real) + $signed(twiddle_factor_table_8_imag));
  assign _zz_14813 = ($signed(_zz_1208) - $signed(_zz_14814));
  assign _zz_14814 = ($signed(_zz_14815) * $signed(twiddle_factor_table_8_imag));
  assign _zz_14815 = ($signed(data_mid_105_real) + $signed(data_mid_105_imag));
  assign _zz_14816 = fixTo_1446_dout;
  assign _zz_14817 = ($signed(_zz_1208) + $signed(_zz_14818));
  assign _zz_14818 = ($signed(_zz_14819) * $signed(twiddle_factor_table_8_real));
  assign _zz_14819 = ($signed(data_mid_105_imag) - $signed(data_mid_105_real));
  assign _zz_14820 = fixTo_1447_dout;
  assign _zz_14821 = _zz_14822[31 : 0];
  assign _zz_14822 = _zz_14823;
  assign _zz_14823 = ($signed(_zz_14824) >>> _zz_1209);
  assign _zz_14824 = _zz_14825;
  assign _zz_14825 = ($signed(_zz_14827) - $signed(_zz_1206));
  assign _zz_14826 = ({8'd0,data_mid_97_real} <<< 8);
  assign _zz_14827 = {{8{_zz_14826[23]}}, _zz_14826};
  assign _zz_14828 = fixTo_1448_dout;
  assign _zz_14829 = _zz_14830[31 : 0];
  assign _zz_14830 = _zz_14831;
  assign _zz_14831 = ($signed(_zz_14832) >>> _zz_1209);
  assign _zz_14832 = _zz_14833;
  assign _zz_14833 = ($signed(_zz_14835) - $signed(_zz_1207));
  assign _zz_14834 = ({8'd0,data_mid_97_imag} <<< 8);
  assign _zz_14835 = {{8{_zz_14834[23]}}, _zz_14834};
  assign _zz_14836 = fixTo_1449_dout;
  assign _zz_14837 = _zz_14838[31 : 0];
  assign _zz_14838 = _zz_14839;
  assign _zz_14839 = ($signed(_zz_14840) >>> _zz_1210);
  assign _zz_14840 = _zz_14841;
  assign _zz_14841 = ($signed(_zz_14843) + $signed(_zz_1206));
  assign _zz_14842 = ({8'd0,data_mid_97_real} <<< 8);
  assign _zz_14843 = {{8{_zz_14842[23]}}, _zz_14842};
  assign _zz_14844 = fixTo_1450_dout;
  assign _zz_14845 = _zz_14846[31 : 0];
  assign _zz_14846 = _zz_14847;
  assign _zz_14847 = ($signed(_zz_14848) >>> _zz_1210);
  assign _zz_14848 = _zz_14849;
  assign _zz_14849 = ($signed(_zz_14851) + $signed(_zz_1207));
  assign _zz_14850 = ({8'd0,data_mid_97_imag} <<< 8);
  assign _zz_14851 = {{8{_zz_14850[23]}}, _zz_14850};
  assign _zz_14852 = fixTo_1451_dout;
  assign _zz_14853 = ($signed(twiddle_factor_table_9_real) + $signed(twiddle_factor_table_9_imag));
  assign _zz_14854 = ($signed(_zz_1213) - $signed(_zz_14855));
  assign _zz_14855 = ($signed(_zz_14856) * $signed(twiddle_factor_table_9_imag));
  assign _zz_14856 = ($signed(data_mid_106_real) + $signed(data_mid_106_imag));
  assign _zz_14857 = fixTo_1452_dout;
  assign _zz_14858 = ($signed(_zz_1213) + $signed(_zz_14859));
  assign _zz_14859 = ($signed(_zz_14860) * $signed(twiddle_factor_table_9_real));
  assign _zz_14860 = ($signed(data_mid_106_imag) - $signed(data_mid_106_real));
  assign _zz_14861 = fixTo_1453_dout;
  assign _zz_14862 = _zz_14863[31 : 0];
  assign _zz_14863 = _zz_14864;
  assign _zz_14864 = ($signed(_zz_14865) >>> _zz_1214);
  assign _zz_14865 = _zz_14866;
  assign _zz_14866 = ($signed(_zz_14868) - $signed(_zz_1211));
  assign _zz_14867 = ({8'd0,data_mid_98_real} <<< 8);
  assign _zz_14868 = {{8{_zz_14867[23]}}, _zz_14867};
  assign _zz_14869 = fixTo_1454_dout;
  assign _zz_14870 = _zz_14871[31 : 0];
  assign _zz_14871 = _zz_14872;
  assign _zz_14872 = ($signed(_zz_14873) >>> _zz_1214);
  assign _zz_14873 = _zz_14874;
  assign _zz_14874 = ($signed(_zz_14876) - $signed(_zz_1212));
  assign _zz_14875 = ({8'd0,data_mid_98_imag} <<< 8);
  assign _zz_14876 = {{8{_zz_14875[23]}}, _zz_14875};
  assign _zz_14877 = fixTo_1455_dout;
  assign _zz_14878 = _zz_14879[31 : 0];
  assign _zz_14879 = _zz_14880;
  assign _zz_14880 = ($signed(_zz_14881) >>> _zz_1215);
  assign _zz_14881 = _zz_14882;
  assign _zz_14882 = ($signed(_zz_14884) + $signed(_zz_1211));
  assign _zz_14883 = ({8'd0,data_mid_98_real} <<< 8);
  assign _zz_14884 = {{8{_zz_14883[23]}}, _zz_14883};
  assign _zz_14885 = fixTo_1456_dout;
  assign _zz_14886 = _zz_14887[31 : 0];
  assign _zz_14887 = _zz_14888;
  assign _zz_14888 = ($signed(_zz_14889) >>> _zz_1215);
  assign _zz_14889 = _zz_14890;
  assign _zz_14890 = ($signed(_zz_14892) + $signed(_zz_1212));
  assign _zz_14891 = ({8'd0,data_mid_98_imag} <<< 8);
  assign _zz_14892 = {{8{_zz_14891[23]}}, _zz_14891};
  assign _zz_14893 = fixTo_1457_dout;
  assign _zz_14894 = ($signed(twiddle_factor_table_10_real) + $signed(twiddle_factor_table_10_imag));
  assign _zz_14895 = ($signed(_zz_1218) - $signed(_zz_14896));
  assign _zz_14896 = ($signed(_zz_14897) * $signed(twiddle_factor_table_10_imag));
  assign _zz_14897 = ($signed(data_mid_107_real) + $signed(data_mid_107_imag));
  assign _zz_14898 = fixTo_1458_dout;
  assign _zz_14899 = ($signed(_zz_1218) + $signed(_zz_14900));
  assign _zz_14900 = ($signed(_zz_14901) * $signed(twiddle_factor_table_10_real));
  assign _zz_14901 = ($signed(data_mid_107_imag) - $signed(data_mid_107_real));
  assign _zz_14902 = fixTo_1459_dout;
  assign _zz_14903 = _zz_14904[31 : 0];
  assign _zz_14904 = _zz_14905;
  assign _zz_14905 = ($signed(_zz_14906) >>> _zz_1219);
  assign _zz_14906 = _zz_14907;
  assign _zz_14907 = ($signed(_zz_14909) - $signed(_zz_1216));
  assign _zz_14908 = ({8'd0,data_mid_99_real} <<< 8);
  assign _zz_14909 = {{8{_zz_14908[23]}}, _zz_14908};
  assign _zz_14910 = fixTo_1460_dout;
  assign _zz_14911 = _zz_14912[31 : 0];
  assign _zz_14912 = _zz_14913;
  assign _zz_14913 = ($signed(_zz_14914) >>> _zz_1219);
  assign _zz_14914 = _zz_14915;
  assign _zz_14915 = ($signed(_zz_14917) - $signed(_zz_1217));
  assign _zz_14916 = ({8'd0,data_mid_99_imag} <<< 8);
  assign _zz_14917 = {{8{_zz_14916[23]}}, _zz_14916};
  assign _zz_14918 = fixTo_1461_dout;
  assign _zz_14919 = _zz_14920[31 : 0];
  assign _zz_14920 = _zz_14921;
  assign _zz_14921 = ($signed(_zz_14922) >>> _zz_1220);
  assign _zz_14922 = _zz_14923;
  assign _zz_14923 = ($signed(_zz_14925) + $signed(_zz_1216));
  assign _zz_14924 = ({8'd0,data_mid_99_real} <<< 8);
  assign _zz_14925 = {{8{_zz_14924[23]}}, _zz_14924};
  assign _zz_14926 = fixTo_1462_dout;
  assign _zz_14927 = _zz_14928[31 : 0];
  assign _zz_14928 = _zz_14929;
  assign _zz_14929 = ($signed(_zz_14930) >>> _zz_1220);
  assign _zz_14930 = _zz_14931;
  assign _zz_14931 = ($signed(_zz_14933) + $signed(_zz_1217));
  assign _zz_14932 = ({8'd0,data_mid_99_imag} <<< 8);
  assign _zz_14933 = {{8{_zz_14932[23]}}, _zz_14932};
  assign _zz_14934 = fixTo_1463_dout;
  assign _zz_14935 = ($signed(twiddle_factor_table_11_real) + $signed(twiddle_factor_table_11_imag));
  assign _zz_14936 = ($signed(_zz_1223) - $signed(_zz_14937));
  assign _zz_14937 = ($signed(_zz_14938) * $signed(twiddle_factor_table_11_imag));
  assign _zz_14938 = ($signed(data_mid_108_real) + $signed(data_mid_108_imag));
  assign _zz_14939 = fixTo_1464_dout;
  assign _zz_14940 = ($signed(_zz_1223) + $signed(_zz_14941));
  assign _zz_14941 = ($signed(_zz_14942) * $signed(twiddle_factor_table_11_real));
  assign _zz_14942 = ($signed(data_mid_108_imag) - $signed(data_mid_108_real));
  assign _zz_14943 = fixTo_1465_dout;
  assign _zz_14944 = _zz_14945[31 : 0];
  assign _zz_14945 = _zz_14946;
  assign _zz_14946 = ($signed(_zz_14947) >>> _zz_1224);
  assign _zz_14947 = _zz_14948;
  assign _zz_14948 = ($signed(_zz_14950) - $signed(_zz_1221));
  assign _zz_14949 = ({8'd0,data_mid_100_real} <<< 8);
  assign _zz_14950 = {{8{_zz_14949[23]}}, _zz_14949};
  assign _zz_14951 = fixTo_1466_dout;
  assign _zz_14952 = _zz_14953[31 : 0];
  assign _zz_14953 = _zz_14954;
  assign _zz_14954 = ($signed(_zz_14955) >>> _zz_1224);
  assign _zz_14955 = _zz_14956;
  assign _zz_14956 = ($signed(_zz_14958) - $signed(_zz_1222));
  assign _zz_14957 = ({8'd0,data_mid_100_imag} <<< 8);
  assign _zz_14958 = {{8{_zz_14957[23]}}, _zz_14957};
  assign _zz_14959 = fixTo_1467_dout;
  assign _zz_14960 = _zz_14961[31 : 0];
  assign _zz_14961 = _zz_14962;
  assign _zz_14962 = ($signed(_zz_14963) >>> _zz_1225);
  assign _zz_14963 = _zz_14964;
  assign _zz_14964 = ($signed(_zz_14966) + $signed(_zz_1221));
  assign _zz_14965 = ({8'd0,data_mid_100_real} <<< 8);
  assign _zz_14966 = {{8{_zz_14965[23]}}, _zz_14965};
  assign _zz_14967 = fixTo_1468_dout;
  assign _zz_14968 = _zz_14969[31 : 0];
  assign _zz_14969 = _zz_14970;
  assign _zz_14970 = ($signed(_zz_14971) >>> _zz_1225);
  assign _zz_14971 = _zz_14972;
  assign _zz_14972 = ($signed(_zz_14974) + $signed(_zz_1222));
  assign _zz_14973 = ({8'd0,data_mid_100_imag} <<< 8);
  assign _zz_14974 = {{8{_zz_14973[23]}}, _zz_14973};
  assign _zz_14975 = fixTo_1469_dout;
  assign _zz_14976 = ($signed(twiddle_factor_table_12_real) + $signed(twiddle_factor_table_12_imag));
  assign _zz_14977 = ($signed(_zz_1228) - $signed(_zz_14978));
  assign _zz_14978 = ($signed(_zz_14979) * $signed(twiddle_factor_table_12_imag));
  assign _zz_14979 = ($signed(data_mid_109_real) + $signed(data_mid_109_imag));
  assign _zz_14980 = fixTo_1470_dout;
  assign _zz_14981 = ($signed(_zz_1228) + $signed(_zz_14982));
  assign _zz_14982 = ($signed(_zz_14983) * $signed(twiddle_factor_table_12_real));
  assign _zz_14983 = ($signed(data_mid_109_imag) - $signed(data_mid_109_real));
  assign _zz_14984 = fixTo_1471_dout;
  assign _zz_14985 = _zz_14986[31 : 0];
  assign _zz_14986 = _zz_14987;
  assign _zz_14987 = ($signed(_zz_14988) >>> _zz_1229);
  assign _zz_14988 = _zz_14989;
  assign _zz_14989 = ($signed(_zz_14991) - $signed(_zz_1226));
  assign _zz_14990 = ({8'd0,data_mid_101_real} <<< 8);
  assign _zz_14991 = {{8{_zz_14990[23]}}, _zz_14990};
  assign _zz_14992 = fixTo_1472_dout;
  assign _zz_14993 = _zz_14994[31 : 0];
  assign _zz_14994 = _zz_14995;
  assign _zz_14995 = ($signed(_zz_14996) >>> _zz_1229);
  assign _zz_14996 = _zz_14997;
  assign _zz_14997 = ($signed(_zz_14999) - $signed(_zz_1227));
  assign _zz_14998 = ({8'd0,data_mid_101_imag} <<< 8);
  assign _zz_14999 = {{8{_zz_14998[23]}}, _zz_14998};
  assign _zz_15000 = fixTo_1473_dout;
  assign _zz_15001 = _zz_15002[31 : 0];
  assign _zz_15002 = _zz_15003;
  assign _zz_15003 = ($signed(_zz_15004) >>> _zz_1230);
  assign _zz_15004 = _zz_15005;
  assign _zz_15005 = ($signed(_zz_15007) + $signed(_zz_1226));
  assign _zz_15006 = ({8'd0,data_mid_101_real} <<< 8);
  assign _zz_15007 = {{8{_zz_15006[23]}}, _zz_15006};
  assign _zz_15008 = fixTo_1474_dout;
  assign _zz_15009 = _zz_15010[31 : 0];
  assign _zz_15010 = _zz_15011;
  assign _zz_15011 = ($signed(_zz_15012) >>> _zz_1230);
  assign _zz_15012 = _zz_15013;
  assign _zz_15013 = ($signed(_zz_15015) + $signed(_zz_1227));
  assign _zz_15014 = ({8'd0,data_mid_101_imag} <<< 8);
  assign _zz_15015 = {{8{_zz_15014[23]}}, _zz_15014};
  assign _zz_15016 = fixTo_1475_dout;
  assign _zz_15017 = ($signed(twiddle_factor_table_13_real) + $signed(twiddle_factor_table_13_imag));
  assign _zz_15018 = ($signed(_zz_1233) - $signed(_zz_15019));
  assign _zz_15019 = ($signed(_zz_15020) * $signed(twiddle_factor_table_13_imag));
  assign _zz_15020 = ($signed(data_mid_110_real) + $signed(data_mid_110_imag));
  assign _zz_15021 = fixTo_1476_dout;
  assign _zz_15022 = ($signed(_zz_1233) + $signed(_zz_15023));
  assign _zz_15023 = ($signed(_zz_15024) * $signed(twiddle_factor_table_13_real));
  assign _zz_15024 = ($signed(data_mid_110_imag) - $signed(data_mid_110_real));
  assign _zz_15025 = fixTo_1477_dout;
  assign _zz_15026 = _zz_15027[31 : 0];
  assign _zz_15027 = _zz_15028;
  assign _zz_15028 = ($signed(_zz_15029) >>> _zz_1234);
  assign _zz_15029 = _zz_15030;
  assign _zz_15030 = ($signed(_zz_15032) - $signed(_zz_1231));
  assign _zz_15031 = ({8'd0,data_mid_102_real} <<< 8);
  assign _zz_15032 = {{8{_zz_15031[23]}}, _zz_15031};
  assign _zz_15033 = fixTo_1478_dout;
  assign _zz_15034 = _zz_15035[31 : 0];
  assign _zz_15035 = _zz_15036;
  assign _zz_15036 = ($signed(_zz_15037) >>> _zz_1234);
  assign _zz_15037 = _zz_15038;
  assign _zz_15038 = ($signed(_zz_15040) - $signed(_zz_1232));
  assign _zz_15039 = ({8'd0,data_mid_102_imag} <<< 8);
  assign _zz_15040 = {{8{_zz_15039[23]}}, _zz_15039};
  assign _zz_15041 = fixTo_1479_dout;
  assign _zz_15042 = _zz_15043[31 : 0];
  assign _zz_15043 = _zz_15044;
  assign _zz_15044 = ($signed(_zz_15045) >>> _zz_1235);
  assign _zz_15045 = _zz_15046;
  assign _zz_15046 = ($signed(_zz_15048) + $signed(_zz_1231));
  assign _zz_15047 = ({8'd0,data_mid_102_real} <<< 8);
  assign _zz_15048 = {{8{_zz_15047[23]}}, _zz_15047};
  assign _zz_15049 = fixTo_1480_dout;
  assign _zz_15050 = _zz_15051[31 : 0];
  assign _zz_15051 = _zz_15052;
  assign _zz_15052 = ($signed(_zz_15053) >>> _zz_1235);
  assign _zz_15053 = _zz_15054;
  assign _zz_15054 = ($signed(_zz_15056) + $signed(_zz_1232));
  assign _zz_15055 = ({8'd0,data_mid_102_imag} <<< 8);
  assign _zz_15056 = {{8{_zz_15055[23]}}, _zz_15055};
  assign _zz_15057 = fixTo_1481_dout;
  assign _zz_15058 = ($signed(twiddle_factor_table_14_real) + $signed(twiddle_factor_table_14_imag));
  assign _zz_15059 = ($signed(_zz_1238) - $signed(_zz_15060));
  assign _zz_15060 = ($signed(_zz_15061) * $signed(twiddle_factor_table_14_imag));
  assign _zz_15061 = ($signed(data_mid_111_real) + $signed(data_mid_111_imag));
  assign _zz_15062 = fixTo_1482_dout;
  assign _zz_15063 = ($signed(_zz_1238) + $signed(_zz_15064));
  assign _zz_15064 = ($signed(_zz_15065) * $signed(twiddle_factor_table_14_real));
  assign _zz_15065 = ($signed(data_mid_111_imag) - $signed(data_mid_111_real));
  assign _zz_15066 = fixTo_1483_dout;
  assign _zz_15067 = _zz_15068[31 : 0];
  assign _zz_15068 = _zz_15069;
  assign _zz_15069 = ($signed(_zz_15070) >>> _zz_1239);
  assign _zz_15070 = _zz_15071;
  assign _zz_15071 = ($signed(_zz_15073) - $signed(_zz_1236));
  assign _zz_15072 = ({8'd0,data_mid_103_real} <<< 8);
  assign _zz_15073 = {{8{_zz_15072[23]}}, _zz_15072};
  assign _zz_15074 = fixTo_1484_dout;
  assign _zz_15075 = _zz_15076[31 : 0];
  assign _zz_15076 = _zz_15077;
  assign _zz_15077 = ($signed(_zz_15078) >>> _zz_1239);
  assign _zz_15078 = _zz_15079;
  assign _zz_15079 = ($signed(_zz_15081) - $signed(_zz_1237));
  assign _zz_15080 = ({8'd0,data_mid_103_imag} <<< 8);
  assign _zz_15081 = {{8{_zz_15080[23]}}, _zz_15080};
  assign _zz_15082 = fixTo_1485_dout;
  assign _zz_15083 = _zz_15084[31 : 0];
  assign _zz_15084 = _zz_15085;
  assign _zz_15085 = ($signed(_zz_15086) >>> _zz_1240);
  assign _zz_15086 = _zz_15087;
  assign _zz_15087 = ($signed(_zz_15089) + $signed(_zz_1236));
  assign _zz_15088 = ({8'd0,data_mid_103_real} <<< 8);
  assign _zz_15089 = {{8{_zz_15088[23]}}, _zz_15088};
  assign _zz_15090 = fixTo_1486_dout;
  assign _zz_15091 = _zz_15092[31 : 0];
  assign _zz_15092 = _zz_15093;
  assign _zz_15093 = ($signed(_zz_15094) >>> _zz_1240);
  assign _zz_15094 = _zz_15095;
  assign _zz_15095 = ($signed(_zz_15097) + $signed(_zz_1237));
  assign _zz_15096 = ({8'd0,data_mid_103_imag} <<< 8);
  assign _zz_15097 = {{8{_zz_15096[23]}}, _zz_15096};
  assign _zz_15098 = fixTo_1487_dout;
  assign _zz_15099 = ($signed(twiddle_factor_table_7_real) + $signed(twiddle_factor_table_7_imag));
  assign _zz_15100 = ($signed(_zz_1243) - $signed(_zz_15101));
  assign _zz_15101 = ($signed(_zz_15102) * $signed(twiddle_factor_table_7_imag));
  assign _zz_15102 = ($signed(data_mid_120_real) + $signed(data_mid_120_imag));
  assign _zz_15103 = fixTo_1488_dout;
  assign _zz_15104 = ($signed(_zz_1243) + $signed(_zz_15105));
  assign _zz_15105 = ($signed(_zz_15106) * $signed(twiddle_factor_table_7_real));
  assign _zz_15106 = ($signed(data_mid_120_imag) - $signed(data_mid_120_real));
  assign _zz_15107 = fixTo_1489_dout;
  assign _zz_15108 = _zz_15109[31 : 0];
  assign _zz_15109 = _zz_15110;
  assign _zz_15110 = ($signed(_zz_15111) >>> _zz_1244);
  assign _zz_15111 = _zz_15112;
  assign _zz_15112 = ($signed(_zz_15114) - $signed(_zz_1241));
  assign _zz_15113 = ({8'd0,data_mid_112_real} <<< 8);
  assign _zz_15114 = {{8{_zz_15113[23]}}, _zz_15113};
  assign _zz_15115 = fixTo_1490_dout;
  assign _zz_15116 = _zz_15117[31 : 0];
  assign _zz_15117 = _zz_15118;
  assign _zz_15118 = ($signed(_zz_15119) >>> _zz_1244);
  assign _zz_15119 = _zz_15120;
  assign _zz_15120 = ($signed(_zz_15122) - $signed(_zz_1242));
  assign _zz_15121 = ({8'd0,data_mid_112_imag} <<< 8);
  assign _zz_15122 = {{8{_zz_15121[23]}}, _zz_15121};
  assign _zz_15123 = fixTo_1491_dout;
  assign _zz_15124 = _zz_15125[31 : 0];
  assign _zz_15125 = _zz_15126;
  assign _zz_15126 = ($signed(_zz_15127) >>> _zz_1245);
  assign _zz_15127 = _zz_15128;
  assign _zz_15128 = ($signed(_zz_15130) + $signed(_zz_1241));
  assign _zz_15129 = ({8'd0,data_mid_112_real} <<< 8);
  assign _zz_15130 = {{8{_zz_15129[23]}}, _zz_15129};
  assign _zz_15131 = fixTo_1492_dout;
  assign _zz_15132 = _zz_15133[31 : 0];
  assign _zz_15133 = _zz_15134;
  assign _zz_15134 = ($signed(_zz_15135) >>> _zz_1245);
  assign _zz_15135 = _zz_15136;
  assign _zz_15136 = ($signed(_zz_15138) + $signed(_zz_1242));
  assign _zz_15137 = ({8'd0,data_mid_112_imag} <<< 8);
  assign _zz_15138 = {{8{_zz_15137[23]}}, _zz_15137};
  assign _zz_15139 = fixTo_1493_dout;
  assign _zz_15140 = ($signed(twiddle_factor_table_8_real) + $signed(twiddle_factor_table_8_imag));
  assign _zz_15141 = ($signed(_zz_1248) - $signed(_zz_15142));
  assign _zz_15142 = ($signed(_zz_15143) * $signed(twiddle_factor_table_8_imag));
  assign _zz_15143 = ($signed(data_mid_121_real) + $signed(data_mid_121_imag));
  assign _zz_15144 = fixTo_1494_dout;
  assign _zz_15145 = ($signed(_zz_1248) + $signed(_zz_15146));
  assign _zz_15146 = ($signed(_zz_15147) * $signed(twiddle_factor_table_8_real));
  assign _zz_15147 = ($signed(data_mid_121_imag) - $signed(data_mid_121_real));
  assign _zz_15148 = fixTo_1495_dout;
  assign _zz_15149 = _zz_15150[31 : 0];
  assign _zz_15150 = _zz_15151;
  assign _zz_15151 = ($signed(_zz_15152) >>> _zz_1249);
  assign _zz_15152 = _zz_15153;
  assign _zz_15153 = ($signed(_zz_15155) - $signed(_zz_1246));
  assign _zz_15154 = ({8'd0,data_mid_113_real} <<< 8);
  assign _zz_15155 = {{8{_zz_15154[23]}}, _zz_15154};
  assign _zz_15156 = fixTo_1496_dout;
  assign _zz_15157 = _zz_15158[31 : 0];
  assign _zz_15158 = _zz_15159;
  assign _zz_15159 = ($signed(_zz_15160) >>> _zz_1249);
  assign _zz_15160 = _zz_15161;
  assign _zz_15161 = ($signed(_zz_15163) - $signed(_zz_1247));
  assign _zz_15162 = ({8'd0,data_mid_113_imag} <<< 8);
  assign _zz_15163 = {{8{_zz_15162[23]}}, _zz_15162};
  assign _zz_15164 = fixTo_1497_dout;
  assign _zz_15165 = _zz_15166[31 : 0];
  assign _zz_15166 = _zz_15167;
  assign _zz_15167 = ($signed(_zz_15168) >>> _zz_1250);
  assign _zz_15168 = _zz_15169;
  assign _zz_15169 = ($signed(_zz_15171) + $signed(_zz_1246));
  assign _zz_15170 = ({8'd0,data_mid_113_real} <<< 8);
  assign _zz_15171 = {{8{_zz_15170[23]}}, _zz_15170};
  assign _zz_15172 = fixTo_1498_dout;
  assign _zz_15173 = _zz_15174[31 : 0];
  assign _zz_15174 = _zz_15175;
  assign _zz_15175 = ($signed(_zz_15176) >>> _zz_1250);
  assign _zz_15176 = _zz_15177;
  assign _zz_15177 = ($signed(_zz_15179) + $signed(_zz_1247));
  assign _zz_15178 = ({8'd0,data_mid_113_imag} <<< 8);
  assign _zz_15179 = {{8{_zz_15178[23]}}, _zz_15178};
  assign _zz_15180 = fixTo_1499_dout;
  assign _zz_15181 = ($signed(twiddle_factor_table_9_real) + $signed(twiddle_factor_table_9_imag));
  assign _zz_15182 = ($signed(_zz_1253) - $signed(_zz_15183));
  assign _zz_15183 = ($signed(_zz_15184) * $signed(twiddle_factor_table_9_imag));
  assign _zz_15184 = ($signed(data_mid_122_real) + $signed(data_mid_122_imag));
  assign _zz_15185 = fixTo_1500_dout;
  assign _zz_15186 = ($signed(_zz_1253) + $signed(_zz_15187));
  assign _zz_15187 = ($signed(_zz_15188) * $signed(twiddle_factor_table_9_real));
  assign _zz_15188 = ($signed(data_mid_122_imag) - $signed(data_mid_122_real));
  assign _zz_15189 = fixTo_1501_dout;
  assign _zz_15190 = _zz_15191[31 : 0];
  assign _zz_15191 = _zz_15192;
  assign _zz_15192 = ($signed(_zz_15193) >>> _zz_1254);
  assign _zz_15193 = _zz_15194;
  assign _zz_15194 = ($signed(_zz_15196) - $signed(_zz_1251));
  assign _zz_15195 = ({8'd0,data_mid_114_real} <<< 8);
  assign _zz_15196 = {{8{_zz_15195[23]}}, _zz_15195};
  assign _zz_15197 = fixTo_1502_dout;
  assign _zz_15198 = _zz_15199[31 : 0];
  assign _zz_15199 = _zz_15200;
  assign _zz_15200 = ($signed(_zz_15201) >>> _zz_1254);
  assign _zz_15201 = _zz_15202;
  assign _zz_15202 = ($signed(_zz_15204) - $signed(_zz_1252));
  assign _zz_15203 = ({8'd0,data_mid_114_imag} <<< 8);
  assign _zz_15204 = {{8{_zz_15203[23]}}, _zz_15203};
  assign _zz_15205 = fixTo_1503_dout;
  assign _zz_15206 = _zz_15207[31 : 0];
  assign _zz_15207 = _zz_15208;
  assign _zz_15208 = ($signed(_zz_15209) >>> _zz_1255);
  assign _zz_15209 = _zz_15210;
  assign _zz_15210 = ($signed(_zz_15212) + $signed(_zz_1251));
  assign _zz_15211 = ({8'd0,data_mid_114_real} <<< 8);
  assign _zz_15212 = {{8{_zz_15211[23]}}, _zz_15211};
  assign _zz_15213 = fixTo_1504_dout;
  assign _zz_15214 = _zz_15215[31 : 0];
  assign _zz_15215 = _zz_15216;
  assign _zz_15216 = ($signed(_zz_15217) >>> _zz_1255);
  assign _zz_15217 = _zz_15218;
  assign _zz_15218 = ($signed(_zz_15220) + $signed(_zz_1252));
  assign _zz_15219 = ({8'd0,data_mid_114_imag} <<< 8);
  assign _zz_15220 = {{8{_zz_15219[23]}}, _zz_15219};
  assign _zz_15221 = fixTo_1505_dout;
  assign _zz_15222 = ($signed(twiddle_factor_table_10_real) + $signed(twiddle_factor_table_10_imag));
  assign _zz_15223 = ($signed(_zz_1258) - $signed(_zz_15224));
  assign _zz_15224 = ($signed(_zz_15225) * $signed(twiddle_factor_table_10_imag));
  assign _zz_15225 = ($signed(data_mid_123_real) + $signed(data_mid_123_imag));
  assign _zz_15226 = fixTo_1506_dout;
  assign _zz_15227 = ($signed(_zz_1258) + $signed(_zz_15228));
  assign _zz_15228 = ($signed(_zz_15229) * $signed(twiddle_factor_table_10_real));
  assign _zz_15229 = ($signed(data_mid_123_imag) - $signed(data_mid_123_real));
  assign _zz_15230 = fixTo_1507_dout;
  assign _zz_15231 = _zz_15232[31 : 0];
  assign _zz_15232 = _zz_15233;
  assign _zz_15233 = ($signed(_zz_15234) >>> _zz_1259);
  assign _zz_15234 = _zz_15235;
  assign _zz_15235 = ($signed(_zz_15237) - $signed(_zz_1256));
  assign _zz_15236 = ({8'd0,data_mid_115_real} <<< 8);
  assign _zz_15237 = {{8{_zz_15236[23]}}, _zz_15236};
  assign _zz_15238 = fixTo_1508_dout;
  assign _zz_15239 = _zz_15240[31 : 0];
  assign _zz_15240 = _zz_15241;
  assign _zz_15241 = ($signed(_zz_15242) >>> _zz_1259);
  assign _zz_15242 = _zz_15243;
  assign _zz_15243 = ($signed(_zz_15245) - $signed(_zz_1257));
  assign _zz_15244 = ({8'd0,data_mid_115_imag} <<< 8);
  assign _zz_15245 = {{8{_zz_15244[23]}}, _zz_15244};
  assign _zz_15246 = fixTo_1509_dout;
  assign _zz_15247 = _zz_15248[31 : 0];
  assign _zz_15248 = _zz_15249;
  assign _zz_15249 = ($signed(_zz_15250) >>> _zz_1260);
  assign _zz_15250 = _zz_15251;
  assign _zz_15251 = ($signed(_zz_15253) + $signed(_zz_1256));
  assign _zz_15252 = ({8'd0,data_mid_115_real} <<< 8);
  assign _zz_15253 = {{8{_zz_15252[23]}}, _zz_15252};
  assign _zz_15254 = fixTo_1510_dout;
  assign _zz_15255 = _zz_15256[31 : 0];
  assign _zz_15256 = _zz_15257;
  assign _zz_15257 = ($signed(_zz_15258) >>> _zz_1260);
  assign _zz_15258 = _zz_15259;
  assign _zz_15259 = ($signed(_zz_15261) + $signed(_zz_1257));
  assign _zz_15260 = ({8'd0,data_mid_115_imag} <<< 8);
  assign _zz_15261 = {{8{_zz_15260[23]}}, _zz_15260};
  assign _zz_15262 = fixTo_1511_dout;
  assign _zz_15263 = ($signed(twiddle_factor_table_11_real) + $signed(twiddle_factor_table_11_imag));
  assign _zz_15264 = ($signed(_zz_1263) - $signed(_zz_15265));
  assign _zz_15265 = ($signed(_zz_15266) * $signed(twiddle_factor_table_11_imag));
  assign _zz_15266 = ($signed(data_mid_124_real) + $signed(data_mid_124_imag));
  assign _zz_15267 = fixTo_1512_dout;
  assign _zz_15268 = ($signed(_zz_1263) + $signed(_zz_15269));
  assign _zz_15269 = ($signed(_zz_15270) * $signed(twiddle_factor_table_11_real));
  assign _zz_15270 = ($signed(data_mid_124_imag) - $signed(data_mid_124_real));
  assign _zz_15271 = fixTo_1513_dout;
  assign _zz_15272 = _zz_15273[31 : 0];
  assign _zz_15273 = _zz_15274;
  assign _zz_15274 = ($signed(_zz_15275) >>> _zz_1264);
  assign _zz_15275 = _zz_15276;
  assign _zz_15276 = ($signed(_zz_15278) - $signed(_zz_1261));
  assign _zz_15277 = ({8'd0,data_mid_116_real} <<< 8);
  assign _zz_15278 = {{8{_zz_15277[23]}}, _zz_15277};
  assign _zz_15279 = fixTo_1514_dout;
  assign _zz_15280 = _zz_15281[31 : 0];
  assign _zz_15281 = _zz_15282;
  assign _zz_15282 = ($signed(_zz_15283) >>> _zz_1264);
  assign _zz_15283 = _zz_15284;
  assign _zz_15284 = ($signed(_zz_15286) - $signed(_zz_1262));
  assign _zz_15285 = ({8'd0,data_mid_116_imag} <<< 8);
  assign _zz_15286 = {{8{_zz_15285[23]}}, _zz_15285};
  assign _zz_15287 = fixTo_1515_dout;
  assign _zz_15288 = _zz_15289[31 : 0];
  assign _zz_15289 = _zz_15290;
  assign _zz_15290 = ($signed(_zz_15291) >>> _zz_1265);
  assign _zz_15291 = _zz_15292;
  assign _zz_15292 = ($signed(_zz_15294) + $signed(_zz_1261));
  assign _zz_15293 = ({8'd0,data_mid_116_real} <<< 8);
  assign _zz_15294 = {{8{_zz_15293[23]}}, _zz_15293};
  assign _zz_15295 = fixTo_1516_dout;
  assign _zz_15296 = _zz_15297[31 : 0];
  assign _zz_15297 = _zz_15298;
  assign _zz_15298 = ($signed(_zz_15299) >>> _zz_1265);
  assign _zz_15299 = _zz_15300;
  assign _zz_15300 = ($signed(_zz_15302) + $signed(_zz_1262));
  assign _zz_15301 = ({8'd0,data_mid_116_imag} <<< 8);
  assign _zz_15302 = {{8{_zz_15301[23]}}, _zz_15301};
  assign _zz_15303 = fixTo_1517_dout;
  assign _zz_15304 = ($signed(twiddle_factor_table_12_real) + $signed(twiddle_factor_table_12_imag));
  assign _zz_15305 = ($signed(_zz_1268) - $signed(_zz_15306));
  assign _zz_15306 = ($signed(_zz_15307) * $signed(twiddle_factor_table_12_imag));
  assign _zz_15307 = ($signed(data_mid_125_real) + $signed(data_mid_125_imag));
  assign _zz_15308 = fixTo_1518_dout;
  assign _zz_15309 = ($signed(_zz_1268) + $signed(_zz_15310));
  assign _zz_15310 = ($signed(_zz_15311) * $signed(twiddle_factor_table_12_real));
  assign _zz_15311 = ($signed(data_mid_125_imag) - $signed(data_mid_125_real));
  assign _zz_15312 = fixTo_1519_dout;
  assign _zz_15313 = _zz_15314[31 : 0];
  assign _zz_15314 = _zz_15315;
  assign _zz_15315 = ($signed(_zz_15316) >>> _zz_1269);
  assign _zz_15316 = _zz_15317;
  assign _zz_15317 = ($signed(_zz_15319) - $signed(_zz_1266));
  assign _zz_15318 = ({8'd0,data_mid_117_real} <<< 8);
  assign _zz_15319 = {{8{_zz_15318[23]}}, _zz_15318};
  assign _zz_15320 = fixTo_1520_dout;
  assign _zz_15321 = _zz_15322[31 : 0];
  assign _zz_15322 = _zz_15323;
  assign _zz_15323 = ($signed(_zz_15324) >>> _zz_1269);
  assign _zz_15324 = _zz_15325;
  assign _zz_15325 = ($signed(_zz_15327) - $signed(_zz_1267));
  assign _zz_15326 = ({8'd0,data_mid_117_imag} <<< 8);
  assign _zz_15327 = {{8{_zz_15326[23]}}, _zz_15326};
  assign _zz_15328 = fixTo_1521_dout;
  assign _zz_15329 = _zz_15330[31 : 0];
  assign _zz_15330 = _zz_15331;
  assign _zz_15331 = ($signed(_zz_15332) >>> _zz_1270);
  assign _zz_15332 = _zz_15333;
  assign _zz_15333 = ($signed(_zz_15335) + $signed(_zz_1266));
  assign _zz_15334 = ({8'd0,data_mid_117_real} <<< 8);
  assign _zz_15335 = {{8{_zz_15334[23]}}, _zz_15334};
  assign _zz_15336 = fixTo_1522_dout;
  assign _zz_15337 = _zz_15338[31 : 0];
  assign _zz_15338 = _zz_15339;
  assign _zz_15339 = ($signed(_zz_15340) >>> _zz_1270);
  assign _zz_15340 = _zz_15341;
  assign _zz_15341 = ($signed(_zz_15343) + $signed(_zz_1267));
  assign _zz_15342 = ({8'd0,data_mid_117_imag} <<< 8);
  assign _zz_15343 = {{8{_zz_15342[23]}}, _zz_15342};
  assign _zz_15344 = fixTo_1523_dout;
  assign _zz_15345 = ($signed(twiddle_factor_table_13_real) + $signed(twiddle_factor_table_13_imag));
  assign _zz_15346 = ($signed(_zz_1273) - $signed(_zz_15347));
  assign _zz_15347 = ($signed(_zz_15348) * $signed(twiddle_factor_table_13_imag));
  assign _zz_15348 = ($signed(data_mid_126_real) + $signed(data_mid_126_imag));
  assign _zz_15349 = fixTo_1524_dout;
  assign _zz_15350 = ($signed(_zz_1273) + $signed(_zz_15351));
  assign _zz_15351 = ($signed(_zz_15352) * $signed(twiddle_factor_table_13_real));
  assign _zz_15352 = ($signed(data_mid_126_imag) - $signed(data_mid_126_real));
  assign _zz_15353 = fixTo_1525_dout;
  assign _zz_15354 = _zz_15355[31 : 0];
  assign _zz_15355 = _zz_15356;
  assign _zz_15356 = ($signed(_zz_15357) >>> _zz_1274);
  assign _zz_15357 = _zz_15358;
  assign _zz_15358 = ($signed(_zz_15360) - $signed(_zz_1271));
  assign _zz_15359 = ({8'd0,data_mid_118_real} <<< 8);
  assign _zz_15360 = {{8{_zz_15359[23]}}, _zz_15359};
  assign _zz_15361 = fixTo_1526_dout;
  assign _zz_15362 = _zz_15363[31 : 0];
  assign _zz_15363 = _zz_15364;
  assign _zz_15364 = ($signed(_zz_15365) >>> _zz_1274);
  assign _zz_15365 = _zz_15366;
  assign _zz_15366 = ($signed(_zz_15368) - $signed(_zz_1272));
  assign _zz_15367 = ({8'd0,data_mid_118_imag} <<< 8);
  assign _zz_15368 = {{8{_zz_15367[23]}}, _zz_15367};
  assign _zz_15369 = fixTo_1527_dout;
  assign _zz_15370 = _zz_15371[31 : 0];
  assign _zz_15371 = _zz_15372;
  assign _zz_15372 = ($signed(_zz_15373) >>> _zz_1275);
  assign _zz_15373 = _zz_15374;
  assign _zz_15374 = ($signed(_zz_15376) + $signed(_zz_1271));
  assign _zz_15375 = ({8'd0,data_mid_118_real} <<< 8);
  assign _zz_15376 = {{8{_zz_15375[23]}}, _zz_15375};
  assign _zz_15377 = fixTo_1528_dout;
  assign _zz_15378 = _zz_15379[31 : 0];
  assign _zz_15379 = _zz_15380;
  assign _zz_15380 = ($signed(_zz_15381) >>> _zz_1275);
  assign _zz_15381 = _zz_15382;
  assign _zz_15382 = ($signed(_zz_15384) + $signed(_zz_1272));
  assign _zz_15383 = ({8'd0,data_mid_118_imag} <<< 8);
  assign _zz_15384 = {{8{_zz_15383[23]}}, _zz_15383};
  assign _zz_15385 = fixTo_1529_dout;
  assign _zz_15386 = ($signed(twiddle_factor_table_14_real) + $signed(twiddle_factor_table_14_imag));
  assign _zz_15387 = ($signed(_zz_1278) - $signed(_zz_15388));
  assign _zz_15388 = ($signed(_zz_15389) * $signed(twiddle_factor_table_14_imag));
  assign _zz_15389 = ($signed(data_mid_127_real) + $signed(data_mid_127_imag));
  assign _zz_15390 = fixTo_1530_dout;
  assign _zz_15391 = ($signed(_zz_1278) + $signed(_zz_15392));
  assign _zz_15392 = ($signed(_zz_15393) * $signed(twiddle_factor_table_14_real));
  assign _zz_15393 = ($signed(data_mid_127_imag) - $signed(data_mid_127_real));
  assign _zz_15394 = fixTo_1531_dout;
  assign _zz_15395 = _zz_15396[31 : 0];
  assign _zz_15396 = _zz_15397;
  assign _zz_15397 = ($signed(_zz_15398) >>> _zz_1279);
  assign _zz_15398 = _zz_15399;
  assign _zz_15399 = ($signed(_zz_15401) - $signed(_zz_1276));
  assign _zz_15400 = ({8'd0,data_mid_119_real} <<< 8);
  assign _zz_15401 = {{8{_zz_15400[23]}}, _zz_15400};
  assign _zz_15402 = fixTo_1532_dout;
  assign _zz_15403 = _zz_15404[31 : 0];
  assign _zz_15404 = _zz_15405;
  assign _zz_15405 = ($signed(_zz_15406) >>> _zz_1279);
  assign _zz_15406 = _zz_15407;
  assign _zz_15407 = ($signed(_zz_15409) - $signed(_zz_1277));
  assign _zz_15408 = ({8'd0,data_mid_119_imag} <<< 8);
  assign _zz_15409 = {{8{_zz_15408[23]}}, _zz_15408};
  assign _zz_15410 = fixTo_1533_dout;
  assign _zz_15411 = _zz_15412[31 : 0];
  assign _zz_15412 = _zz_15413;
  assign _zz_15413 = ($signed(_zz_15414) >>> _zz_1280);
  assign _zz_15414 = _zz_15415;
  assign _zz_15415 = ($signed(_zz_15417) + $signed(_zz_1276));
  assign _zz_15416 = ({8'd0,data_mid_119_real} <<< 8);
  assign _zz_15417 = {{8{_zz_15416[23]}}, _zz_15416};
  assign _zz_15418 = fixTo_1534_dout;
  assign _zz_15419 = _zz_15420[31 : 0];
  assign _zz_15420 = _zz_15421;
  assign _zz_15421 = ($signed(_zz_15422) >>> _zz_1280);
  assign _zz_15422 = _zz_15423;
  assign _zz_15423 = ($signed(_zz_15425) + $signed(_zz_1277));
  assign _zz_15424 = ({8'd0,data_mid_119_imag} <<< 8);
  assign _zz_15425 = {{8{_zz_15424[23]}}, _zz_15424};
  assign _zz_15426 = fixTo_1535_dout;
  assign _zz_15427 = ($signed(twiddle_factor_table_15_real) + $signed(twiddle_factor_table_15_imag));
  assign _zz_15428 = ($signed(_zz_1283) - $signed(_zz_15429));
  assign _zz_15429 = ($signed(_zz_15430) * $signed(twiddle_factor_table_15_imag));
  assign _zz_15430 = ($signed(data_mid_16_real) + $signed(data_mid_16_imag));
  assign _zz_15431 = fixTo_1536_dout;
  assign _zz_15432 = ($signed(_zz_1283) + $signed(_zz_15433));
  assign _zz_15433 = ($signed(_zz_15434) * $signed(twiddle_factor_table_15_real));
  assign _zz_15434 = ($signed(data_mid_16_imag) - $signed(data_mid_16_real));
  assign _zz_15435 = fixTo_1537_dout;
  assign _zz_15436 = _zz_15437[31 : 0];
  assign _zz_15437 = _zz_15438;
  assign _zz_15438 = ($signed(_zz_15439) >>> _zz_1284);
  assign _zz_15439 = _zz_15440;
  assign _zz_15440 = ($signed(_zz_15442) - $signed(_zz_1281));
  assign _zz_15441 = ({8'd0,data_mid_0_real} <<< 8);
  assign _zz_15442 = {{8{_zz_15441[23]}}, _zz_15441};
  assign _zz_15443 = fixTo_1538_dout;
  assign _zz_15444 = _zz_15445[31 : 0];
  assign _zz_15445 = _zz_15446;
  assign _zz_15446 = ($signed(_zz_15447) >>> _zz_1284);
  assign _zz_15447 = _zz_15448;
  assign _zz_15448 = ($signed(_zz_15450) - $signed(_zz_1282));
  assign _zz_15449 = ({8'd0,data_mid_0_imag} <<< 8);
  assign _zz_15450 = {{8{_zz_15449[23]}}, _zz_15449};
  assign _zz_15451 = fixTo_1539_dout;
  assign _zz_15452 = _zz_15453[31 : 0];
  assign _zz_15453 = _zz_15454;
  assign _zz_15454 = ($signed(_zz_15455) >>> _zz_1285);
  assign _zz_15455 = _zz_15456;
  assign _zz_15456 = ($signed(_zz_15458) + $signed(_zz_1281));
  assign _zz_15457 = ({8'd0,data_mid_0_real} <<< 8);
  assign _zz_15458 = {{8{_zz_15457[23]}}, _zz_15457};
  assign _zz_15459 = fixTo_1540_dout;
  assign _zz_15460 = _zz_15461[31 : 0];
  assign _zz_15461 = _zz_15462;
  assign _zz_15462 = ($signed(_zz_15463) >>> _zz_1285);
  assign _zz_15463 = _zz_15464;
  assign _zz_15464 = ($signed(_zz_15466) + $signed(_zz_1282));
  assign _zz_15465 = ({8'd0,data_mid_0_imag} <<< 8);
  assign _zz_15466 = {{8{_zz_15465[23]}}, _zz_15465};
  assign _zz_15467 = fixTo_1541_dout;
  assign _zz_15468 = ($signed(twiddle_factor_table_16_real) + $signed(twiddle_factor_table_16_imag));
  assign _zz_15469 = ($signed(_zz_1288) - $signed(_zz_15470));
  assign _zz_15470 = ($signed(_zz_15471) * $signed(twiddle_factor_table_16_imag));
  assign _zz_15471 = ($signed(data_mid_17_real) + $signed(data_mid_17_imag));
  assign _zz_15472 = fixTo_1542_dout;
  assign _zz_15473 = ($signed(_zz_1288) + $signed(_zz_15474));
  assign _zz_15474 = ($signed(_zz_15475) * $signed(twiddle_factor_table_16_real));
  assign _zz_15475 = ($signed(data_mid_17_imag) - $signed(data_mid_17_real));
  assign _zz_15476 = fixTo_1543_dout;
  assign _zz_15477 = _zz_15478[31 : 0];
  assign _zz_15478 = _zz_15479;
  assign _zz_15479 = ($signed(_zz_15480) >>> _zz_1289);
  assign _zz_15480 = _zz_15481;
  assign _zz_15481 = ($signed(_zz_15483) - $signed(_zz_1286));
  assign _zz_15482 = ({8'd0,data_mid_1_real} <<< 8);
  assign _zz_15483 = {{8{_zz_15482[23]}}, _zz_15482};
  assign _zz_15484 = fixTo_1544_dout;
  assign _zz_15485 = _zz_15486[31 : 0];
  assign _zz_15486 = _zz_15487;
  assign _zz_15487 = ($signed(_zz_15488) >>> _zz_1289);
  assign _zz_15488 = _zz_15489;
  assign _zz_15489 = ($signed(_zz_15491) - $signed(_zz_1287));
  assign _zz_15490 = ({8'd0,data_mid_1_imag} <<< 8);
  assign _zz_15491 = {{8{_zz_15490[23]}}, _zz_15490};
  assign _zz_15492 = fixTo_1545_dout;
  assign _zz_15493 = _zz_15494[31 : 0];
  assign _zz_15494 = _zz_15495;
  assign _zz_15495 = ($signed(_zz_15496) >>> _zz_1290);
  assign _zz_15496 = _zz_15497;
  assign _zz_15497 = ($signed(_zz_15499) + $signed(_zz_1286));
  assign _zz_15498 = ({8'd0,data_mid_1_real} <<< 8);
  assign _zz_15499 = {{8{_zz_15498[23]}}, _zz_15498};
  assign _zz_15500 = fixTo_1546_dout;
  assign _zz_15501 = _zz_15502[31 : 0];
  assign _zz_15502 = _zz_15503;
  assign _zz_15503 = ($signed(_zz_15504) >>> _zz_1290);
  assign _zz_15504 = _zz_15505;
  assign _zz_15505 = ($signed(_zz_15507) + $signed(_zz_1287));
  assign _zz_15506 = ({8'd0,data_mid_1_imag} <<< 8);
  assign _zz_15507 = {{8{_zz_15506[23]}}, _zz_15506};
  assign _zz_15508 = fixTo_1547_dout;
  assign _zz_15509 = ($signed(twiddle_factor_table_17_real) + $signed(twiddle_factor_table_17_imag));
  assign _zz_15510 = ($signed(_zz_1293) - $signed(_zz_15511));
  assign _zz_15511 = ($signed(_zz_15512) * $signed(twiddle_factor_table_17_imag));
  assign _zz_15512 = ($signed(data_mid_18_real) + $signed(data_mid_18_imag));
  assign _zz_15513 = fixTo_1548_dout;
  assign _zz_15514 = ($signed(_zz_1293) + $signed(_zz_15515));
  assign _zz_15515 = ($signed(_zz_15516) * $signed(twiddle_factor_table_17_real));
  assign _zz_15516 = ($signed(data_mid_18_imag) - $signed(data_mid_18_real));
  assign _zz_15517 = fixTo_1549_dout;
  assign _zz_15518 = _zz_15519[31 : 0];
  assign _zz_15519 = _zz_15520;
  assign _zz_15520 = ($signed(_zz_15521) >>> _zz_1294);
  assign _zz_15521 = _zz_15522;
  assign _zz_15522 = ($signed(_zz_15524) - $signed(_zz_1291));
  assign _zz_15523 = ({8'd0,data_mid_2_real} <<< 8);
  assign _zz_15524 = {{8{_zz_15523[23]}}, _zz_15523};
  assign _zz_15525 = fixTo_1550_dout;
  assign _zz_15526 = _zz_15527[31 : 0];
  assign _zz_15527 = _zz_15528;
  assign _zz_15528 = ($signed(_zz_15529) >>> _zz_1294);
  assign _zz_15529 = _zz_15530;
  assign _zz_15530 = ($signed(_zz_15532) - $signed(_zz_1292));
  assign _zz_15531 = ({8'd0,data_mid_2_imag} <<< 8);
  assign _zz_15532 = {{8{_zz_15531[23]}}, _zz_15531};
  assign _zz_15533 = fixTo_1551_dout;
  assign _zz_15534 = _zz_15535[31 : 0];
  assign _zz_15535 = _zz_15536;
  assign _zz_15536 = ($signed(_zz_15537) >>> _zz_1295);
  assign _zz_15537 = _zz_15538;
  assign _zz_15538 = ($signed(_zz_15540) + $signed(_zz_1291));
  assign _zz_15539 = ({8'd0,data_mid_2_real} <<< 8);
  assign _zz_15540 = {{8{_zz_15539[23]}}, _zz_15539};
  assign _zz_15541 = fixTo_1552_dout;
  assign _zz_15542 = _zz_15543[31 : 0];
  assign _zz_15543 = _zz_15544;
  assign _zz_15544 = ($signed(_zz_15545) >>> _zz_1295);
  assign _zz_15545 = _zz_15546;
  assign _zz_15546 = ($signed(_zz_15548) + $signed(_zz_1292));
  assign _zz_15547 = ({8'd0,data_mid_2_imag} <<< 8);
  assign _zz_15548 = {{8{_zz_15547[23]}}, _zz_15547};
  assign _zz_15549 = fixTo_1553_dout;
  assign _zz_15550 = ($signed(twiddle_factor_table_18_real) + $signed(twiddle_factor_table_18_imag));
  assign _zz_15551 = ($signed(_zz_1298) - $signed(_zz_15552));
  assign _zz_15552 = ($signed(_zz_15553) * $signed(twiddle_factor_table_18_imag));
  assign _zz_15553 = ($signed(data_mid_19_real) + $signed(data_mid_19_imag));
  assign _zz_15554 = fixTo_1554_dout;
  assign _zz_15555 = ($signed(_zz_1298) + $signed(_zz_15556));
  assign _zz_15556 = ($signed(_zz_15557) * $signed(twiddle_factor_table_18_real));
  assign _zz_15557 = ($signed(data_mid_19_imag) - $signed(data_mid_19_real));
  assign _zz_15558 = fixTo_1555_dout;
  assign _zz_15559 = _zz_15560[31 : 0];
  assign _zz_15560 = _zz_15561;
  assign _zz_15561 = ($signed(_zz_15562) >>> _zz_1299);
  assign _zz_15562 = _zz_15563;
  assign _zz_15563 = ($signed(_zz_15565) - $signed(_zz_1296));
  assign _zz_15564 = ({8'd0,data_mid_3_real} <<< 8);
  assign _zz_15565 = {{8{_zz_15564[23]}}, _zz_15564};
  assign _zz_15566 = fixTo_1556_dout;
  assign _zz_15567 = _zz_15568[31 : 0];
  assign _zz_15568 = _zz_15569;
  assign _zz_15569 = ($signed(_zz_15570) >>> _zz_1299);
  assign _zz_15570 = _zz_15571;
  assign _zz_15571 = ($signed(_zz_15573) - $signed(_zz_1297));
  assign _zz_15572 = ({8'd0,data_mid_3_imag} <<< 8);
  assign _zz_15573 = {{8{_zz_15572[23]}}, _zz_15572};
  assign _zz_15574 = fixTo_1557_dout;
  assign _zz_15575 = _zz_15576[31 : 0];
  assign _zz_15576 = _zz_15577;
  assign _zz_15577 = ($signed(_zz_15578) >>> _zz_1300);
  assign _zz_15578 = _zz_15579;
  assign _zz_15579 = ($signed(_zz_15581) + $signed(_zz_1296));
  assign _zz_15580 = ({8'd0,data_mid_3_real} <<< 8);
  assign _zz_15581 = {{8{_zz_15580[23]}}, _zz_15580};
  assign _zz_15582 = fixTo_1558_dout;
  assign _zz_15583 = _zz_15584[31 : 0];
  assign _zz_15584 = _zz_15585;
  assign _zz_15585 = ($signed(_zz_15586) >>> _zz_1300);
  assign _zz_15586 = _zz_15587;
  assign _zz_15587 = ($signed(_zz_15589) + $signed(_zz_1297));
  assign _zz_15588 = ({8'd0,data_mid_3_imag} <<< 8);
  assign _zz_15589 = {{8{_zz_15588[23]}}, _zz_15588};
  assign _zz_15590 = fixTo_1559_dout;
  assign _zz_15591 = ($signed(twiddle_factor_table_19_real) + $signed(twiddle_factor_table_19_imag));
  assign _zz_15592 = ($signed(_zz_1303) - $signed(_zz_15593));
  assign _zz_15593 = ($signed(_zz_15594) * $signed(twiddle_factor_table_19_imag));
  assign _zz_15594 = ($signed(data_mid_20_real) + $signed(data_mid_20_imag));
  assign _zz_15595 = fixTo_1560_dout;
  assign _zz_15596 = ($signed(_zz_1303) + $signed(_zz_15597));
  assign _zz_15597 = ($signed(_zz_15598) * $signed(twiddle_factor_table_19_real));
  assign _zz_15598 = ($signed(data_mid_20_imag) - $signed(data_mid_20_real));
  assign _zz_15599 = fixTo_1561_dout;
  assign _zz_15600 = _zz_15601[31 : 0];
  assign _zz_15601 = _zz_15602;
  assign _zz_15602 = ($signed(_zz_15603) >>> _zz_1304);
  assign _zz_15603 = _zz_15604;
  assign _zz_15604 = ($signed(_zz_15606) - $signed(_zz_1301));
  assign _zz_15605 = ({8'd0,data_mid_4_real} <<< 8);
  assign _zz_15606 = {{8{_zz_15605[23]}}, _zz_15605};
  assign _zz_15607 = fixTo_1562_dout;
  assign _zz_15608 = _zz_15609[31 : 0];
  assign _zz_15609 = _zz_15610;
  assign _zz_15610 = ($signed(_zz_15611) >>> _zz_1304);
  assign _zz_15611 = _zz_15612;
  assign _zz_15612 = ($signed(_zz_15614) - $signed(_zz_1302));
  assign _zz_15613 = ({8'd0,data_mid_4_imag} <<< 8);
  assign _zz_15614 = {{8{_zz_15613[23]}}, _zz_15613};
  assign _zz_15615 = fixTo_1563_dout;
  assign _zz_15616 = _zz_15617[31 : 0];
  assign _zz_15617 = _zz_15618;
  assign _zz_15618 = ($signed(_zz_15619) >>> _zz_1305);
  assign _zz_15619 = _zz_15620;
  assign _zz_15620 = ($signed(_zz_15622) + $signed(_zz_1301));
  assign _zz_15621 = ({8'd0,data_mid_4_real} <<< 8);
  assign _zz_15622 = {{8{_zz_15621[23]}}, _zz_15621};
  assign _zz_15623 = fixTo_1564_dout;
  assign _zz_15624 = _zz_15625[31 : 0];
  assign _zz_15625 = _zz_15626;
  assign _zz_15626 = ($signed(_zz_15627) >>> _zz_1305);
  assign _zz_15627 = _zz_15628;
  assign _zz_15628 = ($signed(_zz_15630) + $signed(_zz_1302));
  assign _zz_15629 = ({8'd0,data_mid_4_imag} <<< 8);
  assign _zz_15630 = {{8{_zz_15629[23]}}, _zz_15629};
  assign _zz_15631 = fixTo_1565_dout;
  assign _zz_15632 = ($signed(twiddle_factor_table_20_real) + $signed(twiddle_factor_table_20_imag));
  assign _zz_15633 = ($signed(_zz_1308) - $signed(_zz_15634));
  assign _zz_15634 = ($signed(_zz_15635) * $signed(twiddle_factor_table_20_imag));
  assign _zz_15635 = ($signed(data_mid_21_real) + $signed(data_mid_21_imag));
  assign _zz_15636 = fixTo_1566_dout;
  assign _zz_15637 = ($signed(_zz_1308) + $signed(_zz_15638));
  assign _zz_15638 = ($signed(_zz_15639) * $signed(twiddle_factor_table_20_real));
  assign _zz_15639 = ($signed(data_mid_21_imag) - $signed(data_mid_21_real));
  assign _zz_15640 = fixTo_1567_dout;
  assign _zz_15641 = _zz_15642[31 : 0];
  assign _zz_15642 = _zz_15643;
  assign _zz_15643 = ($signed(_zz_15644) >>> _zz_1309);
  assign _zz_15644 = _zz_15645;
  assign _zz_15645 = ($signed(_zz_15647) - $signed(_zz_1306));
  assign _zz_15646 = ({8'd0,data_mid_5_real} <<< 8);
  assign _zz_15647 = {{8{_zz_15646[23]}}, _zz_15646};
  assign _zz_15648 = fixTo_1568_dout;
  assign _zz_15649 = _zz_15650[31 : 0];
  assign _zz_15650 = _zz_15651;
  assign _zz_15651 = ($signed(_zz_15652) >>> _zz_1309);
  assign _zz_15652 = _zz_15653;
  assign _zz_15653 = ($signed(_zz_15655) - $signed(_zz_1307));
  assign _zz_15654 = ({8'd0,data_mid_5_imag} <<< 8);
  assign _zz_15655 = {{8{_zz_15654[23]}}, _zz_15654};
  assign _zz_15656 = fixTo_1569_dout;
  assign _zz_15657 = _zz_15658[31 : 0];
  assign _zz_15658 = _zz_15659;
  assign _zz_15659 = ($signed(_zz_15660) >>> _zz_1310);
  assign _zz_15660 = _zz_15661;
  assign _zz_15661 = ($signed(_zz_15663) + $signed(_zz_1306));
  assign _zz_15662 = ({8'd0,data_mid_5_real} <<< 8);
  assign _zz_15663 = {{8{_zz_15662[23]}}, _zz_15662};
  assign _zz_15664 = fixTo_1570_dout;
  assign _zz_15665 = _zz_15666[31 : 0];
  assign _zz_15666 = _zz_15667;
  assign _zz_15667 = ($signed(_zz_15668) >>> _zz_1310);
  assign _zz_15668 = _zz_15669;
  assign _zz_15669 = ($signed(_zz_15671) + $signed(_zz_1307));
  assign _zz_15670 = ({8'd0,data_mid_5_imag} <<< 8);
  assign _zz_15671 = {{8{_zz_15670[23]}}, _zz_15670};
  assign _zz_15672 = fixTo_1571_dout;
  assign _zz_15673 = ($signed(twiddle_factor_table_21_real) + $signed(twiddle_factor_table_21_imag));
  assign _zz_15674 = ($signed(_zz_1313) - $signed(_zz_15675));
  assign _zz_15675 = ($signed(_zz_15676) * $signed(twiddle_factor_table_21_imag));
  assign _zz_15676 = ($signed(data_mid_22_real) + $signed(data_mid_22_imag));
  assign _zz_15677 = fixTo_1572_dout;
  assign _zz_15678 = ($signed(_zz_1313) + $signed(_zz_15679));
  assign _zz_15679 = ($signed(_zz_15680) * $signed(twiddle_factor_table_21_real));
  assign _zz_15680 = ($signed(data_mid_22_imag) - $signed(data_mid_22_real));
  assign _zz_15681 = fixTo_1573_dout;
  assign _zz_15682 = _zz_15683[31 : 0];
  assign _zz_15683 = _zz_15684;
  assign _zz_15684 = ($signed(_zz_15685) >>> _zz_1314);
  assign _zz_15685 = _zz_15686;
  assign _zz_15686 = ($signed(_zz_15688) - $signed(_zz_1311));
  assign _zz_15687 = ({8'd0,data_mid_6_real} <<< 8);
  assign _zz_15688 = {{8{_zz_15687[23]}}, _zz_15687};
  assign _zz_15689 = fixTo_1574_dout;
  assign _zz_15690 = _zz_15691[31 : 0];
  assign _zz_15691 = _zz_15692;
  assign _zz_15692 = ($signed(_zz_15693) >>> _zz_1314);
  assign _zz_15693 = _zz_15694;
  assign _zz_15694 = ($signed(_zz_15696) - $signed(_zz_1312));
  assign _zz_15695 = ({8'd0,data_mid_6_imag} <<< 8);
  assign _zz_15696 = {{8{_zz_15695[23]}}, _zz_15695};
  assign _zz_15697 = fixTo_1575_dout;
  assign _zz_15698 = _zz_15699[31 : 0];
  assign _zz_15699 = _zz_15700;
  assign _zz_15700 = ($signed(_zz_15701) >>> _zz_1315);
  assign _zz_15701 = _zz_15702;
  assign _zz_15702 = ($signed(_zz_15704) + $signed(_zz_1311));
  assign _zz_15703 = ({8'd0,data_mid_6_real} <<< 8);
  assign _zz_15704 = {{8{_zz_15703[23]}}, _zz_15703};
  assign _zz_15705 = fixTo_1576_dout;
  assign _zz_15706 = _zz_15707[31 : 0];
  assign _zz_15707 = _zz_15708;
  assign _zz_15708 = ($signed(_zz_15709) >>> _zz_1315);
  assign _zz_15709 = _zz_15710;
  assign _zz_15710 = ($signed(_zz_15712) + $signed(_zz_1312));
  assign _zz_15711 = ({8'd0,data_mid_6_imag} <<< 8);
  assign _zz_15712 = {{8{_zz_15711[23]}}, _zz_15711};
  assign _zz_15713 = fixTo_1577_dout;
  assign _zz_15714 = ($signed(twiddle_factor_table_22_real) + $signed(twiddle_factor_table_22_imag));
  assign _zz_15715 = ($signed(_zz_1318) - $signed(_zz_15716));
  assign _zz_15716 = ($signed(_zz_15717) * $signed(twiddle_factor_table_22_imag));
  assign _zz_15717 = ($signed(data_mid_23_real) + $signed(data_mid_23_imag));
  assign _zz_15718 = fixTo_1578_dout;
  assign _zz_15719 = ($signed(_zz_1318) + $signed(_zz_15720));
  assign _zz_15720 = ($signed(_zz_15721) * $signed(twiddle_factor_table_22_real));
  assign _zz_15721 = ($signed(data_mid_23_imag) - $signed(data_mid_23_real));
  assign _zz_15722 = fixTo_1579_dout;
  assign _zz_15723 = _zz_15724[31 : 0];
  assign _zz_15724 = _zz_15725;
  assign _zz_15725 = ($signed(_zz_15726) >>> _zz_1319);
  assign _zz_15726 = _zz_15727;
  assign _zz_15727 = ($signed(_zz_15729) - $signed(_zz_1316));
  assign _zz_15728 = ({8'd0,data_mid_7_real} <<< 8);
  assign _zz_15729 = {{8{_zz_15728[23]}}, _zz_15728};
  assign _zz_15730 = fixTo_1580_dout;
  assign _zz_15731 = _zz_15732[31 : 0];
  assign _zz_15732 = _zz_15733;
  assign _zz_15733 = ($signed(_zz_15734) >>> _zz_1319);
  assign _zz_15734 = _zz_15735;
  assign _zz_15735 = ($signed(_zz_15737) - $signed(_zz_1317));
  assign _zz_15736 = ({8'd0,data_mid_7_imag} <<< 8);
  assign _zz_15737 = {{8{_zz_15736[23]}}, _zz_15736};
  assign _zz_15738 = fixTo_1581_dout;
  assign _zz_15739 = _zz_15740[31 : 0];
  assign _zz_15740 = _zz_15741;
  assign _zz_15741 = ($signed(_zz_15742) >>> _zz_1320);
  assign _zz_15742 = _zz_15743;
  assign _zz_15743 = ($signed(_zz_15745) + $signed(_zz_1316));
  assign _zz_15744 = ({8'd0,data_mid_7_real} <<< 8);
  assign _zz_15745 = {{8{_zz_15744[23]}}, _zz_15744};
  assign _zz_15746 = fixTo_1582_dout;
  assign _zz_15747 = _zz_15748[31 : 0];
  assign _zz_15748 = _zz_15749;
  assign _zz_15749 = ($signed(_zz_15750) >>> _zz_1320);
  assign _zz_15750 = _zz_15751;
  assign _zz_15751 = ($signed(_zz_15753) + $signed(_zz_1317));
  assign _zz_15752 = ({8'd0,data_mid_7_imag} <<< 8);
  assign _zz_15753 = {{8{_zz_15752[23]}}, _zz_15752};
  assign _zz_15754 = fixTo_1583_dout;
  assign _zz_15755 = ($signed(twiddle_factor_table_23_real) + $signed(twiddle_factor_table_23_imag));
  assign _zz_15756 = ($signed(_zz_1323) - $signed(_zz_15757));
  assign _zz_15757 = ($signed(_zz_15758) * $signed(twiddle_factor_table_23_imag));
  assign _zz_15758 = ($signed(data_mid_24_real) + $signed(data_mid_24_imag));
  assign _zz_15759 = fixTo_1584_dout;
  assign _zz_15760 = ($signed(_zz_1323) + $signed(_zz_15761));
  assign _zz_15761 = ($signed(_zz_15762) * $signed(twiddle_factor_table_23_real));
  assign _zz_15762 = ($signed(data_mid_24_imag) - $signed(data_mid_24_real));
  assign _zz_15763 = fixTo_1585_dout;
  assign _zz_15764 = _zz_15765[31 : 0];
  assign _zz_15765 = _zz_15766;
  assign _zz_15766 = ($signed(_zz_15767) >>> _zz_1324);
  assign _zz_15767 = _zz_15768;
  assign _zz_15768 = ($signed(_zz_15770) - $signed(_zz_1321));
  assign _zz_15769 = ({8'd0,data_mid_8_real} <<< 8);
  assign _zz_15770 = {{8{_zz_15769[23]}}, _zz_15769};
  assign _zz_15771 = fixTo_1586_dout;
  assign _zz_15772 = _zz_15773[31 : 0];
  assign _zz_15773 = _zz_15774;
  assign _zz_15774 = ($signed(_zz_15775) >>> _zz_1324);
  assign _zz_15775 = _zz_15776;
  assign _zz_15776 = ($signed(_zz_15778) - $signed(_zz_1322));
  assign _zz_15777 = ({8'd0,data_mid_8_imag} <<< 8);
  assign _zz_15778 = {{8{_zz_15777[23]}}, _zz_15777};
  assign _zz_15779 = fixTo_1587_dout;
  assign _zz_15780 = _zz_15781[31 : 0];
  assign _zz_15781 = _zz_15782;
  assign _zz_15782 = ($signed(_zz_15783) >>> _zz_1325);
  assign _zz_15783 = _zz_15784;
  assign _zz_15784 = ($signed(_zz_15786) + $signed(_zz_1321));
  assign _zz_15785 = ({8'd0,data_mid_8_real} <<< 8);
  assign _zz_15786 = {{8{_zz_15785[23]}}, _zz_15785};
  assign _zz_15787 = fixTo_1588_dout;
  assign _zz_15788 = _zz_15789[31 : 0];
  assign _zz_15789 = _zz_15790;
  assign _zz_15790 = ($signed(_zz_15791) >>> _zz_1325);
  assign _zz_15791 = _zz_15792;
  assign _zz_15792 = ($signed(_zz_15794) + $signed(_zz_1322));
  assign _zz_15793 = ({8'd0,data_mid_8_imag} <<< 8);
  assign _zz_15794 = {{8{_zz_15793[23]}}, _zz_15793};
  assign _zz_15795 = fixTo_1589_dout;
  assign _zz_15796 = ($signed(twiddle_factor_table_24_real) + $signed(twiddle_factor_table_24_imag));
  assign _zz_15797 = ($signed(_zz_1328) - $signed(_zz_15798));
  assign _zz_15798 = ($signed(_zz_15799) * $signed(twiddle_factor_table_24_imag));
  assign _zz_15799 = ($signed(data_mid_25_real) + $signed(data_mid_25_imag));
  assign _zz_15800 = fixTo_1590_dout;
  assign _zz_15801 = ($signed(_zz_1328) + $signed(_zz_15802));
  assign _zz_15802 = ($signed(_zz_15803) * $signed(twiddle_factor_table_24_real));
  assign _zz_15803 = ($signed(data_mid_25_imag) - $signed(data_mid_25_real));
  assign _zz_15804 = fixTo_1591_dout;
  assign _zz_15805 = _zz_15806[31 : 0];
  assign _zz_15806 = _zz_15807;
  assign _zz_15807 = ($signed(_zz_15808) >>> _zz_1329);
  assign _zz_15808 = _zz_15809;
  assign _zz_15809 = ($signed(_zz_15811) - $signed(_zz_1326));
  assign _zz_15810 = ({8'd0,data_mid_9_real} <<< 8);
  assign _zz_15811 = {{8{_zz_15810[23]}}, _zz_15810};
  assign _zz_15812 = fixTo_1592_dout;
  assign _zz_15813 = _zz_15814[31 : 0];
  assign _zz_15814 = _zz_15815;
  assign _zz_15815 = ($signed(_zz_15816) >>> _zz_1329);
  assign _zz_15816 = _zz_15817;
  assign _zz_15817 = ($signed(_zz_15819) - $signed(_zz_1327));
  assign _zz_15818 = ({8'd0,data_mid_9_imag} <<< 8);
  assign _zz_15819 = {{8{_zz_15818[23]}}, _zz_15818};
  assign _zz_15820 = fixTo_1593_dout;
  assign _zz_15821 = _zz_15822[31 : 0];
  assign _zz_15822 = _zz_15823;
  assign _zz_15823 = ($signed(_zz_15824) >>> _zz_1330);
  assign _zz_15824 = _zz_15825;
  assign _zz_15825 = ($signed(_zz_15827) + $signed(_zz_1326));
  assign _zz_15826 = ({8'd0,data_mid_9_real} <<< 8);
  assign _zz_15827 = {{8{_zz_15826[23]}}, _zz_15826};
  assign _zz_15828 = fixTo_1594_dout;
  assign _zz_15829 = _zz_15830[31 : 0];
  assign _zz_15830 = _zz_15831;
  assign _zz_15831 = ($signed(_zz_15832) >>> _zz_1330);
  assign _zz_15832 = _zz_15833;
  assign _zz_15833 = ($signed(_zz_15835) + $signed(_zz_1327));
  assign _zz_15834 = ({8'd0,data_mid_9_imag} <<< 8);
  assign _zz_15835 = {{8{_zz_15834[23]}}, _zz_15834};
  assign _zz_15836 = fixTo_1595_dout;
  assign _zz_15837 = ($signed(twiddle_factor_table_25_real) + $signed(twiddle_factor_table_25_imag));
  assign _zz_15838 = ($signed(_zz_1333) - $signed(_zz_15839));
  assign _zz_15839 = ($signed(_zz_15840) * $signed(twiddle_factor_table_25_imag));
  assign _zz_15840 = ($signed(data_mid_26_real) + $signed(data_mid_26_imag));
  assign _zz_15841 = fixTo_1596_dout;
  assign _zz_15842 = ($signed(_zz_1333) + $signed(_zz_15843));
  assign _zz_15843 = ($signed(_zz_15844) * $signed(twiddle_factor_table_25_real));
  assign _zz_15844 = ($signed(data_mid_26_imag) - $signed(data_mid_26_real));
  assign _zz_15845 = fixTo_1597_dout;
  assign _zz_15846 = _zz_15847[31 : 0];
  assign _zz_15847 = _zz_15848;
  assign _zz_15848 = ($signed(_zz_15849) >>> _zz_1334);
  assign _zz_15849 = _zz_15850;
  assign _zz_15850 = ($signed(_zz_15852) - $signed(_zz_1331));
  assign _zz_15851 = ({8'd0,data_mid_10_real} <<< 8);
  assign _zz_15852 = {{8{_zz_15851[23]}}, _zz_15851};
  assign _zz_15853 = fixTo_1598_dout;
  assign _zz_15854 = _zz_15855[31 : 0];
  assign _zz_15855 = _zz_15856;
  assign _zz_15856 = ($signed(_zz_15857) >>> _zz_1334);
  assign _zz_15857 = _zz_15858;
  assign _zz_15858 = ($signed(_zz_15860) - $signed(_zz_1332));
  assign _zz_15859 = ({8'd0,data_mid_10_imag} <<< 8);
  assign _zz_15860 = {{8{_zz_15859[23]}}, _zz_15859};
  assign _zz_15861 = fixTo_1599_dout;
  assign _zz_15862 = _zz_15863[31 : 0];
  assign _zz_15863 = _zz_15864;
  assign _zz_15864 = ($signed(_zz_15865) >>> _zz_1335);
  assign _zz_15865 = _zz_15866;
  assign _zz_15866 = ($signed(_zz_15868) + $signed(_zz_1331));
  assign _zz_15867 = ({8'd0,data_mid_10_real} <<< 8);
  assign _zz_15868 = {{8{_zz_15867[23]}}, _zz_15867};
  assign _zz_15869 = fixTo_1600_dout;
  assign _zz_15870 = _zz_15871[31 : 0];
  assign _zz_15871 = _zz_15872;
  assign _zz_15872 = ($signed(_zz_15873) >>> _zz_1335);
  assign _zz_15873 = _zz_15874;
  assign _zz_15874 = ($signed(_zz_15876) + $signed(_zz_1332));
  assign _zz_15875 = ({8'd0,data_mid_10_imag} <<< 8);
  assign _zz_15876 = {{8{_zz_15875[23]}}, _zz_15875};
  assign _zz_15877 = fixTo_1601_dout;
  assign _zz_15878 = ($signed(twiddle_factor_table_26_real) + $signed(twiddle_factor_table_26_imag));
  assign _zz_15879 = ($signed(_zz_1338) - $signed(_zz_15880));
  assign _zz_15880 = ($signed(_zz_15881) * $signed(twiddle_factor_table_26_imag));
  assign _zz_15881 = ($signed(data_mid_27_real) + $signed(data_mid_27_imag));
  assign _zz_15882 = fixTo_1602_dout;
  assign _zz_15883 = ($signed(_zz_1338) + $signed(_zz_15884));
  assign _zz_15884 = ($signed(_zz_15885) * $signed(twiddle_factor_table_26_real));
  assign _zz_15885 = ($signed(data_mid_27_imag) - $signed(data_mid_27_real));
  assign _zz_15886 = fixTo_1603_dout;
  assign _zz_15887 = _zz_15888[31 : 0];
  assign _zz_15888 = _zz_15889;
  assign _zz_15889 = ($signed(_zz_15890) >>> _zz_1339);
  assign _zz_15890 = _zz_15891;
  assign _zz_15891 = ($signed(_zz_15893) - $signed(_zz_1336));
  assign _zz_15892 = ({8'd0,data_mid_11_real} <<< 8);
  assign _zz_15893 = {{8{_zz_15892[23]}}, _zz_15892};
  assign _zz_15894 = fixTo_1604_dout;
  assign _zz_15895 = _zz_15896[31 : 0];
  assign _zz_15896 = _zz_15897;
  assign _zz_15897 = ($signed(_zz_15898) >>> _zz_1339);
  assign _zz_15898 = _zz_15899;
  assign _zz_15899 = ($signed(_zz_15901) - $signed(_zz_1337));
  assign _zz_15900 = ({8'd0,data_mid_11_imag} <<< 8);
  assign _zz_15901 = {{8{_zz_15900[23]}}, _zz_15900};
  assign _zz_15902 = fixTo_1605_dout;
  assign _zz_15903 = _zz_15904[31 : 0];
  assign _zz_15904 = _zz_15905;
  assign _zz_15905 = ($signed(_zz_15906) >>> _zz_1340);
  assign _zz_15906 = _zz_15907;
  assign _zz_15907 = ($signed(_zz_15909) + $signed(_zz_1336));
  assign _zz_15908 = ({8'd0,data_mid_11_real} <<< 8);
  assign _zz_15909 = {{8{_zz_15908[23]}}, _zz_15908};
  assign _zz_15910 = fixTo_1606_dout;
  assign _zz_15911 = _zz_15912[31 : 0];
  assign _zz_15912 = _zz_15913;
  assign _zz_15913 = ($signed(_zz_15914) >>> _zz_1340);
  assign _zz_15914 = _zz_15915;
  assign _zz_15915 = ($signed(_zz_15917) + $signed(_zz_1337));
  assign _zz_15916 = ({8'd0,data_mid_11_imag} <<< 8);
  assign _zz_15917 = {{8{_zz_15916[23]}}, _zz_15916};
  assign _zz_15918 = fixTo_1607_dout;
  assign _zz_15919 = ($signed(twiddle_factor_table_27_real) + $signed(twiddle_factor_table_27_imag));
  assign _zz_15920 = ($signed(_zz_1343) - $signed(_zz_15921));
  assign _zz_15921 = ($signed(_zz_15922) * $signed(twiddle_factor_table_27_imag));
  assign _zz_15922 = ($signed(data_mid_28_real) + $signed(data_mid_28_imag));
  assign _zz_15923 = fixTo_1608_dout;
  assign _zz_15924 = ($signed(_zz_1343) + $signed(_zz_15925));
  assign _zz_15925 = ($signed(_zz_15926) * $signed(twiddle_factor_table_27_real));
  assign _zz_15926 = ($signed(data_mid_28_imag) - $signed(data_mid_28_real));
  assign _zz_15927 = fixTo_1609_dout;
  assign _zz_15928 = _zz_15929[31 : 0];
  assign _zz_15929 = _zz_15930;
  assign _zz_15930 = ($signed(_zz_15931) >>> _zz_1344);
  assign _zz_15931 = _zz_15932;
  assign _zz_15932 = ($signed(_zz_15934) - $signed(_zz_1341));
  assign _zz_15933 = ({8'd0,data_mid_12_real} <<< 8);
  assign _zz_15934 = {{8{_zz_15933[23]}}, _zz_15933};
  assign _zz_15935 = fixTo_1610_dout;
  assign _zz_15936 = _zz_15937[31 : 0];
  assign _zz_15937 = _zz_15938;
  assign _zz_15938 = ($signed(_zz_15939) >>> _zz_1344);
  assign _zz_15939 = _zz_15940;
  assign _zz_15940 = ($signed(_zz_15942) - $signed(_zz_1342));
  assign _zz_15941 = ({8'd0,data_mid_12_imag} <<< 8);
  assign _zz_15942 = {{8{_zz_15941[23]}}, _zz_15941};
  assign _zz_15943 = fixTo_1611_dout;
  assign _zz_15944 = _zz_15945[31 : 0];
  assign _zz_15945 = _zz_15946;
  assign _zz_15946 = ($signed(_zz_15947) >>> _zz_1345);
  assign _zz_15947 = _zz_15948;
  assign _zz_15948 = ($signed(_zz_15950) + $signed(_zz_1341));
  assign _zz_15949 = ({8'd0,data_mid_12_real} <<< 8);
  assign _zz_15950 = {{8{_zz_15949[23]}}, _zz_15949};
  assign _zz_15951 = fixTo_1612_dout;
  assign _zz_15952 = _zz_15953[31 : 0];
  assign _zz_15953 = _zz_15954;
  assign _zz_15954 = ($signed(_zz_15955) >>> _zz_1345);
  assign _zz_15955 = _zz_15956;
  assign _zz_15956 = ($signed(_zz_15958) + $signed(_zz_1342));
  assign _zz_15957 = ({8'd0,data_mid_12_imag} <<< 8);
  assign _zz_15958 = {{8{_zz_15957[23]}}, _zz_15957};
  assign _zz_15959 = fixTo_1613_dout;
  assign _zz_15960 = ($signed(twiddle_factor_table_28_real) + $signed(twiddle_factor_table_28_imag));
  assign _zz_15961 = ($signed(_zz_1348) - $signed(_zz_15962));
  assign _zz_15962 = ($signed(_zz_15963) * $signed(twiddle_factor_table_28_imag));
  assign _zz_15963 = ($signed(data_mid_29_real) + $signed(data_mid_29_imag));
  assign _zz_15964 = fixTo_1614_dout;
  assign _zz_15965 = ($signed(_zz_1348) + $signed(_zz_15966));
  assign _zz_15966 = ($signed(_zz_15967) * $signed(twiddle_factor_table_28_real));
  assign _zz_15967 = ($signed(data_mid_29_imag) - $signed(data_mid_29_real));
  assign _zz_15968 = fixTo_1615_dout;
  assign _zz_15969 = _zz_15970[31 : 0];
  assign _zz_15970 = _zz_15971;
  assign _zz_15971 = ($signed(_zz_15972) >>> _zz_1349);
  assign _zz_15972 = _zz_15973;
  assign _zz_15973 = ($signed(_zz_15975) - $signed(_zz_1346));
  assign _zz_15974 = ({8'd0,data_mid_13_real} <<< 8);
  assign _zz_15975 = {{8{_zz_15974[23]}}, _zz_15974};
  assign _zz_15976 = fixTo_1616_dout;
  assign _zz_15977 = _zz_15978[31 : 0];
  assign _zz_15978 = _zz_15979;
  assign _zz_15979 = ($signed(_zz_15980) >>> _zz_1349);
  assign _zz_15980 = _zz_15981;
  assign _zz_15981 = ($signed(_zz_15983) - $signed(_zz_1347));
  assign _zz_15982 = ({8'd0,data_mid_13_imag} <<< 8);
  assign _zz_15983 = {{8{_zz_15982[23]}}, _zz_15982};
  assign _zz_15984 = fixTo_1617_dout;
  assign _zz_15985 = _zz_15986[31 : 0];
  assign _zz_15986 = _zz_15987;
  assign _zz_15987 = ($signed(_zz_15988) >>> _zz_1350);
  assign _zz_15988 = _zz_15989;
  assign _zz_15989 = ($signed(_zz_15991) + $signed(_zz_1346));
  assign _zz_15990 = ({8'd0,data_mid_13_real} <<< 8);
  assign _zz_15991 = {{8{_zz_15990[23]}}, _zz_15990};
  assign _zz_15992 = fixTo_1618_dout;
  assign _zz_15993 = _zz_15994[31 : 0];
  assign _zz_15994 = _zz_15995;
  assign _zz_15995 = ($signed(_zz_15996) >>> _zz_1350);
  assign _zz_15996 = _zz_15997;
  assign _zz_15997 = ($signed(_zz_15999) + $signed(_zz_1347));
  assign _zz_15998 = ({8'd0,data_mid_13_imag} <<< 8);
  assign _zz_15999 = {{8{_zz_15998[23]}}, _zz_15998};
  assign _zz_16000 = fixTo_1619_dout;
  assign _zz_16001 = ($signed(twiddle_factor_table_29_real) + $signed(twiddle_factor_table_29_imag));
  assign _zz_16002 = ($signed(_zz_1353) - $signed(_zz_16003));
  assign _zz_16003 = ($signed(_zz_16004) * $signed(twiddle_factor_table_29_imag));
  assign _zz_16004 = ($signed(data_mid_30_real) + $signed(data_mid_30_imag));
  assign _zz_16005 = fixTo_1620_dout;
  assign _zz_16006 = ($signed(_zz_1353) + $signed(_zz_16007));
  assign _zz_16007 = ($signed(_zz_16008) * $signed(twiddle_factor_table_29_real));
  assign _zz_16008 = ($signed(data_mid_30_imag) - $signed(data_mid_30_real));
  assign _zz_16009 = fixTo_1621_dout;
  assign _zz_16010 = _zz_16011[31 : 0];
  assign _zz_16011 = _zz_16012;
  assign _zz_16012 = ($signed(_zz_16013) >>> _zz_1354);
  assign _zz_16013 = _zz_16014;
  assign _zz_16014 = ($signed(_zz_16016) - $signed(_zz_1351));
  assign _zz_16015 = ({8'd0,data_mid_14_real} <<< 8);
  assign _zz_16016 = {{8{_zz_16015[23]}}, _zz_16015};
  assign _zz_16017 = fixTo_1622_dout;
  assign _zz_16018 = _zz_16019[31 : 0];
  assign _zz_16019 = _zz_16020;
  assign _zz_16020 = ($signed(_zz_16021) >>> _zz_1354);
  assign _zz_16021 = _zz_16022;
  assign _zz_16022 = ($signed(_zz_16024) - $signed(_zz_1352));
  assign _zz_16023 = ({8'd0,data_mid_14_imag} <<< 8);
  assign _zz_16024 = {{8{_zz_16023[23]}}, _zz_16023};
  assign _zz_16025 = fixTo_1623_dout;
  assign _zz_16026 = _zz_16027[31 : 0];
  assign _zz_16027 = _zz_16028;
  assign _zz_16028 = ($signed(_zz_16029) >>> _zz_1355);
  assign _zz_16029 = _zz_16030;
  assign _zz_16030 = ($signed(_zz_16032) + $signed(_zz_1351));
  assign _zz_16031 = ({8'd0,data_mid_14_real} <<< 8);
  assign _zz_16032 = {{8{_zz_16031[23]}}, _zz_16031};
  assign _zz_16033 = fixTo_1624_dout;
  assign _zz_16034 = _zz_16035[31 : 0];
  assign _zz_16035 = _zz_16036;
  assign _zz_16036 = ($signed(_zz_16037) >>> _zz_1355);
  assign _zz_16037 = _zz_16038;
  assign _zz_16038 = ($signed(_zz_16040) + $signed(_zz_1352));
  assign _zz_16039 = ({8'd0,data_mid_14_imag} <<< 8);
  assign _zz_16040 = {{8{_zz_16039[23]}}, _zz_16039};
  assign _zz_16041 = fixTo_1625_dout;
  assign _zz_16042 = ($signed(twiddle_factor_table_30_real) + $signed(twiddle_factor_table_30_imag));
  assign _zz_16043 = ($signed(_zz_1358) - $signed(_zz_16044));
  assign _zz_16044 = ($signed(_zz_16045) * $signed(twiddle_factor_table_30_imag));
  assign _zz_16045 = ($signed(data_mid_31_real) + $signed(data_mid_31_imag));
  assign _zz_16046 = fixTo_1626_dout;
  assign _zz_16047 = ($signed(_zz_1358) + $signed(_zz_16048));
  assign _zz_16048 = ($signed(_zz_16049) * $signed(twiddle_factor_table_30_real));
  assign _zz_16049 = ($signed(data_mid_31_imag) - $signed(data_mid_31_real));
  assign _zz_16050 = fixTo_1627_dout;
  assign _zz_16051 = _zz_16052[31 : 0];
  assign _zz_16052 = _zz_16053;
  assign _zz_16053 = ($signed(_zz_16054) >>> _zz_1359);
  assign _zz_16054 = _zz_16055;
  assign _zz_16055 = ($signed(_zz_16057) - $signed(_zz_1356));
  assign _zz_16056 = ({8'd0,data_mid_15_real} <<< 8);
  assign _zz_16057 = {{8{_zz_16056[23]}}, _zz_16056};
  assign _zz_16058 = fixTo_1628_dout;
  assign _zz_16059 = _zz_16060[31 : 0];
  assign _zz_16060 = _zz_16061;
  assign _zz_16061 = ($signed(_zz_16062) >>> _zz_1359);
  assign _zz_16062 = _zz_16063;
  assign _zz_16063 = ($signed(_zz_16065) - $signed(_zz_1357));
  assign _zz_16064 = ({8'd0,data_mid_15_imag} <<< 8);
  assign _zz_16065 = {{8{_zz_16064[23]}}, _zz_16064};
  assign _zz_16066 = fixTo_1629_dout;
  assign _zz_16067 = _zz_16068[31 : 0];
  assign _zz_16068 = _zz_16069;
  assign _zz_16069 = ($signed(_zz_16070) >>> _zz_1360);
  assign _zz_16070 = _zz_16071;
  assign _zz_16071 = ($signed(_zz_16073) + $signed(_zz_1356));
  assign _zz_16072 = ({8'd0,data_mid_15_real} <<< 8);
  assign _zz_16073 = {{8{_zz_16072[23]}}, _zz_16072};
  assign _zz_16074 = fixTo_1630_dout;
  assign _zz_16075 = _zz_16076[31 : 0];
  assign _zz_16076 = _zz_16077;
  assign _zz_16077 = ($signed(_zz_16078) >>> _zz_1360);
  assign _zz_16078 = _zz_16079;
  assign _zz_16079 = ($signed(_zz_16081) + $signed(_zz_1357));
  assign _zz_16080 = ({8'd0,data_mid_15_imag} <<< 8);
  assign _zz_16081 = {{8{_zz_16080[23]}}, _zz_16080};
  assign _zz_16082 = fixTo_1631_dout;
  assign _zz_16083 = ($signed(twiddle_factor_table_15_real) + $signed(twiddle_factor_table_15_imag));
  assign _zz_16084 = ($signed(_zz_1363) - $signed(_zz_16085));
  assign _zz_16085 = ($signed(_zz_16086) * $signed(twiddle_factor_table_15_imag));
  assign _zz_16086 = ($signed(data_mid_48_real) + $signed(data_mid_48_imag));
  assign _zz_16087 = fixTo_1632_dout;
  assign _zz_16088 = ($signed(_zz_1363) + $signed(_zz_16089));
  assign _zz_16089 = ($signed(_zz_16090) * $signed(twiddle_factor_table_15_real));
  assign _zz_16090 = ($signed(data_mid_48_imag) - $signed(data_mid_48_real));
  assign _zz_16091 = fixTo_1633_dout;
  assign _zz_16092 = _zz_16093[31 : 0];
  assign _zz_16093 = _zz_16094;
  assign _zz_16094 = ($signed(_zz_16095) >>> _zz_1364);
  assign _zz_16095 = _zz_16096;
  assign _zz_16096 = ($signed(_zz_16098) - $signed(_zz_1361));
  assign _zz_16097 = ({8'd0,data_mid_32_real} <<< 8);
  assign _zz_16098 = {{8{_zz_16097[23]}}, _zz_16097};
  assign _zz_16099 = fixTo_1634_dout;
  assign _zz_16100 = _zz_16101[31 : 0];
  assign _zz_16101 = _zz_16102;
  assign _zz_16102 = ($signed(_zz_16103) >>> _zz_1364);
  assign _zz_16103 = _zz_16104;
  assign _zz_16104 = ($signed(_zz_16106) - $signed(_zz_1362));
  assign _zz_16105 = ({8'd0,data_mid_32_imag} <<< 8);
  assign _zz_16106 = {{8{_zz_16105[23]}}, _zz_16105};
  assign _zz_16107 = fixTo_1635_dout;
  assign _zz_16108 = _zz_16109[31 : 0];
  assign _zz_16109 = _zz_16110;
  assign _zz_16110 = ($signed(_zz_16111) >>> _zz_1365);
  assign _zz_16111 = _zz_16112;
  assign _zz_16112 = ($signed(_zz_16114) + $signed(_zz_1361));
  assign _zz_16113 = ({8'd0,data_mid_32_real} <<< 8);
  assign _zz_16114 = {{8{_zz_16113[23]}}, _zz_16113};
  assign _zz_16115 = fixTo_1636_dout;
  assign _zz_16116 = _zz_16117[31 : 0];
  assign _zz_16117 = _zz_16118;
  assign _zz_16118 = ($signed(_zz_16119) >>> _zz_1365);
  assign _zz_16119 = _zz_16120;
  assign _zz_16120 = ($signed(_zz_16122) + $signed(_zz_1362));
  assign _zz_16121 = ({8'd0,data_mid_32_imag} <<< 8);
  assign _zz_16122 = {{8{_zz_16121[23]}}, _zz_16121};
  assign _zz_16123 = fixTo_1637_dout;
  assign _zz_16124 = ($signed(twiddle_factor_table_16_real) + $signed(twiddle_factor_table_16_imag));
  assign _zz_16125 = ($signed(_zz_1368) - $signed(_zz_16126));
  assign _zz_16126 = ($signed(_zz_16127) * $signed(twiddle_factor_table_16_imag));
  assign _zz_16127 = ($signed(data_mid_49_real) + $signed(data_mid_49_imag));
  assign _zz_16128 = fixTo_1638_dout;
  assign _zz_16129 = ($signed(_zz_1368) + $signed(_zz_16130));
  assign _zz_16130 = ($signed(_zz_16131) * $signed(twiddle_factor_table_16_real));
  assign _zz_16131 = ($signed(data_mid_49_imag) - $signed(data_mid_49_real));
  assign _zz_16132 = fixTo_1639_dout;
  assign _zz_16133 = _zz_16134[31 : 0];
  assign _zz_16134 = _zz_16135;
  assign _zz_16135 = ($signed(_zz_16136) >>> _zz_1369);
  assign _zz_16136 = _zz_16137;
  assign _zz_16137 = ($signed(_zz_16139) - $signed(_zz_1366));
  assign _zz_16138 = ({8'd0,data_mid_33_real} <<< 8);
  assign _zz_16139 = {{8{_zz_16138[23]}}, _zz_16138};
  assign _zz_16140 = fixTo_1640_dout;
  assign _zz_16141 = _zz_16142[31 : 0];
  assign _zz_16142 = _zz_16143;
  assign _zz_16143 = ($signed(_zz_16144) >>> _zz_1369);
  assign _zz_16144 = _zz_16145;
  assign _zz_16145 = ($signed(_zz_16147) - $signed(_zz_1367));
  assign _zz_16146 = ({8'd0,data_mid_33_imag} <<< 8);
  assign _zz_16147 = {{8{_zz_16146[23]}}, _zz_16146};
  assign _zz_16148 = fixTo_1641_dout;
  assign _zz_16149 = _zz_16150[31 : 0];
  assign _zz_16150 = _zz_16151;
  assign _zz_16151 = ($signed(_zz_16152) >>> _zz_1370);
  assign _zz_16152 = _zz_16153;
  assign _zz_16153 = ($signed(_zz_16155) + $signed(_zz_1366));
  assign _zz_16154 = ({8'd0,data_mid_33_real} <<< 8);
  assign _zz_16155 = {{8{_zz_16154[23]}}, _zz_16154};
  assign _zz_16156 = fixTo_1642_dout;
  assign _zz_16157 = _zz_16158[31 : 0];
  assign _zz_16158 = _zz_16159;
  assign _zz_16159 = ($signed(_zz_16160) >>> _zz_1370);
  assign _zz_16160 = _zz_16161;
  assign _zz_16161 = ($signed(_zz_16163) + $signed(_zz_1367));
  assign _zz_16162 = ({8'd0,data_mid_33_imag} <<< 8);
  assign _zz_16163 = {{8{_zz_16162[23]}}, _zz_16162};
  assign _zz_16164 = fixTo_1643_dout;
  assign _zz_16165 = ($signed(twiddle_factor_table_17_real) + $signed(twiddle_factor_table_17_imag));
  assign _zz_16166 = ($signed(_zz_1373) - $signed(_zz_16167));
  assign _zz_16167 = ($signed(_zz_16168) * $signed(twiddle_factor_table_17_imag));
  assign _zz_16168 = ($signed(data_mid_50_real) + $signed(data_mid_50_imag));
  assign _zz_16169 = fixTo_1644_dout;
  assign _zz_16170 = ($signed(_zz_1373) + $signed(_zz_16171));
  assign _zz_16171 = ($signed(_zz_16172) * $signed(twiddle_factor_table_17_real));
  assign _zz_16172 = ($signed(data_mid_50_imag) - $signed(data_mid_50_real));
  assign _zz_16173 = fixTo_1645_dout;
  assign _zz_16174 = _zz_16175[31 : 0];
  assign _zz_16175 = _zz_16176;
  assign _zz_16176 = ($signed(_zz_16177) >>> _zz_1374);
  assign _zz_16177 = _zz_16178;
  assign _zz_16178 = ($signed(_zz_16180) - $signed(_zz_1371));
  assign _zz_16179 = ({8'd0,data_mid_34_real} <<< 8);
  assign _zz_16180 = {{8{_zz_16179[23]}}, _zz_16179};
  assign _zz_16181 = fixTo_1646_dout;
  assign _zz_16182 = _zz_16183[31 : 0];
  assign _zz_16183 = _zz_16184;
  assign _zz_16184 = ($signed(_zz_16185) >>> _zz_1374);
  assign _zz_16185 = _zz_16186;
  assign _zz_16186 = ($signed(_zz_16188) - $signed(_zz_1372));
  assign _zz_16187 = ({8'd0,data_mid_34_imag} <<< 8);
  assign _zz_16188 = {{8{_zz_16187[23]}}, _zz_16187};
  assign _zz_16189 = fixTo_1647_dout;
  assign _zz_16190 = _zz_16191[31 : 0];
  assign _zz_16191 = _zz_16192;
  assign _zz_16192 = ($signed(_zz_16193) >>> _zz_1375);
  assign _zz_16193 = _zz_16194;
  assign _zz_16194 = ($signed(_zz_16196) + $signed(_zz_1371));
  assign _zz_16195 = ({8'd0,data_mid_34_real} <<< 8);
  assign _zz_16196 = {{8{_zz_16195[23]}}, _zz_16195};
  assign _zz_16197 = fixTo_1648_dout;
  assign _zz_16198 = _zz_16199[31 : 0];
  assign _zz_16199 = _zz_16200;
  assign _zz_16200 = ($signed(_zz_16201) >>> _zz_1375);
  assign _zz_16201 = _zz_16202;
  assign _zz_16202 = ($signed(_zz_16204) + $signed(_zz_1372));
  assign _zz_16203 = ({8'd0,data_mid_34_imag} <<< 8);
  assign _zz_16204 = {{8{_zz_16203[23]}}, _zz_16203};
  assign _zz_16205 = fixTo_1649_dout;
  assign _zz_16206 = ($signed(twiddle_factor_table_18_real) + $signed(twiddle_factor_table_18_imag));
  assign _zz_16207 = ($signed(_zz_1378) - $signed(_zz_16208));
  assign _zz_16208 = ($signed(_zz_16209) * $signed(twiddle_factor_table_18_imag));
  assign _zz_16209 = ($signed(data_mid_51_real) + $signed(data_mid_51_imag));
  assign _zz_16210 = fixTo_1650_dout;
  assign _zz_16211 = ($signed(_zz_1378) + $signed(_zz_16212));
  assign _zz_16212 = ($signed(_zz_16213) * $signed(twiddle_factor_table_18_real));
  assign _zz_16213 = ($signed(data_mid_51_imag) - $signed(data_mid_51_real));
  assign _zz_16214 = fixTo_1651_dout;
  assign _zz_16215 = _zz_16216[31 : 0];
  assign _zz_16216 = _zz_16217;
  assign _zz_16217 = ($signed(_zz_16218) >>> _zz_1379);
  assign _zz_16218 = _zz_16219;
  assign _zz_16219 = ($signed(_zz_16221) - $signed(_zz_1376));
  assign _zz_16220 = ({8'd0,data_mid_35_real} <<< 8);
  assign _zz_16221 = {{8{_zz_16220[23]}}, _zz_16220};
  assign _zz_16222 = fixTo_1652_dout;
  assign _zz_16223 = _zz_16224[31 : 0];
  assign _zz_16224 = _zz_16225;
  assign _zz_16225 = ($signed(_zz_16226) >>> _zz_1379);
  assign _zz_16226 = _zz_16227;
  assign _zz_16227 = ($signed(_zz_16229) - $signed(_zz_1377));
  assign _zz_16228 = ({8'd0,data_mid_35_imag} <<< 8);
  assign _zz_16229 = {{8{_zz_16228[23]}}, _zz_16228};
  assign _zz_16230 = fixTo_1653_dout;
  assign _zz_16231 = _zz_16232[31 : 0];
  assign _zz_16232 = _zz_16233;
  assign _zz_16233 = ($signed(_zz_16234) >>> _zz_1380);
  assign _zz_16234 = _zz_16235;
  assign _zz_16235 = ($signed(_zz_16237) + $signed(_zz_1376));
  assign _zz_16236 = ({8'd0,data_mid_35_real} <<< 8);
  assign _zz_16237 = {{8{_zz_16236[23]}}, _zz_16236};
  assign _zz_16238 = fixTo_1654_dout;
  assign _zz_16239 = _zz_16240[31 : 0];
  assign _zz_16240 = _zz_16241;
  assign _zz_16241 = ($signed(_zz_16242) >>> _zz_1380);
  assign _zz_16242 = _zz_16243;
  assign _zz_16243 = ($signed(_zz_16245) + $signed(_zz_1377));
  assign _zz_16244 = ({8'd0,data_mid_35_imag} <<< 8);
  assign _zz_16245 = {{8{_zz_16244[23]}}, _zz_16244};
  assign _zz_16246 = fixTo_1655_dout;
  assign _zz_16247 = ($signed(twiddle_factor_table_19_real) + $signed(twiddle_factor_table_19_imag));
  assign _zz_16248 = ($signed(_zz_1383) - $signed(_zz_16249));
  assign _zz_16249 = ($signed(_zz_16250) * $signed(twiddle_factor_table_19_imag));
  assign _zz_16250 = ($signed(data_mid_52_real) + $signed(data_mid_52_imag));
  assign _zz_16251 = fixTo_1656_dout;
  assign _zz_16252 = ($signed(_zz_1383) + $signed(_zz_16253));
  assign _zz_16253 = ($signed(_zz_16254) * $signed(twiddle_factor_table_19_real));
  assign _zz_16254 = ($signed(data_mid_52_imag) - $signed(data_mid_52_real));
  assign _zz_16255 = fixTo_1657_dout;
  assign _zz_16256 = _zz_16257[31 : 0];
  assign _zz_16257 = _zz_16258;
  assign _zz_16258 = ($signed(_zz_16259) >>> _zz_1384);
  assign _zz_16259 = _zz_16260;
  assign _zz_16260 = ($signed(_zz_16262) - $signed(_zz_1381));
  assign _zz_16261 = ({8'd0,data_mid_36_real} <<< 8);
  assign _zz_16262 = {{8{_zz_16261[23]}}, _zz_16261};
  assign _zz_16263 = fixTo_1658_dout;
  assign _zz_16264 = _zz_16265[31 : 0];
  assign _zz_16265 = _zz_16266;
  assign _zz_16266 = ($signed(_zz_16267) >>> _zz_1384);
  assign _zz_16267 = _zz_16268;
  assign _zz_16268 = ($signed(_zz_16270) - $signed(_zz_1382));
  assign _zz_16269 = ({8'd0,data_mid_36_imag} <<< 8);
  assign _zz_16270 = {{8{_zz_16269[23]}}, _zz_16269};
  assign _zz_16271 = fixTo_1659_dout;
  assign _zz_16272 = _zz_16273[31 : 0];
  assign _zz_16273 = _zz_16274;
  assign _zz_16274 = ($signed(_zz_16275) >>> _zz_1385);
  assign _zz_16275 = _zz_16276;
  assign _zz_16276 = ($signed(_zz_16278) + $signed(_zz_1381));
  assign _zz_16277 = ({8'd0,data_mid_36_real} <<< 8);
  assign _zz_16278 = {{8{_zz_16277[23]}}, _zz_16277};
  assign _zz_16279 = fixTo_1660_dout;
  assign _zz_16280 = _zz_16281[31 : 0];
  assign _zz_16281 = _zz_16282;
  assign _zz_16282 = ($signed(_zz_16283) >>> _zz_1385);
  assign _zz_16283 = _zz_16284;
  assign _zz_16284 = ($signed(_zz_16286) + $signed(_zz_1382));
  assign _zz_16285 = ({8'd0,data_mid_36_imag} <<< 8);
  assign _zz_16286 = {{8{_zz_16285[23]}}, _zz_16285};
  assign _zz_16287 = fixTo_1661_dout;
  assign _zz_16288 = ($signed(twiddle_factor_table_20_real) + $signed(twiddle_factor_table_20_imag));
  assign _zz_16289 = ($signed(_zz_1388) - $signed(_zz_16290));
  assign _zz_16290 = ($signed(_zz_16291) * $signed(twiddle_factor_table_20_imag));
  assign _zz_16291 = ($signed(data_mid_53_real) + $signed(data_mid_53_imag));
  assign _zz_16292 = fixTo_1662_dout;
  assign _zz_16293 = ($signed(_zz_1388) + $signed(_zz_16294));
  assign _zz_16294 = ($signed(_zz_16295) * $signed(twiddle_factor_table_20_real));
  assign _zz_16295 = ($signed(data_mid_53_imag) - $signed(data_mid_53_real));
  assign _zz_16296 = fixTo_1663_dout;
  assign _zz_16297 = _zz_16298[31 : 0];
  assign _zz_16298 = _zz_16299;
  assign _zz_16299 = ($signed(_zz_16300) >>> _zz_1389);
  assign _zz_16300 = _zz_16301;
  assign _zz_16301 = ($signed(_zz_16303) - $signed(_zz_1386));
  assign _zz_16302 = ({8'd0,data_mid_37_real} <<< 8);
  assign _zz_16303 = {{8{_zz_16302[23]}}, _zz_16302};
  assign _zz_16304 = fixTo_1664_dout;
  assign _zz_16305 = _zz_16306[31 : 0];
  assign _zz_16306 = _zz_16307;
  assign _zz_16307 = ($signed(_zz_16308) >>> _zz_1389);
  assign _zz_16308 = _zz_16309;
  assign _zz_16309 = ($signed(_zz_16311) - $signed(_zz_1387));
  assign _zz_16310 = ({8'd0,data_mid_37_imag} <<< 8);
  assign _zz_16311 = {{8{_zz_16310[23]}}, _zz_16310};
  assign _zz_16312 = fixTo_1665_dout;
  assign _zz_16313 = _zz_16314[31 : 0];
  assign _zz_16314 = _zz_16315;
  assign _zz_16315 = ($signed(_zz_16316) >>> _zz_1390);
  assign _zz_16316 = _zz_16317;
  assign _zz_16317 = ($signed(_zz_16319) + $signed(_zz_1386));
  assign _zz_16318 = ({8'd0,data_mid_37_real} <<< 8);
  assign _zz_16319 = {{8{_zz_16318[23]}}, _zz_16318};
  assign _zz_16320 = fixTo_1666_dout;
  assign _zz_16321 = _zz_16322[31 : 0];
  assign _zz_16322 = _zz_16323;
  assign _zz_16323 = ($signed(_zz_16324) >>> _zz_1390);
  assign _zz_16324 = _zz_16325;
  assign _zz_16325 = ($signed(_zz_16327) + $signed(_zz_1387));
  assign _zz_16326 = ({8'd0,data_mid_37_imag} <<< 8);
  assign _zz_16327 = {{8{_zz_16326[23]}}, _zz_16326};
  assign _zz_16328 = fixTo_1667_dout;
  assign _zz_16329 = ($signed(twiddle_factor_table_21_real) + $signed(twiddle_factor_table_21_imag));
  assign _zz_16330 = ($signed(_zz_1393) - $signed(_zz_16331));
  assign _zz_16331 = ($signed(_zz_16332) * $signed(twiddle_factor_table_21_imag));
  assign _zz_16332 = ($signed(data_mid_54_real) + $signed(data_mid_54_imag));
  assign _zz_16333 = fixTo_1668_dout;
  assign _zz_16334 = ($signed(_zz_1393) + $signed(_zz_16335));
  assign _zz_16335 = ($signed(_zz_16336) * $signed(twiddle_factor_table_21_real));
  assign _zz_16336 = ($signed(data_mid_54_imag) - $signed(data_mid_54_real));
  assign _zz_16337 = fixTo_1669_dout;
  assign _zz_16338 = _zz_16339[31 : 0];
  assign _zz_16339 = _zz_16340;
  assign _zz_16340 = ($signed(_zz_16341) >>> _zz_1394);
  assign _zz_16341 = _zz_16342;
  assign _zz_16342 = ($signed(_zz_16344) - $signed(_zz_1391));
  assign _zz_16343 = ({8'd0,data_mid_38_real} <<< 8);
  assign _zz_16344 = {{8{_zz_16343[23]}}, _zz_16343};
  assign _zz_16345 = fixTo_1670_dout;
  assign _zz_16346 = _zz_16347[31 : 0];
  assign _zz_16347 = _zz_16348;
  assign _zz_16348 = ($signed(_zz_16349) >>> _zz_1394);
  assign _zz_16349 = _zz_16350;
  assign _zz_16350 = ($signed(_zz_16352) - $signed(_zz_1392));
  assign _zz_16351 = ({8'd0,data_mid_38_imag} <<< 8);
  assign _zz_16352 = {{8{_zz_16351[23]}}, _zz_16351};
  assign _zz_16353 = fixTo_1671_dout;
  assign _zz_16354 = _zz_16355[31 : 0];
  assign _zz_16355 = _zz_16356;
  assign _zz_16356 = ($signed(_zz_16357) >>> _zz_1395);
  assign _zz_16357 = _zz_16358;
  assign _zz_16358 = ($signed(_zz_16360) + $signed(_zz_1391));
  assign _zz_16359 = ({8'd0,data_mid_38_real} <<< 8);
  assign _zz_16360 = {{8{_zz_16359[23]}}, _zz_16359};
  assign _zz_16361 = fixTo_1672_dout;
  assign _zz_16362 = _zz_16363[31 : 0];
  assign _zz_16363 = _zz_16364;
  assign _zz_16364 = ($signed(_zz_16365) >>> _zz_1395);
  assign _zz_16365 = _zz_16366;
  assign _zz_16366 = ($signed(_zz_16368) + $signed(_zz_1392));
  assign _zz_16367 = ({8'd0,data_mid_38_imag} <<< 8);
  assign _zz_16368 = {{8{_zz_16367[23]}}, _zz_16367};
  assign _zz_16369 = fixTo_1673_dout;
  assign _zz_16370 = ($signed(twiddle_factor_table_22_real) + $signed(twiddle_factor_table_22_imag));
  assign _zz_16371 = ($signed(_zz_1398) - $signed(_zz_16372));
  assign _zz_16372 = ($signed(_zz_16373) * $signed(twiddle_factor_table_22_imag));
  assign _zz_16373 = ($signed(data_mid_55_real) + $signed(data_mid_55_imag));
  assign _zz_16374 = fixTo_1674_dout;
  assign _zz_16375 = ($signed(_zz_1398) + $signed(_zz_16376));
  assign _zz_16376 = ($signed(_zz_16377) * $signed(twiddle_factor_table_22_real));
  assign _zz_16377 = ($signed(data_mid_55_imag) - $signed(data_mid_55_real));
  assign _zz_16378 = fixTo_1675_dout;
  assign _zz_16379 = _zz_16380[31 : 0];
  assign _zz_16380 = _zz_16381;
  assign _zz_16381 = ($signed(_zz_16382) >>> _zz_1399);
  assign _zz_16382 = _zz_16383;
  assign _zz_16383 = ($signed(_zz_16385) - $signed(_zz_1396));
  assign _zz_16384 = ({8'd0,data_mid_39_real} <<< 8);
  assign _zz_16385 = {{8{_zz_16384[23]}}, _zz_16384};
  assign _zz_16386 = fixTo_1676_dout;
  assign _zz_16387 = _zz_16388[31 : 0];
  assign _zz_16388 = _zz_16389;
  assign _zz_16389 = ($signed(_zz_16390) >>> _zz_1399);
  assign _zz_16390 = _zz_16391;
  assign _zz_16391 = ($signed(_zz_16393) - $signed(_zz_1397));
  assign _zz_16392 = ({8'd0,data_mid_39_imag} <<< 8);
  assign _zz_16393 = {{8{_zz_16392[23]}}, _zz_16392};
  assign _zz_16394 = fixTo_1677_dout;
  assign _zz_16395 = _zz_16396[31 : 0];
  assign _zz_16396 = _zz_16397;
  assign _zz_16397 = ($signed(_zz_16398) >>> _zz_1400);
  assign _zz_16398 = _zz_16399;
  assign _zz_16399 = ($signed(_zz_16401) + $signed(_zz_1396));
  assign _zz_16400 = ({8'd0,data_mid_39_real} <<< 8);
  assign _zz_16401 = {{8{_zz_16400[23]}}, _zz_16400};
  assign _zz_16402 = fixTo_1678_dout;
  assign _zz_16403 = _zz_16404[31 : 0];
  assign _zz_16404 = _zz_16405;
  assign _zz_16405 = ($signed(_zz_16406) >>> _zz_1400);
  assign _zz_16406 = _zz_16407;
  assign _zz_16407 = ($signed(_zz_16409) + $signed(_zz_1397));
  assign _zz_16408 = ({8'd0,data_mid_39_imag} <<< 8);
  assign _zz_16409 = {{8{_zz_16408[23]}}, _zz_16408};
  assign _zz_16410 = fixTo_1679_dout;
  assign _zz_16411 = ($signed(twiddle_factor_table_23_real) + $signed(twiddle_factor_table_23_imag));
  assign _zz_16412 = ($signed(_zz_1403) - $signed(_zz_16413));
  assign _zz_16413 = ($signed(_zz_16414) * $signed(twiddle_factor_table_23_imag));
  assign _zz_16414 = ($signed(data_mid_56_real) + $signed(data_mid_56_imag));
  assign _zz_16415 = fixTo_1680_dout;
  assign _zz_16416 = ($signed(_zz_1403) + $signed(_zz_16417));
  assign _zz_16417 = ($signed(_zz_16418) * $signed(twiddle_factor_table_23_real));
  assign _zz_16418 = ($signed(data_mid_56_imag) - $signed(data_mid_56_real));
  assign _zz_16419 = fixTo_1681_dout;
  assign _zz_16420 = _zz_16421[31 : 0];
  assign _zz_16421 = _zz_16422;
  assign _zz_16422 = ($signed(_zz_16423) >>> _zz_1404);
  assign _zz_16423 = _zz_16424;
  assign _zz_16424 = ($signed(_zz_16426) - $signed(_zz_1401));
  assign _zz_16425 = ({8'd0,data_mid_40_real} <<< 8);
  assign _zz_16426 = {{8{_zz_16425[23]}}, _zz_16425};
  assign _zz_16427 = fixTo_1682_dout;
  assign _zz_16428 = _zz_16429[31 : 0];
  assign _zz_16429 = _zz_16430;
  assign _zz_16430 = ($signed(_zz_16431) >>> _zz_1404);
  assign _zz_16431 = _zz_16432;
  assign _zz_16432 = ($signed(_zz_16434) - $signed(_zz_1402));
  assign _zz_16433 = ({8'd0,data_mid_40_imag} <<< 8);
  assign _zz_16434 = {{8{_zz_16433[23]}}, _zz_16433};
  assign _zz_16435 = fixTo_1683_dout;
  assign _zz_16436 = _zz_16437[31 : 0];
  assign _zz_16437 = _zz_16438;
  assign _zz_16438 = ($signed(_zz_16439) >>> _zz_1405);
  assign _zz_16439 = _zz_16440;
  assign _zz_16440 = ($signed(_zz_16442) + $signed(_zz_1401));
  assign _zz_16441 = ({8'd0,data_mid_40_real} <<< 8);
  assign _zz_16442 = {{8{_zz_16441[23]}}, _zz_16441};
  assign _zz_16443 = fixTo_1684_dout;
  assign _zz_16444 = _zz_16445[31 : 0];
  assign _zz_16445 = _zz_16446;
  assign _zz_16446 = ($signed(_zz_16447) >>> _zz_1405);
  assign _zz_16447 = _zz_16448;
  assign _zz_16448 = ($signed(_zz_16450) + $signed(_zz_1402));
  assign _zz_16449 = ({8'd0,data_mid_40_imag} <<< 8);
  assign _zz_16450 = {{8{_zz_16449[23]}}, _zz_16449};
  assign _zz_16451 = fixTo_1685_dout;
  assign _zz_16452 = ($signed(twiddle_factor_table_24_real) + $signed(twiddle_factor_table_24_imag));
  assign _zz_16453 = ($signed(_zz_1408) - $signed(_zz_16454));
  assign _zz_16454 = ($signed(_zz_16455) * $signed(twiddle_factor_table_24_imag));
  assign _zz_16455 = ($signed(data_mid_57_real) + $signed(data_mid_57_imag));
  assign _zz_16456 = fixTo_1686_dout;
  assign _zz_16457 = ($signed(_zz_1408) + $signed(_zz_16458));
  assign _zz_16458 = ($signed(_zz_16459) * $signed(twiddle_factor_table_24_real));
  assign _zz_16459 = ($signed(data_mid_57_imag) - $signed(data_mid_57_real));
  assign _zz_16460 = fixTo_1687_dout;
  assign _zz_16461 = _zz_16462[31 : 0];
  assign _zz_16462 = _zz_16463;
  assign _zz_16463 = ($signed(_zz_16464) >>> _zz_1409);
  assign _zz_16464 = _zz_16465;
  assign _zz_16465 = ($signed(_zz_16467) - $signed(_zz_1406));
  assign _zz_16466 = ({8'd0,data_mid_41_real} <<< 8);
  assign _zz_16467 = {{8{_zz_16466[23]}}, _zz_16466};
  assign _zz_16468 = fixTo_1688_dout;
  assign _zz_16469 = _zz_16470[31 : 0];
  assign _zz_16470 = _zz_16471;
  assign _zz_16471 = ($signed(_zz_16472) >>> _zz_1409);
  assign _zz_16472 = _zz_16473;
  assign _zz_16473 = ($signed(_zz_16475) - $signed(_zz_1407));
  assign _zz_16474 = ({8'd0,data_mid_41_imag} <<< 8);
  assign _zz_16475 = {{8{_zz_16474[23]}}, _zz_16474};
  assign _zz_16476 = fixTo_1689_dout;
  assign _zz_16477 = _zz_16478[31 : 0];
  assign _zz_16478 = _zz_16479;
  assign _zz_16479 = ($signed(_zz_16480) >>> _zz_1410);
  assign _zz_16480 = _zz_16481;
  assign _zz_16481 = ($signed(_zz_16483) + $signed(_zz_1406));
  assign _zz_16482 = ({8'd0,data_mid_41_real} <<< 8);
  assign _zz_16483 = {{8{_zz_16482[23]}}, _zz_16482};
  assign _zz_16484 = fixTo_1690_dout;
  assign _zz_16485 = _zz_16486[31 : 0];
  assign _zz_16486 = _zz_16487;
  assign _zz_16487 = ($signed(_zz_16488) >>> _zz_1410);
  assign _zz_16488 = _zz_16489;
  assign _zz_16489 = ($signed(_zz_16491) + $signed(_zz_1407));
  assign _zz_16490 = ({8'd0,data_mid_41_imag} <<< 8);
  assign _zz_16491 = {{8{_zz_16490[23]}}, _zz_16490};
  assign _zz_16492 = fixTo_1691_dout;
  assign _zz_16493 = ($signed(twiddle_factor_table_25_real) + $signed(twiddle_factor_table_25_imag));
  assign _zz_16494 = ($signed(_zz_1413) - $signed(_zz_16495));
  assign _zz_16495 = ($signed(_zz_16496) * $signed(twiddle_factor_table_25_imag));
  assign _zz_16496 = ($signed(data_mid_58_real) + $signed(data_mid_58_imag));
  assign _zz_16497 = fixTo_1692_dout;
  assign _zz_16498 = ($signed(_zz_1413) + $signed(_zz_16499));
  assign _zz_16499 = ($signed(_zz_16500) * $signed(twiddle_factor_table_25_real));
  assign _zz_16500 = ($signed(data_mid_58_imag) - $signed(data_mid_58_real));
  assign _zz_16501 = fixTo_1693_dout;
  assign _zz_16502 = _zz_16503[31 : 0];
  assign _zz_16503 = _zz_16504;
  assign _zz_16504 = ($signed(_zz_16505) >>> _zz_1414);
  assign _zz_16505 = _zz_16506;
  assign _zz_16506 = ($signed(_zz_16508) - $signed(_zz_1411));
  assign _zz_16507 = ({8'd0,data_mid_42_real} <<< 8);
  assign _zz_16508 = {{8{_zz_16507[23]}}, _zz_16507};
  assign _zz_16509 = fixTo_1694_dout;
  assign _zz_16510 = _zz_16511[31 : 0];
  assign _zz_16511 = _zz_16512;
  assign _zz_16512 = ($signed(_zz_16513) >>> _zz_1414);
  assign _zz_16513 = _zz_16514;
  assign _zz_16514 = ($signed(_zz_16516) - $signed(_zz_1412));
  assign _zz_16515 = ({8'd0,data_mid_42_imag} <<< 8);
  assign _zz_16516 = {{8{_zz_16515[23]}}, _zz_16515};
  assign _zz_16517 = fixTo_1695_dout;
  assign _zz_16518 = _zz_16519[31 : 0];
  assign _zz_16519 = _zz_16520;
  assign _zz_16520 = ($signed(_zz_16521) >>> _zz_1415);
  assign _zz_16521 = _zz_16522;
  assign _zz_16522 = ($signed(_zz_16524) + $signed(_zz_1411));
  assign _zz_16523 = ({8'd0,data_mid_42_real} <<< 8);
  assign _zz_16524 = {{8{_zz_16523[23]}}, _zz_16523};
  assign _zz_16525 = fixTo_1696_dout;
  assign _zz_16526 = _zz_16527[31 : 0];
  assign _zz_16527 = _zz_16528;
  assign _zz_16528 = ($signed(_zz_16529) >>> _zz_1415);
  assign _zz_16529 = _zz_16530;
  assign _zz_16530 = ($signed(_zz_16532) + $signed(_zz_1412));
  assign _zz_16531 = ({8'd0,data_mid_42_imag} <<< 8);
  assign _zz_16532 = {{8{_zz_16531[23]}}, _zz_16531};
  assign _zz_16533 = fixTo_1697_dout;
  assign _zz_16534 = ($signed(twiddle_factor_table_26_real) + $signed(twiddle_factor_table_26_imag));
  assign _zz_16535 = ($signed(_zz_1418) - $signed(_zz_16536));
  assign _zz_16536 = ($signed(_zz_16537) * $signed(twiddle_factor_table_26_imag));
  assign _zz_16537 = ($signed(data_mid_59_real) + $signed(data_mid_59_imag));
  assign _zz_16538 = fixTo_1698_dout;
  assign _zz_16539 = ($signed(_zz_1418) + $signed(_zz_16540));
  assign _zz_16540 = ($signed(_zz_16541) * $signed(twiddle_factor_table_26_real));
  assign _zz_16541 = ($signed(data_mid_59_imag) - $signed(data_mid_59_real));
  assign _zz_16542 = fixTo_1699_dout;
  assign _zz_16543 = _zz_16544[31 : 0];
  assign _zz_16544 = _zz_16545;
  assign _zz_16545 = ($signed(_zz_16546) >>> _zz_1419);
  assign _zz_16546 = _zz_16547;
  assign _zz_16547 = ($signed(_zz_16549) - $signed(_zz_1416));
  assign _zz_16548 = ({8'd0,data_mid_43_real} <<< 8);
  assign _zz_16549 = {{8{_zz_16548[23]}}, _zz_16548};
  assign _zz_16550 = fixTo_1700_dout;
  assign _zz_16551 = _zz_16552[31 : 0];
  assign _zz_16552 = _zz_16553;
  assign _zz_16553 = ($signed(_zz_16554) >>> _zz_1419);
  assign _zz_16554 = _zz_16555;
  assign _zz_16555 = ($signed(_zz_16557) - $signed(_zz_1417));
  assign _zz_16556 = ({8'd0,data_mid_43_imag} <<< 8);
  assign _zz_16557 = {{8{_zz_16556[23]}}, _zz_16556};
  assign _zz_16558 = fixTo_1701_dout;
  assign _zz_16559 = _zz_16560[31 : 0];
  assign _zz_16560 = _zz_16561;
  assign _zz_16561 = ($signed(_zz_16562) >>> _zz_1420);
  assign _zz_16562 = _zz_16563;
  assign _zz_16563 = ($signed(_zz_16565) + $signed(_zz_1416));
  assign _zz_16564 = ({8'd0,data_mid_43_real} <<< 8);
  assign _zz_16565 = {{8{_zz_16564[23]}}, _zz_16564};
  assign _zz_16566 = fixTo_1702_dout;
  assign _zz_16567 = _zz_16568[31 : 0];
  assign _zz_16568 = _zz_16569;
  assign _zz_16569 = ($signed(_zz_16570) >>> _zz_1420);
  assign _zz_16570 = _zz_16571;
  assign _zz_16571 = ($signed(_zz_16573) + $signed(_zz_1417));
  assign _zz_16572 = ({8'd0,data_mid_43_imag} <<< 8);
  assign _zz_16573 = {{8{_zz_16572[23]}}, _zz_16572};
  assign _zz_16574 = fixTo_1703_dout;
  assign _zz_16575 = ($signed(twiddle_factor_table_27_real) + $signed(twiddle_factor_table_27_imag));
  assign _zz_16576 = ($signed(_zz_1423) - $signed(_zz_16577));
  assign _zz_16577 = ($signed(_zz_16578) * $signed(twiddle_factor_table_27_imag));
  assign _zz_16578 = ($signed(data_mid_60_real) + $signed(data_mid_60_imag));
  assign _zz_16579 = fixTo_1704_dout;
  assign _zz_16580 = ($signed(_zz_1423) + $signed(_zz_16581));
  assign _zz_16581 = ($signed(_zz_16582) * $signed(twiddle_factor_table_27_real));
  assign _zz_16582 = ($signed(data_mid_60_imag) - $signed(data_mid_60_real));
  assign _zz_16583 = fixTo_1705_dout;
  assign _zz_16584 = _zz_16585[31 : 0];
  assign _zz_16585 = _zz_16586;
  assign _zz_16586 = ($signed(_zz_16587) >>> _zz_1424);
  assign _zz_16587 = _zz_16588;
  assign _zz_16588 = ($signed(_zz_16590) - $signed(_zz_1421));
  assign _zz_16589 = ({8'd0,data_mid_44_real} <<< 8);
  assign _zz_16590 = {{8{_zz_16589[23]}}, _zz_16589};
  assign _zz_16591 = fixTo_1706_dout;
  assign _zz_16592 = _zz_16593[31 : 0];
  assign _zz_16593 = _zz_16594;
  assign _zz_16594 = ($signed(_zz_16595) >>> _zz_1424);
  assign _zz_16595 = _zz_16596;
  assign _zz_16596 = ($signed(_zz_16598) - $signed(_zz_1422));
  assign _zz_16597 = ({8'd0,data_mid_44_imag} <<< 8);
  assign _zz_16598 = {{8{_zz_16597[23]}}, _zz_16597};
  assign _zz_16599 = fixTo_1707_dout;
  assign _zz_16600 = _zz_16601[31 : 0];
  assign _zz_16601 = _zz_16602;
  assign _zz_16602 = ($signed(_zz_16603) >>> _zz_1425);
  assign _zz_16603 = _zz_16604;
  assign _zz_16604 = ($signed(_zz_16606) + $signed(_zz_1421));
  assign _zz_16605 = ({8'd0,data_mid_44_real} <<< 8);
  assign _zz_16606 = {{8{_zz_16605[23]}}, _zz_16605};
  assign _zz_16607 = fixTo_1708_dout;
  assign _zz_16608 = _zz_16609[31 : 0];
  assign _zz_16609 = _zz_16610;
  assign _zz_16610 = ($signed(_zz_16611) >>> _zz_1425);
  assign _zz_16611 = _zz_16612;
  assign _zz_16612 = ($signed(_zz_16614) + $signed(_zz_1422));
  assign _zz_16613 = ({8'd0,data_mid_44_imag} <<< 8);
  assign _zz_16614 = {{8{_zz_16613[23]}}, _zz_16613};
  assign _zz_16615 = fixTo_1709_dout;
  assign _zz_16616 = ($signed(twiddle_factor_table_28_real) + $signed(twiddle_factor_table_28_imag));
  assign _zz_16617 = ($signed(_zz_1428) - $signed(_zz_16618));
  assign _zz_16618 = ($signed(_zz_16619) * $signed(twiddle_factor_table_28_imag));
  assign _zz_16619 = ($signed(data_mid_61_real) + $signed(data_mid_61_imag));
  assign _zz_16620 = fixTo_1710_dout;
  assign _zz_16621 = ($signed(_zz_1428) + $signed(_zz_16622));
  assign _zz_16622 = ($signed(_zz_16623) * $signed(twiddle_factor_table_28_real));
  assign _zz_16623 = ($signed(data_mid_61_imag) - $signed(data_mid_61_real));
  assign _zz_16624 = fixTo_1711_dout;
  assign _zz_16625 = _zz_16626[31 : 0];
  assign _zz_16626 = _zz_16627;
  assign _zz_16627 = ($signed(_zz_16628) >>> _zz_1429);
  assign _zz_16628 = _zz_16629;
  assign _zz_16629 = ($signed(_zz_16631) - $signed(_zz_1426));
  assign _zz_16630 = ({8'd0,data_mid_45_real} <<< 8);
  assign _zz_16631 = {{8{_zz_16630[23]}}, _zz_16630};
  assign _zz_16632 = fixTo_1712_dout;
  assign _zz_16633 = _zz_16634[31 : 0];
  assign _zz_16634 = _zz_16635;
  assign _zz_16635 = ($signed(_zz_16636) >>> _zz_1429);
  assign _zz_16636 = _zz_16637;
  assign _zz_16637 = ($signed(_zz_16639) - $signed(_zz_1427));
  assign _zz_16638 = ({8'd0,data_mid_45_imag} <<< 8);
  assign _zz_16639 = {{8{_zz_16638[23]}}, _zz_16638};
  assign _zz_16640 = fixTo_1713_dout;
  assign _zz_16641 = _zz_16642[31 : 0];
  assign _zz_16642 = _zz_16643;
  assign _zz_16643 = ($signed(_zz_16644) >>> _zz_1430);
  assign _zz_16644 = _zz_16645;
  assign _zz_16645 = ($signed(_zz_16647) + $signed(_zz_1426));
  assign _zz_16646 = ({8'd0,data_mid_45_real} <<< 8);
  assign _zz_16647 = {{8{_zz_16646[23]}}, _zz_16646};
  assign _zz_16648 = fixTo_1714_dout;
  assign _zz_16649 = _zz_16650[31 : 0];
  assign _zz_16650 = _zz_16651;
  assign _zz_16651 = ($signed(_zz_16652) >>> _zz_1430);
  assign _zz_16652 = _zz_16653;
  assign _zz_16653 = ($signed(_zz_16655) + $signed(_zz_1427));
  assign _zz_16654 = ({8'd0,data_mid_45_imag} <<< 8);
  assign _zz_16655 = {{8{_zz_16654[23]}}, _zz_16654};
  assign _zz_16656 = fixTo_1715_dout;
  assign _zz_16657 = ($signed(twiddle_factor_table_29_real) + $signed(twiddle_factor_table_29_imag));
  assign _zz_16658 = ($signed(_zz_1433) - $signed(_zz_16659));
  assign _zz_16659 = ($signed(_zz_16660) * $signed(twiddle_factor_table_29_imag));
  assign _zz_16660 = ($signed(data_mid_62_real) + $signed(data_mid_62_imag));
  assign _zz_16661 = fixTo_1716_dout;
  assign _zz_16662 = ($signed(_zz_1433) + $signed(_zz_16663));
  assign _zz_16663 = ($signed(_zz_16664) * $signed(twiddle_factor_table_29_real));
  assign _zz_16664 = ($signed(data_mid_62_imag) - $signed(data_mid_62_real));
  assign _zz_16665 = fixTo_1717_dout;
  assign _zz_16666 = _zz_16667[31 : 0];
  assign _zz_16667 = _zz_16668;
  assign _zz_16668 = ($signed(_zz_16669) >>> _zz_1434);
  assign _zz_16669 = _zz_16670;
  assign _zz_16670 = ($signed(_zz_16672) - $signed(_zz_1431));
  assign _zz_16671 = ({8'd0,data_mid_46_real} <<< 8);
  assign _zz_16672 = {{8{_zz_16671[23]}}, _zz_16671};
  assign _zz_16673 = fixTo_1718_dout;
  assign _zz_16674 = _zz_16675[31 : 0];
  assign _zz_16675 = _zz_16676;
  assign _zz_16676 = ($signed(_zz_16677) >>> _zz_1434);
  assign _zz_16677 = _zz_16678;
  assign _zz_16678 = ($signed(_zz_16680) - $signed(_zz_1432));
  assign _zz_16679 = ({8'd0,data_mid_46_imag} <<< 8);
  assign _zz_16680 = {{8{_zz_16679[23]}}, _zz_16679};
  assign _zz_16681 = fixTo_1719_dout;
  assign _zz_16682 = _zz_16683[31 : 0];
  assign _zz_16683 = _zz_16684;
  assign _zz_16684 = ($signed(_zz_16685) >>> _zz_1435);
  assign _zz_16685 = _zz_16686;
  assign _zz_16686 = ($signed(_zz_16688) + $signed(_zz_1431));
  assign _zz_16687 = ({8'd0,data_mid_46_real} <<< 8);
  assign _zz_16688 = {{8{_zz_16687[23]}}, _zz_16687};
  assign _zz_16689 = fixTo_1720_dout;
  assign _zz_16690 = _zz_16691[31 : 0];
  assign _zz_16691 = _zz_16692;
  assign _zz_16692 = ($signed(_zz_16693) >>> _zz_1435);
  assign _zz_16693 = _zz_16694;
  assign _zz_16694 = ($signed(_zz_16696) + $signed(_zz_1432));
  assign _zz_16695 = ({8'd0,data_mid_46_imag} <<< 8);
  assign _zz_16696 = {{8{_zz_16695[23]}}, _zz_16695};
  assign _zz_16697 = fixTo_1721_dout;
  assign _zz_16698 = ($signed(twiddle_factor_table_30_real) + $signed(twiddle_factor_table_30_imag));
  assign _zz_16699 = ($signed(_zz_1438) - $signed(_zz_16700));
  assign _zz_16700 = ($signed(_zz_16701) * $signed(twiddle_factor_table_30_imag));
  assign _zz_16701 = ($signed(data_mid_63_real) + $signed(data_mid_63_imag));
  assign _zz_16702 = fixTo_1722_dout;
  assign _zz_16703 = ($signed(_zz_1438) + $signed(_zz_16704));
  assign _zz_16704 = ($signed(_zz_16705) * $signed(twiddle_factor_table_30_real));
  assign _zz_16705 = ($signed(data_mid_63_imag) - $signed(data_mid_63_real));
  assign _zz_16706 = fixTo_1723_dout;
  assign _zz_16707 = _zz_16708[31 : 0];
  assign _zz_16708 = _zz_16709;
  assign _zz_16709 = ($signed(_zz_16710) >>> _zz_1439);
  assign _zz_16710 = _zz_16711;
  assign _zz_16711 = ($signed(_zz_16713) - $signed(_zz_1436));
  assign _zz_16712 = ({8'd0,data_mid_47_real} <<< 8);
  assign _zz_16713 = {{8{_zz_16712[23]}}, _zz_16712};
  assign _zz_16714 = fixTo_1724_dout;
  assign _zz_16715 = _zz_16716[31 : 0];
  assign _zz_16716 = _zz_16717;
  assign _zz_16717 = ($signed(_zz_16718) >>> _zz_1439);
  assign _zz_16718 = _zz_16719;
  assign _zz_16719 = ($signed(_zz_16721) - $signed(_zz_1437));
  assign _zz_16720 = ({8'd0,data_mid_47_imag} <<< 8);
  assign _zz_16721 = {{8{_zz_16720[23]}}, _zz_16720};
  assign _zz_16722 = fixTo_1725_dout;
  assign _zz_16723 = _zz_16724[31 : 0];
  assign _zz_16724 = _zz_16725;
  assign _zz_16725 = ($signed(_zz_16726) >>> _zz_1440);
  assign _zz_16726 = _zz_16727;
  assign _zz_16727 = ($signed(_zz_16729) + $signed(_zz_1436));
  assign _zz_16728 = ({8'd0,data_mid_47_real} <<< 8);
  assign _zz_16729 = {{8{_zz_16728[23]}}, _zz_16728};
  assign _zz_16730 = fixTo_1726_dout;
  assign _zz_16731 = _zz_16732[31 : 0];
  assign _zz_16732 = _zz_16733;
  assign _zz_16733 = ($signed(_zz_16734) >>> _zz_1440);
  assign _zz_16734 = _zz_16735;
  assign _zz_16735 = ($signed(_zz_16737) + $signed(_zz_1437));
  assign _zz_16736 = ({8'd0,data_mid_47_imag} <<< 8);
  assign _zz_16737 = {{8{_zz_16736[23]}}, _zz_16736};
  assign _zz_16738 = fixTo_1727_dout;
  assign _zz_16739 = ($signed(twiddle_factor_table_15_real) + $signed(twiddle_factor_table_15_imag));
  assign _zz_16740 = ($signed(_zz_1443) - $signed(_zz_16741));
  assign _zz_16741 = ($signed(_zz_16742) * $signed(twiddle_factor_table_15_imag));
  assign _zz_16742 = ($signed(data_mid_80_real) + $signed(data_mid_80_imag));
  assign _zz_16743 = fixTo_1728_dout;
  assign _zz_16744 = ($signed(_zz_1443) + $signed(_zz_16745));
  assign _zz_16745 = ($signed(_zz_16746) * $signed(twiddle_factor_table_15_real));
  assign _zz_16746 = ($signed(data_mid_80_imag) - $signed(data_mid_80_real));
  assign _zz_16747 = fixTo_1729_dout;
  assign _zz_16748 = _zz_16749[31 : 0];
  assign _zz_16749 = _zz_16750;
  assign _zz_16750 = ($signed(_zz_16751) >>> _zz_1444);
  assign _zz_16751 = _zz_16752;
  assign _zz_16752 = ($signed(_zz_16754) - $signed(_zz_1441));
  assign _zz_16753 = ({8'd0,data_mid_64_real} <<< 8);
  assign _zz_16754 = {{8{_zz_16753[23]}}, _zz_16753};
  assign _zz_16755 = fixTo_1730_dout;
  assign _zz_16756 = _zz_16757[31 : 0];
  assign _zz_16757 = _zz_16758;
  assign _zz_16758 = ($signed(_zz_16759) >>> _zz_1444);
  assign _zz_16759 = _zz_16760;
  assign _zz_16760 = ($signed(_zz_16762) - $signed(_zz_1442));
  assign _zz_16761 = ({8'd0,data_mid_64_imag} <<< 8);
  assign _zz_16762 = {{8{_zz_16761[23]}}, _zz_16761};
  assign _zz_16763 = fixTo_1731_dout;
  assign _zz_16764 = _zz_16765[31 : 0];
  assign _zz_16765 = _zz_16766;
  assign _zz_16766 = ($signed(_zz_16767) >>> _zz_1445);
  assign _zz_16767 = _zz_16768;
  assign _zz_16768 = ($signed(_zz_16770) + $signed(_zz_1441));
  assign _zz_16769 = ({8'd0,data_mid_64_real} <<< 8);
  assign _zz_16770 = {{8{_zz_16769[23]}}, _zz_16769};
  assign _zz_16771 = fixTo_1732_dout;
  assign _zz_16772 = _zz_16773[31 : 0];
  assign _zz_16773 = _zz_16774;
  assign _zz_16774 = ($signed(_zz_16775) >>> _zz_1445);
  assign _zz_16775 = _zz_16776;
  assign _zz_16776 = ($signed(_zz_16778) + $signed(_zz_1442));
  assign _zz_16777 = ({8'd0,data_mid_64_imag} <<< 8);
  assign _zz_16778 = {{8{_zz_16777[23]}}, _zz_16777};
  assign _zz_16779 = fixTo_1733_dout;
  assign _zz_16780 = ($signed(twiddle_factor_table_16_real) + $signed(twiddle_factor_table_16_imag));
  assign _zz_16781 = ($signed(_zz_1448) - $signed(_zz_16782));
  assign _zz_16782 = ($signed(_zz_16783) * $signed(twiddle_factor_table_16_imag));
  assign _zz_16783 = ($signed(data_mid_81_real) + $signed(data_mid_81_imag));
  assign _zz_16784 = fixTo_1734_dout;
  assign _zz_16785 = ($signed(_zz_1448) + $signed(_zz_16786));
  assign _zz_16786 = ($signed(_zz_16787) * $signed(twiddle_factor_table_16_real));
  assign _zz_16787 = ($signed(data_mid_81_imag) - $signed(data_mid_81_real));
  assign _zz_16788 = fixTo_1735_dout;
  assign _zz_16789 = _zz_16790[31 : 0];
  assign _zz_16790 = _zz_16791;
  assign _zz_16791 = ($signed(_zz_16792) >>> _zz_1449);
  assign _zz_16792 = _zz_16793;
  assign _zz_16793 = ($signed(_zz_16795) - $signed(_zz_1446));
  assign _zz_16794 = ({8'd0,data_mid_65_real} <<< 8);
  assign _zz_16795 = {{8{_zz_16794[23]}}, _zz_16794};
  assign _zz_16796 = fixTo_1736_dout;
  assign _zz_16797 = _zz_16798[31 : 0];
  assign _zz_16798 = _zz_16799;
  assign _zz_16799 = ($signed(_zz_16800) >>> _zz_1449);
  assign _zz_16800 = _zz_16801;
  assign _zz_16801 = ($signed(_zz_16803) - $signed(_zz_1447));
  assign _zz_16802 = ({8'd0,data_mid_65_imag} <<< 8);
  assign _zz_16803 = {{8{_zz_16802[23]}}, _zz_16802};
  assign _zz_16804 = fixTo_1737_dout;
  assign _zz_16805 = _zz_16806[31 : 0];
  assign _zz_16806 = _zz_16807;
  assign _zz_16807 = ($signed(_zz_16808) >>> _zz_1450);
  assign _zz_16808 = _zz_16809;
  assign _zz_16809 = ($signed(_zz_16811) + $signed(_zz_1446));
  assign _zz_16810 = ({8'd0,data_mid_65_real} <<< 8);
  assign _zz_16811 = {{8{_zz_16810[23]}}, _zz_16810};
  assign _zz_16812 = fixTo_1738_dout;
  assign _zz_16813 = _zz_16814[31 : 0];
  assign _zz_16814 = _zz_16815;
  assign _zz_16815 = ($signed(_zz_16816) >>> _zz_1450);
  assign _zz_16816 = _zz_16817;
  assign _zz_16817 = ($signed(_zz_16819) + $signed(_zz_1447));
  assign _zz_16818 = ({8'd0,data_mid_65_imag} <<< 8);
  assign _zz_16819 = {{8{_zz_16818[23]}}, _zz_16818};
  assign _zz_16820 = fixTo_1739_dout;
  assign _zz_16821 = ($signed(twiddle_factor_table_17_real) + $signed(twiddle_factor_table_17_imag));
  assign _zz_16822 = ($signed(_zz_1453) - $signed(_zz_16823));
  assign _zz_16823 = ($signed(_zz_16824) * $signed(twiddle_factor_table_17_imag));
  assign _zz_16824 = ($signed(data_mid_82_real) + $signed(data_mid_82_imag));
  assign _zz_16825 = fixTo_1740_dout;
  assign _zz_16826 = ($signed(_zz_1453) + $signed(_zz_16827));
  assign _zz_16827 = ($signed(_zz_16828) * $signed(twiddle_factor_table_17_real));
  assign _zz_16828 = ($signed(data_mid_82_imag) - $signed(data_mid_82_real));
  assign _zz_16829 = fixTo_1741_dout;
  assign _zz_16830 = _zz_16831[31 : 0];
  assign _zz_16831 = _zz_16832;
  assign _zz_16832 = ($signed(_zz_16833) >>> _zz_1454);
  assign _zz_16833 = _zz_16834;
  assign _zz_16834 = ($signed(_zz_16836) - $signed(_zz_1451));
  assign _zz_16835 = ({8'd0,data_mid_66_real} <<< 8);
  assign _zz_16836 = {{8{_zz_16835[23]}}, _zz_16835};
  assign _zz_16837 = fixTo_1742_dout;
  assign _zz_16838 = _zz_16839[31 : 0];
  assign _zz_16839 = _zz_16840;
  assign _zz_16840 = ($signed(_zz_16841) >>> _zz_1454);
  assign _zz_16841 = _zz_16842;
  assign _zz_16842 = ($signed(_zz_16844) - $signed(_zz_1452));
  assign _zz_16843 = ({8'd0,data_mid_66_imag} <<< 8);
  assign _zz_16844 = {{8{_zz_16843[23]}}, _zz_16843};
  assign _zz_16845 = fixTo_1743_dout;
  assign _zz_16846 = _zz_16847[31 : 0];
  assign _zz_16847 = _zz_16848;
  assign _zz_16848 = ($signed(_zz_16849) >>> _zz_1455);
  assign _zz_16849 = _zz_16850;
  assign _zz_16850 = ($signed(_zz_16852) + $signed(_zz_1451));
  assign _zz_16851 = ({8'd0,data_mid_66_real} <<< 8);
  assign _zz_16852 = {{8{_zz_16851[23]}}, _zz_16851};
  assign _zz_16853 = fixTo_1744_dout;
  assign _zz_16854 = _zz_16855[31 : 0];
  assign _zz_16855 = _zz_16856;
  assign _zz_16856 = ($signed(_zz_16857) >>> _zz_1455);
  assign _zz_16857 = _zz_16858;
  assign _zz_16858 = ($signed(_zz_16860) + $signed(_zz_1452));
  assign _zz_16859 = ({8'd0,data_mid_66_imag} <<< 8);
  assign _zz_16860 = {{8{_zz_16859[23]}}, _zz_16859};
  assign _zz_16861 = fixTo_1745_dout;
  assign _zz_16862 = ($signed(twiddle_factor_table_18_real) + $signed(twiddle_factor_table_18_imag));
  assign _zz_16863 = ($signed(_zz_1458) - $signed(_zz_16864));
  assign _zz_16864 = ($signed(_zz_16865) * $signed(twiddle_factor_table_18_imag));
  assign _zz_16865 = ($signed(data_mid_83_real) + $signed(data_mid_83_imag));
  assign _zz_16866 = fixTo_1746_dout;
  assign _zz_16867 = ($signed(_zz_1458) + $signed(_zz_16868));
  assign _zz_16868 = ($signed(_zz_16869) * $signed(twiddle_factor_table_18_real));
  assign _zz_16869 = ($signed(data_mid_83_imag) - $signed(data_mid_83_real));
  assign _zz_16870 = fixTo_1747_dout;
  assign _zz_16871 = _zz_16872[31 : 0];
  assign _zz_16872 = _zz_16873;
  assign _zz_16873 = ($signed(_zz_16874) >>> _zz_1459);
  assign _zz_16874 = _zz_16875;
  assign _zz_16875 = ($signed(_zz_16877) - $signed(_zz_1456));
  assign _zz_16876 = ({8'd0,data_mid_67_real} <<< 8);
  assign _zz_16877 = {{8{_zz_16876[23]}}, _zz_16876};
  assign _zz_16878 = fixTo_1748_dout;
  assign _zz_16879 = _zz_16880[31 : 0];
  assign _zz_16880 = _zz_16881;
  assign _zz_16881 = ($signed(_zz_16882) >>> _zz_1459);
  assign _zz_16882 = _zz_16883;
  assign _zz_16883 = ($signed(_zz_16885) - $signed(_zz_1457));
  assign _zz_16884 = ({8'd0,data_mid_67_imag} <<< 8);
  assign _zz_16885 = {{8{_zz_16884[23]}}, _zz_16884};
  assign _zz_16886 = fixTo_1749_dout;
  assign _zz_16887 = _zz_16888[31 : 0];
  assign _zz_16888 = _zz_16889;
  assign _zz_16889 = ($signed(_zz_16890) >>> _zz_1460);
  assign _zz_16890 = _zz_16891;
  assign _zz_16891 = ($signed(_zz_16893) + $signed(_zz_1456));
  assign _zz_16892 = ({8'd0,data_mid_67_real} <<< 8);
  assign _zz_16893 = {{8{_zz_16892[23]}}, _zz_16892};
  assign _zz_16894 = fixTo_1750_dout;
  assign _zz_16895 = _zz_16896[31 : 0];
  assign _zz_16896 = _zz_16897;
  assign _zz_16897 = ($signed(_zz_16898) >>> _zz_1460);
  assign _zz_16898 = _zz_16899;
  assign _zz_16899 = ($signed(_zz_16901) + $signed(_zz_1457));
  assign _zz_16900 = ({8'd0,data_mid_67_imag} <<< 8);
  assign _zz_16901 = {{8{_zz_16900[23]}}, _zz_16900};
  assign _zz_16902 = fixTo_1751_dout;
  assign _zz_16903 = ($signed(twiddle_factor_table_19_real) + $signed(twiddle_factor_table_19_imag));
  assign _zz_16904 = ($signed(_zz_1463) - $signed(_zz_16905));
  assign _zz_16905 = ($signed(_zz_16906) * $signed(twiddle_factor_table_19_imag));
  assign _zz_16906 = ($signed(data_mid_84_real) + $signed(data_mid_84_imag));
  assign _zz_16907 = fixTo_1752_dout;
  assign _zz_16908 = ($signed(_zz_1463) + $signed(_zz_16909));
  assign _zz_16909 = ($signed(_zz_16910) * $signed(twiddle_factor_table_19_real));
  assign _zz_16910 = ($signed(data_mid_84_imag) - $signed(data_mid_84_real));
  assign _zz_16911 = fixTo_1753_dout;
  assign _zz_16912 = _zz_16913[31 : 0];
  assign _zz_16913 = _zz_16914;
  assign _zz_16914 = ($signed(_zz_16915) >>> _zz_1464);
  assign _zz_16915 = _zz_16916;
  assign _zz_16916 = ($signed(_zz_16918) - $signed(_zz_1461));
  assign _zz_16917 = ({8'd0,data_mid_68_real} <<< 8);
  assign _zz_16918 = {{8{_zz_16917[23]}}, _zz_16917};
  assign _zz_16919 = fixTo_1754_dout;
  assign _zz_16920 = _zz_16921[31 : 0];
  assign _zz_16921 = _zz_16922;
  assign _zz_16922 = ($signed(_zz_16923) >>> _zz_1464);
  assign _zz_16923 = _zz_16924;
  assign _zz_16924 = ($signed(_zz_16926) - $signed(_zz_1462));
  assign _zz_16925 = ({8'd0,data_mid_68_imag} <<< 8);
  assign _zz_16926 = {{8{_zz_16925[23]}}, _zz_16925};
  assign _zz_16927 = fixTo_1755_dout;
  assign _zz_16928 = _zz_16929[31 : 0];
  assign _zz_16929 = _zz_16930;
  assign _zz_16930 = ($signed(_zz_16931) >>> _zz_1465);
  assign _zz_16931 = _zz_16932;
  assign _zz_16932 = ($signed(_zz_16934) + $signed(_zz_1461));
  assign _zz_16933 = ({8'd0,data_mid_68_real} <<< 8);
  assign _zz_16934 = {{8{_zz_16933[23]}}, _zz_16933};
  assign _zz_16935 = fixTo_1756_dout;
  assign _zz_16936 = _zz_16937[31 : 0];
  assign _zz_16937 = _zz_16938;
  assign _zz_16938 = ($signed(_zz_16939) >>> _zz_1465);
  assign _zz_16939 = _zz_16940;
  assign _zz_16940 = ($signed(_zz_16942) + $signed(_zz_1462));
  assign _zz_16941 = ({8'd0,data_mid_68_imag} <<< 8);
  assign _zz_16942 = {{8{_zz_16941[23]}}, _zz_16941};
  assign _zz_16943 = fixTo_1757_dout;
  assign _zz_16944 = ($signed(twiddle_factor_table_20_real) + $signed(twiddle_factor_table_20_imag));
  assign _zz_16945 = ($signed(_zz_1468) - $signed(_zz_16946));
  assign _zz_16946 = ($signed(_zz_16947) * $signed(twiddle_factor_table_20_imag));
  assign _zz_16947 = ($signed(data_mid_85_real) + $signed(data_mid_85_imag));
  assign _zz_16948 = fixTo_1758_dout;
  assign _zz_16949 = ($signed(_zz_1468) + $signed(_zz_16950));
  assign _zz_16950 = ($signed(_zz_16951) * $signed(twiddle_factor_table_20_real));
  assign _zz_16951 = ($signed(data_mid_85_imag) - $signed(data_mid_85_real));
  assign _zz_16952 = fixTo_1759_dout;
  assign _zz_16953 = _zz_16954[31 : 0];
  assign _zz_16954 = _zz_16955;
  assign _zz_16955 = ($signed(_zz_16956) >>> _zz_1469);
  assign _zz_16956 = _zz_16957;
  assign _zz_16957 = ($signed(_zz_16959) - $signed(_zz_1466));
  assign _zz_16958 = ({8'd0,data_mid_69_real} <<< 8);
  assign _zz_16959 = {{8{_zz_16958[23]}}, _zz_16958};
  assign _zz_16960 = fixTo_1760_dout;
  assign _zz_16961 = _zz_16962[31 : 0];
  assign _zz_16962 = _zz_16963;
  assign _zz_16963 = ($signed(_zz_16964) >>> _zz_1469);
  assign _zz_16964 = _zz_16965;
  assign _zz_16965 = ($signed(_zz_16967) - $signed(_zz_1467));
  assign _zz_16966 = ({8'd0,data_mid_69_imag} <<< 8);
  assign _zz_16967 = {{8{_zz_16966[23]}}, _zz_16966};
  assign _zz_16968 = fixTo_1761_dout;
  assign _zz_16969 = _zz_16970[31 : 0];
  assign _zz_16970 = _zz_16971;
  assign _zz_16971 = ($signed(_zz_16972) >>> _zz_1470);
  assign _zz_16972 = _zz_16973;
  assign _zz_16973 = ($signed(_zz_16975) + $signed(_zz_1466));
  assign _zz_16974 = ({8'd0,data_mid_69_real} <<< 8);
  assign _zz_16975 = {{8{_zz_16974[23]}}, _zz_16974};
  assign _zz_16976 = fixTo_1762_dout;
  assign _zz_16977 = _zz_16978[31 : 0];
  assign _zz_16978 = _zz_16979;
  assign _zz_16979 = ($signed(_zz_16980) >>> _zz_1470);
  assign _zz_16980 = _zz_16981;
  assign _zz_16981 = ($signed(_zz_16983) + $signed(_zz_1467));
  assign _zz_16982 = ({8'd0,data_mid_69_imag} <<< 8);
  assign _zz_16983 = {{8{_zz_16982[23]}}, _zz_16982};
  assign _zz_16984 = fixTo_1763_dout;
  assign _zz_16985 = ($signed(twiddle_factor_table_21_real) + $signed(twiddle_factor_table_21_imag));
  assign _zz_16986 = ($signed(_zz_1473) - $signed(_zz_16987));
  assign _zz_16987 = ($signed(_zz_16988) * $signed(twiddle_factor_table_21_imag));
  assign _zz_16988 = ($signed(data_mid_86_real) + $signed(data_mid_86_imag));
  assign _zz_16989 = fixTo_1764_dout;
  assign _zz_16990 = ($signed(_zz_1473) + $signed(_zz_16991));
  assign _zz_16991 = ($signed(_zz_16992) * $signed(twiddle_factor_table_21_real));
  assign _zz_16992 = ($signed(data_mid_86_imag) - $signed(data_mid_86_real));
  assign _zz_16993 = fixTo_1765_dout;
  assign _zz_16994 = _zz_16995[31 : 0];
  assign _zz_16995 = _zz_16996;
  assign _zz_16996 = ($signed(_zz_16997) >>> _zz_1474);
  assign _zz_16997 = _zz_16998;
  assign _zz_16998 = ($signed(_zz_17000) - $signed(_zz_1471));
  assign _zz_16999 = ({8'd0,data_mid_70_real} <<< 8);
  assign _zz_17000 = {{8{_zz_16999[23]}}, _zz_16999};
  assign _zz_17001 = fixTo_1766_dout;
  assign _zz_17002 = _zz_17003[31 : 0];
  assign _zz_17003 = _zz_17004;
  assign _zz_17004 = ($signed(_zz_17005) >>> _zz_1474);
  assign _zz_17005 = _zz_17006;
  assign _zz_17006 = ($signed(_zz_17008) - $signed(_zz_1472));
  assign _zz_17007 = ({8'd0,data_mid_70_imag} <<< 8);
  assign _zz_17008 = {{8{_zz_17007[23]}}, _zz_17007};
  assign _zz_17009 = fixTo_1767_dout;
  assign _zz_17010 = _zz_17011[31 : 0];
  assign _zz_17011 = _zz_17012;
  assign _zz_17012 = ($signed(_zz_17013) >>> _zz_1475);
  assign _zz_17013 = _zz_17014;
  assign _zz_17014 = ($signed(_zz_17016) + $signed(_zz_1471));
  assign _zz_17015 = ({8'd0,data_mid_70_real} <<< 8);
  assign _zz_17016 = {{8{_zz_17015[23]}}, _zz_17015};
  assign _zz_17017 = fixTo_1768_dout;
  assign _zz_17018 = _zz_17019[31 : 0];
  assign _zz_17019 = _zz_17020;
  assign _zz_17020 = ($signed(_zz_17021) >>> _zz_1475);
  assign _zz_17021 = _zz_17022;
  assign _zz_17022 = ($signed(_zz_17024) + $signed(_zz_1472));
  assign _zz_17023 = ({8'd0,data_mid_70_imag} <<< 8);
  assign _zz_17024 = {{8{_zz_17023[23]}}, _zz_17023};
  assign _zz_17025 = fixTo_1769_dout;
  assign _zz_17026 = ($signed(twiddle_factor_table_22_real) + $signed(twiddle_factor_table_22_imag));
  assign _zz_17027 = ($signed(_zz_1478) - $signed(_zz_17028));
  assign _zz_17028 = ($signed(_zz_17029) * $signed(twiddle_factor_table_22_imag));
  assign _zz_17029 = ($signed(data_mid_87_real) + $signed(data_mid_87_imag));
  assign _zz_17030 = fixTo_1770_dout;
  assign _zz_17031 = ($signed(_zz_1478) + $signed(_zz_17032));
  assign _zz_17032 = ($signed(_zz_17033) * $signed(twiddle_factor_table_22_real));
  assign _zz_17033 = ($signed(data_mid_87_imag) - $signed(data_mid_87_real));
  assign _zz_17034 = fixTo_1771_dout;
  assign _zz_17035 = _zz_17036[31 : 0];
  assign _zz_17036 = _zz_17037;
  assign _zz_17037 = ($signed(_zz_17038) >>> _zz_1479);
  assign _zz_17038 = _zz_17039;
  assign _zz_17039 = ($signed(_zz_17041) - $signed(_zz_1476));
  assign _zz_17040 = ({8'd0,data_mid_71_real} <<< 8);
  assign _zz_17041 = {{8{_zz_17040[23]}}, _zz_17040};
  assign _zz_17042 = fixTo_1772_dout;
  assign _zz_17043 = _zz_17044[31 : 0];
  assign _zz_17044 = _zz_17045;
  assign _zz_17045 = ($signed(_zz_17046) >>> _zz_1479);
  assign _zz_17046 = _zz_17047;
  assign _zz_17047 = ($signed(_zz_17049) - $signed(_zz_1477));
  assign _zz_17048 = ({8'd0,data_mid_71_imag} <<< 8);
  assign _zz_17049 = {{8{_zz_17048[23]}}, _zz_17048};
  assign _zz_17050 = fixTo_1773_dout;
  assign _zz_17051 = _zz_17052[31 : 0];
  assign _zz_17052 = _zz_17053;
  assign _zz_17053 = ($signed(_zz_17054) >>> _zz_1480);
  assign _zz_17054 = _zz_17055;
  assign _zz_17055 = ($signed(_zz_17057) + $signed(_zz_1476));
  assign _zz_17056 = ({8'd0,data_mid_71_real} <<< 8);
  assign _zz_17057 = {{8{_zz_17056[23]}}, _zz_17056};
  assign _zz_17058 = fixTo_1774_dout;
  assign _zz_17059 = _zz_17060[31 : 0];
  assign _zz_17060 = _zz_17061;
  assign _zz_17061 = ($signed(_zz_17062) >>> _zz_1480);
  assign _zz_17062 = _zz_17063;
  assign _zz_17063 = ($signed(_zz_17065) + $signed(_zz_1477));
  assign _zz_17064 = ({8'd0,data_mid_71_imag} <<< 8);
  assign _zz_17065 = {{8{_zz_17064[23]}}, _zz_17064};
  assign _zz_17066 = fixTo_1775_dout;
  assign _zz_17067 = ($signed(twiddle_factor_table_23_real) + $signed(twiddle_factor_table_23_imag));
  assign _zz_17068 = ($signed(_zz_1483) - $signed(_zz_17069));
  assign _zz_17069 = ($signed(_zz_17070) * $signed(twiddle_factor_table_23_imag));
  assign _zz_17070 = ($signed(data_mid_88_real) + $signed(data_mid_88_imag));
  assign _zz_17071 = fixTo_1776_dout;
  assign _zz_17072 = ($signed(_zz_1483) + $signed(_zz_17073));
  assign _zz_17073 = ($signed(_zz_17074) * $signed(twiddle_factor_table_23_real));
  assign _zz_17074 = ($signed(data_mid_88_imag) - $signed(data_mid_88_real));
  assign _zz_17075 = fixTo_1777_dout;
  assign _zz_17076 = _zz_17077[31 : 0];
  assign _zz_17077 = _zz_17078;
  assign _zz_17078 = ($signed(_zz_17079) >>> _zz_1484);
  assign _zz_17079 = _zz_17080;
  assign _zz_17080 = ($signed(_zz_17082) - $signed(_zz_1481));
  assign _zz_17081 = ({8'd0,data_mid_72_real} <<< 8);
  assign _zz_17082 = {{8{_zz_17081[23]}}, _zz_17081};
  assign _zz_17083 = fixTo_1778_dout;
  assign _zz_17084 = _zz_17085[31 : 0];
  assign _zz_17085 = _zz_17086;
  assign _zz_17086 = ($signed(_zz_17087) >>> _zz_1484);
  assign _zz_17087 = _zz_17088;
  assign _zz_17088 = ($signed(_zz_17090) - $signed(_zz_1482));
  assign _zz_17089 = ({8'd0,data_mid_72_imag} <<< 8);
  assign _zz_17090 = {{8{_zz_17089[23]}}, _zz_17089};
  assign _zz_17091 = fixTo_1779_dout;
  assign _zz_17092 = _zz_17093[31 : 0];
  assign _zz_17093 = _zz_17094;
  assign _zz_17094 = ($signed(_zz_17095) >>> _zz_1485);
  assign _zz_17095 = _zz_17096;
  assign _zz_17096 = ($signed(_zz_17098) + $signed(_zz_1481));
  assign _zz_17097 = ({8'd0,data_mid_72_real} <<< 8);
  assign _zz_17098 = {{8{_zz_17097[23]}}, _zz_17097};
  assign _zz_17099 = fixTo_1780_dout;
  assign _zz_17100 = _zz_17101[31 : 0];
  assign _zz_17101 = _zz_17102;
  assign _zz_17102 = ($signed(_zz_17103) >>> _zz_1485);
  assign _zz_17103 = _zz_17104;
  assign _zz_17104 = ($signed(_zz_17106) + $signed(_zz_1482));
  assign _zz_17105 = ({8'd0,data_mid_72_imag} <<< 8);
  assign _zz_17106 = {{8{_zz_17105[23]}}, _zz_17105};
  assign _zz_17107 = fixTo_1781_dout;
  assign _zz_17108 = ($signed(twiddle_factor_table_24_real) + $signed(twiddle_factor_table_24_imag));
  assign _zz_17109 = ($signed(_zz_1488) - $signed(_zz_17110));
  assign _zz_17110 = ($signed(_zz_17111) * $signed(twiddle_factor_table_24_imag));
  assign _zz_17111 = ($signed(data_mid_89_real) + $signed(data_mid_89_imag));
  assign _zz_17112 = fixTo_1782_dout;
  assign _zz_17113 = ($signed(_zz_1488) + $signed(_zz_17114));
  assign _zz_17114 = ($signed(_zz_17115) * $signed(twiddle_factor_table_24_real));
  assign _zz_17115 = ($signed(data_mid_89_imag) - $signed(data_mid_89_real));
  assign _zz_17116 = fixTo_1783_dout;
  assign _zz_17117 = _zz_17118[31 : 0];
  assign _zz_17118 = _zz_17119;
  assign _zz_17119 = ($signed(_zz_17120) >>> _zz_1489);
  assign _zz_17120 = _zz_17121;
  assign _zz_17121 = ($signed(_zz_17123) - $signed(_zz_1486));
  assign _zz_17122 = ({8'd0,data_mid_73_real} <<< 8);
  assign _zz_17123 = {{8{_zz_17122[23]}}, _zz_17122};
  assign _zz_17124 = fixTo_1784_dout;
  assign _zz_17125 = _zz_17126[31 : 0];
  assign _zz_17126 = _zz_17127;
  assign _zz_17127 = ($signed(_zz_17128) >>> _zz_1489);
  assign _zz_17128 = _zz_17129;
  assign _zz_17129 = ($signed(_zz_17131) - $signed(_zz_1487));
  assign _zz_17130 = ({8'd0,data_mid_73_imag} <<< 8);
  assign _zz_17131 = {{8{_zz_17130[23]}}, _zz_17130};
  assign _zz_17132 = fixTo_1785_dout;
  assign _zz_17133 = _zz_17134[31 : 0];
  assign _zz_17134 = _zz_17135;
  assign _zz_17135 = ($signed(_zz_17136) >>> _zz_1490);
  assign _zz_17136 = _zz_17137;
  assign _zz_17137 = ($signed(_zz_17139) + $signed(_zz_1486));
  assign _zz_17138 = ({8'd0,data_mid_73_real} <<< 8);
  assign _zz_17139 = {{8{_zz_17138[23]}}, _zz_17138};
  assign _zz_17140 = fixTo_1786_dout;
  assign _zz_17141 = _zz_17142[31 : 0];
  assign _zz_17142 = _zz_17143;
  assign _zz_17143 = ($signed(_zz_17144) >>> _zz_1490);
  assign _zz_17144 = _zz_17145;
  assign _zz_17145 = ($signed(_zz_17147) + $signed(_zz_1487));
  assign _zz_17146 = ({8'd0,data_mid_73_imag} <<< 8);
  assign _zz_17147 = {{8{_zz_17146[23]}}, _zz_17146};
  assign _zz_17148 = fixTo_1787_dout;
  assign _zz_17149 = ($signed(twiddle_factor_table_25_real) + $signed(twiddle_factor_table_25_imag));
  assign _zz_17150 = ($signed(_zz_1493) - $signed(_zz_17151));
  assign _zz_17151 = ($signed(_zz_17152) * $signed(twiddle_factor_table_25_imag));
  assign _zz_17152 = ($signed(data_mid_90_real) + $signed(data_mid_90_imag));
  assign _zz_17153 = fixTo_1788_dout;
  assign _zz_17154 = ($signed(_zz_1493) + $signed(_zz_17155));
  assign _zz_17155 = ($signed(_zz_17156) * $signed(twiddle_factor_table_25_real));
  assign _zz_17156 = ($signed(data_mid_90_imag) - $signed(data_mid_90_real));
  assign _zz_17157 = fixTo_1789_dout;
  assign _zz_17158 = _zz_17159[31 : 0];
  assign _zz_17159 = _zz_17160;
  assign _zz_17160 = ($signed(_zz_17161) >>> _zz_1494);
  assign _zz_17161 = _zz_17162;
  assign _zz_17162 = ($signed(_zz_17164) - $signed(_zz_1491));
  assign _zz_17163 = ({8'd0,data_mid_74_real} <<< 8);
  assign _zz_17164 = {{8{_zz_17163[23]}}, _zz_17163};
  assign _zz_17165 = fixTo_1790_dout;
  assign _zz_17166 = _zz_17167[31 : 0];
  assign _zz_17167 = _zz_17168;
  assign _zz_17168 = ($signed(_zz_17169) >>> _zz_1494);
  assign _zz_17169 = _zz_17170;
  assign _zz_17170 = ($signed(_zz_17172) - $signed(_zz_1492));
  assign _zz_17171 = ({8'd0,data_mid_74_imag} <<< 8);
  assign _zz_17172 = {{8{_zz_17171[23]}}, _zz_17171};
  assign _zz_17173 = fixTo_1791_dout;
  assign _zz_17174 = _zz_17175[31 : 0];
  assign _zz_17175 = _zz_17176;
  assign _zz_17176 = ($signed(_zz_17177) >>> _zz_1495);
  assign _zz_17177 = _zz_17178;
  assign _zz_17178 = ($signed(_zz_17180) + $signed(_zz_1491));
  assign _zz_17179 = ({8'd0,data_mid_74_real} <<< 8);
  assign _zz_17180 = {{8{_zz_17179[23]}}, _zz_17179};
  assign _zz_17181 = fixTo_1792_dout;
  assign _zz_17182 = _zz_17183[31 : 0];
  assign _zz_17183 = _zz_17184;
  assign _zz_17184 = ($signed(_zz_17185) >>> _zz_1495);
  assign _zz_17185 = _zz_17186;
  assign _zz_17186 = ($signed(_zz_17188) + $signed(_zz_1492));
  assign _zz_17187 = ({8'd0,data_mid_74_imag} <<< 8);
  assign _zz_17188 = {{8{_zz_17187[23]}}, _zz_17187};
  assign _zz_17189 = fixTo_1793_dout;
  assign _zz_17190 = ($signed(twiddle_factor_table_26_real) + $signed(twiddle_factor_table_26_imag));
  assign _zz_17191 = ($signed(_zz_1498) - $signed(_zz_17192));
  assign _zz_17192 = ($signed(_zz_17193) * $signed(twiddle_factor_table_26_imag));
  assign _zz_17193 = ($signed(data_mid_91_real) + $signed(data_mid_91_imag));
  assign _zz_17194 = fixTo_1794_dout;
  assign _zz_17195 = ($signed(_zz_1498) + $signed(_zz_17196));
  assign _zz_17196 = ($signed(_zz_17197) * $signed(twiddle_factor_table_26_real));
  assign _zz_17197 = ($signed(data_mid_91_imag) - $signed(data_mid_91_real));
  assign _zz_17198 = fixTo_1795_dout;
  assign _zz_17199 = _zz_17200[31 : 0];
  assign _zz_17200 = _zz_17201;
  assign _zz_17201 = ($signed(_zz_17202) >>> _zz_1499);
  assign _zz_17202 = _zz_17203;
  assign _zz_17203 = ($signed(_zz_17205) - $signed(_zz_1496));
  assign _zz_17204 = ({8'd0,data_mid_75_real} <<< 8);
  assign _zz_17205 = {{8{_zz_17204[23]}}, _zz_17204};
  assign _zz_17206 = fixTo_1796_dout;
  assign _zz_17207 = _zz_17208[31 : 0];
  assign _zz_17208 = _zz_17209;
  assign _zz_17209 = ($signed(_zz_17210) >>> _zz_1499);
  assign _zz_17210 = _zz_17211;
  assign _zz_17211 = ($signed(_zz_17213) - $signed(_zz_1497));
  assign _zz_17212 = ({8'd0,data_mid_75_imag} <<< 8);
  assign _zz_17213 = {{8{_zz_17212[23]}}, _zz_17212};
  assign _zz_17214 = fixTo_1797_dout;
  assign _zz_17215 = _zz_17216[31 : 0];
  assign _zz_17216 = _zz_17217;
  assign _zz_17217 = ($signed(_zz_17218) >>> _zz_1500);
  assign _zz_17218 = _zz_17219;
  assign _zz_17219 = ($signed(_zz_17221) + $signed(_zz_1496));
  assign _zz_17220 = ({8'd0,data_mid_75_real} <<< 8);
  assign _zz_17221 = {{8{_zz_17220[23]}}, _zz_17220};
  assign _zz_17222 = fixTo_1798_dout;
  assign _zz_17223 = _zz_17224[31 : 0];
  assign _zz_17224 = _zz_17225;
  assign _zz_17225 = ($signed(_zz_17226) >>> _zz_1500);
  assign _zz_17226 = _zz_17227;
  assign _zz_17227 = ($signed(_zz_17229) + $signed(_zz_1497));
  assign _zz_17228 = ({8'd0,data_mid_75_imag} <<< 8);
  assign _zz_17229 = {{8{_zz_17228[23]}}, _zz_17228};
  assign _zz_17230 = fixTo_1799_dout;
  assign _zz_17231 = ($signed(twiddle_factor_table_27_real) + $signed(twiddle_factor_table_27_imag));
  assign _zz_17232 = ($signed(_zz_1503) - $signed(_zz_17233));
  assign _zz_17233 = ($signed(_zz_17234) * $signed(twiddle_factor_table_27_imag));
  assign _zz_17234 = ($signed(data_mid_92_real) + $signed(data_mid_92_imag));
  assign _zz_17235 = fixTo_1800_dout;
  assign _zz_17236 = ($signed(_zz_1503) + $signed(_zz_17237));
  assign _zz_17237 = ($signed(_zz_17238) * $signed(twiddle_factor_table_27_real));
  assign _zz_17238 = ($signed(data_mid_92_imag) - $signed(data_mid_92_real));
  assign _zz_17239 = fixTo_1801_dout;
  assign _zz_17240 = _zz_17241[31 : 0];
  assign _zz_17241 = _zz_17242;
  assign _zz_17242 = ($signed(_zz_17243) >>> _zz_1504);
  assign _zz_17243 = _zz_17244;
  assign _zz_17244 = ($signed(_zz_17246) - $signed(_zz_1501));
  assign _zz_17245 = ({8'd0,data_mid_76_real} <<< 8);
  assign _zz_17246 = {{8{_zz_17245[23]}}, _zz_17245};
  assign _zz_17247 = fixTo_1802_dout;
  assign _zz_17248 = _zz_17249[31 : 0];
  assign _zz_17249 = _zz_17250;
  assign _zz_17250 = ($signed(_zz_17251) >>> _zz_1504);
  assign _zz_17251 = _zz_17252;
  assign _zz_17252 = ($signed(_zz_17254) - $signed(_zz_1502));
  assign _zz_17253 = ({8'd0,data_mid_76_imag} <<< 8);
  assign _zz_17254 = {{8{_zz_17253[23]}}, _zz_17253};
  assign _zz_17255 = fixTo_1803_dout;
  assign _zz_17256 = _zz_17257[31 : 0];
  assign _zz_17257 = _zz_17258;
  assign _zz_17258 = ($signed(_zz_17259) >>> _zz_1505);
  assign _zz_17259 = _zz_17260;
  assign _zz_17260 = ($signed(_zz_17262) + $signed(_zz_1501));
  assign _zz_17261 = ({8'd0,data_mid_76_real} <<< 8);
  assign _zz_17262 = {{8{_zz_17261[23]}}, _zz_17261};
  assign _zz_17263 = fixTo_1804_dout;
  assign _zz_17264 = _zz_17265[31 : 0];
  assign _zz_17265 = _zz_17266;
  assign _zz_17266 = ($signed(_zz_17267) >>> _zz_1505);
  assign _zz_17267 = _zz_17268;
  assign _zz_17268 = ($signed(_zz_17270) + $signed(_zz_1502));
  assign _zz_17269 = ({8'd0,data_mid_76_imag} <<< 8);
  assign _zz_17270 = {{8{_zz_17269[23]}}, _zz_17269};
  assign _zz_17271 = fixTo_1805_dout;
  assign _zz_17272 = ($signed(twiddle_factor_table_28_real) + $signed(twiddle_factor_table_28_imag));
  assign _zz_17273 = ($signed(_zz_1508) - $signed(_zz_17274));
  assign _zz_17274 = ($signed(_zz_17275) * $signed(twiddle_factor_table_28_imag));
  assign _zz_17275 = ($signed(data_mid_93_real) + $signed(data_mid_93_imag));
  assign _zz_17276 = fixTo_1806_dout;
  assign _zz_17277 = ($signed(_zz_1508) + $signed(_zz_17278));
  assign _zz_17278 = ($signed(_zz_17279) * $signed(twiddle_factor_table_28_real));
  assign _zz_17279 = ($signed(data_mid_93_imag) - $signed(data_mid_93_real));
  assign _zz_17280 = fixTo_1807_dout;
  assign _zz_17281 = _zz_17282[31 : 0];
  assign _zz_17282 = _zz_17283;
  assign _zz_17283 = ($signed(_zz_17284) >>> _zz_1509);
  assign _zz_17284 = _zz_17285;
  assign _zz_17285 = ($signed(_zz_17287) - $signed(_zz_1506));
  assign _zz_17286 = ({8'd0,data_mid_77_real} <<< 8);
  assign _zz_17287 = {{8{_zz_17286[23]}}, _zz_17286};
  assign _zz_17288 = fixTo_1808_dout;
  assign _zz_17289 = _zz_17290[31 : 0];
  assign _zz_17290 = _zz_17291;
  assign _zz_17291 = ($signed(_zz_17292) >>> _zz_1509);
  assign _zz_17292 = _zz_17293;
  assign _zz_17293 = ($signed(_zz_17295) - $signed(_zz_1507));
  assign _zz_17294 = ({8'd0,data_mid_77_imag} <<< 8);
  assign _zz_17295 = {{8{_zz_17294[23]}}, _zz_17294};
  assign _zz_17296 = fixTo_1809_dout;
  assign _zz_17297 = _zz_17298[31 : 0];
  assign _zz_17298 = _zz_17299;
  assign _zz_17299 = ($signed(_zz_17300) >>> _zz_1510);
  assign _zz_17300 = _zz_17301;
  assign _zz_17301 = ($signed(_zz_17303) + $signed(_zz_1506));
  assign _zz_17302 = ({8'd0,data_mid_77_real} <<< 8);
  assign _zz_17303 = {{8{_zz_17302[23]}}, _zz_17302};
  assign _zz_17304 = fixTo_1810_dout;
  assign _zz_17305 = _zz_17306[31 : 0];
  assign _zz_17306 = _zz_17307;
  assign _zz_17307 = ($signed(_zz_17308) >>> _zz_1510);
  assign _zz_17308 = _zz_17309;
  assign _zz_17309 = ($signed(_zz_17311) + $signed(_zz_1507));
  assign _zz_17310 = ({8'd0,data_mid_77_imag} <<< 8);
  assign _zz_17311 = {{8{_zz_17310[23]}}, _zz_17310};
  assign _zz_17312 = fixTo_1811_dout;
  assign _zz_17313 = ($signed(twiddle_factor_table_29_real) + $signed(twiddle_factor_table_29_imag));
  assign _zz_17314 = ($signed(_zz_1513) - $signed(_zz_17315));
  assign _zz_17315 = ($signed(_zz_17316) * $signed(twiddle_factor_table_29_imag));
  assign _zz_17316 = ($signed(data_mid_94_real) + $signed(data_mid_94_imag));
  assign _zz_17317 = fixTo_1812_dout;
  assign _zz_17318 = ($signed(_zz_1513) + $signed(_zz_17319));
  assign _zz_17319 = ($signed(_zz_17320) * $signed(twiddle_factor_table_29_real));
  assign _zz_17320 = ($signed(data_mid_94_imag) - $signed(data_mid_94_real));
  assign _zz_17321 = fixTo_1813_dout;
  assign _zz_17322 = _zz_17323[31 : 0];
  assign _zz_17323 = _zz_17324;
  assign _zz_17324 = ($signed(_zz_17325) >>> _zz_1514);
  assign _zz_17325 = _zz_17326;
  assign _zz_17326 = ($signed(_zz_17328) - $signed(_zz_1511));
  assign _zz_17327 = ({8'd0,data_mid_78_real} <<< 8);
  assign _zz_17328 = {{8{_zz_17327[23]}}, _zz_17327};
  assign _zz_17329 = fixTo_1814_dout;
  assign _zz_17330 = _zz_17331[31 : 0];
  assign _zz_17331 = _zz_17332;
  assign _zz_17332 = ($signed(_zz_17333) >>> _zz_1514);
  assign _zz_17333 = _zz_17334;
  assign _zz_17334 = ($signed(_zz_17336) - $signed(_zz_1512));
  assign _zz_17335 = ({8'd0,data_mid_78_imag} <<< 8);
  assign _zz_17336 = {{8{_zz_17335[23]}}, _zz_17335};
  assign _zz_17337 = fixTo_1815_dout;
  assign _zz_17338 = _zz_17339[31 : 0];
  assign _zz_17339 = _zz_17340;
  assign _zz_17340 = ($signed(_zz_17341) >>> _zz_1515);
  assign _zz_17341 = _zz_17342;
  assign _zz_17342 = ($signed(_zz_17344) + $signed(_zz_1511));
  assign _zz_17343 = ({8'd0,data_mid_78_real} <<< 8);
  assign _zz_17344 = {{8{_zz_17343[23]}}, _zz_17343};
  assign _zz_17345 = fixTo_1816_dout;
  assign _zz_17346 = _zz_17347[31 : 0];
  assign _zz_17347 = _zz_17348;
  assign _zz_17348 = ($signed(_zz_17349) >>> _zz_1515);
  assign _zz_17349 = _zz_17350;
  assign _zz_17350 = ($signed(_zz_17352) + $signed(_zz_1512));
  assign _zz_17351 = ({8'd0,data_mid_78_imag} <<< 8);
  assign _zz_17352 = {{8{_zz_17351[23]}}, _zz_17351};
  assign _zz_17353 = fixTo_1817_dout;
  assign _zz_17354 = ($signed(twiddle_factor_table_30_real) + $signed(twiddle_factor_table_30_imag));
  assign _zz_17355 = ($signed(_zz_1518) - $signed(_zz_17356));
  assign _zz_17356 = ($signed(_zz_17357) * $signed(twiddle_factor_table_30_imag));
  assign _zz_17357 = ($signed(data_mid_95_real) + $signed(data_mid_95_imag));
  assign _zz_17358 = fixTo_1818_dout;
  assign _zz_17359 = ($signed(_zz_1518) + $signed(_zz_17360));
  assign _zz_17360 = ($signed(_zz_17361) * $signed(twiddle_factor_table_30_real));
  assign _zz_17361 = ($signed(data_mid_95_imag) - $signed(data_mid_95_real));
  assign _zz_17362 = fixTo_1819_dout;
  assign _zz_17363 = _zz_17364[31 : 0];
  assign _zz_17364 = _zz_17365;
  assign _zz_17365 = ($signed(_zz_17366) >>> _zz_1519);
  assign _zz_17366 = _zz_17367;
  assign _zz_17367 = ($signed(_zz_17369) - $signed(_zz_1516));
  assign _zz_17368 = ({8'd0,data_mid_79_real} <<< 8);
  assign _zz_17369 = {{8{_zz_17368[23]}}, _zz_17368};
  assign _zz_17370 = fixTo_1820_dout;
  assign _zz_17371 = _zz_17372[31 : 0];
  assign _zz_17372 = _zz_17373;
  assign _zz_17373 = ($signed(_zz_17374) >>> _zz_1519);
  assign _zz_17374 = _zz_17375;
  assign _zz_17375 = ($signed(_zz_17377) - $signed(_zz_1517));
  assign _zz_17376 = ({8'd0,data_mid_79_imag} <<< 8);
  assign _zz_17377 = {{8{_zz_17376[23]}}, _zz_17376};
  assign _zz_17378 = fixTo_1821_dout;
  assign _zz_17379 = _zz_17380[31 : 0];
  assign _zz_17380 = _zz_17381;
  assign _zz_17381 = ($signed(_zz_17382) >>> _zz_1520);
  assign _zz_17382 = _zz_17383;
  assign _zz_17383 = ($signed(_zz_17385) + $signed(_zz_1516));
  assign _zz_17384 = ({8'd0,data_mid_79_real} <<< 8);
  assign _zz_17385 = {{8{_zz_17384[23]}}, _zz_17384};
  assign _zz_17386 = fixTo_1822_dout;
  assign _zz_17387 = _zz_17388[31 : 0];
  assign _zz_17388 = _zz_17389;
  assign _zz_17389 = ($signed(_zz_17390) >>> _zz_1520);
  assign _zz_17390 = _zz_17391;
  assign _zz_17391 = ($signed(_zz_17393) + $signed(_zz_1517));
  assign _zz_17392 = ({8'd0,data_mid_79_imag} <<< 8);
  assign _zz_17393 = {{8{_zz_17392[23]}}, _zz_17392};
  assign _zz_17394 = fixTo_1823_dout;
  assign _zz_17395 = ($signed(twiddle_factor_table_15_real) + $signed(twiddle_factor_table_15_imag));
  assign _zz_17396 = ($signed(_zz_1523) - $signed(_zz_17397));
  assign _zz_17397 = ($signed(_zz_17398) * $signed(twiddle_factor_table_15_imag));
  assign _zz_17398 = ($signed(data_mid_112_real) + $signed(data_mid_112_imag));
  assign _zz_17399 = fixTo_1824_dout;
  assign _zz_17400 = ($signed(_zz_1523) + $signed(_zz_17401));
  assign _zz_17401 = ($signed(_zz_17402) * $signed(twiddle_factor_table_15_real));
  assign _zz_17402 = ($signed(data_mid_112_imag) - $signed(data_mid_112_real));
  assign _zz_17403 = fixTo_1825_dout;
  assign _zz_17404 = _zz_17405[31 : 0];
  assign _zz_17405 = _zz_17406;
  assign _zz_17406 = ($signed(_zz_17407) >>> _zz_1524);
  assign _zz_17407 = _zz_17408;
  assign _zz_17408 = ($signed(_zz_17410) - $signed(_zz_1521));
  assign _zz_17409 = ({8'd0,data_mid_96_real} <<< 8);
  assign _zz_17410 = {{8{_zz_17409[23]}}, _zz_17409};
  assign _zz_17411 = fixTo_1826_dout;
  assign _zz_17412 = _zz_17413[31 : 0];
  assign _zz_17413 = _zz_17414;
  assign _zz_17414 = ($signed(_zz_17415) >>> _zz_1524);
  assign _zz_17415 = _zz_17416;
  assign _zz_17416 = ($signed(_zz_17418) - $signed(_zz_1522));
  assign _zz_17417 = ({8'd0,data_mid_96_imag} <<< 8);
  assign _zz_17418 = {{8{_zz_17417[23]}}, _zz_17417};
  assign _zz_17419 = fixTo_1827_dout;
  assign _zz_17420 = _zz_17421[31 : 0];
  assign _zz_17421 = _zz_17422;
  assign _zz_17422 = ($signed(_zz_17423) >>> _zz_1525);
  assign _zz_17423 = _zz_17424;
  assign _zz_17424 = ($signed(_zz_17426) + $signed(_zz_1521));
  assign _zz_17425 = ({8'd0,data_mid_96_real} <<< 8);
  assign _zz_17426 = {{8{_zz_17425[23]}}, _zz_17425};
  assign _zz_17427 = fixTo_1828_dout;
  assign _zz_17428 = _zz_17429[31 : 0];
  assign _zz_17429 = _zz_17430;
  assign _zz_17430 = ($signed(_zz_17431) >>> _zz_1525);
  assign _zz_17431 = _zz_17432;
  assign _zz_17432 = ($signed(_zz_17434) + $signed(_zz_1522));
  assign _zz_17433 = ({8'd0,data_mid_96_imag} <<< 8);
  assign _zz_17434 = {{8{_zz_17433[23]}}, _zz_17433};
  assign _zz_17435 = fixTo_1829_dout;
  assign _zz_17436 = ($signed(twiddle_factor_table_16_real) + $signed(twiddle_factor_table_16_imag));
  assign _zz_17437 = ($signed(_zz_1528) - $signed(_zz_17438));
  assign _zz_17438 = ($signed(_zz_17439) * $signed(twiddle_factor_table_16_imag));
  assign _zz_17439 = ($signed(data_mid_113_real) + $signed(data_mid_113_imag));
  assign _zz_17440 = fixTo_1830_dout;
  assign _zz_17441 = ($signed(_zz_1528) + $signed(_zz_17442));
  assign _zz_17442 = ($signed(_zz_17443) * $signed(twiddle_factor_table_16_real));
  assign _zz_17443 = ($signed(data_mid_113_imag) - $signed(data_mid_113_real));
  assign _zz_17444 = fixTo_1831_dout;
  assign _zz_17445 = _zz_17446[31 : 0];
  assign _zz_17446 = _zz_17447;
  assign _zz_17447 = ($signed(_zz_17448) >>> _zz_1529);
  assign _zz_17448 = _zz_17449;
  assign _zz_17449 = ($signed(_zz_17451) - $signed(_zz_1526));
  assign _zz_17450 = ({8'd0,data_mid_97_real} <<< 8);
  assign _zz_17451 = {{8{_zz_17450[23]}}, _zz_17450};
  assign _zz_17452 = fixTo_1832_dout;
  assign _zz_17453 = _zz_17454[31 : 0];
  assign _zz_17454 = _zz_17455;
  assign _zz_17455 = ($signed(_zz_17456) >>> _zz_1529);
  assign _zz_17456 = _zz_17457;
  assign _zz_17457 = ($signed(_zz_17459) - $signed(_zz_1527));
  assign _zz_17458 = ({8'd0,data_mid_97_imag} <<< 8);
  assign _zz_17459 = {{8{_zz_17458[23]}}, _zz_17458};
  assign _zz_17460 = fixTo_1833_dout;
  assign _zz_17461 = _zz_17462[31 : 0];
  assign _zz_17462 = _zz_17463;
  assign _zz_17463 = ($signed(_zz_17464) >>> _zz_1530);
  assign _zz_17464 = _zz_17465;
  assign _zz_17465 = ($signed(_zz_17467) + $signed(_zz_1526));
  assign _zz_17466 = ({8'd0,data_mid_97_real} <<< 8);
  assign _zz_17467 = {{8{_zz_17466[23]}}, _zz_17466};
  assign _zz_17468 = fixTo_1834_dout;
  assign _zz_17469 = _zz_17470[31 : 0];
  assign _zz_17470 = _zz_17471;
  assign _zz_17471 = ($signed(_zz_17472) >>> _zz_1530);
  assign _zz_17472 = _zz_17473;
  assign _zz_17473 = ($signed(_zz_17475) + $signed(_zz_1527));
  assign _zz_17474 = ({8'd0,data_mid_97_imag} <<< 8);
  assign _zz_17475 = {{8{_zz_17474[23]}}, _zz_17474};
  assign _zz_17476 = fixTo_1835_dout;
  assign _zz_17477 = ($signed(twiddle_factor_table_17_real) + $signed(twiddle_factor_table_17_imag));
  assign _zz_17478 = ($signed(_zz_1533) - $signed(_zz_17479));
  assign _zz_17479 = ($signed(_zz_17480) * $signed(twiddle_factor_table_17_imag));
  assign _zz_17480 = ($signed(data_mid_114_real) + $signed(data_mid_114_imag));
  assign _zz_17481 = fixTo_1836_dout;
  assign _zz_17482 = ($signed(_zz_1533) + $signed(_zz_17483));
  assign _zz_17483 = ($signed(_zz_17484) * $signed(twiddle_factor_table_17_real));
  assign _zz_17484 = ($signed(data_mid_114_imag) - $signed(data_mid_114_real));
  assign _zz_17485 = fixTo_1837_dout;
  assign _zz_17486 = _zz_17487[31 : 0];
  assign _zz_17487 = _zz_17488;
  assign _zz_17488 = ($signed(_zz_17489) >>> _zz_1534);
  assign _zz_17489 = _zz_17490;
  assign _zz_17490 = ($signed(_zz_17492) - $signed(_zz_1531));
  assign _zz_17491 = ({8'd0,data_mid_98_real} <<< 8);
  assign _zz_17492 = {{8{_zz_17491[23]}}, _zz_17491};
  assign _zz_17493 = fixTo_1838_dout;
  assign _zz_17494 = _zz_17495[31 : 0];
  assign _zz_17495 = _zz_17496;
  assign _zz_17496 = ($signed(_zz_17497) >>> _zz_1534);
  assign _zz_17497 = _zz_17498;
  assign _zz_17498 = ($signed(_zz_17500) - $signed(_zz_1532));
  assign _zz_17499 = ({8'd0,data_mid_98_imag} <<< 8);
  assign _zz_17500 = {{8{_zz_17499[23]}}, _zz_17499};
  assign _zz_17501 = fixTo_1839_dout;
  assign _zz_17502 = _zz_17503[31 : 0];
  assign _zz_17503 = _zz_17504;
  assign _zz_17504 = ($signed(_zz_17505) >>> _zz_1535);
  assign _zz_17505 = _zz_17506;
  assign _zz_17506 = ($signed(_zz_17508) + $signed(_zz_1531));
  assign _zz_17507 = ({8'd0,data_mid_98_real} <<< 8);
  assign _zz_17508 = {{8{_zz_17507[23]}}, _zz_17507};
  assign _zz_17509 = fixTo_1840_dout;
  assign _zz_17510 = _zz_17511[31 : 0];
  assign _zz_17511 = _zz_17512;
  assign _zz_17512 = ($signed(_zz_17513) >>> _zz_1535);
  assign _zz_17513 = _zz_17514;
  assign _zz_17514 = ($signed(_zz_17516) + $signed(_zz_1532));
  assign _zz_17515 = ({8'd0,data_mid_98_imag} <<< 8);
  assign _zz_17516 = {{8{_zz_17515[23]}}, _zz_17515};
  assign _zz_17517 = fixTo_1841_dout;
  assign _zz_17518 = ($signed(twiddle_factor_table_18_real) + $signed(twiddle_factor_table_18_imag));
  assign _zz_17519 = ($signed(_zz_1538) - $signed(_zz_17520));
  assign _zz_17520 = ($signed(_zz_17521) * $signed(twiddle_factor_table_18_imag));
  assign _zz_17521 = ($signed(data_mid_115_real) + $signed(data_mid_115_imag));
  assign _zz_17522 = fixTo_1842_dout;
  assign _zz_17523 = ($signed(_zz_1538) + $signed(_zz_17524));
  assign _zz_17524 = ($signed(_zz_17525) * $signed(twiddle_factor_table_18_real));
  assign _zz_17525 = ($signed(data_mid_115_imag) - $signed(data_mid_115_real));
  assign _zz_17526 = fixTo_1843_dout;
  assign _zz_17527 = _zz_17528[31 : 0];
  assign _zz_17528 = _zz_17529;
  assign _zz_17529 = ($signed(_zz_17530) >>> _zz_1539);
  assign _zz_17530 = _zz_17531;
  assign _zz_17531 = ($signed(_zz_17533) - $signed(_zz_1536));
  assign _zz_17532 = ({8'd0,data_mid_99_real} <<< 8);
  assign _zz_17533 = {{8{_zz_17532[23]}}, _zz_17532};
  assign _zz_17534 = fixTo_1844_dout;
  assign _zz_17535 = _zz_17536[31 : 0];
  assign _zz_17536 = _zz_17537;
  assign _zz_17537 = ($signed(_zz_17538) >>> _zz_1539);
  assign _zz_17538 = _zz_17539;
  assign _zz_17539 = ($signed(_zz_17541) - $signed(_zz_1537));
  assign _zz_17540 = ({8'd0,data_mid_99_imag} <<< 8);
  assign _zz_17541 = {{8{_zz_17540[23]}}, _zz_17540};
  assign _zz_17542 = fixTo_1845_dout;
  assign _zz_17543 = _zz_17544[31 : 0];
  assign _zz_17544 = _zz_17545;
  assign _zz_17545 = ($signed(_zz_17546) >>> _zz_1540);
  assign _zz_17546 = _zz_17547;
  assign _zz_17547 = ($signed(_zz_17549) + $signed(_zz_1536));
  assign _zz_17548 = ({8'd0,data_mid_99_real} <<< 8);
  assign _zz_17549 = {{8{_zz_17548[23]}}, _zz_17548};
  assign _zz_17550 = fixTo_1846_dout;
  assign _zz_17551 = _zz_17552[31 : 0];
  assign _zz_17552 = _zz_17553;
  assign _zz_17553 = ($signed(_zz_17554) >>> _zz_1540);
  assign _zz_17554 = _zz_17555;
  assign _zz_17555 = ($signed(_zz_17557) + $signed(_zz_1537));
  assign _zz_17556 = ({8'd0,data_mid_99_imag} <<< 8);
  assign _zz_17557 = {{8{_zz_17556[23]}}, _zz_17556};
  assign _zz_17558 = fixTo_1847_dout;
  assign _zz_17559 = ($signed(twiddle_factor_table_19_real) + $signed(twiddle_factor_table_19_imag));
  assign _zz_17560 = ($signed(_zz_1543) - $signed(_zz_17561));
  assign _zz_17561 = ($signed(_zz_17562) * $signed(twiddle_factor_table_19_imag));
  assign _zz_17562 = ($signed(data_mid_116_real) + $signed(data_mid_116_imag));
  assign _zz_17563 = fixTo_1848_dout;
  assign _zz_17564 = ($signed(_zz_1543) + $signed(_zz_17565));
  assign _zz_17565 = ($signed(_zz_17566) * $signed(twiddle_factor_table_19_real));
  assign _zz_17566 = ($signed(data_mid_116_imag) - $signed(data_mid_116_real));
  assign _zz_17567 = fixTo_1849_dout;
  assign _zz_17568 = _zz_17569[31 : 0];
  assign _zz_17569 = _zz_17570;
  assign _zz_17570 = ($signed(_zz_17571) >>> _zz_1544);
  assign _zz_17571 = _zz_17572;
  assign _zz_17572 = ($signed(_zz_17574) - $signed(_zz_1541));
  assign _zz_17573 = ({8'd0,data_mid_100_real} <<< 8);
  assign _zz_17574 = {{8{_zz_17573[23]}}, _zz_17573};
  assign _zz_17575 = fixTo_1850_dout;
  assign _zz_17576 = _zz_17577[31 : 0];
  assign _zz_17577 = _zz_17578;
  assign _zz_17578 = ($signed(_zz_17579) >>> _zz_1544);
  assign _zz_17579 = _zz_17580;
  assign _zz_17580 = ($signed(_zz_17582) - $signed(_zz_1542));
  assign _zz_17581 = ({8'd0,data_mid_100_imag} <<< 8);
  assign _zz_17582 = {{8{_zz_17581[23]}}, _zz_17581};
  assign _zz_17583 = fixTo_1851_dout;
  assign _zz_17584 = _zz_17585[31 : 0];
  assign _zz_17585 = _zz_17586;
  assign _zz_17586 = ($signed(_zz_17587) >>> _zz_1545);
  assign _zz_17587 = _zz_17588;
  assign _zz_17588 = ($signed(_zz_17590) + $signed(_zz_1541));
  assign _zz_17589 = ({8'd0,data_mid_100_real} <<< 8);
  assign _zz_17590 = {{8{_zz_17589[23]}}, _zz_17589};
  assign _zz_17591 = fixTo_1852_dout;
  assign _zz_17592 = _zz_17593[31 : 0];
  assign _zz_17593 = _zz_17594;
  assign _zz_17594 = ($signed(_zz_17595) >>> _zz_1545);
  assign _zz_17595 = _zz_17596;
  assign _zz_17596 = ($signed(_zz_17598) + $signed(_zz_1542));
  assign _zz_17597 = ({8'd0,data_mid_100_imag} <<< 8);
  assign _zz_17598 = {{8{_zz_17597[23]}}, _zz_17597};
  assign _zz_17599 = fixTo_1853_dout;
  assign _zz_17600 = ($signed(twiddle_factor_table_20_real) + $signed(twiddle_factor_table_20_imag));
  assign _zz_17601 = ($signed(_zz_1548) - $signed(_zz_17602));
  assign _zz_17602 = ($signed(_zz_17603) * $signed(twiddle_factor_table_20_imag));
  assign _zz_17603 = ($signed(data_mid_117_real) + $signed(data_mid_117_imag));
  assign _zz_17604 = fixTo_1854_dout;
  assign _zz_17605 = ($signed(_zz_1548) + $signed(_zz_17606));
  assign _zz_17606 = ($signed(_zz_17607) * $signed(twiddle_factor_table_20_real));
  assign _zz_17607 = ($signed(data_mid_117_imag) - $signed(data_mid_117_real));
  assign _zz_17608 = fixTo_1855_dout;
  assign _zz_17609 = _zz_17610[31 : 0];
  assign _zz_17610 = _zz_17611;
  assign _zz_17611 = ($signed(_zz_17612) >>> _zz_1549);
  assign _zz_17612 = _zz_17613;
  assign _zz_17613 = ($signed(_zz_17615) - $signed(_zz_1546));
  assign _zz_17614 = ({8'd0,data_mid_101_real} <<< 8);
  assign _zz_17615 = {{8{_zz_17614[23]}}, _zz_17614};
  assign _zz_17616 = fixTo_1856_dout;
  assign _zz_17617 = _zz_17618[31 : 0];
  assign _zz_17618 = _zz_17619;
  assign _zz_17619 = ($signed(_zz_17620) >>> _zz_1549);
  assign _zz_17620 = _zz_17621;
  assign _zz_17621 = ($signed(_zz_17623) - $signed(_zz_1547));
  assign _zz_17622 = ({8'd0,data_mid_101_imag} <<< 8);
  assign _zz_17623 = {{8{_zz_17622[23]}}, _zz_17622};
  assign _zz_17624 = fixTo_1857_dout;
  assign _zz_17625 = _zz_17626[31 : 0];
  assign _zz_17626 = _zz_17627;
  assign _zz_17627 = ($signed(_zz_17628) >>> _zz_1550);
  assign _zz_17628 = _zz_17629;
  assign _zz_17629 = ($signed(_zz_17631) + $signed(_zz_1546));
  assign _zz_17630 = ({8'd0,data_mid_101_real} <<< 8);
  assign _zz_17631 = {{8{_zz_17630[23]}}, _zz_17630};
  assign _zz_17632 = fixTo_1858_dout;
  assign _zz_17633 = _zz_17634[31 : 0];
  assign _zz_17634 = _zz_17635;
  assign _zz_17635 = ($signed(_zz_17636) >>> _zz_1550);
  assign _zz_17636 = _zz_17637;
  assign _zz_17637 = ($signed(_zz_17639) + $signed(_zz_1547));
  assign _zz_17638 = ({8'd0,data_mid_101_imag} <<< 8);
  assign _zz_17639 = {{8{_zz_17638[23]}}, _zz_17638};
  assign _zz_17640 = fixTo_1859_dout;
  assign _zz_17641 = ($signed(twiddle_factor_table_21_real) + $signed(twiddle_factor_table_21_imag));
  assign _zz_17642 = ($signed(_zz_1553) - $signed(_zz_17643));
  assign _zz_17643 = ($signed(_zz_17644) * $signed(twiddle_factor_table_21_imag));
  assign _zz_17644 = ($signed(data_mid_118_real) + $signed(data_mid_118_imag));
  assign _zz_17645 = fixTo_1860_dout;
  assign _zz_17646 = ($signed(_zz_1553) + $signed(_zz_17647));
  assign _zz_17647 = ($signed(_zz_17648) * $signed(twiddle_factor_table_21_real));
  assign _zz_17648 = ($signed(data_mid_118_imag) - $signed(data_mid_118_real));
  assign _zz_17649 = fixTo_1861_dout;
  assign _zz_17650 = _zz_17651[31 : 0];
  assign _zz_17651 = _zz_17652;
  assign _zz_17652 = ($signed(_zz_17653) >>> _zz_1554);
  assign _zz_17653 = _zz_17654;
  assign _zz_17654 = ($signed(_zz_17656) - $signed(_zz_1551));
  assign _zz_17655 = ({8'd0,data_mid_102_real} <<< 8);
  assign _zz_17656 = {{8{_zz_17655[23]}}, _zz_17655};
  assign _zz_17657 = fixTo_1862_dout;
  assign _zz_17658 = _zz_17659[31 : 0];
  assign _zz_17659 = _zz_17660;
  assign _zz_17660 = ($signed(_zz_17661) >>> _zz_1554);
  assign _zz_17661 = _zz_17662;
  assign _zz_17662 = ($signed(_zz_17664) - $signed(_zz_1552));
  assign _zz_17663 = ({8'd0,data_mid_102_imag} <<< 8);
  assign _zz_17664 = {{8{_zz_17663[23]}}, _zz_17663};
  assign _zz_17665 = fixTo_1863_dout;
  assign _zz_17666 = _zz_17667[31 : 0];
  assign _zz_17667 = _zz_17668;
  assign _zz_17668 = ($signed(_zz_17669) >>> _zz_1555);
  assign _zz_17669 = _zz_17670;
  assign _zz_17670 = ($signed(_zz_17672) + $signed(_zz_1551));
  assign _zz_17671 = ({8'd0,data_mid_102_real} <<< 8);
  assign _zz_17672 = {{8{_zz_17671[23]}}, _zz_17671};
  assign _zz_17673 = fixTo_1864_dout;
  assign _zz_17674 = _zz_17675[31 : 0];
  assign _zz_17675 = _zz_17676;
  assign _zz_17676 = ($signed(_zz_17677) >>> _zz_1555);
  assign _zz_17677 = _zz_17678;
  assign _zz_17678 = ($signed(_zz_17680) + $signed(_zz_1552));
  assign _zz_17679 = ({8'd0,data_mid_102_imag} <<< 8);
  assign _zz_17680 = {{8{_zz_17679[23]}}, _zz_17679};
  assign _zz_17681 = fixTo_1865_dout;
  assign _zz_17682 = ($signed(twiddle_factor_table_22_real) + $signed(twiddle_factor_table_22_imag));
  assign _zz_17683 = ($signed(_zz_1558) - $signed(_zz_17684));
  assign _zz_17684 = ($signed(_zz_17685) * $signed(twiddle_factor_table_22_imag));
  assign _zz_17685 = ($signed(data_mid_119_real) + $signed(data_mid_119_imag));
  assign _zz_17686 = fixTo_1866_dout;
  assign _zz_17687 = ($signed(_zz_1558) + $signed(_zz_17688));
  assign _zz_17688 = ($signed(_zz_17689) * $signed(twiddle_factor_table_22_real));
  assign _zz_17689 = ($signed(data_mid_119_imag) - $signed(data_mid_119_real));
  assign _zz_17690 = fixTo_1867_dout;
  assign _zz_17691 = _zz_17692[31 : 0];
  assign _zz_17692 = _zz_17693;
  assign _zz_17693 = ($signed(_zz_17694) >>> _zz_1559);
  assign _zz_17694 = _zz_17695;
  assign _zz_17695 = ($signed(_zz_17697) - $signed(_zz_1556));
  assign _zz_17696 = ({8'd0,data_mid_103_real} <<< 8);
  assign _zz_17697 = {{8{_zz_17696[23]}}, _zz_17696};
  assign _zz_17698 = fixTo_1868_dout;
  assign _zz_17699 = _zz_17700[31 : 0];
  assign _zz_17700 = _zz_17701;
  assign _zz_17701 = ($signed(_zz_17702) >>> _zz_1559);
  assign _zz_17702 = _zz_17703;
  assign _zz_17703 = ($signed(_zz_17705) - $signed(_zz_1557));
  assign _zz_17704 = ({8'd0,data_mid_103_imag} <<< 8);
  assign _zz_17705 = {{8{_zz_17704[23]}}, _zz_17704};
  assign _zz_17706 = fixTo_1869_dout;
  assign _zz_17707 = _zz_17708[31 : 0];
  assign _zz_17708 = _zz_17709;
  assign _zz_17709 = ($signed(_zz_17710) >>> _zz_1560);
  assign _zz_17710 = _zz_17711;
  assign _zz_17711 = ($signed(_zz_17713) + $signed(_zz_1556));
  assign _zz_17712 = ({8'd0,data_mid_103_real} <<< 8);
  assign _zz_17713 = {{8{_zz_17712[23]}}, _zz_17712};
  assign _zz_17714 = fixTo_1870_dout;
  assign _zz_17715 = _zz_17716[31 : 0];
  assign _zz_17716 = _zz_17717;
  assign _zz_17717 = ($signed(_zz_17718) >>> _zz_1560);
  assign _zz_17718 = _zz_17719;
  assign _zz_17719 = ($signed(_zz_17721) + $signed(_zz_1557));
  assign _zz_17720 = ({8'd0,data_mid_103_imag} <<< 8);
  assign _zz_17721 = {{8{_zz_17720[23]}}, _zz_17720};
  assign _zz_17722 = fixTo_1871_dout;
  assign _zz_17723 = ($signed(twiddle_factor_table_23_real) + $signed(twiddle_factor_table_23_imag));
  assign _zz_17724 = ($signed(_zz_1563) - $signed(_zz_17725));
  assign _zz_17725 = ($signed(_zz_17726) * $signed(twiddle_factor_table_23_imag));
  assign _zz_17726 = ($signed(data_mid_120_real) + $signed(data_mid_120_imag));
  assign _zz_17727 = fixTo_1872_dout;
  assign _zz_17728 = ($signed(_zz_1563) + $signed(_zz_17729));
  assign _zz_17729 = ($signed(_zz_17730) * $signed(twiddle_factor_table_23_real));
  assign _zz_17730 = ($signed(data_mid_120_imag) - $signed(data_mid_120_real));
  assign _zz_17731 = fixTo_1873_dout;
  assign _zz_17732 = _zz_17733[31 : 0];
  assign _zz_17733 = _zz_17734;
  assign _zz_17734 = ($signed(_zz_17735) >>> _zz_1564);
  assign _zz_17735 = _zz_17736;
  assign _zz_17736 = ($signed(_zz_17738) - $signed(_zz_1561));
  assign _zz_17737 = ({8'd0,data_mid_104_real} <<< 8);
  assign _zz_17738 = {{8{_zz_17737[23]}}, _zz_17737};
  assign _zz_17739 = fixTo_1874_dout;
  assign _zz_17740 = _zz_17741[31 : 0];
  assign _zz_17741 = _zz_17742;
  assign _zz_17742 = ($signed(_zz_17743) >>> _zz_1564);
  assign _zz_17743 = _zz_17744;
  assign _zz_17744 = ($signed(_zz_17746) - $signed(_zz_1562));
  assign _zz_17745 = ({8'd0,data_mid_104_imag} <<< 8);
  assign _zz_17746 = {{8{_zz_17745[23]}}, _zz_17745};
  assign _zz_17747 = fixTo_1875_dout;
  assign _zz_17748 = _zz_17749[31 : 0];
  assign _zz_17749 = _zz_17750;
  assign _zz_17750 = ($signed(_zz_17751) >>> _zz_1565);
  assign _zz_17751 = _zz_17752;
  assign _zz_17752 = ($signed(_zz_17754) + $signed(_zz_1561));
  assign _zz_17753 = ({8'd0,data_mid_104_real} <<< 8);
  assign _zz_17754 = {{8{_zz_17753[23]}}, _zz_17753};
  assign _zz_17755 = fixTo_1876_dout;
  assign _zz_17756 = _zz_17757[31 : 0];
  assign _zz_17757 = _zz_17758;
  assign _zz_17758 = ($signed(_zz_17759) >>> _zz_1565);
  assign _zz_17759 = _zz_17760;
  assign _zz_17760 = ($signed(_zz_17762) + $signed(_zz_1562));
  assign _zz_17761 = ({8'd0,data_mid_104_imag} <<< 8);
  assign _zz_17762 = {{8{_zz_17761[23]}}, _zz_17761};
  assign _zz_17763 = fixTo_1877_dout;
  assign _zz_17764 = ($signed(twiddle_factor_table_24_real) + $signed(twiddle_factor_table_24_imag));
  assign _zz_17765 = ($signed(_zz_1568) - $signed(_zz_17766));
  assign _zz_17766 = ($signed(_zz_17767) * $signed(twiddle_factor_table_24_imag));
  assign _zz_17767 = ($signed(data_mid_121_real) + $signed(data_mid_121_imag));
  assign _zz_17768 = fixTo_1878_dout;
  assign _zz_17769 = ($signed(_zz_1568) + $signed(_zz_17770));
  assign _zz_17770 = ($signed(_zz_17771) * $signed(twiddle_factor_table_24_real));
  assign _zz_17771 = ($signed(data_mid_121_imag) - $signed(data_mid_121_real));
  assign _zz_17772 = fixTo_1879_dout;
  assign _zz_17773 = _zz_17774[31 : 0];
  assign _zz_17774 = _zz_17775;
  assign _zz_17775 = ($signed(_zz_17776) >>> _zz_1569);
  assign _zz_17776 = _zz_17777;
  assign _zz_17777 = ($signed(_zz_17779) - $signed(_zz_1566));
  assign _zz_17778 = ({8'd0,data_mid_105_real} <<< 8);
  assign _zz_17779 = {{8{_zz_17778[23]}}, _zz_17778};
  assign _zz_17780 = fixTo_1880_dout;
  assign _zz_17781 = _zz_17782[31 : 0];
  assign _zz_17782 = _zz_17783;
  assign _zz_17783 = ($signed(_zz_17784) >>> _zz_1569);
  assign _zz_17784 = _zz_17785;
  assign _zz_17785 = ($signed(_zz_17787) - $signed(_zz_1567));
  assign _zz_17786 = ({8'd0,data_mid_105_imag} <<< 8);
  assign _zz_17787 = {{8{_zz_17786[23]}}, _zz_17786};
  assign _zz_17788 = fixTo_1881_dout;
  assign _zz_17789 = _zz_17790[31 : 0];
  assign _zz_17790 = _zz_17791;
  assign _zz_17791 = ($signed(_zz_17792) >>> _zz_1570);
  assign _zz_17792 = _zz_17793;
  assign _zz_17793 = ($signed(_zz_17795) + $signed(_zz_1566));
  assign _zz_17794 = ({8'd0,data_mid_105_real} <<< 8);
  assign _zz_17795 = {{8{_zz_17794[23]}}, _zz_17794};
  assign _zz_17796 = fixTo_1882_dout;
  assign _zz_17797 = _zz_17798[31 : 0];
  assign _zz_17798 = _zz_17799;
  assign _zz_17799 = ($signed(_zz_17800) >>> _zz_1570);
  assign _zz_17800 = _zz_17801;
  assign _zz_17801 = ($signed(_zz_17803) + $signed(_zz_1567));
  assign _zz_17802 = ({8'd0,data_mid_105_imag} <<< 8);
  assign _zz_17803 = {{8{_zz_17802[23]}}, _zz_17802};
  assign _zz_17804 = fixTo_1883_dout;
  assign _zz_17805 = ($signed(twiddle_factor_table_25_real) + $signed(twiddle_factor_table_25_imag));
  assign _zz_17806 = ($signed(_zz_1573) - $signed(_zz_17807));
  assign _zz_17807 = ($signed(_zz_17808) * $signed(twiddle_factor_table_25_imag));
  assign _zz_17808 = ($signed(data_mid_122_real) + $signed(data_mid_122_imag));
  assign _zz_17809 = fixTo_1884_dout;
  assign _zz_17810 = ($signed(_zz_1573) + $signed(_zz_17811));
  assign _zz_17811 = ($signed(_zz_17812) * $signed(twiddle_factor_table_25_real));
  assign _zz_17812 = ($signed(data_mid_122_imag) - $signed(data_mid_122_real));
  assign _zz_17813 = fixTo_1885_dout;
  assign _zz_17814 = _zz_17815[31 : 0];
  assign _zz_17815 = _zz_17816;
  assign _zz_17816 = ($signed(_zz_17817) >>> _zz_1574);
  assign _zz_17817 = _zz_17818;
  assign _zz_17818 = ($signed(_zz_17820) - $signed(_zz_1571));
  assign _zz_17819 = ({8'd0,data_mid_106_real} <<< 8);
  assign _zz_17820 = {{8{_zz_17819[23]}}, _zz_17819};
  assign _zz_17821 = fixTo_1886_dout;
  assign _zz_17822 = _zz_17823[31 : 0];
  assign _zz_17823 = _zz_17824;
  assign _zz_17824 = ($signed(_zz_17825) >>> _zz_1574);
  assign _zz_17825 = _zz_17826;
  assign _zz_17826 = ($signed(_zz_17828) - $signed(_zz_1572));
  assign _zz_17827 = ({8'd0,data_mid_106_imag} <<< 8);
  assign _zz_17828 = {{8{_zz_17827[23]}}, _zz_17827};
  assign _zz_17829 = fixTo_1887_dout;
  assign _zz_17830 = _zz_17831[31 : 0];
  assign _zz_17831 = _zz_17832;
  assign _zz_17832 = ($signed(_zz_17833) >>> _zz_1575);
  assign _zz_17833 = _zz_17834;
  assign _zz_17834 = ($signed(_zz_17836) + $signed(_zz_1571));
  assign _zz_17835 = ({8'd0,data_mid_106_real} <<< 8);
  assign _zz_17836 = {{8{_zz_17835[23]}}, _zz_17835};
  assign _zz_17837 = fixTo_1888_dout;
  assign _zz_17838 = _zz_17839[31 : 0];
  assign _zz_17839 = _zz_17840;
  assign _zz_17840 = ($signed(_zz_17841) >>> _zz_1575);
  assign _zz_17841 = _zz_17842;
  assign _zz_17842 = ($signed(_zz_17844) + $signed(_zz_1572));
  assign _zz_17843 = ({8'd0,data_mid_106_imag} <<< 8);
  assign _zz_17844 = {{8{_zz_17843[23]}}, _zz_17843};
  assign _zz_17845 = fixTo_1889_dout;
  assign _zz_17846 = ($signed(twiddle_factor_table_26_real) + $signed(twiddle_factor_table_26_imag));
  assign _zz_17847 = ($signed(_zz_1578) - $signed(_zz_17848));
  assign _zz_17848 = ($signed(_zz_17849) * $signed(twiddle_factor_table_26_imag));
  assign _zz_17849 = ($signed(data_mid_123_real) + $signed(data_mid_123_imag));
  assign _zz_17850 = fixTo_1890_dout;
  assign _zz_17851 = ($signed(_zz_1578) + $signed(_zz_17852));
  assign _zz_17852 = ($signed(_zz_17853) * $signed(twiddle_factor_table_26_real));
  assign _zz_17853 = ($signed(data_mid_123_imag) - $signed(data_mid_123_real));
  assign _zz_17854 = fixTo_1891_dout;
  assign _zz_17855 = _zz_17856[31 : 0];
  assign _zz_17856 = _zz_17857;
  assign _zz_17857 = ($signed(_zz_17858) >>> _zz_1579);
  assign _zz_17858 = _zz_17859;
  assign _zz_17859 = ($signed(_zz_17861) - $signed(_zz_1576));
  assign _zz_17860 = ({8'd0,data_mid_107_real} <<< 8);
  assign _zz_17861 = {{8{_zz_17860[23]}}, _zz_17860};
  assign _zz_17862 = fixTo_1892_dout;
  assign _zz_17863 = _zz_17864[31 : 0];
  assign _zz_17864 = _zz_17865;
  assign _zz_17865 = ($signed(_zz_17866) >>> _zz_1579);
  assign _zz_17866 = _zz_17867;
  assign _zz_17867 = ($signed(_zz_17869) - $signed(_zz_1577));
  assign _zz_17868 = ({8'd0,data_mid_107_imag} <<< 8);
  assign _zz_17869 = {{8{_zz_17868[23]}}, _zz_17868};
  assign _zz_17870 = fixTo_1893_dout;
  assign _zz_17871 = _zz_17872[31 : 0];
  assign _zz_17872 = _zz_17873;
  assign _zz_17873 = ($signed(_zz_17874) >>> _zz_1580);
  assign _zz_17874 = _zz_17875;
  assign _zz_17875 = ($signed(_zz_17877) + $signed(_zz_1576));
  assign _zz_17876 = ({8'd0,data_mid_107_real} <<< 8);
  assign _zz_17877 = {{8{_zz_17876[23]}}, _zz_17876};
  assign _zz_17878 = fixTo_1894_dout;
  assign _zz_17879 = _zz_17880[31 : 0];
  assign _zz_17880 = _zz_17881;
  assign _zz_17881 = ($signed(_zz_17882) >>> _zz_1580);
  assign _zz_17882 = _zz_17883;
  assign _zz_17883 = ($signed(_zz_17885) + $signed(_zz_1577));
  assign _zz_17884 = ({8'd0,data_mid_107_imag} <<< 8);
  assign _zz_17885 = {{8{_zz_17884[23]}}, _zz_17884};
  assign _zz_17886 = fixTo_1895_dout;
  assign _zz_17887 = ($signed(twiddle_factor_table_27_real) + $signed(twiddle_factor_table_27_imag));
  assign _zz_17888 = ($signed(_zz_1583) - $signed(_zz_17889));
  assign _zz_17889 = ($signed(_zz_17890) * $signed(twiddle_factor_table_27_imag));
  assign _zz_17890 = ($signed(data_mid_124_real) + $signed(data_mid_124_imag));
  assign _zz_17891 = fixTo_1896_dout;
  assign _zz_17892 = ($signed(_zz_1583) + $signed(_zz_17893));
  assign _zz_17893 = ($signed(_zz_17894) * $signed(twiddle_factor_table_27_real));
  assign _zz_17894 = ($signed(data_mid_124_imag) - $signed(data_mid_124_real));
  assign _zz_17895 = fixTo_1897_dout;
  assign _zz_17896 = _zz_17897[31 : 0];
  assign _zz_17897 = _zz_17898;
  assign _zz_17898 = ($signed(_zz_17899) >>> _zz_1584);
  assign _zz_17899 = _zz_17900;
  assign _zz_17900 = ($signed(_zz_17902) - $signed(_zz_1581));
  assign _zz_17901 = ({8'd0,data_mid_108_real} <<< 8);
  assign _zz_17902 = {{8{_zz_17901[23]}}, _zz_17901};
  assign _zz_17903 = fixTo_1898_dout;
  assign _zz_17904 = _zz_17905[31 : 0];
  assign _zz_17905 = _zz_17906;
  assign _zz_17906 = ($signed(_zz_17907) >>> _zz_1584);
  assign _zz_17907 = _zz_17908;
  assign _zz_17908 = ($signed(_zz_17910) - $signed(_zz_1582));
  assign _zz_17909 = ({8'd0,data_mid_108_imag} <<< 8);
  assign _zz_17910 = {{8{_zz_17909[23]}}, _zz_17909};
  assign _zz_17911 = fixTo_1899_dout;
  assign _zz_17912 = _zz_17913[31 : 0];
  assign _zz_17913 = _zz_17914;
  assign _zz_17914 = ($signed(_zz_17915) >>> _zz_1585);
  assign _zz_17915 = _zz_17916;
  assign _zz_17916 = ($signed(_zz_17918) + $signed(_zz_1581));
  assign _zz_17917 = ({8'd0,data_mid_108_real} <<< 8);
  assign _zz_17918 = {{8{_zz_17917[23]}}, _zz_17917};
  assign _zz_17919 = fixTo_1900_dout;
  assign _zz_17920 = _zz_17921[31 : 0];
  assign _zz_17921 = _zz_17922;
  assign _zz_17922 = ($signed(_zz_17923) >>> _zz_1585);
  assign _zz_17923 = _zz_17924;
  assign _zz_17924 = ($signed(_zz_17926) + $signed(_zz_1582));
  assign _zz_17925 = ({8'd0,data_mid_108_imag} <<< 8);
  assign _zz_17926 = {{8{_zz_17925[23]}}, _zz_17925};
  assign _zz_17927 = fixTo_1901_dout;
  assign _zz_17928 = ($signed(twiddle_factor_table_28_real) + $signed(twiddle_factor_table_28_imag));
  assign _zz_17929 = ($signed(_zz_1588) - $signed(_zz_17930));
  assign _zz_17930 = ($signed(_zz_17931) * $signed(twiddle_factor_table_28_imag));
  assign _zz_17931 = ($signed(data_mid_125_real) + $signed(data_mid_125_imag));
  assign _zz_17932 = fixTo_1902_dout;
  assign _zz_17933 = ($signed(_zz_1588) + $signed(_zz_17934));
  assign _zz_17934 = ($signed(_zz_17935) * $signed(twiddle_factor_table_28_real));
  assign _zz_17935 = ($signed(data_mid_125_imag) - $signed(data_mid_125_real));
  assign _zz_17936 = fixTo_1903_dout;
  assign _zz_17937 = _zz_17938[31 : 0];
  assign _zz_17938 = _zz_17939;
  assign _zz_17939 = ($signed(_zz_17940) >>> _zz_1589);
  assign _zz_17940 = _zz_17941;
  assign _zz_17941 = ($signed(_zz_17943) - $signed(_zz_1586));
  assign _zz_17942 = ({8'd0,data_mid_109_real} <<< 8);
  assign _zz_17943 = {{8{_zz_17942[23]}}, _zz_17942};
  assign _zz_17944 = fixTo_1904_dout;
  assign _zz_17945 = _zz_17946[31 : 0];
  assign _zz_17946 = _zz_17947;
  assign _zz_17947 = ($signed(_zz_17948) >>> _zz_1589);
  assign _zz_17948 = _zz_17949;
  assign _zz_17949 = ($signed(_zz_17951) - $signed(_zz_1587));
  assign _zz_17950 = ({8'd0,data_mid_109_imag} <<< 8);
  assign _zz_17951 = {{8{_zz_17950[23]}}, _zz_17950};
  assign _zz_17952 = fixTo_1905_dout;
  assign _zz_17953 = _zz_17954[31 : 0];
  assign _zz_17954 = _zz_17955;
  assign _zz_17955 = ($signed(_zz_17956) >>> _zz_1590);
  assign _zz_17956 = _zz_17957;
  assign _zz_17957 = ($signed(_zz_17959) + $signed(_zz_1586));
  assign _zz_17958 = ({8'd0,data_mid_109_real} <<< 8);
  assign _zz_17959 = {{8{_zz_17958[23]}}, _zz_17958};
  assign _zz_17960 = fixTo_1906_dout;
  assign _zz_17961 = _zz_17962[31 : 0];
  assign _zz_17962 = _zz_17963;
  assign _zz_17963 = ($signed(_zz_17964) >>> _zz_1590);
  assign _zz_17964 = _zz_17965;
  assign _zz_17965 = ($signed(_zz_17967) + $signed(_zz_1587));
  assign _zz_17966 = ({8'd0,data_mid_109_imag} <<< 8);
  assign _zz_17967 = {{8{_zz_17966[23]}}, _zz_17966};
  assign _zz_17968 = fixTo_1907_dout;
  assign _zz_17969 = ($signed(twiddle_factor_table_29_real) + $signed(twiddle_factor_table_29_imag));
  assign _zz_17970 = ($signed(_zz_1593) - $signed(_zz_17971));
  assign _zz_17971 = ($signed(_zz_17972) * $signed(twiddle_factor_table_29_imag));
  assign _zz_17972 = ($signed(data_mid_126_real) + $signed(data_mid_126_imag));
  assign _zz_17973 = fixTo_1908_dout;
  assign _zz_17974 = ($signed(_zz_1593) + $signed(_zz_17975));
  assign _zz_17975 = ($signed(_zz_17976) * $signed(twiddle_factor_table_29_real));
  assign _zz_17976 = ($signed(data_mid_126_imag) - $signed(data_mid_126_real));
  assign _zz_17977 = fixTo_1909_dout;
  assign _zz_17978 = _zz_17979[31 : 0];
  assign _zz_17979 = _zz_17980;
  assign _zz_17980 = ($signed(_zz_17981) >>> _zz_1594);
  assign _zz_17981 = _zz_17982;
  assign _zz_17982 = ($signed(_zz_17984) - $signed(_zz_1591));
  assign _zz_17983 = ({8'd0,data_mid_110_real} <<< 8);
  assign _zz_17984 = {{8{_zz_17983[23]}}, _zz_17983};
  assign _zz_17985 = fixTo_1910_dout;
  assign _zz_17986 = _zz_17987[31 : 0];
  assign _zz_17987 = _zz_17988;
  assign _zz_17988 = ($signed(_zz_17989) >>> _zz_1594);
  assign _zz_17989 = _zz_17990;
  assign _zz_17990 = ($signed(_zz_17992) - $signed(_zz_1592));
  assign _zz_17991 = ({8'd0,data_mid_110_imag} <<< 8);
  assign _zz_17992 = {{8{_zz_17991[23]}}, _zz_17991};
  assign _zz_17993 = fixTo_1911_dout;
  assign _zz_17994 = _zz_17995[31 : 0];
  assign _zz_17995 = _zz_17996;
  assign _zz_17996 = ($signed(_zz_17997) >>> _zz_1595);
  assign _zz_17997 = _zz_17998;
  assign _zz_17998 = ($signed(_zz_18000) + $signed(_zz_1591));
  assign _zz_17999 = ({8'd0,data_mid_110_real} <<< 8);
  assign _zz_18000 = {{8{_zz_17999[23]}}, _zz_17999};
  assign _zz_18001 = fixTo_1912_dout;
  assign _zz_18002 = _zz_18003[31 : 0];
  assign _zz_18003 = _zz_18004;
  assign _zz_18004 = ($signed(_zz_18005) >>> _zz_1595);
  assign _zz_18005 = _zz_18006;
  assign _zz_18006 = ($signed(_zz_18008) + $signed(_zz_1592));
  assign _zz_18007 = ({8'd0,data_mid_110_imag} <<< 8);
  assign _zz_18008 = {{8{_zz_18007[23]}}, _zz_18007};
  assign _zz_18009 = fixTo_1913_dout;
  assign _zz_18010 = ($signed(twiddle_factor_table_30_real) + $signed(twiddle_factor_table_30_imag));
  assign _zz_18011 = ($signed(_zz_1598) - $signed(_zz_18012));
  assign _zz_18012 = ($signed(_zz_18013) * $signed(twiddle_factor_table_30_imag));
  assign _zz_18013 = ($signed(data_mid_127_real) + $signed(data_mid_127_imag));
  assign _zz_18014 = fixTo_1914_dout;
  assign _zz_18015 = ($signed(_zz_1598) + $signed(_zz_18016));
  assign _zz_18016 = ($signed(_zz_18017) * $signed(twiddle_factor_table_30_real));
  assign _zz_18017 = ($signed(data_mid_127_imag) - $signed(data_mid_127_real));
  assign _zz_18018 = fixTo_1915_dout;
  assign _zz_18019 = _zz_18020[31 : 0];
  assign _zz_18020 = _zz_18021;
  assign _zz_18021 = ($signed(_zz_18022) >>> _zz_1599);
  assign _zz_18022 = _zz_18023;
  assign _zz_18023 = ($signed(_zz_18025) - $signed(_zz_1596));
  assign _zz_18024 = ({8'd0,data_mid_111_real} <<< 8);
  assign _zz_18025 = {{8{_zz_18024[23]}}, _zz_18024};
  assign _zz_18026 = fixTo_1916_dout;
  assign _zz_18027 = _zz_18028[31 : 0];
  assign _zz_18028 = _zz_18029;
  assign _zz_18029 = ($signed(_zz_18030) >>> _zz_1599);
  assign _zz_18030 = _zz_18031;
  assign _zz_18031 = ($signed(_zz_18033) - $signed(_zz_1597));
  assign _zz_18032 = ({8'd0,data_mid_111_imag} <<< 8);
  assign _zz_18033 = {{8{_zz_18032[23]}}, _zz_18032};
  assign _zz_18034 = fixTo_1917_dout;
  assign _zz_18035 = _zz_18036[31 : 0];
  assign _zz_18036 = _zz_18037;
  assign _zz_18037 = ($signed(_zz_18038) >>> _zz_1600);
  assign _zz_18038 = _zz_18039;
  assign _zz_18039 = ($signed(_zz_18041) + $signed(_zz_1596));
  assign _zz_18040 = ({8'd0,data_mid_111_real} <<< 8);
  assign _zz_18041 = {{8{_zz_18040[23]}}, _zz_18040};
  assign _zz_18042 = fixTo_1918_dout;
  assign _zz_18043 = _zz_18044[31 : 0];
  assign _zz_18044 = _zz_18045;
  assign _zz_18045 = ($signed(_zz_18046) >>> _zz_1600);
  assign _zz_18046 = _zz_18047;
  assign _zz_18047 = ($signed(_zz_18049) + $signed(_zz_1597));
  assign _zz_18048 = ({8'd0,data_mid_111_imag} <<< 8);
  assign _zz_18049 = {{8{_zz_18048[23]}}, _zz_18048};
  assign _zz_18050 = fixTo_1919_dout;
  assign _zz_18051 = ($signed(twiddle_factor_table_31_real) + $signed(twiddle_factor_table_31_imag));
  assign _zz_18052 = ($signed(_zz_1603) - $signed(_zz_18053));
  assign _zz_18053 = ($signed(_zz_18054) * $signed(twiddle_factor_table_31_imag));
  assign _zz_18054 = ($signed(data_mid_32_real) + $signed(data_mid_32_imag));
  assign _zz_18055 = fixTo_1920_dout;
  assign _zz_18056 = ($signed(_zz_1603) + $signed(_zz_18057));
  assign _zz_18057 = ($signed(_zz_18058) * $signed(twiddle_factor_table_31_real));
  assign _zz_18058 = ($signed(data_mid_32_imag) - $signed(data_mid_32_real));
  assign _zz_18059 = fixTo_1921_dout;
  assign _zz_18060 = _zz_18061[31 : 0];
  assign _zz_18061 = _zz_18062;
  assign _zz_18062 = ($signed(_zz_18063) >>> _zz_1604);
  assign _zz_18063 = _zz_18064;
  assign _zz_18064 = ($signed(_zz_18066) - $signed(_zz_1601));
  assign _zz_18065 = ({8'd0,data_mid_0_real} <<< 8);
  assign _zz_18066 = {{8{_zz_18065[23]}}, _zz_18065};
  assign _zz_18067 = fixTo_1922_dout;
  assign _zz_18068 = _zz_18069[31 : 0];
  assign _zz_18069 = _zz_18070;
  assign _zz_18070 = ($signed(_zz_18071) >>> _zz_1604);
  assign _zz_18071 = _zz_18072;
  assign _zz_18072 = ($signed(_zz_18074) - $signed(_zz_1602));
  assign _zz_18073 = ({8'd0,data_mid_0_imag} <<< 8);
  assign _zz_18074 = {{8{_zz_18073[23]}}, _zz_18073};
  assign _zz_18075 = fixTo_1923_dout;
  assign _zz_18076 = _zz_18077[31 : 0];
  assign _zz_18077 = _zz_18078;
  assign _zz_18078 = ($signed(_zz_18079) >>> _zz_1605);
  assign _zz_18079 = _zz_18080;
  assign _zz_18080 = ($signed(_zz_18082) + $signed(_zz_1601));
  assign _zz_18081 = ({8'd0,data_mid_0_real} <<< 8);
  assign _zz_18082 = {{8{_zz_18081[23]}}, _zz_18081};
  assign _zz_18083 = fixTo_1924_dout;
  assign _zz_18084 = _zz_18085[31 : 0];
  assign _zz_18085 = _zz_18086;
  assign _zz_18086 = ($signed(_zz_18087) >>> _zz_1605);
  assign _zz_18087 = _zz_18088;
  assign _zz_18088 = ($signed(_zz_18090) + $signed(_zz_1602));
  assign _zz_18089 = ({8'd0,data_mid_0_imag} <<< 8);
  assign _zz_18090 = {{8{_zz_18089[23]}}, _zz_18089};
  assign _zz_18091 = fixTo_1925_dout;
  assign _zz_18092 = ($signed(twiddle_factor_table_32_real) + $signed(twiddle_factor_table_32_imag));
  assign _zz_18093 = ($signed(_zz_1608) - $signed(_zz_18094));
  assign _zz_18094 = ($signed(_zz_18095) * $signed(twiddle_factor_table_32_imag));
  assign _zz_18095 = ($signed(data_mid_33_real) + $signed(data_mid_33_imag));
  assign _zz_18096 = fixTo_1926_dout;
  assign _zz_18097 = ($signed(_zz_1608) + $signed(_zz_18098));
  assign _zz_18098 = ($signed(_zz_18099) * $signed(twiddle_factor_table_32_real));
  assign _zz_18099 = ($signed(data_mid_33_imag) - $signed(data_mid_33_real));
  assign _zz_18100 = fixTo_1927_dout;
  assign _zz_18101 = _zz_18102[31 : 0];
  assign _zz_18102 = _zz_18103;
  assign _zz_18103 = ($signed(_zz_18104) >>> _zz_1609);
  assign _zz_18104 = _zz_18105;
  assign _zz_18105 = ($signed(_zz_18107) - $signed(_zz_1606));
  assign _zz_18106 = ({8'd0,data_mid_1_real} <<< 8);
  assign _zz_18107 = {{8{_zz_18106[23]}}, _zz_18106};
  assign _zz_18108 = fixTo_1928_dout;
  assign _zz_18109 = _zz_18110[31 : 0];
  assign _zz_18110 = _zz_18111;
  assign _zz_18111 = ($signed(_zz_18112) >>> _zz_1609);
  assign _zz_18112 = _zz_18113;
  assign _zz_18113 = ($signed(_zz_18115) - $signed(_zz_1607));
  assign _zz_18114 = ({8'd0,data_mid_1_imag} <<< 8);
  assign _zz_18115 = {{8{_zz_18114[23]}}, _zz_18114};
  assign _zz_18116 = fixTo_1929_dout;
  assign _zz_18117 = _zz_18118[31 : 0];
  assign _zz_18118 = _zz_18119;
  assign _zz_18119 = ($signed(_zz_18120) >>> _zz_1610);
  assign _zz_18120 = _zz_18121;
  assign _zz_18121 = ($signed(_zz_18123) + $signed(_zz_1606));
  assign _zz_18122 = ({8'd0,data_mid_1_real} <<< 8);
  assign _zz_18123 = {{8{_zz_18122[23]}}, _zz_18122};
  assign _zz_18124 = fixTo_1930_dout;
  assign _zz_18125 = _zz_18126[31 : 0];
  assign _zz_18126 = _zz_18127;
  assign _zz_18127 = ($signed(_zz_18128) >>> _zz_1610);
  assign _zz_18128 = _zz_18129;
  assign _zz_18129 = ($signed(_zz_18131) + $signed(_zz_1607));
  assign _zz_18130 = ({8'd0,data_mid_1_imag} <<< 8);
  assign _zz_18131 = {{8{_zz_18130[23]}}, _zz_18130};
  assign _zz_18132 = fixTo_1931_dout;
  assign _zz_18133 = ($signed(twiddle_factor_table_33_real) + $signed(twiddle_factor_table_33_imag));
  assign _zz_18134 = ($signed(_zz_1613) - $signed(_zz_18135));
  assign _zz_18135 = ($signed(_zz_18136) * $signed(twiddle_factor_table_33_imag));
  assign _zz_18136 = ($signed(data_mid_34_real) + $signed(data_mid_34_imag));
  assign _zz_18137 = fixTo_1932_dout;
  assign _zz_18138 = ($signed(_zz_1613) + $signed(_zz_18139));
  assign _zz_18139 = ($signed(_zz_18140) * $signed(twiddle_factor_table_33_real));
  assign _zz_18140 = ($signed(data_mid_34_imag) - $signed(data_mid_34_real));
  assign _zz_18141 = fixTo_1933_dout;
  assign _zz_18142 = _zz_18143[31 : 0];
  assign _zz_18143 = _zz_18144;
  assign _zz_18144 = ($signed(_zz_18145) >>> _zz_1614);
  assign _zz_18145 = _zz_18146;
  assign _zz_18146 = ($signed(_zz_18148) - $signed(_zz_1611));
  assign _zz_18147 = ({8'd0,data_mid_2_real} <<< 8);
  assign _zz_18148 = {{8{_zz_18147[23]}}, _zz_18147};
  assign _zz_18149 = fixTo_1934_dout;
  assign _zz_18150 = _zz_18151[31 : 0];
  assign _zz_18151 = _zz_18152;
  assign _zz_18152 = ($signed(_zz_18153) >>> _zz_1614);
  assign _zz_18153 = _zz_18154;
  assign _zz_18154 = ($signed(_zz_18156) - $signed(_zz_1612));
  assign _zz_18155 = ({8'd0,data_mid_2_imag} <<< 8);
  assign _zz_18156 = {{8{_zz_18155[23]}}, _zz_18155};
  assign _zz_18157 = fixTo_1935_dout;
  assign _zz_18158 = _zz_18159[31 : 0];
  assign _zz_18159 = _zz_18160;
  assign _zz_18160 = ($signed(_zz_18161) >>> _zz_1615);
  assign _zz_18161 = _zz_18162;
  assign _zz_18162 = ($signed(_zz_18164) + $signed(_zz_1611));
  assign _zz_18163 = ({8'd0,data_mid_2_real} <<< 8);
  assign _zz_18164 = {{8{_zz_18163[23]}}, _zz_18163};
  assign _zz_18165 = fixTo_1936_dout;
  assign _zz_18166 = _zz_18167[31 : 0];
  assign _zz_18167 = _zz_18168;
  assign _zz_18168 = ($signed(_zz_18169) >>> _zz_1615);
  assign _zz_18169 = _zz_18170;
  assign _zz_18170 = ($signed(_zz_18172) + $signed(_zz_1612));
  assign _zz_18171 = ({8'd0,data_mid_2_imag} <<< 8);
  assign _zz_18172 = {{8{_zz_18171[23]}}, _zz_18171};
  assign _zz_18173 = fixTo_1937_dout;
  assign _zz_18174 = ($signed(twiddle_factor_table_34_real) + $signed(twiddle_factor_table_34_imag));
  assign _zz_18175 = ($signed(_zz_1618) - $signed(_zz_18176));
  assign _zz_18176 = ($signed(_zz_18177) * $signed(twiddle_factor_table_34_imag));
  assign _zz_18177 = ($signed(data_mid_35_real) + $signed(data_mid_35_imag));
  assign _zz_18178 = fixTo_1938_dout;
  assign _zz_18179 = ($signed(_zz_1618) + $signed(_zz_18180));
  assign _zz_18180 = ($signed(_zz_18181) * $signed(twiddle_factor_table_34_real));
  assign _zz_18181 = ($signed(data_mid_35_imag) - $signed(data_mid_35_real));
  assign _zz_18182 = fixTo_1939_dout;
  assign _zz_18183 = _zz_18184[31 : 0];
  assign _zz_18184 = _zz_18185;
  assign _zz_18185 = ($signed(_zz_18186) >>> _zz_1619);
  assign _zz_18186 = _zz_18187;
  assign _zz_18187 = ($signed(_zz_18189) - $signed(_zz_1616));
  assign _zz_18188 = ({8'd0,data_mid_3_real} <<< 8);
  assign _zz_18189 = {{8{_zz_18188[23]}}, _zz_18188};
  assign _zz_18190 = fixTo_1940_dout;
  assign _zz_18191 = _zz_18192[31 : 0];
  assign _zz_18192 = _zz_18193;
  assign _zz_18193 = ($signed(_zz_18194) >>> _zz_1619);
  assign _zz_18194 = _zz_18195;
  assign _zz_18195 = ($signed(_zz_18197) - $signed(_zz_1617));
  assign _zz_18196 = ({8'd0,data_mid_3_imag} <<< 8);
  assign _zz_18197 = {{8{_zz_18196[23]}}, _zz_18196};
  assign _zz_18198 = fixTo_1941_dout;
  assign _zz_18199 = _zz_18200[31 : 0];
  assign _zz_18200 = _zz_18201;
  assign _zz_18201 = ($signed(_zz_18202) >>> _zz_1620);
  assign _zz_18202 = _zz_18203;
  assign _zz_18203 = ($signed(_zz_18205) + $signed(_zz_1616));
  assign _zz_18204 = ({8'd0,data_mid_3_real} <<< 8);
  assign _zz_18205 = {{8{_zz_18204[23]}}, _zz_18204};
  assign _zz_18206 = fixTo_1942_dout;
  assign _zz_18207 = _zz_18208[31 : 0];
  assign _zz_18208 = _zz_18209;
  assign _zz_18209 = ($signed(_zz_18210) >>> _zz_1620);
  assign _zz_18210 = _zz_18211;
  assign _zz_18211 = ($signed(_zz_18213) + $signed(_zz_1617));
  assign _zz_18212 = ({8'd0,data_mid_3_imag} <<< 8);
  assign _zz_18213 = {{8{_zz_18212[23]}}, _zz_18212};
  assign _zz_18214 = fixTo_1943_dout;
  assign _zz_18215 = ($signed(twiddle_factor_table_35_real) + $signed(twiddle_factor_table_35_imag));
  assign _zz_18216 = ($signed(_zz_1623) - $signed(_zz_18217));
  assign _zz_18217 = ($signed(_zz_18218) * $signed(twiddle_factor_table_35_imag));
  assign _zz_18218 = ($signed(data_mid_36_real) + $signed(data_mid_36_imag));
  assign _zz_18219 = fixTo_1944_dout;
  assign _zz_18220 = ($signed(_zz_1623) + $signed(_zz_18221));
  assign _zz_18221 = ($signed(_zz_18222) * $signed(twiddle_factor_table_35_real));
  assign _zz_18222 = ($signed(data_mid_36_imag) - $signed(data_mid_36_real));
  assign _zz_18223 = fixTo_1945_dout;
  assign _zz_18224 = _zz_18225[31 : 0];
  assign _zz_18225 = _zz_18226;
  assign _zz_18226 = ($signed(_zz_18227) >>> _zz_1624);
  assign _zz_18227 = _zz_18228;
  assign _zz_18228 = ($signed(_zz_18230) - $signed(_zz_1621));
  assign _zz_18229 = ({8'd0,data_mid_4_real} <<< 8);
  assign _zz_18230 = {{8{_zz_18229[23]}}, _zz_18229};
  assign _zz_18231 = fixTo_1946_dout;
  assign _zz_18232 = _zz_18233[31 : 0];
  assign _zz_18233 = _zz_18234;
  assign _zz_18234 = ($signed(_zz_18235) >>> _zz_1624);
  assign _zz_18235 = _zz_18236;
  assign _zz_18236 = ($signed(_zz_18238) - $signed(_zz_1622));
  assign _zz_18237 = ({8'd0,data_mid_4_imag} <<< 8);
  assign _zz_18238 = {{8{_zz_18237[23]}}, _zz_18237};
  assign _zz_18239 = fixTo_1947_dout;
  assign _zz_18240 = _zz_18241[31 : 0];
  assign _zz_18241 = _zz_18242;
  assign _zz_18242 = ($signed(_zz_18243) >>> _zz_1625);
  assign _zz_18243 = _zz_18244;
  assign _zz_18244 = ($signed(_zz_18246) + $signed(_zz_1621));
  assign _zz_18245 = ({8'd0,data_mid_4_real} <<< 8);
  assign _zz_18246 = {{8{_zz_18245[23]}}, _zz_18245};
  assign _zz_18247 = fixTo_1948_dout;
  assign _zz_18248 = _zz_18249[31 : 0];
  assign _zz_18249 = _zz_18250;
  assign _zz_18250 = ($signed(_zz_18251) >>> _zz_1625);
  assign _zz_18251 = _zz_18252;
  assign _zz_18252 = ($signed(_zz_18254) + $signed(_zz_1622));
  assign _zz_18253 = ({8'd0,data_mid_4_imag} <<< 8);
  assign _zz_18254 = {{8{_zz_18253[23]}}, _zz_18253};
  assign _zz_18255 = fixTo_1949_dout;
  assign _zz_18256 = ($signed(twiddle_factor_table_36_real) + $signed(twiddle_factor_table_36_imag));
  assign _zz_18257 = ($signed(_zz_1628) - $signed(_zz_18258));
  assign _zz_18258 = ($signed(_zz_18259) * $signed(twiddle_factor_table_36_imag));
  assign _zz_18259 = ($signed(data_mid_37_real) + $signed(data_mid_37_imag));
  assign _zz_18260 = fixTo_1950_dout;
  assign _zz_18261 = ($signed(_zz_1628) + $signed(_zz_18262));
  assign _zz_18262 = ($signed(_zz_18263) * $signed(twiddle_factor_table_36_real));
  assign _zz_18263 = ($signed(data_mid_37_imag) - $signed(data_mid_37_real));
  assign _zz_18264 = fixTo_1951_dout;
  assign _zz_18265 = _zz_18266[31 : 0];
  assign _zz_18266 = _zz_18267;
  assign _zz_18267 = ($signed(_zz_18268) >>> _zz_1629);
  assign _zz_18268 = _zz_18269;
  assign _zz_18269 = ($signed(_zz_18271) - $signed(_zz_1626));
  assign _zz_18270 = ({8'd0,data_mid_5_real} <<< 8);
  assign _zz_18271 = {{8{_zz_18270[23]}}, _zz_18270};
  assign _zz_18272 = fixTo_1952_dout;
  assign _zz_18273 = _zz_18274[31 : 0];
  assign _zz_18274 = _zz_18275;
  assign _zz_18275 = ($signed(_zz_18276) >>> _zz_1629);
  assign _zz_18276 = _zz_18277;
  assign _zz_18277 = ($signed(_zz_18279) - $signed(_zz_1627));
  assign _zz_18278 = ({8'd0,data_mid_5_imag} <<< 8);
  assign _zz_18279 = {{8{_zz_18278[23]}}, _zz_18278};
  assign _zz_18280 = fixTo_1953_dout;
  assign _zz_18281 = _zz_18282[31 : 0];
  assign _zz_18282 = _zz_18283;
  assign _zz_18283 = ($signed(_zz_18284) >>> _zz_1630);
  assign _zz_18284 = _zz_18285;
  assign _zz_18285 = ($signed(_zz_18287) + $signed(_zz_1626));
  assign _zz_18286 = ({8'd0,data_mid_5_real} <<< 8);
  assign _zz_18287 = {{8{_zz_18286[23]}}, _zz_18286};
  assign _zz_18288 = fixTo_1954_dout;
  assign _zz_18289 = _zz_18290[31 : 0];
  assign _zz_18290 = _zz_18291;
  assign _zz_18291 = ($signed(_zz_18292) >>> _zz_1630);
  assign _zz_18292 = _zz_18293;
  assign _zz_18293 = ($signed(_zz_18295) + $signed(_zz_1627));
  assign _zz_18294 = ({8'd0,data_mid_5_imag} <<< 8);
  assign _zz_18295 = {{8{_zz_18294[23]}}, _zz_18294};
  assign _zz_18296 = fixTo_1955_dout;
  assign _zz_18297 = ($signed(twiddle_factor_table_37_real) + $signed(twiddle_factor_table_37_imag));
  assign _zz_18298 = ($signed(_zz_1633) - $signed(_zz_18299));
  assign _zz_18299 = ($signed(_zz_18300) * $signed(twiddle_factor_table_37_imag));
  assign _zz_18300 = ($signed(data_mid_38_real) + $signed(data_mid_38_imag));
  assign _zz_18301 = fixTo_1956_dout;
  assign _zz_18302 = ($signed(_zz_1633) + $signed(_zz_18303));
  assign _zz_18303 = ($signed(_zz_18304) * $signed(twiddle_factor_table_37_real));
  assign _zz_18304 = ($signed(data_mid_38_imag) - $signed(data_mid_38_real));
  assign _zz_18305 = fixTo_1957_dout;
  assign _zz_18306 = _zz_18307[31 : 0];
  assign _zz_18307 = _zz_18308;
  assign _zz_18308 = ($signed(_zz_18309) >>> _zz_1634);
  assign _zz_18309 = _zz_18310;
  assign _zz_18310 = ($signed(_zz_18312) - $signed(_zz_1631));
  assign _zz_18311 = ({8'd0,data_mid_6_real} <<< 8);
  assign _zz_18312 = {{8{_zz_18311[23]}}, _zz_18311};
  assign _zz_18313 = fixTo_1958_dout;
  assign _zz_18314 = _zz_18315[31 : 0];
  assign _zz_18315 = _zz_18316;
  assign _zz_18316 = ($signed(_zz_18317) >>> _zz_1634);
  assign _zz_18317 = _zz_18318;
  assign _zz_18318 = ($signed(_zz_18320) - $signed(_zz_1632));
  assign _zz_18319 = ({8'd0,data_mid_6_imag} <<< 8);
  assign _zz_18320 = {{8{_zz_18319[23]}}, _zz_18319};
  assign _zz_18321 = fixTo_1959_dout;
  assign _zz_18322 = _zz_18323[31 : 0];
  assign _zz_18323 = _zz_18324;
  assign _zz_18324 = ($signed(_zz_18325) >>> _zz_1635);
  assign _zz_18325 = _zz_18326;
  assign _zz_18326 = ($signed(_zz_18328) + $signed(_zz_1631));
  assign _zz_18327 = ({8'd0,data_mid_6_real} <<< 8);
  assign _zz_18328 = {{8{_zz_18327[23]}}, _zz_18327};
  assign _zz_18329 = fixTo_1960_dout;
  assign _zz_18330 = _zz_18331[31 : 0];
  assign _zz_18331 = _zz_18332;
  assign _zz_18332 = ($signed(_zz_18333) >>> _zz_1635);
  assign _zz_18333 = _zz_18334;
  assign _zz_18334 = ($signed(_zz_18336) + $signed(_zz_1632));
  assign _zz_18335 = ({8'd0,data_mid_6_imag} <<< 8);
  assign _zz_18336 = {{8{_zz_18335[23]}}, _zz_18335};
  assign _zz_18337 = fixTo_1961_dout;
  assign _zz_18338 = ($signed(twiddle_factor_table_38_real) + $signed(twiddle_factor_table_38_imag));
  assign _zz_18339 = ($signed(_zz_1638) - $signed(_zz_18340));
  assign _zz_18340 = ($signed(_zz_18341) * $signed(twiddle_factor_table_38_imag));
  assign _zz_18341 = ($signed(data_mid_39_real) + $signed(data_mid_39_imag));
  assign _zz_18342 = fixTo_1962_dout;
  assign _zz_18343 = ($signed(_zz_1638) + $signed(_zz_18344));
  assign _zz_18344 = ($signed(_zz_18345) * $signed(twiddle_factor_table_38_real));
  assign _zz_18345 = ($signed(data_mid_39_imag) - $signed(data_mid_39_real));
  assign _zz_18346 = fixTo_1963_dout;
  assign _zz_18347 = _zz_18348[31 : 0];
  assign _zz_18348 = _zz_18349;
  assign _zz_18349 = ($signed(_zz_18350) >>> _zz_1639);
  assign _zz_18350 = _zz_18351;
  assign _zz_18351 = ($signed(_zz_18353) - $signed(_zz_1636));
  assign _zz_18352 = ({8'd0,data_mid_7_real} <<< 8);
  assign _zz_18353 = {{8{_zz_18352[23]}}, _zz_18352};
  assign _zz_18354 = fixTo_1964_dout;
  assign _zz_18355 = _zz_18356[31 : 0];
  assign _zz_18356 = _zz_18357;
  assign _zz_18357 = ($signed(_zz_18358) >>> _zz_1639);
  assign _zz_18358 = _zz_18359;
  assign _zz_18359 = ($signed(_zz_18361) - $signed(_zz_1637));
  assign _zz_18360 = ({8'd0,data_mid_7_imag} <<< 8);
  assign _zz_18361 = {{8{_zz_18360[23]}}, _zz_18360};
  assign _zz_18362 = fixTo_1965_dout;
  assign _zz_18363 = _zz_18364[31 : 0];
  assign _zz_18364 = _zz_18365;
  assign _zz_18365 = ($signed(_zz_18366) >>> _zz_1640);
  assign _zz_18366 = _zz_18367;
  assign _zz_18367 = ($signed(_zz_18369) + $signed(_zz_1636));
  assign _zz_18368 = ({8'd0,data_mid_7_real} <<< 8);
  assign _zz_18369 = {{8{_zz_18368[23]}}, _zz_18368};
  assign _zz_18370 = fixTo_1966_dout;
  assign _zz_18371 = _zz_18372[31 : 0];
  assign _zz_18372 = _zz_18373;
  assign _zz_18373 = ($signed(_zz_18374) >>> _zz_1640);
  assign _zz_18374 = _zz_18375;
  assign _zz_18375 = ($signed(_zz_18377) + $signed(_zz_1637));
  assign _zz_18376 = ({8'd0,data_mid_7_imag} <<< 8);
  assign _zz_18377 = {{8{_zz_18376[23]}}, _zz_18376};
  assign _zz_18378 = fixTo_1967_dout;
  assign _zz_18379 = ($signed(twiddle_factor_table_39_real) + $signed(twiddle_factor_table_39_imag));
  assign _zz_18380 = ($signed(_zz_1643) - $signed(_zz_18381));
  assign _zz_18381 = ($signed(_zz_18382) * $signed(twiddle_factor_table_39_imag));
  assign _zz_18382 = ($signed(data_mid_40_real) + $signed(data_mid_40_imag));
  assign _zz_18383 = fixTo_1968_dout;
  assign _zz_18384 = ($signed(_zz_1643) + $signed(_zz_18385));
  assign _zz_18385 = ($signed(_zz_18386) * $signed(twiddle_factor_table_39_real));
  assign _zz_18386 = ($signed(data_mid_40_imag) - $signed(data_mid_40_real));
  assign _zz_18387 = fixTo_1969_dout;
  assign _zz_18388 = _zz_18389[31 : 0];
  assign _zz_18389 = _zz_18390;
  assign _zz_18390 = ($signed(_zz_18391) >>> _zz_1644);
  assign _zz_18391 = _zz_18392;
  assign _zz_18392 = ($signed(_zz_18394) - $signed(_zz_1641));
  assign _zz_18393 = ({8'd0,data_mid_8_real} <<< 8);
  assign _zz_18394 = {{8{_zz_18393[23]}}, _zz_18393};
  assign _zz_18395 = fixTo_1970_dout;
  assign _zz_18396 = _zz_18397[31 : 0];
  assign _zz_18397 = _zz_18398;
  assign _zz_18398 = ($signed(_zz_18399) >>> _zz_1644);
  assign _zz_18399 = _zz_18400;
  assign _zz_18400 = ($signed(_zz_18402) - $signed(_zz_1642));
  assign _zz_18401 = ({8'd0,data_mid_8_imag} <<< 8);
  assign _zz_18402 = {{8{_zz_18401[23]}}, _zz_18401};
  assign _zz_18403 = fixTo_1971_dout;
  assign _zz_18404 = _zz_18405[31 : 0];
  assign _zz_18405 = _zz_18406;
  assign _zz_18406 = ($signed(_zz_18407) >>> _zz_1645);
  assign _zz_18407 = _zz_18408;
  assign _zz_18408 = ($signed(_zz_18410) + $signed(_zz_1641));
  assign _zz_18409 = ({8'd0,data_mid_8_real} <<< 8);
  assign _zz_18410 = {{8{_zz_18409[23]}}, _zz_18409};
  assign _zz_18411 = fixTo_1972_dout;
  assign _zz_18412 = _zz_18413[31 : 0];
  assign _zz_18413 = _zz_18414;
  assign _zz_18414 = ($signed(_zz_18415) >>> _zz_1645);
  assign _zz_18415 = _zz_18416;
  assign _zz_18416 = ($signed(_zz_18418) + $signed(_zz_1642));
  assign _zz_18417 = ({8'd0,data_mid_8_imag} <<< 8);
  assign _zz_18418 = {{8{_zz_18417[23]}}, _zz_18417};
  assign _zz_18419 = fixTo_1973_dout;
  assign _zz_18420 = ($signed(twiddle_factor_table_40_real) + $signed(twiddle_factor_table_40_imag));
  assign _zz_18421 = ($signed(_zz_1648) - $signed(_zz_18422));
  assign _zz_18422 = ($signed(_zz_18423) * $signed(twiddle_factor_table_40_imag));
  assign _zz_18423 = ($signed(data_mid_41_real) + $signed(data_mid_41_imag));
  assign _zz_18424 = fixTo_1974_dout;
  assign _zz_18425 = ($signed(_zz_1648) + $signed(_zz_18426));
  assign _zz_18426 = ($signed(_zz_18427) * $signed(twiddle_factor_table_40_real));
  assign _zz_18427 = ($signed(data_mid_41_imag) - $signed(data_mid_41_real));
  assign _zz_18428 = fixTo_1975_dout;
  assign _zz_18429 = _zz_18430[31 : 0];
  assign _zz_18430 = _zz_18431;
  assign _zz_18431 = ($signed(_zz_18432) >>> _zz_1649);
  assign _zz_18432 = _zz_18433;
  assign _zz_18433 = ($signed(_zz_18435) - $signed(_zz_1646));
  assign _zz_18434 = ({8'd0,data_mid_9_real} <<< 8);
  assign _zz_18435 = {{8{_zz_18434[23]}}, _zz_18434};
  assign _zz_18436 = fixTo_1976_dout;
  assign _zz_18437 = _zz_18438[31 : 0];
  assign _zz_18438 = _zz_18439;
  assign _zz_18439 = ($signed(_zz_18440) >>> _zz_1649);
  assign _zz_18440 = _zz_18441;
  assign _zz_18441 = ($signed(_zz_18443) - $signed(_zz_1647));
  assign _zz_18442 = ({8'd0,data_mid_9_imag} <<< 8);
  assign _zz_18443 = {{8{_zz_18442[23]}}, _zz_18442};
  assign _zz_18444 = fixTo_1977_dout;
  assign _zz_18445 = _zz_18446[31 : 0];
  assign _zz_18446 = _zz_18447;
  assign _zz_18447 = ($signed(_zz_18448) >>> _zz_1650);
  assign _zz_18448 = _zz_18449;
  assign _zz_18449 = ($signed(_zz_18451) + $signed(_zz_1646));
  assign _zz_18450 = ({8'd0,data_mid_9_real} <<< 8);
  assign _zz_18451 = {{8{_zz_18450[23]}}, _zz_18450};
  assign _zz_18452 = fixTo_1978_dout;
  assign _zz_18453 = _zz_18454[31 : 0];
  assign _zz_18454 = _zz_18455;
  assign _zz_18455 = ($signed(_zz_18456) >>> _zz_1650);
  assign _zz_18456 = _zz_18457;
  assign _zz_18457 = ($signed(_zz_18459) + $signed(_zz_1647));
  assign _zz_18458 = ({8'd0,data_mid_9_imag} <<< 8);
  assign _zz_18459 = {{8{_zz_18458[23]}}, _zz_18458};
  assign _zz_18460 = fixTo_1979_dout;
  assign _zz_18461 = ($signed(twiddle_factor_table_41_real) + $signed(twiddle_factor_table_41_imag));
  assign _zz_18462 = ($signed(_zz_1653) - $signed(_zz_18463));
  assign _zz_18463 = ($signed(_zz_18464) * $signed(twiddle_factor_table_41_imag));
  assign _zz_18464 = ($signed(data_mid_42_real) + $signed(data_mid_42_imag));
  assign _zz_18465 = fixTo_1980_dout;
  assign _zz_18466 = ($signed(_zz_1653) + $signed(_zz_18467));
  assign _zz_18467 = ($signed(_zz_18468) * $signed(twiddle_factor_table_41_real));
  assign _zz_18468 = ($signed(data_mid_42_imag) - $signed(data_mid_42_real));
  assign _zz_18469 = fixTo_1981_dout;
  assign _zz_18470 = _zz_18471[31 : 0];
  assign _zz_18471 = _zz_18472;
  assign _zz_18472 = ($signed(_zz_18473) >>> _zz_1654);
  assign _zz_18473 = _zz_18474;
  assign _zz_18474 = ($signed(_zz_18476) - $signed(_zz_1651));
  assign _zz_18475 = ({8'd0,data_mid_10_real} <<< 8);
  assign _zz_18476 = {{8{_zz_18475[23]}}, _zz_18475};
  assign _zz_18477 = fixTo_1982_dout;
  assign _zz_18478 = _zz_18479[31 : 0];
  assign _zz_18479 = _zz_18480;
  assign _zz_18480 = ($signed(_zz_18481) >>> _zz_1654);
  assign _zz_18481 = _zz_18482;
  assign _zz_18482 = ($signed(_zz_18484) - $signed(_zz_1652));
  assign _zz_18483 = ({8'd0,data_mid_10_imag} <<< 8);
  assign _zz_18484 = {{8{_zz_18483[23]}}, _zz_18483};
  assign _zz_18485 = fixTo_1983_dout;
  assign _zz_18486 = _zz_18487[31 : 0];
  assign _zz_18487 = _zz_18488;
  assign _zz_18488 = ($signed(_zz_18489) >>> _zz_1655);
  assign _zz_18489 = _zz_18490;
  assign _zz_18490 = ($signed(_zz_18492) + $signed(_zz_1651));
  assign _zz_18491 = ({8'd0,data_mid_10_real} <<< 8);
  assign _zz_18492 = {{8{_zz_18491[23]}}, _zz_18491};
  assign _zz_18493 = fixTo_1984_dout;
  assign _zz_18494 = _zz_18495[31 : 0];
  assign _zz_18495 = _zz_18496;
  assign _zz_18496 = ($signed(_zz_18497) >>> _zz_1655);
  assign _zz_18497 = _zz_18498;
  assign _zz_18498 = ($signed(_zz_18500) + $signed(_zz_1652));
  assign _zz_18499 = ({8'd0,data_mid_10_imag} <<< 8);
  assign _zz_18500 = {{8{_zz_18499[23]}}, _zz_18499};
  assign _zz_18501 = fixTo_1985_dout;
  assign _zz_18502 = ($signed(twiddle_factor_table_42_real) + $signed(twiddle_factor_table_42_imag));
  assign _zz_18503 = ($signed(_zz_1658) - $signed(_zz_18504));
  assign _zz_18504 = ($signed(_zz_18505) * $signed(twiddle_factor_table_42_imag));
  assign _zz_18505 = ($signed(data_mid_43_real) + $signed(data_mid_43_imag));
  assign _zz_18506 = fixTo_1986_dout;
  assign _zz_18507 = ($signed(_zz_1658) + $signed(_zz_18508));
  assign _zz_18508 = ($signed(_zz_18509) * $signed(twiddle_factor_table_42_real));
  assign _zz_18509 = ($signed(data_mid_43_imag) - $signed(data_mid_43_real));
  assign _zz_18510 = fixTo_1987_dout;
  assign _zz_18511 = _zz_18512[31 : 0];
  assign _zz_18512 = _zz_18513;
  assign _zz_18513 = ($signed(_zz_18514) >>> _zz_1659);
  assign _zz_18514 = _zz_18515;
  assign _zz_18515 = ($signed(_zz_18517) - $signed(_zz_1656));
  assign _zz_18516 = ({8'd0,data_mid_11_real} <<< 8);
  assign _zz_18517 = {{8{_zz_18516[23]}}, _zz_18516};
  assign _zz_18518 = fixTo_1988_dout;
  assign _zz_18519 = _zz_18520[31 : 0];
  assign _zz_18520 = _zz_18521;
  assign _zz_18521 = ($signed(_zz_18522) >>> _zz_1659);
  assign _zz_18522 = _zz_18523;
  assign _zz_18523 = ($signed(_zz_18525) - $signed(_zz_1657));
  assign _zz_18524 = ({8'd0,data_mid_11_imag} <<< 8);
  assign _zz_18525 = {{8{_zz_18524[23]}}, _zz_18524};
  assign _zz_18526 = fixTo_1989_dout;
  assign _zz_18527 = _zz_18528[31 : 0];
  assign _zz_18528 = _zz_18529;
  assign _zz_18529 = ($signed(_zz_18530) >>> _zz_1660);
  assign _zz_18530 = _zz_18531;
  assign _zz_18531 = ($signed(_zz_18533) + $signed(_zz_1656));
  assign _zz_18532 = ({8'd0,data_mid_11_real} <<< 8);
  assign _zz_18533 = {{8{_zz_18532[23]}}, _zz_18532};
  assign _zz_18534 = fixTo_1990_dout;
  assign _zz_18535 = _zz_18536[31 : 0];
  assign _zz_18536 = _zz_18537;
  assign _zz_18537 = ($signed(_zz_18538) >>> _zz_1660);
  assign _zz_18538 = _zz_18539;
  assign _zz_18539 = ($signed(_zz_18541) + $signed(_zz_1657));
  assign _zz_18540 = ({8'd0,data_mid_11_imag} <<< 8);
  assign _zz_18541 = {{8{_zz_18540[23]}}, _zz_18540};
  assign _zz_18542 = fixTo_1991_dout;
  assign _zz_18543 = ($signed(twiddle_factor_table_43_real) + $signed(twiddle_factor_table_43_imag));
  assign _zz_18544 = ($signed(_zz_1663) - $signed(_zz_18545));
  assign _zz_18545 = ($signed(_zz_18546) * $signed(twiddle_factor_table_43_imag));
  assign _zz_18546 = ($signed(data_mid_44_real) + $signed(data_mid_44_imag));
  assign _zz_18547 = fixTo_1992_dout;
  assign _zz_18548 = ($signed(_zz_1663) + $signed(_zz_18549));
  assign _zz_18549 = ($signed(_zz_18550) * $signed(twiddle_factor_table_43_real));
  assign _zz_18550 = ($signed(data_mid_44_imag) - $signed(data_mid_44_real));
  assign _zz_18551 = fixTo_1993_dout;
  assign _zz_18552 = _zz_18553[31 : 0];
  assign _zz_18553 = _zz_18554;
  assign _zz_18554 = ($signed(_zz_18555) >>> _zz_1664);
  assign _zz_18555 = _zz_18556;
  assign _zz_18556 = ($signed(_zz_18558) - $signed(_zz_1661));
  assign _zz_18557 = ({8'd0,data_mid_12_real} <<< 8);
  assign _zz_18558 = {{8{_zz_18557[23]}}, _zz_18557};
  assign _zz_18559 = fixTo_1994_dout;
  assign _zz_18560 = _zz_18561[31 : 0];
  assign _zz_18561 = _zz_18562;
  assign _zz_18562 = ($signed(_zz_18563) >>> _zz_1664);
  assign _zz_18563 = _zz_18564;
  assign _zz_18564 = ($signed(_zz_18566) - $signed(_zz_1662));
  assign _zz_18565 = ({8'd0,data_mid_12_imag} <<< 8);
  assign _zz_18566 = {{8{_zz_18565[23]}}, _zz_18565};
  assign _zz_18567 = fixTo_1995_dout;
  assign _zz_18568 = _zz_18569[31 : 0];
  assign _zz_18569 = _zz_18570;
  assign _zz_18570 = ($signed(_zz_18571) >>> _zz_1665);
  assign _zz_18571 = _zz_18572;
  assign _zz_18572 = ($signed(_zz_18574) + $signed(_zz_1661));
  assign _zz_18573 = ({8'd0,data_mid_12_real} <<< 8);
  assign _zz_18574 = {{8{_zz_18573[23]}}, _zz_18573};
  assign _zz_18575 = fixTo_1996_dout;
  assign _zz_18576 = _zz_18577[31 : 0];
  assign _zz_18577 = _zz_18578;
  assign _zz_18578 = ($signed(_zz_18579) >>> _zz_1665);
  assign _zz_18579 = _zz_18580;
  assign _zz_18580 = ($signed(_zz_18582) + $signed(_zz_1662));
  assign _zz_18581 = ({8'd0,data_mid_12_imag} <<< 8);
  assign _zz_18582 = {{8{_zz_18581[23]}}, _zz_18581};
  assign _zz_18583 = fixTo_1997_dout;
  assign _zz_18584 = ($signed(twiddle_factor_table_44_real) + $signed(twiddle_factor_table_44_imag));
  assign _zz_18585 = ($signed(_zz_1668) - $signed(_zz_18586));
  assign _zz_18586 = ($signed(_zz_18587) * $signed(twiddle_factor_table_44_imag));
  assign _zz_18587 = ($signed(data_mid_45_real) + $signed(data_mid_45_imag));
  assign _zz_18588 = fixTo_1998_dout;
  assign _zz_18589 = ($signed(_zz_1668) + $signed(_zz_18590));
  assign _zz_18590 = ($signed(_zz_18591) * $signed(twiddle_factor_table_44_real));
  assign _zz_18591 = ($signed(data_mid_45_imag) - $signed(data_mid_45_real));
  assign _zz_18592 = fixTo_1999_dout;
  assign _zz_18593 = _zz_18594[31 : 0];
  assign _zz_18594 = _zz_18595;
  assign _zz_18595 = ($signed(_zz_18596) >>> _zz_1669);
  assign _zz_18596 = _zz_18597;
  assign _zz_18597 = ($signed(_zz_18599) - $signed(_zz_1666));
  assign _zz_18598 = ({8'd0,data_mid_13_real} <<< 8);
  assign _zz_18599 = {{8{_zz_18598[23]}}, _zz_18598};
  assign _zz_18600 = fixTo_2000_dout;
  assign _zz_18601 = _zz_18602[31 : 0];
  assign _zz_18602 = _zz_18603;
  assign _zz_18603 = ($signed(_zz_18604) >>> _zz_1669);
  assign _zz_18604 = _zz_18605;
  assign _zz_18605 = ($signed(_zz_18607) - $signed(_zz_1667));
  assign _zz_18606 = ({8'd0,data_mid_13_imag} <<< 8);
  assign _zz_18607 = {{8{_zz_18606[23]}}, _zz_18606};
  assign _zz_18608 = fixTo_2001_dout;
  assign _zz_18609 = _zz_18610[31 : 0];
  assign _zz_18610 = _zz_18611;
  assign _zz_18611 = ($signed(_zz_18612) >>> _zz_1670);
  assign _zz_18612 = _zz_18613;
  assign _zz_18613 = ($signed(_zz_18615) + $signed(_zz_1666));
  assign _zz_18614 = ({8'd0,data_mid_13_real} <<< 8);
  assign _zz_18615 = {{8{_zz_18614[23]}}, _zz_18614};
  assign _zz_18616 = fixTo_2002_dout;
  assign _zz_18617 = _zz_18618[31 : 0];
  assign _zz_18618 = _zz_18619;
  assign _zz_18619 = ($signed(_zz_18620) >>> _zz_1670);
  assign _zz_18620 = _zz_18621;
  assign _zz_18621 = ($signed(_zz_18623) + $signed(_zz_1667));
  assign _zz_18622 = ({8'd0,data_mid_13_imag} <<< 8);
  assign _zz_18623 = {{8{_zz_18622[23]}}, _zz_18622};
  assign _zz_18624 = fixTo_2003_dout;
  assign _zz_18625 = ($signed(twiddle_factor_table_45_real) + $signed(twiddle_factor_table_45_imag));
  assign _zz_18626 = ($signed(_zz_1673) - $signed(_zz_18627));
  assign _zz_18627 = ($signed(_zz_18628) * $signed(twiddle_factor_table_45_imag));
  assign _zz_18628 = ($signed(data_mid_46_real) + $signed(data_mid_46_imag));
  assign _zz_18629 = fixTo_2004_dout;
  assign _zz_18630 = ($signed(_zz_1673) + $signed(_zz_18631));
  assign _zz_18631 = ($signed(_zz_18632) * $signed(twiddle_factor_table_45_real));
  assign _zz_18632 = ($signed(data_mid_46_imag) - $signed(data_mid_46_real));
  assign _zz_18633 = fixTo_2005_dout;
  assign _zz_18634 = _zz_18635[31 : 0];
  assign _zz_18635 = _zz_18636;
  assign _zz_18636 = ($signed(_zz_18637) >>> _zz_1674);
  assign _zz_18637 = _zz_18638;
  assign _zz_18638 = ($signed(_zz_18640) - $signed(_zz_1671));
  assign _zz_18639 = ({8'd0,data_mid_14_real} <<< 8);
  assign _zz_18640 = {{8{_zz_18639[23]}}, _zz_18639};
  assign _zz_18641 = fixTo_2006_dout;
  assign _zz_18642 = _zz_18643[31 : 0];
  assign _zz_18643 = _zz_18644;
  assign _zz_18644 = ($signed(_zz_18645) >>> _zz_1674);
  assign _zz_18645 = _zz_18646;
  assign _zz_18646 = ($signed(_zz_18648) - $signed(_zz_1672));
  assign _zz_18647 = ({8'd0,data_mid_14_imag} <<< 8);
  assign _zz_18648 = {{8{_zz_18647[23]}}, _zz_18647};
  assign _zz_18649 = fixTo_2007_dout;
  assign _zz_18650 = _zz_18651[31 : 0];
  assign _zz_18651 = _zz_18652;
  assign _zz_18652 = ($signed(_zz_18653) >>> _zz_1675);
  assign _zz_18653 = _zz_18654;
  assign _zz_18654 = ($signed(_zz_18656) + $signed(_zz_1671));
  assign _zz_18655 = ({8'd0,data_mid_14_real} <<< 8);
  assign _zz_18656 = {{8{_zz_18655[23]}}, _zz_18655};
  assign _zz_18657 = fixTo_2008_dout;
  assign _zz_18658 = _zz_18659[31 : 0];
  assign _zz_18659 = _zz_18660;
  assign _zz_18660 = ($signed(_zz_18661) >>> _zz_1675);
  assign _zz_18661 = _zz_18662;
  assign _zz_18662 = ($signed(_zz_18664) + $signed(_zz_1672));
  assign _zz_18663 = ({8'd0,data_mid_14_imag} <<< 8);
  assign _zz_18664 = {{8{_zz_18663[23]}}, _zz_18663};
  assign _zz_18665 = fixTo_2009_dout;
  assign _zz_18666 = ($signed(twiddle_factor_table_46_real) + $signed(twiddle_factor_table_46_imag));
  assign _zz_18667 = ($signed(_zz_1678) - $signed(_zz_18668));
  assign _zz_18668 = ($signed(_zz_18669) * $signed(twiddle_factor_table_46_imag));
  assign _zz_18669 = ($signed(data_mid_47_real) + $signed(data_mid_47_imag));
  assign _zz_18670 = fixTo_2010_dout;
  assign _zz_18671 = ($signed(_zz_1678) + $signed(_zz_18672));
  assign _zz_18672 = ($signed(_zz_18673) * $signed(twiddle_factor_table_46_real));
  assign _zz_18673 = ($signed(data_mid_47_imag) - $signed(data_mid_47_real));
  assign _zz_18674 = fixTo_2011_dout;
  assign _zz_18675 = _zz_18676[31 : 0];
  assign _zz_18676 = _zz_18677;
  assign _zz_18677 = ($signed(_zz_18678) >>> _zz_1679);
  assign _zz_18678 = _zz_18679;
  assign _zz_18679 = ($signed(_zz_18681) - $signed(_zz_1676));
  assign _zz_18680 = ({8'd0,data_mid_15_real} <<< 8);
  assign _zz_18681 = {{8{_zz_18680[23]}}, _zz_18680};
  assign _zz_18682 = fixTo_2012_dout;
  assign _zz_18683 = _zz_18684[31 : 0];
  assign _zz_18684 = _zz_18685;
  assign _zz_18685 = ($signed(_zz_18686) >>> _zz_1679);
  assign _zz_18686 = _zz_18687;
  assign _zz_18687 = ($signed(_zz_18689) - $signed(_zz_1677));
  assign _zz_18688 = ({8'd0,data_mid_15_imag} <<< 8);
  assign _zz_18689 = {{8{_zz_18688[23]}}, _zz_18688};
  assign _zz_18690 = fixTo_2013_dout;
  assign _zz_18691 = _zz_18692[31 : 0];
  assign _zz_18692 = _zz_18693;
  assign _zz_18693 = ($signed(_zz_18694) >>> _zz_1680);
  assign _zz_18694 = _zz_18695;
  assign _zz_18695 = ($signed(_zz_18697) + $signed(_zz_1676));
  assign _zz_18696 = ({8'd0,data_mid_15_real} <<< 8);
  assign _zz_18697 = {{8{_zz_18696[23]}}, _zz_18696};
  assign _zz_18698 = fixTo_2014_dout;
  assign _zz_18699 = _zz_18700[31 : 0];
  assign _zz_18700 = _zz_18701;
  assign _zz_18701 = ($signed(_zz_18702) >>> _zz_1680);
  assign _zz_18702 = _zz_18703;
  assign _zz_18703 = ($signed(_zz_18705) + $signed(_zz_1677));
  assign _zz_18704 = ({8'd0,data_mid_15_imag} <<< 8);
  assign _zz_18705 = {{8{_zz_18704[23]}}, _zz_18704};
  assign _zz_18706 = fixTo_2015_dout;
  assign _zz_18707 = ($signed(twiddle_factor_table_47_real) + $signed(twiddle_factor_table_47_imag));
  assign _zz_18708 = ($signed(_zz_1683) - $signed(_zz_18709));
  assign _zz_18709 = ($signed(_zz_18710) * $signed(twiddle_factor_table_47_imag));
  assign _zz_18710 = ($signed(data_mid_48_real) + $signed(data_mid_48_imag));
  assign _zz_18711 = fixTo_2016_dout;
  assign _zz_18712 = ($signed(_zz_1683) + $signed(_zz_18713));
  assign _zz_18713 = ($signed(_zz_18714) * $signed(twiddle_factor_table_47_real));
  assign _zz_18714 = ($signed(data_mid_48_imag) - $signed(data_mid_48_real));
  assign _zz_18715 = fixTo_2017_dout;
  assign _zz_18716 = _zz_18717[31 : 0];
  assign _zz_18717 = _zz_18718;
  assign _zz_18718 = ($signed(_zz_18719) >>> _zz_1684);
  assign _zz_18719 = _zz_18720;
  assign _zz_18720 = ($signed(_zz_18722) - $signed(_zz_1681));
  assign _zz_18721 = ({8'd0,data_mid_16_real} <<< 8);
  assign _zz_18722 = {{8{_zz_18721[23]}}, _zz_18721};
  assign _zz_18723 = fixTo_2018_dout;
  assign _zz_18724 = _zz_18725[31 : 0];
  assign _zz_18725 = _zz_18726;
  assign _zz_18726 = ($signed(_zz_18727) >>> _zz_1684);
  assign _zz_18727 = _zz_18728;
  assign _zz_18728 = ($signed(_zz_18730) - $signed(_zz_1682));
  assign _zz_18729 = ({8'd0,data_mid_16_imag} <<< 8);
  assign _zz_18730 = {{8{_zz_18729[23]}}, _zz_18729};
  assign _zz_18731 = fixTo_2019_dout;
  assign _zz_18732 = _zz_18733[31 : 0];
  assign _zz_18733 = _zz_18734;
  assign _zz_18734 = ($signed(_zz_18735) >>> _zz_1685);
  assign _zz_18735 = _zz_18736;
  assign _zz_18736 = ($signed(_zz_18738) + $signed(_zz_1681));
  assign _zz_18737 = ({8'd0,data_mid_16_real} <<< 8);
  assign _zz_18738 = {{8{_zz_18737[23]}}, _zz_18737};
  assign _zz_18739 = fixTo_2020_dout;
  assign _zz_18740 = _zz_18741[31 : 0];
  assign _zz_18741 = _zz_18742;
  assign _zz_18742 = ($signed(_zz_18743) >>> _zz_1685);
  assign _zz_18743 = _zz_18744;
  assign _zz_18744 = ($signed(_zz_18746) + $signed(_zz_1682));
  assign _zz_18745 = ({8'd0,data_mid_16_imag} <<< 8);
  assign _zz_18746 = {{8{_zz_18745[23]}}, _zz_18745};
  assign _zz_18747 = fixTo_2021_dout;
  assign _zz_18748 = ($signed(twiddle_factor_table_48_real) + $signed(twiddle_factor_table_48_imag));
  assign _zz_18749 = ($signed(_zz_1688) - $signed(_zz_18750));
  assign _zz_18750 = ($signed(_zz_18751) * $signed(twiddle_factor_table_48_imag));
  assign _zz_18751 = ($signed(data_mid_49_real) + $signed(data_mid_49_imag));
  assign _zz_18752 = fixTo_2022_dout;
  assign _zz_18753 = ($signed(_zz_1688) + $signed(_zz_18754));
  assign _zz_18754 = ($signed(_zz_18755) * $signed(twiddle_factor_table_48_real));
  assign _zz_18755 = ($signed(data_mid_49_imag) - $signed(data_mid_49_real));
  assign _zz_18756 = fixTo_2023_dout;
  assign _zz_18757 = _zz_18758[31 : 0];
  assign _zz_18758 = _zz_18759;
  assign _zz_18759 = ($signed(_zz_18760) >>> _zz_1689);
  assign _zz_18760 = _zz_18761;
  assign _zz_18761 = ($signed(_zz_18763) - $signed(_zz_1686));
  assign _zz_18762 = ({8'd0,data_mid_17_real} <<< 8);
  assign _zz_18763 = {{8{_zz_18762[23]}}, _zz_18762};
  assign _zz_18764 = fixTo_2024_dout;
  assign _zz_18765 = _zz_18766[31 : 0];
  assign _zz_18766 = _zz_18767;
  assign _zz_18767 = ($signed(_zz_18768) >>> _zz_1689);
  assign _zz_18768 = _zz_18769;
  assign _zz_18769 = ($signed(_zz_18771) - $signed(_zz_1687));
  assign _zz_18770 = ({8'd0,data_mid_17_imag} <<< 8);
  assign _zz_18771 = {{8{_zz_18770[23]}}, _zz_18770};
  assign _zz_18772 = fixTo_2025_dout;
  assign _zz_18773 = _zz_18774[31 : 0];
  assign _zz_18774 = _zz_18775;
  assign _zz_18775 = ($signed(_zz_18776) >>> _zz_1690);
  assign _zz_18776 = _zz_18777;
  assign _zz_18777 = ($signed(_zz_18779) + $signed(_zz_1686));
  assign _zz_18778 = ({8'd0,data_mid_17_real} <<< 8);
  assign _zz_18779 = {{8{_zz_18778[23]}}, _zz_18778};
  assign _zz_18780 = fixTo_2026_dout;
  assign _zz_18781 = _zz_18782[31 : 0];
  assign _zz_18782 = _zz_18783;
  assign _zz_18783 = ($signed(_zz_18784) >>> _zz_1690);
  assign _zz_18784 = _zz_18785;
  assign _zz_18785 = ($signed(_zz_18787) + $signed(_zz_1687));
  assign _zz_18786 = ({8'd0,data_mid_17_imag} <<< 8);
  assign _zz_18787 = {{8{_zz_18786[23]}}, _zz_18786};
  assign _zz_18788 = fixTo_2027_dout;
  assign _zz_18789 = ($signed(twiddle_factor_table_49_real) + $signed(twiddle_factor_table_49_imag));
  assign _zz_18790 = ($signed(_zz_1693) - $signed(_zz_18791));
  assign _zz_18791 = ($signed(_zz_18792) * $signed(twiddle_factor_table_49_imag));
  assign _zz_18792 = ($signed(data_mid_50_real) + $signed(data_mid_50_imag));
  assign _zz_18793 = fixTo_2028_dout;
  assign _zz_18794 = ($signed(_zz_1693) + $signed(_zz_18795));
  assign _zz_18795 = ($signed(_zz_18796) * $signed(twiddle_factor_table_49_real));
  assign _zz_18796 = ($signed(data_mid_50_imag) - $signed(data_mid_50_real));
  assign _zz_18797 = fixTo_2029_dout;
  assign _zz_18798 = _zz_18799[31 : 0];
  assign _zz_18799 = _zz_18800;
  assign _zz_18800 = ($signed(_zz_18801) >>> _zz_1694);
  assign _zz_18801 = _zz_18802;
  assign _zz_18802 = ($signed(_zz_18804) - $signed(_zz_1691));
  assign _zz_18803 = ({8'd0,data_mid_18_real} <<< 8);
  assign _zz_18804 = {{8{_zz_18803[23]}}, _zz_18803};
  assign _zz_18805 = fixTo_2030_dout;
  assign _zz_18806 = _zz_18807[31 : 0];
  assign _zz_18807 = _zz_18808;
  assign _zz_18808 = ($signed(_zz_18809) >>> _zz_1694);
  assign _zz_18809 = _zz_18810;
  assign _zz_18810 = ($signed(_zz_18812) - $signed(_zz_1692));
  assign _zz_18811 = ({8'd0,data_mid_18_imag} <<< 8);
  assign _zz_18812 = {{8{_zz_18811[23]}}, _zz_18811};
  assign _zz_18813 = fixTo_2031_dout;
  assign _zz_18814 = _zz_18815[31 : 0];
  assign _zz_18815 = _zz_18816;
  assign _zz_18816 = ($signed(_zz_18817) >>> _zz_1695);
  assign _zz_18817 = _zz_18818;
  assign _zz_18818 = ($signed(_zz_18820) + $signed(_zz_1691));
  assign _zz_18819 = ({8'd0,data_mid_18_real} <<< 8);
  assign _zz_18820 = {{8{_zz_18819[23]}}, _zz_18819};
  assign _zz_18821 = fixTo_2032_dout;
  assign _zz_18822 = _zz_18823[31 : 0];
  assign _zz_18823 = _zz_18824;
  assign _zz_18824 = ($signed(_zz_18825) >>> _zz_1695);
  assign _zz_18825 = _zz_18826;
  assign _zz_18826 = ($signed(_zz_18828) + $signed(_zz_1692));
  assign _zz_18827 = ({8'd0,data_mid_18_imag} <<< 8);
  assign _zz_18828 = {{8{_zz_18827[23]}}, _zz_18827};
  assign _zz_18829 = fixTo_2033_dout;
  assign _zz_18830 = ($signed(twiddle_factor_table_50_real) + $signed(twiddle_factor_table_50_imag));
  assign _zz_18831 = ($signed(_zz_1698) - $signed(_zz_18832));
  assign _zz_18832 = ($signed(_zz_18833) * $signed(twiddle_factor_table_50_imag));
  assign _zz_18833 = ($signed(data_mid_51_real) + $signed(data_mid_51_imag));
  assign _zz_18834 = fixTo_2034_dout;
  assign _zz_18835 = ($signed(_zz_1698) + $signed(_zz_18836));
  assign _zz_18836 = ($signed(_zz_18837) * $signed(twiddle_factor_table_50_real));
  assign _zz_18837 = ($signed(data_mid_51_imag) - $signed(data_mid_51_real));
  assign _zz_18838 = fixTo_2035_dout;
  assign _zz_18839 = _zz_18840[31 : 0];
  assign _zz_18840 = _zz_18841;
  assign _zz_18841 = ($signed(_zz_18842) >>> _zz_1699);
  assign _zz_18842 = _zz_18843;
  assign _zz_18843 = ($signed(_zz_18845) - $signed(_zz_1696));
  assign _zz_18844 = ({8'd0,data_mid_19_real} <<< 8);
  assign _zz_18845 = {{8{_zz_18844[23]}}, _zz_18844};
  assign _zz_18846 = fixTo_2036_dout;
  assign _zz_18847 = _zz_18848[31 : 0];
  assign _zz_18848 = _zz_18849;
  assign _zz_18849 = ($signed(_zz_18850) >>> _zz_1699);
  assign _zz_18850 = _zz_18851;
  assign _zz_18851 = ($signed(_zz_18853) - $signed(_zz_1697));
  assign _zz_18852 = ({8'd0,data_mid_19_imag} <<< 8);
  assign _zz_18853 = {{8{_zz_18852[23]}}, _zz_18852};
  assign _zz_18854 = fixTo_2037_dout;
  assign _zz_18855 = _zz_18856[31 : 0];
  assign _zz_18856 = _zz_18857;
  assign _zz_18857 = ($signed(_zz_18858) >>> _zz_1700);
  assign _zz_18858 = _zz_18859;
  assign _zz_18859 = ($signed(_zz_18861) + $signed(_zz_1696));
  assign _zz_18860 = ({8'd0,data_mid_19_real} <<< 8);
  assign _zz_18861 = {{8{_zz_18860[23]}}, _zz_18860};
  assign _zz_18862 = fixTo_2038_dout;
  assign _zz_18863 = _zz_18864[31 : 0];
  assign _zz_18864 = _zz_18865;
  assign _zz_18865 = ($signed(_zz_18866) >>> _zz_1700);
  assign _zz_18866 = _zz_18867;
  assign _zz_18867 = ($signed(_zz_18869) + $signed(_zz_1697));
  assign _zz_18868 = ({8'd0,data_mid_19_imag} <<< 8);
  assign _zz_18869 = {{8{_zz_18868[23]}}, _zz_18868};
  assign _zz_18870 = fixTo_2039_dout;
  assign _zz_18871 = ($signed(twiddle_factor_table_51_real) + $signed(twiddle_factor_table_51_imag));
  assign _zz_18872 = ($signed(_zz_1703) - $signed(_zz_18873));
  assign _zz_18873 = ($signed(_zz_18874) * $signed(twiddle_factor_table_51_imag));
  assign _zz_18874 = ($signed(data_mid_52_real) + $signed(data_mid_52_imag));
  assign _zz_18875 = fixTo_2040_dout;
  assign _zz_18876 = ($signed(_zz_1703) + $signed(_zz_18877));
  assign _zz_18877 = ($signed(_zz_18878) * $signed(twiddle_factor_table_51_real));
  assign _zz_18878 = ($signed(data_mid_52_imag) - $signed(data_mid_52_real));
  assign _zz_18879 = fixTo_2041_dout;
  assign _zz_18880 = _zz_18881[31 : 0];
  assign _zz_18881 = _zz_18882;
  assign _zz_18882 = ($signed(_zz_18883) >>> _zz_1704);
  assign _zz_18883 = _zz_18884;
  assign _zz_18884 = ($signed(_zz_18886) - $signed(_zz_1701));
  assign _zz_18885 = ({8'd0,data_mid_20_real} <<< 8);
  assign _zz_18886 = {{8{_zz_18885[23]}}, _zz_18885};
  assign _zz_18887 = fixTo_2042_dout;
  assign _zz_18888 = _zz_18889[31 : 0];
  assign _zz_18889 = _zz_18890;
  assign _zz_18890 = ($signed(_zz_18891) >>> _zz_1704);
  assign _zz_18891 = _zz_18892;
  assign _zz_18892 = ($signed(_zz_18894) - $signed(_zz_1702));
  assign _zz_18893 = ({8'd0,data_mid_20_imag} <<< 8);
  assign _zz_18894 = {{8{_zz_18893[23]}}, _zz_18893};
  assign _zz_18895 = fixTo_2043_dout;
  assign _zz_18896 = _zz_18897[31 : 0];
  assign _zz_18897 = _zz_18898;
  assign _zz_18898 = ($signed(_zz_18899) >>> _zz_1705);
  assign _zz_18899 = _zz_18900;
  assign _zz_18900 = ($signed(_zz_18902) + $signed(_zz_1701));
  assign _zz_18901 = ({8'd0,data_mid_20_real} <<< 8);
  assign _zz_18902 = {{8{_zz_18901[23]}}, _zz_18901};
  assign _zz_18903 = fixTo_2044_dout;
  assign _zz_18904 = _zz_18905[31 : 0];
  assign _zz_18905 = _zz_18906;
  assign _zz_18906 = ($signed(_zz_18907) >>> _zz_1705);
  assign _zz_18907 = _zz_18908;
  assign _zz_18908 = ($signed(_zz_18910) + $signed(_zz_1702));
  assign _zz_18909 = ({8'd0,data_mid_20_imag} <<< 8);
  assign _zz_18910 = {{8{_zz_18909[23]}}, _zz_18909};
  assign _zz_18911 = fixTo_2045_dout;
  assign _zz_18912 = ($signed(twiddle_factor_table_52_real) + $signed(twiddle_factor_table_52_imag));
  assign _zz_18913 = ($signed(_zz_1708) - $signed(_zz_18914));
  assign _zz_18914 = ($signed(_zz_18915) * $signed(twiddle_factor_table_52_imag));
  assign _zz_18915 = ($signed(data_mid_53_real) + $signed(data_mid_53_imag));
  assign _zz_18916 = fixTo_2046_dout;
  assign _zz_18917 = ($signed(_zz_1708) + $signed(_zz_18918));
  assign _zz_18918 = ($signed(_zz_18919) * $signed(twiddle_factor_table_52_real));
  assign _zz_18919 = ($signed(data_mid_53_imag) - $signed(data_mid_53_real));
  assign _zz_18920 = fixTo_2047_dout;
  assign _zz_18921 = _zz_18922[31 : 0];
  assign _zz_18922 = _zz_18923;
  assign _zz_18923 = ($signed(_zz_18924) >>> _zz_1709);
  assign _zz_18924 = _zz_18925;
  assign _zz_18925 = ($signed(_zz_18927) - $signed(_zz_1706));
  assign _zz_18926 = ({8'd0,data_mid_21_real} <<< 8);
  assign _zz_18927 = {{8{_zz_18926[23]}}, _zz_18926};
  assign _zz_18928 = fixTo_2048_dout;
  assign _zz_18929 = _zz_18930[31 : 0];
  assign _zz_18930 = _zz_18931;
  assign _zz_18931 = ($signed(_zz_18932) >>> _zz_1709);
  assign _zz_18932 = _zz_18933;
  assign _zz_18933 = ($signed(_zz_18935) - $signed(_zz_1707));
  assign _zz_18934 = ({8'd0,data_mid_21_imag} <<< 8);
  assign _zz_18935 = {{8{_zz_18934[23]}}, _zz_18934};
  assign _zz_18936 = fixTo_2049_dout;
  assign _zz_18937 = _zz_18938[31 : 0];
  assign _zz_18938 = _zz_18939;
  assign _zz_18939 = ($signed(_zz_18940) >>> _zz_1710);
  assign _zz_18940 = _zz_18941;
  assign _zz_18941 = ($signed(_zz_18943) + $signed(_zz_1706));
  assign _zz_18942 = ({8'd0,data_mid_21_real} <<< 8);
  assign _zz_18943 = {{8{_zz_18942[23]}}, _zz_18942};
  assign _zz_18944 = fixTo_2050_dout;
  assign _zz_18945 = _zz_18946[31 : 0];
  assign _zz_18946 = _zz_18947;
  assign _zz_18947 = ($signed(_zz_18948) >>> _zz_1710);
  assign _zz_18948 = _zz_18949;
  assign _zz_18949 = ($signed(_zz_18951) + $signed(_zz_1707));
  assign _zz_18950 = ({8'd0,data_mid_21_imag} <<< 8);
  assign _zz_18951 = {{8{_zz_18950[23]}}, _zz_18950};
  assign _zz_18952 = fixTo_2051_dout;
  assign _zz_18953 = ($signed(twiddle_factor_table_53_real) + $signed(twiddle_factor_table_53_imag));
  assign _zz_18954 = ($signed(_zz_1713) - $signed(_zz_18955));
  assign _zz_18955 = ($signed(_zz_18956) * $signed(twiddle_factor_table_53_imag));
  assign _zz_18956 = ($signed(data_mid_54_real) + $signed(data_mid_54_imag));
  assign _zz_18957 = fixTo_2052_dout;
  assign _zz_18958 = ($signed(_zz_1713) + $signed(_zz_18959));
  assign _zz_18959 = ($signed(_zz_18960) * $signed(twiddle_factor_table_53_real));
  assign _zz_18960 = ($signed(data_mid_54_imag) - $signed(data_mid_54_real));
  assign _zz_18961 = fixTo_2053_dout;
  assign _zz_18962 = _zz_18963[31 : 0];
  assign _zz_18963 = _zz_18964;
  assign _zz_18964 = ($signed(_zz_18965) >>> _zz_1714);
  assign _zz_18965 = _zz_18966;
  assign _zz_18966 = ($signed(_zz_18968) - $signed(_zz_1711));
  assign _zz_18967 = ({8'd0,data_mid_22_real} <<< 8);
  assign _zz_18968 = {{8{_zz_18967[23]}}, _zz_18967};
  assign _zz_18969 = fixTo_2054_dout;
  assign _zz_18970 = _zz_18971[31 : 0];
  assign _zz_18971 = _zz_18972;
  assign _zz_18972 = ($signed(_zz_18973) >>> _zz_1714);
  assign _zz_18973 = _zz_18974;
  assign _zz_18974 = ($signed(_zz_18976) - $signed(_zz_1712));
  assign _zz_18975 = ({8'd0,data_mid_22_imag} <<< 8);
  assign _zz_18976 = {{8{_zz_18975[23]}}, _zz_18975};
  assign _zz_18977 = fixTo_2055_dout;
  assign _zz_18978 = _zz_18979[31 : 0];
  assign _zz_18979 = _zz_18980;
  assign _zz_18980 = ($signed(_zz_18981) >>> _zz_1715);
  assign _zz_18981 = _zz_18982;
  assign _zz_18982 = ($signed(_zz_18984) + $signed(_zz_1711));
  assign _zz_18983 = ({8'd0,data_mid_22_real} <<< 8);
  assign _zz_18984 = {{8{_zz_18983[23]}}, _zz_18983};
  assign _zz_18985 = fixTo_2056_dout;
  assign _zz_18986 = _zz_18987[31 : 0];
  assign _zz_18987 = _zz_18988;
  assign _zz_18988 = ($signed(_zz_18989) >>> _zz_1715);
  assign _zz_18989 = _zz_18990;
  assign _zz_18990 = ($signed(_zz_18992) + $signed(_zz_1712));
  assign _zz_18991 = ({8'd0,data_mid_22_imag} <<< 8);
  assign _zz_18992 = {{8{_zz_18991[23]}}, _zz_18991};
  assign _zz_18993 = fixTo_2057_dout;
  assign _zz_18994 = ($signed(twiddle_factor_table_54_real) + $signed(twiddle_factor_table_54_imag));
  assign _zz_18995 = ($signed(_zz_1718) - $signed(_zz_18996));
  assign _zz_18996 = ($signed(_zz_18997) * $signed(twiddle_factor_table_54_imag));
  assign _zz_18997 = ($signed(data_mid_55_real) + $signed(data_mid_55_imag));
  assign _zz_18998 = fixTo_2058_dout;
  assign _zz_18999 = ($signed(_zz_1718) + $signed(_zz_19000));
  assign _zz_19000 = ($signed(_zz_19001) * $signed(twiddle_factor_table_54_real));
  assign _zz_19001 = ($signed(data_mid_55_imag) - $signed(data_mid_55_real));
  assign _zz_19002 = fixTo_2059_dout;
  assign _zz_19003 = _zz_19004[31 : 0];
  assign _zz_19004 = _zz_19005;
  assign _zz_19005 = ($signed(_zz_19006) >>> _zz_1719);
  assign _zz_19006 = _zz_19007;
  assign _zz_19007 = ($signed(_zz_19009) - $signed(_zz_1716));
  assign _zz_19008 = ({8'd0,data_mid_23_real} <<< 8);
  assign _zz_19009 = {{8{_zz_19008[23]}}, _zz_19008};
  assign _zz_19010 = fixTo_2060_dout;
  assign _zz_19011 = _zz_19012[31 : 0];
  assign _zz_19012 = _zz_19013;
  assign _zz_19013 = ($signed(_zz_19014) >>> _zz_1719);
  assign _zz_19014 = _zz_19015;
  assign _zz_19015 = ($signed(_zz_19017) - $signed(_zz_1717));
  assign _zz_19016 = ({8'd0,data_mid_23_imag} <<< 8);
  assign _zz_19017 = {{8{_zz_19016[23]}}, _zz_19016};
  assign _zz_19018 = fixTo_2061_dout;
  assign _zz_19019 = _zz_19020[31 : 0];
  assign _zz_19020 = _zz_19021;
  assign _zz_19021 = ($signed(_zz_19022) >>> _zz_1720);
  assign _zz_19022 = _zz_19023;
  assign _zz_19023 = ($signed(_zz_19025) + $signed(_zz_1716));
  assign _zz_19024 = ({8'd0,data_mid_23_real} <<< 8);
  assign _zz_19025 = {{8{_zz_19024[23]}}, _zz_19024};
  assign _zz_19026 = fixTo_2062_dout;
  assign _zz_19027 = _zz_19028[31 : 0];
  assign _zz_19028 = _zz_19029;
  assign _zz_19029 = ($signed(_zz_19030) >>> _zz_1720);
  assign _zz_19030 = _zz_19031;
  assign _zz_19031 = ($signed(_zz_19033) + $signed(_zz_1717));
  assign _zz_19032 = ({8'd0,data_mid_23_imag} <<< 8);
  assign _zz_19033 = {{8{_zz_19032[23]}}, _zz_19032};
  assign _zz_19034 = fixTo_2063_dout;
  assign _zz_19035 = ($signed(twiddle_factor_table_55_real) + $signed(twiddle_factor_table_55_imag));
  assign _zz_19036 = ($signed(_zz_1723) - $signed(_zz_19037));
  assign _zz_19037 = ($signed(_zz_19038) * $signed(twiddle_factor_table_55_imag));
  assign _zz_19038 = ($signed(data_mid_56_real) + $signed(data_mid_56_imag));
  assign _zz_19039 = fixTo_2064_dout;
  assign _zz_19040 = ($signed(_zz_1723) + $signed(_zz_19041));
  assign _zz_19041 = ($signed(_zz_19042) * $signed(twiddle_factor_table_55_real));
  assign _zz_19042 = ($signed(data_mid_56_imag) - $signed(data_mid_56_real));
  assign _zz_19043 = fixTo_2065_dout;
  assign _zz_19044 = _zz_19045[31 : 0];
  assign _zz_19045 = _zz_19046;
  assign _zz_19046 = ($signed(_zz_19047) >>> _zz_1724);
  assign _zz_19047 = _zz_19048;
  assign _zz_19048 = ($signed(_zz_19050) - $signed(_zz_1721));
  assign _zz_19049 = ({8'd0,data_mid_24_real} <<< 8);
  assign _zz_19050 = {{8{_zz_19049[23]}}, _zz_19049};
  assign _zz_19051 = fixTo_2066_dout;
  assign _zz_19052 = _zz_19053[31 : 0];
  assign _zz_19053 = _zz_19054;
  assign _zz_19054 = ($signed(_zz_19055) >>> _zz_1724);
  assign _zz_19055 = _zz_19056;
  assign _zz_19056 = ($signed(_zz_19058) - $signed(_zz_1722));
  assign _zz_19057 = ({8'd0,data_mid_24_imag} <<< 8);
  assign _zz_19058 = {{8{_zz_19057[23]}}, _zz_19057};
  assign _zz_19059 = fixTo_2067_dout;
  assign _zz_19060 = _zz_19061[31 : 0];
  assign _zz_19061 = _zz_19062;
  assign _zz_19062 = ($signed(_zz_19063) >>> _zz_1725);
  assign _zz_19063 = _zz_19064;
  assign _zz_19064 = ($signed(_zz_19066) + $signed(_zz_1721));
  assign _zz_19065 = ({8'd0,data_mid_24_real} <<< 8);
  assign _zz_19066 = {{8{_zz_19065[23]}}, _zz_19065};
  assign _zz_19067 = fixTo_2068_dout;
  assign _zz_19068 = _zz_19069[31 : 0];
  assign _zz_19069 = _zz_19070;
  assign _zz_19070 = ($signed(_zz_19071) >>> _zz_1725);
  assign _zz_19071 = _zz_19072;
  assign _zz_19072 = ($signed(_zz_19074) + $signed(_zz_1722));
  assign _zz_19073 = ({8'd0,data_mid_24_imag} <<< 8);
  assign _zz_19074 = {{8{_zz_19073[23]}}, _zz_19073};
  assign _zz_19075 = fixTo_2069_dout;
  assign _zz_19076 = ($signed(twiddle_factor_table_56_real) + $signed(twiddle_factor_table_56_imag));
  assign _zz_19077 = ($signed(_zz_1728) - $signed(_zz_19078));
  assign _zz_19078 = ($signed(_zz_19079) * $signed(twiddle_factor_table_56_imag));
  assign _zz_19079 = ($signed(data_mid_57_real) + $signed(data_mid_57_imag));
  assign _zz_19080 = fixTo_2070_dout;
  assign _zz_19081 = ($signed(_zz_1728) + $signed(_zz_19082));
  assign _zz_19082 = ($signed(_zz_19083) * $signed(twiddle_factor_table_56_real));
  assign _zz_19083 = ($signed(data_mid_57_imag) - $signed(data_mid_57_real));
  assign _zz_19084 = fixTo_2071_dout;
  assign _zz_19085 = _zz_19086[31 : 0];
  assign _zz_19086 = _zz_19087;
  assign _zz_19087 = ($signed(_zz_19088) >>> _zz_1729);
  assign _zz_19088 = _zz_19089;
  assign _zz_19089 = ($signed(_zz_19091) - $signed(_zz_1726));
  assign _zz_19090 = ({8'd0,data_mid_25_real} <<< 8);
  assign _zz_19091 = {{8{_zz_19090[23]}}, _zz_19090};
  assign _zz_19092 = fixTo_2072_dout;
  assign _zz_19093 = _zz_19094[31 : 0];
  assign _zz_19094 = _zz_19095;
  assign _zz_19095 = ($signed(_zz_19096) >>> _zz_1729);
  assign _zz_19096 = _zz_19097;
  assign _zz_19097 = ($signed(_zz_19099) - $signed(_zz_1727));
  assign _zz_19098 = ({8'd0,data_mid_25_imag} <<< 8);
  assign _zz_19099 = {{8{_zz_19098[23]}}, _zz_19098};
  assign _zz_19100 = fixTo_2073_dout;
  assign _zz_19101 = _zz_19102[31 : 0];
  assign _zz_19102 = _zz_19103;
  assign _zz_19103 = ($signed(_zz_19104) >>> _zz_1730);
  assign _zz_19104 = _zz_19105;
  assign _zz_19105 = ($signed(_zz_19107) + $signed(_zz_1726));
  assign _zz_19106 = ({8'd0,data_mid_25_real} <<< 8);
  assign _zz_19107 = {{8{_zz_19106[23]}}, _zz_19106};
  assign _zz_19108 = fixTo_2074_dout;
  assign _zz_19109 = _zz_19110[31 : 0];
  assign _zz_19110 = _zz_19111;
  assign _zz_19111 = ($signed(_zz_19112) >>> _zz_1730);
  assign _zz_19112 = _zz_19113;
  assign _zz_19113 = ($signed(_zz_19115) + $signed(_zz_1727));
  assign _zz_19114 = ({8'd0,data_mid_25_imag} <<< 8);
  assign _zz_19115 = {{8{_zz_19114[23]}}, _zz_19114};
  assign _zz_19116 = fixTo_2075_dout;
  assign _zz_19117 = ($signed(twiddle_factor_table_57_real) + $signed(twiddle_factor_table_57_imag));
  assign _zz_19118 = ($signed(_zz_1733) - $signed(_zz_19119));
  assign _zz_19119 = ($signed(_zz_19120) * $signed(twiddle_factor_table_57_imag));
  assign _zz_19120 = ($signed(data_mid_58_real) + $signed(data_mid_58_imag));
  assign _zz_19121 = fixTo_2076_dout;
  assign _zz_19122 = ($signed(_zz_1733) + $signed(_zz_19123));
  assign _zz_19123 = ($signed(_zz_19124) * $signed(twiddle_factor_table_57_real));
  assign _zz_19124 = ($signed(data_mid_58_imag) - $signed(data_mid_58_real));
  assign _zz_19125 = fixTo_2077_dout;
  assign _zz_19126 = _zz_19127[31 : 0];
  assign _zz_19127 = _zz_19128;
  assign _zz_19128 = ($signed(_zz_19129) >>> _zz_1734);
  assign _zz_19129 = _zz_19130;
  assign _zz_19130 = ($signed(_zz_19132) - $signed(_zz_1731));
  assign _zz_19131 = ({8'd0,data_mid_26_real} <<< 8);
  assign _zz_19132 = {{8{_zz_19131[23]}}, _zz_19131};
  assign _zz_19133 = fixTo_2078_dout;
  assign _zz_19134 = _zz_19135[31 : 0];
  assign _zz_19135 = _zz_19136;
  assign _zz_19136 = ($signed(_zz_19137) >>> _zz_1734);
  assign _zz_19137 = _zz_19138;
  assign _zz_19138 = ($signed(_zz_19140) - $signed(_zz_1732));
  assign _zz_19139 = ({8'd0,data_mid_26_imag} <<< 8);
  assign _zz_19140 = {{8{_zz_19139[23]}}, _zz_19139};
  assign _zz_19141 = fixTo_2079_dout;
  assign _zz_19142 = _zz_19143[31 : 0];
  assign _zz_19143 = _zz_19144;
  assign _zz_19144 = ($signed(_zz_19145) >>> _zz_1735);
  assign _zz_19145 = _zz_19146;
  assign _zz_19146 = ($signed(_zz_19148) + $signed(_zz_1731));
  assign _zz_19147 = ({8'd0,data_mid_26_real} <<< 8);
  assign _zz_19148 = {{8{_zz_19147[23]}}, _zz_19147};
  assign _zz_19149 = fixTo_2080_dout;
  assign _zz_19150 = _zz_19151[31 : 0];
  assign _zz_19151 = _zz_19152;
  assign _zz_19152 = ($signed(_zz_19153) >>> _zz_1735);
  assign _zz_19153 = _zz_19154;
  assign _zz_19154 = ($signed(_zz_19156) + $signed(_zz_1732));
  assign _zz_19155 = ({8'd0,data_mid_26_imag} <<< 8);
  assign _zz_19156 = {{8{_zz_19155[23]}}, _zz_19155};
  assign _zz_19157 = fixTo_2081_dout;
  assign _zz_19158 = ($signed(twiddle_factor_table_58_real) + $signed(twiddle_factor_table_58_imag));
  assign _zz_19159 = ($signed(_zz_1738) - $signed(_zz_19160));
  assign _zz_19160 = ($signed(_zz_19161) * $signed(twiddle_factor_table_58_imag));
  assign _zz_19161 = ($signed(data_mid_59_real) + $signed(data_mid_59_imag));
  assign _zz_19162 = fixTo_2082_dout;
  assign _zz_19163 = ($signed(_zz_1738) + $signed(_zz_19164));
  assign _zz_19164 = ($signed(_zz_19165) * $signed(twiddle_factor_table_58_real));
  assign _zz_19165 = ($signed(data_mid_59_imag) - $signed(data_mid_59_real));
  assign _zz_19166 = fixTo_2083_dout;
  assign _zz_19167 = _zz_19168[31 : 0];
  assign _zz_19168 = _zz_19169;
  assign _zz_19169 = ($signed(_zz_19170) >>> _zz_1739);
  assign _zz_19170 = _zz_19171;
  assign _zz_19171 = ($signed(_zz_19173) - $signed(_zz_1736));
  assign _zz_19172 = ({8'd0,data_mid_27_real} <<< 8);
  assign _zz_19173 = {{8{_zz_19172[23]}}, _zz_19172};
  assign _zz_19174 = fixTo_2084_dout;
  assign _zz_19175 = _zz_19176[31 : 0];
  assign _zz_19176 = _zz_19177;
  assign _zz_19177 = ($signed(_zz_19178) >>> _zz_1739);
  assign _zz_19178 = _zz_19179;
  assign _zz_19179 = ($signed(_zz_19181) - $signed(_zz_1737));
  assign _zz_19180 = ({8'd0,data_mid_27_imag} <<< 8);
  assign _zz_19181 = {{8{_zz_19180[23]}}, _zz_19180};
  assign _zz_19182 = fixTo_2085_dout;
  assign _zz_19183 = _zz_19184[31 : 0];
  assign _zz_19184 = _zz_19185;
  assign _zz_19185 = ($signed(_zz_19186) >>> _zz_1740);
  assign _zz_19186 = _zz_19187;
  assign _zz_19187 = ($signed(_zz_19189) + $signed(_zz_1736));
  assign _zz_19188 = ({8'd0,data_mid_27_real} <<< 8);
  assign _zz_19189 = {{8{_zz_19188[23]}}, _zz_19188};
  assign _zz_19190 = fixTo_2086_dout;
  assign _zz_19191 = _zz_19192[31 : 0];
  assign _zz_19192 = _zz_19193;
  assign _zz_19193 = ($signed(_zz_19194) >>> _zz_1740);
  assign _zz_19194 = _zz_19195;
  assign _zz_19195 = ($signed(_zz_19197) + $signed(_zz_1737));
  assign _zz_19196 = ({8'd0,data_mid_27_imag} <<< 8);
  assign _zz_19197 = {{8{_zz_19196[23]}}, _zz_19196};
  assign _zz_19198 = fixTo_2087_dout;
  assign _zz_19199 = ($signed(twiddle_factor_table_59_real) + $signed(twiddle_factor_table_59_imag));
  assign _zz_19200 = ($signed(_zz_1743) - $signed(_zz_19201));
  assign _zz_19201 = ($signed(_zz_19202) * $signed(twiddle_factor_table_59_imag));
  assign _zz_19202 = ($signed(data_mid_60_real) + $signed(data_mid_60_imag));
  assign _zz_19203 = fixTo_2088_dout;
  assign _zz_19204 = ($signed(_zz_1743) + $signed(_zz_19205));
  assign _zz_19205 = ($signed(_zz_19206) * $signed(twiddle_factor_table_59_real));
  assign _zz_19206 = ($signed(data_mid_60_imag) - $signed(data_mid_60_real));
  assign _zz_19207 = fixTo_2089_dout;
  assign _zz_19208 = _zz_19209[31 : 0];
  assign _zz_19209 = _zz_19210;
  assign _zz_19210 = ($signed(_zz_19211) >>> _zz_1744);
  assign _zz_19211 = _zz_19212;
  assign _zz_19212 = ($signed(_zz_19214) - $signed(_zz_1741));
  assign _zz_19213 = ({8'd0,data_mid_28_real} <<< 8);
  assign _zz_19214 = {{8{_zz_19213[23]}}, _zz_19213};
  assign _zz_19215 = fixTo_2090_dout;
  assign _zz_19216 = _zz_19217[31 : 0];
  assign _zz_19217 = _zz_19218;
  assign _zz_19218 = ($signed(_zz_19219) >>> _zz_1744);
  assign _zz_19219 = _zz_19220;
  assign _zz_19220 = ($signed(_zz_19222) - $signed(_zz_1742));
  assign _zz_19221 = ({8'd0,data_mid_28_imag} <<< 8);
  assign _zz_19222 = {{8{_zz_19221[23]}}, _zz_19221};
  assign _zz_19223 = fixTo_2091_dout;
  assign _zz_19224 = _zz_19225[31 : 0];
  assign _zz_19225 = _zz_19226;
  assign _zz_19226 = ($signed(_zz_19227) >>> _zz_1745);
  assign _zz_19227 = _zz_19228;
  assign _zz_19228 = ($signed(_zz_19230) + $signed(_zz_1741));
  assign _zz_19229 = ({8'd0,data_mid_28_real} <<< 8);
  assign _zz_19230 = {{8{_zz_19229[23]}}, _zz_19229};
  assign _zz_19231 = fixTo_2092_dout;
  assign _zz_19232 = _zz_19233[31 : 0];
  assign _zz_19233 = _zz_19234;
  assign _zz_19234 = ($signed(_zz_19235) >>> _zz_1745);
  assign _zz_19235 = _zz_19236;
  assign _zz_19236 = ($signed(_zz_19238) + $signed(_zz_1742));
  assign _zz_19237 = ({8'd0,data_mid_28_imag} <<< 8);
  assign _zz_19238 = {{8{_zz_19237[23]}}, _zz_19237};
  assign _zz_19239 = fixTo_2093_dout;
  assign _zz_19240 = ($signed(twiddle_factor_table_60_real) + $signed(twiddle_factor_table_60_imag));
  assign _zz_19241 = ($signed(_zz_1748) - $signed(_zz_19242));
  assign _zz_19242 = ($signed(_zz_19243) * $signed(twiddle_factor_table_60_imag));
  assign _zz_19243 = ($signed(data_mid_61_real) + $signed(data_mid_61_imag));
  assign _zz_19244 = fixTo_2094_dout;
  assign _zz_19245 = ($signed(_zz_1748) + $signed(_zz_19246));
  assign _zz_19246 = ($signed(_zz_19247) * $signed(twiddle_factor_table_60_real));
  assign _zz_19247 = ($signed(data_mid_61_imag) - $signed(data_mid_61_real));
  assign _zz_19248 = fixTo_2095_dout;
  assign _zz_19249 = _zz_19250[31 : 0];
  assign _zz_19250 = _zz_19251;
  assign _zz_19251 = ($signed(_zz_19252) >>> _zz_1749);
  assign _zz_19252 = _zz_19253;
  assign _zz_19253 = ($signed(_zz_19255) - $signed(_zz_1746));
  assign _zz_19254 = ({8'd0,data_mid_29_real} <<< 8);
  assign _zz_19255 = {{8{_zz_19254[23]}}, _zz_19254};
  assign _zz_19256 = fixTo_2096_dout;
  assign _zz_19257 = _zz_19258[31 : 0];
  assign _zz_19258 = _zz_19259;
  assign _zz_19259 = ($signed(_zz_19260) >>> _zz_1749);
  assign _zz_19260 = _zz_19261;
  assign _zz_19261 = ($signed(_zz_19263) - $signed(_zz_1747));
  assign _zz_19262 = ({8'd0,data_mid_29_imag} <<< 8);
  assign _zz_19263 = {{8{_zz_19262[23]}}, _zz_19262};
  assign _zz_19264 = fixTo_2097_dout;
  assign _zz_19265 = _zz_19266[31 : 0];
  assign _zz_19266 = _zz_19267;
  assign _zz_19267 = ($signed(_zz_19268) >>> _zz_1750);
  assign _zz_19268 = _zz_19269;
  assign _zz_19269 = ($signed(_zz_19271) + $signed(_zz_1746));
  assign _zz_19270 = ({8'd0,data_mid_29_real} <<< 8);
  assign _zz_19271 = {{8{_zz_19270[23]}}, _zz_19270};
  assign _zz_19272 = fixTo_2098_dout;
  assign _zz_19273 = _zz_19274[31 : 0];
  assign _zz_19274 = _zz_19275;
  assign _zz_19275 = ($signed(_zz_19276) >>> _zz_1750);
  assign _zz_19276 = _zz_19277;
  assign _zz_19277 = ($signed(_zz_19279) + $signed(_zz_1747));
  assign _zz_19278 = ({8'd0,data_mid_29_imag} <<< 8);
  assign _zz_19279 = {{8{_zz_19278[23]}}, _zz_19278};
  assign _zz_19280 = fixTo_2099_dout;
  assign _zz_19281 = ($signed(twiddle_factor_table_61_real) + $signed(twiddle_factor_table_61_imag));
  assign _zz_19282 = ($signed(_zz_1753) - $signed(_zz_19283));
  assign _zz_19283 = ($signed(_zz_19284) * $signed(twiddle_factor_table_61_imag));
  assign _zz_19284 = ($signed(data_mid_62_real) + $signed(data_mid_62_imag));
  assign _zz_19285 = fixTo_2100_dout;
  assign _zz_19286 = ($signed(_zz_1753) + $signed(_zz_19287));
  assign _zz_19287 = ($signed(_zz_19288) * $signed(twiddle_factor_table_61_real));
  assign _zz_19288 = ($signed(data_mid_62_imag) - $signed(data_mid_62_real));
  assign _zz_19289 = fixTo_2101_dout;
  assign _zz_19290 = _zz_19291[31 : 0];
  assign _zz_19291 = _zz_19292;
  assign _zz_19292 = ($signed(_zz_19293) >>> _zz_1754);
  assign _zz_19293 = _zz_19294;
  assign _zz_19294 = ($signed(_zz_19296) - $signed(_zz_1751));
  assign _zz_19295 = ({8'd0,data_mid_30_real} <<< 8);
  assign _zz_19296 = {{8{_zz_19295[23]}}, _zz_19295};
  assign _zz_19297 = fixTo_2102_dout;
  assign _zz_19298 = _zz_19299[31 : 0];
  assign _zz_19299 = _zz_19300;
  assign _zz_19300 = ($signed(_zz_19301) >>> _zz_1754);
  assign _zz_19301 = _zz_19302;
  assign _zz_19302 = ($signed(_zz_19304) - $signed(_zz_1752));
  assign _zz_19303 = ({8'd0,data_mid_30_imag} <<< 8);
  assign _zz_19304 = {{8{_zz_19303[23]}}, _zz_19303};
  assign _zz_19305 = fixTo_2103_dout;
  assign _zz_19306 = _zz_19307[31 : 0];
  assign _zz_19307 = _zz_19308;
  assign _zz_19308 = ($signed(_zz_19309) >>> _zz_1755);
  assign _zz_19309 = _zz_19310;
  assign _zz_19310 = ($signed(_zz_19312) + $signed(_zz_1751));
  assign _zz_19311 = ({8'd0,data_mid_30_real} <<< 8);
  assign _zz_19312 = {{8{_zz_19311[23]}}, _zz_19311};
  assign _zz_19313 = fixTo_2104_dout;
  assign _zz_19314 = _zz_19315[31 : 0];
  assign _zz_19315 = _zz_19316;
  assign _zz_19316 = ($signed(_zz_19317) >>> _zz_1755);
  assign _zz_19317 = _zz_19318;
  assign _zz_19318 = ($signed(_zz_19320) + $signed(_zz_1752));
  assign _zz_19319 = ({8'd0,data_mid_30_imag} <<< 8);
  assign _zz_19320 = {{8{_zz_19319[23]}}, _zz_19319};
  assign _zz_19321 = fixTo_2105_dout;
  assign _zz_19322 = ($signed(twiddle_factor_table_62_real) + $signed(twiddle_factor_table_62_imag));
  assign _zz_19323 = ($signed(_zz_1758) - $signed(_zz_19324));
  assign _zz_19324 = ($signed(_zz_19325) * $signed(twiddle_factor_table_62_imag));
  assign _zz_19325 = ($signed(data_mid_63_real) + $signed(data_mid_63_imag));
  assign _zz_19326 = fixTo_2106_dout;
  assign _zz_19327 = ($signed(_zz_1758) + $signed(_zz_19328));
  assign _zz_19328 = ($signed(_zz_19329) * $signed(twiddle_factor_table_62_real));
  assign _zz_19329 = ($signed(data_mid_63_imag) - $signed(data_mid_63_real));
  assign _zz_19330 = fixTo_2107_dout;
  assign _zz_19331 = _zz_19332[31 : 0];
  assign _zz_19332 = _zz_19333;
  assign _zz_19333 = ($signed(_zz_19334) >>> _zz_1759);
  assign _zz_19334 = _zz_19335;
  assign _zz_19335 = ($signed(_zz_19337) - $signed(_zz_1756));
  assign _zz_19336 = ({8'd0,data_mid_31_real} <<< 8);
  assign _zz_19337 = {{8{_zz_19336[23]}}, _zz_19336};
  assign _zz_19338 = fixTo_2108_dout;
  assign _zz_19339 = _zz_19340[31 : 0];
  assign _zz_19340 = _zz_19341;
  assign _zz_19341 = ($signed(_zz_19342) >>> _zz_1759);
  assign _zz_19342 = _zz_19343;
  assign _zz_19343 = ($signed(_zz_19345) - $signed(_zz_1757));
  assign _zz_19344 = ({8'd0,data_mid_31_imag} <<< 8);
  assign _zz_19345 = {{8{_zz_19344[23]}}, _zz_19344};
  assign _zz_19346 = fixTo_2109_dout;
  assign _zz_19347 = _zz_19348[31 : 0];
  assign _zz_19348 = _zz_19349;
  assign _zz_19349 = ($signed(_zz_19350) >>> _zz_1760);
  assign _zz_19350 = _zz_19351;
  assign _zz_19351 = ($signed(_zz_19353) + $signed(_zz_1756));
  assign _zz_19352 = ({8'd0,data_mid_31_real} <<< 8);
  assign _zz_19353 = {{8{_zz_19352[23]}}, _zz_19352};
  assign _zz_19354 = fixTo_2110_dout;
  assign _zz_19355 = _zz_19356[31 : 0];
  assign _zz_19356 = _zz_19357;
  assign _zz_19357 = ($signed(_zz_19358) >>> _zz_1760);
  assign _zz_19358 = _zz_19359;
  assign _zz_19359 = ($signed(_zz_19361) + $signed(_zz_1757));
  assign _zz_19360 = ({8'd0,data_mid_31_imag} <<< 8);
  assign _zz_19361 = {{8{_zz_19360[23]}}, _zz_19360};
  assign _zz_19362 = fixTo_2111_dout;
  assign _zz_19363 = ($signed(twiddle_factor_table_31_real) + $signed(twiddle_factor_table_31_imag));
  assign _zz_19364 = ($signed(_zz_1763) - $signed(_zz_19365));
  assign _zz_19365 = ($signed(_zz_19366) * $signed(twiddle_factor_table_31_imag));
  assign _zz_19366 = ($signed(data_mid_96_real) + $signed(data_mid_96_imag));
  assign _zz_19367 = fixTo_2112_dout;
  assign _zz_19368 = ($signed(_zz_1763) + $signed(_zz_19369));
  assign _zz_19369 = ($signed(_zz_19370) * $signed(twiddle_factor_table_31_real));
  assign _zz_19370 = ($signed(data_mid_96_imag) - $signed(data_mid_96_real));
  assign _zz_19371 = fixTo_2113_dout;
  assign _zz_19372 = _zz_19373[31 : 0];
  assign _zz_19373 = _zz_19374;
  assign _zz_19374 = ($signed(_zz_19375) >>> _zz_1764);
  assign _zz_19375 = _zz_19376;
  assign _zz_19376 = ($signed(_zz_19378) - $signed(_zz_1761));
  assign _zz_19377 = ({8'd0,data_mid_64_real} <<< 8);
  assign _zz_19378 = {{8{_zz_19377[23]}}, _zz_19377};
  assign _zz_19379 = fixTo_2114_dout;
  assign _zz_19380 = _zz_19381[31 : 0];
  assign _zz_19381 = _zz_19382;
  assign _zz_19382 = ($signed(_zz_19383) >>> _zz_1764);
  assign _zz_19383 = _zz_19384;
  assign _zz_19384 = ($signed(_zz_19386) - $signed(_zz_1762));
  assign _zz_19385 = ({8'd0,data_mid_64_imag} <<< 8);
  assign _zz_19386 = {{8{_zz_19385[23]}}, _zz_19385};
  assign _zz_19387 = fixTo_2115_dout;
  assign _zz_19388 = _zz_19389[31 : 0];
  assign _zz_19389 = _zz_19390;
  assign _zz_19390 = ($signed(_zz_19391) >>> _zz_1765);
  assign _zz_19391 = _zz_19392;
  assign _zz_19392 = ($signed(_zz_19394) + $signed(_zz_1761));
  assign _zz_19393 = ({8'd0,data_mid_64_real} <<< 8);
  assign _zz_19394 = {{8{_zz_19393[23]}}, _zz_19393};
  assign _zz_19395 = fixTo_2116_dout;
  assign _zz_19396 = _zz_19397[31 : 0];
  assign _zz_19397 = _zz_19398;
  assign _zz_19398 = ($signed(_zz_19399) >>> _zz_1765);
  assign _zz_19399 = _zz_19400;
  assign _zz_19400 = ($signed(_zz_19402) + $signed(_zz_1762));
  assign _zz_19401 = ({8'd0,data_mid_64_imag} <<< 8);
  assign _zz_19402 = {{8{_zz_19401[23]}}, _zz_19401};
  assign _zz_19403 = fixTo_2117_dout;
  assign _zz_19404 = ($signed(twiddle_factor_table_32_real) + $signed(twiddle_factor_table_32_imag));
  assign _zz_19405 = ($signed(_zz_1768) - $signed(_zz_19406));
  assign _zz_19406 = ($signed(_zz_19407) * $signed(twiddle_factor_table_32_imag));
  assign _zz_19407 = ($signed(data_mid_97_real) + $signed(data_mid_97_imag));
  assign _zz_19408 = fixTo_2118_dout;
  assign _zz_19409 = ($signed(_zz_1768) + $signed(_zz_19410));
  assign _zz_19410 = ($signed(_zz_19411) * $signed(twiddle_factor_table_32_real));
  assign _zz_19411 = ($signed(data_mid_97_imag) - $signed(data_mid_97_real));
  assign _zz_19412 = fixTo_2119_dout;
  assign _zz_19413 = _zz_19414[31 : 0];
  assign _zz_19414 = _zz_19415;
  assign _zz_19415 = ($signed(_zz_19416) >>> _zz_1769);
  assign _zz_19416 = _zz_19417;
  assign _zz_19417 = ($signed(_zz_19419) - $signed(_zz_1766));
  assign _zz_19418 = ({8'd0,data_mid_65_real} <<< 8);
  assign _zz_19419 = {{8{_zz_19418[23]}}, _zz_19418};
  assign _zz_19420 = fixTo_2120_dout;
  assign _zz_19421 = _zz_19422[31 : 0];
  assign _zz_19422 = _zz_19423;
  assign _zz_19423 = ($signed(_zz_19424) >>> _zz_1769);
  assign _zz_19424 = _zz_19425;
  assign _zz_19425 = ($signed(_zz_19427) - $signed(_zz_1767));
  assign _zz_19426 = ({8'd0,data_mid_65_imag} <<< 8);
  assign _zz_19427 = {{8{_zz_19426[23]}}, _zz_19426};
  assign _zz_19428 = fixTo_2121_dout;
  assign _zz_19429 = _zz_19430[31 : 0];
  assign _zz_19430 = _zz_19431;
  assign _zz_19431 = ($signed(_zz_19432) >>> _zz_1770);
  assign _zz_19432 = _zz_19433;
  assign _zz_19433 = ($signed(_zz_19435) + $signed(_zz_1766));
  assign _zz_19434 = ({8'd0,data_mid_65_real} <<< 8);
  assign _zz_19435 = {{8{_zz_19434[23]}}, _zz_19434};
  assign _zz_19436 = fixTo_2122_dout;
  assign _zz_19437 = _zz_19438[31 : 0];
  assign _zz_19438 = _zz_19439;
  assign _zz_19439 = ($signed(_zz_19440) >>> _zz_1770);
  assign _zz_19440 = _zz_19441;
  assign _zz_19441 = ($signed(_zz_19443) + $signed(_zz_1767));
  assign _zz_19442 = ({8'd0,data_mid_65_imag} <<< 8);
  assign _zz_19443 = {{8{_zz_19442[23]}}, _zz_19442};
  assign _zz_19444 = fixTo_2123_dout;
  assign _zz_19445 = ($signed(twiddle_factor_table_33_real) + $signed(twiddle_factor_table_33_imag));
  assign _zz_19446 = ($signed(_zz_1773) - $signed(_zz_19447));
  assign _zz_19447 = ($signed(_zz_19448) * $signed(twiddle_factor_table_33_imag));
  assign _zz_19448 = ($signed(data_mid_98_real) + $signed(data_mid_98_imag));
  assign _zz_19449 = fixTo_2124_dout;
  assign _zz_19450 = ($signed(_zz_1773) + $signed(_zz_19451));
  assign _zz_19451 = ($signed(_zz_19452) * $signed(twiddle_factor_table_33_real));
  assign _zz_19452 = ($signed(data_mid_98_imag) - $signed(data_mid_98_real));
  assign _zz_19453 = fixTo_2125_dout;
  assign _zz_19454 = _zz_19455[31 : 0];
  assign _zz_19455 = _zz_19456;
  assign _zz_19456 = ($signed(_zz_19457) >>> _zz_1774);
  assign _zz_19457 = _zz_19458;
  assign _zz_19458 = ($signed(_zz_19460) - $signed(_zz_1771));
  assign _zz_19459 = ({8'd0,data_mid_66_real} <<< 8);
  assign _zz_19460 = {{8{_zz_19459[23]}}, _zz_19459};
  assign _zz_19461 = fixTo_2126_dout;
  assign _zz_19462 = _zz_19463[31 : 0];
  assign _zz_19463 = _zz_19464;
  assign _zz_19464 = ($signed(_zz_19465) >>> _zz_1774);
  assign _zz_19465 = _zz_19466;
  assign _zz_19466 = ($signed(_zz_19468) - $signed(_zz_1772));
  assign _zz_19467 = ({8'd0,data_mid_66_imag} <<< 8);
  assign _zz_19468 = {{8{_zz_19467[23]}}, _zz_19467};
  assign _zz_19469 = fixTo_2127_dout;
  assign _zz_19470 = _zz_19471[31 : 0];
  assign _zz_19471 = _zz_19472;
  assign _zz_19472 = ($signed(_zz_19473) >>> _zz_1775);
  assign _zz_19473 = _zz_19474;
  assign _zz_19474 = ($signed(_zz_19476) + $signed(_zz_1771));
  assign _zz_19475 = ({8'd0,data_mid_66_real} <<< 8);
  assign _zz_19476 = {{8{_zz_19475[23]}}, _zz_19475};
  assign _zz_19477 = fixTo_2128_dout;
  assign _zz_19478 = _zz_19479[31 : 0];
  assign _zz_19479 = _zz_19480;
  assign _zz_19480 = ($signed(_zz_19481) >>> _zz_1775);
  assign _zz_19481 = _zz_19482;
  assign _zz_19482 = ($signed(_zz_19484) + $signed(_zz_1772));
  assign _zz_19483 = ({8'd0,data_mid_66_imag} <<< 8);
  assign _zz_19484 = {{8{_zz_19483[23]}}, _zz_19483};
  assign _zz_19485 = fixTo_2129_dout;
  assign _zz_19486 = ($signed(twiddle_factor_table_34_real) + $signed(twiddle_factor_table_34_imag));
  assign _zz_19487 = ($signed(_zz_1778) - $signed(_zz_19488));
  assign _zz_19488 = ($signed(_zz_19489) * $signed(twiddle_factor_table_34_imag));
  assign _zz_19489 = ($signed(data_mid_99_real) + $signed(data_mid_99_imag));
  assign _zz_19490 = fixTo_2130_dout;
  assign _zz_19491 = ($signed(_zz_1778) + $signed(_zz_19492));
  assign _zz_19492 = ($signed(_zz_19493) * $signed(twiddle_factor_table_34_real));
  assign _zz_19493 = ($signed(data_mid_99_imag) - $signed(data_mid_99_real));
  assign _zz_19494 = fixTo_2131_dout;
  assign _zz_19495 = _zz_19496[31 : 0];
  assign _zz_19496 = _zz_19497;
  assign _zz_19497 = ($signed(_zz_19498) >>> _zz_1779);
  assign _zz_19498 = _zz_19499;
  assign _zz_19499 = ($signed(_zz_19501) - $signed(_zz_1776));
  assign _zz_19500 = ({8'd0,data_mid_67_real} <<< 8);
  assign _zz_19501 = {{8{_zz_19500[23]}}, _zz_19500};
  assign _zz_19502 = fixTo_2132_dout;
  assign _zz_19503 = _zz_19504[31 : 0];
  assign _zz_19504 = _zz_19505;
  assign _zz_19505 = ($signed(_zz_19506) >>> _zz_1779);
  assign _zz_19506 = _zz_19507;
  assign _zz_19507 = ($signed(_zz_19509) - $signed(_zz_1777));
  assign _zz_19508 = ({8'd0,data_mid_67_imag} <<< 8);
  assign _zz_19509 = {{8{_zz_19508[23]}}, _zz_19508};
  assign _zz_19510 = fixTo_2133_dout;
  assign _zz_19511 = _zz_19512[31 : 0];
  assign _zz_19512 = _zz_19513;
  assign _zz_19513 = ($signed(_zz_19514) >>> _zz_1780);
  assign _zz_19514 = _zz_19515;
  assign _zz_19515 = ($signed(_zz_19517) + $signed(_zz_1776));
  assign _zz_19516 = ({8'd0,data_mid_67_real} <<< 8);
  assign _zz_19517 = {{8{_zz_19516[23]}}, _zz_19516};
  assign _zz_19518 = fixTo_2134_dout;
  assign _zz_19519 = _zz_19520[31 : 0];
  assign _zz_19520 = _zz_19521;
  assign _zz_19521 = ($signed(_zz_19522) >>> _zz_1780);
  assign _zz_19522 = _zz_19523;
  assign _zz_19523 = ($signed(_zz_19525) + $signed(_zz_1777));
  assign _zz_19524 = ({8'd0,data_mid_67_imag} <<< 8);
  assign _zz_19525 = {{8{_zz_19524[23]}}, _zz_19524};
  assign _zz_19526 = fixTo_2135_dout;
  assign _zz_19527 = ($signed(twiddle_factor_table_35_real) + $signed(twiddle_factor_table_35_imag));
  assign _zz_19528 = ($signed(_zz_1783) - $signed(_zz_19529));
  assign _zz_19529 = ($signed(_zz_19530) * $signed(twiddle_factor_table_35_imag));
  assign _zz_19530 = ($signed(data_mid_100_real) + $signed(data_mid_100_imag));
  assign _zz_19531 = fixTo_2136_dout;
  assign _zz_19532 = ($signed(_zz_1783) + $signed(_zz_19533));
  assign _zz_19533 = ($signed(_zz_19534) * $signed(twiddle_factor_table_35_real));
  assign _zz_19534 = ($signed(data_mid_100_imag) - $signed(data_mid_100_real));
  assign _zz_19535 = fixTo_2137_dout;
  assign _zz_19536 = _zz_19537[31 : 0];
  assign _zz_19537 = _zz_19538;
  assign _zz_19538 = ($signed(_zz_19539) >>> _zz_1784);
  assign _zz_19539 = _zz_19540;
  assign _zz_19540 = ($signed(_zz_19542) - $signed(_zz_1781));
  assign _zz_19541 = ({8'd0,data_mid_68_real} <<< 8);
  assign _zz_19542 = {{8{_zz_19541[23]}}, _zz_19541};
  assign _zz_19543 = fixTo_2138_dout;
  assign _zz_19544 = _zz_19545[31 : 0];
  assign _zz_19545 = _zz_19546;
  assign _zz_19546 = ($signed(_zz_19547) >>> _zz_1784);
  assign _zz_19547 = _zz_19548;
  assign _zz_19548 = ($signed(_zz_19550) - $signed(_zz_1782));
  assign _zz_19549 = ({8'd0,data_mid_68_imag} <<< 8);
  assign _zz_19550 = {{8{_zz_19549[23]}}, _zz_19549};
  assign _zz_19551 = fixTo_2139_dout;
  assign _zz_19552 = _zz_19553[31 : 0];
  assign _zz_19553 = _zz_19554;
  assign _zz_19554 = ($signed(_zz_19555) >>> _zz_1785);
  assign _zz_19555 = _zz_19556;
  assign _zz_19556 = ($signed(_zz_19558) + $signed(_zz_1781));
  assign _zz_19557 = ({8'd0,data_mid_68_real} <<< 8);
  assign _zz_19558 = {{8{_zz_19557[23]}}, _zz_19557};
  assign _zz_19559 = fixTo_2140_dout;
  assign _zz_19560 = _zz_19561[31 : 0];
  assign _zz_19561 = _zz_19562;
  assign _zz_19562 = ($signed(_zz_19563) >>> _zz_1785);
  assign _zz_19563 = _zz_19564;
  assign _zz_19564 = ($signed(_zz_19566) + $signed(_zz_1782));
  assign _zz_19565 = ({8'd0,data_mid_68_imag} <<< 8);
  assign _zz_19566 = {{8{_zz_19565[23]}}, _zz_19565};
  assign _zz_19567 = fixTo_2141_dout;
  assign _zz_19568 = ($signed(twiddle_factor_table_36_real) + $signed(twiddle_factor_table_36_imag));
  assign _zz_19569 = ($signed(_zz_1788) - $signed(_zz_19570));
  assign _zz_19570 = ($signed(_zz_19571) * $signed(twiddle_factor_table_36_imag));
  assign _zz_19571 = ($signed(data_mid_101_real) + $signed(data_mid_101_imag));
  assign _zz_19572 = fixTo_2142_dout;
  assign _zz_19573 = ($signed(_zz_1788) + $signed(_zz_19574));
  assign _zz_19574 = ($signed(_zz_19575) * $signed(twiddle_factor_table_36_real));
  assign _zz_19575 = ($signed(data_mid_101_imag) - $signed(data_mid_101_real));
  assign _zz_19576 = fixTo_2143_dout;
  assign _zz_19577 = _zz_19578[31 : 0];
  assign _zz_19578 = _zz_19579;
  assign _zz_19579 = ($signed(_zz_19580) >>> _zz_1789);
  assign _zz_19580 = _zz_19581;
  assign _zz_19581 = ($signed(_zz_19583) - $signed(_zz_1786));
  assign _zz_19582 = ({8'd0,data_mid_69_real} <<< 8);
  assign _zz_19583 = {{8{_zz_19582[23]}}, _zz_19582};
  assign _zz_19584 = fixTo_2144_dout;
  assign _zz_19585 = _zz_19586[31 : 0];
  assign _zz_19586 = _zz_19587;
  assign _zz_19587 = ($signed(_zz_19588) >>> _zz_1789);
  assign _zz_19588 = _zz_19589;
  assign _zz_19589 = ($signed(_zz_19591) - $signed(_zz_1787));
  assign _zz_19590 = ({8'd0,data_mid_69_imag} <<< 8);
  assign _zz_19591 = {{8{_zz_19590[23]}}, _zz_19590};
  assign _zz_19592 = fixTo_2145_dout;
  assign _zz_19593 = _zz_19594[31 : 0];
  assign _zz_19594 = _zz_19595;
  assign _zz_19595 = ($signed(_zz_19596) >>> _zz_1790);
  assign _zz_19596 = _zz_19597;
  assign _zz_19597 = ($signed(_zz_19599) + $signed(_zz_1786));
  assign _zz_19598 = ({8'd0,data_mid_69_real} <<< 8);
  assign _zz_19599 = {{8{_zz_19598[23]}}, _zz_19598};
  assign _zz_19600 = fixTo_2146_dout;
  assign _zz_19601 = _zz_19602[31 : 0];
  assign _zz_19602 = _zz_19603;
  assign _zz_19603 = ($signed(_zz_19604) >>> _zz_1790);
  assign _zz_19604 = _zz_19605;
  assign _zz_19605 = ($signed(_zz_19607) + $signed(_zz_1787));
  assign _zz_19606 = ({8'd0,data_mid_69_imag} <<< 8);
  assign _zz_19607 = {{8{_zz_19606[23]}}, _zz_19606};
  assign _zz_19608 = fixTo_2147_dout;
  assign _zz_19609 = ($signed(twiddle_factor_table_37_real) + $signed(twiddle_factor_table_37_imag));
  assign _zz_19610 = ($signed(_zz_1793) - $signed(_zz_19611));
  assign _zz_19611 = ($signed(_zz_19612) * $signed(twiddle_factor_table_37_imag));
  assign _zz_19612 = ($signed(data_mid_102_real) + $signed(data_mid_102_imag));
  assign _zz_19613 = fixTo_2148_dout;
  assign _zz_19614 = ($signed(_zz_1793) + $signed(_zz_19615));
  assign _zz_19615 = ($signed(_zz_19616) * $signed(twiddle_factor_table_37_real));
  assign _zz_19616 = ($signed(data_mid_102_imag) - $signed(data_mid_102_real));
  assign _zz_19617 = fixTo_2149_dout;
  assign _zz_19618 = _zz_19619[31 : 0];
  assign _zz_19619 = _zz_19620;
  assign _zz_19620 = ($signed(_zz_19621) >>> _zz_1794);
  assign _zz_19621 = _zz_19622;
  assign _zz_19622 = ($signed(_zz_19624) - $signed(_zz_1791));
  assign _zz_19623 = ({8'd0,data_mid_70_real} <<< 8);
  assign _zz_19624 = {{8{_zz_19623[23]}}, _zz_19623};
  assign _zz_19625 = fixTo_2150_dout;
  assign _zz_19626 = _zz_19627[31 : 0];
  assign _zz_19627 = _zz_19628;
  assign _zz_19628 = ($signed(_zz_19629) >>> _zz_1794);
  assign _zz_19629 = _zz_19630;
  assign _zz_19630 = ($signed(_zz_19632) - $signed(_zz_1792));
  assign _zz_19631 = ({8'd0,data_mid_70_imag} <<< 8);
  assign _zz_19632 = {{8{_zz_19631[23]}}, _zz_19631};
  assign _zz_19633 = fixTo_2151_dout;
  assign _zz_19634 = _zz_19635[31 : 0];
  assign _zz_19635 = _zz_19636;
  assign _zz_19636 = ($signed(_zz_19637) >>> _zz_1795);
  assign _zz_19637 = _zz_19638;
  assign _zz_19638 = ($signed(_zz_19640) + $signed(_zz_1791));
  assign _zz_19639 = ({8'd0,data_mid_70_real} <<< 8);
  assign _zz_19640 = {{8{_zz_19639[23]}}, _zz_19639};
  assign _zz_19641 = fixTo_2152_dout;
  assign _zz_19642 = _zz_19643[31 : 0];
  assign _zz_19643 = _zz_19644;
  assign _zz_19644 = ($signed(_zz_19645) >>> _zz_1795);
  assign _zz_19645 = _zz_19646;
  assign _zz_19646 = ($signed(_zz_19648) + $signed(_zz_1792));
  assign _zz_19647 = ({8'd0,data_mid_70_imag} <<< 8);
  assign _zz_19648 = {{8{_zz_19647[23]}}, _zz_19647};
  assign _zz_19649 = fixTo_2153_dout;
  assign _zz_19650 = ($signed(twiddle_factor_table_38_real) + $signed(twiddle_factor_table_38_imag));
  assign _zz_19651 = ($signed(_zz_1798) - $signed(_zz_19652));
  assign _zz_19652 = ($signed(_zz_19653) * $signed(twiddle_factor_table_38_imag));
  assign _zz_19653 = ($signed(data_mid_103_real) + $signed(data_mid_103_imag));
  assign _zz_19654 = fixTo_2154_dout;
  assign _zz_19655 = ($signed(_zz_1798) + $signed(_zz_19656));
  assign _zz_19656 = ($signed(_zz_19657) * $signed(twiddle_factor_table_38_real));
  assign _zz_19657 = ($signed(data_mid_103_imag) - $signed(data_mid_103_real));
  assign _zz_19658 = fixTo_2155_dout;
  assign _zz_19659 = _zz_19660[31 : 0];
  assign _zz_19660 = _zz_19661;
  assign _zz_19661 = ($signed(_zz_19662) >>> _zz_1799);
  assign _zz_19662 = _zz_19663;
  assign _zz_19663 = ($signed(_zz_19665) - $signed(_zz_1796));
  assign _zz_19664 = ({8'd0,data_mid_71_real} <<< 8);
  assign _zz_19665 = {{8{_zz_19664[23]}}, _zz_19664};
  assign _zz_19666 = fixTo_2156_dout;
  assign _zz_19667 = _zz_19668[31 : 0];
  assign _zz_19668 = _zz_19669;
  assign _zz_19669 = ($signed(_zz_19670) >>> _zz_1799);
  assign _zz_19670 = _zz_19671;
  assign _zz_19671 = ($signed(_zz_19673) - $signed(_zz_1797));
  assign _zz_19672 = ({8'd0,data_mid_71_imag} <<< 8);
  assign _zz_19673 = {{8{_zz_19672[23]}}, _zz_19672};
  assign _zz_19674 = fixTo_2157_dout;
  assign _zz_19675 = _zz_19676[31 : 0];
  assign _zz_19676 = _zz_19677;
  assign _zz_19677 = ($signed(_zz_19678) >>> _zz_1800);
  assign _zz_19678 = _zz_19679;
  assign _zz_19679 = ($signed(_zz_19681) + $signed(_zz_1796));
  assign _zz_19680 = ({8'd0,data_mid_71_real} <<< 8);
  assign _zz_19681 = {{8{_zz_19680[23]}}, _zz_19680};
  assign _zz_19682 = fixTo_2158_dout;
  assign _zz_19683 = _zz_19684[31 : 0];
  assign _zz_19684 = _zz_19685;
  assign _zz_19685 = ($signed(_zz_19686) >>> _zz_1800);
  assign _zz_19686 = _zz_19687;
  assign _zz_19687 = ($signed(_zz_19689) + $signed(_zz_1797));
  assign _zz_19688 = ({8'd0,data_mid_71_imag} <<< 8);
  assign _zz_19689 = {{8{_zz_19688[23]}}, _zz_19688};
  assign _zz_19690 = fixTo_2159_dout;
  assign _zz_19691 = ($signed(twiddle_factor_table_39_real) + $signed(twiddle_factor_table_39_imag));
  assign _zz_19692 = ($signed(_zz_1803) - $signed(_zz_19693));
  assign _zz_19693 = ($signed(_zz_19694) * $signed(twiddle_factor_table_39_imag));
  assign _zz_19694 = ($signed(data_mid_104_real) + $signed(data_mid_104_imag));
  assign _zz_19695 = fixTo_2160_dout;
  assign _zz_19696 = ($signed(_zz_1803) + $signed(_zz_19697));
  assign _zz_19697 = ($signed(_zz_19698) * $signed(twiddle_factor_table_39_real));
  assign _zz_19698 = ($signed(data_mid_104_imag) - $signed(data_mid_104_real));
  assign _zz_19699 = fixTo_2161_dout;
  assign _zz_19700 = _zz_19701[31 : 0];
  assign _zz_19701 = _zz_19702;
  assign _zz_19702 = ($signed(_zz_19703) >>> _zz_1804);
  assign _zz_19703 = _zz_19704;
  assign _zz_19704 = ($signed(_zz_19706) - $signed(_zz_1801));
  assign _zz_19705 = ({8'd0,data_mid_72_real} <<< 8);
  assign _zz_19706 = {{8{_zz_19705[23]}}, _zz_19705};
  assign _zz_19707 = fixTo_2162_dout;
  assign _zz_19708 = _zz_19709[31 : 0];
  assign _zz_19709 = _zz_19710;
  assign _zz_19710 = ($signed(_zz_19711) >>> _zz_1804);
  assign _zz_19711 = _zz_19712;
  assign _zz_19712 = ($signed(_zz_19714) - $signed(_zz_1802));
  assign _zz_19713 = ({8'd0,data_mid_72_imag} <<< 8);
  assign _zz_19714 = {{8{_zz_19713[23]}}, _zz_19713};
  assign _zz_19715 = fixTo_2163_dout;
  assign _zz_19716 = _zz_19717[31 : 0];
  assign _zz_19717 = _zz_19718;
  assign _zz_19718 = ($signed(_zz_19719) >>> _zz_1805);
  assign _zz_19719 = _zz_19720;
  assign _zz_19720 = ($signed(_zz_19722) + $signed(_zz_1801));
  assign _zz_19721 = ({8'd0,data_mid_72_real} <<< 8);
  assign _zz_19722 = {{8{_zz_19721[23]}}, _zz_19721};
  assign _zz_19723 = fixTo_2164_dout;
  assign _zz_19724 = _zz_19725[31 : 0];
  assign _zz_19725 = _zz_19726;
  assign _zz_19726 = ($signed(_zz_19727) >>> _zz_1805);
  assign _zz_19727 = _zz_19728;
  assign _zz_19728 = ($signed(_zz_19730) + $signed(_zz_1802));
  assign _zz_19729 = ({8'd0,data_mid_72_imag} <<< 8);
  assign _zz_19730 = {{8{_zz_19729[23]}}, _zz_19729};
  assign _zz_19731 = fixTo_2165_dout;
  assign _zz_19732 = ($signed(twiddle_factor_table_40_real) + $signed(twiddle_factor_table_40_imag));
  assign _zz_19733 = ($signed(_zz_1808) - $signed(_zz_19734));
  assign _zz_19734 = ($signed(_zz_19735) * $signed(twiddle_factor_table_40_imag));
  assign _zz_19735 = ($signed(data_mid_105_real) + $signed(data_mid_105_imag));
  assign _zz_19736 = fixTo_2166_dout;
  assign _zz_19737 = ($signed(_zz_1808) + $signed(_zz_19738));
  assign _zz_19738 = ($signed(_zz_19739) * $signed(twiddle_factor_table_40_real));
  assign _zz_19739 = ($signed(data_mid_105_imag) - $signed(data_mid_105_real));
  assign _zz_19740 = fixTo_2167_dout;
  assign _zz_19741 = _zz_19742[31 : 0];
  assign _zz_19742 = _zz_19743;
  assign _zz_19743 = ($signed(_zz_19744) >>> _zz_1809);
  assign _zz_19744 = _zz_19745;
  assign _zz_19745 = ($signed(_zz_19747) - $signed(_zz_1806));
  assign _zz_19746 = ({8'd0,data_mid_73_real} <<< 8);
  assign _zz_19747 = {{8{_zz_19746[23]}}, _zz_19746};
  assign _zz_19748 = fixTo_2168_dout;
  assign _zz_19749 = _zz_19750[31 : 0];
  assign _zz_19750 = _zz_19751;
  assign _zz_19751 = ($signed(_zz_19752) >>> _zz_1809);
  assign _zz_19752 = _zz_19753;
  assign _zz_19753 = ($signed(_zz_19755) - $signed(_zz_1807));
  assign _zz_19754 = ({8'd0,data_mid_73_imag} <<< 8);
  assign _zz_19755 = {{8{_zz_19754[23]}}, _zz_19754};
  assign _zz_19756 = fixTo_2169_dout;
  assign _zz_19757 = _zz_19758[31 : 0];
  assign _zz_19758 = _zz_19759;
  assign _zz_19759 = ($signed(_zz_19760) >>> _zz_1810);
  assign _zz_19760 = _zz_19761;
  assign _zz_19761 = ($signed(_zz_19763) + $signed(_zz_1806));
  assign _zz_19762 = ({8'd0,data_mid_73_real} <<< 8);
  assign _zz_19763 = {{8{_zz_19762[23]}}, _zz_19762};
  assign _zz_19764 = fixTo_2170_dout;
  assign _zz_19765 = _zz_19766[31 : 0];
  assign _zz_19766 = _zz_19767;
  assign _zz_19767 = ($signed(_zz_19768) >>> _zz_1810);
  assign _zz_19768 = _zz_19769;
  assign _zz_19769 = ($signed(_zz_19771) + $signed(_zz_1807));
  assign _zz_19770 = ({8'd0,data_mid_73_imag} <<< 8);
  assign _zz_19771 = {{8{_zz_19770[23]}}, _zz_19770};
  assign _zz_19772 = fixTo_2171_dout;
  assign _zz_19773 = ($signed(twiddle_factor_table_41_real) + $signed(twiddle_factor_table_41_imag));
  assign _zz_19774 = ($signed(_zz_1813) - $signed(_zz_19775));
  assign _zz_19775 = ($signed(_zz_19776) * $signed(twiddle_factor_table_41_imag));
  assign _zz_19776 = ($signed(data_mid_106_real) + $signed(data_mid_106_imag));
  assign _zz_19777 = fixTo_2172_dout;
  assign _zz_19778 = ($signed(_zz_1813) + $signed(_zz_19779));
  assign _zz_19779 = ($signed(_zz_19780) * $signed(twiddle_factor_table_41_real));
  assign _zz_19780 = ($signed(data_mid_106_imag) - $signed(data_mid_106_real));
  assign _zz_19781 = fixTo_2173_dout;
  assign _zz_19782 = _zz_19783[31 : 0];
  assign _zz_19783 = _zz_19784;
  assign _zz_19784 = ($signed(_zz_19785) >>> _zz_1814);
  assign _zz_19785 = _zz_19786;
  assign _zz_19786 = ($signed(_zz_19788) - $signed(_zz_1811));
  assign _zz_19787 = ({8'd0,data_mid_74_real} <<< 8);
  assign _zz_19788 = {{8{_zz_19787[23]}}, _zz_19787};
  assign _zz_19789 = fixTo_2174_dout;
  assign _zz_19790 = _zz_19791[31 : 0];
  assign _zz_19791 = _zz_19792;
  assign _zz_19792 = ($signed(_zz_19793) >>> _zz_1814);
  assign _zz_19793 = _zz_19794;
  assign _zz_19794 = ($signed(_zz_19796) - $signed(_zz_1812));
  assign _zz_19795 = ({8'd0,data_mid_74_imag} <<< 8);
  assign _zz_19796 = {{8{_zz_19795[23]}}, _zz_19795};
  assign _zz_19797 = fixTo_2175_dout;
  assign _zz_19798 = _zz_19799[31 : 0];
  assign _zz_19799 = _zz_19800;
  assign _zz_19800 = ($signed(_zz_19801) >>> _zz_1815);
  assign _zz_19801 = _zz_19802;
  assign _zz_19802 = ($signed(_zz_19804) + $signed(_zz_1811));
  assign _zz_19803 = ({8'd0,data_mid_74_real} <<< 8);
  assign _zz_19804 = {{8{_zz_19803[23]}}, _zz_19803};
  assign _zz_19805 = fixTo_2176_dout;
  assign _zz_19806 = _zz_19807[31 : 0];
  assign _zz_19807 = _zz_19808;
  assign _zz_19808 = ($signed(_zz_19809) >>> _zz_1815);
  assign _zz_19809 = _zz_19810;
  assign _zz_19810 = ($signed(_zz_19812) + $signed(_zz_1812));
  assign _zz_19811 = ({8'd0,data_mid_74_imag} <<< 8);
  assign _zz_19812 = {{8{_zz_19811[23]}}, _zz_19811};
  assign _zz_19813 = fixTo_2177_dout;
  assign _zz_19814 = ($signed(twiddle_factor_table_42_real) + $signed(twiddle_factor_table_42_imag));
  assign _zz_19815 = ($signed(_zz_1818) - $signed(_zz_19816));
  assign _zz_19816 = ($signed(_zz_19817) * $signed(twiddle_factor_table_42_imag));
  assign _zz_19817 = ($signed(data_mid_107_real) + $signed(data_mid_107_imag));
  assign _zz_19818 = fixTo_2178_dout;
  assign _zz_19819 = ($signed(_zz_1818) + $signed(_zz_19820));
  assign _zz_19820 = ($signed(_zz_19821) * $signed(twiddle_factor_table_42_real));
  assign _zz_19821 = ($signed(data_mid_107_imag) - $signed(data_mid_107_real));
  assign _zz_19822 = fixTo_2179_dout;
  assign _zz_19823 = _zz_19824[31 : 0];
  assign _zz_19824 = _zz_19825;
  assign _zz_19825 = ($signed(_zz_19826) >>> _zz_1819);
  assign _zz_19826 = _zz_19827;
  assign _zz_19827 = ($signed(_zz_19829) - $signed(_zz_1816));
  assign _zz_19828 = ({8'd0,data_mid_75_real} <<< 8);
  assign _zz_19829 = {{8{_zz_19828[23]}}, _zz_19828};
  assign _zz_19830 = fixTo_2180_dout;
  assign _zz_19831 = _zz_19832[31 : 0];
  assign _zz_19832 = _zz_19833;
  assign _zz_19833 = ($signed(_zz_19834) >>> _zz_1819);
  assign _zz_19834 = _zz_19835;
  assign _zz_19835 = ($signed(_zz_19837) - $signed(_zz_1817));
  assign _zz_19836 = ({8'd0,data_mid_75_imag} <<< 8);
  assign _zz_19837 = {{8{_zz_19836[23]}}, _zz_19836};
  assign _zz_19838 = fixTo_2181_dout;
  assign _zz_19839 = _zz_19840[31 : 0];
  assign _zz_19840 = _zz_19841;
  assign _zz_19841 = ($signed(_zz_19842) >>> _zz_1820);
  assign _zz_19842 = _zz_19843;
  assign _zz_19843 = ($signed(_zz_19845) + $signed(_zz_1816));
  assign _zz_19844 = ({8'd0,data_mid_75_real} <<< 8);
  assign _zz_19845 = {{8{_zz_19844[23]}}, _zz_19844};
  assign _zz_19846 = fixTo_2182_dout;
  assign _zz_19847 = _zz_19848[31 : 0];
  assign _zz_19848 = _zz_19849;
  assign _zz_19849 = ($signed(_zz_19850) >>> _zz_1820);
  assign _zz_19850 = _zz_19851;
  assign _zz_19851 = ($signed(_zz_19853) + $signed(_zz_1817));
  assign _zz_19852 = ({8'd0,data_mid_75_imag} <<< 8);
  assign _zz_19853 = {{8{_zz_19852[23]}}, _zz_19852};
  assign _zz_19854 = fixTo_2183_dout;
  assign _zz_19855 = ($signed(twiddle_factor_table_43_real) + $signed(twiddle_factor_table_43_imag));
  assign _zz_19856 = ($signed(_zz_1823) - $signed(_zz_19857));
  assign _zz_19857 = ($signed(_zz_19858) * $signed(twiddle_factor_table_43_imag));
  assign _zz_19858 = ($signed(data_mid_108_real) + $signed(data_mid_108_imag));
  assign _zz_19859 = fixTo_2184_dout;
  assign _zz_19860 = ($signed(_zz_1823) + $signed(_zz_19861));
  assign _zz_19861 = ($signed(_zz_19862) * $signed(twiddle_factor_table_43_real));
  assign _zz_19862 = ($signed(data_mid_108_imag) - $signed(data_mid_108_real));
  assign _zz_19863 = fixTo_2185_dout;
  assign _zz_19864 = _zz_19865[31 : 0];
  assign _zz_19865 = _zz_19866;
  assign _zz_19866 = ($signed(_zz_19867) >>> _zz_1824);
  assign _zz_19867 = _zz_19868;
  assign _zz_19868 = ($signed(_zz_19870) - $signed(_zz_1821));
  assign _zz_19869 = ({8'd0,data_mid_76_real} <<< 8);
  assign _zz_19870 = {{8{_zz_19869[23]}}, _zz_19869};
  assign _zz_19871 = fixTo_2186_dout;
  assign _zz_19872 = _zz_19873[31 : 0];
  assign _zz_19873 = _zz_19874;
  assign _zz_19874 = ($signed(_zz_19875) >>> _zz_1824);
  assign _zz_19875 = _zz_19876;
  assign _zz_19876 = ($signed(_zz_19878) - $signed(_zz_1822));
  assign _zz_19877 = ({8'd0,data_mid_76_imag} <<< 8);
  assign _zz_19878 = {{8{_zz_19877[23]}}, _zz_19877};
  assign _zz_19879 = fixTo_2187_dout;
  assign _zz_19880 = _zz_19881[31 : 0];
  assign _zz_19881 = _zz_19882;
  assign _zz_19882 = ($signed(_zz_19883) >>> _zz_1825);
  assign _zz_19883 = _zz_19884;
  assign _zz_19884 = ($signed(_zz_19886) + $signed(_zz_1821));
  assign _zz_19885 = ({8'd0,data_mid_76_real} <<< 8);
  assign _zz_19886 = {{8{_zz_19885[23]}}, _zz_19885};
  assign _zz_19887 = fixTo_2188_dout;
  assign _zz_19888 = _zz_19889[31 : 0];
  assign _zz_19889 = _zz_19890;
  assign _zz_19890 = ($signed(_zz_19891) >>> _zz_1825);
  assign _zz_19891 = _zz_19892;
  assign _zz_19892 = ($signed(_zz_19894) + $signed(_zz_1822));
  assign _zz_19893 = ({8'd0,data_mid_76_imag} <<< 8);
  assign _zz_19894 = {{8{_zz_19893[23]}}, _zz_19893};
  assign _zz_19895 = fixTo_2189_dout;
  assign _zz_19896 = ($signed(twiddle_factor_table_44_real) + $signed(twiddle_factor_table_44_imag));
  assign _zz_19897 = ($signed(_zz_1828) - $signed(_zz_19898));
  assign _zz_19898 = ($signed(_zz_19899) * $signed(twiddle_factor_table_44_imag));
  assign _zz_19899 = ($signed(data_mid_109_real) + $signed(data_mid_109_imag));
  assign _zz_19900 = fixTo_2190_dout;
  assign _zz_19901 = ($signed(_zz_1828) + $signed(_zz_19902));
  assign _zz_19902 = ($signed(_zz_19903) * $signed(twiddle_factor_table_44_real));
  assign _zz_19903 = ($signed(data_mid_109_imag) - $signed(data_mid_109_real));
  assign _zz_19904 = fixTo_2191_dout;
  assign _zz_19905 = _zz_19906[31 : 0];
  assign _zz_19906 = _zz_19907;
  assign _zz_19907 = ($signed(_zz_19908) >>> _zz_1829);
  assign _zz_19908 = _zz_19909;
  assign _zz_19909 = ($signed(_zz_19911) - $signed(_zz_1826));
  assign _zz_19910 = ({8'd0,data_mid_77_real} <<< 8);
  assign _zz_19911 = {{8{_zz_19910[23]}}, _zz_19910};
  assign _zz_19912 = fixTo_2192_dout;
  assign _zz_19913 = _zz_19914[31 : 0];
  assign _zz_19914 = _zz_19915;
  assign _zz_19915 = ($signed(_zz_19916) >>> _zz_1829);
  assign _zz_19916 = _zz_19917;
  assign _zz_19917 = ($signed(_zz_19919) - $signed(_zz_1827));
  assign _zz_19918 = ({8'd0,data_mid_77_imag} <<< 8);
  assign _zz_19919 = {{8{_zz_19918[23]}}, _zz_19918};
  assign _zz_19920 = fixTo_2193_dout;
  assign _zz_19921 = _zz_19922[31 : 0];
  assign _zz_19922 = _zz_19923;
  assign _zz_19923 = ($signed(_zz_19924) >>> _zz_1830);
  assign _zz_19924 = _zz_19925;
  assign _zz_19925 = ($signed(_zz_19927) + $signed(_zz_1826));
  assign _zz_19926 = ({8'd0,data_mid_77_real} <<< 8);
  assign _zz_19927 = {{8{_zz_19926[23]}}, _zz_19926};
  assign _zz_19928 = fixTo_2194_dout;
  assign _zz_19929 = _zz_19930[31 : 0];
  assign _zz_19930 = _zz_19931;
  assign _zz_19931 = ($signed(_zz_19932) >>> _zz_1830);
  assign _zz_19932 = _zz_19933;
  assign _zz_19933 = ($signed(_zz_19935) + $signed(_zz_1827));
  assign _zz_19934 = ({8'd0,data_mid_77_imag} <<< 8);
  assign _zz_19935 = {{8{_zz_19934[23]}}, _zz_19934};
  assign _zz_19936 = fixTo_2195_dout;
  assign _zz_19937 = ($signed(twiddle_factor_table_45_real) + $signed(twiddle_factor_table_45_imag));
  assign _zz_19938 = ($signed(_zz_1833) - $signed(_zz_19939));
  assign _zz_19939 = ($signed(_zz_19940) * $signed(twiddle_factor_table_45_imag));
  assign _zz_19940 = ($signed(data_mid_110_real) + $signed(data_mid_110_imag));
  assign _zz_19941 = fixTo_2196_dout;
  assign _zz_19942 = ($signed(_zz_1833) + $signed(_zz_19943));
  assign _zz_19943 = ($signed(_zz_19944) * $signed(twiddle_factor_table_45_real));
  assign _zz_19944 = ($signed(data_mid_110_imag) - $signed(data_mid_110_real));
  assign _zz_19945 = fixTo_2197_dout;
  assign _zz_19946 = _zz_19947[31 : 0];
  assign _zz_19947 = _zz_19948;
  assign _zz_19948 = ($signed(_zz_19949) >>> _zz_1834);
  assign _zz_19949 = _zz_19950;
  assign _zz_19950 = ($signed(_zz_19952) - $signed(_zz_1831));
  assign _zz_19951 = ({8'd0,data_mid_78_real} <<< 8);
  assign _zz_19952 = {{8{_zz_19951[23]}}, _zz_19951};
  assign _zz_19953 = fixTo_2198_dout;
  assign _zz_19954 = _zz_19955[31 : 0];
  assign _zz_19955 = _zz_19956;
  assign _zz_19956 = ($signed(_zz_19957) >>> _zz_1834);
  assign _zz_19957 = _zz_19958;
  assign _zz_19958 = ($signed(_zz_19960) - $signed(_zz_1832));
  assign _zz_19959 = ({8'd0,data_mid_78_imag} <<< 8);
  assign _zz_19960 = {{8{_zz_19959[23]}}, _zz_19959};
  assign _zz_19961 = fixTo_2199_dout;
  assign _zz_19962 = _zz_19963[31 : 0];
  assign _zz_19963 = _zz_19964;
  assign _zz_19964 = ($signed(_zz_19965) >>> _zz_1835);
  assign _zz_19965 = _zz_19966;
  assign _zz_19966 = ($signed(_zz_19968) + $signed(_zz_1831));
  assign _zz_19967 = ({8'd0,data_mid_78_real} <<< 8);
  assign _zz_19968 = {{8{_zz_19967[23]}}, _zz_19967};
  assign _zz_19969 = fixTo_2200_dout;
  assign _zz_19970 = _zz_19971[31 : 0];
  assign _zz_19971 = _zz_19972;
  assign _zz_19972 = ($signed(_zz_19973) >>> _zz_1835);
  assign _zz_19973 = _zz_19974;
  assign _zz_19974 = ($signed(_zz_19976) + $signed(_zz_1832));
  assign _zz_19975 = ({8'd0,data_mid_78_imag} <<< 8);
  assign _zz_19976 = {{8{_zz_19975[23]}}, _zz_19975};
  assign _zz_19977 = fixTo_2201_dout;
  assign _zz_19978 = ($signed(twiddle_factor_table_46_real) + $signed(twiddle_factor_table_46_imag));
  assign _zz_19979 = ($signed(_zz_1838) - $signed(_zz_19980));
  assign _zz_19980 = ($signed(_zz_19981) * $signed(twiddle_factor_table_46_imag));
  assign _zz_19981 = ($signed(data_mid_111_real) + $signed(data_mid_111_imag));
  assign _zz_19982 = fixTo_2202_dout;
  assign _zz_19983 = ($signed(_zz_1838) + $signed(_zz_19984));
  assign _zz_19984 = ($signed(_zz_19985) * $signed(twiddle_factor_table_46_real));
  assign _zz_19985 = ($signed(data_mid_111_imag) - $signed(data_mid_111_real));
  assign _zz_19986 = fixTo_2203_dout;
  assign _zz_19987 = _zz_19988[31 : 0];
  assign _zz_19988 = _zz_19989;
  assign _zz_19989 = ($signed(_zz_19990) >>> _zz_1839);
  assign _zz_19990 = _zz_19991;
  assign _zz_19991 = ($signed(_zz_19993) - $signed(_zz_1836));
  assign _zz_19992 = ({8'd0,data_mid_79_real} <<< 8);
  assign _zz_19993 = {{8{_zz_19992[23]}}, _zz_19992};
  assign _zz_19994 = fixTo_2204_dout;
  assign _zz_19995 = _zz_19996[31 : 0];
  assign _zz_19996 = _zz_19997;
  assign _zz_19997 = ($signed(_zz_19998) >>> _zz_1839);
  assign _zz_19998 = _zz_19999;
  assign _zz_19999 = ($signed(_zz_20001) - $signed(_zz_1837));
  assign _zz_20000 = ({8'd0,data_mid_79_imag} <<< 8);
  assign _zz_20001 = {{8{_zz_20000[23]}}, _zz_20000};
  assign _zz_20002 = fixTo_2205_dout;
  assign _zz_20003 = _zz_20004[31 : 0];
  assign _zz_20004 = _zz_20005;
  assign _zz_20005 = ($signed(_zz_20006) >>> _zz_1840);
  assign _zz_20006 = _zz_20007;
  assign _zz_20007 = ($signed(_zz_20009) + $signed(_zz_1836));
  assign _zz_20008 = ({8'd0,data_mid_79_real} <<< 8);
  assign _zz_20009 = {{8{_zz_20008[23]}}, _zz_20008};
  assign _zz_20010 = fixTo_2206_dout;
  assign _zz_20011 = _zz_20012[31 : 0];
  assign _zz_20012 = _zz_20013;
  assign _zz_20013 = ($signed(_zz_20014) >>> _zz_1840);
  assign _zz_20014 = _zz_20015;
  assign _zz_20015 = ($signed(_zz_20017) + $signed(_zz_1837));
  assign _zz_20016 = ({8'd0,data_mid_79_imag} <<< 8);
  assign _zz_20017 = {{8{_zz_20016[23]}}, _zz_20016};
  assign _zz_20018 = fixTo_2207_dout;
  assign _zz_20019 = ($signed(twiddle_factor_table_47_real) + $signed(twiddle_factor_table_47_imag));
  assign _zz_20020 = ($signed(_zz_1843) - $signed(_zz_20021));
  assign _zz_20021 = ($signed(_zz_20022) * $signed(twiddle_factor_table_47_imag));
  assign _zz_20022 = ($signed(data_mid_112_real) + $signed(data_mid_112_imag));
  assign _zz_20023 = fixTo_2208_dout;
  assign _zz_20024 = ($signed(_zz_1843) + $signed(_zz_20025));
  assign _zz_20025 = ($signed(_zz_20026) * $signed(twiddle_factor_table_47_real));
  assign _zz_20026 = ($signed(data_mid_112_imag) - $signed(data_mid_112_real));
  assign _zz_20027 = fixTo_2209_dout;
  assign _zz_20028 = _zz_20029[31 : 0];
  assign _zz_20029 = _zz_20030;
  assign _zz_20030 = ($signed(_zz_20031) >>> _zz_1844);
  assign _zz_20031 = _zz_20032;
  assign _zz_20032 = ($signed(_zz_20034) - $signed(_zz_1841));
  assign _zz_20033 = ({8'd0,data_mid_80_real} <<< 8);
  assign _zz_20034 = {{8{_zz_20033[23]}}, _zz_20033};
  assign _zz_20035 = fixTo_2210_dout;
  assign _zz_20036 = _zz_20037[31 : 0];
  assign _zz_20037 = _zz_20038;
  assign _zz_20038 = ($signed(_zz_20039) >>> _zz_1844);
  assign _zz_20039 = _zz_20040;
  assign _zz_20040 = ($signed(_zz_20042) - $signed(_zz_1842));
  assign _zz_20041 = ({8'd0,data_mid_80_imag} <<< 8);
  assign _zz_20042 = {{8{_zz_20041[23]}}, _zz_20041};
  assign _zz_20043 = fixTo_2211_dout;
  assign _zz_20044 = _zz_20045[31 : 0];
  assign _zz_20045 = _zz_20046;
  assign _zz_20046 = ($signed(_zz_20047) >>> _zz_1845);
  assign _zz_20047 = _zz_20048;
  assign _zz_20048 = ($signed(_zz_20050) + $signed(_zz_1841));
  assign _zz_20049 = ({8'd0,data_mid_80_real} <<< 8);
  assign _zz_20050 = {{8{_zz_20049[23]}}, _zz_20049};
  assign _zz_20051 = fixTo_2212_dout;
  assign _zz_20052 = _zz_20053[31 : 0];
  assign _zz_20053 = _zz_20054;
  assign _zz_20054 = ($signed(_zz_20055) >>> _zz_1845);
  assign _zz_20055 = _zz_20056;
  assign _zz_20056 = ($signed(_zz_20058) + $signed(_zz_1842));
  assign _zz_20057 = ({8'd0,data_mid_80_imag} <<< 8);
  assign _zz_20058 = {{8{_zz_20057[23]}}, _zz_20057};
  assign _zz_20059 = fixTo_2213_dout;
  assign _zz_20060 = ($signed(twiddle_factor_table_48_real) + $signed(twiddle_factor_table_48_imag));
  assign _zz_20061 = ($signed(_zz_1848) - $signed(_zz_20062));
  assign _zz_20062 = ($signed(_zz_20063) * $signed(twiddle_factor_table_48_imag));
  assign _zz_20063 = ($signed(data_mid_113_real) + $signed(data_mid_113_imag));
  assign _zz_20064 = fixTo_2214_dout;
  assign _zz_20065 = ($signed(_zz_1848) + $signed(_zz_20066));
  assign _zz_20066 = ($signed(_zz_20067) * $signed(twiddle_factor_table_48_real));
  assign _zz_20067 = ($signed(data_mid_113_imag) - $signed(data_mid_113_real));
  assign _zz_20068 = fixTo_2215_dout;
  assign _zz_20069 = _zz_20070[31 : 0];
  assign _zz_20070 = _zz_20071;
  assign _zz_20071 = ($signed(_zz_20072) >>> _zz_1849);
  assign _zz_20072 = _zz_20073;
  assign _zz_20073 = ($signed(_zz_20075) - $signed(_zz_1846));
  assign _zz_20074 = ({8'd0,data_mid_81_real} <<< 8);
  assign _zz_20075 = {{8{_zz_20074[23]}}, _zz_20074};
  assign _zz_20076 = fixTo_2216_dout;
  assign _zz_20077 = _zz_20078[31 : 0];
  assign _zz_20078 = _zz_20079;
  assign _zz_20079 = ($signed(_zz_20080) >>> _zz_1849);
  assign _zz_20080 = _zz_20081;
  assign _zz_20081 = ($signed(_zz_20083) - $signed(_zz_1847));
  assign _zz_20082 = ({8'd0,data_mid_81_imag} <<< 8);
  assign _zz_20083 = {{8{_zz_20082[23]}}, _zz_20082};
  assign _zz_20084 = fixTo_2217_dout;
  assign _zz_20085 = _zz_20086[31 : 0];
  assign _zz_20086 = _zz_20087;
  assign _zz_20087 = ($signed(_zz_20088) >>> _zz_1850);
  assign _zz_20088 = _zz_20089;
  assign _zz_20089 = ($signed(_zz_20091) + $signed(_zz_1846));
  assign _zz_20090 = ({8'd0,data_mid_81_real} <<< 8);
  assign _zz_20091 = {{8{_zz_20090[23]}}, _zz_20090};
  assign _zz_20092 = fixTo_2218_dout;
  assign _zz_20093 = _zz_20094[31 : 0];
  assign _zz_20094 = _zz_20095;
  assign _zz_20095 = ($signed(_zz_20096) >>> _zz_1850);
  assign _zz_20096 = _zz_20097;
  assign _zz_20097 = ($signed(_zz_20099) + $signed(_zz_1847));
  assign _zz_20098 = ({8'd0,data_mid_81_imag} <<< 8);
  assign _zz_20099 = {{8{_zz_20098[23]}}, _zz_20098};
  assign _zz_20100 = fixTo_2219_dout;
  assign _zz_20101 = ($signed(twiddle_factor_table_49_real) + $signed(twiddle_factor_table_49_imag));
  assign _zz_20102 = ($signed(_zz_1853) - $signed(_zz_20103));
  assign _zz_20103 = ($signed(_zz_20104) * $signed(twiddle_factor_table_49_imag));
  assign _zz_20104 = ($signed(data_mid_114_real) + $signed(data_mid_114_imag));
  assign _zz_20105 = fixTo_2220_dout;
  assign _zz_20106 = ($signed(_zz_1853) + $signed(_zz_20107));
  assign _zz_20107 = ($signed(_zz_20108) * $signed(twiddle_factor_table_49_real));
  assign _zz_20108 = ($signed(data_mid_114_imag) - $signed(data_mid_114_real));
  assign _zz_20109 = fixTo_2221_dout;
  assign _zz_20110 = _zz_20111[31 : 0];
  assign _zz_20111 = _zz_20112;
  assign _zz_20112 = ($signed(_zz_20113) >>> _zz_1854);
  assign _zz_20113 = _zz_20114;
  assign _zz_20114 = ($signed(_zz_20116) - $signed(_zz_1851));
  assign _zz_20115 = ({8'd0,data_mid_82_real} <<< 8);
  assign _zz_20116 = {{8{_zz_20115[23]}}, _zz_20115};
  assign _zz_20117 = fixTo_2222_dout;
  assign _zz_20118 = _zz_20119[31 : 0];
  assign _zz_20119 = _zz_20120;
  assign _zz_20120 = ($signed(_zz_20121) >>> _zz_1854);
  assign _zz_20121 = _zz_20122;
  assign _zz_20122 = ($signed(_zz_20124) - $signed(_zz_1852));
  assign _zz_20123 = ({8'd0,data_mid_82_imag} <<< 8);
  assign _zz_20124 = {{8{_zz_20123[23]}}, _zz_20123};
  assign _zz_20125 = fixTo_2223_dout;
  assign _zz_20126 = _zz_20127[31 : 0];
  assign _zz_20127 = _zz_20128;
  assign _zz_20128 = ($signed(_zz_20129) >>> _zz_1855);
  assign _zz_20129 = _zz_20130;
  assign _zz_20130 = ($signed(_zz_20132) + $signed(_zz_1851));
  assign _zz_20131 = ({8'd0,data_mid_82_real} <<< 8);
  assign _zz_20132 = {{8{_zz_20131[23]}}, _zz_20131};
  assign _zz_20133 = fixTo_2224_dout;
  assign _zz_20134 = _zz_20135[31 : 0];
  assign _zz_20135 = _zz_20136;
  assign _zz_20136 = ($signed(_zz_20137) >>> _zz_1855);
  assign _zz_20137 = _zz_20138;
  assign _zz_20138 = ($signed(_zz_20140) + $signed(_zz_1852));
  assign _zz_20139 = ({8'd0,data_mid_82_imag} <<< 8);
  assign _zz_20140 = {{8{_zz_20139[23]}}, _zz_20139};
  assign _zz_20141 = fixTo_2225_dout;
  assign _zz_20142 = ($signed(twiddle_factor_table_50_real) + $signed(twiddle_factor_table_50_imag));
  assign _zz_20143 = ($signed(_zz_1858) - $signed(_zz_20144));
  assign _zz_20144 = ($signed(_zz_20145) * $signed(twiddle_factor_table_50_imag));
  assign _zz_20145 = ($signed(data_mid_115_real) + $signed(data_mid_115_imag));
  assign _zz_20146 = fixTo_2226_dout;
  assign _zz_20147 = ($signed(_zz_1858) + $signed(_zz_20148));
  assign _zz_20148 = ($signed(_zz_20149) * $signed(twiddle_factor_table_50_real));
  assign _zz_20149 = ($signed(data_mid_115_imag) - $signed(data_mid_115_real));
  assign _zz_20150 = fixTo_2227_dout;
  assign _zz_20151 = _zz_20152[31 : 0];
  assign _zz_20152 = _zz_20153;
  assign _zz_20153 = ($signed(_zz_20154) >>> _zz_1859);
  assign _zz_20154 = _zz_20155;
  assign _zz_20155 = ($signed(_zz_20157) - $signed(_zz_1856));
  assign _zz_20156 = ({8'd0,data_mid_83_real} <<< 8);
  assign _zz_20157 = {{8{_zz_20156[23]}}, _zz_20156};
  assign _zz_20158 = fixTo_2228_dout;
  assign _zz_20159 = _zz_20160[31 : 0];
  assign _zz_20160 = _zz_20161;
  assign _zz_20161 = ($signed(_zz_20162) >>> _zz_1859);
  assign _zz_20162 = _zz_20163;
  assign _zz_20163 = ($signed(_zz_20165) - $signed(_zz_1857));
  assign _zz_20164 = ({8'd0,data_mid_83_imag} <<< 8);
  assign _zz_20165 = {{8{_zz_20164[23]}}, _zz_20164};
  assign _zz_20166 = fixTo_2229_dout;
  assign _zz_20167 = _zz_20168[31 : 0];
  assign _zz_20168 = _zz_20169;
  assign _zz_20169 = ($signed(_zz_20170) >>> _zz_1860);
  assign _zz_20170 = _zz_20171;
  assign _zz_20171 = ($signed(_zz_20173) + $signed(_zz_1856));
  assign _zz_20172 = ({8'd0,data_mid_83_real} <<< 8);
  assign _zz_20173 = {{8{_zz_20172[23]}}, _zz_20172};
  assign _zz_20174 = fixTo_2230_dout;
  assign _zz_20175 = _zz_20176[31 : 0];
  assign _zz_20176 = _zz_20177;
  assign _zz_20177 = ($signed(_zz_20178) >>> _zz_1860);
  assign _zz_20178 = _zz_20179;
  assign _zz_20179 = ($signed(_zz_20181) + $signed(_zz_1857));
  assign _zz_20180 = ({8'd0,data_mid_83_imag} <<< 8);
  assign _zz_20181 = {{8{_zz_20180[23]}}, _zz_20180};
  assign _zz_20182 = fixTo_2231_dout;
  assign _zz_20183 = ($signed(twiddle_factor_table_51_real) + $signed(twiddle_factor_table_51_imag));
  assign _zz_20184 = ($signed(_zz_1863) - $signed(_zz_20185));
  assign _zz_20185 = ($signed(_zz_20186) * $signed(twiddle_factor_table_51_imag));
  assign _zz_20186 = ($signed(data_mid_116_real) + $signed(data_mid_116_imag));
  assign _zz_20187 = fixTo_2232_dout;
  assign _zz_20188 = ($signed(_zz_1863) + $signed(_zz_20189));
  assign _zz_20189 = ($signed(_zz_20190) * $signed(twiddle_factor_table_51_real));
  assign _zz_20190 = ($signed(data_mid_116_imag) - $signed(data_mid_116_real));
  assign _zz_20191 = fixTo_2233_dout;
  assign _zz_20192 = _zz_20193[31 : 0];
  assign _zz_20193 = _zz_20194;
  assign _zz_20194 = ($signed(_zz_20195) >>> _zz_1864);
  assign _zz_20195 = _zz_20196;
  assign _zz_20196 = ($signed(_zz_20198) - $signed(_zz_1861));
  assign _zz_20197 = ({8'd0,data_mid_84_real} <<< 8);
  assign _zz_20198 = {{8{_zz_20197[23]}}, _zz_20197};
  assign _zz_20199 = fixTo_2234_dout;
  assign _zz_20200 = _zz_20201[31 : 0];
  assign _zz_20201 = _zz_20202;
  assign _zz_20202 = ($signed(_zz_20203) >>> _zz_1864);
  assign _zz_20203 = _zz_20204;
  assign _zz_20204 = ($signed(_zz_20206) - $signed(_zz_1862));
  assign _zz_20205 = ({8'd0,data_mid_84_imag} <<< 8);
  assign _zz_20206 = {{8{_zz_20205[23]}}, _zz_20205};
  assign _zz_20207 = fixTo_2235_dout;
  assign _zz_20208 = _zz_20209[31 : 0];
  assign _zz_20209 = _zz_20210;
  assign _zz_20210 = ($signed(_zz_20211) >>> _zz_1865);
  assign _zz_20211 = _zz_20212;
  assign _zz_20212 = ($signed(_zz_20214) + $signed(_zz_1861));
  assign _zz_20213 = ({8'd0,data_mid_84_real} <<< 8);
  assign _zz_20214 = {{8{_zz_20213[23]}}, _zz_20213};
  assign _zz_20215 = fixTo_2236_dout;
  assign _zz_20216 = _zz_20217[31 : 0];
  assign _zz_20217 = _zz_20218;
  assign _zz_20218 = ($signed(_zz_20219) >>> _zz_1865);
  assign _zz_20219 = _zz_20220;
  assign _zz_20220 = ($signed(_zz_20222) + $signed(_zz_1862));
  assign _zz_20221 = ({8'd0,data_mid_84_imag} <<< 8);
  assign _zz_20222 = {{8{_zz_20221[23]}}, _zz_20221};
  assign _zz_20223 = fixTo_2237_dout;
  assign _zz_20224 = ($signed(twiddle_factor_table_52_real) + $signed(twiddle_factor_table_52_imag));
  assign _zz_20225 = ($signed(_zz_1868) - $signed(_zz_20226));
  assign _zz_20226 = ($signed(_zz_20227) * $signed(twiddle_factor_table_52_imag));
  assign _zz_20227 = ($signed(data_mid_117_real) + $signed(data_mid_117_imag));
  assign _zz_20228 = fixTo_2238_dout;
  assign _zz_20229 = ($signed(_zz_1868) + $signed(_zz_20230));
  assign _zz_20230 = ($signed(_zz_20231) * $signed(twiddle_factor_table_52_real));
  assign _zz_20231 = ($signed(data_mid_117_imag) - $signed(data_mid_117_real));
  assign _zz_20232 = fixTo_2239_dout;
  assign _zz_20233 = _zz_20234[31 : 0];
  assign _zz_20234 = _zz_20235;
  assign _zz_20235 = ($signed(_zz_20236) >>> _zz_1869);
  assign _zz_20236 = _zz_20237;
  assign _zz_20237 = ($signed(_zz_20239) - $signed(_zz_1866));
  assign _zz_20238 = ({8'd0,data_mid_85_real} <<< 8);
  assign _zz_20239 = {{8{_zz_20238[23]}}, _zz_20238};
  assign _zz_20240 = fixTo_2240_dout;
  assign _zz_20241 = _zz_20242[31 : 0];
  assign _zz_20242 = _zz_20243;
  assign _zz_20243 = ($signed(_zz_20244) >>> _zz_1869);
  assign _zz_20244 = _zz_20245;
  assign _zz_20245 = ($signed(_zz_20247) - $signed(_zz_1867));
  assign _zz_20246 = ({8'd0,data_mid_85_imag} <<< 8);
  assign _zz_20247 = {{8{_zz_20246[23]}}, _zz_20246};
  assign _zz_20248 = fixTo_2241_dout;
  assign _zz_20249 = _zz_20250[31 : 0];
  assign _zz_20250 = _zz_20251;
  assign _zz_20251 = ($signed(_zz_20252) >>> _zz_1870);
  assign _zz_20252 = _zz_20253;
  assign _zz_20253 = ($signed(_zz_20255) + $signed(_zz_1866));
  assign _zz_20254 = ({8'd0,data_mid_85_real} <<< 8);
  assign _zz_20255 = {{8{_zz_20254[23]}}, _zz_20254};
  assign _zz_20256 = fixTo_2242_dout;
  assign _zz_20257 = _zz_20258[31 : 0];
  assign _zz_20258 = _zz_20259;
  assign _zz_20259 = ($signed(_zz_20260) >>> _zz_1870);
  assign _zz_20260 = _zz_20261;
  assign _zz_20261 = ($signed(_zz_20263) + $signed(_zz_1867));
  assign _zz_20262 = ({8'd0,data_mid_85_imag} <<< 8);
  assign _zz_20263 = {{8{_zz_20262[23]}}, _zz_20262};
  assign _zz_20264 = fixTo_2243_dout;
  assign _zz_20265 = ($signed(twiddle_factor_table_53_real) + $signed(twiddle_factor_table_53_imag));
  assign _zz_20266 = ($signed(_zz_1873) - $signed(_zz_20267));
  assign _zz_20267 = ($signed(_zz_20268) * $signed(twiddle_factor_table_53_imag));
  assign _zz_20268 = ($signed(data_mid_118_real) + $signed(data_mid_118_imag));
  assign _zz_20269 = fixTo_2244_dout;
  assign _zz_20270 = ($signed(_zz_1873) + $signed(_zz_20271));
  assign _zz_20271 = ($signed(_zz_20272) * $signed(twiddle_factor_table_53_real));
  assign _zz_20272 = ($signed(data_mid_118_imag) - $signed(data_mid_118_real));
  assign _zz_20273 = fixTo_2245_dout;
  assign _zz_20274 = _zz_20275[31 : 0];
  assign _zz_20275 = _zz_20276;
  assign _zz_20276 = ($signed(_zz_20277) >>> _zz_1874);
  assign _zz_20277 = _zz_20278;
  assign _zz_20278 = ($signed(_zz_20280) - $signed(_zz_1871));
  assign _zz_20279 = ({8'd0,data_mid_86_real} <<< 8);
  assign _zz_20280 = {{8{_zz_20279[23]}}, _zz_20279};
  assign _zz_20281 = fixTo_2246_dout;
  assign _zz_20282 = _zz_20283[31 : 0];
  assign _zz_20283 = _zz_20284;
  assign _zz_20284 = ($signed(_zz_20285) >>> _zz_1874);
  assign _zz_20285 = _zz_20286;
  assign _zz_20286 = ($signed(_zz_20288) - $signed(_zz_1872));
  assign _zz_20287 = ({8'd0,data_mid_86_imag} <<< 8);
  assign _zz_20288 = {{8{_zz_20287[23]}}, _zz_20287};
  assign _zz_20289 = fixTo_2247_dout;
  assign _zz_20290 = _zz_20291[31 : 0];
  assign _zz_20291 = _zz_20292;
  assign _zz_20292 = ($signed(_zz_20293) >>> _zz_1875);
  assign _zz_20293 = _zz_20294;
  assign _zz_20294 = ($signed(_zz_20296) + $signed(_zz_1871));
  assign _zz_20295 = ({8'd0,data_mid_86_real} <<< 8);
  assign _zz_20296 = {{8{_zz_20295[23]}}, _zz_20295};
  assign _zz_20297 = fixTo_2248_dout;
  assign _zz_20298 = _zz_20299[31 : 0];
  assign _zz_20299 = _zz_20300;
  assign _zz_20300 = ($signed(_zz_20301) >>> _zz_1875);
  assign _zz_20301 = _zz_20302;
  assign _zz_20302 = ($signed(_zz_20304) + $signed(_zz_1872));
  assign _zz_20303 = ({8'd0,data_mid_86_imag} <<< 8);
  assign _zz_20304 = {{8{_zz_20303[23]}}, _zz_20303};
  assign _zz_20305 = fixTo_2249_dout;
  assign _zz_20306 = ($signed(twiddle_factor_table_54_real) + $signed(twiddle_factor_table_54_imag));
  assign _zz_20307 = ($signed(_zz_1878) - $signed(_zz_20308));
  assign _zz_20308 = ($signed(_zz_20309) * $signed(twiddle_factor_table_54_imag));
  assign _zz_20309 = ($signed(data_mid_119_real) + $signed(data_mid_119_imag));
  assign _zz_20310 = fixTo_2250_dout;
  assign _zz_20311 = ($signed(_zz_1878) + $signed(_zz_20312));
  assign _zz_20312 = ($signed(_zz_20313) * $signed(twiddle_factor_table_54_real));
  assign _zz_20313 = ($signed(data_mid_119_imag) - $signed(data_mid_119_real));
  assign _zz_20314 = fixTo_2251_dout;
  assign _zz_20315 = _zz_20316[31 : 0];
  assign _zz_20316 = _zz_20317;
  assign _zz_20317 = ($signed(_zz_20318) >>> _zz_1879);
  assign _zz_20318 = _zz_20319;
  assign _zz_20319 = ($signed(_zz_20321) - $signed(_zz_1876));
  assign _zz_20320 = ({8'd0,data_mid_87_real} <<< 8);
  assign _zz_20321 = {{8{_zz_20320[23]}}, _zz_20320};
  assign _zz_20322 = fixTo_2252_dout;
  assign _zz_20323 = _zz_20324[31 : 0];
  assign _zz_20324 = _zz_20325;
  assign _zz_20325 = ($signed(_zz_20326) >>> _zz_1879);
  assign _zz_20326 = _zz_20327;
  assign _zz_20327 = ($signed(_zz_20329) - $signed(_zz_1877));
  assign _zz_20328 = ({8'd0,data_mid_87_imag} <<< 8);
  assign _zz_20329 = {{8{_zz_20328[23]}}, _zz_20328};
  assign _zz_20330 = fixTo_2253_dout;
  assign _zz_20331 = _zz_20332[31 : 0];
  assign _zz_20332 = _zz_20333;
  assign _zz_20333 = ($signed(_zz_20334) >>> _zz_1880);
  assign _zz_20334 = _zz_20335;
  assign _zz_20335 = ($signed(_zz_20337) + $signed(_zz_1876));
  assign _zz_20336 = ({8'd0,data_mid_87_real} <<< 8);
  assign _zz_20337 = {{8{_zz_20336[23]}}, _zz_20336};
  assign _zz_20338 = fixTo_2254_dout;
  assign _zz_20339 = _zz_20340[31 : 0];
  assign _zz_20340 = _zz_20341;
  assign _zz_20341 = ($signed(_zz_20342) >>> _zz_1880);
  assign _zz_20342 = _zz_20343;
  assign _zz_20343 = ($signed(_zz_20345) + $signed(_zz_1877));
  assign _zz_20344 = ({8'd0,data_mid_87_imag} <<< 8);
  assign _zz_20345 = {{8{_zz_20344[23]}}, _zz_20344};
  assign _zz_20346 = fixTo_2255_dout;
  assign _zz_20347 = ($signed(twiddle_factor_table_55_real) + $signed(twiddle_factor_table_55_imag));
  assign _zz_20348 = ($signed(_zz_1883) - $signed(_zz_20349));
  assign _zz_20349 = ($signed(_zz_20350) * $signed(twiddle_factor_table_55_imag));
  assign _zz_20350 = ($signed(data_mid_120_real) + $signed(data_mid_120_imag));
  assign _zz_20351 = fixTo_2256_dout;
  assign _zz_20352 = ($signed(_zz_1883) + $signed(_zz_20353));
  assign _zz_20353 = ($signed(_zz_20354) * $signed(twiddle_factor_table_55_real));
  assign _zz_20354 = ($signed(data_mid_120_imag) - $signed(data_mid_120_real));
  assign _zz_20355 = fixTo_2257_dout;
  assign _zz_20356 = _zz_20357[31 : 0];
  assign _zz_20357 = _zz_20358;
  assign _zz_20358 = ($signed(_zz_20359) >>> _zz_1884);
  assign _zz_20359 = _zz_20360;
  assign _zz_20360 = ($signed(_zz_20362) - $signed(_zz_1881));
  assign _zz_20361 = ({8'd0,data_mid_88_real} <<< 8);
  assign _zz_20362 = {{8{_zz_20361[23]}}, _zz_20361};
  assign _zz_20363 = fixTo_2258_dout;
  assign _zz_20364 = _zz_20365[31 : 0];
  assign _zz_20365 = _zz_20366;
  assign _zz_20366 = ($signed(_zz_20367) >>> _zz_1884);
  assign _zz_20367 = _zz_20368;
  assign _zz_20368 = ($signed(_zz_20370) - $signed(_zz_1882));
  assign _zz_20369 = ({8'd0,data_mid_88_imag} <<< 8);
  assign _zz_20370 = {{8{_zz_20369[23]}}, _zz_20369};
  assign _zz_20371 = fixTo_2259_dout;
  assign _zz_20372 = _zz_20373[31 : 0];
  assign _zz_20373 = _zz_20374;
  assign _zz_20374 = ($signed(_zz_20375) >>> _zz_1885);
  assign _zz_20375 = _zz_20376;
  assign _zz_20376 = ($signed(_zz_20378) + $signed(_zz_1881));
  assign _zz_20377 = ({8'd0,data_mid_88_real} <<< 8);
  assign _zz_20378 = {{8{_zz_20377[23]}}, _zz_20377};
  assign _zz_20379 = fixTo_2260_dout;
  assign _zz_20380 = _zz_20381[31 : 0];
  assign _zz_20381 = _zz_20382;
  assign _zz_20382 = ($signed(_zz_20383) >>> _zz_1885);
  assign _zz_20383 = _zz_20384;
  assign _zz_20384 = ($signed(_zz_20386) + $signed(_zz_1882));
  assign _zz_20385 = ({8'd0,data_mid_88_imag} <<< 8);
  assign _zz_20386 = {{8{_zz_20385[23]}}, _zz_20385};
  assign _zz_20387 = fixTo_2261_dout;
  assign _zz_20388 = ($signed(twiddle_factor_table_56_real) + $signed(twiddle_factor_table_56_imag));
  assign _zz_20389 = ($signed(_zz_1888) - $signed(_zz_20390));
  assign _zz_20390 = ($signed(_zz_20391) * $signed(twiddle_factor_table_56_imag));
  assign _zz_20391 = ($signed(data_mid_121_real) + $signed(data_mid_121_imag));
  assign _zz_20392 = fixTo_2262_dout;
  assign _zz_20393 = ($signed(_zz_1888) + $signed(_zz_20394));
  assign _zz_20394 = ($signed(_zz_20395) * $signed(twiddle_factor_table_56_real));
  assign _zz_20395 = ($signed(data_mid_121_imag) - $signed(data_mid_121_real));
  assign _zz_20396 = fixTo_2263_dout;
  assign _zz_20397 = _zz_20398[31 : 0];
  assign _zz_20398 = _zz_20399;
  assign _zz_20399 = ($signed(_zz_20400) >>> _zz_1889);
  assign _zz_20400 = _zz_20401;
  assign _zz_20401 = ($signed(_zz_20403) - $signed(_zz_1886));
  assign _zz_20402 = ({8'd0,data_mid_89_real} <<< 8);
  assign _zz_20403 = {{8{_zz_20402[23]}}, _zz_20402};
  assign _zz_20404 = fixTo_2264_dout;
  assign _zz_20405 = _zz_20406[31 : 0];
  assign _zz_20406 = _zz_20407;
  assign _zz_20407 = ($signed(_zz_20408) >>> _zz_1889);
  assign _zz_20408 = _zz_20409;
  assign _zz_20409 = ($signed(_zz_20411) - $signed(_zz_1887));
  assign _zz_20410 = ({8'd0,data_mid_89_imag} <<< 8);
  assign _zz_20411 = {{8{_zz_20410[23]}}, _zz_20410};
  assign _zz_20412 = fixTo_2265_dout;
  assign _zz_20413 = _zz_20414[31 : 0];
  assign _zz_20414 = _zz_20415;
  assign _zz_20415 = ($signed(_zz_20416) >>> _zz_1890);
  assign _zz_20416 = _zz_20417;
  assign _zz_20417 = ($signed(_zz_20419) + $signed(_zz_1886));
  assign _zz_20418 = ({8'd0,data_mid_89_real} <<< 8);
  assign _zz_20419 = {{8{_zz_20418[23]}}, _zz_20418};
  assign _zz_20420 = fixTo_2266_dout;
  assign _zz_20421 = _zz_20422[31 : 0];
  assign _zz_20422 = _zz_20423;
  assign _zz_20423 = ($signed(_zz_20424) >>> _zz_1890);
  assign _zz_20424 = _zz_20425;
  assign _zz_20425 = ($signed(_zz_20427) + $signed(_zz_1887));
  assign _zz_20426 = ({8'd0,data_mid_89_imag} <<< 8);
  assign _zz_20427 = {{8{_zz_20426[23]}}, _zz_20426};
  assign _zz_20428 = fixTo_2267_dout;
  assign _zz_20429 = ($signed(twiddle_factor_table_57_real) + $signed(twiddle_factor_table_57_imag));
  assign _zz_20430 = ($signed(_zz_1893) - $signed(_zz_20431));
  assign _zz_20431 = ($signed(_zz_20432) * $signed(twiddle_factor_table_57_imag));
  assign _zz_20432 = ($signed(data_mid_122_real) + $signed(data_mid_122_imag));
  assign _zz_20433 = fixTo_2268_dout;
  assign _zz_20434 = ($signed(_zz_1893) + $signed(_zz_20435));
  assign _zz_20435 = ($signed(_zz_20436) * $signed(twiddle_factor_table_57_real));
  assign _zz_20436 = ($signed(data_mid_122_imag) - $signed(data_mid_122_real));
  assign _zz_20437 = fixTo_2269_dout;
  assign _zz_20438 = _zz_20439[31 : 0];
  assign _zz_20439 = _zz_20440;
  assign _zz_20440 = ($signed(_zz_20441) >>> _zz_1894);
  assign _zz_20441 = _zz_20442;
  assign _zz_20442 = ($signed(_zz_20444) - $signed(_zz_1891));
  assign _zz_20443 = ({8'd0,data_mid_90_real} <<< 8);
  assign _zz_20444 = {{8{_zz_20443[23]}}, _zz_20443};
  assign _zz_20445 = fixTo_2270_dout;
  assign _zz_20446 = _zz_20447[31 : 0];
  assign _zz_20447 = _zz_20448;
  assign _zz_20448 = ($signed(_zz_20449) >>> _zz_1894);
  assign _zz_20449 = _zz_20450;
  assign _zz_20450 = ($signed(_zz_20452) - $signed(_zz_1892));
  assign _zz_20451 = ({8'd0,data_mid_90_imag} <<< 8);
  assign _zz_20452 = {{8{_zz_20451[23]}}, _zz_20451};
  assign _zz_20453 = fixTo_2271_dout;
  assign _zz_20454 = _zz_20455[31 : 0];
  assign _zz_20455 = _zz_20456;
  assign _zz_20456 = ($signed(_zz_20457) >>> _zz_1895);
  assign _zz_20457 = _zz_20458;
  assign _zz_20458 = ($signed(_zz_20460) + $signed(_zz_1891));
  assign _zz_20459 = ({8'd0,data_mid_90_real} <<< 8);
  assign _zz_20460 = {{8{_zz_20459[23]}}, _zz_20459};
  assign _zz_20461 = fixTo_2272_dout;
  assign _zz_20462 = _zz_20463[31 : 0];
  assign _zz_20463 = _zz_20464;
  assign _zz_20464 = ($signed(_zz_20465) >>> _zz_1895);
  assign _zz_20465 = _zz_20466;
  assign _zz_20466 = ($signed(_zz_20468) + $signed(_zz_1892));
  assign _zz_20467 = ({8'd0,data_mid_90_imag} <<< 8);
  assign _zz_20468 = {{8{_zz_20467[23]}}, _zz_20467};
  assign _zz_20469 = fixTo_2273_dout;
  assign _zz_20470 = ($signed(twiddle_factor_table_58_real) + $signed(twiddle_factor_table_58_imag));
  assign _zz_20471 = ($signed(_zz_1898) - $signed(_zz_20472));
  assign _zz_20472 = ($signed(_zz_20473) * $signed(twiddle_factor_table_58_imag));
  assign _zz_20473 = ($signed(data_mid_123_real) + $signed(data_mid_123_imag));
  assign _zz_20474 = fixTo_2274_dout;
  assign _zz_20475 = ($signed(_zz_1898) + $signed(_zz_20476));
  assign _zz_20476 = ($signed(_zz_20477) * $signed(twiddle_factor_table_58_real));
  assign _zz_20477 = ($signed(data_mid_123_imag) - $signed(data_mid_123_real));
  assign _zz_20478 = fixTo_2275_dout;
  assign _zz_20479 = _zz_20480[31 : 0];
  assign _zz_20480 = _zz_20481;
  assign _zz_20481 = ($signed(_zz_20482) >>> _zz_1899);
  assign _zz_20482 = _zz_20483;
  assign _zz_20483 = ($signed(_zz_20485) - $signed(_zz_1896));
  assign _zz_20484 = ({8'd0,data_mid_91_real} <<< 8);
  assign _zz_20485 = {{8{_zz_20484[23]}}, _zz_20484};
  assign _zz_20486 = fixTo_2276_dout;
  assign _zz_20487 = _zz_20488[31 : 0];
  assign _zz_20488 = _zz_20489;
  assign _zz_20489 = ($signed(_zz_20490) >>> _zz_1899);
  assign _zz_20490 = _zz_20491;
  assign _zz_20491 = ($signed(_zz_20493) - $signed(_zz_1897));
  assign _zz_20492 = ({8'd0,data_mid_91_imag} <<< 8);
  assign _zz_20493 = {{8{_zz_20492[23]}}, _zz_20492};
  assign _zz_20494 = fixTo_2277_dout;
  assign _zz_20495 = _zz_20496[31 : 0];
  assign _zz_20496 = _zz_20497;
  assign _zz_20497 = ($signed(_zz_20498) >>> _zz_1900);
  assign _zz_20498 = _zz_20499;
  assign _zz_20499 = ($signed(_zz_20501) + $signed(_zz_1896));
  assign _zz_20500 = ({8'd0,data_mid_91_real} <<< 8);
  assign _zz_20501 = {{8{_zz_20500[23]}}, _zz_20500};
  assign _zz_20502 = fixTo_2278_dout;
  assign _zz_20503 = _zz_20504[31 : 0];
  assign _zz_20504 = _zz_20505;
  assign _zz_20505 = ($signed(_zz_20506) >>> _zz_1900);
  assign _zz_20506 = _zz_20507;
  assign _zz_20507 = ($signed(_zz_20509) + $signed(_zz_1897));
  assign _zz_20508 = ({8'd0,data_mid_91_imag} <<< 8);
  assign _zz_20509 = {{8{_zz_20508[23]}}, _zz_20508};
  assign _zz_20510 = fixTo_2279_dout;
  assign _zz_20511 = ($signed(twiddle_factor_table_59_real) + $signed(twiddle_factor_table_59_imag));
  assign _zz_20512 = ($signed(_zz_1903) - $signed(_zz_20513));
  assign _zz_20513 = ($signed(_zz_20514) * $signed(twiddle_factor_table_59_imag));
  assign _zz_20514 = ($signed(data_mid_124_real) + $signed(data_mid_124_imag));
  assign _zz_20515 = fixTo_2280_dout;
  assign _zz_20516 = ($signed(_zz_1903) + $signed(_zz_20517));
  assign _zz_20517 = ($signed(_zz_20518) * $signed(twiddle_factor_table_59_real));
  assign _zz_20518 = ($signed(data_mid_124_imag) - $signed(data_mid_124_real));
  assign _zz_20519 = fixTo_2281_dout;
  assign _zz_20520 = _zz_20521[31 : 0];
  assign _zz_20521 = _zz_20522;
  assign _zz_20522 = ($signed(_zz_20523) >>> _zz_1904);
  assign _zz_20523 = _zz_20524;
  assign _zz_20524 = ($signed(_zz_20526) - $signed(_zz_1901));
  assign _zz_20525 = ({8'd0,data_mid_92_real} <<< 8);
  assign _zz_20526 = {{8{_zz_20525[23]}}, _zz_20525};
  assign _zz_20527 = fixTo_2282_dout;
  assign _zz_20528 = _zz_20529[31 : 0];
  assign _zz_20529 = _zz_20530;
  assign _zz_20530 = ($signed(_zz_20531) >>> _zz_1904);
  assign _zz_20531 = _zz_20532;
  assign _zz_20532 = ($signed(_zz_20534) - $signed(_zz_1902));
  assign _zz_20533 = ({8'd0,data_mid_92_imag} <<< 8);
  assign _zz_20534 = {{8{_zz_20533[23]}}, _zz_20533};
  assign _zz_20535 = fixTo_2283_dout;
  assign _zz_20536 = _zz_20537[31 : 0];
  assign _zz_20537 = _zz_20538;
  assign _zz_20538 = ($signed(_zz_20539) >>> _zz_1905);
  assign _zz_20539 = _zz_20540;
  assign _zz_20540 = ($signed(_zz_20542) + $signed(_zz_1901));
  assign _zz_20541 = ({8'd0,data_mid_92_real} <<< 8);
  assign _zz_20542 = {{8{_zz_20541[23]}}, _zz_20541};
  assign _zz_20543 = fixTo_2284_dout;
  assign _zz_20544 = _zz_20545[31 : 0];
  assign _zz_20545 = _zz_20546;
  assign _zz_20546 = ($signed(_zz_20547) >>> _zz_1905);
  assign _zz_20547 = _zz_20548;
  assign _zz_20548 = ($signed(_zz_20550) + $signed(_zz_1902));
  assign _zz_20549 = ({8'd0,data_mid_92_imag} <<< 8);
  assign _zz_20550 = {{8{_zz_20549[23]}}, _zz_20549};
  assign _zz_20551 = fixTo_2285_dout;
  assign _zz_20552 = ($signed(twiddle_factor_table_60_real) + $signed(twiddle_factor_table_60_imag));
  assign _zz_20553 = ($signed(_zz_1908) - $signed(_zz_20554));
  assign _zz_20554 = ($signed(_zz_20555) * $signed(twiddle_factor_table_60_imag));
  assign _zz_20555 = ($signed(data_mid_125_real) + $signed(data_mid_125_imag));
  assign _zz_20556 = fixTo_2286_dout;
  assign _zz_20557 = ($signed(_zz_1908) + $signed(_zz_20558));
  assign _zz_20558 = ($signed(_zz_20559) * $signed(twiddle_factor_table_60_real));
  assign _zz_20559 = ($signed(data_mid_125_imag) - $signed(data_mid_125_real));
  assign _zz_20560 = fixTo_2287_dout;
  assign _zz_20561 = _zz_20562[31 : 0];
  assign _zz_20562 = _zz_20563;
  assign _zz_20563 = ($signed(_zz_20564) >>> _zz_1909);
  assign _zz_20564 = _zz_20565;
  assign _zz_20565 = ($signed(_zz_20567) - $signed(_zz_1906));
  assign _zz_20566 = ({8'd0,data_mid_93_real} <<< 8);
  assign _zz_20567 = {{8{_zz_20566[23]}}, _zz_20566};
  assign _zz_20568 = fixTo_2288_dout;
  assign _zz_20569 = _zz_20570[31 : 0];
  assign _zz_20570 = _zz_20571;
  assign _zz_20571 = ($signed(_zz_20572) >>> _zz_1909);
  assign _zz_20572 = _zz_20573;
  assign _zz_20573 = ($signed(_zz_20575) - $signed(_zz_1907));
  assign _zz_20574 = ({8'd0,data_mid_93_imag} <<< 8);
  assign _zz_20575 = {{8{_zz_20574[23]}}, _zz_20574};
  assign _zz_20576 = fixTo_2289_dout;
  assign _zz_20577 = _zz_20578[31 : 0];
  assign _zz_20578 = _zz_20579;
  assign _zz_20579 = ($signed(_zz_20580) >>> _zz_1910);
  assign _zz_20580 = _zz_20581;
  assign _zz_20581 = ($signed(_zz_20583) + $signed(_zz_1906));
  assign _zz_20582 = ({8'd0,data_mid_93_real} <<< 8);
  assign _zz_20583 = {{8{_zz_20582[23]}}, _zz_20582};
  assign _zz_20584 = fixTo_2290_dout;
  assign _zz_20585 = _zz_20586[31 : 0];
  assign _zz_20586 = _zz_20587;
  assign _zz_20587 = ($signed(_zz_20588) >>> _zz_1910);
  assign _zz_20588 = _zz_20589;
  assign _zz_20589 = ($signed(_zz_20591) + $signed(_zz_1907));
  assign _zz_20590 = ({8'd0,data_mid_93_imag} <<< 8);
  assign _zz_20591 = {{8{_zz_20590[23]}}, _zz_20590};
  assign _zz_20592 = fixTo_2291_dout;
  assign _zz_20593 = ($signed(twiddle_factor_table_61_real) + $signed(twiddle_factor_table_61_imag));
  assign _zz_20594 = ($signed(_zz_1913) - $signed(_zz_20595));
  assign _zz_20595 = ($signed(_zz_20596) * $signed(twiddle_factor_table_61_imag));
  assign _zz_20596 = ($signed(data_mid_126_real) + $signed(data_mid_126_imag));
  assign _zz_20597 = fixTo_2292_dout;
  assign _zz_20598 = ($signed(_zz_1913) + $signed(_zz_20599));
  assign _zz_20599 = ($signed(_zz_20600) * $signed(twiddle_factor_table_61_real));
  assign _zz_20600 = ($signed(data_mid_126_imag) - $signed(data_mid_126_real));
  assign _zz_20601 = fixTo_2293_dout;
  assign _zz_20602 = _zz_20603[31 : 0];
  assign _zz_20603 = _zz_20604;
  assign _zz_20604 = ($signed(_zz_20605) >>> _zz_1914);
  assign _zz_20605 = _zz_20606;
  assign _zz_20606 = ($signed(_zz_20608) - $signed(_zz_1911));
  assign _zz_20607 = ({8'd0,data_mid_94_real} <<< 8);
  assign _zz_20608 = {{8{_zz_20607[23]}}, _zz_20607};
  assign _zz_20609 = fixTo_2294_dout;
  assign _zz_20610 = _zz_20611[31 : 0];
  assign _zz_20611 = _zz_20612;
  assign _zz_20612 = ($signed(_zz_20613) >>> _zz_1914);
  assign _zz_20613 = _zz_20614;
  assign _zz_20614 = ($signed(_zz_20616) - $signed(_zz_1912));
  assign _zz_20615 = ({8'd0,data_mid_94_imag} <<< 8);
  assign _zz_20616 = {{8{_zz_20615[23]}}, _zz_20615};
  assign _zz_20617 = fixTo_2295_dout;
  assign _zz_20618 = _zz_20619[31 : 0];
  assign _zz_20619 = _zz_20620;
  assign _zz_20620 = ($signed(_zz_20621) >>> _zz_1915);
  assign _zz_20621 = _zz_20622;
  assign _zz_20622 = ($signed(_zz_20624) + $signed(_zz_1911));
  assign _zz_20623 = ({8'd0,data_mid_94_real} <<< 8);
  assign _zz_20624 = {{8{_zz_20623[23]}}, _zz_20623};
  assign _zz_20625 = fixTo_2296_dout;
  assign _zz_20626 = _zz_20627[31 : 0];
  assign _zz_20627 = _zz_20628;
  assign _zz_20628 = ($signed(_zz_20629) >>> _zz_1915);
  assign _zz_20629 = _zz_20630;
  assign _zz_20630 = ($signed(_zz_20632) + $signed(_zz_1912));
  assign _zz_20631 = ({8'd0,data_mid_94_imag} <<< 8);
  assign _zz_20632 = {{8{_zz_20631[23]}}, _zz_20631};
  assign _zz_20633 = fixTo_2297_dout;
  assign _zz_20634 = ($signed(twiddle_factor_table_62_real) + $signed(twiddle_factor_table_62_imag));
  assign _zz_20635 = ($signed(_zz_1918) - $signed(_zz_20636));
  assign _zz_20636 = ($signed(_zz_20637) * $signed(twiddle_factor_table_62_imag));
  assign _zz_20637 = ($signed(data_mid_127_real) + $signed(data_mid_127_imag));
  assign _zz_20638 = fixTo_2298_dout;
  assign _zz_20639 = ($signed(_zz_1918) + $signed(_zz_20640));
  assign _zz_20640 = ($signed(_zz_20641) * $signed(twiddle_factor_table_62_real));
  assign _zz_20641 = ($signed(data_mid_127_imag) - $signed(data_mid_127_real));
  assign _zz_20642 = fixTo_2299_dout;
  assign _zz_20643 = _zz_20644[31 : 0];
  assign _zz_20644 = _zz_20645;
  assign _zz_20645 = ($signed(_zz_20646) >>> _zz_1919);
  assign _zz_20646 = _zz_20647;
  assign _zz_20647 = ($signed(_zz_20649) - $signed(_zz_1916));
  assign _zz_20648 = ({8'd0,data_mid_95_real} <<< 8);
  assign _zz_20649 = {{8{_zz_20648[23]}}, _zz_20648};
  assign _zz_20650 = fixTo_2300_dout;
  assign _zz_20651 = _zz_20652[31 : 0];
  assign _zz_20652 = _zz_20653;
  assign _zz_20653 = ($signed(_zz_20654) >>> _zz_1919);
  assign _zz_20654 = _zz_20655;
  assign _zz_20655 = ($signed(_zz_20657) - $signed(_zz_1917));
  assign _zz_20656 = ({8'd0,data_mid_95_imag} <<< 8);
  assign _zz_20657 = {{8{_zz_20656[23]}}, _zz_20656};
  assign _zz_20658 = fixTo_2301_dout;
  assign _zz_20659 = _zz_20660[31 : 0];
  assign _zz_20660 = _zz_20661;
  assign _zz_20661 = ($signed(_zz_20662) >>> _zz_1920);
  assign _zz_20662 = _zz_20663;
  assign _zz_20663 = ($signed(_zz_20665) + $signed(_zz_1916));
  assign _zz_20664 = ({8'd0,data_mid_95_real} <<< 8);
  assign _zz_20665 = {{8{_zz_20664[23]}}, _zz_20664};
  assign _zz_20666 = fixTo_2302_dout;
  assign _zz_20667 = _zz_20668[31 : 0];
  assign _zz_20668 = _zz_20669;
  assign _zz_20669 = ($signed(_zz_20670) >>> _zz_1920);
  assign _zz_20670 = _zz_20671;
  assign _zz_20671 = ($signed(_zz_20673) + $signed(_zz_1917));
  assign _zz_20672 = ({8'd0,data_mid_95_imag} <<< 8);
  assign _zz_20673 = {{8{_zz_20672[23]}}, _zz_20672};
  assign _zz_20674 = fixTo_2303_dout;
  assign _zz_20675 = ($signed(twiddle_factor_table_63_real) + $signed(twiddle_factor_table_63_imag));
  assign _zz_20676 = ($signed(_zz_1923) - $signed(_zz_20677));
  assign _zz_20677 = ($signed(_zz_20678) * $signed(twiddle_factor_table_63_imag));
  assign _zz_20678 = ($signed(data_mid_64_real) + $signed(data_mid_64_imag));
  assign _zz_20679 = fixTo_2304_dout;
  assign _zz_20680 = ($signed(_zz_1923) + $signed(_zz_20681));
  assign _zz_20681 = ($signed(_zz_20682) * $signed(twiddle_factor_table_63_real));
  assign _zz_20682 = ($signed(data_mid_64_imag) - $signed(data_mid_64_real));
  assign _zz_20683 = fixTo_2305_dout;
  assign _zz_20684 = _zz_20685[31 : 0];
  assign _zz_20685 = _zz_20686;
  assign _zz_20686 = ($signed(_zz_20687) >>> _zz_1924);
  assign _zz_20687 = _zz_20688;
  assign _zz_20688 = ($signed(_zz_20690) - $signed(_zz_1921));
  assign _zz_20689 = ({8'd0,data_mid_0_real} <<< 8);
  assign _zz_20690 = {{8{_zz_20689[23]}}, _zz_20689};
  assign _zz_20691 = fixTo_2306_dout;
  assign _zz_20692 = _zz_20693[31 : 0];
  assign _zz_20693 = _zz_20694;
  assign _zz_20694 = ($signed(_zz_20695) >>> _zz_1924);
  assign _zz_20695 = _zz_20696;
  assign _zz_20696 = ($signed(_zz_20698) - $signed(_zz_1922));
  assign _zz_20697 = ({8'd0,data_mid_0_imag} <<< 8);
  assign _zz_20698 = {{8{_zz_20697[23]}}, _zz_20697};
  assign _zz_20699 = fixTo_2307_dout;
  assign _zz_20700 = _zz_20701[31 : 0];
  assign _zz_20701 = _zz_20702;
  assign _zz_20702 = ($signed(_zz_20703) >>> _zz_1925);
  assign _zz_20703 = _zz_20704;
  assign _zz_20704 = ($signed(_zz_20706) + $signed(_zz_1921));
  assign _zz_20705 = ({8'd0,data_mid_0_real} <<< 8);
  assign _zz_20706 = {{8{_zz_20705[23]}}, _zz_20705};
  assign _zz_20707 = fixTo_2308_dout;
  assign _zz_20708 = _zz_20709[31 : 0];
  assign _zz_20709 = _zz_20710;
  assign _zz_20710 = ($signed(_zz_20711) >>> _zz_1925);
  assign _zz_20711 = _zz_20712;
  assign _zz_20712 = ($signed(_zz_20714) + $signed(_zz_1922));
  assign _zz_20713 = ({8'd0,data_mid_0_imag} <<< 8);
  assign _zz_20714 = {{8{_zz_20713[23]}}, _zz_20713};
  assign _zz_20715 = fixTo_2309_dout;
  assign _zz_20716 = ($signed(twiddle_factor_table_64_real) + $signed(twiddle_factor_table_64_imag));
  assign _zz_20717 = ($signed(_zz_1928) - $signed(_zz_20718));
  assign _zz_20718 = ($signed(_zz_20719) * $signed(twiddle_factor_table_64_imag));
  assign _zz_20719 = ($signed(data_mid_65_real) + $signed(data_mid_65_imag));
  assign _zz_20720 = fixTo_2310_dout;
  assign _zz_20721 = ($signed(_zz_1928) + $signed(_zz_20722));
  assign _zz_20722 = ($signed(_zz_20723) * $signed(twiddle_factor_table_64_real));
  assign _zz_20723 = ($signed(data_mid_65_imag) - $signed(data_mid_65_real));
  assign _zz_20724 = fixTo_2311_dout;
  assign _zz_20725 = _zz_20726[31 : 0];
  assign _zz_20726 = _zz_20727;
  assign _zz_20727 = ($signed(_zz_20728) >>> _zz_1929);
  assign _zz_20728 = _zz_20729;
  assign _zz_20729 = ($signed(_zz_20731) - $signed(_zz_1926));
  assign _zz_20730 = ({8'd0,data_mid_1_real} <<< 8);
  assign _zz_20731 = {{8{_zz_20730[23]}}, _zz_20730};
  assign _zz_20732 = fixTo_2312_dout;
  assign _zz_20733 = _zz_20734[31 : 0];
  assign _zz_20734 = _zz_20735;
  assign _zz_20735 = ($signed(_zz_20736) >>> _zz_1929);
  assign _zz_20736 = _zz_20737;
  assign _zz_20737 = ($signed(_zz_20739) - $signed(_zz_1927));
  assign _zz_20738 = ({8'd0,data_mid_1_imag} <<< 8);
  assign _zz_20739 = {{8{_zz_20738[23]}}, _zz_20738};
  assign _zz_20740 = fixTo_2313_dout;
  assign _zz_20741 = _zz_20742[31 : 0];
  assign _zz_20742 = _zz_20743;
  assign _zz_20743 = ($signed(_zz_20744) >>> _zz_1930);
  assign _zz_20744 = _zz_20745;
  assign _zz_20745 = ($signed(_zz_20747) + $signed(_zz_1926));
  assign _zz_20746 = ({8'd0,data_mid_1_real} <<< 8);
  assign _zz_20747 = {{8{_zz_20746[23]}}, _zz_20746};
  assign _zz_20748 = fixTo_2314_dout;
  assign _zz_20749 = _zz_20750[31 : 0];
  assign _zz_20750 = _zz_20751;
  assign _zz_20751 = ($signed(_zz_20752) >>> _zz_1930);
  assign _zz_20752 = _zz_20753;
  assign _zz_20753 = ($signed(_zz_20755) + $signed(_zz_1927));
  assign _zz_20754 = ({8'd0,data_mid_1_imag} <<< 8);
  assign _zz_20755 = {{8{_zz_20754[23]}}, _zz_20754};
  assign _zz_20756 = fixTo_2315_dout;
  assign _zz_20757 = ($signed(twiddle_factor_table_65_real) + $signed(twiddle_factor_table_65_imag));
  assign _zz_20758 = ($signed(_zz_1933) - $signed(_zz_20759));
  assign _zz_20759 = ($signed(_zz_20760) * $signed(twiddle_factor_table_65_imag));
  assign _zz_20760 = ($signed(data_mid_66_real) + $signed(data_mid_66_imag));
  assign _zz_20761 = fixTo_2316_dout;
  assign _zz_20762 = ($signed(_zz_1933) + $signed(_zz_20763));
  assign _zz_20763 = ($signed(_zz_20764) * $signed(twiddle_factor_table_65_real));
  assign _zz_20764 = ($signed(data_mid_66_imag) - $signed(data_mid_66_real));
  assign _zz_20765 = fixTo_2317_dout;
  assign _zz_20766 = _zz_20767[31 : 0];
  assign _zz_20767 = _zz_20768;
  assign _zz_20768 = ($signed(_zz_20769) >>> _zz_1934);
  assign _zz_20769 = _zz_20770;
  assign _zz_20770 = ($signed(_zz_20772) - $signed(_zz_1931));
  assign _zz_20771 = ({8'd0,data_mid_2_real} <<< 8);
  assign _zz_20772 = {{8{_zz_20771[23]}}, _zz_20771};
  assign _zz_20773 = fixTo_2318_dout;
  assign _zz_20774 = _zz_20775[31 : 0];
  assign _zz_20775 = _zz_20776;
  assign _zz_20776 = ($signed(_zz_20777) >>> _zz_1934);
  assign _zz_20777 = _zz_20778;
  assign _zz_20778 = ($signed(_zz_20780) - $signed(_zz_1932));
  assign _zz_20779 = ({8'd0,data_mid_2_imag} <<< 8);
  assign _zz_20780 = {{8{_zz_20779[23]}}, _zz_20779};
  assign _zz_20781 = fixTo_2319_dout;
  assign _zz_20782 = _zz_20783[31 : 0];
  assign _zz_20783 = _zz_20784;
  assign _zz_20784 = ($signed(_zz_20785) >>> _zz_1935);
  assign _zz_20785 = _zz_20786;
  assign _zz_20786 = ($signed(_zz_20788) + $signed(_zz_1931));
  assign _zz_20787 = ({8'd0,data_mid_2_real} <<< 8);
  assign _zz_20788 = {{8{_zz_20787[23]}}, _zz_20787};
  assign _zz_20789 = fixTo_2320_dout;
  assign _zz_20790 = _zz_20791[31 : 0];
  assign _zz_20791 = _zz_20792;
  assign _zz_20792 = ($signed(_zz_20793) >>> _zz_1935);
  assign _zz_20793 = _zz_20794;
  assign _zz_20794 = ($signed(_zz_20796) + $signed(_zz_1932));
  assign _zz_20795 = ({8'd0,data_mid_2_imag} <<< 8);
  assign _zz_20796 = {{8{_zz_20795[23]}}, _zz_20795};
  assign _zz_20797 = fixTo_2321_dout;
  assign _zz_20798 = ($signed(twiddle_factor_table_66_real) + $signed(twiddle_factor_table_66_imag));
  assign _zz_20799 = ($signed(_zz_1938) - $signed(_zz_20800));
  assign _zz_20800 = ($signed(_zz_20801) * $signed(twiddle_factor_table_66_imag));
  assign _zz_20801 = ($signed(data_mid_67_real) + $signed(data_mid_67_imag));
  assign _zz_20802 = fixTo_2322_dout;
  assign _zz_20803 = ($signed(_zz_1938) + $signed(_zz_20804));
  assign _zz_20804 = ($signed(_zz_20805) * $signed(twiddle_factor_table_66_real));
  assign _zz_20805 = ($signed(data_mid_67_imag) - $signed(data_mid_67_real));
  assign _zz_20806 = fixTo_2323_dout;
  assign _zz_20807 = _zz_20808[31 : 0];
  assign _zz_20808 = _zz_20809;
  assign _zz_20809 = ($signed(_zz_20810) >>> _zz_1939);
  assign _zz_20810 = _zz_20811;
  assign _zz_20811 = ($signed(_zz_20813) - $signed(_zz_1936));
  assign _zz_20812 = ({8'd0,data_mid_3_real} <<< 8);
  assign _zz_20813 = {{8{_zz_20812[23]}}, _zz_20812};
  assign _zz_20814 = fixTo_2324_dout;
  assign _zz_20815 = _zz_20816[31 : 0];
  assign _zz_20816 = _zz_20817;
  assign _zz_20817 = ($signed(_zz_20818) >>> _zz_1939);
  assign _zz_20818 = _zz_20819;
  assign _zz_20819 = ($signed(_zz_20821) - $signed(_zz_1937));
  assign _zz_20820 = ({8'd0,data_mid_3_imag} <<< 8);
  assign _zz_20821 = {{8{_zz_20820[23]}}, _zz_20820};
  assign _zz_20822 = fixTo_2325_dout;
  assign _zz_20823 = _zz_20824[31 : 0];
  assign _zz_20824 = _zz_20825;
  assign _zz_20825 = ($signed(_zz_20826) >>> _zz_1940);
  assign _zz_20826 = _zz_20827;
  assign _zz_20827 = ($signed(_zz_20829) + $signed(_zz_1936));
  assign _zz_20828 = ({8'd0,data_mid_3_real} <<< 8);
  assign _zz_20829 = {{8{_zz_20828[23]}}, _zz_20828};
  assign _zz_20830 = fixTo_2326_dout;
  assign _zz_20831 = _zz_20832[31 : 0];
  assign _zz_20832 = _zz_20833;
  assign _zz_20833 = ($signed(_zz_20834) >>> _zz_1940);
  assign _zz_20834 = _zz_20835;
  assign _zz_20835 = ($signed(_zz_20837) + $signed(_zz_1937));
  assign _zz_20836 = ({8'd0,data_mid_3_imag} <<< 8);
  assign _zz_20837 = {{8{_zz_20836[23]}}, _zz_20836};
  assign _zz_20838 = fixTo_2327_dout;
  assign _zz_20839 = ($signed(twiddle_factor_table_67_real) + $signed(twiddle_factor_table_67_imag));
  assign _zz_20840 = ($signed(_zz_1943) - $signed(_zz_20841));
  assign _zz_20841 = ($signed(_zz_20842) * $signed(twiddle_factor_table_67_imag));
  assign _zz_20842 = ($signed(data_mid_68_real) + $signed(data_mid_68_imag));
  assign _zz_20843 = fixTo_2328_dout;
  assign _zz_20844 = ($signed(_zz_1943) + $signed(_zz_20845));
  assign _zz_20845 = ($signed(_zz_20846) * $signed(twiddle_factor_table_67_real));
  assign _zz_20846 = ($signed(data_mid_68_imag) - $signed(data_mid_68_real));
  assign _zz_20847 = fixTo_2329_dout;
  assign _zz_20848 = _zz_20849[31 : 0];
  assign _zz_20849 = _zz_20850;
  assign _zz_20850 = ($signed(_zz_20851) >>> _zz_1944);
  assign _zz_20851 = _zz_20852;
  assign _zz_20852 = ($signed(_zz_20854) - $signed(_zz_1941));
  assign _zz_20853 = ({8'd0,data_mid_4_real} <<< 8);
  assign _zz_20854 = {{8{_zz_20853[23]}}, _zz_20853};
  assign _zz_20855 = fixTo_2330_dout;
  assign _zz_20856 = _zz_20857[31 : 0];
  assign _zz_20857 = _zz_20858;
  assign _zz_20858 = ($signed(_zz_20859) >>> _zz_1944);
  assign _zz_20859 = _zz_20860;
  assign _zz_20860 = ($signed(_zz_20862) - $signed(_zz_1942));
  assign _zz_20861 = ({8'd0,data_mid_4_imag} <<< 8);
  assign _zz_20862 = {{8{_zz_20861[23]}}, _zz_20861};
  assign _zz_20863 = fixTo_2331_dout;
  assign _zz_20864 = _zz_20865[31 : 0];
  assign _zz_20865 = _zz_20866;
  assign _zz_20866 = ($signed(_zz_20867) >>> _zz_1945);
  assign _zz_20867 = _zz_20868;
  assign _zz_20868 = ($signed(_zz_20870) + $signed(_zz_1941));
  assign _zz_20869 = ({8'd0,data_mid_4_real} <<< 8);
  assign _zz_20870 = {{8{_zz_20869[23]}}, _zz_20869};
  assign _zz_20871 = fixTo_2332_dout;
  assign _zz_20872 = _zz_20873[31 : 0];
  assign _zz_20873 = _zz_20874;
  assign _zz_20874 = ($signed(_zz_20875) >>> _zz_1945);
  assign _zz_20875 = _zz_20876;
  assign _zz_20876 = ($signed(_zz_20878) + $signed(_zz_1942));
  assign _zz_20877 = ({8'd0,data_mid_4_imag} <<< 8);
  assign _zz_20878 = {{8{_zz_20877[23]}}, _zz_20877};
  assign _zz_20879 = fixTo_2333_dout;
  assign _zz_20880 = ($signed(twiddle_factor_table_68_real) + $signed(twiddle_factor_table_68_imag));
  assign _zz_20881 = ($signed(_zz_1948) - $signed(_zz_20882));
  assign _zz_20882 = ($signed(_zz_20883) * $signed(twiddle_factor_table_68_imag));
  assign _zz_20883 = ($signed(data_mid_69_real) + $signed(data_mid_69_imag));
  assign _zz_20884 = fixTo_2334_dout;
  assign _zz_20885 = ($signed(_zz_1948) + $signed(_zz_20886));
  assign _zz_20886 = ($signed(_zz_20887) * $signed(twiddle_factor_table_68_real));
  assign _zz_20887 = ($signed(data_mid_69_imag) - $signed(data_mid_69_real));
  assign _zz_20888 = fixTo_2335_dout;
  assign _zz_20889 = _zz_20890[31 : 0];
  assign _zz_20890 = _zz_20891;
  assign _zz_20891 = ($signed(_zz_20892) >>> _zz_1949);
  assign _zz_20892 = _zz_20893;
  assign _zz_20893 = ($signed(_zz_20895) - $signed(_zz_1946));
  assign _zz_20894 = ({8'd0,data_mid_5_real} <<< 8);
  assign _zz_20895 = {{8{_zz_20894[23]}}, _zz_20894};
  assign _zz_20896 = fixTo_2336_dout;
  assign _zz_20897 = _zz_20898[31 : 0];
  assign _zz_20898 = _zz_20899;
  assign _zz_20899 = ($signed(_zz_20900) >>> _zz_1949);
  assign _zz_20900 = _zz_20901;
  assign _zz_20901 = ($signed(_zz_20903) - $signed(_zz_1947));
  assign _zz_20902 = ({8'd0,data_mid_5_imag} <<< 8);
  assign _zz_20903 = {{8{_zz_20902[23]}}, _zz_20902};
  assign _zz_20904 = fixTo_2337_dout;
  assign _zz_20905 = _zz_20906[31 : 0];
  assign _zz_20906 = _zz_20907;
  assign _zz_20907 = ($signed(_zz_20908) >>> _zz_1950);
  assign _zz_20908 = _zz_20909;
  assign _zz_20909 = ($signed(_zz_20911) + $signed(_zz_1946));
  assign _zz_20910 = ({8'd0,data_mid_5_real} <<< 8);
  assign _zz_20911 = {{8{_zz_20910[23]}}, _zz_20910};
  assign _zz_20912 = fixTo_2338_dout;
  assign _zz_20913 = _zz_20914[31 : 0];
  assign _zz_20914 = _zz_20915;
  assign _zz_20915 = ($signed(_zz_20916) >>> _zz_1950);
  assign _zz_20916 = _zz_20917;
  assign _zz_20917 = ($signed(_zz_20919) + $signed(_zz_1947));
  assign _zz_20918 = ({8'd0,data_mid_5_imag} <<< 8);
  assign _zz_20919 = {{8{_zz_20918[23]}}, _zz_20918};
  assign _zz_20920 = fixTo_2339_dout;
  assign _zz_20921 = ($signed(twiddle_factor_table_69_real) + $signed(twiddle_factor_table_69_imag));
  assign _zz_20922 = ($signed(_zz_1953) - $signed(_zz_20923));
  assign _zz_20923 = ($signed(_zz_20924) * $signed(twiddle_factor_table_69_imag));
  assign _zz_20924 = ($signed(data_mid_70_real) + $signed(data_mid_70_imag));
  assign _zz_20925 = fixTo_2340_dout;
  assign _zz_20926 = ($signed(_zz_1953) + $signed(_zz_20927));
  assign _zz_20927 = ($signed(_zz_20928) * $signed(twiddle_factor_table_69_real));
  assign _zz_20928 = ($signed(data_mid_70_imag) - $signed(data_mid_70_real));
  assign _zz_20929 = fixTo_2341_dout;
  assign _zz_20930 = _zz_20931[31 : 0];
  assign _zz_20931 = _zz_20932;
  assign _zz_20932 = ($signed(_zz_20933) >>> _zz_1954);
  assign _zz_20933 = _zz_20934;
  assign _zz_20934 = ($signed(_zz_20936) - $signed(_zz_1951));
  assign _zz_20935 = ({8'd0,data_mid_6_real} <<< 8);
  assign _zz_20936 = {{8{_zz_20935[23]}}, _zz_20935};
  assign _zz_20937 = fixTo_2342_dout;
  assign _zz_20938 = _zz_20939[31 : 0];
  assign _zz_20939 = _zz_20940;
  assign _zz_20940 = ($signed(_zz_20941) >>> _zz_1954);
  assign _zz_20941 = _zz_20942;
  assign _zz_20942 = ($signed(_zz_20944) - $signed(_zz_1952));
  assign _zz_20943 = ({8'd0,data_mid_6_imag} <<< 8);
  assign _zz_20944 = {{8{_zz_20943[23]}}, _zz_20943};
  assign _zz_20945 = fixTo_2343_dout;
  assign _zz_20946 = _zz_20947[31 : 0];
  assign _zz_20947 = _zz_20948;
  assign _zz_20948 = ($signed(_zz_20949) >>> _zz_1955);
  assign _zz_20949 = _zz_20950;
  assign _zz_20950 = ($signed(_zz_20952) + $signed(_zz_1951));
  assign _zz_20951 = ({8'd0,data_mid_6_real} <<< 8);
  assign _zz_20952 = {{8{_zz_20951[23]}}, _zz_20951};
  assign _zz_20953 = fixTo_2344_dout;
  assign _zz_20954 = _zz_20955[31 : 0];
  assign _zz_20955 = _zz_20956;
  assign _zz_20956 = ($signed(_zz_20957) >>> _zz_1955);
  assign _zz_20957 = _zz_20958;
  assign _zz_20958 = ($signed(_zz_20960) + $signed(_zz_1952));
  assign _zz_20959 = ({8'd0,data_mid_6_imag} <<< 8);
  assign _zz_20960 = {{8{_zz_20959[23]}}, _zz_20959};
  assign _zz_20961 = fixTo_2345_dout;
  assign _zz_20962 = ($signed(twiddle_factor_table_70_real) + $signed(twiddle_factor_table_70_imag));
  assign _zz_20963 = ($signed(_zz_1958) - $signed(_zz_20964));
  assign _zz_20964 = ($signed(_zz_20965) * $signed(twiddle_factor_table_70_imag));
  assign _zz_20965 = ($signed(data_mid_71_real) + $signed(data_mid_71_imag));
  assign _zz_20966 = fixTo_2346_dout;
  assign _zz_20967 = ($signed(_zz_1958) + $signed(_zz_20968));
  assign _zz_20968 = ($signed(_zz_20969) * $signed(twiddle_factor_table_70_real));
  assign _zz_20969 = ($signed(data_mid_71_imag) - $signed(data_mid_71_real));
  assign _zz_20970 = fixTo_2347_dout;
  assign _zz_20971 = _zz_20972[31 : 0];
  assign _zz_20972 = _zz_20973;
  assign _zz_20973 = ($signed(_zz_20974) >>> _zz_1959);
  assign _zz_20974 = _zz_20975;
  assign _zz_20975 = ($signed(_zz_20977) - $signed(_zz_1956));
  assign _zz_20976 = ({8'd0,data_mid_7_real} <<< 8);
  assign _zz_20977 = {{8{_zz_20976[23]}}, _zz_20976};
  assign _zz_20978 = fixTo_2348_dout;
  assign _zz_20979 = _zz_20980[31 : 0];
  assign _zz_20980 = _zz_20981;
  assign _zz_20981 = ($signed(_zz_20982) >>> _zz_1959);
  assign _zz_20982 = _zz_20983;
  assign _zz_20983 = ($signed(_zz_20985) - $signed(_zz_1957));
  assign _zz_20984 = ({8'd0,data_mid_7_imag} <<< 8);
  assign _zz_20985 = {{8{_zz_20984[23]}}, _zz_20984};
  assign _zz_20986 = fixTo_2349_dout;
  assign _zz_20987 = _zz_20988[31 : 0];
  assign _zz_20988 = _zz_20989;
  assign _zz_20989 = ($signed(_zz_20990) >>> _zz_1960);
  assign _zz_20990 = _zz_20991;
  assign _zz_20991 = ($signed(_zz_20993) + $signed(_zz_1956));
  assign _zz_20992 = ({8'd0,data_mid_7_real} <<< 8);
  assign _zz_20993 = {{8{_zz_20992[23]}}, _zz_20992};
  assign _zz_20994 = fixTo_2350_dout;
  assign _zz_20995 = _zz_20996[31 : 0];
  assign _zz_20996 = _zz_20997;
  assign _zz_20997 = ($signed(_zz_20998) >>> _zz_1960);
  assign _zz_20998 = _zz_20999;
  assign _zz_20999 = ($signed(_zz_21001) + $signed(_zz_1957));
  assign _zz_21000 = ({8'd0,data_mid_7_imag} <<< 8);
  assign _zz_21001 = {{8{_zz_21000[23]}}, _zz_21000};
  assign _zz_21002 = fixTo_2351_dout;
  assign _zz_21003 = ($signed(twiddle_factor_table_71_real) + $signed(twiddle_factor_table_71_imag));
  assign _zz_21004 = ($signed(_zz_1963) - $signed(_zz_21005));
  assign _zz_21005 = ($signed(_zz_21006) * $signed(twiddle_factor_table_71_imag));
  assign _zz_21006 = ($signed(data_mid_72_real) + $signed(data_mid_72_imag));
  assign _zz_21007 = fixTo_2352_dout;
  assign _zz_21008 = ($signed(_zz_1963) + $signed(_zz_21009));
  assign _zz_21009 = ($signed(_zz_21010) * $signed(twiddle_factor_table_71_real));
  assign _zz_21010 = ($signed(data_mid_72_imag) - $signed(data_mid_72_real));
  assign _zz_21011 = fixTo_2353_dout;
  assign _zz_21012 = _zz_21013[31 : 0];
  assign _zz_21013 = _zz_21014;
  assign _zz_21014 = ($signed(_zz_21015) >>> _zz_1964);
  assign _zz_21015 = _zz_21016;
  assign _zz_21016 = ($signed(_zz_21018) - $signed(_zz_1961));
  assign _zz_21017 = ({8'd0,data_mid_8_real} <<< 8);
  assign _zz_21018 = {{8{_zz_21017[23]}}, _zz_21017};
  assign _zz_21019 = fixTo_2354_dout;
  assign _zz_21020 = _zz_21021[31 : 0];
  assign _zz_21021 = _zz_21022;
  assign _zz_21022 = ($signed(_zz_21023) >>> _zz_1964);
  assign _zz_21023 = _zz_21024;
  assign _zz_21024 = ($signed(_zz_21026) - $signed(_zz_1962));
  assign _zz_21025 = ({8'd0,data_mid_8_imag} <<< 8);
  assign _zz_21026 = {{8{_zz_21025[23]}}, _zz_21025};
  assign _zz_21027 = fixTo_2355_dout;
  assign _zz_21028 = _zz_21029[31 : 0];
  assign _zz_21029 = _zz_21030;
  assign _zz_21030 = ($signed(_zz_21031) >>> _zz_1965);
  assign _zz_21031 = _zz_21032;
  assign _zz_21032 = ($signed(_zz_21034) + $signed(_zz_1961));
  assign _zz_21033 = ({8'd0,data_mid_8_real} <<< 8);
  assign _zz_21034 = {{8{_zz_21033[23]}}, _zz_21033};
  assign _zz_21035 = fixTo_2356_dout;
  assign _zz_21036 = _zz_21037[31 : 0];
  assign _zz_21037 = _zz_21038;
  assign _zz_21038 = ($signed(_zz_21039) >>> _zz_1965);
  assign _zz_21039 = _zz_21040;
  assign _zz_21040 = ($signed(_zz_21042) + $signed(_zz_1962));
  assign _zz_21041 = ({8'd0,data_mid_8_imag} <<< 8);
  assign _zz_21042 = {{8{_zz_21041[23]}}, _zz_21041};
  assign _zz_21043 = fixTo_2357_dout;
  assign _zz_21044 = ($signed(twiddle_factor_table_72_real) + $signed(twiddle_factor_table_72_imag));
  assign _zz_21045 = ($signed(_zz_1968) - $signed(_zz_21046));
  assign _zz_21046 = ($signed(_zz_21047) * $signed(twiddle_factor_table_72_imag));
  assign _zz_21047 = ($signed(data_mid_73_real) + $signed(data_mid_73_imag));
  assign _zz_21048 = fixTo_2358_dout;
  assign _zz_21049 = ($signed(_zz_1968) + $signed(_zz_21050));
  assign _zz_21050 = ($signed(_zz_21051) * $signed(twiddle_factor_table_72_real));
  assign _zz_21051 = ($signed(data_mid_73_imag) - $signed(data_mid_73_real));
  assign _zz_21052 = fixTo_2359_dout;
  assign _zz_21053 = _zz_21054[31 : 0];
  assign _zz_21054 = _zz_21055;
  assign _zz_21055 = ($signed(_zz_21056) >>> _zz_1969);
  assign _zz_21056 = _zz_21057;
  assign _zz_21057 = ($signed(_zz_21059) - $signed(_zz_1966));
  assign _zz_21058 = ({8'd0,data_mid_9_real} <<< 8);
  assign _zz_21059 = {{8{_zz_21058[23]}}, _zz_21058};
  assign _zz_21060 = fixTo_2360_dout;
  assign _zz_21061 = _zz_21062[31 : 0];
  assign _zz_21062 = _zz_21063;
  assign _zz_21063 = ($signed(_zz_21064) >>> _zz_1969);
  assign _zz_21064 = _zz_21065;
  assign _zz_21065 = ($signed(_zz_21067) - $signed(_zz_1967));
  assign _zz_21066 = ({8'd0,data_mid_9_imag} <<< 8);
  assign _zz_21067 = {{8{_zz_21066[23]}}, _zz_21066};
  assign _zz_21068 = fixTo_2361_dout;
  assign _zz_21069 = _zz_21070[31 : 0];
  assign _zz_21070 = _zz_21071;
  assign _zz_21071 = ($signed(_zz_21072) >>> _zz_1970);
  assign _zz_21072 = _zz_21073;
  assign _zz_21073 = ($signed(_zz_21075) + $signed(_zz_1966));
  assign _zz_21074 = ({8'd0,data_mid_9_real} <<< 8);
  assign _zz_21075 = {{8{_zz_21074[23]}}, _zz_21074};
  assign _zz_21076 = fixTo_2362_dout;
  assign _zz_21077 = _zz_21078[31 : 0];
  assign _zz_21078 = _zz_21079;
  assign _zz_21079 = ($signed(_zz_21080) >>> _zz_1970);
  assign _zz_21080 = _zz_21081;
  assign _zz_21081 = ($signed(_zz_21083) + $signed(_zz_1967));
  assign _zz_21082 = ({8'd0,data_mid_9_imag} <<< 8);
  assign _zz_21083 = {{8{_zz_21082[23]}}, _zz_21082};
  assign _zz_21084 = fixTo_2363_dout;
  assign _zz_21085 = ($signed(twiddle_factor_table_73_real) + $signed(twiddle_factor_table_73_imag));
  assign _zz_21086 = ($signed(_zz_1973) - $signed(_zz_21087));
  assign _zz_21087 = ($signed(_zz_21088) * $signed(twiddle_factor_table_73_imag));
  assign _zz_21088 = ($signed(data_mid_74_real) + $signed(data_mid_74_imag));
  assign _zz_21089 = fixTo_2364_dout;
  assign _zz_21090 = ($signed(_zz_1973) + $signed(_zz_21091));
  assign _zz_21091 = ($signed(_zz_21092) * $signed(twiddle_factor_table_73_real));
  assign _zz_21092 = ($signed(data_mid_74_imag) - $signed(data_mid_74_real));
  assign _zz_21093 = fixTo_2365_dout;
  assign _zz_21094 = _zz_21095[31 : 0];
  assign _zz_21095 = _zz_21096;
  assign _zz_21096 = ($signed(_zz_21097) >>> _zz_1974);
  assign _zz_21097 = _zz_21098;
  assign _zz_21098 = ($signed(_zz_21100) - $signed(_zz_1971));
  assign _zz_21099 = ({8'd0,data_mid_10_real} <<< 8);
  assign _zz_21100 = {{8{_zz_21099[23]}}, _zz_21099};
  assign _zz_21101 = fixTo_2366_dout;
  assign _zz_21102 = _zz_21103[31 : 0];
  assign _zz_21103 = _zz_21104;
  assign _zz_21104 = ($signed(_zz_21105) >>> _zz_1974);
  assign _zz_21105 = _zz_21106;
  assign _zz_21106 = ($signed(_zz_21108) - $signed(_zz_1972));
  assign _zz_21107 = ({8'd0,data_mid_10_imag} <<< 8);
  assign _zz_21108 = {{8{_zz_21107[23]}}, _zz_21107};
  assign _zz_21109 = fixTo_2367_dout;
  assign _zz_21110 = _zz_21111[31 : 0];
  assign _zz_21111 = _zz_21112;
  assign _zz_21112 = ($signed(_zz_21113) >>> _zz_1975);
  assign _zz_21113 = _zz_21114;
  assign _zz_21114 = ($signed(_zz_21116) + $signed(_zz_1971));
  assign _zz_21115 = ({8'd0,data_mid_10_real} <<< 8);
  assign _zz_21116 = {{8{_zz_21115[23]}}, _zz_21115};
  assign _zz_21117 = fixTo_2368_dout;
  assign _zz_21118 = _zz_21119[31 : 0];
  assign _zz_21119 = _zz_21120;
  assign _zz_21120 = ($signed(_zz_21121) >>> _zz_1975);
  assign _zz_21121 = _zz_21122;
  assign _zz_21122 = ($signed(_zz_21124) + $signed(_zz_1972));
  assign _zz_21123 = ({8'd0,data_mid_10_imag} <<< 8);
  assign _zz_21124 = {{8{_zz_21123[23]}}, _zz_21123};
  assign _zz_21125 = fixTo_2369_dout;
  assign _zz_21126 = ($signed(twiddle_factor_table_74_real) + $signed(twiddle_factor_table_74_imag));
  assign _zz_21127 = ($signed(_zz_1978) - $signed(_zz_21128));
  assign _zz_21128 = ($signed(_zz_21129) * $signed(twiddle_factor_table_74_imag));
  assign _zz_21129 = ($signed(data_mid_75_real) + $signed(data_mid_75_imag));
  assign _zz_21130 = fixTo_2370_dout;
  assign _zz_21131 = ($signed(_zz_1978) + $signed(_zz_21132));
  assign _zz_21132 = ($signed(_zz_21133) * $signed(twiddle_factor_table_74_real));
  assign _zz_21133 = ($signed(data_mid_75_imag) - $signed(data_mid_75_real));
  assign _zz_21134 = fixTo_2371_dout;
  assign _zz_21135 = _zz_21136[31 : 0];
  assign _zz_21136 = _zz_21137;
  assign _zz_21137 = ($signed(_zz_21138) >>> _zz_1979);
  assign _zz_21138 = _zz_21139;
  assign _zz_21139 = ($signed(_zz_21141) - $signed(_zz_1976));
  assign _zz_21140 = ({8'd0,data_mid_11_real} <<< 8);
  assign _zz_21141 = {{8{_zz_21140[23]}}, _zz_21140};
  assign _zz_21142 = fixTo_2372_dout;
  assign _zz_21143 = _zz_21144[31 : 0];
  assign _zz_21144 = _zz_21145;
  assign _zz_21145 = ($signed(_zz_21146) >>> _zz_1979);
  assign _zz_21146 = _zz_21147;
  assign _zz_21147 = ($signed(_zz_21149) - $signed(_zz_1977));
  assign _zz_21148 = ({8'd0,data_mid_11_imag} <<< 8);
  assign _zz_21149 = {{8{_zz_21148[23]}}, _zz_21148};
  assign _zz_21150 = fixTo_2373_dout;
  assign _zz_21151 = _zz_21152[31 : 0];
  assign _zz_21152 = _zz_21153;
  assign _zz_21153 = ($signed(_zz_21154) >>> _zz_1980);
  assign _zz_21154 = _zz_21155;
  assign _zz_21155 = ($signed(_zz_21157) + $signed(_zz_1976));
  assign _zz_21156 = ({8'd0,data_mid_11_real} <<< 8);
  assign _zz_21157 = {{8{_zz_21156[23]}}, _zz_21156};
  assign _zz_21158 = fixTo_2374_dout;
  assign _zz_21159 = _zz_21160[31 : 0];
  assign _zz_21160 = _zz_21161;
  assign _zz_21161 = ($signed(_zz_21162) >>> _zz_1980);
  assign _zz_21162 = _zz_21163;
  assign _zz_21163 = ($signed(_zz_21165) + $signed(_zz_1977));
  assign _zz_21164 = ({8'd0,data_mid_11_imag} <<< 8);
  assign _zz_21165 = {{8{_zz_21164[23]}}, _zz_21164};
  assign _zz_21166 = fixTo_2375_dout;
  assign _zz_21167 = ($signed(twiddle_factor_table_75_real) + $signed(twiddle_factor_table_75_imag));
  assign _zz_21168 = ($signed(_zz_1983) - $signed(_zz_21169));
  assign _zz_21169 = ($signed(_zz_21170) * $signed(twiddle_factor_table_75_imag));
  assign _zz_21170 = ($signed(data_mid_76_real) + $signed(data_mid_76_imag));
  assign _zz_21171 = fixTo_2376_dout;
  assign _zz_21172 = ($signed(_zz_1983) + $signed(_zz_21173));
  assign _zz_21173 = ($signed(_zz_21174) * $signed(twiddle_factor_table_75_real));
  assign _zz_21174 = ($signed(data_mid_76_imag) - $signed(data_mid_76_real));
  assign _zz_21175 = fixTo_2377_dout;
  assign _zz_21176 = _zz_21177[31 : 0];
  assign _zz_21177 = _zz_21178;
  assign _zz_21178 = ($signed(_zz_21179) >>> _zz_1984);
  assign _zz_21179 = _zz_21180;
  assign _zz_21180 = ($signed(_zz_21182) - $signed(_zz_1981));
  assign _zz_21181 = ({8'd0,data_mid_12_real} <<< 8);
  assign _zz_21182 = {{8{_zz_21181[23]}}, _zz_21181};
  assign _zz_21183 = fixTo_2378_dout;
  assign _zz_21184 = _zz_21185[31 : 0];
  assign _zz_21185 = _zz_21186;
  assign _zz_21186 = ($signed(_zz_21187) >>> _zz_1984);
  assign _zz_21187 = _zz_21188;
  assign _zz_21188 = ($signed(_zz_21190) - $signed(_zz_1982));
  assign _zz_21189 = ({8'd0,data_mid_12_imag} <<< 8);
  assign _zz_21190 = {{8{_zz_21189[23]}}, _zz_21189};
  assign _zz_21191 = fixTo_2379_dout;
  assign _zz_21192 = _zz_21193[31 : 0];
  assign _zz_21193 = _zz_21194;
  assign _zz_21194 = ($signed(_zz_21195) >>> _zz_1985);
  assign _zz_21195 = _zz_21196;
  assign _zz_21196 = ($signed(_zz_21198) + $signed(_zz_1981));
  assign _zz_21197 = ({8'd0,data_mid_12_real} <<< 8);
  assign _zz_21198 = {{8{_zz_21197[23]}}, _zz_21197};
  assign _zz_21199 = fixTo_2380_dout;
  assign _zz_21200 = _zz_21201[31 : 0];
  assign _zz_21201 = _zz_21202;
  assign _zz_21202 = ($signed(_zz_21203) >>> _zz_1985);
  assign _zz_21203 = _zz_21204;
  assign _zz_21204 = ($signed(_zz_21206) + $signed(_zz_1982));
  assign _zz_21205 = ({8'd0,data_mid_12_imag} <<< 8);
  assign _zz_21206 = {{8{_zz_21205[23]}}, _zz_21205};
  assign _zz_21207 = fixTo_2381_dout;
  assign _zz_21208 = ($signed(twiddle_factor_table_76_real) + $signed(twiddle_factor_table_76_imag));
  assign _zz_21209 = ($signed(_zz_1988) - $signed(_zz_21210));
  assign _zz_21210 = ($signed(_zz_21211) * $signed(twiddle_factor_table_76_imag));
  assign _zz_21211 = ($signed(data_mid_77_real) + $signed(data_mid_77_imag));
  assign _zz_21212 = fixTo_2382_dout;
  assign _zz_21213 = ($signed(_zz_1988) + $signed(_zz_21214));
  assign _zz_21214 = ($signed(_zz_21215) * $signed(twiddle_factor_table_76_real));
  assign _zz_21215 = ($signed(data_mid_77_imag) - $signed(data_mid_77_real));
  assign _zz_21216 = fixTo_2383_dout;
  assign _zz_21217 = _zz_21218[31 : 0];
  assign _zz_21218 = _zz_21219;
  assign _zz_21219 = ($signed(_zz_21220) >>> _zz_1989);
  assign _zz_21220 = _zz_21221;
  assign _zz_21221 = ($signed(_zz_21223) - $signed(_zz_1986));
  assign _zz_21222 = ({8'd0,data_mid_13_real} <<< 8);
  assign _zz_21223 = {{8{_zz_21222[23]}}, _zz_21222};
  assign _zz_21224 = fixTo_2384_dout;
  assign _zz_21225 = _zz_21226[31 : 0];
  assign _zz_21226 = _zz_21227;
  assign _zz_21227 = ($signed(_zz_21228) >>> _zz_1989);
  assign _zz_21228 = _zz_21229;
  assign _zz_21229 = ($signed(_zz_21231) - $signed(_zz_1987));
  assign _zz_21230 = ({8'd0,data_mid_13_imag} <<< 8);
  assign _zz_21231 = {{8{_zz_21230[23]}}, _zz_21230};
  assign _zz_21232 = fixTo_2385_dout;
  assign _zz_21233 = _zz_21234[31 : 0];
  assign _zz_21234 = _zz_21235;
  assign _zz_21235 = ($signed(_zz_21236) >>> _zz_1990);
  assign _zz_21236 = _zz_21237;
  assign _zz_21237 = ($signed(_zz_21239) + $signed(_zz_1986));
  assign _zz_21238 = ({8'd0,data_mid_13_real} <<< 8);
  assign _zz_21239 = {{8{_zz_21238[23]}}, _zz_21238};
  assign _zz_21240 = fixTo_2386_dout;
  assign _zz_21241 = _zz_21242[31 : 0];
  assign _zz_21242 = _zz_21243;
  assign _zz_21243 = ($signed(_zz_21244) >>> _zz_1990);
  assign _zz_21244 = _zz_21245;
  assign _zz_21245 = ($signed(_zz_21247) + $signed(_zz_1987));
  assign _zz_21246 = ({8'd0,data_mid_13_imag} <<< 8);
  assign _zz_21247 = {{8{_zz_21246[23]}}, _zz_21246};
  assign _zz_21248 = fixTo_2387_dout;
  assign _zz_21249 = ($signed(twiddle_factor_table_77_real) + $signed(twiddle_factor_table_77_imag));
  assign _zz_21250 = ($signed(_zz_1993) - $signed(_zz_21251));
  assign _zz_21251 = ($signed(_zz_21252) * $signed(twiddle_factor_table_77_imag));
  assign _zz_21252 = ($signed(data_mid_78_real) + $signed(data_mid_78_imag));
  assign _zz_21253 = fixTo_2388_dout;
  assign _zz_21254 = ($signed(_zz_1993) + $signed(_zz_21255));
  assign _zz_21255 = ($signed(_zz_21256) * $signed(twiddle_factor_table_77_real));
  assign _zz_21256 = ($signed(data_mid_78_imag) - $signed(data_mid_78_real));
  assign _zz_21257 = fixTo_2389_dout;
  assign _zz_21258 = _zz_21259[31 : 0];
  assign _zz_21259 = _zz_21260;
  assign _zz_21260 = ($signed(_zz_21261) >>> _zz_1994);
  assign _zz_21261 = _zz_21262;
  assign _zz_21262 = ($signed(_zz_21264) - $signed(_zz_1991));
  assign _zz_21263 = ({8'd0,data_mid_14_real} <<< 8);
  assign _zz_21264 = {{8{_zz_21263[23]}}, _zz_21263};
  assign _zz_21265 = fixTo_2390_dout;
  assign _zz_21266 = _zz_21267[31 : 0];
  assign _zz_21267 = _zz_21268;
  assign _zz_21268 = ($signed(_zz_21269) >>> _zz_1994);
  assign _zz_21269 = _zz_21270;
  assign _zz_21270 = ($signed(_zz_21272) - $signed(_zz_1992));
  assign _zz_21271 = ({8'd0,data_mid_14_imag} <<< 8);
  assign _zz_21272 = {{8{_zz_21271[23]}}, _zz_21271};
  assign _zz_21273 = fixTo_2391_dout;
  assign _zz_21274 = _zz_21275[31 : 0];
  assign _zz_21275 = _zz_21276;
  assign _zz_21276 = ($signed(_zz_21277) >>> _zz_1995);
  assign _zz_21277 = _zz_21278;
  assign _zz_21278 = ($signed(_zz_21280) + $signed(_zz_1991));
  assign _zz_21279 = ({8'd0,data_mid_14_real} <<< 8);
  assign _zz_21280 = {{8{_zz_21279[23]}}, _zz_21279};
  assign _zz_21281 = fixTo_2392_dout;
  assign _zz_21282 = _zz_21283[31 : 0];
  assign _zz_21283 = _zz_21284;
  assign _zz_21284 = ($signed(_zz_21285) >>> _zz_1995);
  assign _zz_21285 = _zz_21286;
  assign _zz_21286 = ($signed(_zz_21288) + $signed(_zz_1992));
  assign _zz_21287 = ({8'd0,data_mid_14_imag} <<< 8);
  assign _zz_21288 = {{8{_zz_21287[23]}}, _zz_21287};
  assign _zz_21289 = fixTo_2393_dout;
  assign _zz_21290 = ($signed(twiddle_factor_table_78_real) + $signed(twiddle_factor_table_78_imag));
  assign _zz_21291 = ($signed(_zz_1998) - $signed(_zz_21292));
  assign _zz_21292 = ($signed(_zz_21293) * $signed(twiddle_factor_table_78_imag));
  assign _zz_21293 = ($signed(data_mid_79_real) + $signed(data_mid_79_imag));
  assign _zz_21294 = fixTo_2394_dout;
  assign _zz_21295 = ($signed(_zz_1998) + $signed(_zz_21296));
  assign _zz_21296 = ($signed(_zz_21297) * $signed(twiddle_factor_table_78_real));
  assign _zz_21297 = ($signed(data_mid_79_imag) - $signed(data_mid_79_real));
  assign _zz_21298 = fixTo_2395_dout;
  assign _zz_21299 = _zz_21300[31 : 0];
  assign _zz_21300 = _zz_21301;
  assign _zz_21301 = ($signed(_zz_21302) >>> _zz_1999);
  assign _zz_21302 = _zz_21303;
  assign _zz_21303 = ($signed(_zz_21305) - $signed(_zz_1996));
  assign _zz_21304 = ({8'd0,data_mid_15_real} <<< 8);
  assign _zz_21305 = {{8{_zz_21304[23]}}, _zz_21304};
  assign _zz_21306 = fixTo_2396_dout;
  assign _zz_21307 = _zz_21308[31 : 0];
  assign _zz_21308 = _zz_21309;
  assign _zz_21309 = ($signed(_zz_21310) >>> _zz_1999);
  assign _zz_21310 = _zz_21311;
  assign _zz_21311 = ($signed(_zz_21313) - $signed(_zz_1997));
  assign _zz_21312 = ({8'd0,data_mid_15_imag} <<< 8);
  assign _zz_21313 = {{8{_zz_21312[23]}}, _zz_21312};
  assign _zz_21314 = fixTo_2397_dout;
  assign _zz_21315 = _zz_21316[31 : 0];
  assign _zz_21316 = _zz_21317;
  assign _zz_21317 = ($signed(_zz_21318) >>> _zz_2000);
  assign _zz_21318 = _zz_21319;
  assign _zz_21319 = ($signed(_zz_21321) + $signed(_zz_1996));
  assign _zz_21320 = ({8'd0,data_mid_15_real} <<< 8);
  assign _zz_21321 = {{8{_zz_21320[23]}}, _zz_21320};
  assign _zz_21322 = fixTo_2398_dout;
  assign _zz_21323 = _zz_21324[31 : 0];
  assign _zz_21324 = _zz_21325;
  assign _zz_21325 = ($signed(_zz_21326) >>> _zz_2000);
  assign _zz_21326 = _zz_21327;
  assign _zz_21327 = ($signed(_zz_21329) + $signed(_zz_1997));
  assign _zz_21328 = ({8'd0,data_mid_15_imag} <<< 8);
  assign _zz_21329 = {{8{_zz_21328[23]}}, _zz_21328};
  assign _zz_21330 = fixTo_2399_dout;
  assign _zz_21331 = ($signed(twiddle_factor_table_79_real) + $signed(twiddle_factor_table_79_imag));
  assign _zz_21332 = ($signed(_zz_2003) - $signed(_zz_21333));
  assign _zz_21333 = ($signed(_zz_21334) * $signed(twiddle_factor_table_79_imag));
  assign _zz_21334 = ($signed(data_mid_80_real) + $signed(data_mid_80_imag));
  assign _zz_21335 = fixTo_2400_dout;
  assign _zz_21336 = ($signed(_zz_2003) + $signed(_zz_21337));
  assign _zz_21337 = ($signed(_zz_21338) * $signed(twiddle_factor_table_79_real));
  assign _zz_21338 = ($signed(data_mid_80_imag) - $signed(data_mid_80_real));
  assign _zz_21339 = fixTo_2401_dout;
  assign _zz_21340 = _zz_21341[31 : 0];
  assign _zz_21341 = _zz_21342;
  assign _zz_21342 = ($signed(_zz_21343) >>> _zz_2004);
  assign _zz_21343 = _zz_21344;
  assign _zz_21344 = ($signed(_zz_21346) - $signed(_zz_2001));
  assign _zz_21345 = ({8'd0,data_mid_16_real} <<< 8);
  assign _zz_21346 = {{8{_zz_21345[23]}}, _zz_21345};
  assign _zz_21347 = fixTo_2402_dout;
  assign _zz_21348 = _zz_21349[31 : 0];
  assign _zz_21349 = _zz_21350;
  assign _zz_21350 = ($signed(_zz_21351) >>> _zz_2004);
  assign _zz_21351 = _zz_21352;
  assign _zz_21352 = ($signed(_zz_21354) - $signed(_zz_2002));
  assign _zz_21353 = ({8'd0,data_mid_16_imag} <<< 8);
  assign _zz_21354 = {{8{_zz_21353[23]}}, _zz_21353};
  assign _zz_21355 = fixTo_2403_dout;
  assign _zz_21356 = _zz_21357[31 : 0];
  assign _zz_21357 = _zz_21358;
  assign _zz_21358 = ($signed(_zz_21359) >>> _zz_2005);
  assign _zz_21359 = _zz_21360;
  assign _zz_21360 = ($signed(_zz_21362) + $signed(_zz_2001));
  assign _zz_21361 = ({8'd0,data_mid_16_real} <<< 8);
  assign _zz_21362 = {{8{_zz_21361[23]}}, _zz_21361};
  assign _zz_21363 = fixTo_2404_dout;
  assign _zz_21364 = _zz_21365[31 : 0];
  assign _zz_21365 = _zz_21366;
  assign _zz_21366 = ($signed(_zz_21367) >>> _zz_2005);
  assign _zz_21367 = _zz_21368;
  assign _zz_21368 = ($signed(_zz_21370) + $signed(_zz_2002));
  assign _zz_21369 = ({8'd0,data_mid_16_imag} <<< 8);
  assign _zz_21370 = {{8{_zz_21369[23]}}, _zz_21369};
  assign _zz_21371 = fixTo_2405_dout;
  assign _zz_21372 = ($signed(twiddle_factor_table_80_real) + $signed(twiddle_factor_table_80_imag));
  assign _zz_21373 = ($signed(_zz_2008) - $signed(_zz_21374));
  assign _zz_21374 = ($signed(_zz_21375) * $signed(twiddle_factor_table_80_imag));
  assign _zz_21375 = ($signed(data_mid_81_real) + $signed(data_mid_81_imag));
  assign _zz_21376 = fixTo_2406_dout;
  assign _zz_21377 = ($signed(_zz_2008) + $signed(_zz_21378));
  assign _zz_21378 = ($signed(_zz_21379) * $signed(twiddle_factor_table_80_real));
  assign _zz_21379 = ($signed(data_mid_81_imag) - $signed(data_mid_81_real));
  assign _zz_21380 = fixTo_2407_dout;
  assign _zz_21381 = _zz_21382[31 : 0];
  assign _zz_21382 = _zz_21383;
  assign _zz_21383 = ($signed(_zz_21384) >>> _zz_2009);
  assign _zz_21384 = _zz_21385;
  assign _zz_21385 = ($signed(_zz_21387) - $signed(_zz_2006));
  assign _zz_21386 = ({8'd0,data_mid_17_real} <<< 8);
  assign _zz_21387 = {{8{_zz_21386[23]}}, _zz_21386};
  assign _zz_21388 = fixTo_2408_dout;
  assign _zz_21389 = _zz_21390[31 : 0];
  assign _zz_21390 = _zz_21391;
  assign _zz_21391 = ($signed(_zz_21392) >>> _zz_2009);
  assign _zz_21392 = _zz_21393;
  assign _zz_21393 = ($signed(_zz_21395) - $signed(_zz_2007));
  assign _zz_21394 = ({8'd0,data_mid_17_imag} <<< 8);
  assign _zz_21395 = {{8{_zz_21394[23]}}, _zz_21394};
  assign _zz_21396 = fixTo_2409_dout;
  assign _zz_21397 = _zz_21398[31 : 0];
  assign _zz_21398 = _zz_21399;
  assign _zz_21399 = ($signed(_zz_21400) >>> _zz_2010);
  assign _zz_21400 = _zz_21401;
  assign _zz_21401 = ($signed(_zz_21403) + $signed(_zz_2006));
  assign _zz_21402 = ({8'd0,data_mid_17_real} <<< 8);
  assign _zz_21403 = {{8{_zz_21402[23]}}, _zz_21402};
  assign _zz_21404 = fixTo_2410_dout;
  assign _zz_21405 = _zz_21406[31 : 0];
  assign _zz_21406 = _zz_21407;
  assign _zz_21407 = ($signed(_zz_21408) >>> _zz_2010);
  assign _zz_21408 = _zz_21409;
  assign _zz_21409 = ($signed(_zz_21411) + $signed(_zz_2007));
  assign _zz_21410 = ({8'd0,data_mid_17_imag} <<< 8);
  assign _zz_21411 = {{8{_zz_21410[23]}}, _zz_21410};
  assign _zz_21412 = fixTo_2411_dout;
  assign _zz_21413 = ($signed(twiddle_factor_table_81_real) + $signed(twiddle_factor_table_81_imag));
  assign _zz_21414 = ($signed(_zz_2013) - $signed(_zz_21415));
  assign _zz_21415 = ($signed(_zz_21416) * $signed(twiddle_factor_table_81_imag));
  assign _zz_21416 = ($signed(data_mid_82_real) + $signed(data_mid_82_imag));
  assign _zz_21417 = fixTo_2412_dout;
  assign _zz_21418 = ($signed(_zz_2013) + $signed(_zz_21419));
  assign _zz_21419 = ($signed(_zz_21420) * $signed(twiddle_factor_table_81_real));
  assign _zz_21420 = ($signed(data_mid_82_imag) - $signed(data_mid_82_real));
  assign _zz_21421 = fixTo_2413_dout;
  assign _zz_21422 = _zz_21423[31 : 0];
  assign _zz_21423 = _zz_21424;
  assign _zz_21424 = ($signed(_zz_21425) >>> _zz_2014);
  assign _zz_21425 = _zz_21426;
  assign _zz_21426 = ($signed(_zz_21428) - $signed(_zz_2011));
  assign _zz_21427 = ({8'd0,data_mid_18_real} <<< 8);
  assign _zz_21428 = {{8{_zz_21427[23]}}, _zz_21427};
  assign _zz_21429 = fixTo_2414_dout;
  assign _zz_21430 = _zz_21431[31 : 0];
  assign _zz_21431 = _zz_21432;
  assign _zz_21432 = ($signed(_zz_21433) >>> _zz_2014);
  assign _zz_21433 = _zz_21434;
  assign _zz_21434 = ($signed(_zz_21436) - $signed(_zz_2012));
  assign _zz_21435 = ({8'd0,data_mid_18_imag} <<< 8);
  assign _zz_21436 = {{8{_zz_21435[23]}}, _zz_21435};
  assign _zz_21437 = fixTo_2415_dout;
  assign _zz_21438 = _zz_21439[31 : 0];
  assign _zz_21439 = _zz_21440;
  assign _zz_21440 = ($signed(_zz_21441) >>> _zz_2015);
  assign _zz_21441 = _zz_21442;
  assign _zz_21442 = ($signed(_zz_21444) + $signed(_zz_2011));
  assign _zz_21443 = ({8'd0,data_mid_18_real} <<< 8);
  assign _zz_21444 = {{8{_zz_21443[23]}}, _zz_21443};
  assign _zz_21445 = fixTo_2416_dout;
  assign _zz_21446 = _zz_21447[31 : 0];
  assign _zz_21447 = _zz_21448;
  assign _zz_21448 = ($signed(_zz_21449) >>> _zz_2015);
  assign _zz_21449 = _zz_21450;
  assign _zz_21450 = ($signed(_zz_21452) + $signed(_zz_2012));
  assign _zz_21451 = ({8'd0,data_mid_18_imag} <<< 8);
  assign _zz_21452 = {{8{_zz_21451[23]}}, _zz_21451};
  assign _zz_21453 = fixTo_2417_dout;
  assign _zz_21454 = ($signed(twiddle_factor_table_82_real) + $signed(twiddle_factor_table_82_imag));
  assign _zz_21455 = ($signed(_zz_2018) - $signed(_zz_21456));
  assign _zz_21456 = ($signed(_zz_21457) * $signed(twiddle_factor_table_82_imag));
  assign _zz_21457 = ($signed(data_mid_83_real) + $signed(data_mid_83_imag));
  assign _zz_21458 = fixTo_2418_dout;
  assign _zz_21459 = ($signed(_zz_2018) + $signed(_zz_21460));
  assign _zz_21460 = ($signed(_zz_21461) * $signed(twiddle_factor_table_82_real));
  assign _zz_21461 = ($signed(data_mid_83_imag) - $signed(data_mid_83_real));
  assign _zz_21462 = fixTo_2419_dout;
  assign _zz_21463 = _zz_21464[31 : 0];
  assign _zz_21464 = _zz_21465;
  assign _zz_21465 = ($signed(_zz_21466) >>> _zz_2019);
  assign _zz_21466 = _zz_21467;
  assign _zz_21467 = ($signed(_zz_21469) - $signed(_zz_2016));
  assign _zz_21468 = ({8'd0,data_mid_19_real} <<< 8);
  assign _zz_21469 = {{8{_zz_21468[23]}}, _zz_21468};
  assign _zz_21470 = fixTo_2420_dout;
  assign _zz_21471 = _zz_21472[31 : 0];
  assign _zz_21472 = _zz_21473;
  assign _zz_21473 = ($signed(_zz_21474) >>> _zz_2019);
  assign _zz_21474 = _zz_21475;
  assign _zz_21475 = ($signed(_zz_21477) - $signed(_zz_2017));
  assign _zz_21476 = ({8'd0,data_mid_19_imag} <<< 8);
  assign _zz_21477 = {{8{_zz_21476[23]}}, _zz_21476};
  assign _zz_21478 = fixTo_2421_dout;
  assign _zz_21479 = _zz_21480[31 : 0];
  assign _zz_21480 = _zz_21481;
  assign _zz_21481 = ($signed(_zz_21482) >>> _zz_2020);
  assign _zz_21482 = _zz_21483;
  assign _zz_21483 = ($signed(_zz_21485) + $signed(_zz_2016));
  assign _zz_21484 = ({8'd0,data_mid_19_real} <<< 8);
  assign _zz_21485 = {{8{_zz_21484[23]}}, _zz_21484};
  assign _zz_21486 = fixTo_2422_dout;
  assign _zz_21487 = _zz_21488[31 : 0];
  assign _zz_21488 = _zz_21489;
  assign _zz_21489 = ($signed(_zz_21490) >>> _zz_2020);
  assign _zz_21490 = _zz_21491;
  assign _zz_21491 = ($signed(_zz_21493) + $signed(_zz_2017));
  assign _zz_21492 = ({8'd0,data_mid_19_imag} <<< 8);
  assign _zz_21493 = {{8{_zz_21492[23]}}, _zz_21492};
  assign _zz_21494 = fixTo_2423_dout;
  assign _zz_21495 = ($signed(twiddle_factor_table_83_real) + $signed(twiddle_factor_table_83_imag));
  assign _zz_21496 = ($signed(_zz_2023) - $signed(_zz_21497));
  assign _zz_21497 = ($signed(_zz_21498) * $signed(twiddle_factor_table_83_imag));
  assign _zz_21498 = ($signed(data_mid_84_real) + $signed(data_mid_84_imag));
  assign _zz_21499 = fixTo_2424_dout;
  assign _zz_21500 = ($signed(_zz_2023) + $signed(_zz_21501));
  assign _zz_21501 = ($signed(_zz_21502) * $signed(twiddle_factor_table_83_real));
  assign _zz_21502 = ($signed(data_mid_84_imag) - $signed(data_mid_84_real));
  assign _zz_21503 = fixTo_2425_dout;
  assign _zz_21504 = _zz_21505[31 : 0];
  assign _zz_21505 = _zz_21506;
  assign _zz_21506 = ($signed(_zz_21507) >>> _zz_2024);
  assign _zz_21507 = _zz_21508;
  assign _zz_21508 = ($signed(_zz_21510) - $signed(_zz_2021));
  assign _zz_21509 = ({8'd0,data_mid_20_real} <<< 8);
  assign _zz_21510 = {{8{_zz_21509[23]}}, _zz_21509};
  assign _zz_21511 = fixTo_2426_dout;
  assign _zz_21512 = _zz_21513[31 : 0];
  assign _zz_21513 = _zz_21514;
  assign _zz_21514 = ($signed(_zz_21515) >>> _zz_2024);
  assign _zz_21515 = _zz_21516;
  assign _zz_21516 = ($signed(_zz_21518) - $signed(_zz_2022));
  assign _zz_21517 = ({8'd0,data_mid_20_imag} <<< 8);
  assign _zz_21518 = {{8{_zz_21517[23]}}, _zz_21517};
  assign _zz_21519 = fixTo_2427_dout;
  assign _zz_21520 = _zz_21521[31 : 0];
  assign _zz_21521 = _zz_21522;
  assign _zz_21522 = ($signed(_zz_21523) >>> _zz_2025);
  assign _zz_21523 = _zz_21524;
  assign _zz_21524 = ($signed(_zz_21526) + $signed(_zz_2021));
  assign _zz_21525 = ({8'd0,data_mid_20_real} <<< 8);
  assign _zz_21526 = {{8{_zz_21525[23]}}, _zz_21525};
  assign _zz_21527 = fixTo_2428_dout;
  assign _zz_21528 = _zz_21529[31 : 0];
  assign _zz_21529 = _zz_21530;
  assign _zz_21530 = ($signed(_zz_21531) >>> _zz_2025);
  assign _zz_21531 = _zz_21532;
  assign _zz_21532 = ($signed(_zz_21534) + $signed(_zz_2022));
  assign _zz_21533 = ({8'd0,data_mid_20_imag} <<< 8);
  assign _zz_21534 = {{8{_zz_21533[23]}}, _zz_21533};
  assign _zz_21535 = fixTo_2429_dout;
  assign _zz_21536 = ($signed(twiddle_factor_table_84_real) + $signed(twiddle_factor_table_84_imag));
  assign _zz_21537 = ($signed(_zz_2028) - $signed(_zz_21538));
  assign _zz_21538 = ($signed(_zz_21539) * $signed(twiddle_factor_table_84_imag));
  assign _zz_21539 = ($signed(data_mid_85_real) + $signed(data_mid_85_imag));
  assign _zz_21540 = fixTo_2430_dout;
  assign _zz_21541 = ($signed(_zz_2028) + $signed(_zz_21542));
  assign _zz_21542 = ($signed(_zz_21543) * $signed(twiddle_factor_table_84_real));
  assign _zz_21543 = ($signed(data_mid_85_imag) - $signed(data_mid_85_real));
  assign _zz_21544 = fixTo_2431_dout;
  assign _zz_21545 = _zz_21546[31 : 0];
  assign _zz_21546 = _zz_21547;
  assign _zz_21547 = ($signed(_zz_21548) >>> _zz_2029);
  assign _zz_21548 = _zz_21549;
  assign _zz_21549 = ($signed(_zz_21551) - $signed(_zz_2026));
  assign _zz_21550 = ({8'd0,data_mid_21_real} <<< 8);
  assign _zz_21551 = {{8{_zz_21550[23]}}, _zz_21550};
  assign _zz_21552 = fixTo_2432_dout;
  assign _zz_21553 = _zz_21554[31 : 0];
  assign _zz_21554 = _zz_21555;
  assign _zz_21555 = ($signed(_zz_21556) >>> _zz_2029);
  assign _zz_21556 = _zz_21557;
  assign _zz_21557 = ($signed(_zz_21559) - $signed(_zz_2027));
  assign _zz_21558 = ({8'd0,data_mid_21_imag} <<< 8);
  assign _zz_21559 = {{8{_zz_21558[23]}}, _zz_21558};
  assign _zz_21560 = fixTo_2433_dout;
  assign _zz_21561 = _zz_21562[31 : 0];
  assign _zz_21562 = _zz_21563;
  assign _zz_21563 = ($signed(_zz_21564) >>> _zz_2030);
  assign _zz_21564 = _zz_21565;
  assign _zz_21565 = ($signed(_zz_21567) + $signed(_zz_2026));
  assign _zz_21566 = ({8'd0,data_mid_21_real} <<< 8);
  assign _zz_21567 = {{8{_zz_21566[23]}}, _zz_21566};
  assign _zz_21568 = fixTo_2434_dout;
  assign _zz_21569 = _zz_21570[31 : 0];
  assign _zz_21570 = _zz_21571;
  assign _zz_21571 = ($signed(_zz_21572) >>> _zz_2030);
  assign _zz_21572 = _zz_21573;
  assign _zz_21573 = ($signed(_zz_21575) + $signed(_zz_2027));
  assign _zz_21574 = ({8'd0,data_mid_21_imag} <<< 8);
  assign _zz_21575 = {{8{_zz_21574[23]}}, _zz_21574};
  assign _zz_21576 = fixTo_2435_dout;
  assign _zz_21577 = ($signed(twiddle_factor_table_85_real) + $signed(twiddle_factor_table_85_imag));
  assign _zz_21578 = ($signed(_zz_2033) - $signed(_zz_21579));
  assign _zz_21579 = ($signed(_zz_21580) * $signed(twiddle_factor_table_85_imag));
  assign _zz_21580 = ($signed(data_mid_86_real) + $signed(data_mid_86_imag));
  assign _zz_21581 = fixTo_2436_dout;
  assign _zz_21582 = ($signed(_zz_2033) + $signed(_zz_21583));
  assign _zz_21583 = ($signed(_zz_21584) * $signed(twiddle_factor_table_85_real));
  assign _zz_21584 = ($signed(data_mid_86_imag) - $signed(data_mid_86_real));
  assign _zz_21585 = fixTo_2437_dout;
  assign _zz_21586 = _zz_21587[31 : 0];
  assign _zz_21587 = _zz_21588;
  assign _zz_21588 = ($signed(_zz_21589) >>> _zz_2034);
  assign _zz_21589 = _zz_21590;
  assign _zz_21590 = ($signed(_zz_21592) - $signed(_zz_2031));
  assign _zz_21591 = ({8'd0,data_mid_22_real} <<< 8);
  assign _zz_21592 = {{8{_zz_21591[23]}}, _zz_21591};
  assign _zz_21593 = fixTo_2438_dout;
  assign _zz_21594 = _zz_21595[31 : 0];
  assign _zz_21595 = _zz_21596;
  assign _zz_21596 = ($signed(_zz_21597) >>> _zz_2034);
  assign _zz_21597 = _zz_21598;
  assign _zz_21598 = ($signed(_zz_21600) - $signed(_zz_2032));
  assign _zz_21599 = ({8'd0,data_mid_22_imag} <<< 8);
  assign _zz_21600 = {{8{_zz_21599[23]}}, _zz_21599};
  assign _zz_21601 = fixTo_2439_dout;
  assign _zz_21602 = _zz_21603[31 : 0];
  assign _zz_21603 = _zz_21604;
  assign _zz_21604 = ($signed(_zz_21605) >>> _zz_2035);
  assign _zz_21605 = _zz_21606;
  assign _zz_21606 = ($signed(_zz_21608) + $signed(_zz_2031));
  assign _zz_21607 = ({8'd0,data_mid_22_real} <<< 8);
  assign _zz_21608 = {{8{_zz_21607[23]}}, _zz_21607};
  assign _zz_21609 = fixTo_2440_dout;
  assign _zz_21610 = _zz_21611[31 : 0];
  assign _zz_21611 = _zz_21612;
  assign _zz_21612 = ($signed(_zz_21613) >>> _zz_2035);
  assign _zz_21613 = _zz_21614;
  assign _zz_21614 = ($signed(_zz_21616) + $signed(_zz_2032));
  assign _zz_21615 = ({8'd0,data_mid_22_imag} <<< 8);
  assign _zz_21616 = {{8{_zz_21615[23]}}, _zz_21615};
  assign _zz_21617 = fixTo_2441_dout;
  assign _zz_21618 = ($signed(twiddle_factor_table_86_real) + $signed(twiddle_factor_table_86_imag));
  assign _zz_21619 = ($signed(_zz_2038) - $signed(_zz_21620));
  assign _zz_21620 = ($signed(_zz_21621) * $signed(twiddle_factor_table_86_imag));
  assign _zz_21621 = ($signed(data_mid_87_real) + $signed(data_mid_87_imag));
  assign _zz_21622 = fixTo_2442_dout;
  assign _zz_21623 = ($signed(_zz_2038) + $signed(_zz_21624));
  assign _zz_21624 = ($signed(_zz_21625) * $signed(twiddle_factor_table_86_real));
  assign _zz_21625 = ($signed(data_mid_87_imag) - $signed(data_mid_87_real));
  assign _zz_21626 = fixTo_2443_dout;
  assign _zz_21627 = _zz_21628[31 : 0];
  assign _zz_21628 = _zz_21629;
  assign _zz_21629 = ($signed(_zz_21630) >>> _zz_2039);
  assign _zz_21630 = _zz_21631;
  assign _zz_21631 = ($signed(_zz_21633) - $signed(_zz_2036));
  assign _zz_21632 = ({8'd0,data_mid_23_real} <<< 8);
  assign _zz_21633 = {{8{_zz_21632[23]}}, _zz_21632};
  assign _zz_21634 = fixTo_2444_dout;
  assign _zz_21635 = _zz_21636[31 : 0];
  assign _zz_21636 = _zz_21637;
  assign _zz_21637 = ($signed(_zz_21638) >>> _zz_2039);
  assign _zz_21638 = _zz_21639;
  assign _zz_21639 = ($signed(_zz_21641) - $signed(_zz_2037));
  assign _zz_21640 = ({8'd0,data_mid_23_imag} <<< 8);
  assign _zz_21641 = {{8{_zz_21640[23]}}, _zz_21640};
  assign _zz_21642 = fixTo_2445_dout;
  assign _zz_21643 = _zz_21644[31 : 0];
  assign _zz_21644 = _zz_21645;
  assign _zz_21645 = ($signed(_zz_21646) >>> _zz_2040);
  assign _zz_21646 = _zz_21647;
  assign _zz_21647 = ($signed(_zz_21649) + $signed(_zz_2036));
  assign _zz_21648 = ({8'd0,data_mid_23_real} <<< 8);
  assign _zz_21649 = {{8{_zz_21648[23]}}, _zz_21648};
  assign _zz_21650 = fixTo_2446_dout;
  assign _zz_21651 = _zz_21652[31 : 0];
  assign _zz_21652 = _zz_21653;
  assign _zz_21653 = ($signed(_zz_21654) >>> _zz_2040);
  assign _zz_21654 = _zz_21655;
  assign _zz_21655 = ($signed(_zz_21657) + $signed(_zz_2037));
  assign _zz_21656 = ({8'd0,data_mid_23_imag} <<< 8);
  assign _zz_21657 = {{8{_zz_21656[23]}}, _zz_21656};
  assign _zz_21658 = fixTo_2447_dout;
  assign _zz_21659 = ($signed(twiddle_factor_table_87_real) + $signed(twiddle_factor_table_87_imag));
  assign _zz_21660 = ($signed(_zz_2043) - $signed(_zz_21661));
  assign _zz_21661 = ($signed(_zz_21662) * $signed(twiddle_factor_table_87_imag));
  assign _zz_21662 = ($signed(data_mid_88_real) + $signed(data_mid_88_imag));
  assign _zz_21663 = fixTo_2448_dout;
  assign _zz_21664 = ($signed(_zz_2043) + $signed(_zz_21665));
  assign _zz_21665 = ($signed(_zz_21666) * $signed(twiddle_factor_table_87_real));
  assign _zz_21666 = ($signed(data_mid_88_imag) - $signed(data_mid_88_real));
  assign _zz_21667 = fixTo_2449_dout;
  assign _zz_21668 = _zz_21669[31 : 0];
  assign _zz_21669 = _zz_21670;
  assign _zz_21670 = ($signed(_zz_21671) >>> _zz_2044);
  assign _zz_21671 = _zz_21672;
  assign _zz_21672 = ($signed(_zz_21674) - $signed(_zz_2041));
  assign _zz_21673 = ({8'd0,data_mid_24_real} <<< 8);
  assign _zz_21674 = {{8{_zz_21673[23]}}, _zz_21673};
  assign _zz_21675 = fixTo_2450_dout;
  assign _zz_21676 = _zz_21677[31 : 0];
  assign _zz_21677 = _zz_21678;
  assign _zz_21678 = ($signed(_zz_21679) >>> _zz_2044);
  assign _zz_21679 = _zz_21680;
  assign _zz_21680 = ($signed(_zz_21682) - $signed(_zz_2042));
  assign _zz_21681 = ({8'd0,data_mid_24_imag} <<< 8);
  assign _zz_21682 = {{8{_zz_21681[23]}}, _zz_21681};
  assign _zz_21683 = fixTo_2451_dout;
  assign _zz_21684 = _zz_21685[31 : 0];
  assign _zz_21685 = _zz_21686;
  assign _zz_21686 = ($signed(_zz_21687) >>> _zz_2045);
  assign _zz_21687 = _zz_21688;
  assign _zz_21688 = ($signed(_zz_21690) + $signed(_zz_2041));
  assign _zz_21689 = ({8'd0,data_mid_24_real} <<< 8);
  assign _zz_21690 = {{8{_zz_21689[23]}}, _zz_21689};
  assign _zz_21691 = fixTo_2452_dout;
  assign _zz_21692 = _zz_21693[31 : 0];
  assign _zz_21693 = _zz_21694;
  assign _zz_21694 = ($signed(_zz_21695) >>> _zz_2045);
  assign _zz_21695 = _zz_21696;
  assign _zz_21696 = ($signed(_zz_21698) + $signed(_zz_2042));
  assign _zz_21697 = ({8'd0,data_mid_24_imag} <<< 8);
  assign _zz_21698 = {{8{_zz_21697[23]}}, _zz_21697};
  assign _zz_21699 = fixTo_2453_dout;
  assign _zz_21700 = ($signed(twiddle_factor_table_88_real) + $signed(twiddle_factor_table_88_imag));
  assign _zz_21701 = ($signed(_zz_2048) - $signed(_zz_21702));
  assign _zz_21702 = ($signed(_zz_21703) * $signed(twiddle_factor_table_88_imag));
  assign _zz_21703 = ($signed(data_mid_89_real) + $signed(data_mid_89_imag));
  assign _zz_21704 = fixTo_2454_dout;
  assign _zz_21705 = ($signed(_zz_2048) + $signed(_zz_21706));
  assign _zz_21706 = ($signed(_zz_21707) * $signed(twiddle_factor_table_88_real));
  assign _zz_21707 = ($signed(data_mid_89_imag) - $signed(data_mid_89_real));
  assign _zz_21708 = fixTo_2455_dout;
  assign _zz_21709 = _zz_21710[31 : 0];
  assign _zz_21710 = _zz_21711;
  assign _zz_21711 = ($signed(_zz_21712) >>> _zz_2049);
  assign _zz_21712 = _zz_21713;
  assign _zz_21713 = ($signed(_zz_21715) - $signed(_zz_2046));
  assign _zz_21714 = ({8'd0,data_mid_25_real} <<< 8);
  assign _zz_21715 = {{8{_zz_21714[23]}}, _zz_21714};
  assign _zz_21716 = fixTo_2456_dout;
  assign _zz_21717 = _zz_21718[31 : 0];
  assign _zz_21718 = _zz_21719;
  assign _zz_21719 = ($signed(_zz_21720) >>> _zz_2049);
  assign _zz_21720 = _zz_21721;
  assign _zz_21721 = ($signed(_zz_21723) - $signed(_zz_2047));
  assign _zz_21722 = ({8'd0,data_mid_25_imag} <<< 8);
  assign _zz_21723 = {{8{_zz_21722[23]}}, _zz_21722};
  assign _zz_21724 = fixTo_2457_dout;
  assign _zz_21725 = _zz_21726[31 : 0];
  assign _zz_21726 = _zz_21727;
  assign _zz_21727 = ($signed(_zz_21728) >>> _zz_2050);
  assign _zz_21728 = _zz_21729;
  assign _zz_21729 = ($signed(_zz_21731) + $signed(_zz_2046));
  assign _zz_21730 = ({8'd0,data_mid_25_real} <<< 8);
  assign _zz_21731 = {{8{_zz_21730[23]}}, _zz_21730};
  assign _zz_21732 = fixTo_2458_dout;
  assign _zz_21733 = _zz_21734[31 : 0];
  assign _zz_21734 = _zz_21735;
  assign _zz_21735 = ($signed(_zz_21736) >>> _zz_2050);
  assign _zz_21736 = _zz_21737;
  assign _zz_21737 = ($signed(_zz_21739) + $signed(_zz_2047));
  assign _zz_21738 = ({8'd0,data_mid_25_imag} <<< 8);
  assign _zz_21739 = {{8{_zz_21738[23]}}, _zz_21738};
  assign _zz_21740 = fixTo_2459_dout;
  assign _zz_21741 = ($signed(twiddle_factor_table_89_real) + $signed(twiddle_factor_table_89_imag));
  assign _zz_21742 = ($signed(_zz_2053) - $signed(_zz_21743));
  assign _zz_21743 = ($signed(_zz_21744) * $signed(twiddle_factor_table_89_imag));
  assign _zz_21744 = ($signed(data_mid_90_real) + $signed(data_mid_90_imag));
  assign _zz_21745 = fixTo_2460_dout;
  assign _zz_21746 = ($signed(_zz_2053) + $signed(_zz_21747));
  assign _zz_21747 = ($signed(_zz_21748) * $signed(twiddle_factor_table_89_real));
  assign _zz_21748 = ($signed(data_mid_90_imag) - $signed(data_mid_90_real));
  assign _zz_21749 = fixTo_2461_dout;
  assign _zz_21750 = _zz_21751[31 : 0];
  assign _zz_21751 = _zz_21752;
  assign _zz_21752 = ($signed(_zz_21753) >>> _zz_2054);
  assign _zz_21753 = _zz_21754;
  assign _zz_21754 = ($signed(_zz_21756) - $signed(_zz_2051));
  assign _zz_21755 = ({8'd0,data_mid_26_real} <<< 8);
  assign _zz_21756 = {{8{_zz_21755[23]}}, _zz_21755};
  assign _zz_21757 = fixTo_2462_dout;
  assign _zz_21758 = _zz_21759[31 : 0];
  assign _zz_21759 = _zz_21760;
  assign _zz_21760 = ($signed(_zz_21761) >>> _zz_2054);
  assign _zz_21761 = _zz_21762;
  assign _zz_21762 = ($signed(_zz_21764) - $signed(_zz_2052));
  assign _zz_21763 = ({8'd0,data_mid_26_imag} <<< 8);
  assign _zz_21764 = {{8{_zz_21763[23]}}, _zz_21763};
  assign _zz_21765 = fixTo_2463_dout;
  assign _zz_21766 = _zz_21767[31 : 0];
  assign _zz_21767 = _zz_21768;
  assign _zz_21768 = ($signed(_zz_21769) >>> _zz_2055);
  assign _zz_21769 = _zz_21770;
  assign _zz_21770 = ($signed(_zz_21772) + $signed(_zz_2051));
  assign _zz_21771 = ({8'd0,data_mid_26_real} <<< 8);
  assign _zz_21772 = {{8{_zz_21771[23]}}, _zz_21771};
  assign _zz_21773 = fixTo_2464_dout;
  assign _zz_21774 = _zz_21775[31 : 0];
  assign _zz_21775 = _zz_21776;
  assign _zz_21776 = ($signed(_zz_21777) >>> _zz_2055);
  assign _zz_21777 = _zz_21778;
  assign _zz_21778 = ($signed(_zz_21780) + $signed(_zz_2052));
  assign _zz_21779 = ({8'd0,data_mid_26_imag} <<< 8);
  assign _zz_21780 = {{8{_zz_21779[23]}}, _zz_21779};
  assign _zz_21781 = fixTo_2465_dout;
  assign _zz_21782 = ($signed(twiddle_factor_table_90_real) + $signed(twiddle_factor_table_90_imag));
  assign _zz_21783 = ($signed(_zz_2058) - $signed(_zz_21784));
  assign _zz_21784 = ($signed(_zz_21785) * $signed(twiddle_factor_table_90_imag));
  assign _zz_21785 = ($signed(data_mid_91_real) + $signed(data_mid_91_imag));
  assign _zz_21786 = fixTo_2466_dout;
  assign _zz_21787 = ($signed(_zz_2058) + $signed(_zz_21788));
  assign _zz_21788 = ($signed(_zz_21789) * $signed(twiddle_factor_table_90_real));
  assign _zz_21789 = ($signed(data_mid_91_imag) - $signed(data_mid_91_real));
  assign _zz_21790 = fixTo_2467_dout;
  assign _zz_21791 = _zz_21792[31 : 0];
  assign _zz_21792 = _zz_21793;
  assign _zz_21793 = ($signed(_zz_21794) >>> _zz_2059);
  assign _zz_21794 = _zz_21795;
  assign _zz_21795 = ($signed(_zz_21797) - $signed(_zz_2056));
  assign _zz_21796 = ({8'd0,data_mid_27_real} <<< 8);
  assign _zz_21797 = {{8{_zz_21796[23]}}, _zz_21796};
  assign _zz_21798 = fixTo_2468_dout;
  assign _zz_21799 = _zz_21800[31 : 0];
  assign _zz_21800 = _zz_21801;
  assign _zz_21801 = ($signed(_zz_21802) >>> _zz_2059);
  assign _zz_21802 = _zz_21803;
  assign _zz_21803 = ($signed(_zz_21805) - $signed(_zz_2057));
  assign _zz_21804 = ({8'd0,data_mid_27_imag} <<< 8);
  assign _zz_21805 = {{8{_zz_21804[23]}}, _zz_21804};
  assign _zz_21806 = fixTo_2469_dout;
  assign _zz_21807 = _zz_21808[31 : 0];
  assign _zz_21808 = _zz_21809;
  assign _zz_21809 = ($signed(_zz_21810) >>> _zz_2060);
  assign _zz_21810 = _zz_21811;
  assign _zz_21811 = ($signed(_zz_21813) + $signed(_zz_2056));
  assign _zz_21812 = ({8'd0,data_mid_27_real} <<< 8);
  assign _zz_21813 = {{8{_zz_21812[23]}}, _zz_21812};
  assign _zz_21814 = fixTo_2470_dout;
  assign _zz_21815 = _zz_21816[31 : 0];
  assign _zz_21816 = _zz_21817;
  assign _zz_21817 = ($signed(_zz_21818) >>> _zz_2060);
  assign _zz_21818 = _zz_21819;
  assign _zz_21819 = ($signed(_zz_21821) + $signed(_zz_2057));
  assign _zz_21820 = ({8'd0,data_mid_27_imag} <<< 8);
  assign _zz_21821 = {{8{_zz_21820[23]}}, _zz_21820};
  assign _zz_21822 = fixTo_2471_dout;
  assign _zz_21823 = ($signed(twiddle_factor_table_91_real) + $signed(twiddle_factor_table_91_imag));
  assign _zz_21824 = ($signed(_zz_2063) - $signed(_zz_21825));
  assign _zz_21825 = ($signed(_zz_21826) * $signed(twiddle_factor_table_91_imag));
  assign _zz_21826 = ($signed(data_mid_92_real) + $signed(data_mid_92_imag));
  assign _zz_21827 = fixTo_2472_dout;
  assign _zz_21828 = ($signed(_zz_2063) + $signed(_zz_21829));
  assign _zz_21829 = ($signed(_zz_21830) * $signed(twiddle_factor_table_91_real));
  assign _zz_21830 = ($signed(data_mid_92_imag) - $signed(data_mid_92_real));
  assign _zz_21831 = fixTo_2473_dout;
  assign _zz_21832 = _zz_21833[31 : 0];
  assign _zz_21833 = _zz_21834;
  assign _zz_21834 = ($signed(_zz_21835) >>> _zz_2064);
  assign _zz_21835 = _zz_21836;
  assign _zz_21836 = ($signed(_zz_21838) - $signed(_zz_2061));
  assign _zz_21837 = ({8'd0,data_mid_28_real} <<< 8);
  assign _zz_21838 = {{8{_zz_21837[23]}}, _zz_21837};
  assign _zz_21839 = fixTo_2474_dout;
  assign _zz_21840 = _zz_21841[31 : 0];
  assign _zz_21841 = _zz_21842;
  assign _zz_21842 = ($signed(_zz_21843) >>> _zz_2064);
  assign _zz_21843 = _zz_21844;
  assign _zz_21844 = ($signed(_zz_21846) - $signed(_zz_2062));
  assign _zz_21845 = ({8'd0,data_mid_28_imag} <<< 8);
  assign _zz_21846 = {{8{_zz_21845[23]}}, _zz_21845};
  assign _zz_21847 = fixTo_2475_dout;
  assign _zz_21848 = _zz_21849[31 : 0];
  assign _zz_21849 = _zz_21850;
  assign _zz_21850 = ($signed(_zz_21851) >>> _zz_2065);
  assign _zz_21851 = _zz_21852;
  assign _zz_21852 = ($signed(_zz_21854) + $signed(_zz_2061));
  assign _zz_21853 = ({8'd0,data_mid_28_real} <<< 8);
  assign _zz_21854 = {{8{_zz_21853[23]}}, _zz_21853};
  assign _zz_21855 = fixTo_2476_dout;
  assign _zz_21856 = _zz_21857[31 : 0];
  assign _zz_21857 = _zz_21858;
  assign _zz_21858 = ($signed(_zz_21859) >>> _zz_2065);
  assign _zz_21859 = _zz_21860;
  assign _zz_21860 = ($signed(_zz_21862) + $signed(_zz_2062));
  assign _zz_21861 = ({8'd0,data_mid_28_imag} <<< 8);
  assign _zz_21862 = {{8{_zz_21861[23]}}, _zz_21861};
  assign _zz_21863 = fixTo_2477_dout;
  assign _zz_21864 = ($signed(twiddle_factor_table_92_real) + $signed(twiddle_factor_table_92_imag));
  assign _zz_21865 = ($signed(_zz_2068) - $signed(_zz_21866));
  assign _zz_21866 = ($signed(_zz_21867) * $signed(twiddle_factor_table_92_imag));
  assign _zz_21867 = ($signed(data_mid_93_real) + $signed(data_mid_93_imag));
  assign _zz_21868 = fixTo_2478_dout;
  assign _zz_21869 = ($signed(_zz_2068) + $signed(_zz_21870));
  assign _zz_21870 = ($signed(_zz_21871) * $signed(twiddle_factor_table_92_real));
  assign _zz_21871 = ($signed(data_mid_93_imag) - $signed(data_mid_93_real));
  assign _zz_21872 = fixTo_2479_dout;
  assign _zz_21873 = _zz_21874[31 : 0];
  assign _zz_21874 = _zz_21875;
  assign _zz_21875 = ($signed(_zz_21876) >>> _zz_2069);
  assign _zz_21876 = _zz_21877;
  assign _zz_21877 = ($signed(_zz_21879) - $signed(_zz_2066));
  assign _zz_21878 = ({8'd0,data_mid_29_real} <<< 8);
  assign _zz_21879 = {{8{_zz_21878[23]}}, _zz_21878};
  assign _zz_21880 = fixTo_2480_dout;
  assign _zz_21881 = _zz_21882[31 : 0];
  assign _zz_21882 = _zz_21883;
  assign _zz_21883 = ($signed(_zz_21884) >>> _zz_2069);
  assign _zz_21884 = _zz_21885;
  assign _zz_21885 = ($signed(_zz_21887) - $signed(_zz_2067));
  assign _zz_21886 = ({8'd0,data_mid_29_imag} <<< 8);
  assign _zz_21887 = {{8{_zz_21886[23]}}, _zz_21886};
  assign _zz_21888 = fixTo_2481_dout;
  assign _zz_21889 = _zz_21890[31 : 0];
  assign _zz_21890 = _zz_21891;
  assign _zz_21891 = ($signed(_zz_21892) >>> _zz_2070);
  assign _zz_21892 = _zz_21893;
  assign _zz_21893 = ($signed(_zz_21895) + $signed(_zz_2066));
  assign _zz_21894 = ({8'd0,data_mid_29_real} <<< 8);
  assign _zz_21895 = {{8{_zz_21894[23]}}, _zz_21894};
  assign _zz_21896 = fixTo_2482_dout;
  assign _zz_21897 = _zz_21898[31 : 0];
  assign _zz_21898 = _zz_21899;
  assign _zz_21899 = ($signed(_zz_21900) >>> _zz_2070);
  assign _zz_21900 = _zz_21901;
  assign _zz_21901 = ($signed(_zz_21903) + $signed(_zz_2067));
  assign _zz_21902 = ({8'd0,data_mid_29_imag} <<< 8);
  assign _zz_21903 = {{8{_zz_21902[23]}}, _zz_21902};
  assign _zz_21904 = fixTo_2483_dout;
  assign _zz_21905 = ($signed(twiddle_factor_table_93_real) + $signed(twiddle_factor_table_93_imag));
  assign _zz_21906 = ($signed(_zz_2073) - $signed(_zz_21907));
  assign _zz_21907 = ($signed(_zz_21908) * $signed(twiddle_factor_table_93_imag));
  assign _zz_21908 = ($signed(data_mid_94_real) + $signed(data_mid_94_imag));
  assign _zz_21909 = fixTo_2484_dout;
  assign _zz_21910 = ($signed(_zz_2073) + $signed(_zz_21911));
  assign _zz_21911 = ($signed(_zz_21912) * $signed(twiddle_factor_table_93_real));
  assign _zz_21912 = ($signed(data_mid_94_imag) - $signed(data_mid_94_real));
  assign _zz_21913 = fixTo_2485_dout;
  assign _zz_21914 = _zz_21915[31 : 0];
  assign _zz_21915 = _zz_21916;
  assign _zz_21916 = ($signed(_zz_21917) >>> _zz_2074);
  assign _zz_21917 = _zz_21918;
  assign _zz_21918 = ($signed(_zz_21920) - $signed(_zz_2071));
  assign _zz_21919 = ({8'd0,data_mid_30_real} <<< 8);
  assign _zz_21920 = {{8{_zz_21919[23]}}, _zz_21919};
  assign _zz_21921 = fixTo_2486_dout;
  assign _zz_21922 = _zz_21923[31 : 0];
  assign _zz_21923 = _zz_21924;
  assign _zz_21924 = ($signed(_zz_21925) >>> _zz_2074);
  assign _zz_21925 = _zz_21926;
  assign _zz_21926 = ($signed(_zz_21928) - $signed(_zz_2072));
  assign _zz_21927 = ({8'd0,data_mid_30_imag} <<< 8);
  assign _zz_21928 = {{8{_zz_21927[23]}}, _zz_21927};
  assign _zz_21929 = fixTo_2487_dout;
  assign _zz_21930 = _zz_21931[31 : 0];
  assign _zz_21931 = _zz_21932;
  assign _zz_21932 = ($signed(_zz_21933) >>> _zz_2075);
  assign _zz_21933 = _zz_21934;
  assign _zz_21934 = ($signed(_zz_21936) + $signed(_zz_2071));
  assign _zz_21935 = ({8'd0,data_mid_30_real} <<< 8);
  assign _zz_21936 = {{8{_zz_21935[23]}}, _zz_21935};
  assign _zz_21937 = fixTo_2488_dout;
  assign _zz_21938 = _zz_21939[31 : 0];
  assign _zz_21939 = _zz_21940;
  assign _zz_21940 = ($signed(_zz_21941) >>> _zz_2075);
  assign _zz_21941 = _zz_21942;
  assign _zz_21942 = ($signed(_zz_21944) + $signed(_zz_2072));
  assign _zz_21943 = ({8'd0,data_mid_30_imag} <<< 8);
  assign _zz_21944 = {{8{_zz_21943[23]}}, _zz_21943};
  assign _zz_21945 = fixTo_2489_dout;
  assign _zz_21946 = ($signed(twiddle_factor_table_94_real) + $signed(twiddle_factor_table_94_imag));
  assign _zz_21947 = ($signed(_zz_2078) - $signed(_zz_21948));
  assign _zz_21948 = ($signed(_zz_21949) * $signed(twiddle_factor_table_94_imag));
  assign _zz_21949 = ($signed(data_mid_95_real) + $signed(data_mid_95_imag));
  assign _zz_21950 = fixTo_2490_dout;
  assign _zz_21951 = ($signed(_zz_2078) + $signed(_zz_21952));
  assign _zz_21952 = ($signed(_zz_21953) * $signed(twiddle_factor_table_94_real));
  assign _zz_21953 = ($signed(data_mid_95_imag) - $signed(data_mid_95_real));
  assign _zz_21954 = fixTo_2491_dout;
  assign _zz_21955 = _zz_21956[31 : 0];
  assign _zz_21956 = _zz_21957;
  assign _zz_21957 = ($signed(_zz_21958) >>> _zz_2079);
  assign _zz_21958 = _zz_21959;
  assign _zz_21959 = ($signed(_zz_21961) - $signed(_zz_2076));
  assign _zz_21960 = ({8'd0,data_mid_31_real} <<< 8);
  assign _zz_21961 = {{8{_zz_21960[23]}}, _zz_21960};
  assign _zz_21962 = fixTo_2492_dout;
  assign _zz_21963 = _zz_21964[31 : 0];
  assign _zz_21964 = _zz_21965;
  assign _zz_21965 = ($signed(_zz_21966) >>> _zz_2079);
  assign _zz_21966 = _zz_21967;
  assign _zz_21967 = ($signed(_zz_21969) - $signed(_zz_2077));
  assign _zz_21968 = ({8'd0,data_mid_31_imag} <<< 8);
  assign _zz_21969 = {{8{_zz_21968[23]}}, _zz_21968};
  assign _zz_21970 = fixTo_2493_dout;
  assign _zz_21971 = _zz_21972[31 : 0];
  assign _zz_21972 = _zz_21973;
  assign _zz_21973 = ($signed(_zz_21974) >>> _zz_2080);
  assign _zz_21974 = _zz_21975;
  assign _zz_21975 = ($signed(_zz_21977) + $signed(_zz_2076));
  assign _zz_21976 = ({8'd0,data_mid_31_real} <<< 8);
  assign _zz_21977 = {{8{_zz_21976[23]}}, _zz_21976};
  assign _zz_21978 = fixTo_2494_dout;
  assign _zz_21979 = _zz_21980[31 : 0];
  assign _zz_21980 = _zz_21981;
  assign _zz_21981 = ($signed(_zz_21982) >>> _zz_2080);
  assign _zz_21982 = _zz_21983;
  assign _zz_21983 = ($signed(_zz_21985) + $signed(_zz_2077));
  assign _zz_21984 = ({8'd0,data_mid_31_imag} <<< 8);
  assign _zz_21985 = {{8{_zz_21984[23]}}, _zz_21984};
  assign _zz_21986 = fixTo_2495_dout;
  assign _zz_21987 = ($signed(twiddle_factor_table_95_real) + $signed(twiddle_factor_table_95_imag));
  assign _zz_21988 = ($signed(_zz_2083) - $signed(_zz_21989));
  assign _zz_21989 = ($signed(_zz_21990) * $signed(twiddle_factor_table_95_imag));
  assign _zz_21990 = ($signed(data_mid_96_real) + $signed(data_mid_96_imag));
  assign _zz_21991 = fixTo_2496_dout;
  assign _zz_21992 = ($signed(_zz_2083) + $signed(_zz_21993));
  assign _zz_21993 = ($signed(_zz_21994) * $signed(twiddle_factor_table_95_real));
  assign _zz_21994 = ($signed(data_mid_96_imag) - $signed(data_mid_96_real));
  assign _zz_21995 = fixTo_2497_dout;
  assign _zz_21996 = _zz_21997[31 : 0];
  assign _zz_21997 = _zz_21998;
  assign _zz_21998 = ($signed(_zz_21999) >>> _zz_2084);
  assign _zz_21999 = _zz_22000;
  assign _zz_22000 = ($signed(_zz_22002) - $signed(_zz_2081));
  assign _zz_22001 = ({8'd0,data_mid_32_real} <<< 8);
  assign _zz_22002 = {{8{_zz_22001[23]}}, _zz_22001};
  assign _zz_22003 = fixTo_2498_dout;
  assign _zz_22004 = _zz_22005[31 : 0];
  assign _zz_22005 = _zz_22006;
  assign _zz_22006 = ($signed(_zz_22007) >>> _zz_2084);
  assign _zz_22007 = _zz_22008;
  assign _zz_22008 = ($signed(_zz_22010) - $signed(_zz_2082));
  assign _zz_22009 = ({8'd0,data_mid_32_imag} <<< 8);
  assign _zz_22010 = {{8{_zz_22009[23]}}, _zz_22009};
  assign _zz_22011 = fixTo_2499_dout;
  assign _zz_22012 = _zz_22013[31 : 0];
  assign _zz_22013 = _zz_22014;
  assign _zz_22014 = ($signed(_zz_22015) >>> _zz_2085);
  assign _zz_22015 = _zz_22016;
  assign _zz_22016 = ($signed(_zz_22018) + $signed(_zz_2081));
  assign _zz_22017 = ({8'd0,data_mid_32_real} <<< 8);
  assign _zz_22018 = {{8{_zz_22017[23]}}, _zz_22017};
  assign _zz_22019 = fixTo_2500_dout;
  assign _zz_22020 = _zz_22021[31 : 0];
  assign _zz_22021 = _zz_22022;
  assign _zz_22022 = ($signed(_zz_22023) >>> _zz_2085);
  assign _zz_22023 = _zz_22024;
  assign _zz_22024 = ($signed(_zz_22026) + $signed(_zz_2082));
  assign _zz_22025 = ({8'd0,data_mid_32_imag} <<< 8);
  assign _zz_22026 = {{8{_zz_22025[23]}}, _zz_22025};
  assign _zz_22027 = fixTo_2501_dout;
  assign _zz_22028 = ($signed(twiddle_factor_table_96_real) + $signed(twiddle_factor_table_96_imag));
  assign _zz_22029 = ($signed(_zz_2088) - $signed(_zz_22030));
  assign _zz_22030 = ($signed(_zz_22031) * $signed(twiddle_factor_table_96_imag));
  assign _zz_22031 = ($signed(data_mid_97_real) + $signed(data_mid_97_imag));
  assign _zz_22032 = fixTo_2502_dout;
  assign _zz_22033 = ($signed(_zz_2088) + $signed(_zz_22034));
  assign _zz_22034 = ($signed(_zz_22035) * $signed(twiddle_factor_table_96_real));
  assign _zz_22035 = ($signed(data_mid_97_imag) - $signed(data_mid_97_real));
  assign _zz_22036 = fixTo_2503_dout;
  assign _zz_22037 = _zz_22038[31 : 0];
  assign _zz_22038 = _zz_22039;
  assign _zz_22039 = ($signed(_zz_22040) >>> _zz_2089);
  assign _zz_22040 = _zz_22041;
  assign _zz_22041 = ($signed(_zz_22043) - $signed(_zz_2086));
  assign _zz_22042 = ({8'd0,data_mid_33_real} <<< 8);
  assign _zz_22043 = {{8{_zz_22042[23]}}, _zz_22042};
  assign _zz_22044 = fixTo_2504_dout;
  assign _zz_22045 = _zz_22046[31 : 0];
  assign _zz_22046 = _zz_22047;
  assign _zz_22047 = ($signed(_zz_22048) >>> _zz_2089);
  assign _zz_22048 = _zz_22049;
  assign _zz_22049 = ($signed(_zz_22051) - $signed(_zz_2087));
  assign _zz_22050 = ({8'd0,data_mid_33_imag} <<< 8);
  assign _zz_22051 = {{8{_zz_22050[23]}}, _zz_22050};
  assign _zz_22052 = fixTo_2505_dout;
  assign _zz_22053 = _zz_22054[31 : 0];
  assign _zz_22054 = _zz_22055;
  assign _zz_22055 = ($signed(_zz_22056) >>> _zz_2090);
  assign _zz_22056 = _zz_22057;
  assign _zz_22057 = ($signed(_zz_22059) + $signed(_zz_2086));
  assign _zz_22058 = ({8'd0,data_mid_33_real} <<< 8);
  assign _zz_22059 = {{8{_zz_22058[23]}}, _zz_22058};
  assign _zz_22060 = fixTo_2506_dout;
  assign _zz_22061 = _zz_22062[31 : 0];
  assign _zz_22062 = _zz_22063;
  assign _zz_22063 = ($signed(_zz_22064) >>> _zz_2090);
  assign _zz_22064 = _zz_22065;
  assign _zz_22065 = ($signed(_zz_22067) + $signed(_zz_2087));
  assign _zz_22066 = ({8'd0,data_mid_33_imag} <<< 8);
  assign _zz_22067 = {{8{_zz_22066[23]}}, _zz_22066};
  assign _zz_22068 = fixTo_2507_dout;
  assign _zz_22069 = ($signed(twiddle_factor_table_97_real) + $signed(twiddle_factor_table_97_imag));
  assign _zz_22070 = ($signed(_zz_2093) - $signed(_zz_22071));
  assign _zz_22071 = ($signed(_zz_22072) * $signed(twiddle_factor_table_97_imag));
  assign _zz_22072 = ($signed(data_mid_98_real) + $signed(data_mid_98_imag));
  assign _zz_22073 = fixTo_2508_dout;
  assign _zz_22074 = ($signed(_zz_2093) + $signed(_zz_22075));
  assign _zz_22075 = ($signed(_zz_22076) * $signed(twiddle_factor_table_97_real));
  assign _zz_22076 = ($signed(data_mid_98_imag) - $signed(data_mid_98_real));
  assign _zz_22077 = fixTo_2509_dout;
  assign _zz_22078 = _zz_22079[31 : 0];
  assign _zz_22079 = _zz_22080;
  assign _zz_22080 = ($signed(_zz_22081) >>> _zz_2094);
  assign _zz_22081 = _zz_22082;
  assign _zz_22082 = ($signed(_zz_22084) - $signed(_zz_2091));
  assign _zz_22083 = ({8'd0,data_mid_34_real} <<< 8);
  assign _zz_22084 = {{8{_zz_22083[23]}}, _zz_22083};
  assign _zz_22085 = fixTo_2510_dout;
  assign _zz_22086 = _zz_22087[31 : 0];
  assign _zz_22087 = _zz_22088;
  assign _zz_22088 = ($signed(_zz_22089) >>> _zz_2094);
  assign _zz_22089 = _zz_22090;
  assign _zz_22090 = ($signed(_zz_22092) - $signed(_zz_2092));
  assign _zz_22091 = ({8'd0,data_mid_34_imag} <<< 8);
  assign _zz_22092 = {{8{_zz_22091[23]}}, _zz_22091};
  assign _zz_22093 = fixTo_2511_dout;
  assign _zz_22094 = _zz_22095[31 : 0];
  assign _zz_22095 = _zz_22096;
  assign _zz_22096 = ($signed(_zz_22097) >>> _zz_2095);
  assign _zz_22097 = _zz_22098;
  assign _zz_22098 = ($signed(_zz_22100) + $signed(_zz_2091));
  assign _zz_22099 = ({8'd0,data_mid_34_real} <<< 8);
  assign _zz_22100 = {{8{_zz_22099[23]}}, _zz_22099};
  assign _zz_22101 = fixTo_2512_dout;
  assign _zz_22102 = _zz_22103[31 : 0];
  assign _zz_22103 = _zz_22104;
  assign _zz_22104 = ($signed(_zz_22105) >>> _zz_2095);
  assign _zz_22105 = _zz_22106;
  assign _zz_22106 = ($signed(_zz_22108) + $signed(_zz_2092));
  assign _zz_22107 = ({8'd0,data_mid_34_imag} <<< 8);
  assign _zz_22108 = {{8{_zz_22107[23]}}, _zz_22107};
  assign _zz_22109 = fixTo_2513_dout;
  assign _zz_22110 = ($signed(twiddle_factor_table_98_real) + $signed(twiddle_factor_table_98_imag));
  assign _zz_22111 = ($signed(_zz_2098) - $signed(_zz_22112));
  assign _zz_22112 = ($signed(_zz_22113) * $signed(twiddle_factor_table_98_imag));
  assign _zz_22113 = ($signed(data_mid_99_real) + $signed(data_mid_99_imag));
  assign _zz_22114 = fixTo_2514_dout;
  assign _zz_22115 = ($signed(_zz_2098) + $signed(_zz_22116));
  assign _zz_22116 = ($signed(_zz_22117) * $signed(twiddle_factor_table_98_real));
  assign _zz_22117 = ($signed(data_mid_99_imag) - $signed(data_mid_99_real));
  assign _zz_22118 = fixTo_2515_dout;
  assign _zz_22119 = _zz_22120[31 : 0];
  assign _zz_22120 = _zz_22121;
  assign _zz_22121 = ($signed(_zz_22122) >>> _zz_2099);
  assign _zz_22122 = _zz_22123;
  assign _zz_22123 = ($signed(_zz_22125) - $signed(_zz_2096));
  assign _zz_22124 = ({8'd0,data_mid_35_real} <<< 8);
  assign _zz_22125 = {{8{_zz_22124[23]}}, _zz_22124};
  assign _zz_22126 = fixTo_2516_dout;
  assign _zz_22127 = _zz_22128[31 : 0];
  assign _zz_22128 = _zz_22129;
  assign _zz_22129 = ($signed(_zz_22130) >>> _zz_2099);
  assign _zz_22130 = _zz_22131;
  assign _zz_22131 = ($signed(_zz_22133) - $signed(_zz_2097));
  assign _zz_22132 = ({8'd0,data_mid_35_imag} <<< 8);
  assign _zz_22133 = {{8{_zz_22132[23]}}, _zz_22132};
  assign _zz_22134 = fixTo_2517_dout;
  assign _zz_22135 = _zz_22136[31 : 0];
  assign _zz_22136 = _zz_22137;
  assign _zz_22137 = ($signed(_zz_22138) >>> _zz_2100);
  assign _zz_22138 = _zz_22139;
  assign _zz_22139 = ($signed(_zz_22141) + $signed(_zz_2096));
  assign _zz_22140 = ({8'd0,data_mid_35_real} <<< 8);
  assign _zz_22141 = {{8{_zz_22140[23]}}, _zz_22140};
  assign _zz_22142 = fixTo_2518_dout;
  assign _zz_22143 = _zz_22144[31 : 0];
  assign _zz_22144 = _zz_22145;
  assign _zz_22145 = ($signed(_zz_22146) >>> _zz_2100);
  assign _zz_22146 = _zz_22147;
  assign _zz_22147 = ($signed(_zz_22149) + $signed(_zz_2097));
  assign _zz_22148 = ({8'd0,data_mid_35_imag} <<< 8);
  assign _zz_22149 = {{8{_zz_22148[23]}}, _zz_22148};
  assign _zz_22150 = fixTo_2519_dout;
  assign _zz_22151 = ($signed(twiddle_factor_table_99_real) + $signed(twiddle_factor_table_99_imag));
  assign _zz_22152 = ($signed(_zz_2103) - $signed(_zz_22153));
  assign _zz_22153 = ($signed(_zz_22154) * $signed(twiddle_factor_table_99_imag));
  assign _zz_22154 = ($signed(data_mid_100_real) + $signed(data_mid_100_imag));
  assign _zz_22155 = fixTo_2520_dout;
  assign _zz_22156 = ($signed(_zz_2103) + $signed(_zz_22157));
  assign _zz_22157 = ($signed(_zz_22158) * $signed(twiddle_factor_table_99_real));
  assign _zz_22158 = ($signed(data_mid_100_imag) - $signed(data_mid_100_real));
  assign _zz_22159 = fixTo_2521_dout;
  assign _zz_22160 = _zz_22161[31 : 0];
  assign _zz_22161 = _zz_22162;
  assign _zz_22162 = ($signed(_zz_22163) >>> _zz_2104);
  assign _zz_22163 = _zz_22164;
  assign _zz_22164 = ($signed(_zz_22166) - $signed(_zz_2101));
  assign _zz_22165 = ({8'd0,data_mid_36_real} <<< 8);
  assign _zz_22166 = {{8{_zz_22165[23]}}, _zz_22165};
  assign _zz_22167 = fixTo_2522_dout;
  assign _zz_22168 = _zz_22169[31 : 0];
  assign _zz_22169 = _zz_22170;
  assign _zz_22170 = ($signed(_zz_22171) >>> _zz_2104);
  assign _zz_22171 = _zz_22172;
  assign _zz_22172 = ($signed(_zz_22174) - $signed(_zz_2102));
  assign _zz_22173 = ({8'd0,data_mid_36_imag} <<< 8);
  assign _zz_22174 = {{8{_zz_22173[23]}}, _zz_22173};
  assign _zz_22175 = fixTo_2523_dout;
  assign _zz_22176 = _zz_22177[31 : 0];
  assign _zz_22177 = _zz_22178;
  assign _zz_22178 = ($signed(_zz_22179) >>> _zz_2105);
  assign _zz_22179 = _zz_22180;
  assign _zz_22180 = ($signed(_zz_22182) + $signed(_zz_2101));
  assign _zz_22181 = ({8'd0,data_mid_36_real} <<< 8);
  assign _zz_22182 = {{8{_zz_22181[23]}}, _zz_22181};
  assign _zz_22183 = fixTo_2524_dout;
  assign _zz_22184 = _zz_22185[31 : 0];
  assign _zz_22185 = _zz_22186;
  assign _zz_22186 = ($signed(_zz_22187) >>> _zz_2105);
  assign _zz_22187 = _zz_22188;
  assign _zz_22188 = ($signed(_zz_22190) + $signed(_zz_2102));
  assign _zz_22189 = ({8'd0,data_mid_36_imag} <<< 8);
  assign _zz_22190 = {{8{_zz_22189[23]}}, _zz_22189};
  assign _zz_22191 = fixTo_2525_dout;
  assign _zz_22192 = ($signed(twiddle_factor_table_100_real) + $signed(twiddle_factor_table_100_imag));
  assign _zz_22193 = ($signed(_zz_2108) - $signed(_zz_22194));
  assign _zz_22194 = ($signed(_zz_22195) * $signed(twiddle_factor_table_100_imag));
  assign _zz_22195 = ($signed(data_mid_101_real) + $signed(data_mid_101_imag));
  assign _zz_22196 = fixTo_2526_dout;
  assign _zz_22197 = ($signed(_zz_2108) + $signed(_zz_22198));
  assign _zz_22198 = ($signed(_zz_22199) * $signed(twiddle_factor_table_100_real));
  assign _zz_22199 = ($signed(data_mid_101_imag) - $signed(data_mid_101_real));
  assign _zz_22200 = fixTo_2527_dout;
  assign _zz_22201 = _zz_22202[31 : 0];
  assign _zz_22202 = _zz_22203;
  assign _zz_22203 = ($signed(_zz_22204) >>> _zz_2109);
  assign _zz_22204 = _zz_22205;
  assign _zz_22205 = ($signed(_zz_22207) - $signed(_zz_2106));
  assign _zz_22206 = ({8'd0,data_mid_37_real} <<< 8);
  assign _zz_22207 = {{8{_zz_22206[23]}}, _zz_22206};
  assign _zz_22208 = fixTo_2528_dout;
  assign _zz_22209 = _zz_22210[31 : 0];
  assign _zz_22210 = _zz_22211;
  assign _zz_22211 = ($signed(_zz_22212) >>> _zz_2109);
  assign _zz_22212 = _zz_22213;
  assign _zz_22213 = ($signed(_zz_22215) - $signed(_zz_2107));
  assign _zz_22214 = ({8'd0,data_mid_37_imag} <<< 8);
  assign _zz_22215 = {{8{_zz_22214[23]}}, _zz_22214};
  assign _zz_22216 = fixTo_2529_dout;
  assign _zz_22217 = _zz_22218[31 : 0];
  assign _zz_22218 = _zz_22219;
  assign _zz_22219 = ($signed(_zz_22220) >>> _zz_2110);
  assign _zz_22220 = _zz_22221;
  assign _zz_22221 = ($signed(_zz_22223) + $signed(_zz_2106));
  assign _zz_22222 = ({8'd0,data_mid_37_real} <<< 8);
  assign _zz_22223 = {{8{_zz_22222[23]}}, _zz_22222};
  assign _zz_22224 = fixTo_2530_dout;
  assign _zz_22225 = _zz_22226[31 : 0];
  assign _zz_22226 = _zz_22227;
  assign _zz_22227 = ($signed(_zz_22228) >>> _zz_2110);
  assign _zz_22228 = _zz_22229;
  assign _zz_22229 = ($signed(_zz_22231) + $signed(_zz_2107));
  assign _zz_22230 = ({8'd0,data_mid_37_imag} <<< 8);
  assign _zz_22231 = {{8{_zz_22230[23]}}, _zz_22230};
  assign _zz_22232 = fixTo_2531_dout;
  assign _zz_22233 = ($signed(twiddle_factor_table_101_real) + $signed(twiddle_factor_table_101_imag));
  assign _zz_22234 = ($signed(_zz_2113) - $signed(_zz_22235));
  assign _zz_22235 = ($signed(_zz_22236) * $signed(twiddle_factor_table_101_imag));
  assign _zz_22236 = ($signed(data_mid_102_real) + $signed(data_mid_102_imag));
  assign _zz_22237 = fixTo_2532_dout;
  assign _zz_22238 = ($signed(_zz_2113) + $signed(_zz_22239));
  assign _zz_22239 = ($signed(_zz_22240) * $signed(twiddle_factor_table_101_real));
  assign _zz_22240 = ($signed(data_mid_102_imag) - $signed(data_mid_102_real));
  assign _zz_22241 = fixTo_2533_dout;
  assign _zz_22242 = _zz_22243[31 : 0];
  assign _zz_22243 = _zz_22244;
  assign _zz_22244 = ($signed(_zz_22245) >>> _zz_2114);
  assign _zz_22245 = _zz_22246;
  assign _zz_22246 = ($signed(_zz_22248) - $signed(_zz_2111));
  assign _zz_22247 = ({8'd0,data_mid_38_real} <<< 8);
  assign _zz_22248 = {{8{_zz_22247[23]}}, _zz_22247};
  assign _zz_22249 = fixTo_2534_dout;
  assign _zz_22250 = _zz_22251[31 : 0];
  assign _zz_22251 = _zz_22252;
  assign _zz_22252 = ($signed(_zz_22253) >>> _zz_2114);
  assign _zz_22253 = _zz_22254;
  assign _zz_22254 = ($signed(_zz_22256) - $signed(_zz_2112));
  assign _zz_22255 = ({8'd0,data_mid_38_imag} <<< 8);
  assign _zz_22256 = {{8{_zz_22255[23]}}, _zz_22255};
  assign _zz_22257 = fixTo_2535_dout;
  assign _zz_22258 = _zz_22259[31 : 0];
  assign _zz_22259 = _zz_22260;
  assign _zz_22260 = ($signed(_zz_22261) >>> _zz_2115);
  assign _zz_22261 = _zz_22262;
  assign _zz_22262 = ($signed(_zz_22264) + $signed(_zz_2111));
  assign _zz_22263 = ({8'd0,data_mid_38_real} <<< 8);
  assign _zz_22264 = {{8{_zz_22263[23]}}, _zz_22263};
  assign _zz_22265 = fixTo_2536_dout;
  assign _zz_22266 = _zz_22267[31 : 0];
  assign _zz_22267 = _zz_22268;
  assign _zz_22268 = ($signed(_zz_22269) >>> _zz_2115);
  assign _zz_22269 = _zz_22270;
  assign _zz_22270 = ($signed(_zz_22272) + $signed(_zz_2112));
  assign _zz_22271 = ({8'd0,data_mid_38_imag} <<< 8);
  assign _zz_22272 = {{8{_zz_22271[23]}}, _zz_22271};
  assign _zz_22273 = fixTo_2537_dout;
  assign _zz_22274 = ($signed(twiddle_factor_table_102_real) + $signed(twiddle_factor_table_102_imag));
  assign _zz_22275 = ($signed(_zz_2118) - $signed(_zz_22276));
  assign _zz_22276 = ($signed(_zz_22277) * $signed(twiddle_factor_table_102_imag));
  assign _zz_22277 = ($signed(data_mid_103_real) + $signed(data_mid_103_imag));
  assign _zz_22278 = fixTo_2538_dout;
  assign _zz_22279 = ($signed(_zz_2118) + $signed(_zz_22280));
  assign _zz_22280 = ($signed(_zz_22281) * $signed(twiddle_factor_table_102_real));
  assign _zz_22281 = ($signed(data_mid_103_imag) - $signed(data_mid_103_real));
  assign _zz_22282 = fixTo_2539_dout;
  assign _zz_22283 = _zz_22284[31 : 0];
  assign _zz_22284 = _zz_22285;
  assign _zz_22285 = ($signed(_zz_22286) >>> _zz_2119);
  assign _zz_22286 = _zz_22287;
  assign _zz_22287 = ($signed(_zz_22289) - $signed(_zz_2116));
  assign _zz_22288 = ({8'd0,data_mid_39_real} <<< 8);
  assign _zz_22289 = {{8{_zz_22288[23]}}, _zz_22288};
  assign _zz_22290 = fixTo_2540_dout;
  assign _zz_22291 = _zz_22292[31 : 0];
  assign _zz_22292 = _zz_22293;
  assign _zz_22293 = ($signed(_zz_22294) >>> _zz_2119);
  assign _zz_22294 = _zz_22295;
  assign _zz_22295 = ($signed(_zz_22297) - $signed(_zz_2117));
  assign _zz_22296 = ({8'd0,data_mid_39_imag} <<< 8);
  assign _zz_22297 = {{8{_zz_22296[23]}}, _zz_22296};
  assign _zz_22298 = fixTo_2541_dout;
  assign _zz_22299 = _zz_22300[31 : 0];
  assign _zz_22300 = _zz_22301;
  assign _zz_22301 = ($signed(_zz_22302) >>> _zz_2120);
  assign _zz_22302 = _zz_22303;
  assign _zz_22303 = ($signed(_zz_22305) + $signed(_zz_2116));
  assign _zz_22304 = ({8'd0,data_mid_39_real} <<< 8);
  assign _zz_22305 = {{8{_zz_22304[23]}}, _zz_22304};
  assign _zz_22306 = fixTo_2542_dout;
  assign _zz_22307 = _zz_22308[31 : 0];
  assign _zz_22308 = _zz_22309;
  assign _zz_22309 = ($signed(_zz_22310) >>> _zz_2120);
  assign _zz_22310 = _zz_22311;
  assign _zz_22311 = ($signed(_zz_22313) + $signed(_zz_2117));
  assign _zz_22312 = ({8'd0,data_mid_39_imag} <<< 8);
  assign _zz_22313 = {{8{_zz_22312[23]}}, _zz_22312};
  assign _zz_22314 = fixTo_2543_dout;
  assign _zz_22315 = ($signed(twiddle_factor_table_103_real) + $signed(twiddle_factor_table_103_imag));
  assign _zz_22316 = ($signed(_zz_2123) - $signed(_zz_22317));
  assign _zz_22317 = ($signed(_zz_22318) * $signed(twiddle_factor_table_103_imag));
  assign _zz_22318 = ($signed(data_mid_104_real) + $signed(data_mid_104_imag));
  assign _zz_22319 = fixTo_2544_dout;
  assign _zz_22320 = ($signed(_zz_2123) + $signed(_zz_22321));
  assign _zz_22321 = ($signed(_zz_22322) * $signed(twiddle_factor_table_103_real));
  assign _zz_22322 = ($signed(data_mid_104_imag) - $signed(data_mid_104_real));
  assign _zz_22323 = fixTo_2545_dout;
  assign _zz_22324 = _zz_22325[31 : 0];
  assign _zz_22325 = _zz_22326;
  assign _zz_22326 = ($signed(_zz_22327) >>> _zz_2124);
  assign _zz_22327 = _zz_22328;
  assign _zz_22328 = ($signed(_zz_22330) - $signed(_zz_2121));
  assign _zz_22329 = ({8'd0,data_mid_40_real} <<< 8);
  assign _zz_22330 = {{8{_zz_22329[23]}}, _zz_22329};
  assign _zz_22331 = fixTo_2546_dout;
  assign _zz_22332 = _zz_22333[31 : 0];
  assign _zz_22333 = _zz_22334;
  assign _zz_22334 = ($signed(_zz_22335) >>> _zz_2124);
  assign _zz_22335 = _zz_22336;
  assign _zz_22336 = ($signed(_zz_22338) - $signed(_zz_2122));
  assign _zz_22337 = ({8'd0,data_mid_40_imag} <<< 8);
  assign _zz_22338 = {{8{_zz_22337[23]}}, _zz_22337};
  assign _zz_22339 = fixTo_2547_dout;
  assign _zz_22340 = _zz_22341[31 : 0];
  assign _zz_22341 = _zz_22342;
  assign _zz_22342 = ($signed(_zz_22343) >>> _zz_2125);
  assign _zz_22343 = _zz_22344;
  assign _zz_22344 = ($signed(_zz_22346) + $signed(_zz_2121));
  assign _zz_22345 = ({8'd0,data_mid_40_real} <<< 8);
  assign _zz_22346 = {{8{_zz_22345[23]}}, _zz_22345};
  assign _zz_22347 = fixTo_2548_dout;
  assign _zz_22348 = _zz_22349[31 : 0];
  assign _zz_22349 = _zz_22350;
  assign _zz_22350 = ($signed(_zz_22351) >>> _zz_2125);
  assign _zz_22351 = _zz_22352;
  assign _zz_22352 = ($signed(_zz_22354) + $signed(_zz_2122));
  assign _zz_22353 = ({8'd0,data_mid_40_imag} <<< 8);
  assign _zz_22354 = {{8{_zz_22353[23]}}, _zz_22353};
  assign _zz_22355 = fixTo_2549_dout;
  assign _zz_22356 = ($signed(twiddle_factor_table_104_real) + $signed(twiddle_factor_table_104_imag));
  assign _zz_22357 = ($signed(_zz_2128) - $signed(_zz_22358));
  assign _zz_22358 = ($signed(_zz_22359) * $signed(twiddle_factor_table_104_imag));
  assign _zz_22359 = ($signed(data_mid_105_real) + $signed(data_mid_105_imag));
  assign _zz_22360 = fixTo_2550_dout;
  assign _zz_22361 = ($signed(_zz_2128) + $signed(_zz_22362));
  assign _zz_22362 = ($signed(_zz_22363) * $signed(twiddle_factor_table_104_real));
  assign _zz_22363 = ($signed(data_mid_105_imag) - $signed(data_mid_105_real));
  assign _zz_22364 = fixTo_2551_dout;
  assign _zz_22365 = _zz_22366[31 : 0];
  assign _zz_22366 = _zz_22367;
  assign _zz_22367 = ($signed(_zz_22368) >>> _zz_2129);
  assign _zz_22368 = _zz_22369;
  assign _zz_22369 = ($signed(_zz_22371) - $signed(_zz_2126));
  assign _zz_22370 = ({8'd0,data_mid_41_real} <<< 8);
  assign _zz_22371 = {{8{_zz_22370[23]}}, _zz_22370};
  assign _zz_22372 = fixTo_2552_dout;
  assign _zz_22373 = _zz_22374[31 : 0];
  assign _zz_22374 = _zz_22375;
  assign _zz_22375 = ($signed(_zz_22376) >>> _zz_2129);
  assign _zz_22376 = _zz_22377;
  assign _zz_22377 = ($signed(_zz_22379) - $signed(_zz_2127));
  assign _zz_22378 = ({8'd0,data_mid_41_imag} <<< 8);
  assign _zz_22379 = {{8{_zz_22378[23]}}, _zz_22378};
  assign _zz_22380 = fixTo_2553_dout;
  assign _zz_22381 = _zz_22382[31 : 0];
  assign _zz_22382 = _zz_22383;
  assign _zz_22383 = ($signed(_zz_22384) >>> _zz_2130);
  assign _zz_22384 = _zz_22385;
  assign _zz_22385 = ($signed(_zz_22387) + $signed(_zz_2126));
  assign _zz_22386 = ({8'd0,data_mid_41_real} <<< 8);
  assign _zz_22387 = {{8{_zz_22386[23]}}, _zz_22386};
  assign _zz_22388 = fixTo_2554_dout;
  assign _zz_22389 = _zz_22390[31 : 0];
  assign _zz_22390 = _zz_22391;
  assign _zz_22391 = ($signed(_zz_22392) >>> _zz_2130);
  assign _zz_22392 = _zz_22393;
  assign _zz_22393 = ($signed(_zz_22395) + $signed(_zz_2127));
  assign _zz_22394 = ({8'd0,data_mid_41_imag} <<< 8);
  assign _zz_22395 = {{8{_zz_22394[23]}}, _zz_22394};
  assign _zz_22396 = fixTo_2555_dout;
  assign _zz_22397 = ($signed(twiddle_factor_table_105_real) + $signed(twiddle_factor_table_105_imag));
  assign _zz_22398 = ($signed(_zz_2133) - $signed(_zz_22399));
  assign _zz_22399 = ($signed(_zz_22400) * $signed(twiddle_factor_table_105_imag));
  assign _zz_22400 = ($signed(data_mid_106_real) + $signed(data_mid_106_imag));
  assign _zz_22401 = fixTo_2556_dout;
  assign _zz_22402 = ($signed(_zz_2133) + $signed(_zz_22403));
  assign _zz_22403 = ($signed(_zz_22404) * $signed(twiddle_factor_table_105_real));
  assign _zz_22404 = ($signed(data_mid_106_imag) - $signed(data_mid_106_real));
  assign _zz_22405 = fixTo_2557_dout;
  assign _zz_22406 = _zz_22407[31 : 0];
  assign _zz_22407 = _zz_22408;
  assign _zz_22408 = ($signed(_zz_22409) >>> _zz_2134);
  assign _zz_22409 = _zz_22410;
  assign _zz_22410 = ($signed(_zz_22412) - $signed(_zz_2131));
  assign _zz_22411 = ({8'd0,data_mid_42_real} <<< 8);
  assign _zz_22412 = {{8{_zz_22411[23]}}, _zz_22411};
  assign _zz_22413 = fixTo_2558_dout;
  assign _zz_22414 = _zz_22415[31 : 0];
  assign _zz_22415 = _zz_22416;
  assign _zz_22416 = ($signed(_zz_22417) >>> _zz_2134);
  assign _zz_22417 = _zz_22418;
  assign _zz_22418 = ($signed(_zz_22420) - $signed(_zz_2132));
  assign _zz_22419 = ({8'd0,data_mid_42_imag} <<< 8);
  assign _zz_22420 = {{8{_zz_22419[23]}}, _zz_22419};
  assign _zz_22421 = fixTo_2559_dout;
  assign _zz_22422 = _zz_22423[31 : 0];
  assign _zz_22423 = _zz_22424;
  assign _zz_22424 = ($signed(_zz_22425) >>> _zz_2135);
  assign _zz_22425 = _zz_22426;
  assign _zz_22426 = ($signed(_zz_22428) + $signed(_zz_2131));
  assign _zz_22427 = ({8'd0,data_mid_42_real} <<< 8);
  assign _zz_22428 = {{8{_zz_22427[23]}}, _zz_22427};
  assign _zz_22429 = fixTo_2560_dout;
  assign _zz_22430 = _zz_22431[31 : 0];
  assign _zz_22431 = _zz_22432;
  assign _zz_22432 = ($signed(_zz_22433) >>> _zz_2135);
  assign _zz_22433 = _zz_22434;
  assign _zz_22434 = ($signed(_zz_22436) + $signed(_zz_2132));
  assign _zz_22435 = ({8'd0,data_mid_42_imag} <<< 8);
  assign _zz_22436 = {{8{_zz_22435[23]}}, _zz_22435};
  assign _zz_22437 = fixTo_2561_dout;
  assign _zz_22438 = ($signed(twiddle_factor_table_106_real) + $signed(twiddle_factor_table_106_imag));
  assign _zz_22439 = ($signed(_zz_2138) - $signed(_zz_22440));
  assign _zz_22440 = ($signed(_zz_22441) * $signed(twiddle_factor_table_106_imag));
  assign _zz_22441 = ($signed(data_mid_107_real) + $signed(data_mid_107_imag));
  assign _zz_22442 = fixTo_2562_dout;
  assign _zz_22443 = ($signed(_zz_2138) + $signed(_zz_22444));
  assign _zz_22444 = ($signed(_zz_22445) * $signed(twiddle_factor_table_106_real));
  assign _zz_22445 = ($signed(data_mid_107_imag) - $signed(data_mid_107_real));
  assign _zz_22446 = fixTo_2563_dout;
  assign _zz_22447 = _zz_22448[31 : 0];
  assign _zz_22448 = _zz_22449;
  assign _zz_22449 = ($signed(_zz_22450) >>> _zz_2139);
  assign _zz_22450 = _zz_22451;
  assign _zz_22451 = ($signed(_zz_22453) - $signed(_zz_2136));
  assign _zz_22452 = ({8'd0,data_mid_43_real} <<< 8);
  assign _zz_22453 = {{8{_zz_22452[23]}}, _zz_22452};
  assign _zz_22454 = fixTo_2564_dout;
  assign _zz_22455 = _zz_22456[31 : 0];
  assign _zz_22456 = _zz_22457;
  assign _zz_22457 = ($signed(_zz_22458) >>> _zz_2139);
  assign _zz_22458 = _zz_22459;
  assign _zz_22459 = ($signed(_zz_22461) - $signed(_zz_2137));
  assign _zz_22460 = ({8'd0,data_mid_43_imag} <<< 8);
  assign _zz_22461 = {{8{_zz_22460[23]}}, _zz_22460};
  assign _zz_22462 = fixTo_2565_dout;
  assign _zz_22463 = _zz_22464[31 : 0];
  assign _zz_22464 = _zz_22465;
  assign _zz_22465 = ($signed(_zz_22466) >>> _zz_2140);
  assign _zz_22466 = _zz_22467;
  assign _zz_22467 = ($signed(_zz_22469) + $signed(_zz_2136));
  assign _zz_22468 = ({8'd0,data_mid_43_real} <<< 8);
  assign _zz_22469 = {{8{_zz_22468[23]}}, _zz_22468};
  assign _zz_22470 = fixTo_2566_dout;
  assign _zz_22471 = _zz_22472[31 : 0];
  assign _zz_22472 = _zz_22473;
  assign _zz_22473 = ($signed(_zz_22474) >>> _zz_2140);
  assign _zz_22474 = _zz_22475;
  assign _zz_22475 = ($signed(_zz_22477) + $signed(_zz_2137));
  assign _zz_22476 = ({8'd0,data_mid_43_imag} <<< 8);
  assign _zz_22477 = {{8{_zz_22476[23]}}, _zz_22476};
  assign _zz_22478 = fixTo_2567_dout;
  assign _zz_22479 = ($signed(twiddle_factor_table_107_real) + $signed(twiddle_factor_table_107_imag));
  assign _zz_22480 = ($signed(_zz_2143) - $signed(_zz_22481));
  assign _zz_22481 = ($signed(_zz_22482) * $signed(twiddle_factor_table_107_imag));
  assign _zz_22482 = ($signed(data_mid_108_real) + $signed(data_mid_108_imag));
  assign _zz_22483 = fixTo_2568_dout;
  assign _zz_22484 = ($signed(_zz_2143) + $signed(_zz_22485));
  assign _zz_22485 = ($signed(_zz_22486) * $signed(twiddle_factor_table_107_real));
  assign _zz_22486 = ($signed(data_mid_108_imag) - $signed(data_mid_108_real));
  assign _zz_22487 = fixTo_2569_dout;
  assign _zz_22488 = _zz_22489[31 : 0];
  assign _zz_22489 = _zz_22490;
  assign _zz_22490 = ($signed(_zz_22491) >>> _zz_2144);
  assign _zz_22491 = _zz_22492;
  assign _zz_22492 = ($signed(_zz_22494) - $signed(_zz_2141));
  assign _zz_22493 = ({8'd0,data_mid_44_real} <<< 8);
  assign _zz_22494 = {{8{_zz_22493[23]}}, _zz_22493};
  assign _zz_22495 = fixTo_2570_dout;
  assign _zz_22496 = _zz_22497[31 : 0];
  assign _zz_22497 = _zz_22498;
  assign _zz_22498 = ($signed(_zz_22499) >>> _zz_2144);
  assign _zz_22499 = _zz_22500;
  assign _zz_22500 = ($signed(_zz_22502) - $signed(_zz_2142));
  assign _zz_22501 = ({8'd0,data_mid_44_imag} <<< 8);
  assign _zz_22502 = {{8{_zz_22501[23]}}, _zz_22501};
  assign _zz_22503 = fixTo_2571_dout;
  assign _zz_22504 = _zz_22505[31 : 0];
  assign _zz_22505 = _zz_22506;
  assign _zz_22506 = ($signed(_zz_22507) >>> _zz_2145);
  assign _zz_22507 = _zz_22508;
  assign _zz_22508 = ($signed(_zz_22510) + $signed(_zz_2141));
  assign _zz_22509 = ({8'd0,data_mid_44_real} <<< 8);
  assign _zz_22510 = {{8{_zz_22509[23]}}, _zz_22509};
  assign _zz_22511 = fixTo_2572_dout;
  assign _zz_22512 = _zz_22513[31 : 0];
  assign _zz_22513 = _zz_22514;
  assign _zz_22514 = ($signed(_zz_22515) >>> _zz_2145);
  assign _zz_22515 = _zz_22516;
  assign _zz_22516 = ($signed(_zz_22518) + $signed(_zz_2142));
  assign _zz_22517 = ({8'd0,data_mid_44_imag} <<< 8);
  assign _zz_22518 = {{8{_zz_22517[23]}}, _zz_22517};
  assign _zz_22519 = fixTo_2573_dout;
  assign _zz_22520 = ($signed(twiddle_factor_table_108_real) + $signed(twiddle_factor_table_108_imag));
  assign _zz_22521 = ($signed(_zz_2148) - $signed(_zz_22522));
  assign _zz_22522 = ($signed(_zz_22523) * $signed(twiddle_factor_table_108_imag));
  assign _zz_22523 = ($signed(data_mid_109_real) + $signed(data_mid_109_imag));
  assign _zz_22524 = fixTo_2574_dout;
  assign _zz_22525 = ($signed(_zz_2148) + $signed(_zz_22526));
  assign _zz_22526 = ($signed(_zz_22527) * $signed(twiddle_factor_table_108_real));
  assign _zz_22527 = ($signed(data_mid_109_imag) - $signed(data_mid_109_real));
  assign _zz_22528 = fixTo_2575_dout;
  assign _zz_22529 = _zz_22530[31 : 0];
  assign _zz_22530 = _zz_22531;
  assign _zz_22531 = ($signed(_zz_22532) >>> _zz_2149);
  assign _zz_22532 = _zz_22533;
  assign _zz_22533 = ($signed(_zz_22535) - $signed(_zz_2146));
  assign _zz_22534 = ({8'd0,data_mid_45_real} <<< 8);
  assign _zz_22535 = {{8{_zz_22534[23]}}, _zz_22534};
  assign _zz_22536 = fixTo_2576_dout;
  assign _zz_22537 = _zz_22538[31 : 0];
  assign _zz_22538 = _zz_22539;
  assign _zz_22539 = ($signed(_zz_22540) >>> _zz_2149);
  assign _zz_22540 = _zz_22541;
  assign _zz_22541 = ($signed(_zz_22543) - $signed(_zz_2147));
  assign _zz_22542 = ({8'd0,data_mid_45_imag} <<< 8);
  assign _zz_22543 = {{8{_zz_22542[23]}}, _zz_22542};
  assign _zz_22544 = fixTo_2577_dout;
  assign _zz_22545 = _zz_22546[31 : 0];
  assign _zz_22546 = _zz_22547;
  assign _zz_22547 = ($signed(_zz_22548) >>> _zz_2150);
  assign _zz_22548 = _zz_22549;
  assign _zz_22549 = ($signed(_zz_22551) + $signed(_zz_2146));
  assign _zz_22550 = ({8'd0,data_mid_45_real} <<< 8);
  assign _zz_22551 = {{8{_zz_22550[23]}}, _zz_22550};
  assign _zz_22552 = fixTo_2578_dout;
  assign _zz_22553 = _zz_22554[31 : 0];
  assign _zz_22554 = _zz_22555;
  assign _zz_22555 = ($signed(_zz_22556) >>> _zz_2150);
  assign _zz_22556 = _zz_22557;
  assign _zz_22557 = ($signed(_zz_22559) + $signed(_zz_2147));
  assign _zz_22558 = ({8'd0,data_mid_45_imag} <<< 8);
  assign _zz_22559 = {{8{_zz_22558[23]}}, _zz_22558};
  assign _zz_22560 = fixTo_2579_dout;
  assign _zz_22561 = ($signed(twiddle_factor_table_109_real) + $signed(twiddle_factor_table_109_imag));
  assign _zz_22562 = ($signed(_zz_2153) - $signed(_zz_22563));
  assign _zz_22563 = ($signed(_zz_22564) * $signed(twiddle_factor_table_109_imag));
  assign _zz_22564 = ($signed(data_mid_110_real) + $signed(data_mid_110_imag));
  assign _zz_22565 = fixTo_2580_dout;
  assign _zz_22566 = ($signed(_zz_2153) + $signed(_zz_22567));
  assign _zz_22567 = ($signed(_zz_22568) * $signed(twiddle_factor_table_109_real));
  assign _zz_22568 = ($signed(data_mid_110_imag) - $signed(data_mid_110_real));
  assign _zz_22569 = fixTo_2581_dout;
  assign _zz_22570 = _zz_22571[31 : 0];
  assign _zz_22571 = _zz_22572;
  assign _zz_22572 = ($signed(_zz_22573) >>> _zz_2154);
  assign _zz_22573 = _zz_22574;
  assign _zz_22574 = ($signed(_zz_22576) - $signed(_zz_2151));
  assign _zz_22575 = ({8'd0,data_mid_46_real} <<< 8);
  assign _zz_22576 = {{8{_zz_22575[23]}}, _zz_22575};
  assign _zz_22577 = fixTo_2582_dout;
  assign _zz_22578 = _zz_22579[31 : 0];
  assign _zz_22579 = _zz_22580;
  assign _zz_22580 = ($signed(_zz_22581) >>> _zz_2154);
  assign _zz_22581 = _zz_22582;
  assign _zz_22582 = ($signed(_zz_22584) - $signed(_zz_2152));
  assign _zz_22583 = ({8'd0,data_mid_46_imag} <<< 8);
  assign _zz_22584 = {{8{_zz_22583[23]}}, _zz_22583};
  assign _zz_22585 = fixTo_2583_dout;
  assign _zz_22586 = _zz_22587[31 : 0];
  assign _zz_22587 = _zz_22588;
  assign _zz_22588 = ($signed(_zz_22589) >>> _zz_2155);
  assign _zz_22589 = _zz_22590;
  assign _zz_22590 = ($signed(_zz_22592) + $signed(_zz_2151));
  assign _zz_22591 = ({8'd0,data_mid_46_real} <<< 8);
  assign _zz_22592 = {{8{_zz_22591[23]}}, _zz_22591};
  assign _zz_22593 = fixTo_2584_dout;
  assign _zz_22594 = _zz_22595[31 : 0];
  assign _zz_22595 = _zz_22596;
  assign _zz_22596 = ($signed(_zz_22597) >>> _zz_2155);
  assign _zz_22597 = _zz_22598;
  assign _zz_22598 = ($signed(_zz_22600) + $signed(_zz_2152));
  assign _zz_22599 = ({8'd0,data_mid_46_imag} <<< 8);
  assign _zz_22600 = {{8{_zz_22599[23]}}, _zz_22599};
  assign _zz_22601 = fixTo_2585_dout;
  assign _zz_22602 = ($signed(twiddle_factor_table_110_real) + $signed(twiddle_factor_table_110_imag));
  assign _zz_22603 = ($signed(_zz_2158) - $signed(_zz_22604));
  assign _zz_22604 = ($signed(_zz_22605) * $signed(twiddle_factor_table_110_imag));
  assign _zz_22605 = ($signed(data_mid_111_real) + $signed(data_mid_111_imag));
  assign _zz_22606 = fixTo_2586_dout;
  assign _zz_22607 = ($signed(_zz_2158) + $signed(_zz_22608));
  assign _zz_22608 = ($signed(_zz_22609) * $signed(twiddle_factor_table_110_real));
  assign _zz_22609 = ($signed(data_mid_111_imag) - $signed(data_mid_111_real));
  assign _zz_22610 = fixTo_2587_dout;
  assign _zz_22611 = _zz_22612[31 : 0];
  assign _zz_22612 = _zz_22613;
  assign _zz_22613 = ($signed(_zz_22614) >>> _zz_2159);
  assign _zz_22614 = _zz_22615;
  assign _zz_22615 = ($signed(_zz_22617) - $signed(_zz_2156));
  assign _zz_22616 = ({8'd0,data_mid_47_real} <<< 8);
  assign _zz_22617 = {{8{_zz_22616[23]}}, _zz_22616};
  assign _zz_22618 = fixTo_2588_dout;
  assign _zz_22619 = _zz_22620[31 : 0];
  assign _zz_22620 = _zz_22621;
  assign _zz_22621 = ($signed(_zz_22622) >>> _zz_2159);
  assign _zz_22622 = _zz_22623;
  assign _zz_22623 = ($signed(_zz_22625) - $signed(_zz_2157));
  assign _zz_22624 = ({8'd0,data_mid_47_imag} <<< 8);
  assign _zz_22625 = {{8{_zz_22624[23]}}, _zz_22624};
  assign _zz_22626 = fixTo_2589_dout;
  assign _zz_22627 = _zz_22628[31 : 0];
  assign _zz_22628 = _zz_22629;
  assign _zz_22629 = ($signed(_zz_22630) >>> _zz_2160);
  assign _zz_22630 = _zz_22631;
  assign _zz_22631 = ($signed(_zz_22633) + $signed(_zz_2156));
  assign _zz_22632 = ({8'd0,data_mid_47_real} <<< 8);
  assign _zz_22633 = {{8{_zz_22632[23]}}, _zz_22632};
  assign _zz_22634 = fixTo_2590_dout;
  assign _zz_22635 = _zz_22636[31 : 0];
  assign _zz_22636 = _zz_22637;
  assign _zz_22637 = ($signed(_zz_22638) >>> _zz_2160);
  assign _zz_22638 = _zz_22639;
  assign _zz_22639 = ($signed(_zz_22641) + $signed(_zz_2157));
  assign _zz_22640 = ({8'd0,data_mid_47_imag} <<< 8);
  assign _zz_22641 = {{8{_zz_22640[23]}}, _zz_22640};
  assign _zz_22642 = fixTo_2591_dout;
  assign _zz_22643 = ($signed(twiddle_factor_table_111_real) + $signed(twiddle_factor_table_111_imag));
  assign _zz_22644 = ($signed(_zz_2163) - $signed(_zz_22645));
  assign _zz_22645 = ($signed(_zz_22646) * $signed(twiddle_factor_table_111_imag));
  assign _zz_22646 = ($signed(data_mid_112_real) + $signed(data_mid_112_imag));
  assign _zz_22647 = fixTo_2592_dout;
  assign _zz_22648 = ($signed(_zz_2163) + $signed(_zz_22649));
  assign _zz_22649 = ($signed(_zz_22650) * $signed(twiddle_factor_table_111_real));
  assign _zz_22650 = ($signed(data_mid_112_imag) - $signed(data_mid_112_real));
  assign _zz_22651 = fixTo_2593_dout;
  assign _zz_22652 = _zz_22653[31 : 0];
  assign _zz_22653 = _zz_22654;
  assign _zz_22654 = ($signed(_zz_22655) >>> _zz_2164);
  assign _zz_22655 = _zz_22656;
  assign _zz_22656 = ($signed(_zz_22658) - $signed(_zz_2161));
  assign _zz_22657 = ({8'd0,data_mid_48_real} <<< 8);
  assign _zz_22658 = {{8{_zz_22657[23]}}, _zz_22657};
  assign _zz_22659 = fixTo_2594_dout;
  assign _zz_22660 = _zz_22661[31 : 0];
  assign _zz_22661 = _zz_22662;
  assign _zz_22662 = ($signed(_zz_22663) >>> _zz_2164);
  assign _zz_22663 = _zz_22664;
  assign _zz_22664 = ($signed(_zz_22666) - $signed(_zz_2162));
  assign _zz_22665 = ({8'd0,data_mid_48_imag} <<< 8);
  assign _zz_22666 = {{8{_zz_22665[23]}}, _zz_22665};
  assign _zz_22667 = fixTo_2595_dout;
  assign _zz_22668 = _zz_22669[31 : 0];
  assign _zz_22669 = _zz_22670;
  assign _zz_22670 = ($signed(_zz_22671) >>> _zz_2165);
  assign _zz_22671 = _zz_22672;
  assign _zz_22672 = ($signed(_zz_22674) + $signed(_zz_2161));
  assign _zz_22673 = ({8'd0,data_mid_48_real} <<< 8);
  assign _zz_22674 = {{8{_zz_22673[23]}}, _zz_22673};
  assign _zz_22675 = fixTo_2596_dout;
  assign _zz_22676 = _zz_22677[31 : 0];
  assign _zz_22677 = _zz_22678;
  assign _zz_22678 = ($signed(_zz_22679) >>> _zz_2165);
  assign _zz_22679 = _zz_22680;
  assign _zz_22680 = ($signed(_zz_22682) + $signed(_zz_2162));
  assign _zz_22681 = ({8'd0,data_mid_48_imag} <<< 8);
  assign _zz_22682 = {{8{_zz_22681[23]}}, _zz_22681};
  assign _zz_22683 = fixTo_2597_dout;
  assign _zz_22684 = ($signed(twiddle_factor_table_112_real) + $signed(twiddle_factor_table_112_imag));
  assign _zz_22685 = ($signed(_zz_2168) - $signed(_zz_22686));
  assign _zz_22686 = ($signed(_zz_22687) * $signed(twiddle_factor_table_112_imag));
  assign _zz_22687 = ($signed(data_mid_113_real) + $signed(data_mid_113_imag));
  assign _zz_22688 = fixTo_2598_dout;
  assign _zz_22689 = ($signed(_zz_2168) + $signed(_zz_22690));
  assign _zz_22690 = ($signed(_zz_22691) * $signed(twiddle_factor_table_112_real));
  assign _zz_22691 = ($signed(data_mid_113_imag) - $signed(data_mid_113_real));
  assign _zz_22692 = fixTo_2599_dout;
  assign _zz_22693 = _zz_22694[31 : 0];
  assign _zz_22694 = _zz_22695;
  assign _zz_22695 = ($signed(_zz_22696) >>> _zz_2169);
  assign _zz_22696 = _zz_22697;
  assign _zz_22697 = ($signed(_zz_22699) - $signed(_zz_2166));
  assign _zz_22698 = ({8'd0,data_mid_49_real} <<< 8);
  assign _zz_22699 = {{8{_zz_22698[23]}}, _zz_22698};
  assign _zz_22700 = fixTo_2600_dout;
  assign _zz_22701 = _zz_22702[31 : 0];
  assign _zz_22702 = _zz_22703;
  assign _zz_22703 = ($signed(_zz_22704) >>> _zz_2169);
  assign _zz_22704 = _zz_22705;
  assign _zz_22705 = ($signed(_zz_22707) - $signed(_zz_2167));
  assign _zz_22706 = ({8'd0,data_mid_49_imag} <<< 8);
  assign _zz_22707 = {{8{_zz_22706[23]}}, _zz_22706};
  assign _zz_22708 = fixTo_2601_dout;
  assign _zz_22709 = _zz_22710[31 : 0];
  assign _zz_22710 = _zz_22711;
  assign _zz_22711 = ($signed(_zz_22712) >>> _zz_2170);
  assign _zz_22712 = _zz_22713;
  assign _zz_22713 = ($signed(_zz_22715) + $signed(_zz_2166));
  assign _zz_22714 = ({8'd0,data_mid_49_real} <<< 8);
  assign _zz_22715 = {{8{_zz_22714[23]}}, _zz_22714};
  assign _zz_22716 = fixTo_2602_dout;
  assign _zz_22717 = _zz_22718[31 : 0];
  assign _zz_22718 = _zz_22719;
  assign _zz_22719 = ($signed(_zz_22720) >>> _zz_2170);
  assign _zz_22720 = _zz_22721;
  assign _zz_22721 = ($signed(_zz_22723) + $signed(_zz_2167));
  assign _zz_22722 = ({8'd0,data_mid_49_imag} <<< 8);
  assign _zz_22723 = {{8{_zz_22722[23]}}, _zz_22722};
  assign _zz_22724 = fixTo_2603_dout;
  assign _zz_22725 = ($signed(twiddle_factor_table_113_real) + $signed(twiddle_factor_table_113_imag));
  assign _zz_22726 = ($signed(_zz_2173) - $signed(_zz_22727));
  assign _zz_22727 = ($signed(_zz_22728) * $signed(twiddle_factor_table_113_imag));
  assign _zz_22728 = ($signed(data_mid_114_real) + $signed(data_mid_114_imag));
  assign _zz_22729 = fixTo_2604_dout;
  assign _zz_22730 = ($signed(_zz_2173) + $signed(_zz_22731));
  assign _zz_22731 = ($signed(_zz_22732) * $signed(twiddle_factor_table_113_real));
  assign _zz_22732 = ($signed(data_mid_114_imag) - $signed(data_mid_114_real));
  assign _zz_22733 = fixTo_2605_dout;
  assign _zz_22734 = _zz_22735[31 : 0];
  assign _zz_22735 = _zz_22736;
  assign _zz_22736 = ($signed(_zz_22737) >>> _zz_2174);
  assign _zz_22737 = _zz_22738;
  assign _zz_22738 = ($signed(_zz_22740) - $signed(_zz_2171));
  assign _zz_22739 = ({8'd0,data_mid_50_real} <<< 8);
  assign _zz_22740 = {{8{_zz_22739[23]}}, _zz_22739};
  assign _zz_22741 = fixTo_2606_dout;
  assign _zz_22742 = _zz_22743[31 : 0];
  assign _zz_22743 = _zz_22744;
  assign _zz_22744 = ($signed(_zz_22745) >>> _zz_2174);
  assign _zz_22745 = _zz_22746;
  assign _zz_22746 = ($signed(_zz_22748) - $signed(_zz_2172));
  assign _zz_22747 = ({8'd0,data_mid_50_imag} <<< 8);
  assign _zz_22748 = {{8{_zz_22747[23]}}, _zz_22747};
  assign _zz_22749 = fixTo_2607_dout;
  assign _zz_22750 = _zz_22751[31 : 0];
  assign _zz_22751 = _zz_22752;
  assign _zz_22752 = ($signed(_zz_22753) >>> _zz_2175);
  assign _zz_22753 = _zz_22754;
  assign _zz_22754 = ($signed(_zz_22756) + $signed(_zz_2171));
  assign _zz_22755 = ({8'd0,data_mid_50_real} <<< 8);
  assign _zz_22756 = {{8{_zz_22755[23]}}, _zz_22755};
  assign _zz_22757 = fixTo_2608_dout;
  assign _zz_22758 = _zz_22759[31 : 0];
  assign _zz_22759 = _zz_22760;
  assign _zz_22760 = ($signed(_zz_22761) >>> _zz_2175);
  assign _zz_22761 = _zz_22762;
  assign _zz_22762 = ($signed(_zz_22764) + $signed(_zz_2172));
  assign _zz_22763 = ({8'd0,data_mid_50_imag} <<< 8);
  assign _zz_22764 = {{8{_zz_22763[23]}}, _zz_22763};
  assign _zz_22765 = fixTo_2609_dout;
  assign _zz_22766 = ($signed(twiddle_factor_table_114_real) + $signed(twiddle_factor_table_114_imag));
  assign _zz_22767 = ($signed(_zz_2178) - $signed(_zz_22768));
  assign _zz_22768 = ($signed(_zz_22769) * $signed(twiddle_factor_table_114_imag));
  assign _zz_22769 = ($signed(data_mid_115_real) + $signed(data_mid_115_imag));
  assign _zz_22770 = fixTo_2610_dout;
  assign _zz_22771 = ($signed(_zz_2178) + $signed(_zz_22772));
  assign _zz_22772 = ($signed(_zz_22773) * $signed(twiddle_factor_table_114_real));
  assign _zz_22773 = ($signed(data_mid_115_imag) - $signed(data_mid_115_real));
  assign _zz_22774 = fixTo_2611_dout;
  assign _zz_22775 = _zz_22776[31 : 0];
  assign _zz_22776 = _zz_22777;
  assign _zz_22777 = ($signed(_zz_22778) >>> _zz_2179);
  assign _zz_22778 = _zz_22779;
  assign _zz_22779 = ($signed(_zz_22781) - $signed(_zz_2176));
  assign _zz_22780 = ({8'd0,data_mid_51_real} <<< 8);
  assign _zz_22781 = {{8{_zz_22780[23]}}, _zz_22780};
  assign _zz_22782 = fixTo_2612_dout;
  assign _zz_22783 = _zz_22784[31 : 0];
  assign _zz_22784 = _zz_22785;
  assign _zz_22785 = ($signed(_zz_22786) >>> _zz_2179);
  assign _zz_22786 = _zz_22787;
  assign _zz_22787 = ($signed(_zz_22789) - $signed(_zz_2177));
  assign _zz_22788 = ({8'd0,data_mid_51_imag} <<< 8);
  assign _zz_22789 = {{8{_zz_22788[23]}}, _zz_22788};
  assign _zz_22790 = fixTo_2613_dout;
  assign _zz_22791 = _zz_22792[31 : 0];
  assign _zz_22792 = _zz_22793;
  assign _zz_22793 = ($signed(_zz_22794) >>> _zz_2180);
  assign _zz_22794 = _zz_22795;
  assign _zz_22795 = ($signed(_zz_22797) + $signed(_zz_2176));
  assign _zz_22796 = ({8'd0,data_mid_51_real} <<< 8);
  assign _zz_22797 = {{8{_zz_22796[23]}}, _zz_22796};
  assign _zz_22798 = fixTo_2614_dout;
  assign _zz_22799 = _zz_22800[31 : 0];
  assign _zz_22800 = _zz_22801;
  assign _zz_22801 = ($signed(_zz_22802) >>> _zz_2180);
  assign _zz_22802 = _zz_22803;
  assign _zz_22803 = ($signed(_zz_22805) + $signed(_zz_2177));
  assign _zz_22804 = ({8'd0,data_mid_51_imag} <<< 8);
  assign _zz_22805 = {{8{_zz_22804[23]}}, _zz_22804};
  assign _zz_22806 = fixTo_2615_dout;
  assign _zz_22807 = ($signed(twiddle_factor_table_115_real) + $signed(twiddle_factor_table_115_imag));
  assign _zz_22808 = ($signed(_zz_2183) - $signed(_zz_22809));
  assign _zz_22809 = ($signed(_zz_22810) * $signed(twiddle_factor_table_115_imag));
  assign _zz_22810 = ($signed(data_mid_116_real) + $signed(data_mid_116_imag));
  assign _zz_22811 = fixTo_2616_dout;
  assign _zz_22812 = ($signed(_zz_2183) + $signed(_zz_22813));
  assign _zz_22813 = ($signed(_zz_22814) * $signed(twiddle_factor_table_115_real));
  assign _zz_22814 = ($signed(data_mid_116_imag) - $signed(data_mid_116_real));
  assign _zz_22815 = fixTo_2617_dout;
  assign _zz_22816 = _zz_22817[31 : 0];
  assign _zz_22817 = _zz_22818;
  assign _zz_22818 = ($signed(_zz_22819) >>> _zz_2184);
  assign _zz_22819 = _zz_22820;
  assign _zz_22820 = ($signed(_zz_22822) - $signed(_zz_2181));
  assign _zz_22821 = ({8'd0,data_mid_52_real} <<< 8);
  assign _zz_22822 = {{8{_zz_22821[23]}}, _zz_22821};
  assign _zz_22823 = fixTo_2618_dout;
  assign _zz_22824 = _zz_22825[31 : 0];
  assign _zz_22825 = _zz_22826;
  assign _zz_22826 = ($signed(_zz_22827) >>> _zz_2184);
  assign _zz_22827 = _zz_22828;
  assign _zz_22828 = ($signed(_zz_22830) - $signed(_zz_2182));
  assign _zz_22829 = ({8'd0,data_mid_52_imag} <<< 8);
  assign _zz_22830 = {{8{_zz_22829[23]}}, _zz_22829};
  assign _zz_22831 = fixTo_2619_dout;
  assign _zz_22832 = _zz_22833[31 : 0];
  assign _zz_22833 = _zz_22834;
  assign _zz_22834 = ($signed(_zz_22835) >>> _zz_2185);
  assign _zz_22835 = _zz_22836;
  assign _zz_22836 = ($signed(_zz_22838) + $signed(_zz_2181));
  assign _zz_22837 = ({8'd0,data_mid_52_real} <<< 8);
  assign _zz_22838 = {{8{_zz_22837[23]}}, _zz_22837};
  assign _zz_22839 = fixTo_2620_dout;
  assign _zz_22840 = _zz_22841[31 : 0];
  assign _zz_22841 = _zz_22842;
  assign _zz_22842 = ($signed(_zz_22843) >>> _zz_2185);
  assign _zz_22843 = _zz_22844;
  assign _zz_22844 = ($signed(_zz_22846) + $signed(_zz_2182));
  assign _zz_22845 = ({8'd0,data_mid_52_imag} <<< 8);
  assign _zz_22846 = {{8{_zz_22845[23]}}, _zz_22845};
  assign _zz_22847 = fixTo_2621_dout;
  assign _zz_22848 = ($signed(twiddle_factor_table_116_real) + $signed(twiddle_factor_table_116_imag));
  assign _zz_22849 = ($signed(_zz_2188) - $signed(_zz_22850));
  assign _zz_22850 = ($signed(_zz_22851) * $signed(twiddle_factor_table_116_imag));
  assign _zz_22851 = ($signed(data_mid_117_real) + $signed(data_mid_117_imag));
  assign _zz_22852 = fixTo_2622_dout;
  assign _zz_22853 = ($signed(_zz_2188) + $signed(_zz_22854));
  assign _zz_22854 = ($signed(_zz_22855) * $signed(twiddle_factor_table_116_real));
  assign _zz_22855 = ($signed(data_mid_117_imag) - $signed(data_mid_117_real));
  assign _zz_22856 = fixTo_2623_dout;
  assign _zz_22857 = _zz_22858[31 : 0];
  assign _zz_22858 = _zz_22859;
  assign _zz_22859 = ($signed(_zz_22860) >>> _zz_2189);
  assign _zz_22860 = _zz_22861;
  assign _zz_22861 = ($signed(_zz_22863) - $signed(_zz_2186));
  assign _zz_22862 = ({8'd0,data_mid_53_real} <<< 8);
  assign _zz_22863 = {{8{_zz_22862[23]}}, _zz_22862};
  assign _zz_22864 = fixTo_2624_dout;
  assign _zz_22865 = _zz_22866[31 : 0];
  assign _zz_22866 = _zz_22867;
  assign _zz_22867 = ($signed(_zz_22868) >>> _zz_2189);
  assign _zz_22868 = _zz_22869;
  assign _zz_22869 = ($signed(_zz_22871) - $signed(_zz_2187));
  assign _zz_22870 = ({8'd0,data_mid_53_imag} <<< 8);
  assign _zz_22871 = {{8{_zz_22870[23]}}, _zz_22870};
  assign _zz_22872 = fixTo_2625_dout;
  assign _zz_22873 = _zz_22874[31 : 0];
  assign _zz_22874 = _zz_22875;
  assign _zz_22875 = ($signed(_zz_22876) >>> _zz_2190);
  assign _zz_22876 = _zz_22877;
  assign _zz_22877 = ($signed(_zz_22879) + $signed(_zz_2186));
  assign _zz_22878 = ({8'd0,data_mid_53_real} <<< 8);
  assign _zz_22879 = {{8{_zz_22878[23]}}, _zz_22878};
  assign _zz_22880 = fixTo_2626_dout;
  assign _zz_22881 = _zz_22882[31 : 0];
  assign _zz_22882 = _zz_22883;
  assign _zz_22883 = ($signed(_zz_22884) >>> _zz_2190);
  assign _zz_22884 = _zz_22885;
  assign _zz_22885 = ($signed(_zz_22887) + $signed(_zz_2187));
  assign _zz_22886 = ({8'd0,data_mid_53_imag} <<< 8);
  assign _zz_22887 = {{8{_zz_22886[23]}}, _zz_22886};
  assign _zz_22888 = fixTo_2627_dout;
  assign _zz_22889 = ($signed(twiddle_factor_table_117_real) + $signed(twiddle_factor_table_117_imag));
  assign _zz_22890 = ($signed(_zz_2193) - $signed(_zz_22891));
  assign _zz_22891 = ($signed(_zz_22892) * $signed(twiddle_factor_table_117_imag));
  assign _zz_22892 = ($signed(data_mid_118_real) + $signed(data_mid_118_imag));
  assign _zz_22893 = fixTo_2628_dout;
  assign _zz_22894 = ($signed(_zz_2193) + $signed(_zz_22895));
  assign _zz_22895 = ($signed(_zz_22896) * $signed(twiddle_factor_table_117_real));
  assign _zz_22896 = ($signed(data_mid_118_imag) - $signed(data_mid_118_real));
  assign _zz_22897 = fixTo_2629_dout;
  assign _zz_22898 = _zz_22899[31 : 0];
  assign _zz_22899 = _zz_22900;
  assign _zz_22900 = ($signed(_zz_22901) >>> _zz_2194);
  assign _zz_22901 = _zz_22902;
  assign _zz_22902 = ($signed(_zz_22904) - $signed(_zz_2191));
  assign _zz_22903 = ({8'd0,data_mid_54_real} <<< 8);
  assign _zz_22904 = {{8{_zz_22903[23]}}, _zz_22903};
  assign _zz_22905 = fixTo_2630_dout;
  assign _zz_22906 = _zz_22907[31 : 0];
  assign _zz_22907 = _zz_22908;
  assign _zz_22908 = ($signed(_zz_22909) >>> _zz_2194);
  assign _zz_22909 = _zz_22910;
  assign _zz_22910 = ($signed(_zz_22912) - $signed(_zz_2192));
  assign _zz_22911 = ({8'd0,data_mid_54_imag} <<< 8);
  assign _zz_22912 = {{8{_zz_22911[23]}}, _zz_22911};
  assign _zz_22913 = fixTo_2631_dout;
  assign _zz_22914 = _zz_22915[31 : 0];
  assign _zz_22915 = _zz_22916;
  assign _zz_22916 = ($signed(_zz_22917) >>> _zz_2195);
  assign _zz_22917 = _zz_22918;
  assign _zz_22918 = ($signed(_zz_22920) + $signed(_zz_2191));
  assign _zz_22919 = ({8'd0,data_mid_54_real} <<< 8);
  assign _zz_22920 = {{8{_zz_22919[23]}}, _zz_22919};
  assign _zz_22921 = fixTo_2632_dout;
  assign _zz_22922 = _zz_22923[31 : 0];
  assign _zz_22923 = _zz_22924;
  assign _zz_22924 = ($signed(_zz_22925) >>> _zz_2195);
  assign _zz_22925 = _zz_22926;
  assign _zz_22926 = ($signed(_zz_22928) + $signed(_zz_2192));
  assign _zz_22927 = ({8'd0,data_mid_54_imag} <<< 8);
  assign _zz_22928 = {{8{_zz_22927[23]}}, _zz_22927};
  assign _zz_22929 = fixTo_2633_dout;
  assign _zz_22930 = ($signed(twiddle_factor_table_118_real) + $signed(twiddle_factor_table_118_imag));
  assign _zz_22931 = ($signed(_zz_2198) - $signed(_zz_22932));
  assign _zz_22932 = ($signed(_zz_22933) * $signed(twiddle_factor_table_118_imag));
  assign _zz_22933 = ($signed(data_mid_119_real) + $signed(data_mid_119_imag));
  assign _zz_22934 = fixTo_2634_dout;
  assign _zz_22935 = ($signed(_zz_2198) + $signed(_zz_22936));
  assign _zz_22936 = ($signed(_zz_22937) * $signed(twiddle_factor_table_118_real));
  assign _zz_22937 = ($signed(data_mid_119_imag) - $signed(data_mid_119_real));
  assign _zz_22938 = fixTo_2635_dout;
  assign _zz_22939 = _zz_22940[31 : 0];
  assign _zz_22940 = _zz_22941;
  assign _zz_22941 = ($signed(_zz_22942) >>> _zz_2199);
  assign _zz_22942 = _zz_22943;
  assign _zz_22943 = ($signed(_zz_22945) - $signed(_zz_2196));
  assign _zz_22944 = ({8'd0,data_mid_55_real} <<< 8);
  assign _zz_22945 = {{8{_zz_22944[23]}}, _zz_22944};
  assign _zz_22946 = fixTo_2636_dout;
  assign _zz_22947 = _zz_22948[31 : 0];
  assign _zz_22948 = _zz_22949;
  assign _zz_22949 = ($signed(_zz_22950) >>> _zz_2199);
  assign _zz_22950 = _zz_22951;
  assign _zz_22951 = ($signed(_zz_22953) - $signed(_zz_2197));
  assign _zz_22952 = ({8'd0,data_mid_55_imag} <<< 8);
  assign _zz_22953 = {{8{_zz_22952[23]}}, _zz_22952};
  assign _zz_22954 = fixTo_2637_dout;
  assign _zz_22955 = _zz_22956[31 : 0];
  assign _zz_22956 = _zz_22957;
  assign _zz_22957 = ($signed(_zz_22958) >>> _zz_2200);
  assign _zz_22958 = _zz_22959;
  assign _zz_22959 = ($signed(_zz_22961) + $signed(_zz_2196));
  assign _zz_22960 = ({8'd0,data_mid_55_real} <<< 8);
  assign _zz_22961 = {{8{_zz_22960[23]}}, _zz_22960};
  assign _zz_22962 = fixTo_2638_dout;
  assign _zz_22963 = _zz_22964[31 : 0];
  assign _zz_22964 = _zz_22965;
  assign _zz_22965 = ($signed(_zz_22966) >>> _zz_2200);
  assign _zz_22966 = _zz_22967;
  assign _zz_22967 = ($signed(_zz_22969) + $signed(_zz_2197));
  assign _zz_22968 = ({8'd0,data_mid_55_imag} <<< 8);
  assign _zz_22969 = {{8{_zz_22968[23]}}, _zz_22968};
  assign _zz_22970 = fixTo_2639_dout;
  assign _zz_22971 = ($signed(twiddle_factor_table_119_real) + $signed(twiddle_factor_table_119_imag));
  assign _zz_22972 = ($signed(_zz_2203) - $signed(_zz_22973));
  assign _zz_22973 = ($signed(_zz_22974) * $signed(twiddle_factor_table_119_imag));
  assign _zz_22974 = ($signed(data_mid_120_real) + $signed(data_mid_120_imag));
  assign _zz_22975 = fixTo_2640_dout;
  assign _zz_22976 = ($signed(_zz_2203) + $signed(_zz_22977));
  assign _zz_22977 = ($signed(_zz_22978) * $signed(twiddle_factor_table_119_real));
  assign _zz_22978 = ($signed(data_mid_120_imag) - $signed(data_mid_120_real));
  assign _zz_22979 = fixTo_2641_dout;
  assign _zz_22980 = _zz_22981[31 : 0];
  assign _zz_22981 = _zz_22982;
  assign _zz_22982 = ($signed(_zz_22983) >>> _zz_2204);
  assign _zz_22983 = _zz_22984;
  assign _zz_22984 = ($signed(_zz_22986) - $signed(_zz_2201));
  assign _zz_22985 = ({8'd0,data_mid_56_real} <<< 8);
  assign _zz_22986 = {{8{_zz_22985[23]}}, _zz_22985};
  assign _zz_22987 = fixTo_2642_dout;
  assign _zz_22988 = _zz_22989[31 : 0];
  assign _zz_22989 = _zz_22990;
  assign _zz_22990 = ($signed(_zz_22991) >>> _zz_2204);
  assign _zz_22991 = _zz_22992;
  assign _zz_22992 = ($signed(_zz_22994) - $signed(_zz_2202));
  assign _zz_22993 = ({8'd0,data_mid_56_imag} <<< 8);
  assign _zz_22994 = {{8{_zz_22993[23]}}, _zz_22993};
  assign _zz_22995 = fixTo_2643_dout;
  assign _zz_22996 = _zz_22997[31 : 0];
  assign _zz_22997 = _zz_22998;
  assign _zz_22998 = ($signed(_zz_22999) >>> _zz_2205);
  assign _zz_22999 = _zz_23000;
  assign _zz_23000 = ($signed(_zz_23002) + $signed(_zz_2201));
  assign _zz_23001 = ({8'd0,data_mid_56_real} <<< 8);
  assign _zz_23002 = {{8{_zz_23001[23]}}, _zz_23001};
  assign _zz_23003 = fixTo_2644_dout;
  assign _zz_23004 = _zz_23005[31 : 0];
  assign _zz_23005 = _zz_23006;
  assign _zz_23006 = ($signed(_zz_23007) >>> _zz_2205);
  assign _zz_23007 = _zz_23008;
  assign _zz_23008 = ($signed(_zz_23010) + $signed(_zz_2202));
  assign _zz_23009 = ({8'd0,data_mid_56_imag} <<< 8);
  assign _zz_23010 = {{8{_zz_23009[23]}}, _zz_23009};
  assign _zz_23011 = fixTo_2645_dout;
  assign _zz_23012 = ($signed(twiddle_factor_table_120_real) + $signed(twiddle_factor_table_120_imag));
  assign _zz_23013 = ($signed(_zz_2208) - $signed(_zz_23014));
  assign _zz_23014 = ($signed(_zz_23015) * $signed(twiddle_factor_table_120_imag));
  assign _zz_23015 = ($signed(data_mid_121_real) + $signed(data_mid_121_imag));
  assign _zz_23016 = fixTo_2646_dout;
  assign _zz_23017 = ($signed(_zz_2208) + $signed(_zz_23018));
  assign _zz_23018 = ($signed(_zz_23019) * $signed(twiddle_factor_table_120_real));
  assign _zz_23019 = ($signed(data_mid_121_imag) - $signed(data_mid_121_real));
  assign _zz_23020 = fixTo_2647_dout;
  assign _zz_23021 = _zz_23022[31 : 0];
  assign _zz_23022 = _zz_23023;
  assign _zz_23023 = ($signed(_zz_23024) >>> _zz_2209);
  assign _zz_23024 = _zz_23025;
  assign _zz_23025 = ($signed(_zz_23027) - $signed(_zz_2206));
  assign _zz_23026 = ({8'd0,data_mid_57_real} <<< 8);
  assign _zz_23027 = {{8{_zz_23026[23]}}, _zz_23026};
  assign _zz_23028 = fixTo_2648_dout;
  assign _zz_23029 = _zz_23030[31 : 0];
  assign _zz_23030 = _zz_23031;
  assign _zz_23031 = ($signed(_zz_23032) >>> _zz_2209);
  assign _zz_23032 = _zz_23033;
  assign _zz_23033 = ($signed(_zz_23035) - $signed(_zz_2207));
  assign _zz_23034 = ({8'd0,data_mid_57_imag} <<< 8);
  assign _zz_23035 = {{8{_zz_23034[23]}}, _zz_23034};
  assign _zz_23036 = fixTo_2649_dout;
  assign _zz_23037 = _zz_23038[31 : 0];
  assign _zz_23038 = _zz_23039;
  assign _zz_23039 = ($signed(_zz_23040) >>> _zz_2210);
  assign _zz_23040 = _zz_23041;
  assign _zz_23041 = ($signed(_zz_23043) + $signed(_zz_2206));
  assign _zz_23042 = ({8'd0,data_mid_57_real} <<< 8);
  assign _zz_23043 = {{8{_zz_23042[23]}}, _zz_23042};
  assign _zz_23044 = fixTo_2650_dout;
  assign _zz_23045 = _zz_23046[31 : 0];
  assign _zz_23046 = _zz_23047;
  assign _zz_23047 = ($signed(_zz_23048) >>> _zz_2210);
  assign _zz_23048 = _zz_23049;
  assign _zz_23049 = ($signed(_zz_23051) + $signed(_zz_2207));
  assign _zz_23050 = ({8'd0,data_mid_57_imag} <<< 8);
  assign _zz_23051 = {{8{_zz_23050[23]}}, _zz_23050};
  assign _zz_23052 = fixTo_2651_dout;
  assign _zz_23053 = ($signed(twiddle_factor_table_121_real) + $signed(twiddle_factor_table_121_imag));
  assign _zz_23054 = ($signed(_zz_2213) - $signed(_zz_23055));
  assign _zz_23055 = ($signed(_zz_23056) * $signed(twiddle_factor_table_121_imag));
  assign _zz_23056 = ($signed(data_mid_122_real) + $signed(data_mid_122_imag));
  assign _zz_23057 = fixTo_2652_dout;
  assign _zz_23058 = ($signed(_zz_2213) + $signed(_zz_23059));
  assign _zz_23059 = ($signed(_zz_23060) * $signed(twiddle_factor_table_121_real));
  assign _zz_23060 = ($signed(data_mid_122_imag) - $signed(data_mid_122_real));
  assign _zz_23061 = fixTo_2653_dout;
  assign _zz_23062 = _zz_23063[31 : 0];
  assign _zz_23063 = _zz_23064;
  assign _zz_23064 = ($signed(_zz_23065) >>> _zz_2214);
  assign _zz_23065 = _zz_23066;
  assign _zz_23066 = ($signed(_zz_23068) - $signed(_zz_2211));
  assign _zz_23067 = ({8'd0,data_mid_58_real} <<< 8);
  assign _zz_23068 = {{8{_zz_23067[23]}}, _zz_23067};
  assign _zz_23069 = fixTo_2654_dout;
  assign _zz_23070 = _zz_23071[31 : 0];
  assign _zz_23071 = _zz_23072;
  assign _zz_23072 = ($signed(_zz_23073) >>> _zz_2214);
  assign _zz_23073 = _zz_23074;
  assign _zz_23074 = ($signed(_zz_23076) - $signed(_zz_2212));
  assign _zz_23075 = ({8'd0,data_mid_58_imag} <<< 8);
  assign _zz_23076 = {{8{_zz_23075[23]}}, _zz_23075};
  assign _zz_23077 = fixTo_2655_dout;
  assign _zz_23078 = _zz_23079[31 : 0];
  assign _zz_23079 = _zz_23080;
  assign _zz_23080 = ($signed(_zz_23081) >>> _zz_2215);
  assign _zz_23081 = _zz_23082;
  assign _zz_23082 = ($signed(_zz_23084) + $signed(_zz_2211));
  assign _zz_23083 = ({8'd0,data_mid_58_real} <<< 8);
  assign _zz_23084 = {{8{_zz_23083[23]}}, _zz_23083};
  assign _zz_23085 = fixTo_2656_dout;
  assign _zz_23086 = _zz_23087[31 : 0];
  assign _zz_23087 = _zz_23088;
  assign _zz_23088 = ($signed(_zz_23089) >>> _zz_2215);
  assign _zz_23089 = _zz_23090;
  assign _zz_23090 = ($signed(_zz_23092) + $signed(_zz_2212));
  assign _zz_23091 = ({8'd0,data_mid_58_imag} <<< 8);
  assign _zz_23092 = {{8{_zz_23091[23]}}, _zz_23091};
  assign _zz_23093 = fixTo_2657_dout;
  assign _zz_23094 = ($signed(twiddle_factor_table_122_real) + $signed(twiddle_factor_table_122_imag));
  assign _zz_23095 = ($signed(_zz_2218) - $signed(_zz_23096));
  assign _zz_23096 = ($signed(_zz_23097) * $signed(twiddle_factor_table_122_imag));
  assign _zz_23097 = ($signed(data_mid_123_real) + $signed(data_mid_123_imag));
  assign _zz_23098 = fixTo_2658_dout;
  assign _zz_23099 = ($signed(_zz_2218) + $signed(_zz_23100));
  assign _zz_23100 = ($signed(_zz_23101) * $signed(twiddle_factor_table_122_real));
  assign _zz_23101 = ($signed(data_mid_123_imag) - $signed(data_mid_123_real));
  assign _zz_23102 = fixTo_2659_dout;
  assign _zz_23103 = _zz_23104[31 : 0];
  assign _zz_23104 = _zz_23105;
  assign _zz_23105 = ($signed(_zz_23106) >>> _zz_2219);
  assign _zz_23106 = _zz_23107;
  assign _zz_23107 = ($signed(_zz_23109) - $signed(_zz_2216));
  assign _zz_23108 = ({8'd0,data_mid_59_real} <<< 8);
  assign _zz_23109 = {{8{_zz_23108[23]}}, _zz_23108};
  assign _zz_23110 = fixTo_2660_dout;
  assign _zz_23111 = _zz_23112[31 : 0];
  assign _zz_23112 = _zz_23113;
  assign _zz_23113 = ($signed(_zz_23114) >>> _zz_2219);
  assign _zz_23114 = _zz_23115;
  assign _zz_23115 = ($signed(_zz_23117) - $signed(_zz_2217));
  assign _zz_23116 = ({8'd0,data_mid_59_imag} <<< 8);
  assign _zz_23117 = {{8{_zz_23116[23]}}, _zz_23116};
  assign _zz_23118 = fixTo_2661_dout;
  assign _zz_23119 = _zz_23120[31 : 0];
  assign _zz_23120 = _zz_23121;
  assign _zz_23121 = ($signed(_zz_23122) >>> _zz_2220);
  assign _zz_23122 = _zz_23123;
  assign _zz_23123 = ($signed(_zz_23125) + $signed(_zz_2216));
  assign _zz_23124 = ({8'd0,data_mid_59_real} <<< 8);
  assign _zz_23125 = {{8{_zz_23124[23]}}, _zz_23124};
  assign _zz_23126 = fixTo_2662_dout;
  assign _zz_23127 = _zz_23128[31 : 0];
  assign _zz_23128 = _zz_23129;
  assign _zz_23129 = ($signed(_zz_23130) >>> _zz_2220);
  assign _zz_23130 = _zz_23131;
  assign _zz_23131 = ($signed(_zz_23133) + $signed(_zz_2217));
  assign _zz_23132 = ({8'd0,data_mid_59_imag} <<< 8);
  assign _zz_23133 = {{8{_zz_23132[23]}}, _zz_23132};
  assign _zz_23134 = fixTo_2663_dout;
  assign _zz_23135 = ($signed(twiddle_factor_table_123_real) + $signed(twiddle_factor_table_123_imag));
  assign _zz_23136 = ($signed(_zz_2223) - $signed(_zz_23137));
  assign _zz_23137 = ($signed(_zz_23138) * $signed(twiddle_factor_table_123_imag));
  assign _zz_23138 = ($signed(data_mid_124_real) + $signed(data_mid_124_imag));
  assign _zz_23139 = fixTo_2664_dout;
  assign _zz_23140 = ($signed(_zz_2223) + $signed(_zz_23141));
  assign _zz_23141 = ($signed(_zz_23142) * $signed(twiddle_factor_table_123_real));
  assign _zz_23142 = ($signed(data_mid_124_imag) - $signed(data_mid_124_real));
  assign _zz_23143 = fixTo_2665_dout;
  assign _zz_23144 = _zz_23145[31 : 0];
  assign _zz_23145 = _zz_23146;
  assign _zz_23146 = ($signed(_zz_23147) >>> _zz_2224);
  assign _zz_23147 = _zz_23148;
  assign _zz_23148 = ($signed(_zz_23150) - $signed(_zz_2221));
  assign _zz_23149 = ({8'd0,data_mid_60_real} <<< 8);
  assign _zz_23150 = {{8{_zz_23149[23]}}, _zz_23149};
  assign _zz_23151 = fixTo_2666_dout;
  assign _zz_23152 = _zz_23153[31 : 0];
  assign _zz_23153 = _zz_23154;
  assign _zz_23154 = ($signed(_zz_23155) >>> _zz_2224);
  assign _zz_23155 = _zz_23156;
  assign _zz_23156 = ($signed(_zz_23158) - $signed(_zz_2222));
  assign _zz_23157 = ({8'd0,data_mid_60_imag} <<< 8);
  assign _zz_23158 = {{8{_zz_23157[23]}}, _zz_23157};
  assign _zz_23159 = fixTo_2667_dout;
  assign _zz_23160 = _zz_23161[31 : 0];
  assign _zz_23161 = _zz_23162;
  assign _zz_23162 = ($signed(_zz_23163) >>> _zz_2225);
  assign _zz_23163 = _zz_23164;
  assign _zz_23164 = ($signed(_zz_23166) + $signed(_zz_2221));
  assign _zz_23165 = ({8'd0,data_mid_60_real} <<< 8);
  assign _zz_23166 = {{8{_zz_23165[23]}}, _zz_23165};
  assign _zz_23167 = fixTo_2668_dout;
  assign _zz_23168 = _zz_23169[31 : 0];
  assign _zz_23169 = _zz_23170;
  assign _zz_23170 = ($signed(_zz_23171) >>> _zz_2225);
  assign _zz_23171 = _zz_23172;
  assign _zz_23172 = ($signed(_zz_23174) + $signed(_zz_2222));
  assign _zz_23173 = ({8'd0,data_mid_60_imag} <<< 8);
  assign _zz_23174 = {{8{_zz_23173[23]}}, _zz_23173};
  assign _zz_23175 = fixTo_2669_dout;
  assign _zz_23176 = ($signed(twiddle_factor_table_124_real) + $signed(twiddle_factor_table_124_imag));
  assign _zz_23177 = ($signed(_zz_2228) - $signed(_zz_23178));
  assign _zz_23178 = ($signed(_zz_23179) * $signed(twiddle_factor_table_124_imag));
  assign _zz_23179 = ($signed(data_mid_125_real) + $signed(data_mid_125_imag));
  assign _zz_23180 = fixTo_2670_dout;
  assign _zz_23181 = ($signed(_zz_2228) + $signed(_zz_23182));
  assign _zz_23182 = ($signed(_zz_23183) * $signed(twiddle_factor_table_124_real));
  assign _zz_23183 = ($signed(data_mid_125_imag) - $signed(data_mid_125_real));
  assign _zz_23184 = fixTo_2671_dout;
  assign _zz_23185 = _zz_23186[31 : 0];
  assign _zz_23186 = _zz_23187;
  assign _zz_23187 = ($signed(_zz_23188) >>> _zz_2229);
  assign _zz_23188 = _zz_23189;
  assign _zz_23189 = ($signed(_zz_23191) - $signed(_zz_2226));
  assign _zz_23190 = ({8'd0,data_mid_61_real} <<< 8);
  assign _zz_23191 = {{8{_zz_23190[23]}}, _zz_23190};
  assign _zz_23192 = fixTo_2672_dout;
  assign _zz_23193 = _zz_23194[31 : 0];
  assign _zz_23194 = _zz_23195;
  assign _zz_23195 = ($signed(_zz_23196) >>> _zz_2229);
  assign _zz_23196 = _zz_23197;
  assign _zz_23197 = ($signed(_zz_23199) - $signed(_zz_2227));
  assign _zz_23198 = ({8'd0,data_mid_61_imag} <<< 8);
  assign _zz_23199 = {{8{_zz_23198[23]}}, _zz_23198};
  assign _zz_23200 = fixTo_2673_dout;
  assign _zz_23201 = _zz_23202[31 : 0];
  assign _zz_23202 = _zz_23203;
  assign _zz_23203 = ($signed(_zz_23204) >>> _zz_2230);
  assign _zz_23204 = _zz_23205;
  assign _zz_23205 = ($signed(_zz_23207) + $signed(_zz_2226));
  assign _zz_23206 = ({8'd0,data_mid_61_real} <<< 8);
  assign _zz_23207 = {{8{_zz_23206[23]}}, _zz_23206};
  assign _zz_23208 = fixTo_2674_dout;
  assign _zz_23209 = _zz_23210[31 : 0];
  assign _zz_23210 = _zz_23211;
  assign _zz_23211 = ($signed(_zz_23212) >>> _zz_2230);
  assign _zz_23212 = _zz_23213;
  assign _zz_23213 = ($signed(_zz_23215) + $signed(_zz_2227));
  assign _zz_23214 = ({8'd0,data_mid_61_imag} <<< 8);
  assign _zz_23215 = {{8{_zz_23214[23]}}, _zz_23214};
  assign _zz_23216 = fixTo_2675_dout;
  assign _zz_23217 = ($signed(twiddle_factor_table_125_real) + $signed(twiddle_factor_table_125_imag));
  assign _zz_23218 = ($signed(_zz_2233) - $signed(_zz_23219));
  assign _zz_23219 = ($signed(_zz_23220) * $signed(twiddle_factor_table_125_imag));
  assign _zz_23220 = ($signed(data_mid_126_real) + $signed(data_mid_126_imag));
  assign _zz_23221 = fixTo_2676_dout;
  assign _zz_23222 = ($signed(_zz_2233) + $signed(_zz_23223));
  assign _zz_23223 = ($signed(_zz_23224) * $signed(twiddle_factor_table_125_real));
  assign _zz_23224 = ($signed(data_mid_126_imag) - $signed(data_mid_126_real));
  assign _zz_23225 = fixTo_2677_dout;
  assign _zz_23226 = _zz_23227[31 : 0];
  assign _zz_23227 = _zz_23228;
  assign _zz_23228 = ($signed(_zz_23229) >>> _zz_2234);
  assign _zz_23229 = _zz_23230;
  assign _zz_23230 = ($signed(_zz_23232) - $signed(_zz_2231));
  assign _zz_23231 = ({8'd0,data_mid_62_real} <<< 8);
  assign _zz_23232 = {{8{_zz_23231[23]}}, _zz_23231};
  assign _zz_23233 = fixTo_2678_dout;
  assign _zz_23234 = _zz_23235[31 : 0];
  assign _zz_23235 = _zz_23236;
  assign _zz_23236 = ($signed(_zz_23237) >>> _zz_2234);
  assign _zz_23237 = _zz_23238;
  assign _zz_23238 = ($signed(_zz_23240) - $signed(_zz_2232));
  assign _zz_23239 = ({8'd0,data_mid_62_imag} <<< 8);
  assign _zz_23240 = {{8{_zz_23239[23]}}, _zz_23239};
  assign _zz_23241 = fixTo_2679_dout;
  assign _zz_23242 = _zz_23243[31 : 0];
  assign _zz_23243 = _zz_23244;
  assign _zz_23244 = ($signed(_zz_23245) >>> _zz_2235);
  assign _zz_23245 = _zz_23246;
  assign _zz_23246 = ($signed(_zz_23248) + $signed(_zz_2231));
  assign _zz_23247 = ({8'd0,data_mid_62_real} <<< 8);
  assign _zz_23248 = {{8{_zz_23247[23]}}, _zz_23247};
  assign _zz_23249 = fixTo_2680_dout;
  assign _zz_23250 = _zz_23251[31 : 0];
  assign _zz_23251 = _zz_23252;
  assign _zz_23252 = ($signed(_zz_23253) >>> _zz_2235);
  assign _zz_23253 = _zz_23254;
  assign _zz_23254 = ($signed(_zz_23256) + $signed(_zz_2232));
  assign _zz_23255 = ({8'd0,data_mid_62_imag} <<< 8);
  assign _zz_23256 = {{8{_zz_23255[23]}}, _zz_23255};
  assign _zz_23257 = fixTo_2681_dout;
  assign _zz_23258 = ($signed(twiddle_factor_table_126_real) + $signed(twiddle_factor_table_126_imag));
  assign _zz_23259 = ($signed(_zz_2238) - $signed(_zz_23260));
  assign _zz_23260 = ($signed(_zz_23261) * $signed(twiddle_factor_table_126_imag));
  assign _zz_23261 = ($signed(data_mid_127_real) + $signed(data_mid_127_imag));
  assign _zz_23262 = fixTo_2682_dout;
  assign _zz_23263 = ($signed(_zz_2238) + $signed(_zz_23264));
  assign _zz_23264 = ($signed(_zz_23265) * $signed(twiddle_factor_table_126_real));
  assign _zz_23265 = ($signed(data_mid_127_imag) - $signed(data_mid_127_real));
  assign _zz_23266 = fixTo_2683_dout;
  assign _zz_23267 = _zz_23268[31 : 0];
  assign _zz_23268 = _zz_23269;
  assign _zz_23269 = ($signed(_zz_23270) >>> _zz_2239);
  assign _zz_23270 = _zz_23271;
  assign _zz_23271 = ($signed(_zz_23273) - $signed(_zz_2236));
  assign _zz_23272 = ({8'd0,data_mid_63_real} <<< 8);
  assign _zz_23273 = {{8{_zz_23272[23]}}, _zz_23272};
  assign _zz_23274 = fixTo_2684_dout;
  assign _zz_23275 = _zz_23276[31 : 0];
  assign _zz_23276 = _zz_23277;
  assign _zz_23277 = ($signed(_zz_23278) >>> _zz_2239);
  assign _zz_23278 = _zz_23279;
  assign _zz_23279 = ($signed(_zz_23281) - $signed(_zz_2237));
  assign _zz_23280 = ({8'd0,data_mid_63_imag} <<< 8);
  assign _zz_23281 = {{8{_zz_23280[23]}}, _zz_23280};
  assign _zz_23282 = fixTo_2685_dout;
  assign _zz_23283 = _zz_23284[31 : 0];
  assign _zz_23284 = _zz_23285;
  assign _zz_23285 = ($signed(_zz_23286) >>> _zz_2240);
  assign _zz_23286 = _zz_23287;
  assign _zz_23287 = ($signed(_zz_23289) + $signed(_zz_2236));
  assign _zz_23288 = ({8'd0,data_mid_63_real} <<< 8);
  assign _zz_23289 = {{8{_zz_23288[23]}}, _zz_23288};
  assign _zz_23290 = fixTo_2686_dout;
  assign _zz_23291 = _zz_23292[31 : 0];
  assign _zz_23292 = _zz_23293;
  assign _zz_23293 = ($signed(_zz_23294) >>> _zz_2240);
  assign _zz_23294 = _zz_23295;
  assign _zz_23295 = ($signed(_zz_23297) + $signed(_zz_2237));
  assign _zz_23296 = ({8'd0,data_mid_63_imag} <<< 8);
  assign _zz_23297 = {{8{_zz_23296[23]}}, _zz_23296};
  assign _zz_23298 = fixTo_2687_dout;
  SInt32fixTo31_0_ROUNDTOINF fixTo (
    .din     (_zz_2241[31:0]    ), //i
    .dout    (fixTo_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_1 (
    .din     (_zz_2242[31:0]      ), //i
    .dout    (fixTo_1_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_2 (
    .din     (_zz_2243[31:0]      ), //i
    .dout    (fixTo_2_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_3 (
    .din     (_zz_2244[31:0]      ), //i
    .dout    (fixTo_3_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_4 (
    .din     (_zz_2245[31:0]      ), //i
    .dout    (fixTo_4_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_5 (
    .din     (_zz_2246[31:0]      ), //i
    .dout    (fixTo_5_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_6 (
    .din     (_zz_2247[31:0]      ), //i
    .dout    (fixTo_6_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_7 (
    .din     (_zz_2248[31:0]      ), //i
    .dout    (fixTo_7_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_8 (
    .din     (_zz_2249[31:0]      ), //i
    .dout    (fixTo_8_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_9 (
    .din     (_zz_2250[31:0]      ), //i
    .dout    (fixTo_9_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_10 (
    .din     (_zz_2251[31:0]       ), //i
    .dout    (fixTo_10_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_11 (
    .din     (_zz_2252[31:0]       ), //i
    .dout    (fixTo_11_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_12 (
    .din     (_zz_2253[31:0]       ), //i
    .dout    (fixTo_12_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_13 (
    .din     (_zz_2254[31:0]       ), //i
    .dout    (fixTo_13_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_14 (
    .din     (_zz_2255[31:0]       ), //i
    .dout    (fixTo_14_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_15 (
    .din     (_zz_2256[31:0]       ), //i
    .dout    (fixTo_15_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_16 (
    .din     (_zz_2257[31:0]       ), //i
    .dout    (fixTo_16_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_17 (
    .din     (_zz_2258[31:0]       ), //i
    .dout    (fixTo_17_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_18 (
    .din     (_zz_2259[31:0]       ), //i
    .dout    (fixTo_18_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_19 (
    .din     (_zz_2260[31:0]       ), //i
    .dout    (fixTo_19_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_20 (
    .din     (_zz_2261[31:0]       ), //i
    .dout    (fixTo_20_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_21 (
    .din     (_zz_2262[31:0]       ), //i
    .dout    (fixTo_21_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_22 (
    .din     (_zz_2263[31:0]       ), //i
    .dout    (fixTo_22_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_23 (
    .din     (_zz_2264[31:0]       ), //i
    .dout    (fixTo_23_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_24 (
    .din     (_zz_2265[31:0]       ), //i
    .dout    (fixTo_24_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_25 (
    .din     (_zz_2266[31:0]       ), //i
    .dout    (fixTo_25_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_26 (
    .din     (_zz_2267[31:0]       ), //i
    .dout    (fixTo_26_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_27 (
    .din     (_zz_2268[31:0]       ), //i
    .dout    (fixTo_27_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_28 (
    .din     (_zz_2269[31:0]       ), //i
    .dout    (fixTo_28_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_29 (
    .din     (_zz_2270[31:0]       ), //i
    .dout    (fixTo_29_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_30 (
    .din     (_zz_2271[31:0]       ), //i
    .dout    (fixTo_30_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_31 (
    .din     (_zz_2272[31:0]       ), //i
    .dout    (fixTo_31_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_32 (
    .din     (_zz_2273[31:0]       ), //i
    .dout    (fixTo_32_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_33 (
    .din     (_zz_2274[31:0]       ), //i
    .dout    (fixTo_33_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_34 (
    .din     (_zz_2275[31:0]       ), //i
    .dout    (fixTo_34_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_35 (
    .din     (_zz_2276[31:0]       ), //i
    .dout    (fixTo_35_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_36 (
    .din     (_zz_2277[31:0]       ), //i
    .dout    (fixTo_36_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_37 (
    .din     (_zz_2278[31:0]       ), //i
    .dout    (fixTo_37_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_38 (
    .din     (_zz_2279[31:0]       ), //i
    .dout    (fixTo_38_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_39 (
    .din     (_zz_2280[31:0]       ), //i
    .dout    (fixTo_39_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_40 (
    .din     (_zz_2281[31:0]       ), //i
    .dout    (fixTo_40_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_41 (
    .din     (_zz_2282[31:0]       ), //i
    .dout    (fixTo_41_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_42 (
    .din     (_zz_2283[31:0]       ), //i
    .dout    (fixTo_42_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_43 (
    .din     (_zz_2284[31:0]       ), //i
    .dout    (fixTo_43_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_44 (
    .din     (_zz_2285[31:0]       ), //i
    .dout    (fixTo_44_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_45 (
    .din     (_zz_2286[31:0]       ), //i
    .dout    (fixTo_45_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_46 (
    .din     (_zz_2287[31:0]       ), //i
    .dout    (fixTo_46_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_47 (
    .din     (_zz_2288[31:0]       ), //i
    .dout    (fixTo_47_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_48 (
    .din     (_zz_2289[31:0]       ), //i
    .dout    (fixTo_48_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_49 (
    .din     (_zz_2290[31:0]       ), //i
    .dout    (fixTo_49_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_50 (
    .din     (_zz_2291[31:0]       ), //i
    .dout    (fixTo_50_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_51 (
    .din     (_zz_2292[31:0]       ), //i
    .dout    (fixTo_51_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_52 (
    .din     (_zz_2293[31:0]       ), //i
    .dout    (fixTo_52_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_53 (
    .din     (_zz_2294[31:0]       ), //i
    .dout    (fixTo_53_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_54 (
    .din     (_zz_2295[31:0]       ), //i
    .dout    (fixTo_54_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_55 (
    .din     (_zz_2296[31:0]       ), //i
    .dout    (fixTo_55_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_56 (
    .din     (_zz_2297[31:0]       ), //i
    .dout    (fixTo_56_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_57 (
    .din     (_zz_2298[31:0]       ), //i
    .dout    (fixTo_57_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_58 (
    .din     (_zz_2299[31:0]       ), //i
    .dout    (fixTo_58_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_59 (
    .din     (_zz_2300[31:0]       ), //i
    .dout    (fixTo_59_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_60 (
    .din     (_zz_2301[31:0]       ), //i
    .dout    (fixTo_60_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_61 (
    .din     (_zz_2302[31:0]       ), //i
    .dout    (fixTo_61_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_62 (
    .din     (_zz_2303[31:0]       ), //i
    .dout    (fixTo_62_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_63 (
    .din     (_zz_2304[31:0]       ), //i
    .dout    (fixTo_63_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_64 (
    .din     (_zz_2305[31:0]       ), //i
    .dout    (fixTo_64_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_65 (
    .din     (_zz_2306[31:0]       ), //i
    .dout    (fixTo_65_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_66 (
    .din     (_zz_2307[31:0]       ), //i
    .dout    (fixTo_66_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_67 (
    .din     (_zz_2308[31:0]       ), //i
    .dout    (fixTo_67_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_68 (
    .din     (_zz_2309[31:0]       ), //i
    .dout    (fixTo_68_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_69 (
    .din     (_zz_2310[31:0]       ), //i
    .dout    (fixTo_69_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_70 (
    .din     (_zz_2311[31:0]       ), //i
    .dout    (fixTo_70_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_71 (
    .din     (_zz_2312[31:0]       ), //i
    .dout    (fixTo_71_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_72 (
    .din     (_zz_2313[31:0]       ), //i
    .dout    (fixTo_72_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_73 (
    .din     (_zz_2314[31:0]       ), //i
    .dout    (fixTo_73_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_74 (
    .din     (_zz_2315[31:0]       ), //i
    .dout    (fixTo_74_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_75 (
    .din     (_zz_2316[31:0]       ), //i
    .dout    (fixTo_75_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_76 (
    .din     (_zz_2317[31:0]       ), //i
    .dout    (fixTo_76_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_77 (
    .din     (_zz_2318[31:0]       ), //i
    .dout    (fixTo_77_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_78 (
    .din     (_zz_2319[31:0]       ), //i
    .dout    (fixTo_78_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_79 (
    .din     (_zz_2320[31:0]       ), //i
    .dout    (fixTo_79_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_80 (
    .din     (_zz_2321[31:0]       ), //i
    .dout    (fixTo_80_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_81 (
    .din     (_zz_2322[31:0]       ), //i
    .dout    (fixTo_81_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_82 (
    .din     (_zz_2323[31:0]       ), //i
    .dout    (fixTo_82_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_83 (
    .din     (_zz_2324[31:0]       ), //i
    .dout    (fixTo_83_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_84 (
    .din     (_zz_2325[31:0]       ), //i
    .dout    (fixTo_84_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_85 (
    .din     (_zz_2326[31:0]       ), //i
    .dout    (fixTo_85_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_86 (
    .din     (_zz_2327[31:0]       ), //i
    .dout    (fixTo_86_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_87 (
    .din     (_zz_2328[31:0]       ), //i
    .dout    (fixTo_87_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_88 (
    .din     (_zz_2329[31:0]       ), //i
    .dout    (fixTo_88_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_89 (
    .din     (_zz_2330[31:0]       ), //i
    .dout    (fixTo_89_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_90 (
    .din     (_zz_2331[31:0]       ), //i
    .dout    (fixTo_90_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_91 (
    .din     (_zz_2332[31:0]       ), //i
    .dout    (fixTo_91_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_92 (
    .din     (_zz_2333[31:0]       ), //i
    .dout    (fixTo_92_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_93 (
    .din     (_zz_2334[31:0]       ), //i
    .dout    (fixTo_93_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_94 (
    .din     (_zz_2335[31:0]       ), //i
    .dout    (fixTo_94_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_95 (
    .din     (_zz_2336[31:0]       ), //i
    .dout    (fixTo_95_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_96 (
    .din     (_zz_2337[31:0]       ), //i
    .dout    (fixTo_96_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_97 (
    .din     (_zz_2338[31:0]       ), //i
    .dout    (fixTo_97_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_98 (
    .din     (_zz_2339[31:0]       ), //i
    .dout    (fixTo_98_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_99 (
    .din     (_zz_2340[31:0]       ), //i
    .dout    (fixTo_99_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_100 (
    .din     (_zz_2341[31:0]        ), //i
    .dout    (fixTo_100_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_101 (
    .din     (_zz_2342[31:0]        ), //i
    .dout    (fixTo_101_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_102 (
    .din     (_zz_2343[31:0]        ), //i
    .dout    (fixTo_102_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_103 (
    .din     (_zz_2344[31:0]        ), //i
    .dout    (fixTo_103_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_104 (
    .din     (_zz_2345[31:0]        ), //i
    .dout    (fixTo_104_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_105 (
    .din     (_zz_2346[31:0]        ), //i
    .dout    (fixTo_105_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_106 (
    .din     (_zz_2347[31:0]        ), //i
    .dout    (fixTo_106_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_107 (
    .din     (_zz_2348[31:0]        ), //i
    .dout    (fixTo_107_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_108 (
    .din     (_zz_2349[31:0]        ), //i
    .dout    (fixTo_108_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_109 (
    .din     (_zz_2350[31:0]        ), //i
    .dout    (fixTo_109_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_110 (
    .din     (_zz_2351[31:0]        ), //i
    .dout    (fixTo_110_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_111 (
    .din     (_zz_2352[31:0]        ), //i
    .dout    (fixTo_111_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_112 (
    .din     (_zz_2353[31:0]        ), //i
    .dout    (fixTo_112_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_113 (
    .din     (_zz_2354[31:0]        ), //i
    .dout    (fixTo_113_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_114 (
    .din     (_zz_2355[31:0]        ), //i
    .dout    (fixTo_114_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_115 (
    .din     (_zz_2356[31:0]        ), //i
    .dout    (fixTo_115_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_116 (
    .din     (_zz_2357[31:0]        ), //i
    .dout    (fixTo_116_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_117 (
    .din     (_zz_2358[31:0]        ), //i
    .dout    (fixTo_117_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_118 (
    .din     (_zz_2359[31:0]        ), //i
    .dout    (fixTo_118_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_119 (
    .din     (_zz_2360[31:0]        ), //i
    .dout    (fixTo_119_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_120 (
    .din     (_zz_2361[31:0]        ), //i
    .dout    (fixTo_120_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_121 (
    .din     (_zz_2362[31:0]        ), //i
    .dout    (fixTo_121_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_122 (
    .din     (_zz_2363[31:0]        ), //i
    .dout    (fixTo_122_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_123 (
    .din     (_zz_2364[31:0]        ), //i
    .dout    (fixTo_123_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_124 (
    .din     (_zz_2365[31:0]        ), //i
    .dout    (fixTo_124_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_125 (
    .din     (_zz_2366[31:0]        ), //i
    .dout    (fixTo_125_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_126 (
    .din     (_zz_2367[31:0]        ), //i
    .dout    (fixTo_126_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_127 (
    .din     (_zz_2368[31:0]        ), //i
    .dout    (fixTo_127_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_128 (
    .din     (_zz_2369[31:0]        ), //i
    .dout    (fixTo_128_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_129 (
    .din     (_zz_2370[31:0]        ), //i
    .dout    (fixTo_129_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_130 (
    .din     (_zz_2371[31:0]        ), //i
    .dout    (fixTo_130_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_131 (
    .din     (_zz_2372[31:0]        ), //i
    .dout    (fixTo_131_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_132 (
    .din     (_zz_2373[31:0]        ), //i
    .dout    (fixTo_132_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_133 (
    .din     (_zz_2374[31:0]        ), //i
    .dout    (fixTo_133_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_134 (
    .din     (_zz_2375[31:0]        ), //i
    .dout    (fixTo_134_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_135 (
    .din     (_zz_2376[31:0]        ), //i
    .dout    (fixTo_135_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_136 (
    .din     (_zz_2377[31:0]        ), //i
    .dout    (fixTo_136_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_137 (
    .din     (_zz_2378[31:0]        ), //i
    .dout    (fixTo_137_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_138 (
    .din     (_zz_2379[31:0]        ), //i
    .dout    (fixTo_138_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_139 (
    .din     (_zz_2380[31:0]        ), //i
    .dout    (fixTo_139_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_140 (
    .din     (_zz_2381[31:0]        ), //i
    .dout    (fixTo_140_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_141 (
    .din     (_zz_2382[31:0]        ), //i
    .dout    (fixTo_141_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_142 (
    .din     (_zz_2383[31:0]        ), //i
    .dout    (fixTo_142_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_143 (
    .din     (_zz_2384[31:0]        ), //i
    .dout    (fixTo_143_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_144 (
    .din     (_zz_2385[31:0]        ), //i
    .dout    (fixTo_144_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_145 (
    .din     (_zz_2386[31:0]        ), //i
    .dout    (fixTo_145_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_146 (
    .din     (_zz_2387[31:0]        ), //i
    .dout    (fixTo_146_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_147 (
    .din     (_zz_2388[31:0]        ), //i
    .dout    (fixTo_147_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_148 (
    .din     (_zz_2389[31:0]        ), //i
    .dout    (fixTo_148_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_149 (
    .din     (_zz_2390[31:0]        ), //i
    .dout    (fixTo_149_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_150 (
    .din     (_zz_2391[31:0]        ), //i
    .dout    (fixTo_150_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_151 (
    .din     (_zz_2392[31:0]        ), //i
    .dout    (fixTo_151_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_152 (
    .din     (_zz_2393[31:0]        ), //i
    .dout    (fixTo_152_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_153 (
    .din     (_zz_2394[31:0]        ), //i
    .dout    (fixTo_153_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_154 (
    .din     (_zz_2395[31:0]        ), //i
    .dout    (fixTo_154_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_155 (
    .din     (_zz_2396[31:0]        ), //i
    .dout    (fixTo_155_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_156 (
    .din     (_zz_2397[31:0]        ), //i
    .dout    (fixTo_156_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_157 (
    .din     (_zz_2398[31:0]        ), //i
    .dout    (fixTo_157_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_158 (
    .din     (_zz_2399[31:0]        ), //i
    .dout    (fixTo_158_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_159 (
    .din     (_zz_2400[31:0]        ), //i
    .dout    (fixTo_159_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_160 (
    .din     (_zz_2401[31:0]        ), //i
    .dout    (fixTo_160_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_161 (
    .din     (_zz_2402[31:0]        ), //i
    .dout    (fixTo_161_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_162 (
    .din     (_zz_2403[31:0]        ), //i
    .dout    (fixTo_162_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_163 (
    .din     (_zz_2404[31:0]        ), //i
    .dout    (fixTo_163_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_164 (
    .din     (_zz_2405[31:0]        ), //i
    .dout    (fixTo_164_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_165 (
    .din     (_zz_2406[31:0]        ), //i
    .dout    (fixTo_165_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_166 (
    .din     (_zz_2407[31:0]        ), //i
    .dout    (fixTo_166_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_167 (
    .din     (_zz_2408[31:0]        ), //i
    .dout    (fixTo_167_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_168 (
    .din     (_zz_2409[31:0]        ), //i
    .dout    (fixTo_168_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_169 (
    .din     (_zz_2410[31:0]        ), //i
    .dout    (fixTo_169_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_170 (
    .din     (_zz_2411[31:0]        ), //i
    .dout    (fixTo_170_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_171 (
    .din     (_zz_2412[31:0]        ), //i
    .dout    (fixTo_171_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_172 (
    .din     (_zz_2413[31:0]        ), //i
    .dout    (fixTo_172_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_173 (
    .din     (_zz_2414[31:0]        ), //i
    .dout    (fixTo_173_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_174 (
    .din     (_zz_2415[31:0]        ), //i
    .dout    (fixTo_174_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_175 (
    .din     (_zz_2416[31:0]        ), //i
    .dout    (fixTo_175_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_176 (
    .din     (_zz_2417[31:0]        ), //i
    .dout    (fixTo_176_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_177 (
    .din     (_zz_2418[31:0]        ), //i
    .dout    (fixTo_177_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_178 (
    .din     (_zz_2419[31:0]        ), //i
    .dout    (fixTo_178_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_179 (
    .din     (_zz_2420[31:0]        ), //i
    .dout    (fixTo_179_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_180 (
    .din     (_zz_2421[31:0]        ), //i
    .dout    (fixTo_180_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_181 (
    .din     (_zz_2422[31:0]        ), //i
    .dout    (fixTo_181_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_182 (
    .din     (_zz_2423[31:0]        ), //i
    .dout    (fixTo_182_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_183 (
    .din     (_zz_2424[31:0]        ), //i
    .dout    (fixTo_183_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_184 (
    .din     (_zz_2425[31:0]        ), //i
    .dout    (fixTo_184_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_185 (
    .din     (_zz_2426[31:0]        ), //i
    .dout    (fixTo_185_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_186 (
    .din     (_zz_2427[31:0]        ), //i
    .dout    (fixTo_186_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_187 (
    .din     (_zz_2428[31:0]        ), //i
    .dout    (fixTo_187_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_188 (
    .din     (_zz_2429[31:0]        ), //i
    .dout    (fixTo_188_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_189 (
    .din     (_zz_2430[31:0]        ), //i
    .dout    (fixTo_189_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_190 (
    .din     (_zz_2431[31:0]        ), //i
    .dout    (fixTo_190_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_191 (
    .din     (_zz_2432[31:0]        ), //i
    .dout    (fixTo_191_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_192 (
    .din     (_zz_2433[31:0]        ), //i
    .dout    (fixTo_192_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_193 (
    .din     (_zz_2434[31:0]        ), //i
    .dout    (fixTo_193_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_194 (
    .din     (_zz_2435[31:0]        ), //i
    .dout    (fixTo_194_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_195 (
    .din     (_zz_2436[31:0]        ), //i
    .dout    (fixTo_195_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_196 (
    .din     (_zz_2437[31:0]        ), //i
    .dout    (fixTo_196_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_197 (
    .din     (_zz_2438[31:0]        ), //i
    .dout    (fixTo_197_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_198 (
    .din     (_zz_2439[31:0]        ), //i
    .dout    (fixTo_198_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_199 (
    .din     (_zz_2440[31:0]        ), //i
    .dout    (fixTo_199_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_200 (
    .din     (_zz_2441[31:0]        ), //i
    .dout    (fixTo_200_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_201 (
    .din     (_zz_2442[31:0]        ), //i
    .dout    (fixTo_201_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_202 (
    .din     (_zz_2443[31:0]        ), //i
    .dout    (fixTo_202_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_203 (
    .din     (_zz_2444[31:0]        ), //i
    .dout    (fixTo_203_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_204 (
    .din     (_zz_2445[31:0]        ), //i
    .dout    (fixTo_204_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_205 (
    .din     (_zz_2446[31:0]        ), //i
    .dout    (fixTo_205_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_206 (
    .din     (_zz_2447[31:0]        ), //i
    .dout    (fixTo_206_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_207 (
    .din     (_zz_2448[31:0]        ), //i
    .dout    (fixTo_207_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_208 (
    .din     (_zz_2449[31:0]        ), //i
    .dout    (fixTo_208_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_209 (
    .din     (_zz_2450[31:0]        ), //i
    .dout    (fixTo_209_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_210 (
    .din     (_zz_2451[31:0]        ), //i
    .dout    (fixTo_210_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_211 (
    .din     (_zz_2452[31:0]        ), //i
    .dout    (fixTo_211_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_212 (
    .din     (_zz_2453[31:0]        ), //i
    .dout    (fixTo_212_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_213 (
    .din     (_zz_2454[31:0]        ), //i
    .dout    (fixTo_213_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_214 (
    .din     (_zz_2455[31:0]        ), //i
    .dout    (fixTo_214_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_215 (
    .din     (_zz_2456[31:0]        ), //i
    .dout    (fixTo_215_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_216 (
    .din     (_zz_2457[31:0]        ), //i
    .dout    (fixTo_216_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_217 (
    .din     (_zz_2458[31:0]        ), //i
    .dout    (fixTo_217_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_218 (
    .din     (_zz_2459[31:0]        ), //i
    .dout    (fixTo_218_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_219 (
    .din     (_zz_2460[31:0]        ), //i
    .dout    (fixTo_219_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_220 (
    .din     (_zz_2461[31:0]        ), //i
    .dout    (fixTo_220_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_221 (
    .din     (_zz_2462[31:0]        ), //i
    .dout    (fixTo_221_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_222 (
    .din     (_zz_2463[31:0]        ), //i
    .dout    (fixTo_222_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_223 (
    .din     (_zz_2464[31:0]        ), //i
    .dout    (fixTo_223_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_224 (
    .din     (_zz_2465[31:0]        ), //i
    .dout    (fixTo_224_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_225 (
    .din     (_zz_2466[31:0]        ), //i
    .dout    (fixTo_225_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_226 (
    .din     (_zz_2467[31:0]        ), //i
    .dout    (fixTo_226_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_227 (
    .din     (_zz_2468[31:0]        ), //i
    .dout    (fixTo_227_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_228 (
    .din     (_zz_2469[31:0]        ), //i
    .dout    (fixTo_228_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_229 (
    .din     (_zz_2470[31:0]        ), //i
    .dout    (fixTo_229_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_230 (
    .din     (_zz_2471[31:0]        ), //i
    .dout    (fixTo_230_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_231 (
    .din     (_zz_2472[31:0]        ), //i
    .dout    (fixTo_231_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_232 (
    .din     (_zz_2473[31:0]        ), //i
    .dout    (fixTo_232_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_233 (
    .din     (_zz_2474[31:0]        ), //i
    .dout    (fixTo_233_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_234 (
    .din     (_zz_2475[31:0]        ), //i
    .dout    (fixTo_234_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_235 (
    .din     (_zz_2476[31:0]        ), //i
    .dout    (fixTo_235_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_236 (
    .din     (_zz_2477[31:0]        ), //i
    .dout    (fixTo_236_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_237 (
    .din     (_zz_2478[31:0]        ), //i
    .dout    (fixTo_237_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_238 (
    .din     (_zz_2479[31:0]        ), //i
    .dout    (fixTo_238_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_239 (
    .din     (_zz_2480[31:0]        ), //i
    .dout    (fixTo_239_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_240 (
    .din     (_zz_2481[31:0]        ), //i
    .dout    (fixTo_240_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_241 (
    .din     (_zz_2482[31:0]        ), //i
    .dout    (fixTo_241_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_242 (
    .din     (_zz_2483[31:0]        ), //i
    .dout    (fixTo_242_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_243 (
    .din     (_zz_2484[31:0]        ), //i
    .dout    (fixTo_243_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_244 (
    .din     (_zz_2485[31:0]        ), //i
    .dout    (fixTo_244_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_245 (
    .din     (_zz_2486[31:0]        ), //i
    .dout    (fixTo_245_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_246 (
    .din     (_zz_2487[31:0]        ), //i
    .dout    (fixTo_246_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_247 (
    .din     (_zz_2488[31:0]        ), //i
    .dout    (fixTo_247_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_248 (
    .din     (_zz_2489[31:0]        ), //i
    .dout    (fixTo_248_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_249 (
    .din     (_zz_2490[31:0]        ), //i
    .dout    (fixTo_249_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_250 (
    .din     (_zz_2491[31:0]        ), //i
    .dout    (fixTo_250_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_251 (
    .din     (_zz_2492[31:0]        ), //i
    .dout    (fixTo_251_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_252 (
    .din     (_zz_2493[31:0]        ), //i
    .dout    (fixTo_252_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_253 (
    .din     (_zz_2494[31:0]        ), //i
    .dout    (fixTo_253_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_254 (
    .din     (_zz_2495[31:0]        ), //i
    .dout    (fixTo_254_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_255 (
    .din     (_zz_2496[31:0]        ), //i
    .dout    (fixTo_255_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_256 (
    .din     (_zz_2497[31:0]        ), //i
    .dout    (fixTo_256_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_257 (
    .din     (_zz_2498[31:0]        ), //i
    .dout    (fixTo_257_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_258 (
    .din     (_zz_2499[31:0]        ), //i
    .dout    (fixTo_258_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_259 (
    .din     (_zz_2500[31:0]        ), //i
    .dout    (fixTo_259_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_260 (
    .din     (_zz_2501[31:0]        ), //i
    .dout    (fixTo_260_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_261 (
    .din     (_zz_2502[31:0]        ), //i
    .dout    (fixTo_261_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_262 (
    .din     (_zz_2503[31:0]        ), //i
    .dout    (fixTo_262_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_263 (
    .din     (_zz_2504[31:0]        ), //i
    .dout    (fixTo_263_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_264 (
    .din     (_zz_2505[31:0]        ), //i
    .dout    (fixTo_264_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_265 (
    .din     (_zz_2506[31:0]        ), //i
    .dout    (fixTo_265_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_266 (
    .din     (_zz_2507[31:0]        ), //i
    .dout    (fixTo_266_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_267 (
    .din     (_zz_2508[31:0]        ), //i
    .dout    (fixTo_267_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_268 (
    .din     (_zz_2509[31:0]        ), //i
    .dout    (fixTo_268_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_269 (
    .din     (_zz_2510[31:0]        ), //i
    .dout    (fixTo_269_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_270 (
    .din     (_zz_2511[31:0]        ), //i
    .dout    (fixTo_270_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_271 (
    .din     (_zz_2512[31:0]        ), //i
    .dout    (fixTo_271_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_272 (
    .din     (_zz_2513[31:0]        ), //i
    .dout    (fixTo_272_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_273 (
    .din     (_zz_2514[31:0]        ), //i
    .dout    (fixTo_273_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_274 (
    .din     (_zz_2515[31:0]        ), //i
    .dout    (fixTo_274_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_275 (
    .din     (_zz_2516[31:0]        ), //i
    .dout    (fixTo_275_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_276 (
    .din     (_zz_2517[31:0]        ), //i
    .dout    (fixTo_276_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_277 (
    .din     (_zz_2518[31:0]        ), //i
    .dout    (fixTo_277_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_278 (
    .din     (_zz_2519[31:0]        ), //i
    .dout    (fixTo_278_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_279 (
    .din     (_zz_2520[31:0]        ), //i
    .dout    (fixTo_279_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_280 (
    .din     (_zz_2521[31:0]        ), //i
    .dout    (fixTo_280_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_281 (
    .din     (_zz_2522[31:0]        ), //i
    .dout    (fixTo_281_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_282 (
    .din     (_zz_2523[31:0]        ), //i
    .dout    (fixTo_282_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_283 (
    .din     (_zz_2524[31:0]        ), //i
    .dout    (fixTo_283_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_284 (
    .din     (_zz_2525[31:0]        ), //i
    .dout    (fixTo_284_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_285 (
    .din     (_zz_2526[31:0]        ), //i
    .dout    (fixTo_285_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_286 (
    .din     (_zz_2527[31:0]        ), //i
    .dout    (fixTo_286_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_287 (
    .din     (_zz_2528[31:0]        ), //i
    .dout    (fixTo_287_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_288 (
    .din     (_zz_2529[31:0]        ), //i
    .dout    (fixTo_288_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_289 (
    .din     (_zz_2530[31:0]        ), //i
    .dout    (fixTo_289_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_290 (
    .din     (_zz_2531[31:0]        ), //i
    .dout    (fixTo_290_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_291 (
    .din     (_zz_2532[31:0]        ), //i
    .dout    (fixTo_291_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_292 (
    .din     (_zz_2533[31:0]        ), //i
    .dout    (fixTo_292_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_293 (
    .din     (_zz_2534[31:0]        ), //i
    .dout    (fixTo_293_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_294 (
    .din     (_zz_2535[31:0]        ), //i
    .dout    (fixTo_294_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_295 (
    .din     (_zz_2536[31:0]        ), //i
    .dout    (fixTo_295_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_296 (
    .din     (_zz_2537[31:0]        ), //i
    .dout    (fixTo_296_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_297 (
    .din     (_zz_2538[31:0]        ), //i
    .dout    (fixTo_297_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_298 (
    .din     (_zz_2539[31:0]        ), //i
    .dout    (fixTo_298_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_299 (
    .din     (_zz_2540[31:0]        ), //i
    .dout    (fixTo_299_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_300 (
    .din     (_zz_2541[31:0]        ), //i
    .dout    (fixTo_300_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_301 (
    .din     (_zz_2542[31:0]        ), //i
    .dout    (fixTo_301_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_302 (
    .din     (_zz_2543[31:0]        ), //i
    .dout    (fixTo_302_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_303 (
    .din     (_zz_2544[31:0]        ), //i
    .dout    (fixTo_303_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_304 (
    .din     (_zz_2545[31:0]        ), //i
    .dout    (fixTo_304_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_305 (
    .din     (_zz_2546[31:0]        ), //i
    .dout    (fixTo_305_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_306 (
    .din     (_zz_2547[31:0]        ), //i
    .dout    (fixTo_306_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_307 (
    .din     (_zz_2548[31:0]        ), //i
    .dout    (fixTo_307_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_308 (
    .din     (_zz_2549[31:0]        ), //i
    .dout    (fixTo_308_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_309 (
    .din     (_zz_2550[31:0]        ), //i
    .dout    (fixTo_309_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_310 (
    .din     (_zz_2551[31:0]        ), //i
    .dout    (fixTo_310_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_311 (
    .din     (_zz_2552[31:0]        ), //i
    .dout    (fixTo_311_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_312 (
    .din     (_zz_2553[31:0]        ), //i
    .dout    (fixTo_312_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_313 (
    .din     (_zz_2554[31:0]        ), //i
    .dout    (fixTo_313_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_314 (
    .din     (_zz_2555[31:0]        ), //i
    .dout    (fixTo_314_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_315 (
    .din     (_zz_2556[31:0]        ), //i
    .dout    (fixTo_315_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_316 (
    .din     (_zz_2557[31:0]        ), //i
    .dout    (fixTo_316_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_317 (
    .din     (_zz_2558[31:0]        ), //i
    .dout    (fixTo_317_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_318 (
    .din     (_zz_2559[31:0]        ), //i
    .dout    (fixTo_318_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_319 (
    .din     (_zz_2560[31:0]        ), //i
    .dout    (fixTo_319_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_320 (
    .din     (_zz_2561[31:0]        ), //i
    .dout    (fixTo_320_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_321 (
    .din     (_zz_2562[31:0]        ), //i
    .dout    (fixTo_321_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_322 (
    .din     (_zz_2563[31:0]        ), //i
    .dout    (fixTo_322_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_323 (
    .din     (_zz_2564[31:0]        ), //i
    .dout    (fixTo_323_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_324 (
    .din     (_zz_2565[31:0]        ), //i
    .dout    (fixTo_324_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_325 (
    .din     (_zz_2566[31:0]        ), //i
    .dout    (fixTo_325_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_326 (
    .din     (_zz_2567[31:0]        ), //i
    .dout    (fixTo_326_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_327 (
    .din     (_zz_2568[31:0]        ), //i
    .dout    (fixTo_327_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_328 (
    .din     (_zz_2569[31:0]        ), //i
    .dout    (fixTo_328_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_329 (
    .din     (_zz_2570[31:0]        ), //i
    .dout    (fixTo_329_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_330 (
    .din     (_zz_2571[31:0]        ), //i
    .dout    (fixTo_330_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_331 (
    .din     (_zz_2572[31:0]        ), //i
    .dout    (fixTo_331_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_332 (
    .din     (_zz_2573[31:0]        ), //i
    .dout    (fixTo_332_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_333 (
    .din     (_zz_2574[31:0]        ), //i
    .dout    (fixTo_333_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_334 (
    .din     (_zz_2575[31:0]        ), //i
    .dout    (fixTo_334_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_335 (
    .din     (_zz_2576[31:0]        ), //i
    .dout    (fixTo_335_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_336 (
    .din     (_zz_2577[31:0]        ), //i
    .dout    (fixTo_336_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_337 (
    .din     (_zz_2578[31:0]        ), //i
    .dout    (fixTo_337_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_338 (
    .din     (_zz_2579[31:0]        ), //i
    .dout    (fixTo_338_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_339 (
    .din     (_zz_2580[31:0]        ), //i
    .dout    (fixTo_339_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_340 (
    .din     (_zz_2581[31:0]        ), //i
    .dout    (fixTo_340_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_341 (
    .din     (_zz_2582[31:0]        ), //i
    .dout    (fixTo_341_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_342 (
    .din     (_zz_2583[31:0]        ), //i
    .dout    (fixTo_342_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_343 (
    .din     (_zz_2584[31:0]        ), //i
    .dout    (fixTo_343_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_344 (
    .din     (_zz_2585[31:0]        ), //i
    .dout    (fixTo_344_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_345 (
    .din     (_zz_2586[31:0]        ), //i
    .dout    (fixTo_345_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_346 (
    .din     (_zz_2587[31:0]        ), //i
    .dout    (fixTo_346_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_347 (
    .din     (_zz_2588[31:0]        ), //i
    .dout    (fixTo_347_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_348 (
    .din     (_zz_2589[31:0]        ), //i
    .dout    (fixTo_348_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_349 (
    .din     (_zz_2590[31:0]        ), //i
    .dout    (fixTo_349_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_350 (
    .din     (_zz_2591[31:0]        ), //i
    .dout    (fixTo_350_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_351 (
    .din     (_zz_2592[31:0]        ), //i
    .dout    (fixTo_351_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_352 (
    .din     (_zz_2593[31:0]        ), //i
    .dout    (fixTo_352_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_353 (
    .din     (_zz_2594[31:0]        ), //i
    .dout    (fixTo_353_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_354 (
    .din     (_zz_2595[31:0]        ), //i
    .dout    (fixTo_354_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_355 (
    .din     (_zz_2596[31:0]        ), //i
    .dout    (fixTo_355_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_356 (
    .din     (_zz_2597[31:0]        ), //i
    .dout    (fixTo_356_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_357 (
    .din     (_zz_2598[31:0]        ), //i
    .dout    (fixTo_357_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_358 (
    .din     (_zz_2599[31:0]        ), //i
    .dout    (fixTo_358_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_359 (
    .din     (_zz_2600[31:0]        ), //i
    .dout    (fixTo_359_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_360 (
    .din     (_zz_2601[31:0]        ), //i
    .dout    (fixTo_360_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_361 (
    .din     (_zz_2602[31:0]        ), //i
    .dout    (fixTo_361_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_362 (
    .din     (_zz_2603[31:0]        ), //i
    .dout    (fixTo_362_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_363 (
    .din     (_zz_2604[31:0]        ), //i
    .dout    (fixTo_363_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_364 (
    .din     (_zz_2605[31:0]        ), //i
    .dout    (fixTo_364_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_365 (
    .din     (_zz_2606[31:0]        ), //i
    .dout    (fixTo_365_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_366 (
    .din     (_zz_2607[31:0]        ), //i
    .dout    (fixTo_366_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_367 (
    .din     (_zz_2608[31:0]        ), //i
    .dout    (fixTo_367_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_368 (
    .din     (_zz_2609[31:0]        ), //i
    .dout    (fixTo_368_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_369 (
    .din     (_zz_2610[31:0]        ), //i
    .dout    (fixTo_369_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_370 (
    .din     (_zz_2611[31:0]        ), //i
    .dout    (fixTo_370_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_371 (
    .din     (_zz_2612[31:0]        ), //i
    .dout    (fixTo_371_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_372 (
    .din     (_zz_2613[31:0]        ), //i
    .dout    (fixTo_372_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_373 (
    .din     (_zz_2614[31:0]        ), //i
    .dout    (fixTo_373_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_374 (
    .din     (_zz_2615[31:0]        ), //i
    .dout    (fixTo_374_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_375 (
    .din     (_zz_2616[31:0]        ), //i
    .dout    (fixTo_375_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_376 (
    .din     (_zz_2617[31:0]        ), //i
    .dout    (fixTo_376_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_377 (
    .din     (_zz_2618[31:0]        ), //i
    .dout    (fixTo_377_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_378 (
    .din     (_zz_2619[31:0]        ), //i
    .dout    (fixTo_378_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_379 (
    .din     (_zz_2620[31:0]        ), //i
    .dout    (fixTo_379_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_380 (
    .din     (_zz_2621[31:0]        ), //i
    .dout    (fixTo_380_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_381 (
    .din     (_zz_2622[31:0]        ), //i
    .dout    (fixTo_381_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_382 (
    .din     (_zz_2623[31:0]        ), //i
    .dout    (fixTo_382_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_383 (
    .din     (_zz_2624[31:0]        ), //i
    .dout    (fixTo_383_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_384 (
    .din     (_zz_2625[31:0]        ), //i
    .dout    (fixTo_384_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_385 (
    .din     (_zz_2626[31:0]        ), //i
    .dout    (fixTo_385_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_386 (
    .din     (_zz_2627[31:0]        ), //i
    .dout    (fixTo_386_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_387 (
    .din     (_zz_2628[31:0]        ), //i
    .dout    (fixTo_387_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_388 (
    .din     (_zz_2629[31:0]        ), //i
    .dout    (fixTo_388_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_389 (
    .din     (_zz_2630[31:0]        ), //i
    .dout    (fixTo_389_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_390 (
    .din     (_zz_2631[31:0]        ), //i
    .dout    (fixTo_390_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_391 (
    .din     (_zz_2632[31:0]        ), //i
    .dout    (fixTo_391_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_392 (
    .din     (_zz_2633[31:0]        ), //i
    .dout    (fixTo_392_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_393 (
    .din     (_zz_2634[31:0]        ), //i
    .dout    (fixTo_393_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_394 (
    .din     (_zz_2635[31:0]        ), //i
    .dout    (fixTo_394_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_395 (
    .din     (_zz_2636[31:0]        ), //i
    .dout    (fixTo_395_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_396 (
    .din     (_zz_2637[31:0]        ), //i
    .dout    (fixTo_396_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_397 (
    .din     (_zz_2638[31:0]        ), //i
    .dout    (fixTo_397_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_398 (
    .din     (_zz_2639[31:0]        ), //i
    .dout    (fixTo_398_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_399 (
    .din     (_zz_2640[31:0]        ), //i
    .dout    (fixTo_399_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_400 (
    .din     (_zz_2641[31:0]        ), //i
    .dout    (fixTo_400_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_401 (
    .din     (_zz_2642[31:0]        ), //i
    .dout    (fixTo_401_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_402 (
    .din     (_zz_2643[31:0]        ), //i
    .dout    (fixTo_402_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_403 (
    .din     (_zz_2644[31:0]        ), //i
    .dout    (fixTo_403_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_404 (
    .din     (_zz_2645[31:0]        ), //i
    .dout    (fixTo_404_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_405 (
    .din     (_zz_2646[31:0]        ), //i
    .dout    (fixTo_405_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_406 (
    .din     (_zz_2647[31:0]        ), //i
    .dout    (fixTo_406_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_407 (
    .din     (_zz_2648[31:0]        ), //i
    .dout    (fixTo_407_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_408 (
    .din     (_zz_2649[31:0]        ), //i
    .dout    (fixTo_408_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_409 (
    .din     (_zz_2650[31:0]        ), //i
    .dout    (fixTo_409_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_410 (
    .din     (_zz_2651[31:0]        ), //i
    .dout    (fixTo_410_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_411 (
    .din     (_zz_2652[31:0]        ), //i
    .dout    (fixTo_411_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_412 (
    .din     (_zz_2653[31:0]        ), //i
    .dout    (fixTo_412_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_413 (
    .din     (_zz_2654[31:0]        ), //i
    .dout    (fixTo_413_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_414 (
    .din     (_zz_2655[31:0]        ), //i
    .dout    (fixTo_414_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_415 (
    .din     (_zz_2656[31:0]        ), //i
    .dout    (fixTo_415_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_416 (
    .din     (_zz_2657[31:0]        ), //i
    .dout    (fixTo_416_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_417 (
    .din     (_zz_2658[31:0]        ), //i
    .dout    (fixTo_417_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_418 (
    .din     (_zz_2659[31:0]        ), //i
    .dout    (fixTo_418_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_419 (
    .din     (_zz_2660[31:0]        ), //i
    .dout    (fixTo_419_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_420 (
    .din     (_zz_2661[31:0]        ), //i
    .dout    (fixTo_420_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_421 (
    .din     (_zz_2662[31:0]        ), //i
    .dout    (fixTo_421_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_422 (
    .din     (_zz_2663[31:0]        ), //i
    .dout    (fixTo_422_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_423 (
    .din     (_zz_2664[31:0]        ), //i
    .dout    (fixTo_423_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_424 (
    .din     (_zz_2665[31:0]        ), //i
    .dout    (fixTo_424_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_425 (
    .din     (_zz_2666[31:0]        ), //i
    .dout    (fixTo_425_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_426 (
    .din     (_zz_2667[31:0]        ), //i
    .dout    (fixTo_426_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_427 (
    .din     (_zz_2668[31:0]        ), //i
    .dout    (fixTo_427_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_428 (
    .din     (_zz_2669[31:0]        ), //i
    .dout    (fixTo_428_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_429 (
    .din     (_zz_2670[31:0]        ), //i
    .dout    (fixTo_429_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_430 (
    .din     (_zz_2671[31:0]        ), //i
    .dout    (fixTo_430_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_431 (
    .din     (_zz_2672[31:0]        ), //i
    .dout    (fixTo_431_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_432 (
    .din     (_zz_2673[31:0]        ), //i
    .dout    (fixTo_432_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_433 (
    .din     (_zz_2674[31:0]        ), //i
    .dout    (fixTo_433_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_434 (
    .din     (_zz_2675[31:0]        ), //i
    .dout    (fixTo_434_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_435 (
    .din     (_zz_2676[31:0]        ), //i
    .dout    (fixTo_435_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_436 (
    .din     (_zz_2677[31:0]        ), //i
    .dout    (fixTo_436_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_437 (
    .din     (_zz_2678[31:0]        ), //i
    .dout    (fixTo_437_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_438 (
    .din     (_zz_2679[31:0]        ), //i
    .dout    (fixTo_438_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_439 (
    .din     (_zz_2680[31:0]        ), //i
    .dout    (fixTo_439_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_440 (
    .din     (_zz_2681[31:0]        ), //i
    .dout    (fixTo_440_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_441 (
    .din     (_zz_2682[31:0]        ), //i
    .dout    (fixTo_441_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_442 (
    .din     (_zz_2683[31:0]        ), //i
    .dout    (fixTo_442_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_443 (
    .din     (_zz_2684[31:0]        ), //i
    .dout    (fixTo_443_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_444 (
    .din     (_zz_2685[31:0]        ), //i
    .dout    (fixTo_444_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_445 (
    .din     (_zz_2686[31:0]        ), //i
    .dout    (fixTo_445_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_446 (
    .din     (_zz_2687[31:0]        ), //i
    .dout    (fixTo_446_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_447 (
    .din     (_zz_2688[31:0]        ), //i
    .dout    (fixTo_447_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_448 (
    .din     (_zz_2689[31:0]        ), //i
    .dout    (fixTo_448_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_449 (
    .din     (_zz_2690[31:0]        ), //i
    .dout    (fixTo_449_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_450 (
    .din     (_zz_2691[31:0]        ), //i
    .dout    (fixTo_450_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_451 (
    .din     (_zz_2692[31:0]        ), //i
    .dout    (fixTo_451_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_452 (
    .din     (_zz_2693[31:0]        ), //i
    .dout    (fixTo_452_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_453 (
    .din     (_zz_2694[31:0]        ), //i
    .dout    (fixTo_453_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_454 (
    .din     (_zz_2695[31:0]        ), //i
    .dout    (fixTo_454_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_455 (
    .din     (_zz_2696[31:0]        ), //i
    .dout    (fixTo_455_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_456 (
    .din     (_zz_2697[31:0]        ), //i
    .dout    (fixTo_456_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_457 (
    .din     (_zz_2698[31:0]        ), //i
    .dout    (fixTo_457_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_458 (
    .din     (_zz_2699[31:0]        ), //i
    .dout    (fixTo_458_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_459 (
    .din     (_zz_2700[31:0]        ), //i
    .dout    (fixTo_459_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_460 (
    .din     (_zz_2701[31:0]        ), //i
    .dout    (fixTo_460_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_461 (
    .din     (_zz_2702[31:0]        ), //i
    .dout    (fixTo_461_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_462 (
    .din     (_zz_2703[31:0]        ), //i
    .dout    (fixTo_462_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_463 (
    .din     (_zz_2704[31:0]        ), //i
    .dout    (fixTo_463_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_464 (
    .din     (_zz_2705[31:0]        ), //i
    .dout    (fixTo_464_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_465 (
    .din     (_zz_2706[31:0]        ), //i
    .dout    (fixTo_465_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_466 (
    .din     (_zz_2707[31:0]        ), //i
    .dout    (fixTo_466_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_467 (
    .din     (_zz_2708[31:0]        ), //i
    .dout    (fixTo_467_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_468 (
    .din     (_zz_2709[31:0]        ), //i
    .dout    (fixTo_468_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_469 (
    .din     (_zz_2710[31:0]        ), //i
    .dout    (fixTo_469_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_470 (
    .din     (_zz_2711[31:0]        ), //i
    .dout    (fixTo_470_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_471 (
    .din     (_zz_2712[31:0]        ), //i
    .dout    (fixTo_471_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_472 (
    .din     (_zz_2713[31:0]        ), //i
    .dout    (fixTo_472_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_473 (
    .din     (_zz_2714[31:0]        ), //i
    .dout    (fixTo_473_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_474 (
    .din     (_zz_2715[31:0]        ), //i
    .dout    (fixTo_474_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_475 (
    .din     (_zz_2716[31:0]        ), //i
    .dout    (fixTo_475_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_476 (
    .din     (_zz_2717[31:0]        ), //i
    .dout    (fixTo_476_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_477 (
    .din     (_zz_2718[31:0]        ), //i
    .dout    (fixTo_477_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_478 (
    .din     (_zz_2719[31:0]        ), //i
    .dout    (fixTo_478_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_479 (
    .din     (_zz_2720[31:0]        ), //i
    .dout    (fixTo_479_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_480 (
    .din     (_zz_2721[31:0]        ), //i
    .dout    (fixTo_480_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_481 (
    .din     (_zz_2722[31:0]        ), //i
    .dout    (fixTo_481_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_482 (
    .din     (_zz_2723[31:0]        ), //i
    .dout    (fixTo_482_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_483 (
    .din     (_zz_2724[31:0]        ), //i
    .dout    (fixTo_483_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_484 (
    .din     (_zz_2725[31:0]        ), //i
    .dout    (fixTo_484_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_485 (
    .din     (_zz_2726[31:0]        ), //i
    .dout    (fixTo_485_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_486 (
    .din     (_zz_2727[31:0]        ), //i
    .dout    (fixTo_486_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_487 (
    .din     (_zz_2728[31:0]        ), //i
    .dout    (fixTo_487_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_488 (
    .din     (_zz_2729[31:0]        ), //i
    .dout    (fixTo_488_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_489 (
    .din     (_zz_2730[31:0]        ), //i
    .dout    (fixTo_489_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_490 (
    .din     (_zz_2731[31:0]        ), //i
    .dout    (fixTo_490_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_491 (
    .din     (_zz_2732[31:0]        ), //i
    .dout    (fixTo_491_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_492 (
    .din     (_zz_2733[31:0]        ), //i
    .dout    (fixTo_492_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_493 (
    .din     (_zz_2734[31:0]        ), //i
    .dout    (fixTo_493_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_494 (
    .din     (_zz_2735[31:0]        ), //i
    .dout    (fixTo_494_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_495 (
    .din     (_zz_2736[31:0]        ), //i
    .dout    (fixTo_495_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_496 (
    .din     (_zz_2737[31:0]        ), //i
    .dout    (fixTo_496_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_497 (
    .din     (_zz_2738[31:0]        ), //i
    .dout    (fixTo_497_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_498 (
    .din     (_zz_2739[31:0]        ), //i
    .dout    (fixTo_498_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_499 (
    .din     (_zz_2740[31:0]        ), //i
    .dout    (fixTo_499_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_500 (
    .din     (_zz_2741[31:0]        ), //i
    .dout    (fixTo_500_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_501 (
    .din     (_zz_2742[31:0]        ), //i
    .dout    (fixTo_501_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_502 (
    .din     (_zz_2743[31:0]        ), //i
    .dout    (fixTo_502_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_503 (
    .din     (_zz_2744[31:0]        ), //i
    .dout    (fixTo_503_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_504 (
    .din     (_zz_2745[31:0]        ), //i
    .dout    (fixTo_504_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_505 (
    .din     (_zz_2746[31:0]        ), //i
    .dout    (fixTo_505_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_506 (
    .din     (_zz_2747[31:0]        ), //i
    .dout    (fixTo_506_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_507 (
    .din     (_zz_2748[31:0]        ), //i
    .dout    (fixTo_507_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_508 (
    .din     (_zz_2749[31:0]        ), //i
    .dout    (fixTo_508_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_509 (
    .din     (_zz_2750[31:0]        ), //i
    .dout    (fixTo_509_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_510 (
    .din     (_zz_2751[31:0]        ), //i
    .dout    (fixTo_510_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_511 (
    .din     (_zz_2752[31:0]        ), //i
    .dout    (fixTo_511_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_512 (
    .din     (_zz_2753[31:0]        ), //i
    .dout    (fixTo_512_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_513 (
    .din     (_zz_2754[31:0]        ), //i
    .dout    (fixTo_513_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_514 (
    .din     (_zz_2755[31:0]        ), //i
    .dout    (fixTo_514_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_515 (
    .din     (_zz_2756[31:0]        ), //i
    .dout    (fixTo_515_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_516 (
    .din     (_zz_2757[31:0]        ), //i
    .dout    (fixTo_516_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_517 (
    .din     (_zz_2758[31:0]        ), //i
    .dout    (fixTo_517_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_518 (
    .din     (_zz_2759[31:0]        ), //i
    .dout    (fixTo_518_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_519 (
    .din     (_zz_2760[31:0]        ), //i
    .dout    (fixTo_519_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_520 (
    .din     (_zz_2761[31:0]        ), //i
    .dout    (fixTo_520_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_521 (
    .din     (_zz_2762[31:0]        ), //i
    .dout    (fixTo_521_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_522 (
    .din     (_zz_2763[31:0]        ), //i
    .dout    (fixTo_522_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_523 (
    .din     (_zz_2764[31:0]        ), //i
    .dout    (fixTo_523_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_524 (
    .din     (_zz_2765[31:0]        ), //i
    .dout    (fixTo_524_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_525 (
    .din     (_zz_2766[31:0]        ), //i
    .dout    (fixTo_525_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_526 (
    .din     (_zz_2767[31:0]        ), //i
    .dout    (fixTo_526_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_527 (
    .din     (_zz_2768[31:0]        ), //i
    .dout    (fixTo_527_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_528 (
    .din     (_zz_2769[31:0]        ), //i
    .dout    (fixTo_528_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_529 (
    .din     (_zz_2770[31:0]        ), //i
    .dout    (fixTo_529_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_530 (
    .din     (_zz_2771[31:0]        ), //i
    .dout    (fixTo_530_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_531 (
    .din     (_zz_2772[31:0]        ), //i
    .dout    (fixTo_531_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_532 (
    .din     (_zz_2773[31:0]        ), //i
    .dout    (fixTo_532_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_533 (
    .din     (_zz_2774[31:0]        ), //i
    .dout    (fixTo_533_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_534 (
    .din     (_zz_2775[31:0]        ), //i
    .dout    (fixTo_534_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_535 (
    .din     (_zz_2776[31:0]        ), //i
    .dout    (fixTo_535_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_536 (
    .din     (_zz_2777[31:0]        ), //i
    .dout    (fixTo_536_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_537 (
    .din     (_zz_2778[31:0]        ), //i
    .dout    (fixTo_537_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_538 (
    .din     (_zz_2779[31:0]        ), //i
    .dout    (fixTo_538_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_539 (
    .din     (_zz_2780[31:0]        ), //i
    .dout    (fixTo_539_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_540 (
    .din     (_zz_2781[31:0]        ), //i
    .dout    (fixTo_540_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_541 (
    .din     (_zz_2782[31:0]        ), //i
    .dout    (fixTo_541_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_542 (
    .din     (_zz_2783[31:0]        ), //i
    .dout    (fixTo_542_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_543 (
    .din     (_zz_2784[31:0]        ), //i
    .dout    (fixTo_543_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_544 (
    .din     (_zz_2785[31:0]        ), //i
    .dout    (fixTo_544_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_545 (
    .din     (_zz_2786[31:0]        ), //i
    .dout    (fixTo_545_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_546 (
    .din     (_zz_2787[31:0]        ), //i
    .dout    (fixTo_546_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_547 (
    .din     (_zz_2788[31:0]        ), //i
    .dout    (fixTo_547_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_548 (
    .din     (_zz_2789[31:0]        ), //i
    .dout    (fixTo_548_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_549 (
    .din     (_zz_2790[31:0]        ), //i
    .dout    (fixTo_549_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_550 (
    .din     (_zz_2791[31:0]        ), //i
    .dout    (fixTo_550_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_551 (
    .din     (_zz_2792[31:0]        ), //i
    .dout    (fixTo_551_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_552 (
    .din     (_zz_2793[31:0]        ), //i
    .dout    (fixTo_552_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_553 (
    .din     (_zz_2794[31:0]        ), //i
    .dout    (fixTo_553_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_554 (
    .din     (_zz_2795[31:0]        ), //i
    .dout    (fixTo_554_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_555 (
    .din     (_zz_2796[31:0]        ), //i
    .dout    (fixTo_555_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_556 (
    .din     (_zz_2797[31:0]        ), //i
    .dout    (fixTo_556_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_557 (
    .din     (_zz_2798[31:0]        ), //i
    .dout    (fixTo_557_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_558 (
    .din     (_zz_2799[31:0]        ), //i
    .dout    (fixTo_558_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_559 (
    .din     (_zz_2800[31:0]        ), //i
    .dout    (fixTo_559_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_560 (
    .din     (_zz_2801[31:0]        ), //i
    .dout    (fixTo_560_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_561 (
    .din     (_zz_2802[31:0]        ), //i
    .dout    (fixTo_561_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_562 (
    .din     (_zz_2803[31:0]        ), //i
    .dout    (fixTo_562_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_563 (
    .din     (_zz_2804[31:0]        ), //i
    .dout    (fixTo_563_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_564 (
    .din     (_zz_2805[31:0]        ), //i
    .dout    (fixTo_564_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_565 (
    .din     (_zz_2806[31:0]        ), //i
    .dout    (fixTo_565_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_566 (
    .din     (_zz_2807[31:0]        ), //i
    .dout    (fixTo_566_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_567 (
    .din     (_zz_2808[31:0]        ), //i
    .dout    (fixTo_567_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_568 (
    .din     (_zz_2809[31:0]        ), //i
    .dout    (fixTo_568_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_569 (
    .din     (_zz_2810[31:0]        ), //i
    .dout    (fixTo_569_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_570 (
    .din     (_zz_2811[31:0]        ), //i
    .dout    (fixTo_570_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_571 (
    .din     (_zz_2812[31:0]        ), //i
    .dout    (fixTo_571_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_572 (
    .din     (_zz_2813[31:0]        ), //i
    .dout    (fixTo_572_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_573 (
    .din     (_zz_2814[31:0]        ), //i
    .dout    (fixTo_573_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_574 (
    .din     (_zz_2815[31:0]        ), //i
    .dout    (fixTo_574_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_575 (
    .din     (_zz_2816[31:0]        ), //i
    .dout    (fixTo_575_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_576 (
    .din     (_zz_2817[31:0]        ), //i
    .dout    (fixTo_576_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_577 (
    .din     (_zz_2818[31:0]        ), //i
    .dout    (fixTo_577_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_578 (
    .din     (_zz_2819[31:0]        ), //i
    .dout    (fixTo_578_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_579 (
    .din     (_zz_2820[31:0]        ), //i
    .dout    (fixTo_579_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_580 (
    .din     (_zz_2821[31:0]        ), //i
    .dout    (fixTo_580_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_581 (
    .din     (_zz_2822[31:0]        ), //i
    .dout    (fixTo_581_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_582 (
    .din     (_zz_2823[31:0]        ), //i
    .dout    (fixTo_582_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_583 (
    .din     (_zz_2824[31:0]        ), //i
    .dout    (fixTo_583_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_584 (
    .din     (_zz_2825[31:0]        ), //i
    .dout    (fixTo_584_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_585 (
    .din     (_zz_2826[31:0]        ), //i
    .dout    (fixTo_585_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_586 (
    .din     (_zz_2827[31:0]        ), //i
    .dout    (fixTo_586_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_587 (
    .din     (_zz_2828[31:0]        ), //i
    .dout    (fixTo_587_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_588 (
    .din     (_zz_2829[31:0]        ), //i
    .dout    (fixTo_588_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_589 (
    .din     (_zz_2830[31:0]        ), //i
    .dout    (fixTo_589_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_590 (
    .din     (_zz_2831[31:0]        ), //i
    .dout    (fixTo_590_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_591 (
    .din     (_zz_2832[31:0]        ), //i
    .dout    (fixTo_591_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_592 (
    .din     (_zz_2833[31:0]        ), //i
    .dout    (fixTo_592_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_593 (
    .din     (_zz_2834[31:0]        ), //i
    .dout    (fixTo_593_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_594 (
    .din     (_zz_2835[31:0]        ), //i
    .dout    (fixTo_594_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_595 (
    .din     (_zz_2836[31:0]        ), //i
    .dout    (fixTo_595_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_596 (
    .din     (_zz_2837[31:0]        ), //i
    .dout    (fixTo_596_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_597 (
    .din     (_zz_2838[31:0]        ), //i
    .dout    (fixTo_597_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_598 (
    .din     (_zz_2839[31:0]        ), //i
    .dout    (fixTo_598_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_599 (
    .din     (_zz_2840[31:0]        ), //i
    .dout    (fixTo_599_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_600 (
    .din     (_zz_2841[31:0]        ), //i
    .dout    (fixTo_600_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_601 (
    .din     (_zz_2842[31:0]        ), //i
    .dout    (fixTo_601_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_602 (
    .din     (_zz_2843[31:0]        ), //i
    .dout    (fixTo_602_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_603 (
    .din     (_zz_2844[31:0]        ), //i
    .dout    (fixTo_603_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_604 (
    .din     (_zz_2845[31:0]        ), //i
    .dout    (fixTo_604_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_605 (
    .din     (_zz_2846[31:0]        ), //i
    .dout    (fixTo_605_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_606 (
    .din     (_zz_2847[31:0]        ), //i
    .dout    (fixTo_606_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_607 (
    .din     (_zz_2848[31:0]        ), //i
    .dout    (fixTo_607_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_608 (
    .din     (_zz_2849[31:0]        ), //i
    .dout    (fixTo_608_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_609 (
    .din     (_zz_2850[31:0]        ), //i
    .dout    (fixTo_609_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_610 (
    .din     (_zz_2851[31:0]        ), //i
    .dout    (fixTo_610_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_611 (
    .din     (_zz_2852[31:0]        ), //i
    .dout    (fixTo_611_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_612 (
    .din     (_zz_2853[31:0]        ), //i
    .dout    (fixTo_612_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_613 (
    .din     (_zz_2854[31:0]        ), //i
    .dout    (fixTo_613_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_614 (
    .din     (_zz_2855[31:0]        ), //i
    .dout    (fixTo_614_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_615 (
    .din     (_zz_2856[31:0]        ), //i
    .dout    (fixTo_615_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_616 (
    .din     (_zz_2857[31:0]        ), //i
    .dout    (fixTo_616_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_617 (
    .din     (_zz_2858[31:0]        ), //i
    .dout    (fixTo_617_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_618 (
    .din     (_zz_2859[31:0]        ), //i
    .dout    (fixTo_618_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_619 (
    .din     (_zz_2860[31:0]        ), //i
    .dout    (fixTo_619_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_620 (
    .din     (_zz_2861[31:0]        ), //i
    .dout    (fixTo_620_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_621 (
    .din     (_zz_2862[31:0]        ), //i
    .dout    (fixTo_621_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_622 (
    .din     (_zz_2863[31:0]        ), //i
    .dout    (fixTo_622_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_623 (
    .din     (_zz_2864[31:0]        ), //i
    .dout    (fixTo_623_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_624 (
    .din     (_zz_2865[31:0]        ), //i
    .dout    (fixTo_624_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_625 (
    .din     (_zz_2866[31:0]        ), //i
    .dout    (fixTo_625_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_626 (
    .din     (_zz_2867[31:0]        ), //i
    .dout    (fixTo_626_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_627 (
    .din     (_zz_2868[31:0]        ), //i
    .dout    (fixTo_627_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_628 (
    .din     (_zz_2869[31:0]        ), //i
    .dout    (fixTo_628_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_629 (
    .din     (_zz_2870[31:0]        ), //i
    .dout    (fixTo_629_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_630 (
    .din     (_zz_2871[31:0]        ), //i
    .dout    (fixTo_630_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_631 (
    .din     (_zz_2872[31:0]        ), //i
    .dout    (fixTo_631_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_632 (
    .din     (_zz_2873[31:0]        ), //i
    .dout    (fixTo_632_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_633 (
    .din     (_zz_2874[31:0]        ), //i
    .dout    (fixTo_633_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_634 (
    .din     (_zz_2875[31:0]        ), //i
    .dout    (fixTo_634_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_635 (
    .din     (_zz_2876[31:0]        ), //i
    .dout    (fixTo_635_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_636 (
    .din     (_zz_2877[31:0]        ), //i
    .dout    (fixTo_636_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_637 (
    .din     (_zz_2878[31:0]        ), //i
    .dout    (fixTo_637_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_638 (
    .din     (_zz_2879[31:0]        ), //i
    .dout    (fixTo_638_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_639 (
    .din     (_zz_2880[31:0]        ), //i
    .dout    (fixTo_639_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_640 (
    .din     (_zz_2881[31:0]        ), //i
    .dout    (fixTo_640_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_641 (
    .din     (_zz_2882[31:0]        ), //i
    .dout    (fixTo_641_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_642 (
    .din     (_zz_2883[31:0]        ), //i
    .dout    (fixTo_642_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_643 (
    .din     (_zz_2884[31:0]        ), //i
    .dout    (fixTo_643_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_644 (
    .din     (_zz_2885[31:0]        ), //i
    .dout    (fixTo_644_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_645 (
    .din     (_zz_2886[31:0]        ), //i
    .dout    (fixTo_645_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_646 (
    .din     (_zz_2887[31:0]        ), //i
    .dout    (fixTo_646_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_647 (
    .din     (_zz_2888[31:0]        ), //i
    .dout    (fixTo_647_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_648 (
    .din     (_zz_2889[31:0]        ), //i
    .dout    (fixTo_648_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_649 (
    .din     (_zz_2890[31:0]        ), //i
    .dout    (fixTo_649_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_650 (
    .din     (_zz_2891[31:0]        ), //i
    .dout    (fixTo_650_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_651 (
    .din     (_zz_2892[31:0]        ), //i
    .dout    (fixTo_651_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_652 (
    .din     (_zz_2893[31:0]        ), //i
    .dout    (fixTo_652_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_653 (
    .din     (_zz_2894[31:0]        ), //i
    .dout    (fixTo_653_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_654 (
    .din     (_zz_2895[31:0]        ), //i
    .dout    (fixTo_654_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_655 (
    .din     (_zz_2896[31:0]        ), //i
    .dout    (fixTo_655_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_656 (
    .din     (_zz_2897[31:0]        ), //i
    .dout    (fixTo_656_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_657 (
    .din     (_zz_2898[31:0]        ), //i
    .dout    (fixTo_657_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_658 (
    .din     (_zz_2899[31:0]        ), //i
    .dout    (fixTo_658_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_659 (
    .din     (_zz_2900[31:0]        ), //i
    .dout    (fixTo_659_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_660 (
    .din     (_zz_2901[31:0]        ), //i
    .dout    (fixTo_660_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_661 (
    .din     (_zz_2902[31:0]        ), //i
    .dout    (fixTo_661_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_662 (
    .din     (_zz_2903[31:0]        ), //i
    .dout    (fixTo_662_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_663 (
    .din     (_zz_2904[31:0]        ), //i
    .dout    (fixTo_663_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_664 (
    .din     (_zz_2905[31:0]        ), //i
    .dout    (fixTo_664_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_665 (
    .din     (_zz_2906[31:0]        ), //i
    .dout    (fixTo_665_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_666 (
    .din     (_zz_2907[31:0]        ), //i
    .dout    (fixTo_666_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_667 (
    .din     (_zz_2908[31:0]        ), //i
    .dout    (fixTo_667_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_668 (
    .din     (_zz_2909[31:0]        ), //i
    .dout    (fixTo_668_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_669 (
    .din     (_zz_2910[31:0]        ), //i
    .dout    (fixTo_669_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_670 (
    .din     (_zz_2911[31:0]        ), //i
    .dout    (fixTo_670_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_671 (
    .din     (_zz_2912[31:0]        ), //i
    .dout    (fixTo_671_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_672 (
    .din     (_zz_2913[31:0]        ), //i
    .dout    (fixTo_672_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_673 (
    .din     (_zz_2914[31:0]        ), //i
    .dout    (fixTo_673_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_674 (
    .din     (_zz_2915[31:0]        ), //i
    .dout    (fixTo_674_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_675 (
    .din     (_zz_2916[31:0]        ), //i
    .dout    (fixTo_675_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_676 (
    .din     (_zz_2917[31:0]        ), //i
    .dout    (fixTo_676_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_677 (
    .din     (_zz_2918[31:0]        ), //i
    .dout    (fixTo_677_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_678 (
    .din     (_zz_2919[31:0]        ), //i
    .dout    (fixTo_678_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_679 (
    .din     (_zz_2920[31:0]        ), //i
    .dout    (fixTo_679_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_680 (
    .din     (_zz_2921[31:0]        ), //i
    .dout    (fixTo_680_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_681 (
    .din     (_zz_2922[31:0]        ), //i
    .dout    (fixTo_681_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_682 (
    .din     (_zz_2923[31:0]        ), //i
    .dout    (fixTo_682_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_683 (
    .din     (_zz_2924[31:0]        ), //i
    .dout    (fixTo_683_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_684 (
    .din     (_zz_2925[31:0]        ), //i
    .dout    (fixTo_684_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_685 (
    .din     (_zz_2926[31:0]        ), //i
    .dout    (fixTo_685_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_686 (
    .din     (_zz_2927[31:0]        ), //i
    .dout    (fixTo_686_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_687 (
    .din     (_zz_2928[31:0]        ), //i
    .dout    (fixTo_687_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_688 (
    .din     (_zz_2929[31:0]        ), //i
    .dout    (fixTo_688_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_689 (
    .din     (_zz_2930[31:0]        ), //i
    .dout    (fixTo_689_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_690 (
    .din     (_zz_2931[31:0]        ), //i
    .dout    (fixTo_690_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_691 (
    .din     (_zz_2932[31:0]        ), //i
    .dout    (fixTo_691_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_692 (
    .din     (_zz_2933[31:0]        ), //i
    .dout    (fixTo_692_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_693 (
    .din     (_zz_2934[31:0]        ), //i
    .dout    (fixTo_693_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_694 (
    .din     (_zz_2935[31:0]        ), //i
    .dout    (fixTo_694_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_695 (
    .din     (_zz_2936[31:0]        ), //i
    .dout    (fixTo_695_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_696 (
    .din     (_zz_2937[31:0]        ), //i
    .dout    (fixTo_696_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_697 (
    .din     (_zz_2938[31:0]        ), //i
    .dout    (fixTo_697_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_698 (
    .din     (_zz_2939[31:0]        ), //i
    .dout    (fixTo_698_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_699 (
    .din     (_zz_2940[31:0]        ), //i
    .dout    (fixTo_699_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_700 (
    .din     (_zz_2941[31:0]        ), //i
    .dout    (fixTo_700_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_701 (
    .din     (_zz_2942[31:0]        ), //i
    .dout    (fixTo_701_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_702 (
    .din     (_zz_2943[31:0]        ), //i
    .dout    (fixTo_702_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_703 (
    .din     (_zz_2944[31:0]        ), //i
    .dout    (fixTo_703_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_704 (
    .din     (_zz_2945[31:0]        ), //i
    .dout    (fixTo_704_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_705 (
    .din     (_zz_2946[31:0]        ), //i
    .dout    (fixTo_705_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_706 (
    .din     (_zz_2947[31:0]        ), //i
    .dout    (fixTo_706_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_707 (
    .din     (_zz_2948[31:0]        ), //i
    .dout    (fixTo_707_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_708 (
    .din     (_zz_2949[31:0]        ), //i
    .dout    (fixTo_708_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_709 (
    .din     (_zz_2950[31:0]        ), //i
    .dout    (fixTo_709_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_710 (
    .din     (_zz_2951[31:0]        ), //i
    .dout    (fixTo_710_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_711 (
    .din     (_zz_2952[31:0]        ), //i
    .dout    (fixTo_711_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_712 (
    .din     (_zz_2953[31:0]        ), //i
    .dout    (fixTo_712_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_713 (
    .din     (_zz_2954[31:0]        ), //i
    .dout    (fixTo_713_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_714 (
    .din     (_zz_2955[31:0]        ), //i
    .dout    (fixTo_714_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_715 (
    .din     (_zz_2956[31:0]        ), //i
    .dout    (fixTo_715_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_716 (
    .din     (_zz_2957[31:0]        ), //i
    .dout    (fixTo_716_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_717 (
    .din     (_zz_2958[31:0]        ), //i
    .dout    (fixTo_717_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_718 (
    .din     (_zz_2959[31:0]        ), //i
    .dout    (fixTo_718_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_719 (
    .din     (_zz_2960[31:0]        ), //i
    .dout    (fixTo_719_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_720 (
    .din     (_zz_2961[31:0]        ), //i
    .dout    (fixTo_720_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_721 (
    .din     (_zz_2962[31:0]        ), //i
    .dout    (fixTo_721_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_722 (
    .din     (_zz_2963[31:0]        ), //i
    .dout    (fixTo_722_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_723 (
    .din     (_zz_2964[31:0]        ), //i
    .dout    (fixTo_723_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_724 (
    .din     (_zz_2965[31:0]        ), //i
    .dout    (fixTo_724_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_725 (
    .din     (_zz_2966[31:0]        ), //i
    .dout    (fixTo_725_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_726 (
    .din     (_zz_2967[31:0]        ), //i
    .dout    (fixTo_726_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_727 (
    .din     (_zz_2968[31:0]        ), //i
    .dout    (fixTo_727_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_728 (
    .din     (_zz_2969[31:0]        ), //i
    .dout    (fixTo_728_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_729 (
    .din     (_zz_2970[31:0]        ), //i
    .dout    (fixTo_729_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_730 (
    .din     (_zz_2971[31:0]        ), //i
    .dout    (fixTo_730_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_731 (
    .din     (_zz_2972[31:0]        ), //i
    .dout    (fixTo_731_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_732 (
    .din     (_zz_2973[31:0]        ), //i
    .dout    (fixTo_732_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_733 (
    .din     (_zz_2974[31:0]        ), //i
    .dout    (fixTo_733_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_734 (
    .din     (_zz_2975[31:0]        ), //i
    .dout    (fixTo_734_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_735 (
    .din     (_zz_2976[31:0]        ), //i
    .dout    (fixTo_735_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_736 (
    .din     (_zz_2977[31:0]        ), //i
    .dout    (fixTo_736_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_737 (
    .din     (_zz_2978[31:0]        ), //i
    .dout    (fixTo_737_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_738 (
    .din     (_zz_2979[31:0]        ), //i
    .dout    (fixTo_738_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_739 (
    .din     (_zz_2980[31:0]        ), //i
    .dout    (fixTo_739_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_740 (
    .din     (_zz_2981[31:0]        ), //i
    .dout    (fixTo_740_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_741 (
    .din     (_zz_2982[31:0]        ), //i
    .dout    (fixTo_741_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_742 (
    .din     (_zz_2983[31:0]        ), //i
    .dout    (fixTo_742_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_743 (
    .din     (_zz_2984[31:0]        ), //i
    .dout    (fixTo_743_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_744 (
    .din     (_zz_2985[31:0]        ), //i
    .dout    (fixTo_744_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_745 (
    .din     (_zz_2986[31:0]        ), //i
    .dout    (fixTo_745_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_746 (
    .din     (_zz_2987[31:0]        ), //i
    .dout    (fixTo_746_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_747 (
    .din     (_zz_2988[31:0]        ), //i
    .dout    (fixTo_747_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_748 (
    .din     (_zz_2989[31:0]        ), //i
    .dout    (fixTo_748_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_749 (
    .din     (_zz_2990[31:0]        ), //i
    .dout    (fixTo_749_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_750 (
    .din     (_zz_2991[31:0]        ), //i
    .dout    (fixTo_750_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_751 (
    .din     (_zz_2992[31:0]        ), //i
    .dout    (fixTo_751_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_752 (
    .din     (_zz_2993[31:0]        ), //i
    .dout    (fixTo_752_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_753 (
    .din     (_zz_2994[31:0]        ), //i
    .dout    (fixTo_753_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_754 (
    .din     (_zz_2995[31:0]        ), //i
    .dout    (fixTo_754_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_755 (
    .din     (_zz_2996[31:0]        ), //i
    .dout    (fixTo_755_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_756 (
    .din     (_zz_2997[31:0]        ), //i
    .dout    (fixTo_756_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_757 (
    .din     (_zz_2998[31:0]        ), //i
    .dout    (fixTo_757_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_758 (
    .din     (_zz_2999[31:0]        ), //i
    .dout    (fixTo_758_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_759 (
    .din     (_zz_3000[31:0]        ), //i
    .dout    (fixTo_759_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_760 (
    .din     (_zz_3001[31:0]        ), //i
    .dout    (fixTo_760_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_761 (
    .din     (_zz_3002[31:0]        ), //i
    .dout    (fixTo_761_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_762 (
    .din     (_zz_3003[31:0]        ), //i
    .dout    (fixTo_762_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_763 (
    .din     (_zz_3004[31:0]        ), //i
    .dout    (fixTo_763_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_764 (
    .din     (_zz_3005[31:0]        ), //i
    .dout    (fixTo_764_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_765 (
    .din     (_zz_3006[31:0]        ), //i
    .dout    (fixTo_765_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_766 (
    .din     (_zz_3007[31:0]        ), //i
    .dout    (fixTo_766_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_767 (
    .din     (_zz_3008[31:0]        ), //i
    .dout    (fixTo_767_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_768 (
    .din     (_zz_3009[31:0]        ), //i
    .dout    (fixTo_768_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_769 (
    .din     (_zz_3010[31:0]        ), //i
    .dout    (fixTo_769_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_770 (
    .din     (_zz_3011[31:0]        ), //i
    .dout    (fixTo_770_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_771 (
    .din     (_zz_3012[31:0]        ), //i
    .dout    (fixTo_771_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_772 (
    .din     (_zz_3013[31:0]        ), //i
    .dout    (fixTo_772_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_773 (
    .din     (_zz_3014[31:0]        ), //i
    .dout    (fixTo_773_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_774 (
    .din     (_zz_3015[31:0]        ), //i
    .dout    (fixTo_774_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_775 (
    .din     (_zz_3016[31:0]        ), //i
    .dout    (fixTo_775_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_776 (
    .din     (_zz_3017[31:0]        ), //i
    .dout    (fixTo_776_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_777 (
    .din     (_zz_3018[31:0]        ), //i
    .dout    (fixTo_777_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_778 (
    .din     (_zz_3019[31:0]        ), //i
    .dout    (fixTo_778_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_779 (
    .din     (_zz_3020[31:0]        ), //i
    .dout    (fixTo_779_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_780 (
    .din     (_zz_3021[31:0]        ), //i
    .dout    (fixTo_780_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_781 (
    .din     (_zz_3022[31:0]        ), //i
    .dout    (fixTo_781_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_782 (
    .din     (_zz_3023[31:0]        ), //i
    .dout    (fixTo_782_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_783 (
    .din     (_zz_3024[31:0]        ), //i
    .dout    (fixTo_783_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_784 (
    .din     (_zz_3025[31:0]        ), //i
    .dout    (fixTo_784_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_785 (
    .din     (_zz_3026[31:0]        ), //i
    .dout    (fixTo_785_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_786 (
    .din     (_zz_3027[31:0]        ), //i
    .dout    (fixTo_786_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_787 (
    .din     (_zz_3028[31:0]        ), //i
    .dout    (fixTo_787_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_788 (
    .din     (_zz_3029[31:0]        ), //i
    .dout    (fixTo_788_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_789 (
    .din     (_zz_3030[31:0]        ), //i
    .dout    (fixTo_789_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_790 (
    .din     (_zz_3031[31:0]        ), //i
    .dout    (fixTo_790_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_791 (
    .din     (_zz_3032[31:0]        ), //i
    .dout    (fixTo_791_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_792 (
    .din     (_zz_3033[31:0]        ), //i
    .dout    (fixTo_792_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_793 (
    .din     (_zz_3034[31:0]        ), //i
    .dout    (fixTo_793_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_794 (
    .din     (_zz_3035[31:0]        ), //i
    .dout    (fixTo_794_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_795 (
    .din     (_zz_3036[31:0]        ), //i
    .dout    (fixTo_795_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_796 (
    .din     (_zz_3037[31:0]        ), //i
    .dout    (fixTo_796_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_797 (
    .din     (_zz_3038[31:0]        ), //i
    .dout    (fixTo_797_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_798 (
    .din     (_zz_3039[31:0]        ), //i
    .dout    (fixTo_798_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_799 (
    .din     (_zz_3040[31:0]        ), //i
    .dout    (fixTo_799_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_800 (
    .din     (_zz_3041[31:0]        ), //i
    .dout    (fixTo_800_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_801 (
    .din     (_zz_3042[31:0]        ), //i
    .dout    (fixTo_801_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_802 (
    .din     (_zz_3043[31:0]        ), //i
    .dout    (fixTo_802_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_803 (
    .din     (_zz_3044[31:0]        ), //i
    .dout    (fixTo_803_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_804 (
    .din     (_zz_3045[31:0]        ), //i
    .dout    (fixTo_804_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_805 (
    .din     (_zz_3046[31:0]        ), //i
    .dout    (fixTo_805_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_806 (
    .din     (_zz_3047[31:0]        ), //i
    .dout    (fixTo_806_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_807 (
    .din     (_zz_3048[31:0]        ), //i
    .dout    (fixTo_807_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_808 (
    .din     (_zz_3049[31:0]        ), //i
    .dout    (fixTo_808_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_809 (
    .din     (_zz_3050[31:0]        ), //i
    .dout    (fixTo_809_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_810 (
    .din     (_zz_3051[31:0]        ), //i
    .dout    (fixTo_810_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_811 (
    .din     (_zz_3052[31:0]        ), //i
    .dout    (fixTo_811_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_812 (
    .din     (_zz_3053[31:0]        ), //i
    .dout    (fixTo_812_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_813 (
    .din     (_zz_3054[31:0]        ), //i
    .dout    (fixTo_813_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_814 (
    .din     (_zz_3055[31:0]        ), //i
    .dout    (fixTo_814_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_815 (
    .din     (_zz_3056[31:0]        ), //i
    .dout    (fixTo_815_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_816 (
    .din     (_zz_3057[31:0]        ), //i
    .dout    (fixTo_816_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_817 (
    .din     (_zz_3058[31:0]        ), //i
    .dout    (fixTo_817_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_818 (
    .din     (_zz_3059[31:0]        ), //i
    .dout    (fixTo_818_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_819 (
    .din     (_zz_3060[31:0]        ), //i
    .dout    (fixTo_819_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_820 (
    .din     (_zz_3061[31:0]        ), //i
    .dout    (fixTo_820_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_821 (
    .din     (_zz_3062[31:0]        ), //i
    .dout    (fixTo_821_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_822 (
    .din     (_zz_3063[31:0]        ), //i
    .dout    (fixTo_822_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_823 (
    .din     (_zz_3064[31:0]        ), //i
    .dout    (fixTo_823_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_824 (
    .din     (_zz_3065[31:0]        ), //i
    .dout    (fixTo_824_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_825 (
    .din     (_zz_3066[31:0]        ), //i
    .dout    (fixTo_825_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_826 (
    .din     (_zz_3067[31:0]        ), //i
    .dout    (fixTo_826_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_827 (
    .din     (_zz_3068[31:0]        ), //i
    .dout    (fixTo_827_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_828 (
    .din     (_zz_3069[31:0]        ), //i
    .dout    (fixTo_828_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_829 (
    .din     (_zz_3070[31:0]        ), //i
    .dout    (fixTo_829_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_830 (
    .din     (_zz_3071[31:0]        ), //i
    .dout    (fixTo_830_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_831 (
    .din     (_zz_3072[31:0]        ), //i
    .dout    (fixTo_831_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_832 (
    .din     (_zz_3073[31:0]        ), //i
    .dout    (fixTo_832_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_833 (
    .din     (_zz_3074[31:0]        ), //i
    .dout    (fixTo_833_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_834 (
    .din     (_zz_3075[31:0]        ), //i
    .dout    (fixTo_834_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_835 (
    .din     (_zz_3076[31:0]        ), //i
    .dout    (fixTo_835_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_836 (
    .din     (_zz_3077[31:0]        ), //i
    .dout    (fixTo_836_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_837 (
    .din     (_zz_3078[31:0]        ), //i
    .dout    (fixTo_837_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_838 (
    .din     (_zz_3079[31:0]        ), //i
    .dout    (fixTo_838_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_839 (
    .din     (_zz_3080[31:0]        ), //i
    .dout    (fixTo_839_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_840 (
    .din     (_zz_3081[31:0]        ), //i
    .dout    (fixTo_840_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_841 (
    .din     (_zz_3082[31:0]        ), //i
    .dout    (fixTo_841_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_842 (
    .din     (_zz_3083[31:0]        ), //i
    .dout    (fixTo_842_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_843 (
    .din     (_zz_3084[31:0]        ), //i
    .dout    (fixTo_843_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_844 (
    .din     (_zz_3085[31:0]        ), //i
    .dout    (fixTo_844_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_845 (
    .din     (_zz_3086[31:0]        ), //i
    .dout    (fixTo_845_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_846 (
    .din     (_zz_3087[31:0]        ), //i
    .dout    (fixTo_846_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_847 (
    .din     (_zz_3088[31:0]        ), //i
    .dout    (fixTo_847_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_848 (
    .din     (_zz_3089[31:0]        ), //i
    .dout    (fixTo_848_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_849 (
    .din     (_zz_3090[31:0]        ), //i
    .dout    (fixTo_849_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_850 (
    .din     (_zz_3091[31:0]        ), //i
    .dout    (fixTo_850_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_851 (
    .din     (_zz_3092[31:0]        ), //i
    .dout    (fixTo_851_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_852 (
    .din     (_zz_3093[31:0]        ), //i
    .dout    (fixTo_852_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_853 (
    .din     (_zz_3094[31:0]        ), //i
    .dout    (fixTo_853_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_854 (
    .din     (_zz_3095[31:0]        ), //i
    .dout    (fixTo_854_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_855 (
    .din     (_zz_3096[31:0]        ), //i
    .dout    (fixTo_855_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_856 (
    .din     (_zz_3097[31:0]        ), //i
    .dout    (fixTo_856_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_857 (
    .din     (_zz_3098[31:0]        ), //i
    .dout    (fixTo_857_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_858 (
    .din     (_zz_3099[31:0]        ), //i
    .dout    (fixTo_858_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_859 (
    .din     (_zz_3100[31:0]        ), //i
    .dout    (fixTo_859_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_860 (
    .din     (_zz_3101[31:0]        ), //i
    .dout    (fixTo_860_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_861 (
    .din     (_zz_3102[31:0]        ), //i
    .dout    (fixTo_861_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_862 (
    .din     (_zz_3103[31:0]        ), //i
    .dout    (fixTo_862_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_863 (
    .din     (_zz_3104[31:0]        ), //i
    .dout    (fixTo_863_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_864 (
    .din     (_zz_3105[31:0]        ), //i
    .dout    (fixTo_864_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_865 (
    .din     (_zz_3106[31:0]        ), //i
    .dout    (fixTo_865_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_866 (
    .din     (_zz_3107[31:0]        ), //i
    .dout    (fixTo_866_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_867 (
    .din     (_zz_3108[31:0]        ), //i
    .dout    (fixTo_867_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_868 (
    .din     (_zz_3109[31:0]        ), //i
    .dout    (fixTo_868_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_869 (
    .din     (_zz_3110[31:0]        ), //i
    .dout    (fixTo_869_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_870 (
    .din     (_zz_3111[31:0]        ), //i
    .dout    (fixTo_870_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_871 (
    .din     (_zz_3112[31:0]        ), //i
    .dout    (fixTo_871_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_872 (
    .din     (_zz_3113[31:0]        ), //i
    .dout    (fixTo_872_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_873 (
    .din     (_zz_3114[31:0]        ), //i
    .dout    (fixTo_873_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_874 (
    .din     (_zz_3115[31:0]        ), //i
    .dout    (fixTo_874_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_875 (
    .din     (_zz_3116[31:0]        ), //i
    .dout    (fixTo_875_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_876 (
    .din     (_zz_3117[31:0]        ), //i
    .dout    (fixTo_876_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_877 (
    .din     (_zz_3118[31:0]        ), //i
    .dout    (fixTo_877_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_878 (
    .din     (_zz_3119[31:0]        ), //i
    .dout    (fixTo_878_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_879 (
    .din     (_zz_3120[31:0]        ), //i
    .dout    (fixTo_879_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_880 (
    .din     (_zz_3121[31:0]        ), //i
    .dout    (fixTo_880_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_881 (
    .din     (_zz_3122[31:0]        ), //i
    .dout    (fixTo_881_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_882 (
    .din     (_zz_3123[31:0]        ), //i
    .dout    (fixTo_882_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_883 (
    .din     (_zz_3124[31:0]        ), //i
    .dout    (fixTo_883_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_884 (
    .din     (_zz_3125[31:0]        ), //i
    .dout    (fixTo_884_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_885 (
    .din     (_zz_3126[31:0]        ), //i
    .dout    (fixTo_885_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_886 (
    .din     (_zz_3127[31:0]        ), //i
    .dout    (fixTo_886_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_887 (
    .din     (_zz_3128[31:0]        ), //i
    .dout    (fixTo_887_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_888 (
    .din     (_zz_3129[31:0]        ), //i
    .dout    (fixTo_888_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_889 (
    .din     (_zz_3130[31:0]        ), //i
    .dout    (fixTo_889_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_890 (
    .din     (_zz_3131[31:0]        ), //i
    .dout    (fixTo_890_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_891 (
    .din     (_zz_3132[31:0]        ), //i
    .dout    (fixTo_891_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_892 (
    .din     (_zz_3133[31:0]        ), //i
    .dout    (fixTo_892_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_893 (
    .din     (_zz_3134[31:0]        ), //i
    .dout    (fixTo_893_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_894 (
    .din     (_zz_3135[31:0]        ), //i
    .dout    (fixTo_894_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_895 (
    .din     (_zz_3136[31:0]        ), //i
    .dout    (fixTo_895_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_896 (
    .din     (_zz_3137[31:0]        ), //i
    .dout    (fixTo_896_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_897 (
    .din     (_zz_3138[31:0]        ), //i
    .dout    (fixTo_897_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_898 (
    .din     (_zz_3139[31:0]        ), //i
    .dout    (fixTo_898_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_899 (
    .din     (_zz_3140[31:0]        ), //i
    .dout    (fixTo_899_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_900 (
    .din     (_zz_3141[31:0]        ), //i
    .dout    (fixTo_900_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_901 (
    .din     (_zz_3142[31:0]        ), //i
    .dout    (fixTo_901_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_902 (
    .din     (_zz_3143[31:0]        ), //i
    .dout    (fixTo_902_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_903 (
    .din     (_zz_3144[31:0]        ), //i
    .dout    (fixTo_903_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_904 (
    .din     (_zz_3145[31:0]        ), //i
    .dout    (fixTo_904_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_905 (
    .din     (_zz_3146[31:0]        ), //i
    .dout    (fixTo_905_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_906 (
    .din     (_zz_3147[31:0]        ), //i
    .dout    (fixTo_906_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_907 (
    .din     (_zz_3148[31:0]        ), //i
    .dout    (fixTo_907_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_908 (
    .din     (_zz_3149[31:0]        ), //i
    .dout    (fixTo_908_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_909 (
    .din     (_zz_3150[31:0]        ), //i
    .dout    (fixTo_909_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_910 (
    .din     (_zz_3151[31:0]        ), //i
    .dout    (fixTo_910_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_911 (
    .din     (_zz_3152[31:0]        ), //i
    .dout    (fixTo_911_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_912 (
    .din     (_zz_3153[31:0]        ), //i
    .dout    (fixTo_912_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_913 (
    .din     (_zz_3154[31:0]        ), //i
    .dout    (fixTo_913_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_914 (
    .din     (_zz_3155[31:0]        ), //i
    .dout    (fixTo_914_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_915 (
    .din     (_zz_3156[31:0]        ), //i
    .dout    (fixTo_915_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_916 (
    .din     (_zz_3157[31:0]        ), //i
    .dout    (fixTo_916_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_917 (
    .din     (_zz_3158[31:0]        ), //i
    .dout    (fixTo_917_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_918 (
    .din     (_zz_3159[31:0]        ), //i
    .dout    (fixTo_918_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_919 (
    .din     (_zz_3160[31:0]        ), //i
    .dout    (fixTo_919_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_920 (
    .din     (_zz_3161[31:0]        ), //i
    .dout    (fixTo_920_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_921 (
    .din     (_zz_3162[31:0]        ), //i
    .dout    (fixTo_921_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_922 (
    .din     (_zz_3163[31:0]        ), //i
    .dout    (fixTo_922_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_923 (
    .din     (_zz_3164[31:0]        ), //i
    .dout    (fixTo_923_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_924 (
    .din     (_zz_3165[31:0]        ), //i
    .dout    (fixTo_924_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_925 (
    .din     (_zz_3166[31:0]        ), //i
    .dout    (fixTo_925_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_926 (
    .din     (_zz_3167[31:0]        ), //i
    .dout    (fixTo_926_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_927 (
    .din     (_zz_3168[31:0]        ), //i
    .dout    (fixTo_927_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_928 (
    .din     (_zz_3169[31:0]        ), //i
    .dout    (fixTo_928_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_929 (
    .din     (_zz_3170[31:0]        ), //i
    .dout    (fixTo_929_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_930 (
    .din     (_zz_3171[31:0]        ), //i
    .dout    (fixTo_930_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_931 (
    .din     (_zz_3172[31:0]        ), //i
    .dout    (fixTo_931_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_932 (
    .din     (_zz_3173[31:0]        ), //i
    .dout    (fixTo_932_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_933 (
    .din     (_zz_3174[31:0]        ), //i
    .dout    (fixTo_933_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_934 (
    .din     (_zz_3175[31:0]        ), //i
    .dout    (fixTo_934_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_935 (
    .din     (_zz_3176[31:0]        ), //i
    .dout    (fixTo_935_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_936 (
    .din     (_zz_3177[31:0]        ), //i
    .dout    (fixTo_936_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_937 (
    .din     (_zz_3178[31:0]        ), //i
    .dout    (fixTo_937_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_938 (
    .din     (_zz_3179[31:0]        ), //i
    .dout    (fixTo_938_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_939 (
    .din     (_zz_3180[31:0]        ), //i
    .dout    (fixTo_939_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_940 (
    .din     (_zz_3181[31:0]        ), //i
    .dout    (fixTo_940_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_941 (
    .din     (_zz_3182[31:0]        ), //i
    .dout    (fixTo_941_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_942 (
    .din     (_zz_3183[31:0]        ), //i
    .dout    (fixTo_942_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_943 (
    .din     (_zz_3184[31:0]        ), //i
    .dout    (fixTo_943_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_944 (
    .din     (_zz_3185[31:0]        ), //i
    .dout    (fixTo_944_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_945 (
    .din     (_zz_3186[31:0]        ), //i
    .dout    (fixTo_945_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_946 (
    .din     (_zz_3187[31:0]        ), //i
    .dout    (fixTo_946_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_947 (
    .din     (_zz_3188[31:0]        ), //i
    .dout    (fixTo_947_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_948 (
    .din     (_zz_3189[31:0]        ), //i
    .dout    (fixTo_948_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_949 (
    .din     (_zz_3190[31:0]        ), //i
    .dout    (fixTo_949_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_950 (
    .din     (_zz_3191[31:0]        ), //i
    .dout    (fixTo_950_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_951 (
    .din     (_zz_3192[31:0]        ), //i
    .dout    (fixTo_951_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_952 (
    .din     (_zz_3193[31:0]        ), //i
    .dout    (fixTo_952_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_953 (
    .din     (_zz_3194[31:0]        ), //i
    .dout    (fixTo_953_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_954 (
    .din     (_zz_3195[31:0]        ), //i
    .dout    (fixTo_954_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_955 (
    .din     (_zz_3196[31:0]        ), //i
    .dout    (fixTo_955_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_956 (
    .din     (_zz_3197[31:0]        ), //i
    .dout    (fixTo_956_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_957 (
    .din     (_zz_3198[31:0]        ), //i
    .dout    (fixTo_957_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_958 (
    .din     (_zz_3199[31:0]        ), //i
    .dout    (fixTo_958_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_959 (
    .din     (_zz_3200[31:0]        ), //i
    .dout    (fixTo_959_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_960 (
    .din     (_zz_3201[31:0]        ), //i
    .dout    (fixTo_960_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_961 (
    .din     (_zz_3202[31:0]        ), //i
    .dout    (fixTo_961_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_962 (
    .din     (_zz_3203[31:0]        ), //i
    .dout    (fixTo_962_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_963 (
    .din     (_zz_3204[31:0]        ), //i
    .dout    (fixTo_963_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_964 (
    .din     (_zz_3205[31:0]        ), //i
    .dout    (fixTo_964_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_965 (
    .din     (_zz_3206[31:0]        ), //i
    .dout    (fixTo_965_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_966 (
    .din     (_zz_3207[31:0]        ), //i
    .dout    (fixTo_966_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_967 (
    .din     (_zz_3208[31:0]        ), //i
    .dout    (fixTo_967_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_968 (
    .din     (_zz_3209[31:0]        ), //i
    .dout    (fixTo_968_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_969 (
    .din     (_zz_3210[31:0]        ), //i
    .dout    (fixTo_969_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_970 (
    .din     (_zz_3211[31:0]        ), //i
    .dout    (fixTo_970_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_971 (
    .din     (_zz_3212[31:0]        ), //i
    .dout    (fixTo_971_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_972 (
    .din     (_zz_3213[31:0]        ), //i
    .dout    (fixTo_972_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_973 (
    .din     (_zz_3214[31:0]        ), //i
    .dout    (fixTo_973_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_974 (
    .din     (_zz_3215[31:0]        ), //i
    .dout    (fixTo_974_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_975 (
    .din     (_zz_3216[31:0]        ), //i
    .dout    (fixTo_975_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_976 (
    .din     (_zz_3217[31:0]        ), //i
    .dout    (fixTo_976_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_977 (
    .din     (_zz_3218[31:0]        ), //i
    .dout    (fixTo_977_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_978 (
    .din     (_zz_3219[31:0]        ), //i
    .dout    (fixTo_978_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_979 (
    .din     (_zz_3220[31:0]        ), //i
    .dout    (fixTo_979_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_980 (
    .din     (_zz_3221[31:0]        ), //i
    .dout    (fixTo_980_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_981 (
    .din     (_zz_3222[31:0]        ), //i
    .dout    (fixTo_981_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_982 (
    .din     (_zz_3223[31:0]        ), //i
    .dout    (fixTo_982_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_983 (
    .din     (_zz_3224[31:0]        ), //i
    .dout    (fixTo_983_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_984 (
    .din     (_zz_3225[31:0]        ), //i
    .dout    (fixTo_984_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_985 (
    .din     (_zz_3226[31:0]        ), //i
    .dout    (fixTo_985_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_986 (
    .din     (_zz_3227[31:0]        ), //i
    .dout    (fixTo_986_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_987 (
    .din     (_zz_3228[31:0]        ), //i
    .dout    (fixTo_987_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_988 (
    .din     (_zz_3229[31:0]        ), //i
    .dout    (fixTo_988_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_989 (
    .din     (_zz_3230[31:0]        ), //i
    .dout    (fixTo_989_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_990 (
    .din     (_zz_3231[31:0]        ), //i
    .dout    (fixTo_990_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_991 (
    .din     (_zz_3232[31:0]        ), //i
    .dout    (fixTo_991_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_992 (
    .din     (_zz_3233[31:0]        ), //i
    .dout    (fixTo_992_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_993 (
    .din     (_zz_3234[31:0]        ), //i
    .dout    (fixTo_993_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_994 (
    .din     (_zz_3235[31:0]        ), //i
    .dout    (fixTo_994_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_995 (
    .din     (_zz_3236[31:0]        ), //i
    .dout    (fixTo_995_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_996 (
    .din     (_zz_3237[31:0]        ), //i
    .dout    (fixTo_996_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_997 (
    .din     (_zz_3238[31:0]        ), //i
    .dout    (fixTo_997_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_998 (
    .din     (_zz_3239[31:0]        ), //i
    .dout    (fixTo_998_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_999 (
    .din     (_zz_3240[31:0]        ), //i
    .dout    (fixTo_999_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1000 (
    .din     (_zz_3241[31:0]         ), //i
    .dout    (fixTo_1000_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1001 (
    .din     (_zz_3242[31:0]         ), //i
    .dout    (fixTo_1001_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_1002 (
    .din     (_zz_3243[31:0]         ), //i
    .dout    (fixTo_1002_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_1003 (
    .din     (_zz_3244[31:0]         ), //i
    .dout    (fixTo_1003_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1004 (
    .din     (_zz_3245[31:0]         ), //i
    .dout    (fixTo_1004_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1005 (
    .din     (_zz_3246[31:0]         ), //i
    .dout    (fixTo_1005_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1006 (
    .din     (_zz_3247[31:0]         ), //i
    .dout    (fixTo_1006_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1007 (
    .din     (_zz_3248[31:0]         ), //i
    .dout    (fixTo_1007_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_1008 (
    .din     (_zz_3249[31:0]         ), //i
    .dout    (fixTo_1008_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_1009 (
    .din     (_zz_3250[31:0]         ), //i
    .dout    (fixTo_1009_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1010 (
    .din     (_zz_3251[31:0]         ), //i
    .dout    (fixTo_1010_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1011 (
    .din     (_zz_3252[31:0]         ), //i
    .dout    (fixTo_1011_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1012 (
    .din     (_zz_3253[31:0]         ), //i
    .dout    (fixTo_1012_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1013 (
    .din     (_zz_3254[31:0]         ), //i
    .dout    (fixTo_1013_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_1014 (
    .din     (_zz_3255[31:0]         ), //i
    .dout    (fixTo_1014_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_1015 (
    .din     (_zz_3256[31:0]         ), //i
    .dout    (fixTo_1015_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1016 (
    .din     (_zz_3257[31:0]         ), //i
    .dout    (fixTo_1016_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1017 (
    .din     (_zz_3258[31:0]         ), //i
    .dout    (fixTo_1017_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1018 (
    .din     (_zz_3259[31:0]         ), //i
    .dout    (fixTo_1018_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1019 (
    .din     (_zz_3260[31:0]         ), //i
    .dout    (fixTo_1019_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_1020 (
    .din     (_zz_3261[31:0]         ), //i
    .dout    (fixTo_1020_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_1021 (
    .din     (_zz_3262[31:0]         ), //i
    .dout    (fixTo_1021_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1022 (
    .din     (_zz_3263[31:0]         ), //i
    .dout    (fixTo_1022_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1023 (
    .din     (_zz_3264[31:0]         ), //i
    .dout    (fixTo_1023_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1024 (
    .din     (_zz_3265[31:0]         ), //i
    .dout    (fixTo_1024_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1025 (
    .din     (_zz_3266[31:0]         ), //i
    .dout    (fixTo_1025_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_1026 (
    .din     (_zz_3267[31:0]         ), //i
    .dout    (fixTo_1026_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_1027 (
    .din     (_zz_3268[31:0]         ), //i
    .dout    (fixTo_1027_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1028 (
    .din     (_zz_3269[31:0]         ), //i
    .dout    (fixTo_1028_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1029 (
    .din     (_zz_3270[31:0]         ), //i
    .dout    (fixTo_1029_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1030 (
    .din     (_zz_3271[31:0]         ), //i
    .dout    (fixTo_1030_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1031 (
    .din     (_zz_3272[31:0]         ), //i
    .dout    (fixTo_1031_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_1032 (
    .din     (_zz_3273[31:0]         ), //i
    .dout    (fixTo_1032_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_1033 (
    .din     (_zz_3274[31:0]         ), //i
    .dout    (fixTo_1033_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1034 (
    .din     (_zz_3275[31:0]         ), //i
    .dout    (fixTo_1034_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1035 (
    .din     (_zz_3276[31:0]         ), //i
    .dout    (fixTo_1035_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1036 (
    .din     (_zz_3277[31:0]         ), //i
    .dout    (fixTo_1036_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1037 (
    .din     (_zz_3278[31:0]         ), //i
    .dout    (fixTo_1037_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_1038 (
    .din     (_zz_3279[31:0]         ), //i
    .dout    (fixTo_1038_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_1039 (
    .din     (_zz_3280[31:0]         ), //i
    .dout    (fixTo_1039_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1040 (
    .din     (_zz_3281[31:0]         ), //i
    .dout    (fixTo_1040_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1041 (
    .din     (_zz_3282[31:0]         ), //i
    .dout    (fixTo_1041_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1042 (
    .din     (_zz_3283[31:0]         ), //i
    .dout    (fixTo_1042_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1043 (
    .din     (_zz_3284[31:0]         ), //i
    .dout    (fixTo_1043_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_1044 (
    .din     (_zz_3285[31:0]         ), //i
    .dout    (fixTo_1044_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_1045 (
    .din     (_zz_3286[31:0]         ), //i
    .dout    (fixTo_1045_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1046 (
    .din     (_zz_3287[31:0]         ), //i
    .dout    (fixTo_1046_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1047 (
    .din     (_zz_3288[31:0]         ), //i
    .dout    (fixTo_1047_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1048 (
    .din     (_zz_3289[31:0]         ), //i
    .dout    (fixTo_1048_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1049 (
    .din     (_zz_3290[31:0]         ), //i
    .dout    (fixTo_1049_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_1050 (
    .din     (_zz_3291[31:0]         ), //i
    .dout    (fixTo_1050_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_1051 (
    .din     (_zz_3292[31:0]         ), //i
    .dout    (fixTo_1051_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1052 (
    .din     (_zz_3293[31:0]         ), //i
    .dout    (fixTo_1052_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1053 (
    .din     (_zz_3294[31:0]         ), //i
    .dout    (fixTo_1053_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1054 (
    .din     (_zz_3295[31:0]         ), //i
    .dout    (fixTo_1054_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1055 (
    .din     (_zz_3296[31:0]         ), //i
    .dout    (fixTo_1055_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_1056 (
    .din     (_zz_3297[31:0]         ), //i
    .dout    (fixTo_1056_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_1057 (
    .din     (_zz_3298[31:0]         ), //i
    .dout    (fixTo_1057_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1058 (
    .din     (_zz_3299[31:0]         ), //i
    .dout    (fixTo_1058_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1059 (
    .din     (_zz_3300[31:0]         ), //i
    .dout    (fixTo_1059_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1060 (
    .din     (_zz_3301[31:0]         ), //i
    .dout    (fixTo_1060_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1061 (
    .din     (_zz_3302[31:0]         ), //i
    .dout    (fixTo_1061_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_1062 (
    .din     (_zz_3303[31:0]         ), //i
    .dout    (fixTo_1062_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_1063 (
    .din     (_zz_3304[31:0]         ), //i
    .dout    (fixTo_1063_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1064 (
    .din     (_zz_3305[31:0]         ), //i
    .dout    (fixTo_1064_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1065 (
    .din     (_zz_3306[31:0]         ), //i
    .dout    (fixTo_1065_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1066 (
    .din     (_zz_3307[31:0]         ), //i
    .dout    (fixTo_1066_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1067 (
    .din     (_zz_3308[31:0]         ), //i
    .dout    (fixTo_1067_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_1068 (
    .din     (_zz_3309[31:0]         ), //i
    .dout    (fixTo_1068_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_1069 (
    .din     (_zz_3310[31:0]         ), //i
    .dout    (fixTo_1069_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1070 (
    .din     (_zz_3311[31:0]         ), //i
    .dout    (fixTo_1070_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1071 (
    .din     (_zz_3312[31:0]         ), //i
    .dout    (fixTo_1071_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1072 (
    .din     (_zz_3313[31:0]         ), //i
    .dout    (fixTo_1072_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1073 (
    .din     (_zz_3314[31:0]         ), //i
    .dout    (fixTo_1073_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_1074 (
    .din     (_zz_3315[31:0]         ), //i
    .dout    (fixTo_1074_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_1075 (
    .din     (_zz_3316[31:0]         ), //i
    .dout    (fixTo_1075_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1076 (
    .din     (_zz_3317[31:0]         ), //i
    .dout    (fixTo_1076_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1077 (
    .din     (_zz_3318[31:0]         ), //i
    .dout    (fixTo_1077_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1078 (
    .din     (_zz_3319[31:0]         ), //i
    .dout    (fixTo_1078_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1079 (
    .din     (_zz_3320[31:0]         ), //i
    .dout    (fixTo_1079_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_1080 (
    .din     (_zz_3321[31:0]         ), //i
    .dout    (fixTo_1080_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_1081 (
    .din     (_zz_3322[31:0]         ), //i
    .dout    (fixTo_1081_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1082 (
    .din     (_zz_3323[31:0]         ), //i
    .dout    (fixTo_1082_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1083 (
    .din     (_zz_3324[31:0]         ), //i
    .dout    (fixTo_1083_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1084 (
    .din     (_zz_3325[31:0]         ), //i
    .dout    (fixTo_1084_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1085 (
    .din     (_zz_3326[31:0]         ), //i
    .dout    (fixTo_1085_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_1086 (
    .din     (_zz_3327[31:0]         ), //i
    .dout    (fixTo_1086_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_1087 (
    .din     (_zz_3328[31:0]         ), //i
    .dout    (fixTo_1087_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1088 (
    .din     (_zz_3329[31:0]         ), //i
    .dout    (fixTo_1088_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1089 (
    .din     (_zz_3330[31:0]         ), //i
    .dout    (fixTo_1089_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1090 (
    .din     (_zz_3331[31:0]         ), //i
    .dout    (fixTo_1090_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1091 (
    .din     (_zz_3332[31:0]         ), //i
    .dout    (fixTo_1091_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_1092 (
    .din     (_zz_3333[31:0]         ), //i
    .dout    (fixTo_1092_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_1093 (
    .din     (_zz_3334[31:0]         ), //i
    .dout    (fixTo_1093_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1094 (
    .din     (_zz_3335[31:0]         ), //i
    .dout    (fixTo_1094_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1095 (
    .din     (_zz_3336[31:0]         ), //i
    .dout    (fixTo_1095_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1096 (
    .din     (_zz_3337[31:0]         ), //i
    .dout    (fixTo_1096_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1097 (
    .din     (_zz_3338[31:0]         ), //i
    .dout    (fixTo_1097_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_1098 (
    .din     (_zz_3339[31:0]         ), //i
    .dout    (fixTo_1098_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_1099 (
    .din     (_zz_3340[31:0]         ), //i
    .dout    (fixTo_1099_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1100 (
    .din     (_zz_3341[31:0]         ), //i
    .dout    (fixTo_1100_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1101 (
    .din     (_zz_3342[31:0]         ), //i
    .dout    (fixTo_1101_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1102 (
    .din     (_zz_3343[31:0]         ), //i
    .dout    (fixTo_1102_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1103 (
    .din     (_zz_3344[31:0]         ), //i
    .dout    (fixTo_1103_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_1104 (
    .din     (_zz_3345[31:0]         ), //i
    .dout    (fixTo_1104_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_1105 (
    .din     (_zz_3346[31:0]         ), //i
    .dout    (fixTo_1105_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1106 (
    .din     (_zz_3347[31:0]         ), //i
    .dout    (fixTo_1106_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1107 (
    .din     (_zz_3348[31:0]         ), //i
    .dout    (fixTo_1107_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1108 (
    .din     (_zz_3349[31:0]         ), //i
    .dout    (fixTo_1108_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1109 (
    .din     (_zz_3350[31:0]         ), //i
    .dout    (fixTo_1109_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_1110 (
    .din     (_zz_3351[31:0]         ), //i
    .dout    (fixTo_1110_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_1111 (
    .din     (_zz_3352[31:0]         ), //i
    .dout    (fixTo_1111_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1112 (
    .din     (_zz_3353[31:0]         ), //i
    .dout    (fixTo_1112_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1113 (
    .din     (_zz_3354[31:0]         ), //i
    .dout    (fixTo_1113_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1114 (
    .din     (_zz_3355[31:0]         ), //i
    .dout    (fixTo_1114_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1115 (
    .din     (_zz_3356[31:0]         ), //i
    .dout    (fixTo_1115_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_1116 (
    .din     (_zz_3357[31:0]         ), //i
    .dout    (fixTo_1116_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_1117 (
    .din     (_zz_3358[31:0]         ), //i
    .dout    (fixTo_1117_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1118 (
    .din     (_zz_3359[31:0]         ), //i
    .dout    (fixTo_1118_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1119 (
    .din     (_zz_3360[31:0]         ), //i
    .dout    (fixTo_1119_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1120 (
    .din     (_zz_3361[31:0]         ), //i
    .dout    (fixTo_1120_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1121 (
    .din     (_zz_3362[31:0]         ), //i
    .dout    (fixTo_1121_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_1122 (
    .din     (_zz_3363[31:0]         ), //i
    .dout    (fixTo_1122_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_1123 (
    .din     (_zz_3364[31:0]         ), //i
    .dout    (fixTo_1123_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1124 (
    .din     (_zz_3365[31:0]         ), //i
    .dout    (fixTo_1124_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1125 (
    .din     (_zz_3366[31:0]         ), //i
    .dout    (fixTo_1125_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1126 (
    .din     (_zz_3367[31:0]         ), //i
    .dout    (fixTo_1126_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1127 (
    .din     (_zz_3368[31:0]         ), //i
    .dout    (fixTo_1127_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_1128 (
    .din     (_zz_3369[31:0]         ), //i
    .dout    (fixTo_1128_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_1129 (
    .din     (_zz_3370[31:0]         ), //i
    .dout    (fixTo_1129_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1130 (
    .din     (_zz_3371[31:0]         ), //i
    .dout    (fixTo_1130_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1131 (
    .din     (_zz_3372[31:0]         ), //i
    .dout    (fixTo_1131_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1132 (
    .din     (_zz_3373[31:0]         ), //i
    .dout    (fixTo_1132_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1133 (
    .din     (_zz_3374[31:0]         ), //i
    .dout    (fixTo_1133_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_1134 (
    .din     (_zz_3375[31:0]         ), //i
    .dout    (fixTo_1134_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_1135 (
    .din     (_zz_3376[31:0]         ), //i
    .dout    (fixTo_1135_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1136 (
    .din     (_zz_3377[31:0]         ), //i
    .dout    (fixTo_1136_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1137 (
    .din     (_zz_3378[31:0]         ), //i
    .dout    (fixTo_1137_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1138 (
    .din     (_zz_3379[31:0]         ), //i
    .dout    (fixTo_1138_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1139 (
    .din     (_zz_3380[31:0]         ), //i
    .dout    (fixTo_1139_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_1140 (
    .din     (_zz_3381[31:0]         ), //i
    .dout    (fixTo_1140_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_1141 (
    .din     (_zz_3382[31:0]         ), //i
    .dout    (fixTo_1141_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1142 (
    .din     (_zz_3383[31:0]         ), //i
    .dout    (fixTo_1142_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1143 (
    .din     (_zz_3384[31:0]         ), //i
    .dout    (fixTo_1143_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1144 (
    .din     (_zz_3385[31:0]         ), //i
    .dout    (fixTo_1144_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1145 (
    .din     (_zz_3386[31:0]         ), //i
    .dout    (fixTo_1145_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_1146 (
    .din     (_zz_3387[31:0]         ), //i
    .dout    (fixTo_1146_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_1147 (
    .din     (_zz_3388[31:0]         ), //i
    .dout    (fixTo_1147_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1148 (
    .din     (_zz_3389[31:0]         ), //i
    .dout    (fixTo_1148_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1149 (
    .din     (_zz_3390[31:0]         ), //i
    .dout    (fixTo_1149_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1150 (
    .din     (_zz_3391[31:0]         ), //i
    .dout    (fixTo_1150_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1151 (
    .din     (_zz_3392[31:0]         ), //i
    .dout    (fixTo_1151_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_1152 (
    .din     (_zz_3393[31:0]         ), //i
    .dout    (fixTo_1152_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_1153 (
    .din     (_zz_3394[31:0]         ), //i
    .dout    (fixTo_1153_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1154 (
    .din     (_zz_3395[31:0]         ), //i
    .dout    (fixTo_1154_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1155 (
    .din     (_zz_3396[31:0]         ), //i
    .dout    (fixTo_1155_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1156 (
    .din     (_zz_3397[31:0]         ), //i
    .dout    (fixTo_1156_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1157 (
    .din     (_zz_3398[31:0]         ), //i
    .dout    (fixTo_1157_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_1158 (
    .din     (_zz_3399[31:0]         ), //i
    .dout    (fixTo_1158_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_1159 (
    .din     (_zz_3400[31:0]         ), //i
    .dout    (fixTo_1159_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1160 (
    .din     (_zz_3401[31:0]         ), //i
    .dout    (fixTo_1160_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1161 (
    .din     (_zz_3402[31:0]         ), //i
    .dout    (fixTo_1161_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1162 (
    .din     (_zz_3403[31:0]         ), //i
    .dout    (fixTo_1162_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1163 (
    .din     (_zz_3404[31:0]         ), //i
    .dout    (fixTo_1163_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_1164 (
    .din     (_zz_3405[31:0]         ), //i
    .dout    (fixTo_1164_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_1165 (
    .din     (_zz_3406[31:0]         ), //i
    .dout    (fixTo_1165_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1166 (
    .din     (_zz_3407[31:0]         ), //i
    .dout    (fixTo_1166_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1167 (
    .din     (_zz_3408[31:0]         ), //i
    .dout    (fixTo_1167_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1168 (
    .din     (_zz_3409[31:0]         ), //i
    .dout    (fixTo_1168_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1169 (
    .din     (_zz_3410[31:0]         ), //i
    .dout    (fixTo_1169_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_1170 (
    .din     (_zz_3411[31:0]         ), //i
    .dout    (fixTo_1170_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_1171 (
    .din     (_zz_3412[31:0]         ), //i
    .dout    (fixTo_1171_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1172 (
    .din     (_zz_3413[31:0]         ), //i
    .dout    (fixTo_1172_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1173 (
    .din     (_zz_3414[31:0]         ), //i
    .dout    (fixTo_1173_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1174 (
    .din     (_zz_3415[31:0]         ), //i
    .dout    (fixTo_1174_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1175 (
    .din     (_zz_3416[31:0]         ), //i
    .dout    (fixTo_1175_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_1176 (
    .din     (_zz_3417[31:0]         ), //i
    .dout    (fixTo_1176_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_1177 (
    .din     (_zz_3418[31:0]         ), //i
    .dout    (fixTo_1177_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1178 (
    .din     (_zz_3419[31:0]         ), //i
    .dout    (fixTo_1178_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1179 (
    .din     (_zz_3420[31:0]         ), //i
    .dout    (fixTo_1179_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1180 (
    .din     (_zz_3421[31:0]         ), //i
    .dout    (fixTo_1180_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1181 (
    .din     (_zz_3422[31:0]         ), //i
    .dout    (fixTo_1181_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_1182 (
    .din     (_zz_3423[31:0]         ), //i
    .dout    (fixTo_1182_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_1183 (
    .din     (_zz_3424[31:0]         ), //i
    .dout    (fixTo_1183_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1184 (
    .din     (_zz_3425[31:0]         ), //i
    .dout    (fixTo_1184_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1185 (
    .din     (_zz_3426[31:0]         ), //i
    .dout    (fixTo_1185_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1186 (
    .din     (_zz_3427[31:0]         ), //i
    .dout    (fixTo_1186_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1187 (
    .din     (_zz_3428[31:0]         ), //i
    .dout    (fixTo_1187_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_1188 (
    .din     (_zz_3429[31:0]         ), //i
    .dout    (fixTo_1188_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_1189 (
    .din     (_zz_3430[31:0]         ), //i
    .dout    (fixTo_1189_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1190 (
    .din     (_zz_3431[31:0]         ), //i
    .dout    (fixTo_1190_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1191 (
    .din     (_zz_3432[31:0]         ), //i
    .dout    (fixTo_1191_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1192 (
    .din     (_zz_3433[31:0]         ), //i
    .dout    (fixTo_1192_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1193 (
    .din     (_zz_3434[31:0]         ), //i
    .dout    (fixTo_1193_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_1194 (
    .din     (_zz_3435[31:0]         ), //i
    .dout    (fixTo_1194_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_1195 (
    .din     (_zz_3436[31:0]         ), //i
    .dout    (fixTo_1195_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1196 (
    .din     (_zz_3437[31:0]         ), //i
    .dout    (fixTo_1196_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1197 (
    .din     (_zz_3438[31:0]         ), //i
    .dout    (fixTo_1197_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1198 (
    .din     (_zz_3439[31:0]         ), //i
    .dout    (fixTo_1198_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1199 (
    .din     (_zz_3440[31:0]         ), //i
    .dout    (fixTo_1199_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_1200 (
    .din     (_zz_3441[31:0]         ), //i
    .dout    (fixTo_1200_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_1201 (
    .din     (_zz_3442[31:0]         ), //i
    .dout    (fixTo_1201_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1202 (
    .din     (_zz_3443[31:0]         ), //i
    .dout    (fixTo_1202_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1203 (
    .din     (_zz_3444[31:0]         ), //i
    .dout    (fixTo_1203_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1204 (
    .din     (_zz_3445[31:0]         ), //i
    .dout    (fixTo_1204_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1205 (
    .din     (_zz_3446[31:0]         ), //i
    .dout    (fixTo_1205_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_1206 (
    .din     (_zz_3447[31:0]         ), //i
    .dout    (fixTo_1206_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_1207 (
    .din     (_zz_3448[31:0]         ), //i
    .dout    (fixTo_1207_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1208 (
    .din     (_zz_3449[31:0]         ), //i
    .dout    (fixTo_1208_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1209 (
    .din     (_zz_3450[31:0]         ), //i
    .dout    (fixTo_1209_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1210 (
    .din     (_zz_3451[31:0]         ), //i
    .dout    (fixTo_1210_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1211 (
    .din     (_zz_3452[31:0]         ), //i
    .dout    (fixTo_1211_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_1212 (
    .din     (_zz_3453[31:0]         ), //i
    .dout    (fixTo_1212_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_1213 (
    .din     (_zz_3454[31:0]         ), //i
    .dout    (fixTo_1213_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1214 (
    .din     (_zz_3455[31:0]         ), //i
    .dout    (fixTo_1214_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1215 (
    .din     (_zz_3456[31:0]         ), //i
    .dout    (fixTo_1215_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1216 (
    .din     (_zz_3457[31:0]         ), //i
    .dout    (fixTo_1216_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1217 (
    .din     (_zz_3458[31:0]         ), //i
    .dout    (fixTo_1217_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_1218 (
    .din     (_zz_3459[31:0]         ), //i
    .dout    (fixTo_1218_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_1219 (
    .din     (_zz_3460[31:0]         ), //i
    .dout    (fixTo_1219_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1220 (
    .din     (_zz_3461[31:0]         ), //i
    .dout    (fixTo_1220_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1221 (
    .din     (_zz_3462[31:0]         ), //i
    .dout    (fixTo_1221_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1222 (
    .din     (_zz_3463[31:0]         ), //i
    .dout    (fixTo_1222_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1223 (
    .din     (_zz_3464[31:0]         ), //i
    .dout    (fixTo_1223_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_1224 (
    .din     (_zz_3465[31:0]         ), //i
    .dout    (fixTo_1224_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_1225 (
    .din     (_zz_3466[31:0]         ), //i
    .dout    (fixTo_1225_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1226 (
    .din     (_zz_3467[31:0]         ), //i
    .dout    (fixTo_1226_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1227 (
    .din     (_zz_3468[31:0]         ), //i
    .dout    (fixTo_1227_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1228 (
    .din     (_zz_3469[31:0]         ), //i
    .dout    (fixTo_1228_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1229 (
    .din     (_zz_3470[31:0]         ), //i
    .dout    (fixTo_1229_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_1230 (
    .din     (_zz_3471[31:0]         ), //i
    .dout    (fixTo_1230_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_1231 (
    .din     (_zz_3472[31:0]         ), //i
    .dout    (fixTo_1231_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1232 (
    .din     (_zz_3473[31:0]         ), //i
    .dout    (fixTo_1232_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1233 (
    .din     (_zz_3474[31:0]         ), //i
    .dout    (fixTo_1233_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1234 (
    .din     (_zz_3475[31:0]         ), //i
    .dout    (fixTo_1234_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1235 (
    .din     (_zz_3476[31:0]         ), //i
    .dout    (fixTo_1235_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_1236 (
    .din     (_zz_3477[31:0]         ), //i
    .dout    (fixTo_1236_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_1237 (
    .din     (_zz_3478[31:0]         ), //i
    .dout    (fixTo_1237_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1238 (
    .din     (_zz_3479[31:0]         ), //i
    .dout    (fixTo_1238_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1239 (
    .din     (_zz_3480[31:0]         ), //i
    .dout    (fixTo_1239_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1240 (
    .din     (_zz_3481[31:0]         ), //i
    .dout    (fixTo_1240_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1241 (
    .din     (_zz_3482[31:0]         ), //i
    .dout    (fixTo_1241_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_1242 (
    .din     (_zz_3483[31:0]         ), //i
    .dout    (fixTo_1242_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_1243 (
    .din     (_zz_3484[31:0]         ), //i
    .dout    (fixTo_1243_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1244 (
    .din     (_zz_3485[31:0]         ), //i
    .dout    (fixTo_1244_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1245 (
    .din     (_zz_3486[31:0]         ), //i
    .dout    (fixTo_1245_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1246 (
    .din     (_zz_3487[31:0]         ), //i
    .dout    (fixTo_1246_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1247 (
    .din     (_zz_3488[31:0]         ), //i
    .dout    (fixTo_1247_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_1248 (
    .din     (_zz_3489[31:0]         ), //i
    .dout    (fixTo_1248_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_1249 (
    .din     (_zz_3490[31:0]         ), //i
    .dout    (fixTo_1249_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1250 (
    .din     (_zz_3491[31:0]         ), //i
    .dout    (fixTo_1250_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1251 (
    .din     (_zz_3492[31:0]         ), //i
    .dout    (fixTo_1251_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1252 (
    .din     (_zz_3493[31:0]         ), //i
    .dout    (fixTo_1252_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1253 (
    .din     (_zz_3494[31:0]         ), //i
    .dout    (fixTo_1253_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_1254 (
    .din     (_zz_3495[31:0]         ), //i
    .dout    (fixTo_1254_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_1255 (
    .din     (_zz_3496[31:0]         ), //i
    .dout    (fixTo_1255_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1256 (
    .din     (_zz_3497[31:0]         ), //i
    .dout    (fixTo_1256_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1257 (
    .din     (_zz_3498[31:0]         ), //i
    .dout    (fixTo_1257_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1258 (
    .din     (_zz_3499[31:0]         ), //i
    .dout    (fixTo_1258_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1259 (
    .din     (_zz_3500[31:0]         ), //i
    .dout    (fixTo_1259_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_1260 (
    .din     (_zz_3501[31:0]         ), //i
    .dout    (fixTo_1260_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_1261 (
    .din     (_zz_3502[31:0]         ), //i
    .dout    (fixTo_1261_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1262 (
    .din     (_zz_3503[31:0]         ), //i
    .dout    (fixTo_1262_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1263 (
    .din     (_zz_3504[31:0]         ), //i
    .dout    (fixTo_1263_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1264 (
    .din     (_zz_3505[31:0]         ), //i
    .dout    (fixTo_1264_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1265 (
    .din     (_zz_3506[31:0]         ), //i
    .dout    (fixTo_1265_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_1266 (
    .din     (_zz_3507[31:0]         ), //i
    .dout    (fixTo_1266_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_1267 (
    .din     (_zz_3508[31:0]         ), //i
    .dout    (fixTo_1267_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1268 (
    .din     (_zz_3509[31:0]         ), //i
    .dout    (fixTo_1268_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1269 (
    .din     (_zz_3510[31:0]         ), //i
    .dout    (fixTo_1269_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1270 (
    .din     (_zz_3511[31:0]         ), //i
    .dout    (fixTo_1270_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1271 (
    .din     (_zz_3512[31:0]         ), //i
    .dout    (fixTo_1271_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_1272 (
    .din     (_zz_3513[31:0]         ), //i
    .dout    (fixTo_1272_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_1273 (
    .din     (_zz_3514[31:0]         ), //i
    .dout    (fixTo_1273_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1274 (
    .din     (_zz_3515[31:0]         ), //i
    .dout    (fixTo_1274_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1275 (
    .din     (_zz_3516[31:0]         ), //i
    .dout    (fixTo_1275_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1276 (
    .din     (_zz_3517[31:0]         ), //i
    .dout    (fixTo_1276_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1277 (
    .din     (_zz_3518[31:0]         ), //i
    .dout    (fixTo_1277_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_1278 (
    .din     (_zz_3519[31:0]         ), //i
    .dout    (fixTo_1278_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_1279 (
    .din     (_zz_3520[31:0]         ), //i
    .dout    (fixTo_1279_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1280 (
    .din     (_zz_3521[31:0]         ), //i
    .dout    (fixTo_1280_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1281 (
    .din     (_zz_3522[31:0]         ), //i
    .dout    (fixTo_1281_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1282 (
    .din     (_zz_3523[31:0]         ), //i
    .dout    (fixTo_1282_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1283 (
    .din     (_zz_3524[31:0]         ), //i
    .dout    (fixTo_1283_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_1284 (
    .din     (_zz_3525[31:0]         ), //i
    .dout    (fixTo_1284_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_1285 (
    .din     (_zz_3526[31:0]         ), //i
    .dout    (fixTo_1285_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1286 (
    .din     (_zz_3527[31:0]         ), //i
    .dout    (fixTo_1286_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1287 (
    .din     (_zz_3528[31:0]         ), //i
    .dout    (fixTo_1287_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1288 (
    .din     (_zz_3529[31:0]         ), //i
    .dout    (fixTo_1288_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1289 (
    .din     (_zz_3530[31:0]         ), //i
    .dout    (fixTo_1289_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_1290 (
    .din     (_zz_3531[31:0]         ), //i
    .dout    (fixTo_1290_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_1291 (
    .din     (_zz_3532[31:0]         ), //i
    .dout    (fixTo_1291_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1292 (
    .din     (_zz_3533[31:0]         ), //i
    .dout    (fixTo_1292_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1293 (
    .din     (_zz_3534[31:0]         ), //i
    .dout    (fixTo_1293_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1294 (
    .din     (_zz_3535[31:0]         ), //i
    .dout    (fixTo_1294_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1295 (
    .din     (_zz_3536[31:0]         ), //i
    .dout    (fixTo_1295_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_1296 (
    .din     (_zz_3537[31:0]         ), //i
    .dout    (fixTo_1296_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_1297 (
    .din     (_zz_3538[31:0]         ), //i
    .dout    (fixTo_1297_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1298 (
    .din     (_zz_3539[31:0]         ), //i
    .dout    (fixTo_1298_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1299 (
    .din     (_zz_3540[31:0]         ), //i
    .dout    (fixTo_1299_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1300 (
    .din     (_zz_3541[31:0]         ), //i
    .dout    (fixTo_1300_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1301 (
    .din     (_zz_3542[31:0]         ), //i
    .dout    (fixTo_1301_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_1302 (
    .din     (_zz_3543[31:0]         ), //i
    .dout    (fixTo_1302_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_1303 (
    .din     (_zz_3544[31:0]         ), //i
    .dout    (fixTo_1303_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1304 (
    .din     (_zz_3545[31:0]         ), //i
    .dout    (fixTo_1304_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1305 (
    .din     (_zz_3546[31:0]         ), //i
    .dout    (fixTo_1305_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1306 (
    .din     (_zz_3547[31:0]         ), //i
    .dout    (fixTo_1306_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1307 (
    .din     (_zz_3548[31:0]         ), //i
    .dout    (fixTo_1307_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_1308 (
    .din     (_zz_3549[31:0]         ), //i
    .dout    (fixTo_1308_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_1309 (
    .din     (_zz_3550[31:0]         ), //i
    .dout    (fixTo_1309_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1310 (
    .din     (_zz_3551[31:0]         ), //i
    .dout    (fixTo_1310_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1311 (
    .din     (_zz_3552[31:0]         ), //i
    .dout    (fixTo_1311_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1312 (
    .din     (_zz_3553[31:0]         ), //i
    .dout    (fixTo_1312_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1313 (
    .din     (_zz_3554[31:0]         ), //i
    .dout    (fixTo_1313_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_1314 (
    .din     (_zz_3555[31:0]         ), //i
    .dout    (fixTo_1314_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_1315 (
    .din     (_zz_3556[31:0]         ), //i
    .dout    (fixTo_1315_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1316 (
    .din     (_zz_3557[31:0]         ), //i
    .dout    (fixTo_1316_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1317 (
    .din     (_zz_3558[31:0]         ), //i
    .dout    (fixTo_1317_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1318 (
    .din     (_zz_3559[31:0]         ), //i
    .dout    (fixTo_1318_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1319 (
    .din     (_zz_3560[31:0]         ), //i
    .dout    (fixTo_1319_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_1320 (
    .din     (_zz_3561[31:0]         ), //i
    .dout    (fixTo_1320_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_1321 (
    .din     (_zz_3562[31:0]         ), //i
    .dout    (fixTo_1321_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1322 (
    .din     (_zz_3563[31:0]         ), //i
    .dout    (fixTo_1322_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1323 (
    .din     (_zz_3564[31:0]         ), //i
    .dout    (fixTo_1323_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1324 (
    .din     (_zz_3565[31:0]         ), //i
    .dout    (fixTo_1324_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1325 (
    .din     (_zz_3566[31:0]         ), //i
    .dout    (fixTo_1325_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_1326 (
    .din     (_zz_3567[31:0]         ), //i
    .dout    (fixTo_1326_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_1327 (
    .din     (_zz_3568[31:0]         ), //i
    .dout    (fixTo_1327_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1328 (
    .din     (_zz_3569[31:0]         ), //i
    .dout    (fixTo_1328_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1329 (
    .din     (_zz_3570[31:0]         ), //i
    .dout    (fixTo_1329_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1330 (
    .din     (_zz_3571[31:0]         ), //i
    .dout    (fixTo_1330_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1331 (
    .din     (_zz_3572[31:0]         ), //i
    .dout    (fixTo_1331_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_1332 (
    .din     (_zz_3573[31:0]         ), //i
    .dout    (fixTo_1332_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_1333 (
    .din     (_zz_3574[31:0]         ), //i
    .dout    (fixTo_1333_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1334 (
    .din     (_zz_3575[31:0]         ), //i
    .dout    (fixTo_1334_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1335 (
    .din     (_zz_3576[31:0]         ), //i
    .dout    (fixTo_1335_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1336 (
    .din     (_zz_3577[31:0]         ), //i
    .dout    (fixTo_1336_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1337 (
    .din     (_zz_3578[31:0]         ), //i
    .dout    (fixTo_1337_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_1338 (
    .din     (_zz_3579[31:0]         ), //i
    .dout    (fixTo_1338_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_1339 (
    .din     (_zz_3580[31:0]         ), //i
    .dout    (fixTo_1339_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1340 (
    .din     (_zz_3581[31:0]         ), //i
    .dout    (fixTo_1340_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1341 (
    .din     (_zz_3582[31:0]         ), //i
    .dout    (fixTo_1341_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1342 (
    .din     (_zz_3583[31:0]         ), //i
    .dout    (fixTo_1342_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1343 (
    .din     (_zz_3584[31:0]         ), //i
    .dout    (fixTo_1343_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_1344 (
    .din     (_zz_3585[31:0]         ), //i
    .dout    (fixTo_1344_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_1345 (
    .din     (_zz_3586[31:0]         ), //i
    .dout    (fixTo_1345_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1346 (
    .din     (_zz_3587[31:0]         ), //i
    .dout    (fixTo_1346_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1347 (
    .din     (_zz_3588[31:0]         ), //i
    .dout    (fixTo_1347_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1348 (
    .din     (_zz_3589[31:0]         ), //i
    .dout    (fixTo_1348_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1349 (
    .din     (_zz_3590[31:0]         ), //i
    .dout    (fixTo_1349_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_1350 (
    .din     (_zz_3591[31:0]         ), //i
    .dout    (fixTo_1350_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_1351 (
    .din     (_zz_3592[31:0]         ), //i
    .dout    (fixTo_1351_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1352 (
    .din     (_zz_3593[31:0]         ), //i
    .dout    (fixTo_1352_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1353 (
    .din     (_zz_3594[31:0]         ), //i
    .dout    (fixTo_1353_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1354 (
    .din     (_zz_3595[31:0]         ), //i
    .dout    (fixTo_1354_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1355 (
    .din     (_zz_3596[31:0]         ), //i
    .dout    (fixTo_1355_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_1356 (
    .din     (_zz_3597[31:0]         ), //i
    .dout    (fixTo_1356_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_1357 (
    .din     (_zz_3598[31:0]         ), //i
    .dout    (fixTo_1357_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1358 (
    .din     (_zz_3599[31:0]         ), //i
    .dout    (fixTo_1358_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1359 (
    .din     (_zz_3600[31:0]         ), //i
    .dout    (fixTo_1359_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1360 (
    .din     (_zz_3601[31:0]         ), //i
    .dout    (fixTo_1360_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1361 (
    .din     (_zz_3602[31:0]         ), //i
    .dout    (fixTo_1361_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_1362 (
    .din     (_zz_3603[31:0]         ), //i
    .dout    (fixTo_1362_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_1363 (
    .din     (_zz_3604[31:0]         ), //i
    .dout    (fixTo_1363_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1364 (
    .din     (_zz_3605[31:0]         ), //i
    .dout    (fixTo_1364_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1365 (
    .din     (_zz_3606[31:0]         ), //i
    .dout    (fixTo_1365_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1366 (
    .din     (_zz_3607[31:0]         ), //i
    .dout    (fixTo_1366_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1367 (
    .din     (_zz_3608[31:0]         ), //i
    .dout    (fixTo_1367_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_1368 (
    .din     (_zz_3609[31:0]         ), //i
    .dout    (fixTo_1368_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_1369 (
    .din     (_zz_3610[31:0]         ), //i
    .dout    (fixTo_1369_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1370 (
    .din     (_zz_3611[31:0]         ), //i
    .dout    (fixTo_1370_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1371 (
    .din     (_zz_3612[31:0]         ), //i
    .dout    (fixTo_1371_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1372 (
    .din     (_zz_3613[31:0]         ), //i
    .dout    (fixTo_1372_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1373 (
    .din     (_zz_3614[31:0]         ), //i
    .dout    (fixTo_1373_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_1374 (
    .din     (_zz_3615[31:0]         ), //i
    .dout    (fixTo_1374_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_1375 (
    .din     (_zz_3616[31:0]         ), //i
    .dout    (fixTo_1375_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1376 (
    .din     (_zz_3617[31:0]         ), //i
    .dout    (fixTo_1376_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1377 (
    .din     (_zz_3618[31:0]         ), //i
    .dout    (fixTo_1377_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1378 (
    .din     (_zz_3619[31:0]         ), //i
    .dout    (fixTo_1378_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1379 (
    .din     (_zz_3620[31:0]         ), //i
    .dout    (fixTo_1379_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_1380 (
    .din     (_zz_3621[31:0]         ), //i
    .dout    (fixTo_1380_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_1381 (
    .din     (_zz_3622[31:0]         ), //i
    .dout    (fixTo_1381_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1382 (
    .din     (_zz_3623[31:0]         ), //i
    .dout    (fixTo_1382_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1383 (
    .din     (_zz_3624[31:0]         ), //i
    .dout    (fixTo_1383_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1384 (
    .din     (_zz_3625[31:0]         ), //i
    .dout    (fixTo_1384_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1385 (
    .din     (_zz_3626[31:0]         ), //i
    .dout    (fixTo_1385_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_1386 (
    .din     (_zz_3627[31:0]         ), //i
    .dout    (fixTo_1386_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_1387 (
    .din     (_zz_3628[31:0]         ), //i
    .dout    (fixTo_1387_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1388 (
    .din     (_zz_3629[31:0]         ), //i
    .dout    (fixTo_1388_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1389 (
    .din     (_zz_3630[31:0]         ), //i
    .dout    (fixTo_1389_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1390 (
    .din     (_zz_3631[31:0]         ), //i
    .dout    (fixTo_1390_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1391 (
    .din     (_zz_3632[31:0]         ), //i
    .dout    (fixTo_1391_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_1392 (
    .din     (_zz_3633[31:0]         ), //i
    .dout    (fixTo_1392_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_1393 (
    .din     (_zz_3634[31:0]         ), //i
    .dout    (fixTo_1393_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1394 (
    .din     (_zz_3635[31:0]         ), //i
    .dout    (fixTo_1394_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1395 (
    .din     (_zz_3636[31:0]         ), //i
    .dout    (fixTo_1395_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1396 (
    .din     (_zz_3637[31:0]         ), //i
    .dout    (fixTo_1396_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1397 (
    .din     (_zz_3638[31:0]         ), //i
    .dout    (fixTo_1397_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_1398 (
    .din     (_zz_3639[31:0]         ), //i
    .dout    (fixTo_1398_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_1399 (
    .din     (_zz_3640[31:0]         ), //i
    .dout    (fixTo_1399_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1400 (
    .din     (_zz_3641[31:0]         ), //i
    .dout    (fixTo_1400_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1401 (
    .din     (_zz_3642[31:0]         ), //i
    .dout    (fixTo_1401_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1402 (
    .din     (_zz_3643[31:0]         ), //i
    .dout    (fixTo_1402_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1403 (
    .din     (_zz_3644[31:0]         ), //i
    .dout    (fixTo_1403_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_1404 (
    .din     (_zz_3645[31:0]         ), //i
    .dout    (fixTo_1404_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_1405 (
    .din     (_zz_3646[31:0]         ), //i
    .dout    (fixTo_1405_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1406 (
    .din     (_zz_3647[31:0]         ), //i
    .dout    (fixTo_1406_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1407 (
    .din     (_zz_3648[31:0]         ), //i
    .dout    (fixTo_1407_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1408 (
    .din     (_zz_3649[31:0]         ), //i
    .dout    (fixTo_1408_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1409 (
    .din     (_zz_3650[31:0]         ), //i
    .dout    (fixTo_1409_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_1410 (
    .din     (_zz_3651[31:0]         ), //i
    .dout    (fixTo_1410_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_1411 (
    .din     (_zz_3652[31:0]         ), //i
    .dout    (fixTo_1411_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1412 (
    .din     (_zz_3653[31:0]         ), //i
    .dout    (fixTo_1412_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1413 (
    .din     (_zz_3654[31:0]         ), //i
    .dout    (fixTo_1413_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1414 (
    .din     (_zz_3655[31:0]         ), //i
    .dout    (fixTo_1414_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1415 (
    .din     (_zz_3656[31:0]         ), //i
    .dout    (fixTo_1415_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_1416 (
    .din     (_zz_3657[31:0]         ), //i
    .dout    (fixTo_1416_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_1417 (
    .din     (_zz_3658[31:0]         ), //i
    .dout    (fixTo_1417_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1418 (
    .din     (_zz_3659[31:0]         ), //i
    .dout    (fixTo_1418_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1419 (
    .din     (_zz_3660[31:0]         ), //i
    .dout    (fixTo_1419_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1420 (
    .din     (_zz_3661[31:0]         ), //i
    .dout    (fixTo_1420_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1421 (
    .din     (_zz_3662[31:0]         ), //i
    .dout    (fixTo_1421_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_1422 (
    .din     (_zz_3663[31:0]         ), //i
    .dout    (fixTo_1422_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_1423 (
    .din     (_zz_3664[31:0]         ), //i
    .dout    (fixTo_1423_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1424 (
    .din     (_zz_3665[31:0]         ), //i
    .dout    (fixTo_1424_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1425 (
    .din     (_zz_3666[31:0]         ), //i
    .dout    (fixTo_1425_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1426 (
    .din     (_zz_3667[31:0]         ), //i
    .dout    (fixTo_1426_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1427 (
    .din     (_zz_3668[31:0]         ), //i
    .dout    (fixTo_1427_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_1428 (
    .din     (_zz_3669[31:0]         ), //i
    .dout    (fixTo_1428_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_1429 (
    .din     (_zz_3670[31:0]         ), //i
    .dout    (fixTo_1429_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1430 (
    .din     (_zz_3671[31:0]         ), //i
    .dout    (fixTo_1430_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1431 (
    .din     (_zz_3672[31:0]         ), //i
    .dout    (fixTo_1431_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1432 (
    .din     (_zz_3673[31:0]         ), //i
    .dout    (fixTo_1432_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1433 (
    .din     (_zz_3674[31:0]         ), //i
    .dout    (fixTo_1433_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_1434 (
    .din     (_zz_3675[31:0]         ), //i
    .dout    (fixTo_1434_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_1435 (
    .din     (_zz_3676[31:0]         ), //i
    .dout    (fixTo_1435_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1436 (
    .din     (_zz_3677[31:0]         ), //i
    .dout    (fixTo_1436_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1437 (
    .din     (_zz_3678[31:0]         ), //i
    .dout    (fixTo_1437_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1438 (
    .din     (_zz_3679[31:0]         ), //i
    .dout    (fixTo_1438_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1439 (
    .din     (_zz_3680[31:0]         ), //i
    .dout    (fixTo_1439_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_1440 (
    .din     (_zz_3681[31:0]         ), //i
    .dout    (fixTo_1440_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_1441 (
    .din     (_zz_3682[31:0]         ), //i
    .dout    (fixTo_1441_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1442 (
    .din     (_zz_3683[31:0]         ), //i
    .dout    (fixTo_1442_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1443 (
    .din     (_zz_3684[31:0]         ), //i
    .dout    (fixTo_1443_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1444 (
    .din     (_zz_3685[31:0]         ), //i
    .dout    (fixTo_1444_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1445 (
    .din     (_zz_3686[31:0]         ), //i
    .dout    (fixTo_1445_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_1446 (
    .din     (_zz_3687[31:0]         ), //i
    .dout    (fixTo_1446_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_1447 (
    .din     (_zz_3688[31:0]         ), //i
    .dout    (fixTo_1447_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1448 (
    .din     (_zz_3689[31:0]         ), //i
    .dout    (fixTo_1448_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1449 (
    .din     (_zz_3690[31:0]         ), //i
    .dout    (fixTo_1449_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1450 (
    .din     (_zz_3691[31:0]         ), //i
    .dout    (fixTo_1450_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1451 (
    .din     (_zz_3692[31:0]         ), //i
    .dout    (fixTo_1451_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_1452 (
    .din     (_zz_3693[31:0]         ), //i
    .dout    (fixTo_1452_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_1453 (
    .din     (_zz_3694[31:0]         ), //i
    .dout    (fixTo_1453_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1454 (
    .din     (_zz_3695[31:0]         ), //i
    .dout    (fixTo_1454_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1455 (
    .din     (_zz_3696[31:0]         ), //i
    .dout    (fixTo_1455_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1456 (
    .din     (_zz_3697[31:0]         ), //i
    .dout    (fixTo_1456_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1457 (
    .din     (_zz_3698[31:0]         ), //i
    .dout    (fixTo_1457_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_1458 (
    .din     (_zz_3699[31:0]         ), //i
    .dout    (fixTo_1458_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_1459 (
    .din     (_zz_3700[31:0]         ), //i
    .dout    (fixTo_1459_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1460 (
    .din     (_zz_3701[31:0]         ), //i
    .dout    (fixTo_1460_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1461 (
    .din     (_zz_3702[31:0]         ), //i
    .dout    (fixTo_1461_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1462 (
    .din     (_zz_3703[31:0]         ), //i
    .dout    (fixTo_1462_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1463 (
    .din     (_zz_3704[31:0]         ), //i
    .dout    (fixTo_1463_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_1464 (
    .din     (_zz_3705[31:0]         ), //i
    .dout    (fixTo_1464_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_1465 (
    .din     (_zz_3706[31:0]         ), //i
    .dout    (fixTo_1465_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1466 (
    .din     (_zz_3707[31:0]         ), //i
    .dout    (fixTo_1466_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1467 (
    .din     (_zz_3708[31:0]         ), //i
    .dout    (fixTo_1467_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1468 (
    .din     (_zz_3709[31:0]         ), //i
    .dout    (fixTo_1468_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1469 (
    .din     (_zz_3710[31:0]         ), //i
    .dout    (fixTo_1469_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_1470 (
    .din     (_zz_3711[31:0]         ), //i
    .dout    (fixTo_1470_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_1471 (
    .din     (_zz_3712[31:0]         ), //i
    .dout    (fixTo_1471_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1472 (
    .din     (_zz_3713[31:0]         ), //i
    .dout    (fixTo_1472_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1473 (
    .din     (_zz_3714[31:0]         ), //i
    .dout    (fixTo_1473_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1474 (
    .din     (_zz_3715[31:0]         ), //i
    .dout    (fixTo_1474_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1475 (
    .din     (_zz_3716[31:0]         ), //i
    .dout    (fixTo_1475_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_1476 (
    .din     (_zz_3717[31:0]         ), //i
    .dout    (fixTo_1476_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_1477 (
    .din     (_zz_3718[31:0]         ), //i
    .dout    (fixTo_1477_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1478 (
    .din     (_zz_3719[31:0]         ), //i
    .dout    (fixTo_1478_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1479 (
    .din     (_zz_3720[31:0]         ), //i
    .dout    (fixTo_1479_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1480 (
    .din     (_zz_3721[31:0]         ), //i
    .dout    (fixTo_1480_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1481 (
    .din     (_zz_3722[31:0]         ), //i
    .dout    (fixTo_1481_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_1482 (
    .din     (_zz_3723[31:0]         ), //i
    .dout    (fixTo_1482_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_1483 (
    .din     (_zz_3724[31:0]         ), //i
    .dout    (fixTo_1483_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1484 (
    .din     (_zz_3725[31:0]         ), //i
    .dout    (fixTo_1484_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1485 (
    .din     (_zz_3726[31:0]         ), //i
    .dout    (fixTo_1485_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1486 (
    .din     (_zz_3727[31:0]         ), //i
    .dout    (fixTo_1486_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1487 (
    .din     (_zz_3728[31:0]         ), //i
    .dout    (fixTo_1487_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_1488 (
    .din     (_zz_3729[31:0]         ), //i
    .dout    (fixTo_1488_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_1489 (
    .din     (_zz_3730[31:0]         ), //i
    .dout    (fixTo_1489_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1490 (
    .din     (_zz_3731[31:0]         ), //i
    .dout    (fixTo_1490_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1491 (
    .din     (_zz_3732[31:0]         ), //i
    .dout    (fixTo_1491_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1492 (
    .din     (_zz_3733[31:0]         ), //i
    .dout    (fixTo_1492_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1493 (
    .din     (_zz_3734[31:0]         ), //i
    .dout    (fixTo_1493_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_1494 (
    .din     (_zz_3735[31:0]         ), //i
    .dout    (fixTo_1494_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_1495 (
    .din     (_zz_3736[31:0]         ), //i
    .dout    (fixTo_1495_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1496 (
    .din     (_zz_3737[31:0]         ), //i
    .dout    (fixTo_1496_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1497 (
    .din     (_zz_3738[31:0]         ), //i
    .dout    (fixTo_1497_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1498 (
    .din     (_zz_3739[31:0]         ), //i
    .dout    (fixTo_1498_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1499 (
    .din     (_zz_3740[31:0]         ), //i
    .dout    (fixTo_1499_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_1500 (
    .din     (_zz_3741[31:0]         ), //i
    .dout    (fixTo_1500_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_1501 (
    .din     (_zz_3742[31:0]         ), //i
    .dout    (fixTo_1501_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1502 (
    .din     (_zz_3743[31:0]         ), //i
    .dout    (fixTo_1502_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1503 (
    .din     (_zz_3744[31:0]         ), //i
    .dout    (fixTo_1503_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1504 (
    .din     (_zz_3745[31:0]         ), //i
    .dout    (fixTo_1504_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1505 (
    .din     (_zz_3746[31:0]         ), //i
    .dout    (fixTo_1505_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_1506 (
    .din     (_zz_3747[31:0]         ), //i
    .dout    (fixTo_1506_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_1507 (
    .din     (_zz_3748[31:0]         ), //i
    .dout    (fixTo_1507_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1508 (
    .din     (_zz_3749[31:0]         ), //i
    .dout    (fixTo_1508_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1509 (
    .din     (_zz_3750[31:0]         ), //i
    .dout    (fixTo_1509_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1510 (
    .din     (_zz_3751[31:0]         ), //i
    .dout    (fixTo_1510_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1511 (
    .din     (_zz_3752[31:0]         ), //i
    .dout    (fixTo_1511_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_1512 (
    .din     (_zz_3753[31:0]         ), //i
    .dout    (fixTo_1512_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_1513 (
    .din     (_zz_3754[31:0]         ), //i
    .dout    (fixTo_1513_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1514 (
    .din     (_zz_3755[31:0]         ), //i
    .dout    (fixTo_1514_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1515 (
    .din     (_zz_3756[31:0]         ), //i
    .dout    (fixTo_1515_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1516 (
    .din     (_zz_3757[31:0]         ), //i
    .dout    (fixTo_1516_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1517 (
    .din     (_zz_3758[31:0]         ), //i
    .dout    (fixTo_1517_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_1518 (
    .din     (_zz_3759[31:0]         ), //i
    .dout    (fixTo_1518_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_1519 (
    .din     (_zz_3760[31:0]         ), //i
    .dout    (fixTo_1519_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1520 (
    .din     (_zz_3761[31:0]         ), //i
    .dout    (fixTo_1520_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1521 (
    .din     (_zz_3762[31:0]         ), //i
    .dout    (fixTo_1521_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1522 (
    .din     (_zz_3763[31:0]         ), //i
    .dout    (fixTo_1522_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1523 (
    .din     (_zz_3764[31:0]         ), //i
    .dout    (fixTo_1523_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_1524 (
    .din     (_zz_3765[31:0]         ), //i
    .dout    (fixTo_1524_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_1525 (
    .din     (_zz_3766[31:0]         ), //i
    .dout    (fixTo_1525_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1526 (
    .din     (_zz_3767[31:0]         ), //i
    .dout    (fixTo_1526_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1527 (
    .din     (_zz_3768[31:0]         ), //i
    .dout    (fixTo_1527_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1528 (
    .din     (_zz_3769[31:0]         ), //i
    .dout    (fixTo_1528_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1529 (
    .din     (_zz_3770[31:0]         ), //i
    .dout    (fixTo_1529_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_1530 (
    .din     (_zz_3771[31:0]         ), //i
    .dout    (fixTo_1530_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_1531 (
    .din     (_zz_3772[31:0]         ), //i
    .dout    (fixTo_1531_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1532 (
    .din     (_zz_3773[31:0]         ), //i
    .dout    (fixTo_1532_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1533 (
    .din     (_zz_3774[31:0]         ), //i
    .dout    (fixTo_1533_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1534 (
    .din     (_zz_3775[31:0]         ), //i
    .dout    (fixTo_1534_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1535 (
    .din     (_zz_3776[31:0]         ), //i
    .dout    (fixTo_1535_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_1536 (
    .din     (_zz_3777[31:0]         ), //i
    .dout    (fixTo_1536_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_1537 (
    .din     (_zz_3778[31:0]         ), //i
    .dout    (fixTo_1537_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1538 (
    .din     (_zz_3779[31:0]         ), //i
    .dout    (fixTo_1538_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1539 (
    .din     (_zz_3780[31:0]         ), //i
    .dout    (fixTo_1539_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1540 (
    .din     (_zz_3781[31:0]         ), //i
    .dout    (fixTo_1540_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1541 (
    .din     (_zz_3782[31:0]         ), //i
    .dout    (fixTo_1541_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_1542 (
    .din     (_zz_3783[31:0]         ), //i
    .dout    (fixTo_1542_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_1543 (
    .din     (_zz_3784[31:0]         ), //i
    .dout    (fixTo_1543_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1544 (
    .din     (_zz_3785[31:0]         ), //i
    .dout    (fixTo_1544_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1545 (
    .din     (_zz_3786[31:0]         ), //i
    .dout    (fixTo_1545_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1546 (
    .din     (_zz_3787[31:0]         ), //i
    .dout    (fixTo_1546_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1547 (
    .din     (_zz_3788[31:0]         ), //i
    .dout    (fixTo_1547_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_1548 (
    .din     (_zz_3789[31:0]         ), //i
    .dout    (fixTo_1548_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_1549 (
    .din     (_zz_3790[31:0]         ), //i
    .dout    (fixTo_1549_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1550 (
    .din     (_zz_3791[31:0]         ), //i
    .dout    (fixTo_1550_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1551 (
    .din     (_zz_3792[31:0]         ), //i
    .dout    (fixTo_1551_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1552 (
    .din     (_zz_3793[31:0]         ), //i
    .dout    (fixTo_1552_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1553 (
    .din     (_zz_3794[31:0]         ), //i
    .dout    (fixTo_1553_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_1554 (
    .din     (_zz_3795[31:0]         ), //i
    .dout    (fixTo_1554_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_1555 (
    .din     (_zz_3796[31:0]         ), //i
    .dout    (fixTo_1555_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1556 (
    .din     (_zz_3797[31:0]         ), //i
    .dout    (fixTo_1556_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1557 (
    .din     (_zz_3798[31:0]         ), //i
    .dout    (fixTo_1557_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1558 (
    .din     (_zz_3799[31:0]         ), //i
    .dout    (fixTo_1558_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1559 (
    .din     (_zz_3800[31:0]         ), //i
    .dout    (fixTo_1559_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_1560 (
    .din     (_zz_3801[31:0]         ), //i
    .dout    (fixTo_1560_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_1561 (
    .din     (_zz_3802[31:0]         ), //i
    .dout    (fixTo_1561_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1562 (
    .din     (_zz_3803[31:0]         ), //i
    .dout    (fixTo_1562_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1563 (
    .din     (_zz_3804[31:0]         ), //i
    .dout    (fixTo_1563_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1564 (
    .din     (_zz_3805[31:0]         ), //i
    .dout    (fixTo_1564_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1565 (
    .din     (_zz_3806[31:0]         ), //i
    .dout    (fixTo_1565_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_1566 (
    .din     (_zz_3807[31:0]         ), //i
    .dout    (fixTo_1566_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_1567 (
    .din     (_zz_3808[31:0]         ), //i
    .dout    (fixTo_1567_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1568 (
    .din     (_zz_3809[31:0]         ), //i
    .dout    (fixTo_1568_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1569 (
    .din     (_zz_3810[31:0]         ), //i
    .dout    (fixTo_1569_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1570 (
    .din     (_zz_3811[31:0]         ), //i
    .dout    (fixTo_1570_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1571 (
    .din     (_zz_3812[31:0]         ), //i
    .dout    (fixTo_1571_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_1572 (
    .din     (_zz_3813[31:0]         ), //i
    .dout    (fixTo_1572_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_1573 (
    .din     (_zz_3814[31:0]         ), //i
    .dout    (fixTo_1573_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1574 (
    .din     (_zz_3815[31:0]         ), //i
    .dout    (fixTo_1574_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1575 (
    .din     (_zz_3816[31:0]         ), //i
    .dout    (fixTo_1575_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1576 (
    .din     (_zz_3817[31:0]         ), //i
    .dout    (fixTo_1576_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1577 (
    .din     (_zz_3818[31:0]         ), //i
    .dout    (fixTo_1577_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_1578 (
    .din     (_zz_3819[31:0]         ), //i
    .dout    (fixTo_1578_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_1579 (
    .din     (_zz_3820[31:0]         ), //i
    .dout    (fixTo_1579_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1580 (
    .din     (_zz_3821[31:0]         ), //i
    .dout    (fixTo_1580_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1581 (
    .din     (_zz_3822[31:0]         ), //i
    .dout    (fixTo_1581_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1582 (
    .din     (_zz_3823[31:0]         ), //i
    .dout    (fixTo_1582_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1583 (
    .din     (_zz_3824[31:0]         ), //i
    .dout    (fixTo_1583_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_1584 (
    .din     (_zz_3825[31:0]         ), //i
    .dout    (fixTo_1584_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_1585 (
    .din     (_zz_3826[31:0]         ), //i
    .dout    (fixTo_1585_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1586 (
    .din     (_zz_3827[31:0]         ), //i
    .dout    (fixTo_1586_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1587 (
    .din     (_zz_3828[31:0]         ), //i
    .dout    (fixTo_1587_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1588 (
    .din     (_zz_3829[31:0]         ), //i
    .dout    (fixTo_1588_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1589 (
    .din     (_zz_3830[31:0]         ), //i
    .dout    (fixTo_1589_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_1590 (
    .din     (_zz_3831[31:0]         ), //i
    .dout    (fixTo_1590_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_1591 (
    .din     (_zz_3832[31:0]         ), //i
    .dout    (fixTo_1591_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1592 (
    .din     (_zz_3833[31:0]         ), //i
    .dout    (fixTo_1592_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1593 (
    .din     (_zz_3834[31:0]         ), //i
    .dout    (fixTo_1593_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1594 (
    .din     (_zz_3835[31:0]         ), //i
    .dout    (fixTo_1594_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1595 (
    .din     (_zz_3836[31:0]         ), //i
    .dout    (fixTo_1595_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_1596 (
    .din     (_zz_3837[31:0]         ), //i
    .dout    (fixTo_1596_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_1597 (
    .din     (_zz_3838[31:0]         ), //i
    .dout    (fixTo_1597_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1598 (
    .din     (_zz_3839[31:0]         ), //i
    .dout    (fixTo_1598_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1599 (
    .din     (_zz_3840[31:0]         ), //i
    .dout    (fixTo_1599_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1600 (
    .din     (_zz_3841[31:0]         ), //i
    .dout    (fixTo_1600_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1601 (
    .din     (_zz_3842[31:0]         ), //i
    .dout    (fixTo_1601_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_1602 (
    .din     (_zz_3843[31:0]         ), //i
    .dout    (fixTo_1602_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_1603 (
    .din     (_zz_3844[31:0]         ), //i
    .dout    (fixTo_1603_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1604 (
    .din     (_zz_3845[31:0]         ), //i
    .dout    (fixTo_1604_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1605 (
    .din     (_zz_3846[31:0]         ), //i
    .dout    (fixTo_1605_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1606 (
    .din     (_zz_3847[31:0]         ), //i
    .dout    (fixTo_1606_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1607 (
    .din     (_zz_3848[31:0]         ), //i
    .dout    (fixTo_1607_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_1608 (
    .din     (_zz_3849[31:0]         ), //i
    .dout    (fixTo_1608_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_1609 (
    .din     (_zz_3850[31:0]         ), //i
    .dout    (fixTo_1609_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1610 (
    .din     (_zz_3851[31:0]         ), //i
    .dout    (fixTo_1610_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1611 (
    .din     (_zz_3852[31:0]         ), //i
    .dout    (fixTo_1611_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1612 (
    .din     (_zz_3853[31:0]         ), //i
    .dout    (fixTo_1612_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1613 (
    .din     (_zz_3854[31:0]         ), //i
    .dout    (fixTo_1613_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_1614 (
    .din     (_zz_3855[31:0]         ), //i
    .dout    (fixTo_1614_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_1615 (
    .din     (_zz_3856[31:0]         ), //i
    .dout    (fixTo_1615_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1616 (
    .din     (_zz_3857[31:0]         ), //i
    .dout    (fixTo_1616_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1617 (
    .din     (_zz_3858[31:0]         ), //i
    .dout    (fixTo_1617_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1618 (
    .din     (_zz_3859[31:0]         ), //i
    .dout    (fixTo_1618_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1619 (
    .din     (_zz_3860[31:0]         ), //i
    .dout    (fixTo_1619_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_1620 (
    .din     (_zz_3861[31:0]         ), //i
    .dout    (fixTo_1620_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_1621 (
    .din     (_zz_3862[31:0]         ), //i
    .dout    (fixTo_1621_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1622 (
    .din     (_zz_3863[31:0]         ), //i
    .dout    (fixTo_1622_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1623 (
    .din     (_zz_3864[31:0]         ), //i
    .dout    (fixTo_1623_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1624 (
    .din     (_zz_3865[31:0]         ), //i
    .dout    (fixTo_1624_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1625 (
    .din     (_zz_3866[31:0]         ), //i
    .dout    (fixTo_1625_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_1626 (
    .din     (_zz_3867[31:0]         ), //i
    .dout    (fixTo_1626_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_1627 (
    .din     (_zz_3868[31:0]         ), //i
    .dout    (fixTo_1627_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1628 (
    .din     (_zz_3869[31:0]         ), //i
    .dout    (fixTo_1628_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1629 (
    .din     (_zz_3870[31:0]         ), //i
    .dout    (fixTo_1629_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1630 (
    .din     (_zz_3871[31:0]         ), //i
    .dout    (fixTo_1630_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1631 (
    .din     (_zz_3872[31:0]         ), //i
    .dout    (fixTo_1631_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_1632 (
    .din     (_zz_3873[31:0]         ), //i
    .dout    (fixTo_1632_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_1633 (
    .din     (_zz_3874[31:0]         ), //i
    .dout    (fixTo_1633_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1634 (
    .din     (_zz_3875[31:0]         ), //i
    .dout    (fixTo_1634_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1635 (
    .din     (_zz_3876[31:0]         ), //i
    .dout    (fixTo_1635_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1636 (
    .din     (_zz_3877[31:0]         ), //i
    .dout    (fixTo_1636_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1637 (
    .din     (_zz_3878[31:0]         ), //i
    .dout    (fixTo_1637_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_1638 (
    .din     (_zz_3879[31:0]         ), //i
    .dout    (fixTo_1638_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_1639 (
    .din     (_zz_3880[31:0]         ), //i
    .dout    (fixTo_1639_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1640 (
    .din     (_zz_3881[31:0]         ), //i
    .dout    (fixTo_1640_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1641 (
    .din     (_zz_3882[31:0]         ), //i
    .dout    (fixTo_1641_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1642 (
    .din     (_zz_3883[31:0]         ), //i
    .dout    (fixTo_1642_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1643 (
    .din     (_zz_3884[31:0]         ), //i
    .dout    (fixTo_1643_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_1644 (
    .din     (_zz_3885[31:0]         ), //i
    .dout    (fixTo_1644_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_1645 (
    .din     (_zz_3886[31:0]         ), //i
    .dout    (fixTo_1645_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1646 (
    .din     (_zz_3887[31:0]         ), //i
    .dout    (fixTo_1646_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1647 (
    .din     (_zz_3888[31:0]         ), //i
    .dout    (fixTo_1647_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1648 (
    .din     (_zz_3889[31:0]         ), //i
    .dout    (fixTo_1648_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1649 (
    .din     (_zz_3890[31:0]         ), //i
    .dout    (fixTo_1649_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_1650 (
    .din     (_zz_3891[31:0]         ), //i
    .dout    (fixTo_1650_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_1651 (
    .din     (_zz_3892[31:0]         ), //i
    .dout    (fixTo_1651_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1652 (
    .din     (_zz_3893[31:0]         ), //i
    .dout    (fixTo_1652_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1653 (
    .din     (_zz_3894[31:0]         ), //i
    .dout    (fixTo_1653_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1654 (
    .din     (_zz_3895[31:0]         ), //i
    .dout    (fixTo_1654_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1655 (
    .din     (_zz_3896[31:0]         ), //i
    .dout    (fixTo_1655_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_1656 (
    .din     (_zz_3897[31:0]         ), //i
    .dout    (fixTo_1656_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_1657 (
    .din     (_zz_3898[31:0]         ), //i
    .dout    (fixTo_1657_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1658 (
    .din     (_zz_3899[31:0]         ), //i
    .dout    (fixTo_1658_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1659 (
    .din     (_zz_3900[31:0]         ), //i
    .dout    (fixTo_1659_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1660 (
    .din     (_zz_3901[31:0]         ), //i
    .dout    (fixTo_1660_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1661 (
    .din     (_zz_3902[31:0]         ), //i
    .dout    (fixTo_1661_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_1662 (
    .din     (_zz_3903[31:0]         ), //i
    .dout    (fixTo_1662_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_1663 (
    .din     (_zz_3904[31:0]         ), //i
    .dout    (fixTo_1663_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1664 (
    .din     (_zz_3905[31:0]         ), //i
    .dout    (fixTo_1664_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1665 (
    .din     (_zz_3906[31:0]         ), //i
    .dout    (fixTo_1665_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1666 (
    .din     (_zz_3907[31:0]         ), //i
    .dout    (fixTo_1666_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1667 (
    .din     (_zz_3908[31:0]         ), //i
    .dout    (fixTo_1667_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_1668 (
    .din     (_zz_3909[31:0]         ), //i
    .dout    (fixTo_1668_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_1669 (
    .din     (_zz_3910[31:0]         ), //i
    .dout    (fixTo_1669_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1670 (
    .din     (_zz_3911[31:0]         ), //i
    .dout    (fixTo_1670_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1671 (
    .din     (_zz_3912[31:0]         ), //i
    .dout    (fixTo_1671_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1672 (
    .din     (_zz_3913[31:0]         ), //i
    .dout    (fixTo_1672_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1673 (
    .din     (_zz_3914[31:0]         ), //i
    .dout    (fixTo_1673_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_1674 (
    .din     (_zz_3915[31:0]         ), //i
    .dout    (fixTo_1674_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_1675 (
    .din     (_zz_3916[31:0]         ), //i
    .dout    (fixTo_1675_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1676 (
    .din     (_zz_3917[31:0]         ), //i
    .dout    (fixTo_1676_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1677 (
    .din     (_zz_3918[31:0]         ), //i
    .dout    (fixTo_1677_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1678 (
    .din     (_zz_3919[31:0]         ), //i
    .dout    (fixTo_1678_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1679 (
    .din     (_zz_3920[31:0]         ), //i
    .dout    (fixTo_1679_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_1680 (
    .din     (_zz_3921[31:0]         ), //i
    .dout    (fixTo_1680_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_1681 (
    .din     (_zz_3922[31:0]         ), //i
    .dout    (fixTo_1681_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1682 (
    .din     (_zz_3923[31:0]         ), //i
    .dout    (fixTo_1682_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1683 (
    .din     (_zz_3924[31:0]         ), //i
    .dout    (fixTo_1683_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1684 (
    .din     (_zz_3925[31:0]         ), //i
    .dout    (fixTo_1684_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1685 (
    .din     (_zz_3926[31:0]         ), //i
    .dout    (fixTo_1685_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_1686 (
    .din     (_zz_3927[31:0]         ), //i
    .dout    (fixTo_1686_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_1687 (
    .din     (_zz_3928[31:0]         ), //i
    .dout    (fixTo_1687_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1688 (
    .din     (_zz_3929[31:0]         ), //i
    .dout    (fixTo_1688_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1689 (
    .din     (_zz_3930[31:0]         ), //i
    .dout    (fixTo_1689_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1690 (
    .din     (_zz_3931[31:0]         ), //i
    .dout    (fixTo_1690_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1691 (
    .din     (_zz_3932[31:0]         ), //i
    .dout    (fixTo_1691_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_1692 (
    .din     (_zz_3933[31:0]         ), //i
    .dout    (fixTo_1692_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_1693 (
    .din     (_zz_3934[31:0]         ), //i
    .dout    (fixTo_1693_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1694 (
    .din     (_zz_3935[31:0]         ), //i
    .dout    (fixTo_1694_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1695 (
    .din     (_zz_3936[31:0]         ), //i
    .dout    (fixTo_1695_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1696 (
    .din     (_zz_3937[31:0]         ), //i
    .dout    (fixTo_1696_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1697 (
    .din     (_zz_3938[31:0]         ), //i
    .dout    (fixTo_1697_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_1698 (
    .din     (_zz_3939[31:0]         ), //i
    .dout    (fixTo_1698_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_1699 (
    .din     (_zz_3940[31:0]         ), //i
    .dout    (fixTo_1699_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1700 (
    .din     (_zz_3941[31:0]         ), //i
    .dout    (fixTo_1700_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1701 (
    .din     (_zz_3942[31:0]         ), //i
    .dout    (fixTo_1701_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1702 (
    .din     (_zz_3943[31:0]         ), //i
    .dout    (fixTo_1702_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1703 (
    .din     (_zz_3944[31:0]         ), //i
    .dout    (fixTo_1703_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_1704 (
    .din     (_zz_3945[31:0]         ), //i
    .dout    (fixTo_1704_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_1705 (
    .din     (_zz_3946[31:0]         ), //i
    .dout    (fixTo_1705_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1706 (
    .din     (_zz_3947[31:0]         ), //i
    .dout    (fixTo_1706_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1707 (
    .din     (_zz_3948[31:0]         ), //i
    .dout    (fixTo_1707_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1708 (
    .din     (_zz_3949[31:0]         ), //i
    .dout    (fixTo_1708_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1709 (
    .din     (_zz_3950[31:0]         ), //i
    .dout    (fixTo_1709_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_1710 (
    .din     (_zz_3951[31:0]         ), //i
    .dout    (fixTo_1710_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_1711 (
    .din     (_zz_3952[31:0]         ), //i
    .dout    (fixTo_1711_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1712 (
    .din     (_zz_3953[31:0]         ), //i
    .dout    (fixTo_1712_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1713 (
    .din     (_zz_3954[31:0]         ), //i
    .dout    (fixTo_1713_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1714 (
    .din     (_zz_3955[31:0]         ), //i
    .dout    (fixTo_1714_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1715 (
    .din     (_zz_3956[31:0]         ), //i
    .dout    (fixTo_1715_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_1716 (
    .din     (_zz_3957[31:0]         ), //i
    .dout    (fixTo_1716_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_1717 (
    .din     (_zz_3958[31:0]         ), //i
    .dout    (fixTo_1717_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1718 (
    .din     (_zz_3959[31:0]         ), //i
    .dout    (fixTo_1718_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1719 (
    .din     (_zz_3960[31:0]         ), //i
    .dout    (fixTo_1719_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1720 (
    .din     (_zz_3961[31:0]         ), //i
    .dout    (fixTo_1720_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1721 (
    .din     (_zz_3962[31:0]         ), //i
    .dout    (fixTo_1721_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_1722 (
    .din     (_zz_3963[31:0]         ), //i
    .dout    (fixTo_1722_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_1723 (
    .din     (_zz_3964[31:0]         ), //i
    .dout    (fixTo_1723_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1724 (
    .din     (_zz_3965[31:0]         ), //i
    .dout    (fixTo_1724_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1725 (
    .din     (_zz_3966[31:0]         ), //i
    .dout    (fixTo_1725_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1726 (
    .din     (_zz_3967[31:0]         ), //i
    .dout    (fixTo_1726_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1727 (
    .din     (_zz_3968[31:0]         ), //i
    .dout    (fixTo_1727_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_1728 (
    .din     (_zz_3969[31:0]         ), //i
    .dout    (fixTo_1728_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_1729 (
    .din     (_zz_3970[31:0]         ), //i
    .dout    (fixTo_1729_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1730 (
    .din     (_zz_3971[31:0]         ), //i
    .dout    (fixTo_1730_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1731 (
    .din     (_zz_3972[31:0]         ), //i
    .dout    (fixTo_1731_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1732 (
    .din     (_zz_3973[31:0]         ), //i
    .dout    (fixTo_1732_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1733 (
    .din     (_zz_3974[31:0]         ), //i
    .dout    (fixTo_1733_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_1734 (
    .din     (_zz_3975[31:0]         ), //i
    .dout    (fixTo_1734_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_1735 (
    .din     (_zz_3976[31:0]         ), //i
    .dout    (fixTo_1735_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1736 (
    .din     (_zz_3977[31:0]         ), //i
    .dout    (fixTo_1736_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1737 (
    .din     (_zz_3978[31:0]         ), //i
    .dout    (fixTo_1737_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1738 (
    .din     (_zz_3979[31:0]         ), //i
    .dout    (fixTo_1738_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1739 (
    .din     (_zz_3980[31:0]         ), //i
    .dout    (fixTo_1739_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_1740 (
    .din     (_zz_3981[31:0]         ), //i
    .dout    (fixTo_1740_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_1741 (
    .din     (_zz_3982[31:0]         ), //i
    .dout    (fixTo_1741_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1742 (
    .din     (_zz_3983[31:0]         ), //i
    .dout    (fixTo_1742_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1743 (
    .din     (_zz_3984[31:0]         ), //i
    .dout    (fixTo_1743_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1744 (
    .din     (_zz_3985[31:0]         ), //i
    .dout    (fixTo_1744_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1745 (
    .din     (_zz_3986[31:0]         ), //i
    .dout    (fixTo_1745_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_1746 (
    .din     (_zz_3987[31:0]         ), //i
    .dout    (fixTo_1746_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_1747 (
    .din     (_zz_3988[31:0]         ), //i
    .dout    (fixTo_1747_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1748 (
    .din     (_zz_3989[31:0]         ), //i
    .dout    (fixTo_1748_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1749 (
    .din     (_zz_3990[31:0]         ), //i
    .dout    (fixTo_1749_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1750 (
    .din     (_zz_3991[31:0]         ), //i
    .dout    (fixTo_1750_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1751 (
    .din     (_zz_3992[31:0]         ), //i
    .dout    (fixTo_1751_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_1752 (
    .din     (_zz_3993[31:0]         ), //i
    .dout    (fixTo_1752_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_1753 (
    .din     (_zz_3994[31:0]         ), //i
    .dout    (fixTo_1753_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1754 (
    .din     (_zz_3995[31:0]         ), //i
    .dout    (fixTo_1754_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1755 (
    .din     (_zz_3996[31:0]         ), //i
    .dout    (fixTo_1755_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1756 (
    .din     (_zz_3997[31:0]         ), //i
    .dout    (fixTo_1756_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1757 (
    .din     (_zz_3998[31:0]         ), //i
    .dout    (fixTo_1757_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_1758 (
    .din     (_zz_3999[31:0]         ), //i
    .dout    (fixTo_1758_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_1759 (
    .din     (_zz_4000[31:0]         ), //i
    .dout    (fixTo_1759_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1760 (
    .din     (_zz_4001[31:0]         ), //i
    .dout    (fixTo_1760_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1761 (
    .din     (_zz_4002[31:0]         ), //i
    .dout    (fixTo_1761_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1762 (
    .din     (_zz_4003[31:0]         ), //i
    .dout    (fixTo_1762_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1763 (
    .din     (_zz_4004[31:0]         ), //i
    .dout    (fixTo_1763_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_1764 (
    .din     (_zz_4005[31:0]         ), //i
    .dout    (fixTo_1764_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_1765 (
    .din     (_zz_4006[31:0]         ), //i
    .dout    (fixTo_1765_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1766 (
    .din     (_zz_4007[31:0]         ), //i
    .dout    (fixTo_1766_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1767 (
    .din     (_zz_4008[31:0]         ), //i
    .dout    (fixTo_1767_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1768 (
    .din     (_zz_4009[31:0]         ), //i
    .dout    (fixTo_1768_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1769 (
    .din     (_zz_4010[31:0]         ), //i
    .dout    (fixTo_1769_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_1770 (
    .din     (_zz_4011[31:0]         ), //i
    .dout    (fixTo_1770_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_1771 (
    .din     (_zz_4012[31:0]         ), //i
    .dout    (fixTo_1771_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1772 (
    .din     (_zz_4013[31:0]         ), //i
    .dout    (fixTo_1772_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1773 (
    .din     (_zz_4014[31:0]         ), //i
    .dout    (fixTo_1773_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1774 (
    .din     (_zz_4015[31:0]         ), //i
    .dout    (fixTo_1774_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1775 (
    .din     (_zz_4016[31:0]         ), //i
    .dout    (fixTo_1775_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_1776 (
    .din     (_zz_4017[31:0]         ), //i
    .dout    (fixTo_1776_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_1777 (
    .din     (_zz_4018[31:0]         ), //i
    .dout    (fixTo_1777_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1778 (
    .din     (_zz_4019[31:0]         ), //i
    .dout    (fixTo_1778_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1779 (
    .din     (_zz_4020[31:0]         ), //i
    .dout    (fixTo_1779_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1780 (
    .din     (_zz_4021[31:0]         ), //i
    .dout    (fixTo_1780_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1781 (
    .din     (_zz_4022[31:0]         ), //i
    .dout    (fixTo_1781_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_1782 (
    .din     (_zz_4023[31:0]         ), //i
    .dout    (fixTo_1782_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_1783 (
    .din     (_zz_4024[31:0]         ), //i
    .dout    (fixTo_1783_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1784 (
    .din     (_zz_4025[31:0]         ), //i
    .dout    (fixTo_1784_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1785 (
    .din     (_zz_4026[31:0]         ), //i
    .dout    (fixTo_1785_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1786 (
    .din     (_zz_4027[31:0]         ), //i
    .dout    (fixTo_1786_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1787 (
    .din     (_zz_4028[31:0]         ), //i
    .dout    (fixTo_1787_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_1788 (
    .din     (_zz_4029[31:0]         ), //i
    .dout    (fixTo_1788_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_1789 (
    .din     (_zz_4030[31:0]         ), //i
    .dout    (fixTo_1789_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1790 (
    .din     (_zz_4031[31:0]         ), //i
    .dout    (fixTo_1790_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1791 (
    .din     (_zz_4032[31:0]         ), //i
    .dout    (fixTo_1791_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1792 (
    .din     (_zz_4033[31:0]         ), //i
    .dout    (fixTo_1792_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1793 (
    .din     (_zz_4034[31:0]         ), //i
    .dout    (fixTo_1793_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_1794 (
    .din     (_zz_4035[31:0]         ), //i
    .dout    (fixTo_1794_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_1795 (
    .din     (_zz_4036[31:0]         ), //i
    .dout    (fixTo_1795_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1796 (
    .din     (_zz_4037[31:0]         ), //i
    .dout    (fixTo_1796_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1797 (
    .din     (_zz_4038[31:0]         ), //i
    .dout    (fixTo_1797_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1798 (
    .din     (_zz_4039[31:0]         ), //i
    .dout    (fixTo_1798_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1799 (
    .din     (_zz_4040[31:0]         ), //i
    .dout    (fixTo_1799_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_1800 (
    .din     (_zz_4041[31:0]         ), //i
    .dout    (fixTo_1800_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_1801 (
    .din     (_zz_4042[31:0]         ), //i
    .dout    (fixTo_1801_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1802 (
    .din     (_zz_4043[31:0]         ), //i
    .dout    (fixTo_1802_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1803 (
    .din     (_zz_4044[31:0]         ), //i
    .dout    (fixTo_1803_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1804 (
    .din     (_zz_4045[31:0]         ), //i
    .dout    (fixTo_1804_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1805 (
    .din     (_zz_4046[31:0]         ), //i
    .dout    (fixTo_1805_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_1806 (
    .din     (_zz_4047[31:0]         ), //i
    .dout    (fixTo_1806_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_1807 (
    .din     (_zz_4048[31:0]         ), //i
    .dout    (fixTo_1807_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1808 (
    .din     (_zz_4049[31:0]         ), //i
    .dout    (fixTo_1808_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1809 (
    .din     (_zz_4050[31:0]         ), //i
    .dout    (fixTo_1809_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1810 (
    .din     (_zz_4051[31:0]         ), //i
    .dout    (fixTo_1810_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1811 (
    .din     (_zz_4052[31:0]         ), //i
    .dout    (fixTo_1811_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_1812 (
    .din     (_zz_4053[31:0]         ), //i
    .dout    (fixTo_1812_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_1813 (
    .din     (_zz_4054[31:0]         ), //i
    .dout    (fixTo_1813_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1814 (
    .din     (_zz_4055[31:0]         ), //i
    .dout    (fixTo_1814_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1815 (
    .din     (_zz_4056[31:0]         ), //i
    .dout    (fixTo_1815_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1816 (
    .din     (_zz_4057[31:0]         ), //i
    .dout    (fixTo_1816_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1817 (
    .din     (_zz_4058[31:0]         ), //i
    .dout    (fixTo_1817_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_1818 (
    .din     (_zz_4059[31:0]         ), //i
    .dout    (fixTo_1818_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_1819 (
    .din     (_zz_4060[31:0]         ), //i
    .dout    (fixTo_1819_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1820 (
    .din     (_zz_4061[31:0]         ), //i
    .dout    (fixTo_1820_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1821 (
    .din     (_zz_4062[31:0]         ), //i
    .dout    (fixTo_1821_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1822 (
    .din     (_zz_4063[31:0]         ), //i
    .dout    (fixTo_1822_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1823 (
    .din     (_zz_4064[31:0]         ), //i
    .dout    (fixTo_1823_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_1824 (
    .din     (_zz_4065[31:0]         ), //i
    .dout    (fixTo_1824_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_1825 (
    .din     (_zz_4066[31:0]         ), //i
    .dout    (fixTo_1825_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1826 (
    .din     (_zz_4067[31:0]         ), //i
    .dout    (fixTo_1826_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1827 (
    .din     (_zz_4068[31:0]         ), //i
    .dout    (fixTo_1827_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1828 (
    .din     (_zz_4069[31:0]         ), //i
    .dout    (fixTo_1828_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1829 (
    .din     (_zz_4070[31:0]         ), //i
    .dout    (fixTo_1829_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_1830 (
    .din     (_zz_4071[31:0]         ), //i
    .dout    (fixTo_1830_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_1831 (
    .din     (_zz_4072[31:0]         ), //i
    .dout    (fixTo_1831_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1832 (
    .din     (_zz_4073[31:0]         ), //i
    .dout    (fixTo_1832_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1833 (
    .din     (_zz_4074[31:0]         ), //i
    .dout    (fixTo_1833_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1834 (
    .din     (_zz_4075[31:0]         ), //i
    .dout    (fixTo_1834_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1835 (
    .din     (_zz_4076[31:0]         ), //i
    .dout    (fixTo_1835_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_1836 (
    .din     (_zz_4077[31:0]         ), //i
    .dout    (fixTo_1836_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_1837 (
    .din     (_zz_4078[31:0]         ), //i
    .dout    (fixTo_1837_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1838 (
    .din     (_zz_4079[31:0]         ), //i
    .dout    (fixTo_1838_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1839 (
    .din     (_zz_4080[31:0]         ), //i
    .dout    (fixTo_1839_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1840 (
    .din     (_zz_4081[31:0]         ), //i
    .dout    (fixTo_1840_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1841 (
    .din     (_zz_4082[31:0]         ), //i
    .dout    (fixTo_1841_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_1842 (
    .din     (_zz_4083[31:0]         ), //i
    .dout    (fixTo_1842_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_1843 (
    .din     (_zz_4084[31:0]         ), //i
    .dout    (fixTo_1843_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1844 (
    .din     (_zz_4085[31:0]         ), //i
    .dout    (fixTo_1844_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1845 (
    .din     (_zz_4086[31:0]         ), //i
    .dout    (fixTo_1845_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1846 (
    .din     (_zz_4087[31:0]         ), //i
    .dout    (fixTo_1846_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1847 (
    .din     (_zz_4088[31:0]         ), //i
    .dout    (fixTo_1847_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_1848 (
    .din     (_zz_4089[31:0]         ), //i
    .dout    (fixTo_1848_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_1849 (
    .din     (_zz_4090[31:0]         ), //i
    .dout    (fixTo_1849_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1850 (
    .din     (_zz_4091[31:0]         ), //i
    .dout    (fixTo_1850_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1851 (
    .din     (_zz_4092[31:0]         ), //i
    .dout    (fixTo_1851_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1852 (
    .din     (_zz_4093[31:0]         ), //i
    .dout    (fixTo_1852_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1853 (
    .din     (_zz_4094[31:0]         ), //i
    .dout    (fixTo_1853_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_1854 (
    .din     (_zz_4095[31:0]         ), //i
    .dout    (fixTo_1854_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_1855 (
    .din     (_zz_4096[31:0]         ), //i
    .dout    (fixTo_1855_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1856 (
    .din     (_zz_4097[31:0]         ), //i
    .dout    (fixTo_1856_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1857 (
    .din     (_zz_4098[31:0]         ), //i
    .dout    (fixTo_1857_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1858 (
    .din     (_zz_4099[31:0]         ), //i
    .dout    (fixTo_1858_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1859 (
    .din     (_zz_4100[31:0]         ), //i
    .dout    (fixTo_1859_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_1860 (
    .din     (_zz_4101[31:0]         ), //i
    .dout    (fixTo_1860_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_1861 (
    .din     (_zz_4102[31:0]         ), //i
    .dout    (fixTo_1861_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1862 (
    .din     (_zz_4103[31:0]         ), //i
    .dout    (fixTo_1862_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1863 (
    .din     (_zz_4104[31:0]         ), //i
    .dout    (fixTo_1863_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1864 (
    .din     (_zz_4105[31:0]         ), //i
    .dout    (fixTo_1864_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1865 (
    .din     (_zz_4106[31:0]         ), //i
    .dout    (fixTo_1865_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_1866 (
    .din     (_zz_4107[31:0]         ), //i
    .dout    (fixTo_1866_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_1867 (
    .din     (_zz_4108[31:0]         ), //i
    .dout    (fixTo_1867_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1868 (
    .din     (_zz_4109[31:0]         ), //i
    .dout    (fixTo_1868_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1869 (
    .din     (_zz_4110[31:0]         ), //i
    .dout    (fixTo_1869_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1870 (
    .din     (_zz_4111[31:0]         ), //i
    .dout    (fixTo_1870_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1871 (
    .din     (_zz_4112[31:0]         ), //i
    .dout    (fixTo_1871_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_1872 (
    .din     (_zz_4113[31:0]         ), //i
    .dout    (fixTo_1872_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_1873 (
    .din     (_zz_4114[31:0]         ), //i
    .dout    (fixTo_1873_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1874 (
    .din     (_zz_4115[31:0]         ), //i
    .dout    (fixTo_1874_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1875 (
    .din     (_zz_4116[31:0]         ), //i
    .dout    (fixTo_1875_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1876 (
    .din     (_zz_4117[31:0]         ), //i
    .dout    (fixTo_1876_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1877 (
    .din     (_zz_4118[31:0]         ), //i
    .dout    (fixTo_1877_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_1878 (
    .din     (_zz_4119[31:0]         ), //i
    .dout    (fixTo_1878_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_1879 (
    .din     (_zz_4120[31:0]         ), //i
    .dout    (fixTo_1879_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1880 (
    .din     (_zz_4121[31:0]         ), //i
    .dout    (fixTo_1880_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1881 (
    .din     (_zz_4122[31:0]         ), //i
    .dout    (fixTo_1881_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1882 (
    .din     (_zz_4123[31:0]         ), //i
    .dout    (fixTo_1882_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1883 (
    .din     (_zz_4124[31:0]         ), //i
    .dout    (fixTo_1883_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_1884 (
    .din     (_zz_4125[31:0]         ), //i
    .dout    (fixTo_1884_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_1885 (
    .din     (_zz_4126[31:0]         ), //i
    .dout    (fixTo_1885_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1886 (
    .din     (_zz_4127[31:0]         ), //i
    .dout    (fixTo_1886_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1887 (
    .din     (_zz_4128[31:0]         ), //i
    .dout    (fixTo_1887_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1888 (
    .din     (_zz_4129[31:0]         ), //i
    .dout    (fixTo_1888_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1889 (
    .din     (_zz_4130[31:0]         ), //i
    .dout    (fixTo_1889_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_1890 (
    .din     (_zz_4131[31:0]         ), //i
    .dout    (fixTo_1890_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_1891 (
    .din     (_zz_4132[31:0]         ), //i
    .dout    (fixTo_1891_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1892 (
    .din     (_zz_4133[31:0]         ), //i
    .dout    (fixTo_1892_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1893 (
    .din     (_zz_4134[31:0]         ), //i
    .dout    (fixTo_1893_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1894 (
    .din     (_zz_4135[31:0]         ), //i
    .dout    (fixTo_1894_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1895 (
    .din     (_zz_4136[31:0]         ), //i
    .dout    (fixTo_1895_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_1896 (
    .din     (_zz_4137[31:0]         ), //i
    .dout    (fixTo_1896_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_1897 (
    .din     (_zz_4138[31:0]         ), //i
    .dout    (fixTo_1897_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1898 (
    .din     (_zz_4139[31:0]         ), //i
    .dout    (fixTo_1898_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1899 (
    .din     (_zz_4140[31:0]         ), //i
    .dout    (fixTo_1899_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1900 (
    .din     (_zz_4141[31:0]         ), //i
    .dout    (fixTo_1900_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1901 (
    .din     (_zz_4142[31:0]         ), //i
    .dout    (fixTo_1901_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_1902 (
    .din     (_zz_4143[31:0]         ), //i
    .dout    (fixTo_1902_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_1903 (
    .din     (_zz_4144[31:0]         ), //i
    .dout    (fixTo_1903_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1904 (
    .din     (_zz_4145[31:0]         ), //i
    .dout    (fixTo_1904_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1905 (
    .din     (_zz_4146[31:0]         ), //i
    .dout    (fixTo_1905_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1906 (
    .din     (_zz_4147[31:0]         ), //i
    .dout    (fixTo_1906_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1907 (
    .din     (_zz_4148[31:0]         ), //i
    .dout    (fixTo_1907_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_1908 (
    .din     (_zz_4149[31:0]         ), //i
    .dout    (fixTo_1908_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_1909 (
    .din     (_zz_4150[31:0]         ), //i
    .dout    (fixTo_1909_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1910 (
    .din     (_zz_4151[31:0]         ), //i
    .dout    (fixTo_1910_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1911 (
    .din     (_zz_4152[31:0]         ), //i
    .dout    (fixTo_1911_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1912 (
    .din     (_zz_4153[31:0]         ), //i
    .dout    (fixTo_1912_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1913 (
    .din     (_zz_4154[31:0]         ), //i
    .dout    (fixTo_1913_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_1914 (
    .din     (_zz_4155[31:0]         ), //i
    .dout    (fixTo_1914_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_1915 (
    .din     (_zz_4156[31:0]         ), //i
    .dout    (fixTo_1915_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1916 (
    .din     (_zz_4157[31:0]         ), //i
    .dout    (fixTo_1916_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1917 (
    .din     (_zz_4158[31:0]         ), //i
    .dout    (fixTo_1917_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1918 (
    .din     (_zz_4159[31:0]         ), //i
    .dout    (fixTo_1918_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1919 (
    .din     (_zz_4160[31:0]         ), //i
    .dout    (fixTo_1919_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_1920 (
    .din     (_zz_4161[31:0]         ), //i
    .dout    (fixTo_1920_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_1921 (
    .din     (_zz_4162[31:0]         ), //i
    .dout    (fixTo_1921_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1922 (
    .din     (_zz_4163[31:0]         ), //i
    .dout    (fixTo_1922_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1923 (
    .din     (_zz_4164[31:0]         ), //i
    .dout    (fixTo_1923_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1924 (
    .din     (_zz_4165[31:0]         ), //i
    .dout    (fixTo_1924_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1925 (
    .din     (_zz_4166[31:0]         ), //i
    .dout    (fixTo_1925_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_1926 (
    .din     (_zz_4167[31:0]         ), //i
    .dout    (fixTo_1926_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_1927 (
    .din     (_zz_4168[31:0]         ), //i
    .dout    (fixTo_1927_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1928 (
    .din     (_zz_4169[31:0]         ), //i
    .dout    (fixTo_1928_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1929 (
    .din     (_zz_4170[31:0]         ), //i
    .dout    (fixTo_1929_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1930 (
    .din     (_zz_4171[31:0]         ), //i
    .dout    (fixTo_1930_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1931 (
    .din     (_zz_4172[31:0]         ), //i
    .dout    (fixTo_1931_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_1932 (
    .din     (_zz_4173[31:0]         ), //i
    .dout    (fixTo_1932_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_1933 (
    .din     (_zz_4174[31:0]         ), //i
    .dout    (fixTo_1933_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1934 (
    .din     (_zz_4175[31:0]         ), //i
    .dout    (fixTo_1934_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1935 (
    .din     (_zz_4176[31:0]         ), //i
    .dout    (fixTo_1935_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1936 (
    .din     (_zz_4177[31:0]         ), //i
    .dout    (fixTo_1936_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1937 (
    .din     (_zz_4178[31:0]         ), //i
    .dout    (fixTo_1937_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_1938 (
    .din     (_zz_4179[31:0]         ), //i
    .dout    (fixTo_1938_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_1939 (
    .din     (_zz_4180[31:0]         ), //i
    .dout    (fixTo_1939_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1940 (
    .din     (_zz_4181[31:0]         ), //i
    .dout    (fixTo_1940_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1941 (
    .din     (_zz_4182[31:0]         ), //i
    .dout    (fixTo_1941_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1942 (
    .din     (_zz_4183[31:0]         ), //i
    .dout    (fixTo_1942_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1943 (
    .din     (_zz_4184[31:0]         ), //i
    .dout    (fixTo_1943_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_1944 (
    .din     (_zz_4185[31:0]         ), //i
    .dout    (fixTo_1944_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_1945 (
    .din     (_zz_4186[31:0]         ), //i
    .dout    (fixTo_1945_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1946 (
    .din     (_zz_4187[31:0]         ), //i
    .dout    (fixTo_1946_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1947 (
    .din     (_zz_4188[31:0]         ), //i
    .dout    (fixTo_1947_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1948 (
    .din     (_zz_4189[31:0]         ), //i
    .dout    (fixTo_1948_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1949 (
    .din     (_zz_4190[31:0]         ), //i
    .dout    (fixTo_1949_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_1950 (
    .din     (_zz_4191[31:0]         ), //i
    .dout    (fixTo_1950_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_1951 (
    .din     (_zz_4192[31:0]         ), //i
    .dout    (fixTo_1951_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1952 (
    .din     (_zz_4193[31:0]         ), //i
    .dout    (fixTo_1952_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1953 (
    .din     (_zz_4194[31:0]         ), //i
    .dout    (fixTo_1953_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1954 (
    .din     (_zz_4195[31:0]         ), //i
    .dout    (fixTo_1954_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1955 (
    .din     (_zz_4196[31:0]         ), //i
    .dout    (fixTo_1955_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_1956 (
    .din     (_zz_4197[31:0]         ), //i
    .dout    (fixTo_1956_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_1957 (
    .din     (_zz_4198[31:0]         ), //i
    .dout    (fixTo_1957_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1958 (
    .din     (_zz_4199[31:0]         ), //i
    .dout    (fixTo_1958_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1959 (
    .din     (_zz_4200[31:0]         ), //i
    .dout    (fixTo_1959_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1960 (
    .din     (_zz_4201[31:0]         ), //i
    .dout    (fixTo_1960_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1961 (
    .din     (_zz_4202[31:0]         ), //i
    .dout    (fixTo_1961_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_1962 (
    .din     (_zz_4203[31:0]         ), //i
    .dout    (fixTo_1962_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_1963 (
    .din     (_zz_4204[31:0]         ), //i
    .dout    (fixTo_1963_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1964 (
    .din     (_zz_4205[31:0]         ), //i
    .dout    (fixTo_1964_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1965 (
    .din     (_zz_4206[31:0]         ), //i
    .dout    (fixTo_1965_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1966 (
    .din     (_zz_4207[31:0]         ), //i
    .dout    (fixTo_1966_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1967 (
    .din     (_zz_4208[31:0]         ), //i
    .dout    (fixTo_1967_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_1968 (
    .din     (_zz_4209[31:0]         ), //i
    .dout    (fixTo_1968_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_1969 (
    .din     (_zz_4210[31:0]         ), //i
    .dout    (fixTo_1969_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1970 (
    .din     (_zz_4211[31:0]         ), //i
    .dout    (fixTo_1970_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1971 (
    .din     (_zz_4212[31:0]         ), //i
    .dout    (fixTo_1971_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1972 (
    .din     (_zz_4213[31:0]         ), //i
    .dout    (fixTo_1972_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1973 (
    .din     (_zz_4214[31:0]         ), //i
    .dout    (fixTo_1973_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_1974 (
    .din     (_zz_4215[31:0]         ), //i
    .dout    (fixTo_1974_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_1975 (
    .din     (_zz_4216[31:0]         ), //i
    .dout    (fixTo_1975_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1976 (
    .din     (_zz_4217[31:0]         ), //i
    .dout    (fixTo_1976_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1977 (
    .din     (_zz_4218[31:0]         ), //i
    .dout    (fixTo_1977_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1978 (
    .din     (_zz_4219[31:0]         ), //i
    .dout    (fixTo_1978_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1979 (
    .din     (_zz_4220[31:0]         ), //i
    .dout    (fixTo_1979_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_1980 (
    .din     (_zz_4221[31:0]         ), //i
    .dout    (fixTo_1980_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_1981 (
    .din     (_zz_4222[31:0]         ), //i
    .dout    (fixTo_1981_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1982 (
    .din     (_zz_4223[31:0]         ), //i
    .dout    (fixTo_1982_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1983 (
    .din     (_zz_4224[31:0]         ), //i
    .dout    (fixTo_1983_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1984 (
    .din     (_zz_4225[31:0]         ), //i
    .dout    (fixTo_1984_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1985 (
    .din     (_zz_4226[31:0]         ), //i
    .dout    (fixTo_1985_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_1986 (
    .din     (_zz_4227[31:0]         ), //i
    .dout    (fixTo_1986_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_1987 (
    .din     (_zz_4228[31:0]         ), //i
    .dout    (fixTo_1987_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1988 (
    .din     (_zz_4229[31:0]         ), //i
    .dout    (fixTo_1988_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1989 (
    .din     (_zz_4230[31:0]         ), //i
    .dout    (fixTo_1989_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1990 (
    .din     (_zz_4231[31:0]         ), //i
    .dout    (fixTo_1990_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1991 (
    .din     (_zz_4232[31:0]         ), //i
    .dout    (fixTo_1991_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_1992 (
    .din     (_zz_4233[31:0]         ), //i
    .dout    (fixTo_1992_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_1993 (
    .din     (_zz_4234[31:0]         ), //i
    .dout    (fixTo_1993_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1994 (
    .din     (_zz_4235[31:0]         ), //i
    .dout    (fixTo_1994_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1995 (
    .din     (_zz_4236[31:0]         ), //i
    .dout    (fixTo_1995_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1996 (
    .din     (_zz_4237[31:0]         ), //i
    .dout    (fixTo_1996_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_1997 (
    .din     (_zz_4238[31:0]         ), //i
    .dout    (fixTo_1997_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_1998 (
    .din     (_zz_4239[31:0]         ), //i
    .dout    (fixTo_1998_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_1999 (
    .din     (_zz_4240[31:0]         ), //i
    .dout    (fixTo_1999_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_2000 (
    .din     (_zz_4241[31:0]         ), //i
    .dout    (fixTo_2000_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_2001 (
    .din     (_zz_4242[31:0]         ), //i
    .dout    (fixTo_2001_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_2002 (
    .din     (_zz_4243[31:0]         ), //i
    .dout    (fixTo_2002_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_2003 (
    .din     (_zz_4244[31:0]         ), //i
    .dout    (fixTo_2003_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_2004 (
    .din     (_zz_4245[31:0]         ), //i
    .dout    (fixTo_2004_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_2005 (
    .din     (_zz_4246[31:0]         ), //i
    .dout    (fixTo_2005_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_2006 (
    .din     (_zz_4247[31:0]         ), //i
    .dout    (fixTo_2006_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_2007 (
    .din     (_zz_4248[31:0]         ), //i
    .dout    (fixTo_2007_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_2008 (
    .din     (_zz_4249[31:0]         ), //i
    .dout    (fixTo_2008_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_2009 (
    .din     (_zz_4250[31:0]         ), //i
    .dout    (fixTo_2009_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_2010 (
    .din     (_zz_4251[31:0]         ), //i
    .dout    (fixTo_2010_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_2011 (
    .din     (_zz_4252[31:0]         ), //i
    .dout    (fixTo_2011_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_2012 (
    .din     (_zz_4253[31:0]         ), //i
    .dout    (fixTo_2012_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_2013 (
    .din     (_zz_4254[31:0]         ), //i
    .dout    (fixTo_2013_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_2014 (
    .din     (_zz_4255[31:0]         ), //i
    .dout    (fixTo_2014_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_2015 (
    .din     (_zz_4256[31:0]         ), //i
    .dout    (fixTo_2015_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_2016 (
    .din     (_zz_4257[31:0]         ), //i
    .dout    (fixTo_2016_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_2017 (
    .din     (_zz_4258[31:0]         ), //i
    .dout    (fixTo_2017_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_2018 (
    .din     (_zz_4259[31:0]         ), //i
    .dout    (fixTo_2018_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_2019 (
    .din     (_zz_4260[31:0]         ), //i
    .dout    (fixTo_2019_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_2020 (
    .din     (_zz_4261[31:0]         ), //i
    .dout    (fixTo_2020_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_2021 (
    .din     (_zz_4262[31:0]         ), //i
    .dout    (fixTo_2021_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_2022 (
    .din     (_zz_4263[31:0]         ), //i
    .dout    (fixTo_2022_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_2023 (
    .din     (_zz_4264[31:0]         ), //i
    .dout    (fixTo_2023_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_2024 (
    .din     (_zz_4265[31:0]         ), //i
    .dout    (fixTo_2024_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_2025 (
    .din     (_zz_4266[31:0]         ), //i
    .dout    (fixTo_2025_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_2026 (
    .din     (_zz_4267[31:0]         ), //i
    .dout    (fixTo_2026_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_2027 (
    .din     (_zz_4268[31:0]         ), //i
    .dout    (fixTo_2027_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_2028 (
    .din     (_zz_4269[31:0]         ), //i
    .dout    (fixTo_2028_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_2029 (
    .din     (_zz_4270[31:0]         ), //i
    .dout    (fixTo_2029_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_2030 (
    .din     (_zz_4271[31:0]         ), //i
    .dout    (fixTo_2030_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_2031 (
    .din     (_zz_4272[31:0]         ), //i
    .dout    (fixTo_2031_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_2032 (
    .din     (_zz_4273[31:0]         ), //i
    .dout    (fixTo_2032_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_2033 (
    .din     (_zz_4274[31:0]         ), //i
    .dout    (fixTo_2033_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_2034 (
    .din     (_zz_4275[31:0]         ), //i
    .dout    (fixTo_2034_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_2035 (
    .din     (_zz_4276[31:0]         ), //i
    .dout    (fixTo_2035_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_2036 (
    .din     (_zz_4277[31:0]         ), //i
    .dout    (fixTo_2036_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_2037 (
    .din     (_zz_4278[31:0]         ), //i
    .dout    (fixTo_2037_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_2038 (
    .din     (_zz_4279[31:0]         ), //i
    .dout    (fixTo_2038_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_2039 (
    .din     (_zz_4280[31:0]         ), //i
    .dout    (fixTo_2039_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_2040 (
    .din     (_zz_4281[31:0]         ), //i
    .dout    (fixTo_2040_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_2041 (
    .din     (_zz_4282[31:0]         ), //i
    .dout    (fixTo_2041_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_2042 (
    .din     (_zz_4283[31:0]         ), //i
    .dout    (fixTo_2042_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_2043 (
    .din     (_zz_4284[31:0]         ), //i
    .dout    (fixTo_2043_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_2044 (
    .din     (_zz_4285[31:0]         ), //i
    .dout    (fixTo_2044_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_2045 (
    .din     (_zz_4286[31:0]         ), //i
    .dout    (fixTo_2045_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_2046 (
    .din     (_zz_4287[31:0]         ), //i
    .dout    (fixTo_2046_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_2047 (
    .din     (_zz_4288[31:0]         ), //i
    .dout    (fixTo_2047_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_2048 (
    .din     (_zz_4289[31:0]         ), //i
    .dout    (fixTo_2048_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_2049 (
    .din     (_zz_4290[31:0]         ), //i
    .dout    (fixTo_2049_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_2050 (
    .din     (_zz_4291[31:0]         ), //i
    .dout    (fixTo_2050_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_2051 (
    .din     (_zz_4292[31:0]         ), //i
    .dout    (fixTo_2051_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_2052 (
    .din     (_zz_4293[31:0]         ), //i
    .dout    (fixTo_2052_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_2053 (
    .din     (_zz_4294[31:0]         ), //i
    .dout    (fixTo_2053_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_2054 (
    .din     (_zz_4295[31:0]         ), //i
    .dout    (fixTo_2054_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_2055 (
    .din     (_zz_4296[31:0]         ), //i
    .dout    (fixTo_2055_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_2056 (
    .din     (_zz_4297[31:0]         ), //i
    .dout    (fixTo_2056_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_2057 (
    .din     (_zz_4298[31:0]         ), //i
    .dout    (fixTo_2057_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_2058 (
    .din     (_zz_4299[31:0]         ), //i
    .dout    (fixTo_2058_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_2059 (
    .din     (_zz_4300[31:0]         ), //i
    .dout    (fixTo_2059_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_2060 (
    .din     (_zz_4301[31:0]         ), //i
    .dout    (fixTo_2060_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_2061 (
    .din     (_zz_4302[31:0]         ), //i
    .dout    (fixTo_2061_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_2062 (
    .din     (_zz_4303[31:0]         ), //i
    .dout    (fixTo_2062_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_2063 (
    .din     (_zz_4304[31:0]         ), //i
    .dout    (fixTo_2063_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_2064 (
    .din     (_zz_4305[31:0]         ), //i
    .dout    (fixTo_2064_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_2065 (
    .din     (_zz_4306[31:0]         ), //i
    .dout    (fixTo_2065_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_2066 (
    .din     (_zz_4307[31:0]         ), //i
    .dout    (fixTo_2066_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_2067 (
    .din     (_zz_4308[31:0]         ), //i
    .dout    (fixTo_2067_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_2068 (
    .din     (_zz_4309[31:0]         ), //i
    .dout    (fixTo_2068_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_2069 (
    .din     (_zz_4310[31:0]         ), //i
    .dout    (fixTo_2069_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_2070 (
    .din     (_zz_4311[31:0]         ), //i
    .dout    (fixTo_2070_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_2071 (
    .din     (_zz_4312[31:0]         ), //i
    .dout    (fixTo_2071_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_2072 (
    .din     (_zz_4313[31:0]         ), //i
    .dout    (fixTo_2072_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_2073 (
    .din     (_zz_4314[31:0]         ), //i
    .dout    (fixTo_2073_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_2074 (
    .din     (_zz_4315[31:0]         ), //i
    .dout    (fixTo_2074_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_2075 (
    .din     (_zz_4316[31:0]         ), //i
    .dout    (fixTo_2075_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_2076 (
    .din     (_zz_4317[31:0]         ), //i
    .dout    (fixTo_2076_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_2077 (
    .din     (_zz_4318[31:0]         ), //i
    .dout    (fixTo_2077_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_2078 (
    .din     (_zz_4319[31:0]         ), //i
    .dout    (fixTo_2078_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_2079 (
    .din     (_zz_4320[31:0]         ), //i
    .dout    (fixTo_2079_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_2080 (
    .din     (_zz_4321[31:0]         ), //i
    .dout    (fixTo_2080_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_2081 (
    .din     (_zz_4322[31:0]         ), //i
    .dout    (fixTo_2081_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_2082 (
    .din     (_zz_4323[31:0]         ), //i
    .dout    (fixTo_2082_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_2083 (
    .din     (_zz_4324[31:0]         ), //i
    .dout    (fixTo_2083_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_2084 (
    .din     (_zz_4325[31:0]         ), //i
    .dout    (fixTo_2084_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_2085 (
    .din     (_zz_4326[31:0]         ), //i
    .dout    (fixTo_2085_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_2086 (
    .din     (_zz_4327[31:0]         ), //i
    .dout    (fixTo_2086_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_2087 (
    .din     (_zz_4328[31:0]         ), //i
    .dout    (fixTo_2087_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_2088 (
    .din     (_zz_4329[31:0]         ), //i
    .dout    (fixTo_2088_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_2089 (
    .din     (_zz_4330[31:0]         ), //i
    .dout    (fixTo_2089_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_2090 (
    .din     (_zz_4331[31:0]         ), //i
    .dout    (fixTo_2090_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_2091 (
    .din     (_zz_4332[31:0]         ), //i
    .dout    (fixTo_2091_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_2092 (
    .din     (_zz_4333[31:0]         ), //i
    .dout    (fixTo_2092_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_2093 (
    .din     (_zz_4334[31:0]         ), //i
    .dout    (fixTo_2093_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_2094 (
    .din     (_zz_4335[31:0]         ), //i
    .dout    (fixTo_2094_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_2095 (
    .din     (_zz_4336[31:0]         ), //i
    .dout    (fixTo_2095_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_2096 (
    .din     (_zz_4337[31:0]         ), //i
    .dout    (fixTo_2096_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_2097 (
    .din     (_zz_4338[31:0]         ), //i
    .dout    (fixTo_2097_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_2098 (
    .din     (_zz_4339[31:0]         ), //i
    .dout    (fixTo_2098_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_2099 (
    .din     (_zz_4340[31:0]         ), //i
    .dout    (fixTo_2099_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_2100 (
    .din     (_zz_4341[31:0]         ), //i
    .dout    (fixTo_2100_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_2101 (
    .din     (_zz_4342[31:0]         ), //i
    .dout    (fixTo_2101_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_2102 (
    .din     (_zz_4343[31:0]         ), //i
    .dout    (fixTo_2102_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_2103 (
    .din     (_zz_4344[31:0]         ), //i
    .dout    (fixTo_2103_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_2104 (
    .din     (_zz_4345[31:0]         ), //i
    .dout    (fixTo_2104_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_2105 (
    .din     (_zz_4346[31:0]         ), //i
    .dout    (fixTo_2105_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_2106 (
    .din     (_zz_4347[31:0]         ), //i
    .dout    (fixTo_2106_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_2107 (
    .din     (_zz_4348[31:0]         ), //i
    .dout    (fixTo_2107_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_2108 (
    .din     (_zz_4349[31:0]         ), //i
    .dout    (fixTo_2108_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_2109 (
    .din     (_zz_4350[31:0]         ), //i
    .dout    (fixTo_2109_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_2110 (
    .din     (_zz_4351[31:0]         ), //i
    .dout    (fixTo_2110_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_2111 (
    .din     (_zz_4352[31:0]         ), //i
    .dout    (fixTo_2111_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_2112 (
    .din     (_zz_4353[31:0]         ), //i
    .dout    (fixTo_2112_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_2113 (
    .din     (_zz_4354[31:0]         ), //i
    .dout    (fixTo_2113_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_2114 (
    .din     (_zz_4355[31:0]         ), //i
    .dout    (fixTo_2114_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_2115 (
    .din     (_zz_4356[31:0]         ), //i
    .dout    (fixTo_2115_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_2116 (
    .din     (_zz_4357[31:0]         ), //i
    .dout    (fixTo_2116_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_2117 (
    .din     (_zz_4358[31:0]         ), //i
    .dout    (fixTo_2117_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_2118 (
    .din     (_zz_4359[31:0]         ), //i
    .dout    (fixTo_2118_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_2119 (
    .din     (_zz_4360[31:0]         ), //i
    .dout    (fixTo_2119_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_2120 (
    .din     (_zz_4361[31:0]         ), //i
    .dout    (fixTo_2120_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_2121 (
    .din     (_zz_4362[31:0]         ), //i
    .dout    (fixTo_2121_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_2122 (
    .din     (_zz_4363[31:0]         ), //i
    .dout    (fixTo_2122_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_2123 (
    .din     (_zz_4364[31:0]         ), //i
    .dout    (fixTo_2123_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_2124 (
    .din     (_zz_4365[31:0]         ), //i
    .dout    (fixTo_2124_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_2125 (
    .din     (_zz_4366[31:0]         ), //i
    .dout    (fixTo_2125_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_2126 (
    .din     (_zz_4367[31:0]         ), //i
    .dout    (fixTo_2126_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_2127 (
    .din     (_zz_4368[31:0]         ), //i
    .dout    (fixTo_2127_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_2128 (
    .din     (_zz_4369[31:0]         ), //i
    .dout    (fixTo_2128_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_2129 (
    .din     (_zz_4370[31:0]         ), //i
    .dout    (fixTo_2129_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_2130 (
    .din     (_zz_4371[31:0]         ), //i
    .dout    (fixTo_2130_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_2131 (
    .din     (_zz_4372[31:0]         ), //i
    .dout    (fixTo_2131_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_2132 (
    .din     (_zz_4373[31:0]         ), //i
    .dout    (fixTo_2132_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_2133 (
    .din     (_zz_4374[31:0]         ), //i
    .dout    (fixTo_2133_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_2134 (
    .din     (_zz_4375[31:0]         ), //i
    .dout    (fixTo_2134_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_2135 (
    .din     (_zz_4376[31:0]         ), //i
    .dout    (fixTo_2135_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_2136 (
    .din     (_zz_4377[31:0]         ), //i
    .dout    (fixTo_2136_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_2137 (
    .din     (_zz_4378[31:0]         ), //i
    .dout    (fixTo_2137_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_2138 (
    .din     (_zz_4379[31:0]         ), //i
    .dout    (fixTo_2138_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_2139 (
    .din     (_zz_4380[31:0]         ), //i
    .dout    (fixTo_2139_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_2140 (
    .din     (_zz_4381[31:0]         ), //i
    .dout    (fixTo_2140_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_2141 (
    .din     (_zz_4382[31:0]         ), //i
    .dout    (fixTo_2141_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_2142 (
    .din     (_zz_4383[31:0]         ), //i
    .dout    (fixTo_2142_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_2143 (
    .din     (_zz_4384[31:0]         ), //i
    .dout    (fixTo_2143_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_2144 (
    .din     (_zz_4385[31:0]         ), //i
    .dout    (fixTo_2144_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_2145 (
    .din     (_zz_4386[31:0]         ), //i
    .dout    (fixTo_2145_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_2146 (
    .din     (_zz_4387[31:0]         ), //i
    .dout    (fixTo_2146_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_2147 (
    .din     (_zz_4388[31:0]         ), //i
    .dout    (fixTo_2147_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_2148 (
    .din     (_zz_4389[31:0]         ), //i
    .dout    (fixTo_2148_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_2149 (
    .din     (_zz_4390[31:0]         ), //i
    .dout    (fixTo_2149_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_2150 (
    .din     (_zz_4391[31:0]         ), //i
    .dout    (fixTo_2150_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_2151 (
    .din     (_zz_4392[31:0]         ), //i
    .dout    (fixTo_2151_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_2152 (
    .din     (_zz_4393[31:0]         ), //i
    .dout    (fixTo_2152_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_2153 (
    .din     (_zz_4394[31:0]         ), //i
    .dout    (fixTo_2153_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_2154 (
    .din     (_zz_4395[31:0]         ), //i
    .dout    (fixTo_2154_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_2155 (
    .din     (_zz_4396[31:0]         ), //i
    .dout    (fixTo_2155_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_2156 (
    .din     (_zz_4397[31:0]         ), //i
    .dout    (fixTo_2156_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_2157 (
    .din     (_zz_4398[31:0]         ), //i
    .dout    (fixTo_2157_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_2158 (
    .din     (_zz_4399[31:0]         ), //i
    .dout    (fixTo_2158_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_2159 (
    .din     (_zz_4400[31:0]         ), //i
    .dout    (fixTo_2159_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_2160 (
    .din     (_zz_4401[31:0]         ), //i
    .dout    (fixTo_2160_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_2161 (
    .din     (_zz_4402[31:0]         ), //i
    .dout    (fixTo_2161_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_2162 (
    .din     (_zz_4403[31:0]         ), //i
    .dout    (fixTo_2162_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_2163 (
    .din     (_zz_4404[31:0]         ), //i
    .dout    (fixTo_2163_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_2164 (
    .din     (_zz_4405[31:0]         ), //i
    .dout    (fixTo_2164_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_2165 (
    .din     (_zz_4406[31:0]         ), //i
    .dout    (fixTo_2165_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_2166 (
    .din     (_zz_4407[31:0]         ), //i
    .dout    (fixTo_2166_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_2167 (
    .din     (_zz_4408[31:0]         ), //i
    .dout    (fixTo_2167_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_2168 (
    .din     (_zz_4409[31:0]         ), //i
    .dout    (fixTo_2168_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_2169 (
    .din     (_zz_4410[31:0]         ), //i
    .dout    (fixTo_2169_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_2170 (
    .din     (_zz_4411[31:0]         ), //i
    .dout    (fixTo_2170_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_2171 (
    .din     (_zz_4412[31:0]         ), //i
    .dout    (fixTo_2171_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_2172 (
    .din     (_zz_4413[31:0]         ), //i
    .dout    (fixTo_2172_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_2173 (
    .din     (_zz_4414[31:0]         ), //i
    .dout    (fixTo_2173_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_2174 (
    .din     (_zz_4415[31:0]         ), //i
    .dout    (fixTo_2174_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_2175 (
    .din     (_zz_4416[31:0]         ), //i
    .dout    (fixTo_2175_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_2176 (
    .din     (_zz_4417[31:0]         ), //i
    .dout    (fixTo_2176_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_2177 (
    .din     (_zz_4418[31:0]         ), //i
    .dout    (fixTo_2177_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_2178 (
    .din     (_zz_4419[31:0]         ), //i
    .dout    (fixTo_2178_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_2179 (
    .din     (_zz_4420[31:0]         ), //i
    .dout    (fixTo_2179_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_2180 (
    .din     (_zz_4421[31:0]         ), //i
    .dout    (fixTo_2180_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_2181 (
    .din     (_zz_4422[31:0]         ), //i
    .dout    (fixTo_2181_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_2182 (
    .din     (_zz_4423[31:0]         ), //i
    .dout    (fixTo_2182_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_2183 (
    .din     (_zz_4424[31:0]         ), //i
    .dout    (fixTo_2183_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_2184 (
    .din     (_zz_4425[31:0]         ), //i
    .dout    (fixTo_2184_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_2185 (
    .din     (_zz_4426[31:0]         ), //i
    .dout    (fixTo_2185_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_2186 (
    .din     (_zz_4427[31:0]         ), //i
    .dout    (fixTo_2186_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_2187 (
    .din     (_zz_4428[31:0]         ), //i
    .dout    (fixTo_2187_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_2188 (
    .din     (_zz_4429[31:0]         ), //i
    .dout    (fixTo_2188_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_2189 (
    .din     (_zz_4430[31:0]         ), //i
    .dout    (fixTo_2189_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_2190 (
    .din     (_zz_4431[31:0]         ), //i
    .dout    (fixTo_2190_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_2191 (
    .din     (_zz_4432[31:0]         ), //i
    .dout    (fixTo_2191_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_2192 (
    .din     (_zz_4433[31:0]         ), //i
    .dout    (fixTo_2192_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_2193 (
    .din     (_zz_4434[31:0]         ), //i
    .dout    (fixTo_2193_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_2194 (
    .din     (_zz_4435[31:0]         ), //i
    .dout    (fixTo_2194_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_2195 (
    .din     (_zz_4436[31:0]         ), //i
    .dout    (fixTo_2195_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_2196 (
    .din     (_zz_4437[31:0]         ), //i
    .dout    (fixTo_2196_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_2197 (
    .din     (_zz_4438[31:0]         ), //i
    .dout    (fixTo_2197_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_2198 (
    .din     (_zz_4439[31:0]         ), //i
    .dout    (fixTo_2198_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_2199 (
    .din     (_zz_4440[31:0]         ), //i
    .dout    (fixTo_2199_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_2200 (
    .din     (_zz_4441[31:0]         ), //i
    .dout    (fixTo_2200_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_2201 (
    .din     (_zz_4442[31:0]         ), //i
    .dout    (fixTo_2201_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_2202 (
    .din     (_zz_4443[31:0]         ), //i
    .dout    (fixTo_2202_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_2203 (
    .din     (_zz_4444[31:0]         ), //i
    .dout    (fixTo_2203_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_2204 (
    .din     (_zz_4445[31:0]         ), //i
    .dout    (fixTo_2204_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_2205 (
    .din     (_zz_4446[31:0]         ), //i
    .dout    (fixTo_2205_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_2206 (
    .din     (_zz_4447[31:0]         ), //i
    .dout    (fixTo_2206_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_2207 (
    .din     (_zz_4448[31:0]         ), //i
    .dout    (fixTo_2207_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_2208 (
    .din     (_zz_4449[31:0]         ), //i
    .dout    (fixTo_2208_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_2209 (
    .din     (_zz_4450[31:0]         ), //i
    .dout    (fixTo_2209_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_2210 (
    .din     (_zz_4451[31:0]         ), //i
    .dout    (fixTo_2210_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_2211 (
    .din     (_zz_4452[31:0]         ), //i
    .dout    (fixTo_2211_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_2212 (
    .din     (_zz_4453[31:0]         ), //i
    .dout    (fixTo_2212_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_2213 (
    .din     (_zz_4454[31:0]         ), //i
    .dout    (fixTo_2213_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_2214 (
    .din     (_zz_4455[31:0]         ), //i
    .dout    (fixTo_2214_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_2215 (
    .din     (_zz_4456[31:0]         ), //i
    .dout    (fixTo_2215_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_2216 (
    .din     (_zz_4457[31:0]         ), //i
    .dout    (fixTo_2216_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_2217 (
    .din     (_zz_4458[31:0]         ), //i
    .dout    (fixTo_2217_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_2218 (
    .din     (_zz_4459[31:0]         ), //i
    .dout    (fixTo_2218_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_2219 (
    .din     (_zz_4460[31:0]         ), //i
    .dout    (fixTo_2219_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_2220 (
    .din     (_zz_4461[31:0]         ), //i
    .dout    (fixTo_2220_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_2221 (
    .din     (_zz_4462[31:0]         ), //i
    .dout    (fixTo_2221_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_2222 (
    .din     (_zz_4463[31:0]         ), //i
    .dout    (fixTo_2222_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_2223 (
    .din     (_zz_4464[31:0]         ), //i
    .dout    (fixTo_2223_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_2224 (
    .din     (_zz_4465[31:0]         ), //i
    .dout    (fixTo_2224_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_2225 (
    .din     (_zz_4466[31:0]         ), //i
    .dout    (fixTo_2225_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_2226 (
    .din     (_zz_4467[31:0]         ), //i
    .dout    (fixTo_2226_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_2227 (
    .din     (_zz_4468[31:0]         ), //i
    .dout    (fixTo_2227_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_2228 (
    .din     (_zz_4469[31:0]         ), //i
    .dout    (fixTo_2228_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_2229 (
    .din     (_zz_4470[31:0]         ), //i
    .dout    (fixTo_2229_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_2230 (
    .din     (_zz_4471[31:0]         ), //i
    .dout    (fixTo_2230_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_2231 (
    .din     (_zz_4472[31:0]         ), //i
    .dout    (fixTo_2231_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_2232 (
    .din     (_zz_4473[31:0]         ), //i
    .dout    (fixTo_2232_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_2233 (
    .din     (_zz_4474[31:0]         ), //i
    .dout    (fixTo_2233_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_2234 (
    .din     (_zz_4475[31:0]         ), //i
    .dout    (fixTo_2234_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_2235 (
    .din     (_zz_4476[31:0]         ), //i
    .dout    (fixTo_2235_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_2236 (
    .din     (_zz_4477[31:0]         ), //i
    .dout    (fixTo_2236_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_2237 (
    .din     (_zz_4478[31:0]         ), //i
    .dout    (fixTo_2237_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_2238 (
    .din     (_zz_4479[31:0]         ), //i
    .dout    (fixTo_2238_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_2239 (
    .din     (_zz_4480[31:0]         ), //i
    .dout    (fixTo_2239_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_2240 (
    .din     (_zz_4481[31:0]         ), //i
    .dout    (fixTo_2240_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_2241 (
    .din     (_zz_4482[31:0]         ), //i
    .dout    (fixTo_2241_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_2242 (
    .din     (_zz_4483[31:0]         ), //i
    .dout    (fixTo_2242_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_2243 (
    .din     (_zz_4484[31:0]         ), //i
    .dout    (fixTo_2243_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_2244 (
    .din     (_zz_4485[31:0]         ), //i
    .dout    (fixTo_2244_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_2245 (
    .din     (_zz_4486[31:0]         ), //i
    .dout    (fixTo_2245_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_2246 (
    .din     (_zz_4487[31:0]         ), //i
    .dout    (fixTo_2246_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_2247 (
    .din     (_zz_4488[31:0]         ), //i
    .dout    (fixTo_2247_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_2248 (
    .din     (_zz_4489[31:0]         ), //i
    .dout    (fixTo_2248_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_2249 (
    .din     (_zz_4490[31:0]         ), //i
    .dout    (fixTo_2249_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_2250 (
    .din     (_zz_4491[31:0]         ), //i
    .dout    (fixTo_2250_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_2251 (
    .din     (_zz_4492[31:0]         ), //i
    .dout    (fixTo_2251_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_2252 (
    .din     (_zz_4493[31:0]         ), //i
    .dout    (fixTo_2252_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_2253 (
    .din     (_zz_4494[31:0]         ), //i
    .dout    (fixTo_2253_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_2254 (
    .din     (_zz_4495[31:0]         ), //i
    .dout    (fixTo_2254_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_2255 (
    .din     (_zz_4496[31:0]         ), //i
    .dout    (fixTo_2255_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_2256 (
    .din     (_zz_4497[31:0]         ), //i
    .dout    (fixTo_2256_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_2257 (
    .din     (_zz_4498[31:0]         ), //i
    .dout    (fixTo_2257_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_2258 (
    .din     (_zz_4499[31:0]         ), //i
    .dout    (fixTo_2258_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_2259 (
    .din     (_zz_4500[31:0]         ), //i
    .dout    (fixTo_2259_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_2260 (
    .din     (_zz_4501[31:0]         ), //i
    .dout    (fixTo_2260_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_2261 (
    .din     (_zz_4502[31:0]         ), //i
    .dout    (fixTo_2261_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_2262 (
    .din     (_zz_4503[31:0]         ), //i
    .dout    (fixTo_2262_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_2263 (
    .din     (_zz_4504[31:0]         ), //i
    .dout    (fixTo_2263_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_2264 (
    .din     (_zz_4505[31:0]         ), //i
    .dout    (fixTo_2264_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_2265 (
    .din     (_zz_4506[31:0]         ), //i
    .dout    (fixTo_2265_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_2266 (
    .din     (_zz_4507[31:0]         ), //i
    .dout    (fixTo_2266_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_2267 (
    .din     (_zz_4508[31:0]         ), //i
    .dout    (fixTo_2267_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_2268 (
    .din     (_zz_4509[31:0]         ), //i
    .dout    (fixTo_2268_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_2269 (
    .din     (_zz_4510[31:0]         ), //i
    .dout    (fixTo_2269_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_2270 (
    .din     (_zz_4511[31:0]         ), //i
    .dout    (fixTo_2270_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_2271 (
    .din     (_zz_4512[31:0]         ), //i
    .dout    (fixTo_2271_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_2272 (
    .din     (_zz_4513[31:0]         ), //i
    .dout    (fixTo_2272_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_2273 (
    .din     (_zz_4514[31:0]         ), //i
    .dout    (fixTo_2273_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_2274 (
    .din     (_zz_4515[31:0]         ), //i
    .dout    (fixTo_2274_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_2275 (
    .din     (_zz_4516[31:0]         ), //i
    .dout    (fixTo_2275_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_2276 (
    .din     (_zz_4517[31:0]         ), //i
    .dout    (fixTo_2276_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_2277 (
    .din     (_zz_4518[31:0]         ), //i
    .dout    (fixTo_2277_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_2278 (
    .din     (_zz_4519[31:0]         ), //i
    .dout    (fixTo_2278_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_2279 (
    .din     (_zz_4520[31:0]         ), //i
    .dout    (fixTo_2279_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_2280 (
    .din     (_zz_4521[31:0]         ), //i
    .dout    (fixTo_2280_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_2281 (
    .din     (_zz_4522[31:0]         ), //i
    .dout    (fixTo_2281_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_2282 (
    .din     (_zz_4523[31:0]         ), //i
    .dout    (fixTo_2282_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_2283 (
    .din     (_zz_4524[31:0]         ), //i
    .dout    (fixTo_2283_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_2284 (
    .din     (_zz_4525[31:0]         ), //i
    .dout    (fixTo_2284_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_2285 (
    .din     (_zz_4526[31:0]         ), //i
    .dout    (fixTo_2285_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_2286 (
    .din     (_zz_4527[31:0]         ), //i
    .dout    (fixTo_2286_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_2287 (
    .din     (_zz_4528[31:0]         ), //i
    .dout    (fixTo_2287_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_2288 (
    .din     (_zz_4529[31:0]         ), //i
    .dout    (fixTo_2288_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_2289 (
    .din     (_zz_4530[31:0]         ), //i
    .dout    (fixTo_2289_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_2290 (
    .din     (_zz_4531[31:0]         ), //i
    .dout    (fixTo_2290_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_2291 (
    .din     (_zz_4532[31:0]         ), //i
    .dout    (fixTo_2291_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_2292 (
    .din     (_zz_4533[31:0]         ), //i
    .dout    (fixTo_2292_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_2293 (
    .din     (_zz_4534[31:0]         ), //i
    .dout    (fixTo_2293_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_2294 (
    .din     (_zz_4535[31:0]         ), //i
    .dout    (fixTo_2294_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_2295 (
    .din     (_zz_4536[31:0]         ), //i
    .dout    (fixTo_2295_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_2296 (
    .din     (_zz_4537[31:0]         ), //i
    .dout    (fixTo_2296_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_2297 (
    .din     (_zz_4538[31:0]         ), //i
    .dout    (fixTo_2297_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_2298 (
    .din     (_zz_4539[31:0]         ), //i
    .dout    (fixTo_2298_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_2299 (
    .din     (_zz_4540[31:0]         ), //i
    .dout    (fixTo_2299_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_2300 (
    .din     (_zz_4541[31:0]         ), //i
    .dout    (fixTo_2300_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_2301 (
    .din     (_zz_4542[31:0]         ), //i
    .dout    (fixTo_2301_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_2302 (
    .din     (_zz_4543[31:0]         ), //i
    .dout    (fixTo_2302_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_2303 (
    .din     (_zz_4544[31:0]         ), //i
    .dout    (fixTo_2303_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_2304 (
    .din     (_zz_4545[31:0]         ), //i
    .dout    (fixTo_2304_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_2305 (
    .din     (_zz_4546[31:0]         ), //i
    .dout    (fixTo_2305_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_2306 (
    .din     (_zz_4547[31:0]         ), //i
    .dout    (fixTo_2306_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_2307 (
    .din     (_zz_4548[31:0]         ), //i
    .dout    (fixTo_2307_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_2308 (
    .din     (_zz_4549[31:0]         ), //i
    .dout    (fixTo_2308_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_2309 (
    .din     (_zz_4550[31:0]         ), //i
    .dout    (fixTo_2309_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_2310 (
    .din     (_zz_4551[31:0]         ), //i
    .dout    (fixTo_2310_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_2311 (
    .din     (_zz_4552[31:0]         ), //i
    .dout    (fixTo_2311_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_2312 (
    .din     (_zz_4553[31:0]         ), //i
    .dout    (fixTo_2312_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_2313 (
    .din     (_zz_4554[31:0]         ), //i
    .dout    (fixTo_2313_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_2314 (
    .din     (_zz_4555[31:0]         ), //i
    .dout    (fixTo_2314_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_2315 (
    .din     (_zz_4556[31:0]         ), //i
    .dout    (fixTo_2315_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_2316 (
    .din     (_zz_4557[31:0]         ), //i
    .dout    (fixTo_2316_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_2317 (
    .din     (_zz_4558[31:0]         ), //i
    .dout    (fixTo_2317_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_2318 (
    .din     (_zz_4559[31:0]         ), //i
    .dout    (fixTo_2318_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_2319 (
    .din     (_zz_4560[31:0]         ), //i
    .dout    (fixTo_2319_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_2320 (
    .din     (_zz_4561[31:0]         ), //i
    .dout    (fixTo_2320_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_2321 (
    .din     (_zz_4562[31:0]         ), //i
    .dout    (fixTo_2321_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_2322 (
    .din     (_zz_4563[31:0]         ), //i
    .dout    (fixTo_2322_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_2323 (
    .din     (_zz_4564[31:0]         ), //i
    .dout    (fixTo_2323_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_2324 (
    .din     (_zz_4565[31:0]         ), //i
    .dout    (fixTo_2324_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_2325 (
    .din     (_zz_4566[31:0]         ), //i
    .dout    (fixTo_2325_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_2326 (
    .din     (_zz_4567[31:0]         ), //i
    .dout    (fixTo_2326_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_2327 (
    .din     (_zz_4568[31:0]         ), //i
    .dout    (fixTo_2327_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_2328 (
    .din     (_zz_4569[31:0]         ), //i
    .dout    (fixTo_2328_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_2329 (
    .din     (_zz_4570[31:0]         ), //i
    .dout    (fixTo_2329_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_2330 (
    .din     (_zz_4571[31:0]         ), //i
    .dout    (fixTo_2330_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_2331 (
    .din     (_zz_4572[31:0]         ), //i
    .dout    (fixTo_2331_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_2332 (
    .din     (_zz_4573[31:0]         ), //i
    .dout    (fixTo_2332_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_2333 (
    .din     (_zz_4574[31:0]         ), //i
    .dout    (fixTo_2333_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_2334 (
    .din     (_zz_4575[31:0]         ), //i
    .dout    (fixTo_2334_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_2335 (
    .din     (_zz_4576[31:0]         ), //i
    .dout    (fixTo_2335_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_2336 (
    .din     (_zz_4577[31:0]         ), //i
    .dout    (fixTo_2336_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_2337 (
    .din     (_zz_4578[31:0]         ), //i
    .dout    (fixTo_2337_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_2338 (
    .din     (_zz_4579[31:0]         ), //i
    .dout    (fixTo_2338_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_2339 (
    .din     (_zz_4580[31:0]         ), //i
    .dout    (fixTo_2339_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_2340 (
    .din     (_zz_4581[31:0]         ), //i
    .dout    (fixTo_2340_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_2341 (
    .din     (_zz_4582[31:0]         ), //i
    .dout    (fixTo_2341_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_2342 (
    .din     (_zz_4583[31:0]         ), //i
    .dout    (fixTo_2342_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_2343 (
    .din     (_zz_4584[31:0]         ), //i
    .dout    (fixTo_2343_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_2344 (
    .din     (_zz_4585[31:0]         ), //i
    .dout    (fixTo_2344_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_2345 (
    .din     (_zz_4586[31:0]         ), //i
    .dout    (fixTo_2345_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_2346 (
    .din     (_zz_4587[31:0]         ), //i
    .dout    (fixTo_2346_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_2347 (
    .din     (_zz_4588[31:0]         ), //i
    .dout    (fixTo_2347_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_2348 (
    .din     (_zz_4589[31:0]         ), //i
    .dout    (fixTo_2348_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_2349 (
    .din     (_zz_4590[31:0]         ), //i
    .dout    (fixTo_2349_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_2350 (
    .din     (_zz_4591[31:0]         ), //i
    .dout    (fixTo_2350_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_2351 (
    .din     (_zz_4592[31:0]         ), //i
    .dout    (fixTo_2351_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_2352 (
    .din     (_zz_4593[31:0]         ), //i
    .dout    (fixTo_2352_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_2353 (
    .din     (_zz_4594[31:0]         ), //i
    .dout    (fixTo_2353_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_2354 (
    .din     (_zz_4595[31:0]         ), //i
    .dout    (fixTo_2354_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_2355 (
    .din     (_zz_4596[31:0]         ), //i
    .dout    (fixTo_2355_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_2356 (
    .din     (_zz_4597[31:0]         ), //i
    .dout    (fixTo_2356_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_2357 (
    .din     (_zz_4598[31:0]         ), //i
    .dout    (fixTo_2357_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_2358 (
    .din     (_zz_4599[31:0]         ), //i
    .dout    (fixTo_2358_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_2359 (
    .din     (_zz_4600[31:0]         ), //i
    .dout    (fixTo_2359_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_2360 (
    .din     (_zz_4601[31:0]         ), //i
    .dout    (fixTo_2360_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_2361 (
    .din     (_zz_4602[31:0]         ), //i
    .dout    (fixTo_2361_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_2362 (
    .din     (_zz_4603[31:0]         ), //i
    .dout    (fixTo_2362_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_2363 (
    .din     (_zz_4604[31:0]         ), //i
    .dout    (fixTo_2363_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_2364 (
    .din     (_zz_4605[31:0]         ), //i
    .dout    (fixTo_2364_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_2365 (
    .din     (_zz_4606[31:0]         ), //i
    .dout    (fixTo_2365_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_2366 (
    .din     (_zz_4607[31:0]         ), //i
    .dout    (fixTo_2366_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_2367 (
    .din     (_zz_4608[31:0]         ), //i
    .dout    (fixTo_2367_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_2368 (
    .din     (_zz_4609[31:0]         ), //i
    .dout    (fixTo_2368_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_2369 (
    .din     (_zz_4610[31:0]         ), //i
    .dout    (fixTo_2369_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_2370 (
    .din     (_zz_4611[31:0]         ), //i
    .dout    (fixTo_2370_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_2371 (
    .din     (_zz_4612[31:0]         ), //i
    .dout    (fixTo_2371_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_2372 (
    .din     (_zz_4613[31:0]         ), //i
    .dout    (fixTo_2372_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_2373 (
    .din     (_zz_4614[31:0]         ), //i
    .dout    (fixTo_2373_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_2374 (
    .din     (_zz_4615[31:0]         ), //i
    .dout    (fixTo_2374_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_2375 (
    .din     (_zz_4616[31:0]         ), //i
    .dout    (fixTo_2375_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_2376 (
    .din     (_zz_4617[31:0]         ), //i
    .dout    (fixTo_2376_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_2377 (
    .din     (_zz_4618[31:0]         ), //i
    .dout    (fixTo_2377_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_2378 (
    .din     (_zz_4619[31:0]         ), //i
    .dout    (fixTo_2378_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_2379 (
    .din     (_zz_4620[31:0]         ), //i
    .dout    (fixTo_2379_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_2380 (
    .din     (_zz_4621[31:0]         ), //i
    .dout    (fixTo_2380_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_2381 (
    .din     (_zz_4622[31:0]         ), //i
    .dout    (fixTo_2381_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_2382 (
    .din     (_zz_4623[31:0]         ), //i
    .dout    (fixTo_2382_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_2383 (
    .din     (_zz_4624[31:0]         ), //i
    .dout    (fixTo_2383_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_2384 (
    .din     (_zz_4625[31:0]         ), //i
    .dout    (fixTo_2384_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_2385 (
    .din     (_zz_4626[31:0]         ), //i
    .dout    (fixTo_2385_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_2386 (
    .din     (_zz_4627[31:0]         ), //i
    .dout    (fixTo_2386_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_2387 (
    .din     (_zz_4628[31:0]         ), //i
    .dout    (fixTo_2387_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_2388 (
    .din     (_zz_4629[31:0]         ), //i
    .dout    (fixTo_2388_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_2389 (
    .din     (_zz_4630[31:0]         ), //i
    .dout    (fixTo_2389_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_2390 (
    .din     (_zz_4631[31:0]         ), //i
    .dout    (fixTo_2390_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_2391 (
    .din     (_zz_4632[31:0]         ), //i
    .dout    (fixTo_2391_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_2392 (
    .din     (_zz_4633[31:0]         ), //i
    .dout    (fixTo_2392_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_2393 (
    .din     (_zz_4634[31:0]         ), //i
    .dout    (fixTo_2393_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_2394 (
    .din     (_zz_4635[31:0]         ), //i
    .dout    (fixTo_2394_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_2395 (
    .din     (_zz_4636[31:0]         ), //i
    .dout    (fixTo_2395_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_2396 (
    .din     (_zz_4637[31:0]         ), //i
    .dout    (fixTo_2396_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_2397 (
    .din     (_zz_4638[31:0]         ), //i
    .dout    (fixTo_2397_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_2398 (
    .din     (_zz_4639[31:0]         ), //i
    .dout    (fixTo_2398_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_2399 (
    .din     (_zz_4640[31:0]         ), //i
    .dout    (fixTo_2399_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_2400 (
    .din     (_zz_4641[31:0]         ), //i
    .dout    (fixTo_2400_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_2401 (
    .din     (_zz_4642[31:0]         ), //i
    .dout    (fixTo_2401_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_2402 (
    .din     (_zz_4643[31:0]         ), //i
    .dout    (fixTo_2402_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_2403 (
    .din     (_zz_4644[31:0]         ), //i
    .dout    (fixTo_2403_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_2404 (
    .din     (_zz_4645[31:0]         ), //i
    .dout    (fixTo_2404_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_2405 (
    .din     (_zz_4646[31:0]         ), //i
    .dout    (fixTo_2405_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_2406 (
    .din     (_zz_4647[31:0]         ), //i
    .dout    (fixTo_2406_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_2407 (
    .din     (_zz_4648[31:0]         ), //i
    .dout    (fixTo_2407_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_2408 (
    .din     (_zz_4649[31:0]         ), //i
    .dout    (fixTo_2408_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_2409 (
    .din     (_zz_4650[31:0]         ), //i
    .dout    (fixTo_2409_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_2410 (
    .din     (_zz_4651[31:0]         ), //i
    .dout    (fixTo_2410_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_2411 (
    .din     (_zz_4652[31:0]         ), //i
    .dout    (fixTo_2411_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_2412 (
    .din     (_zz_4653[31:0]         ), //i
    .dout    (fixTo_2412_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_2413 (
    .din     (_zz_4654[31:0]         ), //i
    .dout    (fixTo_2413_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_2414 (
    .din     (_zz_4655[31:0]         ), //i
    .dout    (fixTo_2414_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_2415 (
    .din     (_zz_4656[31:0]         ), //i
    .dout    (fixTo_2415_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_2416 (
    .din     (_zz_4657[31:0]         ), //i
    .dout    (fixTo_2416_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_2417 (
    .din     (_zz_4658[31:0]         ), //i
    .dout    (fixTo_2417_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_2418 (
    .din     (_zz_4659[31:0]         ), //i
    .dout    (fixTo_2418_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_2419 (
    .din     (_zz_4660[31:0]         ), //i
    .dout    (fixTo_2419_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_2420 (
    .din     (_zz_4661[31:0]         ), //i
    .dout    (fixTo_2420_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_2421 (
    .din     (_zz_4662[31:0]         ), //i
    .dout    (fixTo_2421_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_2422 (
    .din     (_zz_4663[31:0]         ), //i
    .dout    (fixTo_2422_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_2423 (
    .din     (_zz_4664[31:0]         ), //i
    .dout    (fixTo_2423_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_2424 (
    .din     (_zz_4665[31:0]         ), //i
    .dout    (fixTo_2424_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_2425 (
    .din     (_zz_4666[31:0]         ), //i
    .dout    (fixTo_2425_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_2426 (
    .din     (_zz_4667[31:0]         ), //i
    .dout    (fixTo_2426_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_2427 (
    .din     (_zz_4668[31:0]         ), //i
    .dout    (fixTo_2427_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_2428 (
    .din     (_zz_4669[31:0]         ), //i
    .dout    (fixTo_2428_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_2429 (
    .din     (_zz_4670[31:0]         ), //i
    .dout    (fixTo_2429_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_2430 (
    .din     (_zz_4671[31:0]         ), //i
    .dout    (fixTo_2430_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_2431 (
    .din     (_zz_4672[31:0]         ), //i
    .dout    (fixTo_2431_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_2432 (
    .din     (_zz_4673[31:0]         ), //i
    .dout    (fixTo_2432_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_2433 (
    .din     (_zz_4674[31:0]         ), //i
    .dout    (fixTo_2433_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_2434 (
    .din     (_zz_4675[31:0]         ), //i
    .dout    (fixTo_2434_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_2435 (
    .din     (_zz_4676[31:0]         ), //i
    .dout    (fixTo_2435_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_2436 (
    .din     (_zz_4677[31:0]         ), //i
    .dout    (fixTo_2436_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_2437 (
    .din     (_zz_4678[31:0]         ), //i
    .dout    (fixTo_2437_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_2438 (
    .din     (_zz_4679[31:0]         ), //i
    .dout    (fixTo_2438_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_2439 (
    .din     (_zz_4680[31:0]         ), //i
    .dout    (fixTo_2439_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_2440 (
    .din     (_zz_4681[31:0]         ), //i
    .dout    (fixTo_2440_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_2441 (
    .din     (_zz_4682[31:0]         ), //i
    .dout    (fixTo_2441_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_2442 (
    .din     (_zz_4683[31:0]         ), //i
    .dout    (fixTo_2442_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_2443 (
    .din     (_zz_4684[31:0]         ), //i
    .dout    (fixTo_2443_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_2444 (
    .din     (_zz_4685[31:0]         ), //i
    .dout    (fixTo_2444_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_2445 (
    .din     (_zz_4686[31:0]         ), //i
    .dout    (fixTo_2445_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_2446 (
    .din     (_zz_4687[31:0]         ), //i
    .dout    (fixTo_2446_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_2447 (
    .din     (_zz_4688[31:0]         ), //i
    .dout    (fixTo_2447_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_2448 (
    .din     (_zz_4689[31:0]         ), //i
    .dout    (fixTo_2448_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_2449 (
    .din     (_zz_4690[31:0]         ), //i
    .dout    (fixTo_2449_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_2450 (
    .din     (_zz_4691[31:0]         ), //i
    .dout    (fixTo_2450_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_2451 (
    .din     (_zz_4692[31:0]         ), //i
    .dout    (fixTo_2451_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_2452 (
    .din     (_zz_4693[31:0]         ), //i
    .dout    (fixTo_2452_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_2453 (
    .din     (_zz_4694[31:0]         ), //i
    .dout    (fixTo_2453_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_2454 (
    .din     (_zz_4695[31:0]         ), //i
    .dout    (fixTo_2454_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_2455 (
    .din     (_zz_4696[31:0]         ), //i
    .dout    (fixTo_2455_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_2456 (
    .din     (_zz_4697[31:0]         ), //i
    .dout    (fixTo_2456_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_2457 (
    .din     (_zz_4698[31:0]         ), //i
    .dout    (fixTo_2457_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_2458 (
    .din     (_zz_4699[31:0]         ), //i
    .dout    (fixTo_2458_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_2459 (
    .din     (_zz_4700[31:0]         ), //i
    .dout    (fixTo_2459_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_2460 (
    .din     (_zz_4701[31:0]         ), //i
    .dout    (fixTo_2460_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_2461 (
    .din     (_zz_4702[31:0]         ), //i
    .dout    (fixTo_2461_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_2462 (
    .din     (_zz_4703[31:0]         ), //i
    .dout    (fixTo_2462_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_2463 (
    .din     (_zz_4704[31:0]         ), //i
    .dout    (fixTo_2463_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_2464 (
    .din     (_zz_4705[31:0]         ), //i
    .dout    (fixTo_2464_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_2465 (
    .din     (_zz_4706[31:0]         ), //i
    .dout    (fixTo_2465_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_2466 (
    .din     (_zz_4707[31:0]         ), //i
    .dout    (fixTo_2466_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_2467 (
    .din     (_zz_4708[31:0]         ), //i
    .dout    (fixTo_2467_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_2468 (
    .din     (_zz_4709[31:0]         ), //i
    .dout    (fixTo_2468_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_2469 (
    .din     (_zz_4710[31:0]         ), //i
    .dout    (fixTo_2469_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_2470 (
    .din     (_zz_4711[31:0]         ), //i
    .dout    (fixTo_2470_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_2471 (
    .din     (_zz_4712[31:0]         ), //i
    .dout    (fixTo_2471_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_2472 (
    .din     (_zz_4713[31:0]         ), //i
    .dout    (fixTo_2472_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_2473 (
    .din     (_zz_4714[31:0]         ), //i
    .dout    (fixTo_2473_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_2474 (
    .din     (_zz_4715[31:0]         ), //i
    .dout    (fixTo_2474_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_2475 (
    .din     (_zz_4716[31:0]         ), //i
    .dout    (fixTo_2475_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_2476 (
    .din     (_zz_4717[31:0]         ), //i
    .dout    (fixTo_2476_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_2477 (
    .din     (_zz_4718[31:0]         ), //i
    .dout    (fixTo_2477_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_2478 (
    .din     (_zz_4719[31:0]         ), //i
    .dout    (fixTo_2478_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_2479 (
    .din     (_zz_4720[31:0]         ), //i
    .dout    (fixTo_2479_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_2480 (
    .din     (_zz_4721[31:0]         ), //i
    .dout    (fixTo_2480_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_2481 (
    .din     (_zz_4722[31:0]         ), //i
    .dout    (fixTo_2481_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_2482 (
    .din     (_zz_4723[31:0]         ), //i
    .dout    (fixTo_2482_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_2483 (
    .din     (_zz_4724[31:0]         ), //i
    .dout    (fixTo_2483_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_2484 (
    .din     (_zz_4725[31:0]         ), //i
    .dout    (fixTo_2484_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_2485 (
    .din     (_zz_4726[31:0]         ), //i
    .dout    (fixTo_2485_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_2486 (
    .din     (_zz_4727[31:0]         ), //i
    .dout    (fixTo_2486_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_2487 (
    .din     (_zz_4728[31:0]         ), //i
    .dout    (fixTo_2487_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_2488 (
    .din     (_zz_4729[31:0]         ), //i
    .dout    (fixTo_2488_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_2489 (
    .din     (_zz_4730[31:0]         ), //i
    .dout    (fixTo_2489_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_2490 (
    .din     (_zz_4731[31:0]         ), //i
    .dout    (fixTo_2490_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_2491 (
    .din     (_zz_4732[31:0]         ), //i
    .dout    (fixTo_2491_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_2492 (
    .din     (_zz_4733[31:0]         ), //i
    .dout    (fixTo_2492_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_2493 (
    .din     (_zz_4734[31:0]         ), //i
    .dout    (fixTo_2493_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_2494 (
    .din     (_zz_4735[31:0]         ), //i
    .dout    (fixTo_2494_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_2495 (
    .din     (_zz_4736[31:0]         ), //i
    .dout    (fixTo_2495_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_2496 (
    .din     (_zz_4737[31:0]         ), //i
    .dout    (fixTo_2496_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_2497 (
    .din     (_zz_4738[31:0]         ), //i
    .dout    (fixTo_2497_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_2498 (
    .din     (_zz_4739[31:0]         ), //i
    .dout    (fixTo_2498_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_2499 (
    .din     (_zz_4740[31:0]         ), //i
    .dout    (fixTo_2499_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_2500 (
    .din     (_zz_4741[31:0]         ), //i
    .dout    (fixTo_2500_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_2501 (
    .din     (_zz_4742[31:0]         ), //i
    .dout    (fixTo_2501_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_2502 (
    .din     (_zz_4743[31:0]         ), //i
    .dout    (fixTo_2502_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_2503 (
    .din     (_zz_4744[31:0]         ), //i
    .dout    (fixTo_2503_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_2504 (
    .din     (_zz_4745[31:0]         ), //i
    .dout    (fixTo_2504_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_2505 (
    .din     (_zz_4746[31:0]         ), //i
    .dout    (fixTo_2505_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_2506 (
    .din     (_zz_4747[31:0]         ), //i
    .dout    (fixTo_2506_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_2507 (
    .din     (_zz_4748[31:0]         ), //i
    .dout    (fixTo_2507_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_2508 (
    .din     (_zz_4749[31:0]         ), //i
    .dout    (fixTo_2508_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_2509 (
    .din     (_zz_4750[31:0]         ), //i
    .dout    (fixTo_2509_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_2510 (
    .din     (_zz_4751[31:0]         ), //i
    .dout    (fixTo_2510_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_2511 (
    .din     (_zz_4752[31:0]         ), //i
    .dout    (fixTo_2511_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_2512 (
    .din     (_zz_4753[31:0]         ), //i
    .dout    (fixTo_2512_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_2513 (
    .din     (_zz_4754[31:0]         ), //i
    .dout    (fixTo_2513_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_2514 (
    .din     (_zz_4755[31:0]         ), //i
    .dout    (fixTo_2514_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_2515 (
    .din     (_zz_4756[31:0]         ), //i
    .dout    (fixTo_2515_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_2516 (
    .din     (_zz_4757[31:0]         ), //i
    .dout    (fixTo_2516_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_2517 (
    .din     (_zz_4758[31:0]         ), //i
    .dout    (fixTo_2517_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_2518 (
    .din     (_zz_4759[31:0]         ), //i
    .dout    (fixTo_2518_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_2519 (
    .din     (_zz_4760[31:0]         ), //i
    .dout    (fixTo_2519_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_2520 (
    .din     (_zz_4761[31:0]         ), //i
    .dout    (fixTo_2520_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_2521 (
    .din     (_zz_4762[31:0]         ), //i
    .dout    (fixTo_2521_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_2522 (
    .din     (_zz_4763[31:0]         ), //i
    .dout    (fixTo_2522_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_2523 (
    .din     (_zz_4764[31:0]         ), //i
    .dout    (fixTo_2523_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_2524 (
    .din     (_zz_4765[31:0]         ), //i
    .dout    (fixTo_2524_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_2525 (
    .din     (_zz_4766[31:0]         ), //i
    .dout    (fixTo_2525_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_2526 (
    .din     (_zz_4767[31:0]         ), //i
    .dout    (fixTo_2526_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_2527 (
    .din     (_zz_4768[31:0]         ), //i
    .dout    (fixTo_2527_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_2528 (
    .din     (_zz_4769[31:0]         ), //i
    .dout    (fixTo_2528_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_2529 (
    .din     (_zz_4770[31:0]         ), //i
    .dout    (fixTo_2529_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_2530 (
    .din     (_zz_4771[31:0]         ), //i
    .dout    (fixTo_2530_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_2531 (
    .din     (_zz_4772[31:0]         ), //i
    .dout    (fixTo_2531_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_2532 (
    .din     (_zz_4773[31:0]         ), //i
    .dout    (fixTo_2532_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_2533 (
    .din     (_zz_4774[31:0]         ), //i
    .dout    (fixTo_2533_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_2534 (
    .din     (_zz_4775[31:0]         ), //i
    .dout    (fixTo_2534_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_2535 (
    .din     (_zz_4776[31:0]         ), //i
    .dout    (fixTo_2535_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_2536 (
    .din     (_zz_4777[31:0]         ), //i
    .dout    (fixTo_2536_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_2537 (
    .din     (_zz_4778[31:0]         ), //i
    .dout    (fixTo_2537_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_2538 (
    .din     (_zz_4779[31:0]         ), //i
    .dout    (fixTo_2538_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_2539 (
    .din     (_zz_4780[31:0]         ), //i
    .dout    (fixTo_2539_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_2540 (
    .din     (_zz_4781[31:0]         ), //i
    .dout    (fixTo_2540_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_2541 (
    .din     (_zz_4782[31:0]         ), //i
    .dout    (fixTo_2541_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_2542 (
    .din     (_zz_4783[31:0]         ), //i
    .dout    (fixTo_2542_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_2543 (
    .din     (_zz_4784[31:0]         ), //i
    .dout    (fixTo_2543_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_2544 (
    .din     (_zz_4785[31:0]         ), //i
    .dout    (fixTo_2544_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_2545 (
    .din     (_zz_4786[31:0]         ), //i
    .dout    (fixTo_2545_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_2546 (
    .din     (_zz_4787[31:0]         ), //i
    .dout    (fixTo_2546_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_2547 (
    .din     (_zz_4788[31:0]         ), //i
    .dout    (fixTo_2547_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_2548 (
    .din     (_zz_4789[31:0]         ), //i
    .dout    (fixTo_2548_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_2549 (
    .din     (_zz_4790[31:0]         ), //i
    .dout    (fixTo_2549_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_2550 (
    .din     (_zz_4791[31:0]         ), //i
    .dout    (fixTo_2550_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_2551 (
    .din     (_zz_4792[31:0]         ), //i
    .dout    (fixTo_2551_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_2552 (
    .din     (_zz_4793[31:0]         ), //i
    .dout    (fixTo_2552_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_2553 (
    .din     (_zz_4794[31:0]         ), //i
    .dout    (fixTo_2553_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_2554 (
    .din     (_zz_4795[31:0]         ), //i
    .dout    (fixTo_2554_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_2555 (
    .din     (_zz_4796[31:0]         ), //i
    .dout    (fixTo_2555_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_2556 (
    .din     (_zz_4797[31:0]         ), //i
    .dout    (fixTo_2556_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_2557 (
    .din     (_zz_4798[31:0]         ), //i
    .dout    (fixTo_2557_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_2558 (
    .din     (_zz_4799[31:0]         ), //i
    .dout    (fixTo_2558_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_2559 (
    .din     (_zz_4800[31:0]         ), //i
    .dout    (fixTo_2559_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_2560 (
    .din     (_zz_4801[31:0]         ), //i
    .dout    (fixTo_2560_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_2561 (
    .din     (_zz_4802[31:0]         ), //i
    .dout    (fixTo_2561_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_2562 (
    .din     (_zz_4803[31:0]         ), //i
    .dout    (fixTo_2562_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_2563 (
    .din     (_zz_4804[31:0]         ), //i
    .dout    (fixTo_2563_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_2564 (
    .din     (_zz_4805[31:0]         ), //i
    .dout    (fixTo_2564_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_2565 (
    .din     (_zz_4806[31:0]         ), //i
    .dout    (fixTo_2565_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_2566 (
    .din     (_zz_4807[31:0]         ), //i
    .dout    (fixTo_2566_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_2567 (
    .din     (_zz_4808[31:0]         ), //i
    .dout    (fixTo_2567_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_2568 (
    .din     (_zz_4809[31:0]         ), //i
    .dout    (fixTo_2568_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_2569 (
    .din     (_zz_4810[31:0]         ), //i
    .dout    (fixTo_2569_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_2570 (
    .din     (_zz_4811[31:0]         ), //i
    .dout    (fixTo_2570_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_2571 (
    .din     (_zz_4812[31:0]         ), //i
    .dout    (fixTo_2571_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_2572 (
    .din     (_zz_4813[31:0]         ), //i
    .dout    (fixTo_2572_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_2573 (
    .din     (_zz_4814[31:0]         ), //i
    .dout    (fixTo_2573_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_2574 (
    .din     (_zz_4815[31:0]         ), //i
    .dout    (fixTo_2574_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_2575 (
    .din     (_zz_4816[31:0]         ), //i
    .dout    (fixTo_2575_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_2576 (
    .din     (_zz_4817[31:0]         ), //i
    .dout    (fixTo_2576_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_2577 (
    .din     (_zz_4818[31:0]         ), //i
    .dout    (fixTo_2577_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_2578 (
    .din     (_zz_4819[31:0]         ), //i
    .dout    (fixTo_2578_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_2579 (
    .din     (_zz_4820[31:0]         ), //i
    .dout    (fixTo_2579_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_2580 (
    .din     (_zz_4821[31:0]         ), //i
    .dout    (fixTo_2580_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_2581 (
    .din     (_zz_4822[31:0]         ), //i
    .dout    (fixTo_2581_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_2582 (
    .din     (_zz_4823[31:0]         ), //i
    .dout    (fixTo_2582_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_2583 (
    .din     (_zz_4824[31:0]         ), //i
    .dout    (fixTo_2583_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_2584 (
    .din     (_zz_4825[31:0]         ), //i
    .dout    (fixTo_2584_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_2585 (
    .din     (_zz_4826[31:0]         ), //i
    .dout    (fixTo_2585_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_2586 (
    .din     (_zz_4827[31:0]         ), //i
    .dout    (fixTo_2586_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_2587 (
    .din     (_zz_4828[31:0]         ), //i
    .dout    (fixTo_2587_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_2588 (
    .din     (_zz_4829[31:0]         ), //i
    .dout    (fixTo_2588_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_2589 (
    .din     (_zz_4830[31:0]         ), //i
    .dout    (fixTo_2589_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_2590 (
    .din     (_zz_4831[31:0]         ), //i
    .dout    (fixTo_2590_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_2591 (
    .din     (_zz_4832[31:0]         ), //i
    .dout    (fixTo_2591_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_2592 (
    .din     (_zz_4833[31:0]         ), //i
    .dout    (fixTo_2592_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_2593 (
    .din     (_zz_4834[31:0]         ), //i
    .dout    (fixTo_2593_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_2594 (
    .din     (_zz_4835[31:0]         ), //i
    .dout    (fixTo_2594_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_2595 (
    .din     (_zz_4836[31:0]         ), //i
    .dout    (fixTo_2595_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_2596 (
    .din     (_zz_4837[31:0]         ), //i
    .dout    (fixTo_2596_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_2597 (
    .din     (_zz_4838[31:0]         ), //i
    .dout    (fixTo_2597_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_2598 (
    .din     (_zz_4839[31:0]         ), //i
    .dout    (fixTo_2598_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_2599 (
    .din     (_zz_4840[31:0]         ), //i
    .dout    (fixTo_2599_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_2600 (
    .din     (_zz_4841[31:0]         ), //i
    .dout    (fixTo_2600_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_2601 (
    .din     (_zz_4842[31:0]         ), //i
    .dout    (fixTo_2601_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_2602 (
    .din     (_zz_4843[31:0]         ), //i
    .dout    (fixTo_2602_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_2603 (
    .din     (_zz_4844[31:0]         ), //i
    .dout    (fixTo_2603_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_2604 (
    .din     (_zz_4845[31:0]         ), //i
    .dout    (fixTo_2604_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_2605 (
    .din     (_zz_4846[31:0]         ), //i
    .dout    (fixTo_2605_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_2606 (
    .din     (_zz_4847[31:0]         ), //i
    .dout    (fixTo_2606_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_2607 (
    .din     (_zz_4848[31:0]         ), //i
    .dout    (fixTo_2607_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_2608 (
    .din     (_zz_4849[31:0]         ), //i
    .dout    (fixTo_2608_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_2609 (
    .din     (_zz_4850[31:0]         ), //i
    .dout    (fixTo_2609_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_2610 (
    .din     (_zz_4851[31:0]         ), //i
    .dout    (fixTo_2610_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_2611 (
    .din     (_zz_4852[31:0]         ), //i
    .dout    (fixTo_2611_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_2612 (
    .din     (_zz_4853[31:0]         ), //i
    .dout    (fixTo_2612_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_2613 (
    .din     (_zz_4854[31:0]         ), //i
    .dout    (fixTo_2613_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_2614 (
    .din     (_zz_4855[31:0]         ), //i
    .dout    (fixTo_2614_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_2615 (
    .din     (_zz_4856[31:0]         ), //i
    .dout    (fixTo_2615_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_2616 (
    .din     (_zz_4857[31:0]         ), //i
    .dout    (fixTo_2616_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_2617 (
    .din     (_zz_4858[31:0]         ), //i
    .dout    (fixTo_2617_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_2618 (
    .din     (_zz_4859[31:0]         ), //i
    .dout    (fixTo_2618_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_2619 (
    .din     (_zz_4860[31:0]         ), //i
    .dout    (fixTo_2619_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_2620 (
    .din     (_zz_4861[31:0]         ), //i
    .dout    (fixTo_2620_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_2621 (
    .din     (_zz_4862[31:0]         ), //i
    .dout    (fixTo_2621_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_2622 (
    .din     (_zz_4863[31:0]         ), //i
    .dout    (fixTo_2622_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_2623 (
    .din     (_zz_4864[31:0]         ), //i
    .dout    (fixTo_2623_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_2624 (
    .din     (_zz_4865[31:0]         ), //i
    .dout    (fixTo_2624_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_2625 (
    .din     (_zz_4866[31:0]         ), //i
    .dout    (fixTo_2625_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_2626 (
    .din     (_zz_4867[31:0]         ), //i
    .dout    (fixTo_2626_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_2627 (
    .din     (_zz_4868[31:0]         ), //i
    .dout    (fixTo_2627_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_2628 (
    .din     (_zz_4869[31:0]         ), //i
    .dout    (fixTo_2628_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_2629 (
    .din     (_zz_4870[31:0]         ), //i
    .dout    (fixTo_2629_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_2630 (
    .din     (_zz_4871[31:0]         ), //i
    .dout    (fixTo_2630_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_2631 (
    .din     (_zz_4872[31:0]         ), //i
    .dout    (fixTo_2631_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_2632 (
    .din     (_zz_4873[31:0]         ), //i
    .dout    (fixTo_2632_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_2633 (
    .din     (_zz_4874[31:0]         ), //i
    .dout    (fixTo_2633_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_2634 (
    .din     (_zz_4875[31:0]         ), //i
    .dout    (fixTo_2634_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_2635 (
    .din     (_zz_4876[31:0]         ), //i
    .dout    (fixTo_2635_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_2636 (
    .din     (_zz_4877[31:0]         ), //i
    .dout    (fixTo_2636_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_2637 (
    .din     (_zz_4878[31:0]         ), //i
    .dout    (fixTo_2637_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_2638 (
    .din     (_zz_4879[31:0]         ), //i
    .dout    (fixTo_2638_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_2639 (
    .din     (_zz_4880[31:0]         ), //i
    .dout    (fixTo_2639_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_2640 (
    .din     (_zz_4881[31:0]         ), //i
    .dout    (fixTo_2640_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_2641 (
    .din     (_zz_4882[31:0]         ), //i
    .dout    (fixTo_2641_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_2642 (
    .din     (_zz_4883[31:0]         ), //i
    .dout    (fixTo_2642_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_2643 (
    .din     (_zz_4884[31:0]         ), //i
    .dout    (fixTo_2643_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_2644 (
    .din     (_zz_4885[31:0]         ), //i
    .dout    (fixTo_2644_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_2645 (
    .din     (_zz_4886[31:0]         ), //i
    .dout    (fixTo_2645_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_2646 (
    .din     (_zz_4887[31:0]         ), //i
    .dout    (fixTo_2646_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_2647 (
    .din     (_zz_4888[31:0]         ), //i
    .dout    (fixTo_2647_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_2648 (
    .din     (_zz_4889[31:0]         ), //i
    .dout    (fixTo_2648_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_2649 (
    .din     (_zz_4890[31:0]         ), //i
    .dout    (fixTo_2649_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_2650 (
    .din     (_zz_4891[31:0]         ), //i
    .dout    (fixTo_2650_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_2651 (
    .din     (_zz_4892[31:0]         ), //i
    .dout    (fixTo_2651_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_2652 (
    .din     (_zz_4893[31:0]         ), //i
    .dout    (fixTo_2652_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_2653 (
    .din     (_zz_4894[31:0]         ), //i
    .dout    (fixTo_2653_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_2654 (
    .din     (_zz_4895[31:0]         ), //i
    .dout    (fixTo_2654_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_2655 (
    .din     (_zz_4896[31:0]         ), //i
    .dout    (fixTo_2655_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_2656 (
    .din     (_zz_4897[31:0]         ), //i
    .dout    (fixTo_2656_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_2657 (
    .din     (_zz_4898[31:0]         ), //i
    .dout    (fixTo_2657_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_2658 (
    .din     (_zz_4899[31:0]         ), //i
    .dout    (fixTo_2658_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_2659 (
    .din     (_zz_4900[31:0]         ), //i
    .dout    (fixTo_2659_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_2660 (
    .din     (_zz_4901[31:0]         ), //i
    .dout    (fixTo_2660_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_2661 (
    .din     (_zz_4902[31:0]         ), //i
    .dout    (fixTo_2661_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_2662 (
    .din     (_zz_4903[31:0]         ), //i
    .dout    (fixTo_2662_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_2663 (
    .din     (_zz_4904[31:0]         ), //i
    .dout    (fixTo_2663_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_2664 (
    .din     (_zz_4905[31:0]         ), //i
    .dout    (fixTo_2664_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_2665 (
    .din     (_zz_4906[31:0]         ), //i
    .dout    (fixTo_2665_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_2666 (
    .din     (_zz_4907[31:0]         ), //i
    .dout    (fixTo_2666_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_2667 (
    .din     (_zz_4908[31:0]         ), //i
    .dout    (fixTo_2667_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_2668 (
    .din     (_zz_4909[31:0]         ), //i
    .dout    (fixTo_2668_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_2669 (
    .din     (_zz_4910[31:0]         ), //i
    .dout    (fixTo_2669_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_2670 (
    .din     (_zz_4911[31:0]         ), //i
    .dout    (fixTo_2670_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_2671 (
    .din     (_zz_4912[31:0]         ), //i
    .dout    (fixTo_2671_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_2672 (
    .din     (_zz_4913[31:0]         ), //i
    .dout    (fixTo_2672_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_2673 (
    .din     (_zz_4914[31:0]         ), //i
    .dout    (fixTo_2673_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_2674 (
    .din     (_zz_4915[31:0]         ), //i
    .dout    (fixTo_2674_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_2675 (
    .din     (_zz_4916[31:0]         ), //i
    .dout    (fixTo_2675_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_2676 (
    .din     (_zz_4917[31:0]         ), //i
    .dout    (fixTo_2676_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_2677 (
    .din     (_zz_4918[31:0]         ), //i
    .dout    (fixTo_2677_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_2678 (
    .din     (_zz_4919[31:0]         ), //i
    .dout    (fixTo_2678_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_2679 (
    .din     (_zz_4920[31:0]         ), //i
    .dout    (fixTo_2679_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_2680 (
    .din     (_zz_4921[31:0]         ), //i
    .dout    (fixTo_2680_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_2681 (
    .din     (_zz_4922[31:0]         ), //i
    .dout    (fixTo_2681_dout[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_2682 (
    .din     (_zz_4923[31:0]         ), //i
    .dout    (fixTo_2682_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_2683 (
    .din     (_zz_4924[31:0]         ), //i
    .dout    (fixTo_2683_dout[31:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_2684 (
    .din     (_zz_4925[31:0]         ), //i
    .dout    (fixTo_2684_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_2685 (
    .din     (_zz_4926[31:0]         ), //i
    .dout    (fixTo_2685_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_2686 (
    .din     (_zz_4927[31:0]         ), //i
    .dout    (fixTo_2686_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_2687 (
    .din     (_zz_4928[31:0]         ), //i
    .dout    (fixTo_2687_dout[15:0]  )  //o
  );
  assign twiddle_factor_table_0_real = 16'h0100;
  assign twiddle_factor_table_0_imag = 16'h0;
  assign twiddle_factor_table_1_real = 16'h0100;
  assign twiddle_factor_table_1_imag = 16'h0;
  assign twiddle_factor_table_2_real = 16'h0;
  assign twiddle_factor_table_2_imag = 16'hff00;
  assign twiddle_factor_table_3_real = 16'h0100;
  assign twiddle_factor_table_3_imag = 16'h0;
  assign twiddle_factor_table_4_real = 16'h00b5;
  assign twiddle_factor_table_4_imag = 16'hff4b;
  assign twiddle_factor_table_5_real = 16'h0;
  assign twiddle_factor_table_5_imag = 16'hff00;
  assign twiddle_factor_table_6_real = 16'hff4b;
  assign twiddle_factor_table_6_imag = 16'hff4b;
  assign twiddle_factor_table_7_real = 16'h0100;
  assign twiddle_factor_table_7_imag = 16'h0;
  assign twiddle_factor_table_8_real = 16'h00ec;
  assign twiddle_factor_table_8_imag = 16'hff9f;
  assign twiddle_factor_table_9_real = 16'h00b5;
  assign twiddle_factor_table_9_imag = 16'hff4b;
  assign twiddle_factor_table_10_real = 16'h0061;
  assign twiddle_factor_table_10_imag = 16'hff14;
  assign twiddle_factor_table_11_real = 16'h0;
  assign twiddle_factor_table_11_imag = 16'hff00;
  assign twiddle_factor_table_12_real = 16'hff9f;
  assign twiddle_factor_table_12_imag = 16'hff14;
  assign twiddle_factor_table_13_real = 16'hff4b;
  assign twiddle_factor_table_13_imag = 16'hff4b;
  assign twiddle_factor_table_14_real = 16'hff14;
  assign twiddle_factor_table_14_imag = 16'hff9f;
  assign twiddle_factor_table_15_real = 16'h0100;
  assign twiddle_factor_table_15_imag = 16'h0;
  assign twiddle_factor_table_16_real = 16'h00fb;
  assign twiddle_factor_table_16_imag = 16'hffcf;
  assign twiddle_factor_table_17_real = 16'h00ec;
  assign twiddle_factor_table_17_imag = 16'hff9f;
  assign twiddle_factor_table_18_real = 16'h00d4;
  assign twiddle_factor_table_18_imag = 16'hff72;
  assign twiddle_factor_table_19_real = 16'h00b5;
  assign twiddle_factor_table_19_imag = 16'hff4b;
  assign twiddle_factor_table_20_real = 16'h008e;
  assign twiddle_factor_table_20_imag = 16'hff2c;
  assign twiddle_factor_table_21_real = 16'h0061;
  assign twiddle_factor_table_21_imag = 16'hff14;
  assign twiddle_factor_table_22_real = 16'h0031;
  assign twiddle_factor_table_22_imag = 16'hff05;
  assign twiddle_factor_table_23_real = 16'h0;
  assign twiddle_factor_table_23_imag = 16'hff00;
  assign twiddle_factor_table_24_real = 16'hffcf;
  assign twiddle_factor_table_24_imag = 16'hff05;
  assign twiddle_factor_table_25_real = 16'hff9f;
  assign twiddle_factor_table_25_imag = 16'hff14;
  assign twiddle_factor_table_26_real = 16'hff72;
  assign twiddle_factor_table_26_imag = 16'hff2c;
  assign twiddle_factor_table_27_real = 16'hff4b;
  assign twiddle_factor_table_27_imag = 16'hff4b;
  assign twiddle_factor_table_28_real = 16'hff2c;
  assign twiddle_factor_table_28_imag = 16'hff72;
  assign twiddle_factor_table_29_real = 16'hff14;
  assign twiddle_factor_table_29_imag = 16'hff9f;
  assign twiddle_factor_table_30_real = 16'hff05;
  assign twiddle_factor_table_30_imag = 16'hffcf;
  assign twiddle_factor_table_31_real = 16'h0100;
  assign twiddle_factor_table_31_imag = 16'h0;
  assign twiddle_factor_table_32_real = 16'h00fe;
  assign twiddle_factor_table_32_imag = 16'hffe7;
  assign twiddle_factor_table_33_real = 16'h00fb;
  assign twiddle_factor_table_33_imag = 16'hffcf;
  assign twiddle_factor_table_34_real = 16'h00f4;
  assign twiddle_factor_table_34_imag = 16'hffb6;
  assign twiddle_factor_table_35_real = 16'h00ec;
  assign twiddle_factor_table_35_imag = 16'hff9f;
  assign twiddle_factor_table_36_real = 16'h00e1;
  assign twiddle_factor_table_36_imag = 16'hff88;
  assign twiddle_factor_table_37_real = 16'h00d4;
  assign twiddle_factor_table_37_imag = 16'hff72;
  assign twiddle_factor_table_38_real = 16'h00c5;
  assign twiddle_factor_table_38_imag = 16'hff5e;
  assign twiddle_factor_table_39_real = 16'h00b5;
  assign twiddle_factor_table_39_imag = 16'hff4b;
  assign twiddle_factor_table_40_real = 16'h00a2;
  assign twiddle_factor_table_40_imag = 16'hff3b;
  assign twiddle_factor_table_41_real = 16'h008e;
  assign twiddle_factor_table_41_imag = 16'hff2c;
  assign twiddle_factor_table_42_real = 16'h0078;
  assign twiddle_factor_table_42_imag = 16'hff1f;
  assign twiddle_factor_table_43_real = 16'h0061;
  assign twiddle_factor_table_43_imag = 16'hff14;
  assign twiddle_factor_table_44_real = 16'h004a;
  assign twiddle_factor_table_44_imag = 16'hff0c;
  assign twiddle_factor_table_45_real = 16'h0031;
  assign twiddle_factor_table_45_imag = 16'hff05;
  assign twiddle_factor_table_46_real = 16'h0019;
  assign twiddle_factor_table_46_imag = 16'hff02;
  assign twiddle_factor_table_47_real = 16'h0;
  assign twiddle_factor_table_47_imag = 16'hff00;
  assign twiddle_factor_table_48_real = 16'hffe7;
  assign twiddle_factor_table_48_imag = 16'hff02;
  assign twiddle_factor_table_49_real = 16'hffcf;
  assign twiddle_factor_table_49_imag = 16'hff05;
  assign twiddle_factor_table_50_real = 16'hffb6;
  assign twiddle_factor_table_50_imag = 16'hff0c;
  assign twiddle_factor_table_51_real = 16'hff9f;
  assign twiddle_factor_table_51_imag = 16'hff14;
  assign twiddle_factor_table_52_real = 16'hff88;
  assign twiddle_factor_table_52_imag = 16'hff1f;
  assign twiddle_factor_table_53_real = 16'hff72;
  assign twiddle_factor_table_53_imag = 16'hff2c;
  assign twiddle_factor_table_54_real = 16'hff5e;
  assign twiddle_factor_table_54_imag = 16'hff3b;
  assign twiddle_factor_table_55_real = 16'hff4b;
  assign twiddle_factor_table_55_imag = 16'hff4b;
  assign twiddle_factor_table_56_real = 16'hff3b;
  assign twiddle_factor_table_56_imag = 16'hff5e;
  assign twiddle_factor_table_57_real = 16'hff2c;
  assign twiddle_factor_table_57_imag = 16'hff72;
  assign twiddle_factor_table_58_real = 16'hff1f;
  assign twiddle_factor_table_58_imag = 16'hff88;
  assign twiddle_factor_table_59_real = 16'hff14;
  assign twiddle_factor_table_59_imag = 16'hff9f;
  assign twiddle_factor_table_60_real = 16'hff0c;
  assign twiddle_factor_table_60_imag = 16'hffb6;
  assign twiddle_factor_table_61_real = 16'hff05;
  assign twiddle_factor_table_61_imag = 16'hffcf;
  assign twiddle_factor_table_62_real = 16'hff02;
  assign twiddle_factor_table_62_imag = 16'hffe7;
  assign twiddle_factor_table_63_real = 16'h0100;
  assign twiddle_factor_table_63_imag = 16'h0;
  assign twiddle_factor_table_64_real = 16'h00ff;
  assign twiddle_factor_table_64_imag = 16'hfff4;
  assign twiddle_factor_table_65_real = 16'h00fe;
  assign twiddle_factor_table_65_imag = 16'hffe7;
  assign twiddle_factor_table_66_real = 16'h00fd;
  assign twiddle_factor_table_66_imag = 16'hffdb;
  assign twiddle_factor_table_67_real = 16'h00fb;
  assign twiddle_factor_table_67_imag = 16'hffcf;
  assign twiddle_factor_table_68_real = 16'h00f8;
  assign twiddle_factor_table_68_imag = 16'hffc2;
  assign twiddle_factor_table_69_real = 16'h00f4;
  assign twiddle_factor_table_69_imag = 16'hffb6;
  assign twiddle_factor_table_70_real = 16'h00f1;
  assign twiddle_factor_table_70_imag = 16'hffaa;
  assign twiddle_factor_table_71_real = 16'h00ec;
  assign twiddle_factor_table_71_imag = 16'hff9f;
  assign twiddle_factor_table_72_real = 16'h00e7;
  assign twiddle_factor_table_72_imag = 16'hff93;
  assign twiddle_factor_table_73_real = 16'h00e1;
  assign twiddle_factor_table_73_imag = 16'hff88;
  assign twiddle_factor_table_74_real = 16'h00db;
  assign twiddle_factor_table_74_imag = 16'hff7d;
  assign twiddle_factor_table_75_real = 16'h00d4;
  assign twiddle_factor_table_75_imag = 16'hff72;
  assign twiddle_factor_table_76_real = 16'h00cd;
  assign twiddle_factor_table_76_imag = 16'hff68;
  assign twiddle_factor_table_77_real = 16'h00c5;
  assign twiddle_factor_table_77_imag = 16'hff5e;
  assign twiddle_factor_table_78_real = 16'h00bd;
  assign twiddle_factor_table_78_imag = 16'hff55;
  assign twiddle_factor_table_79_real = 16'h00b5;
  assign twiddle_factor_table_79_imag = 16'hff4b;
  assign twiddle_factor_table_80_real = 16'h00ab;
  assign twiddle_factor_table_80_imag = 16'hff43;
  assign twiddle_factor_table_81_real = 16'h00a2;
  assign twiddle_factor_table_81_imag = 16'hff3b;
  assign twiddle_factor_table_82_real = 16'h0098;
  assign twiddle_factor_table_82_imag = 16'hff33;
  assign twiddle_factor_table_83_real = 16'h008e;
  assign twiddle_factor_table_83_imag = 16'hff2c;
  assign twiddle_factor_table_84_real = 16'h0083;
  assign twiddle_factor_table_84_imag = 16'hff25;
  assign twiddle_factor_table_85_real = 16'h0078;
  assign twiddle_factor_table_85_imag = 16'hff1f;
  assign twiddle_factor_table_86_real = 16'h006d;
  assign twiddle_factor_table_86_imag = 16'hff19;
  assign twiddle_factor_table_87_real = 16'h0061;
  assign twiddle_factor_table_87_imag = 16'hff14;
  assign twiddle_factor_table_88_real = 16'h0056;
  assign twiddle_factor_table_88_imag = 16'hff0f;
  assign twiddle_factor_table_89_real = 16'h004a;
  assign twiddle_factor_table_89_imag = 16'hff0c;
  assign twiddle_factor_table_90_real = 16'h003e;
  assign twiddle_factor_table_90_imag = 16'hff08;
  assign twiddle_factor_table_91_real = 16'h0031;
  assign twiddle_factor_table_91_imag = 16'hff05;
  assign twiddle_factor_table_92_real = 16'h0025;
  assign twiddle_factor_table_92_imag = 16'hff03;
  assign twiddle_factor_table_93_real = 16'h0019;
  assign twiddle_factor_table_93_imag = 16'hff02;
  assign twiddle_factor_table_94_real = 16'h000c;
  assign twiddle_factor_table_94_imag = 16'hff01;
  assign twiddle_factor_table_95_real = 16'h0;
  assign twiddle_factor_table_95_imag = 16'hff00;
  assign twiddle_factor_table_96_real = 16'hfff4;
  assign twiddle_factor_table_96_imag = 16'hff01;
  assign twiddle_factor_table_97_real = 16'hffe7;
  assign twiddle_factor_table_97_imag = 16'hff02;
  assign twiddle_factor_table_98_real = 16'hffdb;
  assign twiddle_factor_table_98_imag = 16'hff03;
  assign twiddle_factor_table_99_real = 16'hffcf;
  assign twiddle_factor_table_99_imag = 16'hff05;
  assign twiddle_factor_table_100_real = 16'hffc2;
  assign twiddle_factor_table_100_imag = 16'hff08;
  assign twiddle_factor_table_101_real = 16'hffb6;
  assign twiddle_factor_table_101_imag = 16'hff0c;
  assign twiddle_factor_table_102_real = 16'hffaa;
  assign twiddle_factor_table_102_imag = 16'hff0f;
  assign twiddle_factor_table_103_real = 16'hff9f;
  assign twiddle_factor_table_103_imag = 16'hff14;
  assign twiddle_factor_table_104_real = 16'hff93;
  assign twiddle_factor_table_104_imag = 16'hff19;
  assign twiddle_factor_table_105_real = 16'hff88;
  assign twiddle_factor_table_105_imag = 16'hff1f;
  assign twiddle_factor_table_106_real = 16'hff7d;
  assign twiddle_factor_table_106_imag = 16'hff25;
  assign twiddle_factor_table_107_real = 16'hff72;
  assign twiddle_factor_table_107_imag = 16'hff2c;
  assign twiddle_factor_table_108_real = 16'hff68;
  assign twiddle_factor_table_108_imag = 16'hff33;
  assign twiddle_factor_table_109_real = 16'hff5e;
  assign twiddle_factor_table_109_imag = 16'hff3b;
  assign twiddle_factor_table_110_real = 16'hff55;
  assign twiddle_factor_table_110_imag = 16'hff43;
  assign twiddle_factor_table_111_real = 16'hff4b;
  assign twiddle_factor_table_111_imag = 16'hff4b;
  assign twiddle_factor_table_112_real = 16'hff43;
  assign twiddle_factor_table_112_imag = 16'hff55;
  assign twiddle_factor_table_113_real = 16'hff3b;
  assign twiddle_factor_table_113_imag = 16'hff5e;
  assign twiddle_factor_table_114_real = 16'hff33;
  assign twiddle_factor_table_114_imag = 16'hff68;
  assign twiddle_factor_table_115_real = 16'hff2c;
  assign twiddle_factor_table_115_imag = 16'hff72;
  assign twiddle_factor_table_116_real = 16'hff25;
  assign twiddle_factor_table_116_imag = 16'hff7d;
  assign twiddle_factor_table_117_real = 16'hff1f;
  assign twiddle_factor_table_117_imag = 16'hff88;
  assign twiddle_factor_table_118_real = 16'hff19;
  assign twiddle_factor_table_118_imag = 16'hff93;
  assign twiddle_factor_table_119_real = 16'hff14;
  assign twiddle_factor_table_119_imag = 16'hff9f;
  assign twiddle_factor_table_120_real = 16'hff0f;
  assign twiddle_factor_table_120_imag = 16'hffaa;
  assign twiddle_factor_table_121_real = 16'hff0c;
  assign twiddle_factor_table_121_imag = 16'hffb6;
  assign twiddle_factor_table_122_real = 16'hff08;
  assign twiddle_factor_table_122_imag = 16'hffc2;
  assign twiddle_factor_table_123_real = 16'hff05;
  assign twiddle_factor_table_123_imag = 16'hffcf;
  assign twiddle_factor_table_124_real = 16'hff03;
  assign twiddle_factor_table_124_imag = 16'hffdb;
  assign twiddle_factor_table_125_real = 16'hff02;
  assign twiddle_factor_table_125_imag = 16'hffe7;
  assign twiddle_factor_table_126_real = 16'hff01;
  assign twiddle_factor_table_126_imag = 16'hfff4;
  assign data_reorder_0_real = data_in_0_real;
  assign data_reorder_0_imag = data_in_0_imag;
  assign data_reorder_64_real = data_in_1_real;
  assign data_reorder_64_imag = data_in_1_imag;
  assign data_reorder_32_real = data_in_2_real;
  assign data_reorder_32_imag = data_in_2_imag;
  assign data_reorder_96_real = data_in_3_real;
  assign data_reorder_96_imag = data_in_3_imag;
  assign data_reorder_16_real = data_in_4_real;
  assign data_reorder_16_imag = data_in_4_imag;
  assign data_reorder_80_real = data_in_5_real;
  assign data_reorder_80_imag = data_in_5_imag;
  assign data_reorder_48_real = data_in_6_real;
  assign data_reorder_48_imag = data_in_6_imag;
  assign data_reorder_112_real = data_in_7_real;
  assign data_reorder_112_imag = data_in_7_imag;
  assign data_reorder_8_real = data_in_8_real;
  assign data_reorder_8_imag = data_in_8_imag;
  assign data_reorder_72_real = data_in_9_real;
  assign data_reorder_72_imag = data_in_9_imag;
  assign data_reorder_40_real = data_in_10_real;
  assign data_reorder_40_imag = data_in_10_imag;
  assign data_reorder_104_real = data_in_11_real;
  assign data_reorder_104_imag = data_in_11_imag;
  assign data_reorder_24_real = data_in_12_real;
  assign data_reorder_24_imag = data_in_12_imag;
  assign data_reorder_88_real = data_in_13_real;
  assign data_reorder_88_imag = data_in_13_imag;
  assign data_reorder_56_real = data_in_14_real;
  assign data_reorder_56_imag = data_in_14_imag;
  assign data_reorder_120_real = data_in_15_real;
  assign data_reorder_120_imag = data_in_15_imag;
  assign data_reorder_4_real = data_in_16_real;
  assign data_reorder_4_imag = data_in_16_imag;
  assign data_reorder_68_real = data_in_17_real;
  assign data_reorder_68_imag = data_in_17_imag;
  assign data_reorder_36_real = data_in_18_real;
  assign data_reorder_36_imag = data_in_18_imag;
  assign data_reorder_100_real = data_in_19_real;
  assign data_reorder_100_imag = data_in_19_imag;
  assign data_reorder_20_real = data_in_20_real;
  assign data_reorder_20_imag = data_in_20_imag;
  assign data_reorder_84_real = data_in_21_real;
  assign data_reorder_84_imag = data_in_21_imag;
  assign data_reorder_52_real = data_in_22_real;
  assign data_reorder_52_imag = data_in_22_imag;
  assign data_reorder_116_real = data_in_23_real;
  assign data_reorder_116_imag = data_in_23_imag;
  assign data_reorder_12_real = data_in_24_real;
  assign data_reorder_12_imag = data_in_24_imag;
  assign data_reorder_76_real = data_in_25_real;
  assign data_reorder_76_imag = data_in_25_imag;
  assign data_reorder_44_real = data_in_26_real;
  assign data_reorder_44_imag = data_in_26_imag;
  assign data_reorder_108_real = data_in_27_real;
  assign data_reorder_108_imag = data_in_27_imag;
  assign data_reorder_28_real = data_in_28_real;
  assign data_reorder_28_imag = data_in_28_imag;
  assign data_reorder_92_real = data_in_29_real;
  assign data_reorder_92_imag = data_in_29_imag;
  assign data_reorder_60_real = data_in_30_real;
  assign data_reorder_60_imag = data_in_30_imag;
  assign data_reorder_124_real = data_in_31_real;
  assign data_reorder_124_imag = data_in_31_imag;
  assign data_reorder_2_real = data_in_32_real;
  assign data_reorder_2_imag = data_in_32_imag;
  assign data_reorder_66_real = data_in_33_real;
  assign data_reorder_66_imag = data_in_33_imag;
  assign data_reorder_34_real = data_in_34_real;
  assign data_reorder_34_imag = data_in_34_imag;
  assign data_reorder_98_real = data_in_35_real;
  assign data_reorder_98_imag = data_in_35_imag;
  assign data_reorder_18_real = data_in_36_real;
  assign data_reorder_18_imag = data_in_36_imag;
  assign data_reorder_82_real = data_in_37_real;
  assign data_reorder_82_imag = data_in_37_imag;
  assign data_reorder_50_real = data_in_38_real;
  assign data_reorder_50_imag = data_in_38_imag;
  assign data_reorder_114_real = data_in_39_real;
  assign data_reorder_114_imag = data_in_39_imag;
  assign data_reorder_10_real = data_in_40_real;
  assign data_reorder_10_imag = data_in_40_imag;
  assign data_reorder_74_real = data_in_41_real;
  assign data_reorder_74_imag = data_in_41_imag;
  assign data_reorder_42_real = data_in_42_real;
  assign data_reorder_42_imag = data_in_42_imag;
  assign data_reorder_106_real = data_in_43_real;
  assign data_reorder_106_imag = data_in_43_imag;
  assign data_reorder_26_real = data_in_44_real;
  assign data_reorder_26_imag = data_in_44_imag;
  assign data_reorder_90_real = data_in_45_real;
  assign data_reorder_90_imag = data_in_45_imag;
  assign data_reorder_58_real = data_in_46_real;
  assign data_reorder_58_imag = data_in_46_imag;
  assign data_reorder_122_real = data_in_47_real;
  assign data_reorder_122_imag = data_in_47_imag;
  assign data_reorder_6_real = data_in_48_real;
  assign data_reorder_6_imag = data_in_48_imag;
  assign data_reorder_70_real = data_in_49_real;
  assign data_reorder_70_imag = data_in_49_imag;
  assign data_reorder_38_real = data_in_50_real;
  assign data_reorder_38_imag = data_in_50_imag;
  assign data_reorder_102_real = data_in_51_real;
  assign data_reorder_102_imag = data_in_51_imag;
  assign data_reorder_22_real = data_in_52_real;
  assign data_reorder_22_imag = data_in_52_imag;
  assign data_reorder_86_real = data_in_53_real;
  assign data_reorder_86_imag = data_in_53_imag;
  assign data_reorder_54_real = data_in_54_real;
  assign data_reorder_54_imag = data_in_54_imag;
  assign data_reorder_118_real = data_in_55_real;
  assign data_reorder_118_imag = data_in_55_imag;
  assign data_reorder_14_real = data_in_56_real;
  assign data_reorder_14_imag = data_in_56_imag;
  assign data_reorder_78_real = data_in_57_real;
  assign data_reorder_78_imag = data_in_57_imag;
  assign data_reorder_46_real = data_in_58_real;
  assign data_reorder_46_imag = data_in_58_imag;
  assign data_reorder_110_real = data_in_59_real;
  assign data_reorder_110_imag = data_in_59_imag;
  assign data_reorder_30_real = data_in_60_real;
  assign data_reorder_30_imag = data_in_60_imag;
  assign data_reorder_94_real = data_in_61_real;
  assign data_reorder_94_imag = data_in_61_imag;
  assign data_reorder_62_real = data_in_62_real;
  assign data_reorder_62_imag = data_in_62_imag;
  assign data_reorder_126_real = data_in_63_real;
  assign data_reorder_126_imag = data_in_63_imag;
  assign data_reorder_1_real = data_in_64_real;
  assign data_reorder_1_imag = data_in_64_imag;
  assign data_reorder_65_real = data_in_65_real;
  assign data_reorder_65_imag = data_in_65_imag;
  assign data_reorder_33_real = data_in_66_real;
  assign data_reorder_33_imag = data_in_66_imag;
  assign data_reorder_97_real = data_in_67_real;
  assign data_reorder_97_imag = data_in_67_imag;
  assign data_reorder_17_real = data_in_68_real;
  assign data_reorder_17_imag = data_in_68_imag;
  assign data_reorder_81_real = data_in_69_real;
  assign data_reorder_81_imag = data_in_69_imag;
  assign data_reorder_49_real = data_in_70_real;
  assign data_reorder_49_imag = data_in_70_imag;
  assign data_reorder_113_real = data_in_71_real;
  assign data_reorder_113_imag = data_in_71_imag;
  assign data_reorder_9_real = data_in_72_real;
  assign data_reorder_9_imag = data_in_72_imag;
  assign data_reorder_73_real = data_in_73_real;
  assign data_reorder_73_imag = data_in_73_imag;
  assign data_reorder_41_real = data_in_74_real;
  assign data_reorder_41_imag = data_in_74_imag;
  assign data_reorder_105_real = data_in_75_real;
  assign data_reorder_105_imag = data_in_75_imag;
  assign data_reorder_25_real = data_in_76_real;
  assign data_reorder_25_imag = data_in_76_imag;
  assign data_reorder_89_real = data_in_77_real;
  assign data_reorder_89_imag = data_in_77_imag;
  assign data_reorder_57_real = data_in_78_real;
  assign data_reorder_57_imag = data_in_78_imag;
  assign data_reorder_121_real = data_in_79_real;
  assign data_reorder_121_imag = data_in_79_imag;
  assign data_reorder_5_real = data_in_80_real;
  assign data_reorder_5_imag = data_in_80_imag;
  assign data_reorder_69_real = data_in_81_real;
  assign data_reorder_69_imag = data_in_81_imag;
  assign data_reorder_37_real = data_in_82_real;
  assign data_reorder_37_imag = data_in_82_imag;
  assign data_reorder_101_real = data_in_83_real;
  assign data_reorder_101_imag = data_in_83_imag;
  assign data_reorder_21_real = data_in_84_real;
  assign data_reorder_21_imag = data_in_84_imag;
  assign data_reorder_85_real = data_in_85_real;
  assign data_reorder_85_imag = data_in_85_imag;
  assign data_reorder_53_real = data_in_86_real;
  assign data_reorder_53_imag = data_in_86_imag;
  assign data_reorder_117_real = data_in_87_real;
  assign data_reorder_117_imag = data_in_87_imag;
  assign data_reorder_13_real = data_in_88_real;
  assign data_reorder_13_imag = data_in_88_imag;
  assign data_reorder_77_real = data_in_89_real;
  assign data_reorder_77_imag = data_in_89_imag;
  assign data_reorder_45_real = data_in_90_real;
  assign data_reorder_45_imag = data_in_90_imag;
  assign data_reorder_109_real = data_in_91_real;
  assign data_reorder_109_imag = data_in_91_imag;
  assign data_reorder_29_real = data_in_92_real;
  assign data_reorder_29_imag = data_in_92_imag;
  assign data_reorder_93_real = data_in_93_real;
  assign data_reorder_93_imag = data_in_93_imag;
  assign data_reorder_61_real = data_in_94_real;
  assign data_reorder_61_imag = data_in_94_imag;
  assign data_reorder_125_real = data_in_95_real;
  assign data_reorder_125_imag = data_in_95_imag;
  assign data_reorder_3_real = data_in_96_real;
  assign data_reorder_3_imag = data_in_96_imag;
  assign data_reorder_67_real = data_in_97_real;
  assign data_reorder_67_imag = data_in_97_imag;
  assign data_reorder_35_real = data_in_98_real;
  assign data_reorder_35_imag = data_in_98_imag;
  assign data_reorder_99_real = data_in_99_real;
  assign data_reorder_99_imag = data_in_99_imag;
  assign data_reorder_19_real = data_in_100_real;
  assign data_reorder_19_imag = data_in_100_imag;
  assign data_reorder_83_real = data_in_101_real;
  assign data_reorder_83_imag = data_in_101_imag;
  assign data_reorder_51_real = data_in_102_real;
  assign data_reorder_51_imag = data_in_102_imag;
  assign data_reorder_115_real = data_in_103_real;
  assign data_reorder_115_imag = data_in_103_imag;
  assign data_reorder_11_real = data_in_104_real;
  assign data_reorder_11_imag = data_in_104_imag;
  assign data_reorder_75_real = data_in_105_real;
  assign data_reorder_75_imag = data_in_105_imag;
  assign data_reorder_43_real = data_in_106_real;
  assign data_reorder_43_imag = data_in_106_imag;
  assign data_reorder_107_real = data_in_107_real;
  assign data_reorder_107_imag = data_in_107_imag;
  assign data_reorder_27_real = data_in_108_real;
  assign data_reorder_27_imag = data_in_108_imag;
  assign data_reorder_91_real = data_in_109_real;
  assign data_reorder_91_imag = data_in_109_imag;
  assign data_reorder_59_real = data_in_110_real;
  assign data_reorder_59_imag = data_in_110_imag;
  assign data_reorder_123_real = data_in_111_real;
  assign data_reorder_123_imag = data_in_111_imag;
  assign data_reorder_7_real = data_in_112_real;
  assign data_reorder_7_imag = data_in_112_imag;
  assign data_reorder_71_real = data_in_113_real;
  assign data_reorder_71_imag = data_in_113_imag;
  assign data_reorder_39_real = data_in_114_real;
  assign data_reorder_39_imag = data_in_114_imag;
  assign data_reorder_103_real = data_in_115_real;
  assign data_reorder_103_imag = data_in_115_imag;
  assign data_reorder_23_real = data_in_116_real;
  assign data_reorder_23_imag = data_in_116_imag;
  assign data_reorder_87_real = data_in_117_real;
  assign data_reorder_87_imag = data_in_117_imag;
  assign data_reorder_55_real = data_in_118_real;
  assign data_reorder_55_imag = data_in_118_imag;
  assign data_reorder_119_real = data_in_119_real;
  assign data_reorder_119_imag = data_in_119_imag;
  assign data_reorder_15_real = data_in_120_real;
  assign data_reorder_15_imag = data_in_120_imag;
  assign data_reorder_79_real = data_in_121_real;
  assign data_reorder_79_imag = data_in_121_imag;
  assign data_reorder_47_real = data_in_122_real;
  assign data_reorder_47_imag = data_in_122_imag;
  assign data_reorder_111_real = data_in_123_real;
  assign data_reorder_111_imag = data_in_123_imag;
  assign data_reorder_31_real = data_in_124_real;
  assign data_reorder_31_imag = data_in_124_imag;
  assign data_reorder_95_real = data_in_125_real;
  assign data_reorder_95_imag = data_in_125_imag;
  assign data_reorder_63_real = data_in_126_real;
  assign data_reorder_63_imag = data_in_126_imag;
  assign data_reorder_127_real = data_in_127_real;
  assign data_reorder_127_imag = data_in_127_imag;
  always @ (*) begin
    current_level_willIncrement = 1'b0;
    if(null_cond_period)begin
      current_level_willIncrement = 1'b1;
    end
  end

  assign current_level_willClear = 1'b0;
  assign current_level_willOverflowIfInc = (current_level_value == 3'b111);
  assign current_level_willOverflow = (current_level_willOverflowIfInc && current_level_willIncrement);
  always @ (*) begin
    current_level_valueNext = (current_level_value + _zz_4930);
    if(current_level_willClear)begin
      current_level_valueNext = 3'b000;
    end
  end

  assign null_cond_period = (io_data_in_valid_regNext || null_cond_period_minus_1);
  assign _zz_3 = ($signed(_zz_4931) * $signed(data_mid_1_real));
  assign _zz_2241 = _zz_4932;
  assign _zz_1 = _zz_4935[31 : 0];
  assign _zz_2242 = _zz_4936;
  assign _zz_2 = _zz_4939[31 : 0];
  assign _zz_4 = 1'b1;
  assign _zz_2243 = _zz_4940;
  assign _zz_2244 = _zz_4948;
  assign _zz_5 = 1'b1;
  assign _zz_2245 = _zz_4956;
  assign _zz_2246 = _zz_4964;
  assign _zz_8 = ($signed(_zz_4972) * $signed(data_mid_3_real));
  assign _zz_2247 = _zz_4973;
  assign _zz_6 = _zz_4976[31 : 0];
  assign _zz_2248 = _zz_4977;
  assign _zz_7 = _zz_4980[31 : 0];
  assign _zz_9 = 1'b1;
  assign _zz_2249 = _zz_4981;
  assign _zz_2250 = _zz_4989;
  assign _zz_10 = 1'b1;
  assign _zz_2251 = _zz_4997;
  assign _zz_2252 = _zz_5005;
  assign _zz_13 = ($signed(_zz_5013) * $signed(data_mid_5_real));
  assign _zz_2253 = _zz_5014;
  assign _zz_11 = _zz_5017[31 : 0];
  assign _zz_2254 = _zz_5018;
  assign _zz_12 = _zz_5021[31 : 0];
  assign _zz_14 = 1'b1;
  assign _zz_2255 = _zz_5022;
  assign _zz_2256 = _zz_5030;
  assign _zz_15 = 1'b1;
  assign _zz_2257 = _zz_5038;
  assign _zz_2258 = _zz_5046;
  assign _zz_18 = ($signed(_zz_5054) * $signed(data_mid_7_real));
  assign _zz_2259 = _zz_5055;
  assign _zz_16 = _zz_5058[31 : 0];
  assign _zz_2260 = _zz_5059;
  assign _zz_17 = _zz_5062[31 : 0];
  assign _zz_19 = 1'b1;
  assign _zz_2261 = _zz_5063;
  assign _zz_2262 = _zz_5071;
  assign _zz_20 = 1'b1;
  assign _zz_2263 = _zz_5079;
  assign _zz_2264 = _zz_5087;
  assign _zz_23 = ($signed(_zz_5095) * $signed(data_mid_9_real));
  assign _zz_2265 = _zz_5096;
  assign _zz_21 = _zz_5099[31 : 0];
  assign _zz_2266 = _zz_5100;
  assign _zz_22 = _zz_5103[31 : 0];
  assign _zz_24 = 1'b1;
  assign _zz_2267 = _zz_5104;
  assign _zz_2268 = _zz_5112;
  assign _zz_25 = 1'b1;
  assign _zz_2269 = _zz_5120;
  assign _zz_2270 = _zz_5128;
  assign _zz_28 = ($signed(_zz_5136) * $signed(data_mid_11_real));
  assign _zz_2271 = _zz_5137;
  assign _zz_26 = _zz_5140[31 : 0];
  assign _zz_2272 = _zz_5141;
  assign _zz_27 = _zz_5144[31 : 0];
  assign _zz_29 = 1'b1;
  assign _zz_2273 = _zz_5145;
  assign _zz_2274 = _zz_5153;
  assign _zz_30 = 1'b1;
  assign _zz_2275 = _zz_5161;
  assign _zz_2276 = _zz_5169;
  assign _zz_33 = ($signed(_zz_5177) * $signed(data_mid_13_real));
  assign _zz_2277 = _zz_5178;
  assign _zz_31 = _zz_5181[31 : 0];
  assign _zz_2278 = _zz_5182;
  assign _zz_32 = _zz_5185[31 : 0];
  assign _zz_34 = 1'b1;
  assign _zz_2279 = _zz_5186;
  assign _zz_2280 = _zz_5194;
  assign _zz_35 = 1'b1;
  assign _zz_2281 = _zz_5202;
  assign _zz_2282 = _zz_5210;
  assign _zz_38 = ($signed(_zz_5218) * $signed(data_mid_15_real));
  assign _zz_2283 = _zz_5219;
  assign _zz_36 = _zz_5222[31 : 0];
  assign _zz_2284 = _zz_5223;
  assign _zz_37 = _zz_5226[31 : 0];
  assign _zz_39 = 1'b1;
  assign _zz_2285 = _zz_5227;
  assign _zz_2286 = _zz_5235;
  assign _zz_40 = 1'b1;
  assign _zz_2287 = _zz_5243;
  assign _zz_2288 = _zz_5251;
  assign _zz_43 = ($signed(_zz_5259) * $signed(data_mid_17_real));
  assign _zz_2289 = _zz_5260;
  assign _zz_41 = _zz_5263[31 : 0];
  assign _zz_2290 = _zz_5264;
  assign _zz_42 = _zz_5267[31 : 0];
  assign _zz_44 = 1'b1;
  assign _zz_2291 = _zz_5268;
  assign _zz_2292 = _zz_5276;
  assign _zz_45 = 1'b1;
  assign _zz_2293 = _zz_5284;
  assign _zz_2294 = _zz_5292;
  assign _zz_48 = ($signed(_zz_5300) * $signed(data_mid_19_real));
  assign _zz_2295 = _zz_5301;
  assign _zz_46 = _zz_5304[31 : 0];
  assign _zz_2296 = _zz_5305;
  assign _zz_47 = _zz_5308[31 : 0];
  assign _zz_49 = 1'b1;
  assign _zz_2297 = _zz_5309;
  assign _zz_2298 = _zz_5317;
  assign _zz_50 = 1'b1;
  assign _zz_2299 = _zz_5325;
  assign _zz_2300 = _zz_5333;
  assign _zz_53 = ($signed(_zz_5341) * $signed(data_mid_21_real));
  assign _zz_2301 = _zz_5342;
  assign _zz_51 = _zz_5345[31 : 0];
  assign _zz_2302 = _zz_5346;
  assign _zz_52 = _zz_5349[31 : 0];
  assign _zz_54 = 1'b1;
  assign _zz_2303 = _zz_5350;
  assign _zz_2304 = _zz_5358;
  assign _zz_55 = 1'b1;
  assign _zz_2305 = _zz_5366;
  assign _zz_2306 = _zz_5374;
  assign _zz_58 = ($signed(_zz_5382) * $signed(data_mid_23_real));
  assign _zz_2307 = _zz_5383;
  assign _zz_56 = _zz_5386[31 : 0];
  assign _zz_2308 = _zz_5387;
  assign _zz_57 = _zz_5390[31 : 0];
  assign _zz_59 = 1'b1;
  assign _zz_2309 = _zz_5391;
  assign _zz_2310 = _zz_5399;
  assign _zz_60 = 1'b1;
  assign _zz_2311 = _zz_5407;
  assign _zz_2312 = _zz_5415;
  assign _zz_63 = ($signed(_zz_5423) * $signed(data_mid_25_real));
  assign _zz_2313 = _zz_5424;
  assign _zz_61 = _zz_5427[31 : 0];
  assign _zz_2314 = _zz_5428;
  assign _zz_62 = _zz_5431[31 : 0];
  assign _zz_64 = 1'b1;
  assign _zz_2315 = _zz_5432;
  assign _zz_2316 = _zz_5440;
  assign _zz_65 = 1'b1;
  assign _zz_2317 = _zz_5448;
  assign _zz_2318 = _zz_5456;
  assign _zz_68 = ($signed(_zz_5464) * $signed(data_mid_27_real));
  assign _zz_2319 = _zz_5465;
  assign _zz_66 = _zz_5468[31 : 0];
  assign _zz_2320 = _zz_5469;
  assign _zz_67 = _zz_5472[31 : 0];
  assign _zz_69 = 1'b1;
  assign _zz_2321 = _zz_5473;
  assign _zz_2322 = _zz_5481;
  assign _zz_70 = 1'b1;
  assign _zz_2323 = _zz_5489;
  assign _zz_2324 = _zz_5497;
  assign _zz_73 = ($signed(_zz_5505) * $signed(data_mid_29_real));
  assign _zz_2325 = _zz_5506;
  assign _zz_71 = _zz_5509[31 : 0];
  assign _zz_2326 = _zz_5510;
  assign _zz_72 = _zz_5513[31 : 0];
  assign _zz_74 = 1'b1;
  assign _zz_2327 = _zz_5514;
  assign _zz_2328 = _zz_5522;
  assign _zz_75 = 1'b1;
  assign _zz_2329 = _zz_5530;
  assign _zz_2330 = _zz_5538;
  assign _zz_78 = ($signed(_zz_5546) * $signed(data_mid_31_real));
  assign _zz_2331 = _zz_5547;
  assign _zz_76 = _zz_5550[31 : 0];
  assign _zz_2332 = _zz_5551;
  assign _zz_77 = _zz_5554[31 : 0];
  assign _zz_79 = 1'b1;
  assign _zz_2333 = _zz_5555;
  assign _zz_2334 = _zz_5563;
  assign _zz_80 = 1'b1;
  assign _zz_2335 = _zz_5571;
  assign _zz_2336 = _zz_5579;
  assign _zz_83 = ($signed(_zz_5587) * $signed(data_mid_33_real));
  assign _zz_2337 = _zz_5588;
  assign _zz_81 = _zz_5591[31 : 0];
  assign _zz_2338 = _zz_5592;
  assign _zz_82 = _zz_5595[31 : 0];
  assign _zz_84 = 1'b1;
  assign _zz_2339 = _zz_5596;
  assign _zz_2340 = _zz_5604;
  assign _zz_85 = 1'b1;
  assign _zz_2341 = _zz_5612;
  assign _zz_2342 = _zz_5620;
  assign _zz_88 = ($signed(_zz_5628) * $signed(data_mid_35_real));
  assign _zz_2343 = _zz_5629;
  assign _zz_86 = _zz_5632[31 : 0];
  assign _zz_2344 = _zz_5633;
  assign _zz_87 = _zz_5636[31 : 0];
  assign _zz_89 = 1'b1;
  assign _zz_2345 = _zz_5637;
  assign _zz_2346 = _zz_5645;
  assign _zz_90 = 1'b1;
  assign _zz_2347 = _zz_5653;
  assign _zz_2348 = _zz_5661;
  assign _zz_93 = ($signed(_zz_5669) * $signed(data_mid_37_real));
  assign _zz_2349 = _zz_5670;
  assign _zz_91 = _zz_5673[31 : 0];
  assign _zz_2350 = _zz_5674;
  assign _zz_92 = _zz_5677[31 : 0];
  assign _zz_94 = 1'b1;
  assign _zz_2351 = _zz_5678;
  assign _zz_2352 = _zz_5686;
  assign _zz_95 = 1'b1;
  assign _zz_2353 = _zz_5694;
  assign _zz_2354 = _zz_5702;
  assign _zz_98 = ($signed(_zz_5710) * $signed(data_mid_39_real));
  assign _zz_2355 = _zz_5711;
  assign _zz_96 = _zz_5714[31 : 0];
  assign _zz_2356 = _zz_5715;
  assign _zz_97 = _zz_5718[31 : 0];
  assign _zz_99 = 1'b1;
  assign _zz_2357 = _zz_5719;
  assign _zz_2358 = _zz_5727;
  assign _zz_100 = 1'b1;
  assign _zz_2359 = _zz_5735;
  assign _zz_2360 = _zz_5743;
  assign _zz_103 = ($signed(_zz_5751) * $signed(data_mid_41_real));
  assign _zz_2361 = _zz_5752;
  assign _zz_101 = _zz_5755[31 : 0];
  assign _zz_2362 = _zz_5756;
  assign _zz_102 = _zz_5759[31 : 0];
  assign _zz_104 = 1'b1;
  assign _zz_2363 = _zz_5760;
  assign _zz_2364 = _zz_5768;
  assign _zz_105 = 1'b1;
  assign _zz_2365 = _zz_5776;
  assign _zz_2366 = _zz_5784;
  assign _zz_108 = ($signed(_zz_5792) * $signed(data_mid_43_real));
  assign _zz_2367 = _zz_5793;
  assign _zz_106 = _zz_5796[31 : 0];
  assign _zz_2368 = _zz_5797;
  assign _zz_107 = _zz_5800[31 : 0];
  assign _zz_109 = 1'b1;
  assign _zz_2369 = _zz_5801;
  assign _zz_2370 = _zz_5809;
  assign _zz_110 = 1'b1;
  assign _zz_2371 = _zz_5817;
  assign _zz_2372 = _zz_5825;
  assign _zz_113 = ($signed(_zz_5833) * $signed(data_mid_45_real));
  assign _zz_2373 = _zz_5834;
  assign _zz_111 = _zz_5837[31 : 0];
  assign _zz_2374 = _zz_5838;
  assign _zz_112 = _zz_5841[31 : 0];
  assign _zz_114 = 1'b1;
  assign _zz_2375 = _zz_5842;
  assign _zz_2376 = _zz_5850;
  assign _zz_115 = 1'b1;
  assign _zz_2377 = _zz_5858;
  assign _zz_2378 = _zz_5866;
  assign _zz_118 = ($signed(_zz_5874) * $signed(data_mid_47_real));
  assign _zz_2379 = _zz_5875;
  assign _zz_116 = _zz_5878[31 : 0];
  assign _zz_2380 = _zz_5879;
  assign _zz_117 = _zz_5882[31 : 0];
  assign _zz_119 = 1'b1;
  assign _zz_2381 = _zz_5883;
  assign _zz_2382 = _zz_5891;
  assign _zz_120 = 1'b1;
  assign _zz_2383 = _zz_5899;
  assign _zz_2384 = _zz_5907;
  assign _zz_123 = ($signed(_zz_5915) * $signed(data_mid_49_real));
  assign _zz_2385 = _zz_5916;
  assign _zz_121 = _zz_5919[31 : 0];
  assign _zz_2386 = _zz_5920;
  assign _zz_122 = _zz_5923[31 : 0];
  assign _zz_124 = 1'b1;
  assign _zz_2387 = _zz_5924;
  assign _zz_2388 = _zz_5932;
  assign _zz_125 = 1'b1;
  assign _zz_2389 = _zz_5940;
  assign _zz_2390 = _zz_5948;
  assign _zz_128 = ($signed(_zz_5956) * $signed(data_mid_51_real));
  assign _zz_2391 = _zz_5957;
  assign _zz_126 = _zz_5960[31 : 0];
  assign _zz_2392 = _zz_5961;
  assign _zz_127 = _zz_5964[31 : 0];
  assign _zz_129 = 1'b1;
  assign _zz_2393 = _zz_5965;
  assign _zz_2394 = _zz_5973;
  assign _zz_130 = 1'b1;
  assign _zz_2395 = _zz_5981;
  assign _zz_2396 = _zz_5989;
  assign _zz_133 = ($signed(_zz_5997) * $signed(data_mid_53_real));
  assign _zz_2397 = _zz_5998;
  assign _zz_131 = _zz_6001[31 : 0];
  assign _zz_2398 = _zz_6002;
  assign _zz_132 = _zz_6005[31 : 0];
  assign _zz_134 = 1'b1;
  assign _zz_2399 = _zz_6006;
  assign _zz_2400 = _zz_6014;
  assign _zz_135 = 1'b1;
  assign _zz_2401 = _zz_6022;
  assign _zz_2402 = _zz_6030;
  assign _zz_138 = ($signed(_zz_6038) * $signed(data_mid_55_real));
  assign _zz_2403 = _zz_6039;
  assign _zz_136 = _zz_6042[31 : 0];
  assign _zz_2404 = _zz_6043;
  assign _zz_137 = _zz_6046[31 : 0];
  assign _zz_139 = 1'b1;
  assign _zz_2405 = _zz_6047;
  assign _zz_2406 = _zz_6055;
  assign _zz_140 = 1'b1;
  assign _zz_2407 = _zz_6063;
  assign _zz_2408 = _zz_6071;
  assign _zz_143 = ($signed(_zz_6079) * $signed(data_mid_57_real));
  assign _zz_2409 = _zz_6080;
  assign _zz_141 = _zz_6083[31 : 0];
  assign _zz_2410 = _zz_6084;
  assign _zz_142 = _zz_6087[31 : 0];
  assign _zz_144 = 1'b1;
  assign _zz_2411 = _zz_6088;
  assign _zz_2412 = _zz_6096;
  assign _zz_145 = 1'b1;
  assign _zz_2413 = _zz_6104;
  assign _zz_2414 = _zz_6112;
  assign _zz_148 = ($signed(_zz_6120) * $signed(data_mid_59_real));
  assign _zz_2415 = _zz_6121;
  assign _zz_146 = _zz_6124[31 : 0];
  assign _zz_2416 = _zz_6125;
  assign _zz_147 = _zz_6128[31 : 0];
  assign _zz_149 = 1'b1;
  assign _zz_2417 = _zz_6129;
  assign _zz_2418 = _zz_6137;
  assign _zz_150 = 1'b1;
  assign _zz_2419 = _zz_6145;
  assign _zz_2420 = _zz_6153;
  assign _zz_153 = ($signed(_zz_6161) * $signed(data_mid_61_real));
  assign _zz_2421 = _zz_6162;
  assign _zz_151 = _zz_6165[31 : 0];
  assign _zz_2422 = _zz_6166;
  assign _zz_152 = _zz_6169[31 : 0];
  assign _zz_154 = 1'b1;
  assign _zz_2423 = _zz_6170;
  assign _zz_2424 = _zz_6178;
  assign _zz_155 = 1'b1;
  assign _zz_2425 = _zz_6186;
  assign _zz_2426 = _zz_6194;
  assign _zz_158 = ($signed(_zz_6202) * $signed(data_mid_63_real));
  assign _zz_2427 = _zz_6203;
  assign _zz_156 = _zz_6206[31 : 0];
  assign _zz_2428 = _zz_6207;
  assign _zz_157 = _zz_6210[31 : 0];
  assign _zz_159 = 1'b1;
  assign _zz_2429 = _zz_6211;
  assign _zz_2430 = _zz_6219;
  assign _zz_160 = 1'b1;
  assign _zz_2431 = _zz_6227;
  assign _zz_2432 = _zz_6235;
  assign _zz_163 = ($signed(_zz_6243) * $signed(data_mid_65_real));
  assign _zz_2433 = _zz_6244;
  assign _zz_161 = _zz_6247[31 : 0];
  assign _zz_2434 = _zz_6248;
  assign _zz_162 = _zz_6251[31 : 0];
  assign _zz_164 = 1'b1;
  assign _zz_2435 = _zz_6252;
  assign _zz_2436 = _zz_6260;
  assign _zz_165 = 1'b1;
  assign _zz_2437 = _zz_6268;
  assign _zz_2438 = _zz_6276;
  assign _zz_168 = ($signed(_zz_6284) * $signed(data_mid_67_real));
  assign _zz_2439 = _zz_6285;
  assign _zz_166 = _zz_6288[31 : 0];
  assign _zz_2440 = _zz_6289;
  assign _zz_167 = _zz_6292[31 : 0];
  assign _zz_169 = 1'b1;
  assign _zz_2441 = _zz_6293;
  assign _zz_2442 = _zz_6301;
  assign _zz_170 = 1'b1;
  assign _zz_2443 = _zz_6309;
  assign _zz_2444 = _zz_6317;
  assign _zz_173 = ($signed(_zz_6325) * $signed(data_mid_69_real));
  assign _zz_2445 = _zz_6326;
  assign _zz_171 = _zz_6329[31 : 0];
  assign _zz_2446 = _zz_6330;
  assign _zz_172 = _zz_6333[31 : 0];
  assign _zz_174 = 1'b1;
  assign _zz_2447 = _zz_6334;
  assign _zz_2448 = _zz_6342;
  assign _zz_175 = 1'b1;
  assign _zz_2449 = _zz_6350;
  assign _zz_2450 = _zz_6358;
  assign _zz_178 = ($signed(_zz_6366) * $signed(data_mid_71_real));
  assign _zz_2451 = _zz_6367;
  assign _zz_176 = _zz_6370[31 : 0];
  assign _zz_2452 = _zz_6371;
  assign _zz_177 = _zz_6374[31 : 0];
  assign _zz_179 = 1'b1;
  assign _zz_2453 = _zz_6375;
  assign _zz_2454 = _zz_6383;
  assign _zz_180 = 1'b1;
  assign _zz_2455 = _zz_6391;
  assign _zz_2456 = _zz_6399;
  assign _zz_183 = ($signed(_zz_6407) * $signed(data_mid_73_real));
  assign _zz_2457 = _zz_6408;
  assign _zz_181 = _zz_6411[31 : 0];
  assign _zz_2458 = _zz_6412;
  assign _zz_182 = _zz_6415[31 : 0];
  assign _zz_184 = 1'b1;
  assign _zz_2459 = _zz_6416;
  assign _zz_2460 = _zz_6424;
  assign _zz_185 = 1'b1;
  assign _zz_2461 = _zz_6432;
  assign _zz_2462 = _zz_6440;
  assign _zz_188 = ($signed(_zz_6448) * $signed(data_mid_75_real));
  assign _zz_2463 = _zz_6449;
  assign _zz_186 = _zz_6452[31 : 0];
  assign _zz_2464 = _zz_6453;
  assign _zz_187 = _zz_6456[31 : 0];
  assign _zz_189 = 1'b1;
  assign _zz_2465 = _zz_6457;
  assign _zz_2466 = _zz_6465;
  assign _zz_190 = 1'b1;
  assign _zz_2467 = _zz_6473;
  assign _zz_2468 = _zz_6481;
  assign _zz_193 = ($signed(_zz_6489) * $signed(data_mid_77_real));
  assign _zz_2469 = _zz_6490;
  assign _zz_191 = _zz_6493[31 : 0];
  assign _zz_2470 = _zz_6494;
  assign _zz_192 = _zz_6497[31 : 0];
  assign _zz_194 = 1'b1;
  assign _zz_2471 = _zz_6498;
  assign _zz_2472 = _zz_6506;
  assign _zz_195 = 1'b1;
  assign _zz_2473 = _zz_6514;
  assign _zz_2474 = _zz_6522;
  assign _zz_198 = ($signed(_zz_6530) * $signed(data_mid_79_real));
  assign _zz_2475 = _zz_6531;
  assign _zz_196 = _zz_6534[31 : 0];
  assign _zz_2476 = _zz_6535;
  assign _zz_197 = _zz_6538[31 : 0];
  assign _zz_199 = 1'b1;
  assign _zz_2477 = _zz_6539;
  assign _zz_2478 = _zz_6547;
  assign _zz_200 = 1'b1;
  assign _zz_2479 = _zz_6555;
  assign _zz_2480 = _zz_6563;
  assign _zz_203 = ($signed(_zz_6571) * $signed(data_mid_81_real));
  assign _zz_2481 = _zz_6572;
  assign _zz_201 = _zz_6575[31 : 0];
  assign _zz_2482 = _zz_6576;
  assign _zz_202 = _zz_6579[31 : 0];
  assign _zz_204 = 1'b1;
  assign _zz_2483 = _zz_6580;
  assign _zz_2484 = _zz_6588;
  assign _zz_205 = 1'b1;
  assign _zz_2485 = _zz_6596;
  assign _zz_2486 = _zz_6604;
  assign _zz_208 = ($signed(_zz_6612) * $signed(data_mid_83_real));
  assign _zz_2487 = _zz_6613;
  assign _zz_206 = _zz_6616[31 : 0];
  assign _zz_2488 = _zz_6617;
  assign _zz_207 = _zz_6620[31 : 0];
  assign _zz_209 = 1'b1;
  assign _zz_2489 = _zz_6621;
  assign _zz_2490 = _zz_6629;
  assign _zz_210 = 1'b1;
  assign _zz_2491 = _zz_6637;
  assign _zz_2492 = _zz_6645;
  assign _zz_213 = ($signed(_zz_6653) * $signed(data_mid_85_real));
  assign _zz_2493 = _zz_6654;
  assign _zz_211 = _zz_6657[31 : 0];
  assign _zz_2494 = _zz_6658;
  assign _zz_212 = _zz_6661[31 : 0];
  assign _zz_214 = 1'b1;
  assign _zz_2495 = _zz_6662;
  assign _zz_2496 = _zz_6670;
  assign _zz_215 = 1'b1;
  assign _zz_2497 = _zz_6678;
  assign _zz_2498 = _zz_6686;
  assign _zz_218 = ($signed(_zz_6694) * $signed(data_mid_87_real));
  assign _zz_2499 = _zz_6695;
  assign _zz_216 = _zz_6698[31 : 0];
  assign _zz_2500 = _zz_6699;
  assign _zz_217 = _zz_6702[31 : 0];
  assign _zz_219 = 1'b1;
  assign _zz_2501 = _zz_6703;
  assign _zz_2502 = _zz_6711;
  assign _zz_220 = 1'b1;
  assign _zz_2503 = _zz_6719;
  assign _zz_2504 = _zz_6727;
  assign _zz_223 = ($signed(_zz_6735) * $signed(data_mid_89_real));
  assign _zz_2505 = _zz_6736;
  assign _zz_221 = _zz_6739[31 : 0];
  assign _zz_2506 = _zz_6740;
  assign _zz_222 = _zz_6743[31 : 0];
  assign _zz_224 = 1'b1;
  assign _zz_2507 = _zz_6744;
  assign _zz_2508 = _zz_6752;
  assign _zz_225 = 1'b1;
  assign _zz_2509 = _zz_6760;
  assign _zz_2510 = _zz_6768;
  assign _zz_228 = ($signed(_zz_6776) * $signed(data_mid_91_real));
  assign _zz_2511 = _zz_6777;
  assign _zz_226 = _zz_6780[31 : 0];
  assign _zz_2512 = _zz_6781;
  assign _zz_227 = _zz_6784[31 : 0];
  assign _zz_229 = 1'b1;
  assign _zz_2513 = _zz_6785;
  assign _zz_2514 = _zz_6793;
  assign _zz_230 = 1'b1;
  assign _zz_2515 = _zz_6801;
  assign _zz_2516 = _zz_6809;
  assign _zz_233 = ($signed(_zz_6817) * $signed(data_mid_93_real));
  assign _zz_2517 = _zz_6818;
  assign _zz_231 = _zz_6821[31 : 0];
  assign _zz_2518 = _zz_6822;
  assign _zz_232 = _zz_6825[31 : 0];
  assign _zz_234 = 1'b1;
  assign _zz_2519 = _zz_6826;
  assign _zz_2520 = _zz_6834;
  assign _zz_235 = 1'b1;
  assign _zz_2521 = _zz_6842;
  assign _zz_2522 = _zz_6850;
  assign _zz_238 = ($signed(_zz_6858) * $signed(data_mid_95_real));
  assign _zz_2523 = _zz_6859;
  assign _zz_236 = _zz_6862[31 : 0];
  assign _zz_2524 = _zz_6863;
  assign _zz_237 = _zz_6866[31 : 0];
  assign _zz_239 = 1'b1;
  assign _zz_2525 = _zz_6867;
  assign _zz_2526 = _zz_6875;
  assign _zz_240 = 1'b1;
  assign _zz_2527 = _zz_6883;
  assign _zz_2528 = _zz_6891;
  assign _zz_243 = ($signed(_zz_6899) * $signed(data_mid_97_real));
  assign _zz_2529 = _zz_6900;
  assign _zz_241 = _zz_6903[31 : 0];
  assign _zz_2530 = _zz_6904;
  assign _zz_242 = _zz_6907[31 : 0];
  assign _zz_244 = 1'b1;
  assign _zz_2531 = _zz_6908;
  assign _zz_2532 = _zz_6916;
  assign _zz_245 = 1'b1;
  assign _zz_2533 = _zz_6924;
  assign _zz_2534 = _zz_6932;
  assign _zz_248 = ($signed(_zz_6940) * $signed(data_mid_99_real));
  assign _zz_2535 = _zz_6941;
  assign _zz_246 = _zz_6944[31 : 0];
  assign _zz_2536 = _zz_6945;
  assign _zz_247 = _zz_6948[31 : 0];
  assign _zz_249 = 1'b1;
  assign _zz_2537 = _zz_6949;
  assign _zz_2538 = _zz_6957;
  assign _zz_250 = 1'b1;
  assign _zz_2539 = _zz_6965;
  assign _zz_2540 = _zz_6973;
  assign _zz_253 = ($signed(_zz_6981) * $signed(data_mid_101_real));
  assign _zz_2541 = _zz_6982;
  assign _zz_251 = _zz_6985[31 : 0];
  assign _zz_2542 = _zz_6986;
  assign _zz_252 = _zz_6989[31 : 0];
  assign _zz_254 = 1'b1;
  assign _zz_2543 = _zz_6990;
  assign _zz_2544 = _zz_6998;
  assign _zz_255 = 1'b1;
  assign _zz_2545 = _zz_7006;
  assign _zz_2546 = _zz_7014;
  assign _zz_258 = ($signed(_zz_7022) * $signed(data_mid_103_real));
  assign _zz_2547 = _zz_7023;
  assign _zz_256 = _zz_7026[31 : 0];
  assign _zz_2548 = _zz_7027;
  assign _zz_257 = _zz_7030[31 : 0];
  assign _zz_259 = 1'b1;
  assign _zz_2549 = _zz_7031;
  assign _zz_2550 = _zz_7039;
  assign _zz_260 = 1'b1;
  assign _zz_2551 = _zz_7047;
  assign _zz_2552 = _zz_7055;
  assign _zz_263 = ($signed(_zz_7063) * $signed(data_mid_105_real));
  assign _zz_2553 = _zz_7064;
  assign _zz_261 = _zz_7067[31 : 0];
  assign _zz_2554 = _zz_7068;
  assign _zz_262 = _zz_7071[31 : 0];
  assign _zz_264 = 1'b1;
  assign _zz_2555 = _zz_7072;
  assign _zz_2556 = _zz_7080;
  assign _zz_265 = 1'b1;
  assign _zz_2557 = _zz_7088;
  assign _zz_2558 = _zz_7096;
  assign _zz_268 = ($signed(_zz_7104) * $signed(data_mid_107_real));
  assign _zz_2559 = _zz_7105;
  assign _zz_266 = _zz_7108[31 : 0];
  assign _zz_2560 = _zz_7109;
  assign _zz_267 = _zz_7112[31 : 0];
  assign _zz_269 = 1'b1;
  assign _zz_2561 = _zz_7113;
  assign _zz_2562 = _zz_7121;
  assign _zz_270 = 1'b1;
  assign _zz_2563 = _zz_7129;
  assign _zz_2564 = _zz_7137;
  assign _zz_273 = ($signed(_zz_7145) * $signed(data_mid_109_real));
  assign _zz_2565 = _zz_7146;
  assign _zz_271 = _zz_7149[31 : 0];
  assign _zz_2566 = _zz_7150;
  assign _zz_272 = _zz_7153[31 : 0];
  assign _zz_274 = 1'b1;
  assign _zz_2567 = _zz_7154;
  assign _zz_2568 = _zz_7162;
  assign _zz_275 = 1'b1;
  assign _zz_2569 = _zz_7170;
  assign _zz_2570 = _zz_7178;
  assign _zz_278 = ($signed(_zz_7186) * $signed(data_mid_111_real));
  assign _zz_2571 = _zz_7187;
  assign _zz_276 = _zz_7190[31 : 0];
  assign _zz_2572 = _zz_7191;
  assign _zz_277 = _zz_7194[31 : 0];
  assign _zz_279 = 1'b1;
  assign _zz_2573 = _zz_7195;
  assign _zz_2574 = _zz_7203;
  assign _zz_280 = 1'b1;
  assign _zz_2575 = _zz_7211;
  assign _zz_2576 = _zz_7219;
  assign _zz_283 = ($signed(_zz_7227) * $signed(data_mid_113_real));
  assign _zz_2577 = _zz_7228;
  assign _zz_281 = _zz_7231[31 : 0];
  assign _zz_2578 = _zz_7232;
  assign _zz_282 = _zz_7235[31 : 0];
  assign _zz_284 = 1'b1;
  assign _zz_2579 = _zz_7236;
  assign _zz_2580 = _zz_7244;
  assign _zz_285 = 1'b1;
  assign _zz_2581 = _zz_7252;
  assign _zz_2582 = _zz_7260;
  assign _zz_288 = ($signed(_zz_7268) * $signed(data_mid_115_real));
  assign _zz_2583 = _zz_7269;
  assign _zz_286 = _zz_7272[31 : 0];
  assign _zz_2584 = _zz_7273;
  assign _zz_287 = _zz_7276[31 : 0];
  assign _zz_289 = 1'b1;
  assign _zz_2585 = _zz_7277;
  assign _zz_2586 = _zz_7285;
  assign _zz_290 = 1'b1;
  assign _zz_2587 = _zz_7293;
  assign _zz_2588 = _zz_7301;
  assign _zz_293 = ($signed(_zz_7309) * $signed(data_mid_117_real));
  assign _zz_2589 = _zz_7310;
  assign _zz_291 = _zz_7313[31 : 0];
  assign _zz_2590 = _zz_7314;
  assign _zz_292 = _zz_7317[31 : 0];
  assign _zz_294 = 1'b1;
  assign _zz_2591 = _zz_7318;
  assign _zz_2592 = _zz_7326;
  assign _zz_295 = 1'b1;
  assign _zz_2593 = _zz_7334;
  assign _zz_2594 = _zz_7342;
  assign _zz_298 = ($signed(_zz_7350) * $signed(data_mid_119_real));
  assign _zz_2595 = _zz_7351;
  assign _zz_296 = _zz_7354[31 : 0];
  assign _zz_2596 = _zz_7355;
  assign _zz_297 = _zz_7358[31 : 0];
  assign _zz_299 = 1'b1;
  assign _zz_2597 = _zz_7359;
  assign _zz_2598 = _zz_7367;
  assign _zz_300 = 1'b1;
  assign _zz_2599 = _zz_7375;
  assign _zz_2600 = _zz_7383;
  assign _zz_303 = ($signed(_zz_7391) * $signed(data_mid_121_real));
  assign _zz_2601 = _zz_7392;
  assign _zz_301 = _zz_7395[31 : 0];
  assign _zz_2602 = _zz_7396;
  assign _zz_302 = _zz_7399[31 : 0];
  assign _zz_304 = 1'b1;
  assign _zz_2603 = _zz_7400;
  assign _zz_2604 = _zz_7408;
  assign _zz_305 = 1'b1;
  assign _zz_2605 = _zz_7416;
  assign _zz_2606 = _zz_7424;
  assign _zz_308 = ($signed(_zz_7432) * $signed(data_mid_123_real));
  assign _zz_2607 = _zz_7433;
  assign _zz_306 = _zz_7436[31 : 0];
  assign _zz_2608 = _zz_7437;
  assign _zz_307 = _zz_7440[31 : 0];
  assign _zz_309 = 1'b1;
  assign _zz_2609 = _zz_7441;
  assign _zz_2610 = _zz_7449;
  assign _zz_310 = 1'b1;
  assign _zz_2611 = _zz_7457;
  assign _zz_2612 = _zz_7465;
  assign _zz_313 = ($signed(_zz_7473) * $signed(data_mid_125_real));
  assign _zz_2613 = _zz_7474;
  assign _zz_311 = _zz_7477[31 : 0];
  assign _zz_2614 = _zz_7478;
  assign _zz_312 = _zz_7481[31 : 0];
  assign _zz_314 = 1'b1;
  assign _zz_2615 = _zz_7482;
  assign _zz_2616 = _zz_7490;
  assign _zz_315 = 1'b1;
  assign _zz_2617 = _zz_7498;
  assign _zz_2618 = _zz_7506;
  assign _zz_318 = ($signed(_zz_7514) * $signed(data_mid_127_real));
  assign _zz_2619 = _zz_7515;
  assign _zz_316 = _zz_7518[31 : 0];
  assign _zz_2620 = _zz_7519;
  assign _zz_317 = _zz_7522[31 : 0];
  assign _zz_319 = 1'b1;
  assign _zz_2621 = _zz_7523;
  assign _zz_2622 = _zz_7531;
  assign _zz_320 = 1'b1;
  assign _zz_2623 = _zz_7539;
  assign _zz_2624 = _zz_7547;
  assign _zz_323 = ($signed(_zz_7555) * $signed(data_mid_2_real));
  assign _zz_2625 = _zz_7556;
  assign _zz_321 = _zz_7559[31 : 0];
  assign _zz_2626 = _zz_7560;
  assign _zz_322 = _zz_7563[31 : 0];
  assign _zz_324 = 1'b1;
  assign _zz_2627 = _zz_7564;
  assign _zz_2628 = _zz_7572;
  assign _zz_325 = 1'b1;
  assign _zz_2629 = _zz_7580;
  assign _zz_2630 = _zz_7588;
  assign _zz_328 = ($signed(_zz_7596) * $signed(data_mid_3_real));
  assign _zz_2631 = _zz_7597;
  assign _zz_326 = _zz_7600[31 : 0];
  assign _zz_2632 = _zz_7601;
  assign _zz_327 = _zz_7604[31 : 0];
  assign _zz_329 = 1'b1;
  assign _zz_2633 = _zz_7605;
  assign _zz_2634 = _zz_7613;
  assign _zz_330 = 1'b1;
  assign _zz_2635 = _zz_7621;
  assign _zz_2636 = _zz_7629;
  assign _zz_333 = ($signed(_zz_7637) * $signed(data_mid_6_real));
  assign _zz_2637 = _zz_7638;
  assign _zz_331 = _zz_7641[31 : 0];
  assign _zz_2638 = _zz_7642;
  assign _zz_332 = _zz_7645[31 : 0];
  assign _zz_334 = 1'b1;
  assign _zz_2639 = _zz_7646;
  assign _zz_2640 = _zz_7654;
  assign _zz_335 = 1'b1;
  assign _zz_2641 = _zz_7662;
  assign _zz_2642 = _zz_7670;
  assign _zz_338 = ($signed(_zz_7678) * $signed(data_mid_7_real));
  assign _zz_2643 = _zz_7679;
  assign _zz_336 = _zz_7682[31 : 0];
  assign _zz_2644 = _zz_7683;
  assign _zz_337 = _zz_7686[31 : 0];
  assign _zz_339 = 1'b1;
  assign _zz_2645 = _zz_7687;
  assign _zz_2646 = _zz_7695;
  assign _zz_340 = 1'b1;
  assign _zz_2647 = _zz_7703;
  assign _zz_2648 = _zz_7711;
  assign _zz_343 = ($signed(_zz_7719) * $signed(data_mid_10_real));
  assign _zz_2649 = _zz_7720;
  assign _zz_341 = _zz_7723[31 : 0];
  assign _zz_2650 = _zz_7724;
  assign _zz_342 = _zz_7727[31 : 0];
  assign _zz_344 = 1'b1;
  assign _zz_2651 = _zz_7728;
  assign _zz_2652 = _zz_7736;
  assign _zz_345 = 1'b1;
  assign _zz_2653 = _zz_7744;
  assign _zz_2654 = _zz_7752;
  assign _zz_348 = ($signed(_zz_7760) * $signed(data_mid_11_real));
  assign _zz_2655 = _zz_7761;
  assign _zz_346 = _zz_7764[31 : 0];
  assign _zz_2656 = _zz_7765;
  assign _zz_347 = _zz_7768[31 : 0];
  assign _zz_349 = 1'b1;
  assign _zz_2657 = _zz_7769;
  assign _zz_2658 = _zz_7777;
  assign _zz_350 = 1'b1;
  assign _zz_2659 = _zz_7785;
  assign _zz_2660 = _zz_7793;
  assign _zz_353 = ($signed(_zz_7801) * $signed(data_mid_14_real));
  assign _zz_2661 = _zz_7802;
  assign _zz_351 = _zz_7805[31 : 0];
  assign _zz_2662 = _zz_7806;
  assign _zz_352 = _zz_7809[31 : 0];
  assign _zz_354 = 1'b1;
  assign _zz_2663 = _zz_7810;
  assign _zz_2664 = _zz_7818;
  assign _zz_355 = 1'b1;
  assign _zz_2665 = _zz_7826;
  assign _zz_2666 = _zz_7834;
  assign _zz_358 = ($signed(_zz_7842) * $signed(data_mid_15_real));
  assign _zz_2667 = _zz_7843;
  assign _zz_356 = _zz_7846[31 : 0];
  assign _zz_2668 = _zz_7847;
  assign _zz_357 = _zz_7850[31 : 0];
  assign _zz_359 = 1'b1;
  assign _zz_2669 = _zz_7851;
  assign _zz_2670 = _zz_7859;
  assign _zz_360 = 1'b1;
  assign _zz_2671 = _zz_7867;
  assign _zz_2672 = _zz_7875;
  assign _zz_363 = ($signed(_zz_7883) * $signed(data_mid_18_real));
  assign _zz_2673 = _zz_7884;
  assign _zz_361 = _zz_7887[31 : 0];
  assign _zz_2674 = _zz_7888;
  assign _zz_362 = _zz_7891[31 : 0];
  assign _zz_364 = 1'b1;
  assign _zz_2675 = _zz_7892;
  assign _zz_2676 = _zz_7900;
  assign _zz_365 = 1'b1;
  assign _zz_2677 = _zz_7908;
  assign _zz_2678 = _zz_7916;
  assign _zz_368 = ($signed(_zz_7924) * $signed(data_mid_19_real));
  assign _zz_2679 = _zz_7925;
  assign _zz_366 = _zz_7928[31 : 0];
  assign _zz_2680 = _zz_7929;
  assign _zz_367 = _zz_7932[31 : 0];
  assign _zz_369 = 1'b1;
  assign _zz_2681 = _zz_7933;
  assign _zz_2682 = _zz_7941;
  assign _zz_370 = 1'b1;
  assign _zz_2683 = _zz_7949;
  assign _zz_2684 = _zz_7957;
  assign _zz_373 = ($signed(_zz_7965) * $signed(data_mid_22_real));
  assign _zz_2685 = _zz_7966;
  assign _zz_371 = _zz_7969[31 : 0];
  assign _zz_2686 = _zz_7970;
  assign _zz_372 = _zz_7973[31 : 0];
  assign _zz_374 = 1'b1;
  assign _zz_2687 = _zz_7974;
  assign _zz_2688 = _zz_7982;
  assign _zz_375 = 1'b1;
  assign _zz_2689 = _zz_7990;
  assign _zz_2690 = _zz_7998;
  assign _zz_378 = ($signed(_zz_8006) * $signed(data_mid_23_real));
  assign _zz_2691 = _zz_8007;
  assign _zz_376 = _zz_8010[31 : 0];
  assign _zz_2692 = _zz_8011;
  assign _zz_377 = _zz_8014[31 : 0];
  assign _zz_379 = 1'b1;
  assign _zz_2693 = _zz_8015;
  assign _zz_2694 = _zz_8023;
  assign _zz_380 = 1'b1;
  assign _zz_2695 = _zz_8031;
  assign _zz_2696 = _zz_8039;
  assign _zz_383 = ($signed(_zz_8047) * $signed(data_mid_26_real));
  assign _zz_2697 = _zz_8048;
  assign _zz_381 = _zz_8051[31 : 0];
  assign _zz_2698 = _zz_8052;
  assign _zz_382 = _zz_8055[31 : 0];
  assign _zz_384 = 1'b1;
  assign _zz_2699 = _zz_8056;
  assign _zz_2700 = _zz_8064;
  assign _zz_385 = 1'b1;
  assign _zz_2701 = _zz_8072;
  assign _zz_2702 = _zz_8080;
  assign _zz_388 = ($signed(_zz_8088) * $signed(data_mid_27_real));
  assign _zz_2703 = _zz_8089;
  assign _zz_386 = _zz_8092[31 : 0];
  assign _zz_2704 = _zz_8093;
  assign _zz_387 = _zz_8096[31 : 0];
  assign _zz_389 = 1'b1;
  assign _zz_2705 = _zz_8097;
  assign _zz_2706 = _zz_8105;
  assign _zz_390 = 1'b1;
  assign _zz_2707 = _zz_8113;
  assign _zz_2708 = _zz_8121;
  assign _zz_393 = ($signed(_zz_8129) * $signed(data_mid_30_real));
  assign _zz_2709 = _zz_8130;
  assign _zz_391 = _zz_8133[31 : 0];
  assign _zz_2710 = _zz_8134;
  assign _zz_392 = _zz_8137[31 : 0];
  assign _zz_394 = 1'b1;
  assign _zz_2711 = _zz_8138;
  assign _zz_2712 = _zz_8146;
  assign _zz_395 = 1'b1;
  assign _zz_2713 = _zz_8154;
  assign _zz_2714 = _zz_8162;
  assign _zz_398 = ($signed(_zz_8170) * $signed(data_mid_31_real));
  assign _zz_2715 = _zz_8171;
  assign _zz_396 = _zz_8174[31 : 0];
  assign _zz_2716 = _zz_8175;
  assign _zz_397 = _zz_8178[31 : 0];
  assign _zz_399 = 1'b1;
  assign _zz_2717 = _zz_8179;
  assign _zz_2718 = _zz_8187;
  assign _zz_400 = 1'b1;
  assign _zz_2719 = _zz_8195;
  assign _zz_2720 = _zz_8203;
  assign _zz_403 = ($signed(_zz_8211) * $signed(data_mid_34_real));
  assign _zz_2721 = _zz_8212;
  assign _zz_401 = _zz_8215[31 : 0];
  assign _zz_2722 = _zz_8216;
  assign _zz_402 = _zz_8219[31 : 0];
  assign _zz_404 = 1'b1;
  assign _zz_2723 = _zz_8220;
  assign _zz_2724 = _zz_8228;
  assign _zz_405 = 1'b1;
  assign _zz_2725 = _zz_8236;
  assign _zz_2726 = _zz_8244;
  assign _zz_408 = ($signed(_zz_8252) * $signed(data_mid_35_real));
  assign _zz_2727 = _zz_8253;
  assign _zz_406 = _zz_8256[31 : 0];
  assign _zz_2728 = _zz_8257;
  assign _zz_407 = _zz_8260[31 : 0];
  assign _zz_409 = 1'b1;
  assign _zz_2729 = _zz_8261;
  assign _zz_2730 = _zz_8269;
  assign _zz_410 = 1'b1;
  assign _zz_2731 = _zz_8277;
  assign _zz_2732 = _zz_8285;
  assign _zz_413 = ($signed(_zz_8293) * $signed(data_mid_38_real));
  assign _zz_2733 = _zz_8294;
  assign _zz_411 = _zz_8297[31 : 0];
  assign _zz_2734 = _zz_8298;
  assign _zz_412 = _zz_8301[31 : 0];
  assign _zz_414 = 1'b1;
  assign _zz_2735 = _zz_8302;
  assign _zz_2736 = _zz_8310;
  assign _zz_415 = 1'b1;
  assign _zz_2737 = _zz_8318;
  assign _zz_2738 = _zz_8326;
  assign _zz_418 = ($signed(_zz_8334) * $signed(data_mid_39_real));
  assign _zz_2739 = _zz_8335;
  assign _zz_416 = _zz_8338[31 : 0];
  assign _zz_2740 = _zz_8339;
  assign _zz_417 = _zz_8342[31 : 0];
  assign _zz_419 = 1'b1;
  assign _zz_2741 = _zz_8343;
  assign _zz_2742 = _zz_8351;
  assign _zz_420 = 1'b1;
  assign _zz_2743 = _zz_8359;
  assign _zz_2744 = _zz_8367;
  assign _zz_423 = ($signed(_zz_8375) * $signed(data_mid_42_real));
  assign _zz_2745 = _zz_8376;
  assign _zz_421 = _zz_8379[31 : 0];
  assign _zz_2746 = _zz_8380;
  assign _zz_422 = _zz_8383[31 : 0];
  assign _zz_424 = 1'b1;
  assign _zz_2747 = _zz_8384;
  assign _zz_2748 = _zz_8392;
  assign _zz_425 = 1'b1;
  assign _zz_2749 = _zz_8400;
  assign _zz_2750 = _zz_8408;
  assign _zz_428 = ($signed(_zz_8416) * $signed(data_mid_43_real));
  assign _zz_2751 = _zz_8417;
  assign _zz_426 = _zz_8420[31 : 0];
  assign _zz_2752 = _zz_8421;
  assign _zz_427 = _zz_8424[31 : 0];
  assign _zz_429 = 1'b1;
  assign _zz_2753 = _zz_8425;
  assign _zz_2754 = _zz_8433;
  assign _zz_430 = 1'b1;
  assign _zz_2755 = _zz_8441;
  assign _zz_2756 = _zz_8449;
  assign _zz_433 = ($signed(_zz_8457) * $signed(data_mid_46_real));
  assign _zz_2757 = _zz_8458;
  assign _zz_431 = _zz_8461[31 : 0];
  assign _zz_2758 = _zz_8462;
  assign _zz_432 = _zz_8465[31 : 0];
  assign _zz_434 = 1'b1;
  assign _zz_2759 = _zz_8466;
  assign _zz_2760 = _zz_8474;
  assign _zz_435 = 1'b1;
  assign _zz_2761 = _zz_8482;
  assign _zz_2762 = _zz_8490;
  assign _zz_438 = ($signed(_zz_8498) * $signed(data_mid_47_real));
  assign _zz_2763 = _zz_8499;
  assign _zz_436 = _zz_8502[31 : 0];
  assign _zz_2764 = _zz_8503;
  assign _zz_437 = _zz_8506[31 : 0];
  assign _zz_439 = 1'b1;
  assign _zz_2765 = _zz_8507;
  assign _zz_2766 = _zz_8515;
  assign _zz_440 = 1'b1;
  assign _zz_2767 = _zz_8523;
  assign _zz_2768 = _zz_8531;
  assign _zz_443 = ($signed(_zz_8539) * $signed(data_mid_50_real));
  assign _zz_2769 = _zz_8540;
  assign _zz_441 = _zz_8543[31 : 0];
  assign _zz_2770 = _zz_8544;
  assign _zz_442 = _zz_8547[31 : 0];
  assign _zz_444 = 1'b1;
  assign _zz_2771 = _zz_8548;
  assign _zz_2772 = _zz_8556;
  assign _zz_445 = 1'b1;
  assign _zz_2773 = _zz_8564;
  assign _zz_2774 = _zz_8572;
  assign _zz_448 = ($signed(_zz_8580) * $signed(data_mid_51_real));
  assign _zz_2775 = _zz_8581;
  assign _zz_446 = _zz_8584[31 : 0];
  assign _zz_2776 = _zz_8585;
  assign _zz_447 = _zz_8588[31 : 0];
  assign _zz_449 = 1'b1;
  assign _zz_2777 = _zz_8589;
  assign _zz_2778 = _zz_8597;
  assign _zz_450 = 1'b1;
  assign _zz_2779 = _zz_8605;
  assign _zz_2780 = _zz_8613;
  assign _zz_453 = ($signed(_zz_8621) * $signed(data_mid_54_real));
  assign _zz_2781 = _zz_8622;
  assign _zz_451 = _zz_8625[31 : 0];
  assign _zz_2782 = _zz_8626;
  assign _zz_452 = _zz_8629[31 : 0];
  assign _zz_454 = 1'b1;
  assign _zz_2783 = _zz_8630;
  assign _zz_2784 = _zz_8638;
  assign _zz_455 = 1'b1;
  assign _zz_2785 = _zz_8646;
  assign _zz_2786 = _zz_8654;
  assign _zz_458 = ($signed(_zz_8662) * $signed(data_mid_55_real));
  assign _zz_2787 = _zz_8663;
  assign _zz_456 = _zz_8666[31 : 0];
  assign _zz_2788 = _zz_8667;
  assign _zz_457 = _zz_8670[31 : 0];
  assign _zz_459 = 1'b1;
  assign _zz_2789 = _zz_8671;
  assign _zz_2790 = _zz_8679;
  assign _zz_460 = 1'b1;
  assign _zz_2791 = _zz_8687;
  assign _zz_2792 = _zz_8695;
  assign _zz_463 = ($signed(_zz_8703) * $signed(data_mid_58_real));
  assign _zz_2793 = _zz_8704;
  assign _zz_461 = _zz_8707[31 : 0];
  assign _zz_2794 = _zz_8708;
  assign _zz_462 = _zz_8711[31 : 0];
  assign _zz_464 = 1'b1;
  assign _zz_2795 = _zz_8712;
  assign _zz_2796 = _zz_8720;
  assign _zz_465 = 1'b1;
  assign _zz_2797 = _zz_8728;
  assign _zz_2798 = _zz_8736;
  assign _zz_468 = ($signed(_zz_8744) * $signed(data_mid_59_real));
  assign _zz_2799 = _zz_8745;
  assign _zz_466 = _zz_8748[31 : 0];
  assign _zz_2800 = _zz_8749;
  assign _zz_467 = _zz_8752[31 : 0];
  assign _zz_469 = 1'b1;
  assign _zz_2801 = _zz_8753;
  assign _zz_2802 = _zz_8761;
  assign _zz_470 = 1'b1;
  assign _zz_2803 = _zz_8769;
  assign _zz_2804 = _zz_8777;
  assign _zz_473 = ($signed(_zz_8785) * $signed(data_mid_62_real));
  assign _zz_2805 = _zz_8786;
  assign _zz_471 = _zz_8789[31 : 0];
  assign _zz_2806 = _zz_8790;
  assign _zz_472 = _zz_8793[31 : 0];
  assign _zz_474 = 1'b1;
  assign _zz_2807 = _zz_8794;
  assign _zz_2808 = _zz_8802;
  assign _zz_475 = 1'b1;
  assign _zz_2809 = _zz_8810;
  assign _zz_2810 = _zz_8818;
  assign _zz_478 = ($signed(_zz_8826) * $signed(data_mid_63_real));
  assign _zz_2811 = _zz_8827;
  assign _zz_476 = _zz_8830[31 : 0];
  assign _zz_2812 = _zz_8831;
  assign _zz_477 = _zz_8834[31 : 0];
  assign _zz_479 = 1'b1;
  assign _zz_2813 = _zz_8835;
  assign _zz_2814 = _zz_8843;
  assign _zz_480 = 1'b1;
  assign _zz_2815 = _zz_8851;
  assign _zz_2816 = _zz_8859;
  assign _zz_483 = ($signed(_zz_8867) * $signed(data_mid_66_real));
  assign _zz_2817 = _zz_8868;
  assign _zz_481 = _zz_8871[31 : 0];
  assign _zz_2818 = _zz_8872;
  assign _zz_482 = _zz_8875[31 : 0];
  assign _zz_484 = 1'b1;
  assign _zz_2819 = _zz_8876;
  assign _zz_2820 = _zz_8884;
  assign _zz_485 = 1'b1;
  assign _zz_2821 = _zz_8892;
  assign _zz_2822 = _zz_8900;
  assign _zz_488 = ($signed(_zz_8908) * $signed(data_mid_67_real));
  assign _zz_2823 = _zz_8909;
  assign _zz_486 = _zz_8912[31 : 0];
  assign _zz_2824 = _zz_8913;
  assign _zz_487 = _zz_8916[31 : 0];
  assign _zz_489 = 1'b1;
  assign _zz_2825 = _zz_8917;
  assign _zz_2826 = _zz_8925;
  assign _zz_490 = 1'b1;
  assign _zz_2827 = _zz_8933;
  assign _zz_2828 = _zz_8941;
  assign _zz_493 = ($signed(_zz_8949) * $signed(data_mid_70_real));
  assign _zz_2829 = _zz_8950;
  assign _zz_491 = _zz_8953[31 : 0];
  assign _zz_2830 = _zz_8954;
  assign _zz_492 = _zz_8957[31 : 0];
  assign _zz_494 = 1'b1;
  assign _zz_2831 = _zz_8958;
  assign _zz_2832 = _zz_8966;
  assign _zz_495 = 1'b1;
  assign _zz_2833 = _zz_8974;
  assign _zz_2834 = _zz_8982;
  assign _zz_498 = ($signed(_zz_8990) * $signed(data_mid_71_real));
  assign _zz_2835 = _zz_8991;
  assign _zz_496 = _zz_8994[31 : 0];
  assign _zz_2836 = _zz_8995;
  assign _zz_497 = _zz_8998[31 : 0];
  assign _zz_499 = 1'b1;
  assign _zz_2837 = _zz_8999;
  assign _zz_2838 = _zz_9007;
  assign _zz_500 = 1'b1;
  assign _zz_2839 = _zz_9015;
  assign _zz_2840 = _zz_9023;
  assign _zz_503 = ($signed(_zz_9031) * $signed(data_mid_74_real));
  assign _zz_2841 = _zz_9032;
  assign _zz_501 = _zz_9035[31 : 0];
  assign _zz_2842 = _zz_9036;
  assign _zz_502 = _zz_9039[31 : 0];
  assign _zz_504 = 1'b1;
  assign _zz_2843 = _zz_9040;
  assign _zz_2844 = _zz_9048;
  assign _zz_505 = 1'b1;
  assign _zz_2845 = _zz_9056;
  assign _zz_2846 = _zz_9064;
  assign _zz_508 = ($signed(_zz_9072) * $signed(data_mid_75_real));
  assign _zz_2847 = _zz_9073;
  assign _zz_506 = _zz_9076[31 : 0];
  assign _zz_2848 = _zz_9077;
  assign _zz_507 = _zz_9080[31 : 0];
  assign _zz_509 = 1'b1;
  assign _zz_2849 = _zz_9081;
  assign _zz_2850 = _zz_9089;
  assign _zz_510 = 1'b1;
  assign _zz_2851 = _zz_9097;
  assign _zz_2852 = _zz_9105;
  assign _zz_513 = ($signed(_zz_9113) * $signed(data_mid_78_real));
  assign _zz_2853 = _zz_9114;
  assign _zz_511 = _zz_9117[31 : 0];
  assign _zz_2854 = _zz_9118;
  assign _zz_512 = _zz_9121[31 : 0];
  assign _zz_514 = 1'b1;
  assign _zz_2855 = _zz_9122;
  assign _zz_2856 = _zz_9130;
  assign _zz_515 = 1'b1;
  assign _zz_2857 = _zz_9138;
  assign _zz_2858 = _zz_9146;
  assign _zz_518 = ($signed(_zz_9154) * $signed(data_mid_79_real));
  assign _zz_2859 = _zz_9155;
  assign _zz_516 = _zz_9158[31 : 0];
  assign _zz_2860 = _zz_9159;
  assign _zz_517 = _zz_9162[31 : 0];
  assign _zz_519 = 1'b1;
  assign _zz_2861 = _zz_9163;
  assign _zz_2862 = _zz_9171;
  assign _zz_520 = 1'b1;
  assign _zz_2863 = _zz_9179;
  assign _zz_2864 = _zz_9187;
  assign _zz_523 = ($signed(_zz_9195) * $signed(data_mid_82_real));
  assign _zz_2865 = _zz_9196;
  assign _zz_521 = _zz_9199[31 : 0];
  assign _zz_2866 = _zz_9200;
  assign _zz_522 = _zz_9203[31 : 0];
  assign _zz_524 = 1'b1;
  assign _zz_2867 = _zz_9204;
  assign _zz_2868 = _zz_9212;
  assign _zz_525 = 1'b1;
  assign _zz_2869 = _zz_9220;
  assign _zz_2870 = _zz_9228;
  assign _zz_528 = ($signed(_zz_9236) * $signed(data_mid_83_real));
  assign _zz_2871 = _zz_9237;
  assign _zz_526 = _zz_9240[31 : 0];
  assign _zz_2872 = _zz_9241;
  assign _zz_527 = _zz_9244[31 : 0];
  assign _zz_529 = 1'b1;
  assign _zz_2873 = _zz_9245;
  assign _zz_2874 = _zz_9253;
  assign _zz_530 = 1'b1;
  assign _zz_2875 = _zz_9261;
  assign _zz_2876 = _zz_9269;
  assign _zz_533 = ($signed(_zz_9277) * $signed(data_mid_86_real));
  assign _zz_2877 = _zz_9278;
  assign _zz_531 = _zz_9281[31 : 0];
  assign _zz_2878 = _zz_9282;
  assign _zz_532 = _zz_9285[31 : 0];
  assign _zz_534 = 1'b1;
  assign _zz_2879 = _zz_9286;
  assign _zz_2880 = _zz_9294;
  assign _zz_535 = 1'b1;
  assign _zz_2881 = _zz_9302;
  assign _zz_2882 = _zz_9310;
  assign _zz_538 = ($signed(_zz_9318) * $signed(data_mid_87_real));
  assign _zz_2883 = _zz_9319;
  assign _zz_536 = _zz_9322[31 : 0];
  assign _zz_2884 = _zz_9323;
  assign _zz_537 = _zz_9326[31 : 0];
  assign _zz_539 = 1'b1;
  assign _zz_2885 = _zz_9327;
  assign _zz_2886 = _zz_9335;
  assign _zz_540 = 1'b1;
  assign _zz_2887 = _zz_9343;
  assign _zz_2888 = _zz_9351;
  assign _zz_543 = ($signed(_zz_9359) * $signed(data_mid_90_real));
  assign _zz_2889 = _zz_9360;
  assign _zz_541 = _zz_9363[31 : 0];
  assign _zz_2890 = _zz_9364;
  assign _zz_542 = _zz_9367[31 : 0];
  assign _zz_544 = 1'b1;
  assign _zz_2891 = _zz_9368;
  assign _zz_2892 = _zz_9376;
  assign _zz_545 = 1'b1;
  assign _zz_2893 = _zz_9384;
  assign _zz_2894 = _zz_9392;
  assign _zz_548 = ($signed(_zz_9400) * $signed(data_mid_91_real));
  assign _zz_2895 = _zz_9401;
  assign _zz_546 = _zz_9404[31 : 0];
  assign _zz_2896 = _zz_9405;
  assign _zz_547 = _zz_9408[31 : 0];
  assign _zz_549 = 1'b1;
  assign _zz_2897 = _zz_9409;
  assign _zz_2898 = _zz_9417;
  assign _zz_550 = 1'b1;
  assign _zz_2899 = _zz_9425;
  assign _zz_2900 = _zz_9433;
  assign _zz_553 = ($signed(_zz_9441) * $signed(data_mid_94_real));
  assign _zz_2901 = _zz_9442;
  assign _zz_551 = _zz_9445[31 : 0];
  assign _zz_2902 = _zz_9446;
  assign _zz_552 = _zz_9449[31 : 0];
  assign _zz_554 = 1'b1;
  assign _zz_2903 = _zz_9450;
  assign _zz_2904 = _zz_9458;
  assign _zz_555 = 1'b1;
  assign _zz_2905 = _zz_9466;
  assign _zz_2906 = _zz_9474;
  assign _zz_558 = ($signed(_zz_9482) * $signed(data_mid_95_real));
  assign _zz_2907 = _zz_9483;
  assign _zz_556 = _zz_9486[31 : 0];
  assign _zz_2908 = _zz_9487;
  assign _zz_557 = _zz_9490[31 : 0];
  assign _zz_559 = 1'b1;
  assign _zz_2909 = _zz_9491;
  assign _zz_2910 = _zz_9499;
  assign _zz_560 = 1'b1;
  assign _zz_2911 = _zz_9507;
  assign _zz_2912 = _zz_9515;
  assign _zz_563 = ($signed(_zz_9523) * $signed(data_mid_98_real));
  assign _zz_2913 = _zz_9524;
  assign _zz_561 = _zz_9527[31 : 0];
  assign _zz_2914 = _zz_9528;
  assign _zz_562 = _zz_9531[31 : 0];
  assign _zz_564 = 1'b1;
  assign _zz_2915 = _zz_9532;
  assign _zz_2916 = _zz_9540;
  assign _zz_565 = 1'b1;
  assign _zz_2917 = _zz_9548;
  assign _zz_2918 = _zz_9556;
  assign _zz_568 = ($signed(_zz_9564) * $signed(data_mid_99_real));
  assign _zz_2919 = _zz_9565;
  assign _zz_566 = _zz_9568[31 : 0];
  assign _zz_2920 = _zz_9569;
  assign _zz_567 = _zz_9572[31 : 0];
  assign _zz_569 = 1'b1;
  assign _zz_2921 = _zz_9573;
  assign _zz_2922 = _zz_9581;
  assign _zz_570 = 1'b1;
  assign _zz_2923 = _zz_9589;
  assign _zz_2924 = _zz_9597;
  assign _zz_573 = ($signed(_zz_9605) * $signed(data_mid_102_real));
  assign _zz_2925 = _zz_9606;
  assign _zz_571 = _zz_9609[31 : 0];
  assign _zz_2926 = _zz_9610;
  assign _zz_572 = _zz_9613[31 : 0];
  assign _zz_574 = 1'b1;
  assign _zz_2927 = _zz_9614;
  assign _zz_2928 = _zz_9622;
  assign _zz_575 = 1'b1;
  assign _zz_2929 = _zz_9630;
  assign _zz_2930 = _zz_9638;
  assign _zz_578 = ($signed(_zz_9646) * $signed(data_mid_103_real));
  assign _zz_2931 = _zz_9647;
  assign _zz_576 = _zz_9650[31 : 0];
  assign _zz_2932 = _zz_9651;
  assign _zz_577 = _zz_9654[31 : 0];
  assign _zz_579 = 1'b1;
  assign _zz_2933 = _zz_9655;
  assign _zz_2934 = _zz_9663;
  assign _zz_580 = 1'b1;
  assign _zz_2935 = _zz_9671;
  assign _zz_2936 = _zz_9679;
  assign _zz_583 = ($signed(_zz_9687) * $signed(data_mid_106_real));
  assign _zz_2937 = _zz_9688;
  assign _zz_581 = _zz_9691[31 : 0];
  assign _zz_2938 = _zz_9692;
  assign _zz_582 = _zz_9695[31 : 0];
  assign _zz_584 = 1'b1;
  assign _zz_2939 = _zz_9696;
  assign _zz_2940 = _zz_9704;
  assign _zz_585 = 1'b1;
  assign _zz_2941 = _zz_9712;
  assign _zz_2942 = _zz_9720;
  assign _zz_588 = ($signed(_zz_9728) * $signed(data_mid_107_real));
  assign _zz_2943 = _zz_9729;
  assign _zz_586 = _zz_9732[31 : 0];
  assign _zz_2944 = _zz_9733;
  assign _zz_587 = _zz_9736[31 : 0];
  assign _zz_589 = 1'b1;
  assign _zz_2945 = _zz_9737;
  assign _zz_2946 = _zz_9745;
  assign _zz_590 = 1'b1;
  assign _zz_2947 = _zz_9753;
  assign _zz_2948 = _zz_9761;
  assign _zz_593 = ($signed(_zz_9769) * $signed(data_mid_110_real));
  assign _zz_2949 = _zz_9770;
  assign _zz_591 = _zz_9773[31 : 0];
  assign _zz_2950 = _zz_9774;
  assign _zz_592 = _zz_9777[31 : 0];
  assign _zz_594 = 1'b1;
  assign _zz_2951 = _zz_9778;
  assign _zz_2952 = _zz_9786;
  assign _zz_595 = 1'b1;
  assign _zz_2953 = _zz_9794;
  assign _zz_2954 = _zz_9802;
  assign _zz_598 = ($signed(_zz_9810) * $signed(data_mid_111_real));
  assign _zz_2955 = _zz_9811;
  assign _zz_596 = _zz_9814[31 : 0];
  assign _zz_2956 = _zz_9815;
  assign _zz_597 = _zz_9818[31 : 0];
  assign _zz_599 = 1'b1;
  assign _zz_2957 = _zz_9819;
  assign _zz_2958 = _zz_9827;
  assign _zz_600 = 1'b1;
  assign _zz_2959 = _zz_9835;
  assign _zz_2960 = _zz_9843;
  assign _zz_603 = ($signed(_zz_9851) * $signed(data_mid_114_real));
  assign _zz_2961 = _zz_9852;
  assign _zz_601 = _zz_9855[31 : 0];
  assign _zz_2962 = _zz_9856;
  assign _zz_602 = _zz_9859[31 : 0];
  assign _zz_604 = 1'b1;
  assign _zz_2963 = _zz_9860;
  assign _zz_2964 = _zz_9868;
  assign _zz_605 = 1'b1;
  assign _zz_2965 = _zz_9876;
  assign _zz_2966 = _zz_9884;
  assign _zz_608 = ($signed(_zz_9892) * $signed(data_mid_115_real));
  assign _zz_2967 = _zz_9893;
  assign _zz_606 = _zz_9896[31 : 0];
  assign _zz_2968 = _zz_9897;
  assign _zz_607 = _zz_9900[31 : 0];
  assign _zz_609 = 1'b1;
  assign _zz_2969 = _zz_9901;
  assign _zz_2970 = _zz_9909;
  assign _zz_610 = 1'b1;
  assign _zz_2971 = _zz_9917;
  assign _zz_2972 = _zz_9925;
  assign _zz_613 = ($signed(_zz_9933) * $signed(data_mid_118_real));
  assign _zz_2973 = _zz_9934;
  assign _zz_611 = _zz_9937[31 : 0];
  assign _zz_2974 = _zz_9938;
  assign _zz_612 = _zz_9941[31 : 0];
  assign _zz_614 = 1'b1;
  assign _zz_2975 = _zz_9942;
  assign _zz_2976 = _zz_9950;
  assign _zz_615 = 1'b1;
  assign _zz_2977 = _zz_9958;
  assign _zz_2978 = _zz_9966;
  assign _zz_618 = ($signed(_zz_9974) * $signed(data_mid_119_real));
  assign _zz_2979 = _zz_9975;
  assign _zz_616 = _zz_9978[31 : 0];
  assign _zz_2980 = _zz_9979;
  assign _zz_617 = _zz_9982[31 : 0];
  assign _zz_619 = 1'b1;
  assign _zz_2981 = _zz_9983;
  assign _zz_2982 = _zz_9991;
  assign _zz_620 = 1'b1;
  assign _zz_2983 = _zz_9999;
  assign _zz_2984 = _zz_10007;
  assign _zz_623 = ($signed(_zz_10015) * $signed(data_mid_122_real));
  assign _zz_2985 = _zz_10016;
  assign _zz_621 = _zz_10019[31 : 0];
  assign _zz_2986 = _zz_10020;
  assign _zz_622 = _zz_10023[31 : 0];
  assign _zz_624 = 1'b1;
  assign _zz_2987 = _zz_10024;
  assign _zz_2988 = _zz_10032;
  assign _zz_625 = 1'b1;
  assign _zz_2989 = _zz_10040;
  assign _zz_2990 = _zz_10048;
  assign _zz_628 = ($signed(_zz_10056) * $signed(data_mid_123_real));
  assign _zz_2991 = _zz_10057;
  assign _zz_626 = _zz_10060[31 : 0];
  assign _zz_2992 = _zz_10061;
  assign _zz_627 = _zz_10064[31 : 0];
  assign _zz_629 = 1'b1;
  assign _zz_2993 = _zz_10065;
  assign _zz_2994 = _zz_10073;
  assign _zz_630 = 1'b1;
  assign _zz_2995 = _zz_10081;
  assign _zz_2996 = _zz_10089;
  assign _zz_633 = ($signed(_zz_10097) * $signed(data_mid_126_real));
  assign _zz_2997 = _zz_10098;
  assign _zz_631 = _zz_10101[31 : 0];
  assign _zz_2998 = _zz_10102;
  assign _zz_632 = _zz_10105[31 : 0];
  assign _zz_634 = 1'b1;
  assign _zz_2999 = _zz_10106;
  assign _zz_3000 = _zz_10114;
  assign _zz_635 = 1'b1;
  assign _zz_3001 = _zz_10122;
  assign _zz_3002 = _zz_10130;
  assign _zz_638 = ($signed(_zz_10138) * $signed(data_mid_127_real));
  assign _zz_3003 = _zz_10139;
  assign _zz_636 = _zz_10142[31 : 0];
  assign _zz_3004 = _zz_10143;
  assign _zz_637 = _zz_10146[31 : 0];
  assign _zz_639 = 1'b1;
  assign _zz_3005 = _zz_10147;
  assign _zz_3006 = _zz_10155;
  assign _zz_640 = 1'b1;
  assign _zz_3007 = _zz_10163;
  assign _zz_3008 = _zz_10171;
  assign _zz_643 = ($signed(_zz_10179) * $signed(data_mid_4_real));
  assign _zz_3009 = _zz_10180;
  assign _zz_641 = _zz_10183[31 : 0];
  assign _zz_3010 = _zz_10184;
  assign _zz_642 = _zz_10187[31 : 0];
  assign _zz_644 = 1'b1;
  assign _zz_3011 = _zz_10188;
  assign _zz_3012 = _zz_10196;
  assign _zz_645 = 1'b1;
  assign _zz_3013 = _zz_10204;
  assign _zz_3014 = _zz_10212;
  assign _zz_648 = ($signed(_zz_10220) * $signed(data_mid_5_real));
  assign _zz_3015 = _zz_10221;
  assign _zz_646 = _zz_10224[31 : 0];
  assign _zz_3016 = _zz_10225;
  assign _zz_647 = _zz_10228[31 : 0];
  assign _zz_649 = 1'b1;
  assign _zz_3017 = _zz_10229;
  assign _zz_3018 = _zz_10237;
  assign _zz_650 = 1'b1;
  assign _zz_3019 = _zz_10245;
  assign _zz_3020 = _zz_10253;
  assign _zz_653 = ($signed(_zz_10261) * $signed(data_mid_6_real));
  assign _zz_3021 = _zz_10262;
  assign _zz_651 = _zz_10265[31 : 0];
  assign _zz_3022 = _zz_10266;
  assign _zz_652 = _zz_10269[31 : 0];
  assign _zz_654 = 1'b1;
  assign _zz_3023 = _zz_10270;
  assign _zz_3024 = _zz_10278;
  assign _zz_655 = 1'b1;
  assign _zz_3025 = _zz_10286;
  assign _zz_3026 = _zz_10294;
  assign _zz_658 = ($signed(_zz_10302) * $signed(data_mid_7_real));
  assign _zz_3027 = _zz_10303;
  assign _zz_656 = _zz_10306[31 : 0];
  assign _zz_3028 = _zz_10307;
  assign _zz_657 = _zz_10310[31 : 0];
  assign _zz_659 = 1'b1;
  assign _zz_3029 = _zz_10311;
  assign _zz_3030 = _zz_10319;
  assign _zz_660 = 1'b1;
  assign _zz_3031 = _zz_10327;
  assign _zz_3032 = _zz_10335;
  assign _zz_663 = ($signed(_zz_10343) * $signed(data_mid_12_real));
  assign _zz_3033 = _zz_10344;
  assign _zz_661 = _zz_10347[31 : 0];
  assign _zz_3034 = _zz_10348;
  assign _zz_662 = _zz_10351[31 : 0];
  assign _zz_664 = 1'b1;
  assign _zz_3035 = _zz_10352;
  assign _zz_3036 = _zz_10360;
  assign _zz_665 = 1'b1;
  assign _zz_3037 = _zz_10368;
  assign _zz_3038 = _zz_10376;
  assign _zz_668 = ($signed(_zz_10384) * $signed(data_mid_13_real));
  assign _zz_3039 = _zz_10385;
  assign _zz_666 = _zz_10388[31 : 0];
  assign _zz_3040 = _zz_10389;
  assign _zz_667 = _zz_10392[31 : 0];
  assign _zz_669 = 1'b1;
  assign _zz_3041 = _zz_10393;
  assign _zz_3042 = _zz_10401;
  assign _zz_670 = 1'b1;
  assign _zz_3043 = _zz_10409;
  assign _zz_3044 = _zz_10417;
  assign _zz_673 = ($signed(_zz_10425) * $signed(data_mid_14_real));
  assign _zz_3045 = _zz_10426;
  assign _zz_671 = _zz_10429[31 : 0];
  assign _zz_3046 = _zz_10430;
  assign _zz_672 = _zz_10433[31 : 0];
  assign _zz_674 = 1'b1;
  assign _zz_3047 = _zz_10434;
  assign _zz_3048 = _zz_10442;
  assign _zz_675 = 1'b1;
  assign _zz_3049 = _zz_10450;
  assign _zz_3050 = _zz_10458;
  assign _zz_678 = ($signed(_zz_10466) * $signed(data_mid_15_real));
  assign _zz_3051 = _zz_10467;
  assign _zz_676 = _zz_10470[31 : 0];
  assign _zz_3052 = _zz_10471;
  assign _zz_677 = _zz_10474[31 : 0];
  assign _zz_679 = 1'b1;
  assign _zz_3053 = _zz_10475;
  assign _zz_3054 = _zz_10483;
  assign _zz_680 = 1'b1;
  assign _zz_3055 = _zz_10491;
  assign _zz_3056 = _zz_10499;
  assign _zz_683 = ($signed(_zz_10507) * $signed(data_mid_20_real));
  assign _zz_3057 = _zz_10508;
  assign _zz_681 = _zz_10511[31 : 0];
  assign _zz_3058 = _zz_10512;
  assign _zz_682 = _zz_10515[31 : 0];
  assign _zz_684 = 1'b1;
  assign _zz_3059 = _zz_10516;
  assign _zz_3060 = _zz_10524;
  assign _zz_685 = 1'b1;
  assign _zz_3061 = _zz_10532;
  assign _zz_3062 = _zz_10540;
  assign _zz_688 = ($signed(_zz_10548) * $signed(data_mid_21_real));
  assign _zz_3063 = _zz_10549;
  assign _zz_686 = _zz_10552[31 : 0];
  assign _zz_3064 = _zz_10553;
  assign _zz_687 = _zz_10556[31 : 0];
  assign _zz_689 = 1'b1;
  assign _zz_3065 = _zz_10557;
  assign _zz_3066 = _zz_10565;
  assign _zz_690 = 1'b1;
  assign _zz_3067 = _zz_10573;
  assign _zz_3068 = _zz_10581;
  assign _zz_693 = ($signed(_zz_10589) * $signed(data_mid_22_real));
  assign _zz_3069 = _zz_10590;
  assign _zz_691 = _zz_10593[31 : 0];
  assign _zz_3070 = _zz_10594;
  assign _zz_692 = _zz_10597[31 : 0];
  assign _zz_694 = 1'b1;
  assign _zz_3071 = _zz_10598;
  assign _zz_3072 = _zz_10606;
  assign _zz_695 = 1'b1;
  assign _zz_3073 = _zz_10614;
  assign _zz_3074 = _zz_10622;
  assign _zz_698 = ($signed(_zz_10630) * $signed(data_mid_23_real));
  assign _zz_3075 = _zz_10631;
  assign _zz_696 = _zz_10634[31 : 0];
  assign _zz_3076 = _zz_10635;
  assign _zz_697 = _zz_10638[31 : 0];
  assign _zz_699 = 1'b1;
  assign _zz_3077 = _zz_10639;
  assign _zz_3078 = _zz_10647;
  assign _zz_700 = 1'b1;
  assign _zz_3079 = _zz_10655;
  assign _zz_3080 = _zz_10663;
  assign _zz_703 = ($signed(_zz_10671) * $signed(data_mid_28_real));
  assign _zz_3081 = _zz_10672;
  assign _zz_701 = _zz_10675[31 : 0];
  assign _zz_3082 = _zz_10676;
  assign _zz_702 = _zz_10679[31 : 0];
  assign _zz_704 = 1'b1;
  assign _zz_3083 = _zz_10680;
  assign _zz_3084 = _zz_10688;
  assign _zz_705 = 1'b1;
  assign _zz_3085 = _zz_10696;
  assign _zz_3086 = _zz_10704;
  assign _zz_708 = ($signed(_zz_10712) * $signed(data_mid_29_real));
  assign _zz_3087 = _zz_10713;
  assign _zz_706 = _zz_10716[31 : 0];
  assign _zz_3088 = _zz_10717;
  assign _zz_707 = _zz_10720[31 : 0];
  assign _zz_709 = 1'b1;
  assign _zz_3089 = _zz_10721;
  assign _zz_3090 = _zz_10729;
  assign _zz_710 = 1'b1;
  assign _zz_3091 = _zz_10737;
  assign _zz_3092 = _zz_10745;
  assign _zz_713 = ($signed(_zz_10753) * $signed(data_mid_30_real));
  assign _zz_3093 = _zz_10754;
  assign _zz_711 = _zz_10757[31 : 0];
  assign _zz_3094 = _zz_10758;
  assign _zz_712 = _zz_10761[31 : 0];
  assign _zz_714 = 1'b1;
  assign _zz_3095 = _zz_10762;
  assign _zz_3096 = _zz_10770;
  assign _zz_715 = 1'b1;
  assign _zz_3097 = _zz_10778;
  assign _zz_3098 = _zz_10786;
  assign _zz_718 = ($signed(_zz_10794) * $signed(data_mid_31_real));
  assign _zz_3099 = _zz_10795;
  assign _zz_716 = _zz_10798[31 : 0];
  assign _zz_3100 = _zz_10799;
  assign _zz_717 = _zz_10802[31 : 0];
  assign _zz_719 = 1'b1;
  assign _zz_3101 = _zz_10803;
  assign _zz_3102 = _zz_10811;
  assign _zz_720 = 1'b1;
  assign _zz_3103 = _zz_10819;
  assign _zz_3104 = _zz_10827;
  assign _zz_723 = ($signed(_zz_10835) * $signed(data_mid_36_real));
  assign _zz_3105 = _zz_10836;
  assign _zz_721 = _zz_10839[31 : 0];
  assign _zz_3106 = _zz_10840;
  assign _zz_722 = _zz_10843[31 : 0];
  assign _zz_724 = 1'b1;
  assign _zz_3107 = _zz_10844;
  assign _zz_3108 = _zz_10852;
  assign _zz_725 = 1'b1;
  assign _zz_3109 = _zz_10860;
  assign _zz_3110 = _zz_10868;
  assign _zz_728 = ($signed(_zz_10876) * $signed(data_mid_37_real));
  assign _zz_3111 = _zz_10877;
  assign _zz_726 = _zz_10880[31 : 0];
  assign _zz_3112 = _zz_10881;
  assign _zz_727 = _zz_10884[31 : 0];
  assign _zz_729 = 1'b1;
  assign _zz_3113 = _zz_10885;
  assign _zz_3114 = _zz_10893;
  assign _zz_730 = 1'b1;
  assign _zz_3115 = _zz_10901;
  assign _zz_3116 = _zz_10909;
  assign _zz_733 = ($signed(_zz_10917) * $signed(data_mid_38_real));
  assign _zz_3117 = _zz_10918;
  assign _zz_731 = _zz_10921[31 : 0];
  assign _zz_3118 = _zz_10922;
  assign _zz_732 = _zz_10925[31 : 0];
  assign _zz_734 = 1'b1;
  assign _zz_3119 = _zz_10926;
  assign _zz_3120 = _zz_10934;
  assign _zz_735 = 1'b1;
  assign _zz_3121 = _zz_10942;
  assign _zz_3122 = _zz_10950;
  assign _zz_738 = ($signed(_zz_10958) * $signed(data_mid_39_real));
  assign _zz_3123 = _zz_10959;
  assign _zz_736 = _zz_10962[31 : 0];
  assign _zz_3124 = _zz_10963;
  assign _zz_737 = _zz_10966[31 : 0];
  assign _zz_739 = 1'b1;
  assign _zz_3125 = _zz_10967;
  assign _zz_3126 = _zz_10975;
  assign _zz_740 = 1'b1;
  assign _zz_3127 = _zz_10983;
  assign _zz_3128 = _zz_10991;
  assign _zz_743 = ($signed(_zz_10999) * $signed(data_mid_44_real));
  assign _zz_3129 = _zz_11000;
  assign _zz_741 = _zz_11003[31 : 0];
  assign _zz_3130 = _zz_11004;
  assign _zz_742 = _zz_11007[31 : 0];
  assign _zz_744 = 1'b1;
  assign _zz_3131 = _zz_11008;
  assign _zz_3132 = _zz_11016;
  assign _zz_745 = 1'b1;
  assign _zz_3133 = _zz_11024;
  assign _zz_3134 = _zz_11032;
  assign _zz_748 = ($signed(_zz_11040) * $signed(data_mid_45_real));
  assign _zz_3135 = _zz_11041;
  assign _zz_746 = _zz_11044[31 : 0];
  assign _zz_3136 = _zz_11045;
  assign _zz_747 = _zz_11048[31 : 0];
  assign _zz_749 = 1'b1;
  assign _zz_3137 = _zz_11049;
  assign _zz_3138 = _zz_11057;
  assign _zz_750 = 1'b1;
  assign _zz_3139 = _zz_11065;
  assign _zz_3140 = _zz_11073;
  assign _zz_753 = ($signed(_zz_11081) * $signed(data_mid_46_real));
  assign _zz_3141 = _zz_11082;
  assign _zz_751 = _zz_11085[31 : 0];
  assign _zz_3142 = _zz_11086;
  assign _zz_752 = _zz_11089[31 : 0];
  assign _zz_754 = 1'b1;
  assign _zz_3143 = _zz_11090;
  assign _zz_3144 = _zz_11098;
  assign _zz_755 = 1'b1;
  assign _zz_3145 = _zz_11106;
  assign _zz_3146 = _zz_11114;
  assign _zz_758 = ($signed(_zz_11122) * $signed(data_mid_47_real));
  assign _zz_3147 = _zz_11123;
  assign _zz_756 = _zz_11126[31 : 0];
  assign _zz_3148 = _zz_11127;
  assign _zz_757 = _zz_11130[31 : 0];
  assign _zz_759 = 1'b1;
  assign _zz_3149 = _zz_11131;
  assign _zz_3150 = _zz_11139;
  assign _zz_760 = 1'b1;
  assign _zz_3151 = _zz_11147;
  assign _zz_3152 = _zz_11155;
  assign _zz_763 = ($signed(_zz_11163) * $signed(data_mid_52_real));
  assign _zz_3153 = _zz_11164;
  assign _zz_761 = _zz_11167[31 : 0];
  assign _zz_3154 = _zz_11168;
  assign _zz_762 = _zz_11171[31 : 0];
  assign _zz_764 = 1'b1;
  assign _zz_3155 = _zz_11172;
  assign _zz_3156 = _zz_11180;
  assign _zz_765 = 1'b1;
  assign _zz_3157 = _zz_11188;
  assign _zz_3158 = _zz_11196;
  assign _zz_768 = ($signed(_zz_11204) * $signed(data_mid_53_real));
  assign _zz_3159 = _zz_11205;
  assign _zz_766 = _zz_11208[31 : 0];
  assign _zz_3160 = _zz_11209;
  assign _zz_767 = _zz_11212[31 : 0];
  assign _zz_769 = 1'b1;
  assign _zz_3161 = _zz_11213;
  assign _zz_3162 = _zz_11221;
  assign _zz_770 = 1'b1;
  assign _zz_3163 = _zz_11229;
  assign _zz_3164 = _zz_11237;
  assign _zz_773 = ($signed(_zz_11245) * $signed(data_mid_54_real));
  assign _zz_3165 = _zz_11246;
  assign _zz_771 = _zz_11249[31 : 0];
  assign _zz_3166 = _zz_11250;
  assign _zz_772 = _zz_11253[31 : 0];
  assign _zz_774 = 1'b1;
  assign _zz_3167 = _zz_11254;
  assign _zz_3168 = _zz_11262;
  assign _zz_775 = 1'b1;
  assign _zz_3169 = _zz_11270;
  assign _zz_3170 = _zz_11278;
  assign _zz_778 = ($signed(_zz_11286) * $signed(data_mid_55_real));
  assign _zz_3171 = _zz_11287;
  assign _zz_776 = _zz_11290[31 : 0];
  assign _zz_3172 = _zz_11291;
  assign _zz_777 = _zz_11294[31 : 0];
  assign _zz_779 = 1'b1;
  assign _zz_3173 = _zz_11295;
  assign _zz_3174 = _zz_11303;
  assign _zz_780 = 1'b1;
  assign _zz_3175 = _zz_11311;
  assign _zz_3176 = _zz_11319;
  assign _zz_783 = ($signed(_zz_11327) * $signed(data_mid_60_real));
  assign _zz_3177 = _zz_11328;
  assign _zz_781 = _zz_11331[31 : 0];
  assign _zz_3178 = _zz_11332;
  assign _zz_782 = _zz_11335[31 : 0];
  assign _zz_784 = 1'b1;
  assign _zz_3179 = _zz_11336;
  assign _zz_3180 = _zz_11344;
  assign _zz_785 = 1'b1;
  assign _zz_3181 = _zz_11352;
  assign _zz_3182 = _zz_11360;
  assign _zz_788 = ($signed(_zz_11368) * $signed(data_mid_61_real));
  assign _zz_3183 = _zz_11369;
  assign _zz_786 = _zz_11372[31 : 0];
  assign _zz_3184 = _zz_11373;
  assign _zz_787 = _zz_11376[31 : 0];
  assign _zz_789 = 1'b1;
  assign _zz_3185 = _zz_11377;
  assign _zz_3186 = _zz_11385;
  assign _zz_790 = 1'b1;
  assign _zz_3187 = _zz_11393;
  assign _zz_3188 = _zz_11401;
  assign _zz_793 = ($signed(_zz_11409) * $signed(data_mid_62_real));
  assign _zz_3189 = _zz_11410;
  assign _zz_791 = _zz_11413[31 : 0];
  assign _zz_3190 = _zz_11414;
  assign _zz_792 = _zz_11417[31 : 0];
  assign _zz_794 = 1'b1;
  assign _zz_3191 = _zz_11418;
  assign _zz_3192 = _zz_11426;
  assign _zz_795 = 1'b1;
  assign _zz_3193 = _zz_11434;
  assign _zz_3194 = _zz_11442;
  assign _zz_798 = ($signed(_zz_11450) * $signed(data_mid_63_real));
  assign _zz_3195 = _zz_11451;
  assign _zz_796 = _zz_11454[31 : 0];
  assign _zz_3196 = _zz_11455;
  assign _zz_797 = _zz_11458[31 : 0];
  assign _zz_799 = 1'b1;
  assign _zz_3197 = _zz_11459;
  assign _zz_3198 = _zz_11467;
  assign _zz_800 = 1'b1;
  assign _zz_3199 = _zz_11475;
  assign _zz_3200 = _zz_11483;
  assign _zz_803 = ($signed(_zz_11491) * $signed(data_mid_68_real));
  assign _zz_3201 = _zz_11492;
  assign _zz_801 = _zz_11495[31 : 0];
  assign _zz_3202 = _zz_11496;
  assign _zz_802 = _zz_11499[31 : 0];
  assign _zz_804 = 1'b1;
  assign _zz_3203 = _zz_11500;
  assign _zz_3204 = _zz_11508;
  assign _zz_805 = 1'b1;
  assign _zz_3205 = _zz_11516;
  assign _zz_3206 = _zz_11524;
  assign _zz_808 = ($signed(_zz_11532) * $signed(data_mid_69_real));
  assign _zz_3207 = _zz_11533;
  assign _zz_806 = _zz_11536[31 : 0];
  assign _zz_3208 = _zz_11537;
  assign _zz_807 = _zz_11540[31 : 0];
  assign _zz_809 = 1'b1;
  assign _zz_3209 = _zz_11541;
  assign _zz_3210 = _zz_11549;
  assign _zz_810 = 1'b1;
  assign _zz_3211 = _zz_11557;
  assign _zz_3212 = _zz_11565;
  assign _zz_813 = ($signed(_zz_11573) * $signed(data_mid_70_real));
  assign _zz_3213 = _zz_11574;
  assign _zz_811 = _zz_11577[31 : 0];
  assign _zz_3214 = _zz_11578;
  assign _zz_812 = _zz_11581[31 : 0];
  assign _zz_814 = 1'b1;
  assign _zz_3215 = _zz_11582;
  assign _zz_3216 = _zz_11590;
  assign _zz_815 = 1'b1;
  assign _zz_3217 = _zz_11598;
  assign _zz_3218 = _zz_11606;
  assign _zz_818 = ($signed(_zz_11614) * $signed(data_mid_71_real));
  assign _zz_3219 = _zz_11615;
  assign _zz_816 = _zz_11618[31 : 0];
  assign _zz_3220 = _zz_11619;
  assign _zz_817 = _zz_11622[31 : 0];
  assign _zz_819 = 1'b1;
  assign _zz_3221 = _zz_11623;
  assign _zz_3222 = _zz_11631;
  assign _zz_820 = 1'b1;
  assign _zz_3223 = _zz_11639;
  assign _zz_3224 = _zz_11647;
  assign _zz_823 = ($signed(_zz_11655) * $signed(data_mid_76_real));
  assign _zz_3225 = _zz_11656;
  assign _zz_821 = _zz_11659[31 : 0];
  assign _zz_3226 = _zz_11660;
  assign _zz_822 = _zz_11663[31 : 0];
  assign _zz_824 = 1'b1;
  assign _zz_3227 = _zz_11664;
  assign _zz_3228 = _zz_11672;
  assign _zz_825 = 1'b1;
  assign _zz_3229 = _zz_11680;
  assign _zz_3230 = _zz_11688;
  assign _zz_828 = ($signed(_zz_11696) * $signed(data_mid_77_real));
  assign _zz_3231 = _zz_11697;
  assign _zz_826 = _zz_11700[31 : 0];
  assign _zz_3232 = _zz_11701;
  assign _zz_827 = _zz_11704[31 : 0];
  assign _zz_829 = 1'b1;
  assign _zz_3233 = _zz_11705;
  assign _zz_3234 = _zz_11713;
  assign _zz_830 = 1'b1;
  assign _zz_3235 = _zz_11721;
  assign _zz_3236 = _zz_11729;
  assign _zz_833 = ($signed(_zz_11737) * $signed(data_mid_78_real));
  assign _zz_3237 = _zz_11738;
  assign _zz_831 = _zz_11741[31 : 0];
  assign _zz_3238 = _zz_11742;
  assign _zz_832 = _zz_11745[31 : 0];
  assign _zz_834 = 1'b1;
  assign _zz_3239 = _zz_11746;
  assign _zz_3240 = _zz_11754;
  assign _zz_835 = 1'b1;
  assign _zz_3241 = _zz_11762;
  assign _zz_3242 = _zz_11770;
  assign _zz_838 = ($signed(_zz_11778) * $signed(data_mid_79_real));
  assign _zz_3243 = _zz_11779;
  assign _zz_836 = _zz_11782[31 : 0];
  assign _zz_3244 = _zz_11783;
  assign _zz_837 = _zz_11786[31 : 0];
  assign _zz_839 = 1'b1;
  assign _zz_3245 = _zz_11787;
  assign _zz_3246 = _zz_11795;
  assign _zz_840 = 1'b1;
  assign _zz_3247 = _zz_11803;
  assign _zz_3248 = _zz_11811;
  assign _zz_843 = ($signed(_zz_11819) * $signed(data_mid_84_real));
  assign _zz_3249 = _zz_11820;
  assign _zz_841 = _zz_11823[31 : 0];
  assign _zz_3250 = _zz_11824;
  assign _zz_842 = _zz_11827[31 : 0];
  assign _zz_844 = 1'b1;
  assign _zz_3251 = _zz_11828;
  assign _zz_3252 = _zz_11836;
  assign _zz_845 = 1'b1;
  assign _zz_3253 = _zz_11844;
  assign _zz_3254 = _zz_11852;
  assign _zz_848 = ($signed(_zz_11860) * $signed(data_mid_85_real));
  assign _zz_3255 = _zz_11861;
  assign _zz_846 = _zz_11864[31 : 0];
  assign _zz_3256 = _zz_11865;
  assign _zz_847 = _zz_11868[31 : 0];
  assign _zz_849 = 1'b1;
  assign _zz_3257 = _zz_11869;
  assign _zz_3258 = _zz_11877;
  assign _zz_850 = 1'b1;
  assign _zz_3259 = _zz_11885;
  assign _zz_3260 = _zz_11893;
  assign _zz_853 = ($signed(_zz_11901) * $signed(data_mid_86_real));
  assign _zz_3261 = _zz_11902;
  assign _zz_851 = _zz_11905[31 : 0];
  assign _zz_3262 = _zz_11906;
  assign _zz_852 = _zz_11909[31 : 0];
  assign _zz_854 = 1'b1;
  assign _zz_3263 = _zz_11910;
  assign _zz_3264 = _zz_11918;
  assign _zz_855 = 1'b1;
  assign _zz_3265 = _zz_11926;
  assign _zz_3266 = _zz_11934;
  assign _zz_858 = ($signed(_zz_11942) * $signed(data_mid_87_real));
  assign _zz_3267 = _zz_11943;
  assign _zz_856 = _zz_11946[31 : 0];
  assign _zz_3268 = _zz_11947;
  assign _zz_857 = _zz_11950[31 : 0];
  assign _zz_859 = 1'b1;
  assign _zz_3269 = _zz_11951;
  assign _zz_3270 = _zz_11959;
  assign _zz_860 = 1'b1;
  assign _zz_3271 = _zz_11967;
  assign _zz_3272 = _zz_11975;
  assign _zz_863 = ($signed(_zz_11983) * $signed(data_mid_92_real));
  assign _zz_3273 = _zz_11984;
  assign _zz_861 = _zz_11987[31 : 0];
  assign _zz_3274 = _zz_11988;
  assign _zz_862 = _zz_11991[31 : 0];
  assign _zz_864 = 1'b1;
  assign _zz_3275 = _zz_11992;
  assign _zz_3276 = _zz_12000;
  assign _zz_865 = 1'b1;
  assign _zz_3277 = _zz_12008;
  assign _zz_3278 = _zz_12016;
  assign _zz_868 = ($signed(_zz_12024) * $signed(data_mid_93_real));
  assign _zz_3279 = _zz_12025;
  assign _zz_866 = _zz_12028[31 : 0];
  assign _zz_3280 = _zz_12029;
  assign _zz_867 = _zz_12032[31 : 0];
  assign _zz_869 = 1'b1;
  assign _zz_3281 = _zz_12033;
  assign _zz_3282 = _zz_12041;
  assign _zz_870 = 1'b1;
  assign _zz_3283 = _zz_12049;
  assign _zz_3284 = _zz_12057;
  assign _zz_873 = ($signed(_zz_12065) * $signed(data_mid_94_real));
  assign _zz_3285 = _zz_12066;
  assign _zz_871 = _zz_12069[31 : 0];
  assign _zz_3286 = _zz_12070;
  assign _zz_872 = _zz_12073[31 : 0];
  assign _zz_874 = 1'b1;
  assign _zz_3287 = _zz_12074;
  assign _zz_3288 = _zz_12082;
  assign _zz_875 = 1'b1;
  assign _zz_3289 = _zz_12090;
  assign _zz_3290 = _zz_12098;
  assign _zz_878 = ($signed(_zz_12106) * $signed(data_mid_95_real));
  assign _zz_3291 = _zz_12107;
  assign _zz_876 = _zz_12110[31 : 0];
  assign _zz_3292 = _zz_12111;
  assign _zz_877 = _zz_12114[31 : 0];
  assign _zz_879 = 1'b1;
  assign _zz_3293 = _zz_12115;
  assign _zz_3294 = _zz_12123;
  assign _zz_880 = 1'b1;
  assign _zz_3295 = _zz_12131;
  assign _zz_3296 = _zz_12139;
  assign _zz_883 = ($signed(_zz_12147) * $signed(data_mid_100_real));
  assign _zz_3297 = _zz_12148;
  assign _zz_881 = _zz_12151[31 : 0];
  assign _zz_3298 = _zz_12152;
  assign _zz_882 = _zz_12155[31 : 0];
  assign _zz_884 = 1'b1;
  assign _zz_3299 = _zz_12156;
  assign _zz_3300 = _zz_12164;
  assign _zz_885 = 1'b1;
  assign _zz_3301 = _zz_12172;
  assign _zz_3302 = _zz_12180;
  assign _zz_888 = ($signed(_zz_12188) * $signed(data_mid_101_real));
  assign _zz_3303 = _zz_12189;
  assign _zz_886 = _zz_12192[31 : 0];
  assign _zz_3304 = _zz_12193;
  assign _zz_887 = _zz_12196[31 : 0];
  assign _zz_889 = 1'b1;
  assign _zz_3305 = _zz_12197;
  assign _zz_3306 = _zz_12205;
  assign _zz_890 = 1'b1;
  assign _zz_3307 = _zz_12213;
  assign _zz_3308 = _zz_12221;
  assign _zz_893 = ($signed(_zz_12229) * $signed(data_mid_102_real));
  assign _zz_3309 = _zz_12230;
  assign _zz_891 = _zz_12233[31 : 0];
  assign _zz_3310 = _zz_12234;
  assign _zz_892 = _zz_12237[31 : 0];
  assign _zz_894 = 1'b1;
  assign _zz_3311 = _zz_12238;
  assign _zz_3312 = _zz_12246;
  assign _zz_895 = 1'b1;
  assign _zz_3313 = _zz_12254;
  assign _zz_3314 = _zz_12262;
  assign _zz_898 = ($signed(_zz_12270) * $signed(data_mid_103_real));
  assign _zz_3315 = _zz_12271;
  assign _zz_896 = _zz_12274[31 : 0];
  assign _zz_3316 = _zz_12275;
  assign _zz_897 = _zz_12278[31 : 0];
  assign _zz_899 = 1'b1;
  assign _zz_3317 = _zz_12279;
  assign _zz_3318 = _zz_12287;
  assign _zz_900 = 1'b1;
  assign _zz_3319 = _zz_12295;
  assign _zz_3320 = _zz_12303;
  assign _zz_903 = ($signed(_zz_12311) * $signed(data_mid_108_real));
  assign _zz_3321 = _zz_12312;
  assign _zz_901 = _zz_12315[31 : 0];
  assign _zz_3322 = _zz_12316;
  assign _zz_902 = _zz_12319[31 : 0];
  assign _zz_904 = 1'b1;
  assign _zz_3323 = _zz_12320;
  assign _zz_3324 = _zz_12328;
  assign _zz_905 = 1'b1;
  assign _zz_3325 = _zz_12336;
  assign _zz_3326 = _zz_12344;
  assign _zz_908 = ($signed(_zz_12352) * $signed(data_mid_109_real));
  assign _zz_3327 = _zz_12353;
  assign _zz_906 = _zz_12356[31 : 0];
  assign _zz_3328 = _zz_12357;
  assign _zz_907 = _zz_12360[31 : 0];
  assign _zz_909 = 1'b1;
  assign _zz_3329 = _zz_12361;
  assign _zz_3330 = _zz_12369;
  assign _zz_910 = 1'b1;
  assign _zz_3331 = _zz_12377;
  assign _zz_3332 = _zz_12385;
  assign _zz_913 = ($signed(_zz_12393) * $signed(data_mid_110_real));
  assign _zz_3333 = _zz_12394;
  assign _zz_911 = _zz_12397[31 : 0];
  assign _zz_3334 = _zz_12398;
  assign _zz_912 = _zz_12401[31 : 0];
  assign _zz_914 = 1'b1;
  assign _zz_3335 = _zz_12402;
  assign _zz_3336 = _zz_12410;
  assign _zz_915 = 1'b1;
  assign _zz_3337 = _zz_12418;
  assign _zz_3338 = _zz_12426;
  assign _zz_918 = ($signed(_zz_12434) * $signed(data_mid_111_real));
  assign _zz_3339 = _zz_12435;
  assign _zz_916 = _zz_12438[31 : 0];
  assign _zz_3340 = _zz_12439;
  assign _zz_917 = _zz_12442[31 : 0];
  assign _zz_919 = 1'b1;
  assign _zz_3341 = _zz_12443;
  assign _zz_3342 = _zz_12451;
  assign _zz_920 = 1'b1;
  assign _zz_3343 = _zz_12459;
  assign _zz_3344 = _zz_12467;
  assign _zz_923 = ($signed(_zz_12475) * $signed(data_mid_116_real));
  assign _zz_3345 = _zz_12476;
  assign _zz_921 = _zz_12479[31 : 0];
  assign _zz_3346 = _zz_12480;
  assign _zz_922 = _zz_12483[31 : 0];
  assign _zz_924 = 1'b1;
  assign _zz_3347 = _zz_12484;
  assign _zz_3348 = _zz_12492;
  assign _zz_925 = 1'b1;
  assign _zz_3349 = _zz_12500;
  assign _zz_3350 = _zz_12508;
  assign _zz_928 = ($signed(_zz_12516) * $signed(data_mid_117_real));
  assign _zz_3351 = _zz_12517;
  assign _zz_926 = _zz_12520[31 : 0];
  assign _zz_3352 = _zz_12521;
  assign _zz_927 = _zz_12524[31 : 0];
  assign _zz_929 = 1'b1;
  assign _zz_3353 = _zz_12525;
  assign _zz_3354 = _zz_12533;
  assign _zz_930 = 1'b1;
  assign _zz_3355 = _zz_12541;
  assign _zz_3356 = _zz_12549;
  assign _zz_933 = ($signed(_zz_12557) * $signed(data_mid_118_real));
  assign _zz_3357 = _zz_12558;
  assign _zz_931 = _zz_12561[31 : 0];
  assign _zz_3358 = _zz_12562;
  assign _zz_932 = _zz_12565[31 : 0];
  assign _zz_934 = 1'b1;
  assign _zz_3359 = _zz_12566;
  assign _zz_3360 = _zz_12574;
  assign _zz_935 = 1'b1;
  assign _zz_3361 = _zz_12582;
  assign _zz_3362 = _zz_12590;
  assign _zz_938 = ($signed(_zz_12598) * $signed(data_mid_119_real));
  assign _zz_3363 = _zz_12599;
  assign _zz_936 = _zz_12602[31 : 0];
  assign _zz_3364 = _zz_12603;
  assign _zz_937 = _zz_12606[31 : 0];
  assign _zz_939 = 1'b1;
  assign _zz_3365 = _zz_12607;
  assign _zz_3366 = _zz_12615;
  assign _zz_940 = 1'b1;
  assign _zz_3367 = _zz_12623;
  assign _zz_3368 = _zz_12631;
  assign _zz_943 = ($signed(_zz_12639) * $signed(data_mid_124_real));
  assign _zz_3369 = _zz_12640;
  assign _zz_941 = _zz_12643[31 : 0];
  assign _zz_3370 = _zz_12644;
  assign _zz_942 = _zz_12647[31 : 0];
  assign _zz_944 = 1'b1;
  assign _zz_3371 = _zz_12648;
  assign _zz_3372 = _zz_12656;
  assign _zz_945 = 1'b1;
  assign _zz_3373 = _zz_12664;
  assign _zz_3374 = _zz_12672;
  assign _zz_948 = ($signed(_zz_12680) * $signed(data_mid_125_real));
  assign _zz_3375 = _zz_12681;
  assign _zz_946 = _zz_12684[31 : 0];
  assign _zz_3376 = _zz_12685;
  assign _zz_947 = _zz_12688[31 : 0];
  assign _zz_949 = 1'b1;
  assign _zz_3377 = _zz_12689;
  assign _zz_3378 = _zz_12697;
  assign _zz_950 = 1'b1;
  assign _zz_3379 = _zz_12705;
  assign _zz_3380 = _zz_12713;
  assign _zz_953 = ($signed(_zz_12721) * $signed(data_mid_126_real));
  assign _zz_3381 = _zz_12722;
  assign _zz_951 = _zz_12725[31 : 0];
  assign _zz_3382 = _zz_12726;
  assign _zz_952 = _zz_12729[31 : 0];
  assign _zz_954 = 1'b1;
  assign _zz_3383 = _zz_12730;
  assign _zz_3384 = _zz_12738;
  assign _zz_955 = 1'b1;
  assign _zz_3385 = _zz_12746;
  assign _zz_3386 = _zz_12754;
  assign _zz_958 = ($signed(_zz_12762) * $signed(data_mid_127_real));
  assign _zz_3387 = _zz_12763;
  assign _zz_956 = _zz_12766[31 : 0];
  assign _zz_3388 = _zz_12767;
  assign _zz_957 = _zz_12770[31 : 0];
  assign _zz_959 = 1'b1;
  assign _zz_3389 = _zz_12771;
  assign _zz_3390 = _zz_12779;
  assign _zz_960 = 1'b1;
  assign _zz_3391 = _zz_12787;
  assign _zz_3392 = _zz_12795;
  assign _zz_963 = ($signed(_zz_12803) * $signed(data_mid_8_real));
  assign _zz_3393 = _zz_12804;
  assign _zz_961 = _zz_12807[31 : 0];
  assign _zz_3394 = _zz_12808;
  assign _zz_962 = _zz_12811[31 : 0];
  assign _zz_964 = 1'b1;
  assign _zz_3395 = _zz_12812;
  assign _zz_3396 = _zz_12820;
  assign _zz_965 = 1'b1;
  assign _zz_3397 = _zz_12828;
  assign _zz_3398 = _zz_12836;
  assign _zz_968 = ($signed(_zz_12844) * $signed(data_mid_9_real));
  assign _zz_3399 = _zz_12845;
  assign _zz_966 = _zz_12848[31 : 0];
  assign _zz_3400 = _zz_12849;
  assign _zz_967 = _zz_12852[31 : 0];
  assign _zz_969 = 1'b1;
  assign _zz_3401 = _zz_12853;
  assign _zz_3402 = _zz_12861;
  assign _zz_970 = 1'b1;
  assign _zz_3403 = _zz_12869;
  assign _zz_3404 = _zz_12877;
  assign _zz_973 = ($signed(_zz_12885) * $signed(data_mid_10_real));
  assign _zz_3405 = _zz_12886;
  assign _zz_971 = _zz_12889[31 : 0];
  assign _zz_3406 = _zz_12890;
  assign _zz_972 = _zz_12893[31 : 0];
  assign _zz_974 = 1'b1;
  assign _zz_3407 = _zz_12894;
  assign _zz_3408 = _zz_12902;
  assign _zz_975 = 1'b1;
  assign _zz_3409 = _zz_12910;
  assign _zz_3410 = _zz_12918;
  assign _zz_978 = ($signed(_zz_12926) * $signed(data_mid_11_real));
  assign _zz_3411 = _zz_12927;
  assign _zz_976 = _zz_12930[31 : 0];
  assign _zz_3412 = _zz_12931;
  assign _zz_977 = _zz_12934[31 : 0];
  assign _zz_979 = 1'b1;
  assign _zz_3413 = _zz_12935;
  assign _zz_3414 = _zz_12943;
  assign _zz_980 = 1'b1;
  assign _zz_3415 = _zz_12951;
  assign _zz_3416 = _zz_12959;
  assign _zz_983 = ($signed(_zz_12967) * $signed(data_mid_12_real));
  assign _zz_3417 = _zz_12968;
  assign _zz_981 = _zz_12971[31 : 0];
  assign _zz_3418 = _zz_12972;
  assign _zz_982 = _zz_12975[31 : 0];
  assign _zz_984 = 1'b1;
  assign _zz_3419 = _zz_12976;
  assign _zz_3420 = _zz_12984;
  assign _zz_985 = 1'b1;
  assign _zz_3421 = _zz_12992;
  assign _zz_3422 = _zz_13000;
  assign _zz_988 = ($signed(_zz_13008) * $signed(data_mid_13_real));
  assign _zz_3423 = _zz_13009;
  assign _zz_986 = _zz_13012[31 : 0];
  assign _zz_3424 = _zz_13013;
  assign _zz_987 = _zz_13016[31 : 0];
  assign _zz_989 = 1'b1;
  assign _zz_3425 = _zz_13017;
  assign _zz_3426 = _zz_13025;
  assign _zz_990 = 1'b1;
  assign _zz_3427 = _zz_13033;
  assign _zz_3428 = _zz_13041;
  assign _zz_993 = ($signed(_zz_13049) * $signed(data_mid_14_real));
  assign _zz_3429 = _zz_13050;
  assign _zz_991 = _zz_13053[31 : 0];
  assign _zz_3430 = _zz_13054;
  assign _zz_992 = _zz_13057[31 : 0];
  assign _zz_994 = 1'b1;
  assign _zz_3431 = _zz_13058;
  assign _zz_3432 = _zz_13066;
  assign _zz_995 = 1'b1;
  assign _zz_3433 = _zz_13074;
  assign _zz_3434 = _zz_13082;
  assign _zz_998 = ($signed(_zz_13090) * $signed(data_mid_15_real));
  assign _zz_3435 = _zz_13091;
  assign _zz_996 = _zz_13094[31 : 0];
  assign _zz_3436 = _zz_13095;
  assign _zz_997 = _zz_13098[31 : 0];
  assign _zz_999 = 1'b1;
  assign _zz_3437 = _zz_13099;
  assign _zz_3438 = _zz_13107;
  assign _zz_1000 = 1'b1;
  assign _zz_3439 = _zz_13115;
  assign _zz_3440 = _zz_13123;
  assign _zz_1003 = ($signed(_zz_13131) * $signed(data_mid_24_real));
  assign _zz_3441 = _zz_13132;
  assign _zz_1001 = _zz_13135[31 : 0];
  assign _zz_3442 = _zz_13136;
  assign _zz_1002 = _zz_13139[31 : 0];
  assign _zz_1004 = 1'b1;
  assign _zz_3443 = _zz_13140;
  assign _zz_3444 = _zz_13148;
  assign _zz_1005 = 1'b1;
  assign _zz_3445 = _zz_13156;
  assign _zz_3446 = _zz_13164;
  assign _zz_1008 = ($signed(_zz_13172) * $signed(data_mid_25_real));
  assign _zz_3447 = _zz_13173;
  assign _zz_1006 = _zz_13176[31 : 0];
  assign _zz_3448 = _zz_13177;
  assign _zz_1007 = _zz_13180[31 : 0];
  assign _zz_1009 = 1'b1;
  assign _zz_3449 = _zz_13181;
  assign _zz_3450 = _zz_13189;
  assign _zz_1010 = 1'b1;
  assign _zz_3451 = _zz_13197;
  assign _zz_3452 = _zz_13205;
  assign _zz_1013 = ($signed(_zz_13213) * $signed(data_mid_26_real));
  assign _zz_3453 = _zz_13214;
  assign _zz_1011 = _zz_13217[31 : 0];
  assign _zz_3454 = _zz_13218;
  assign _zz_1012 = _zz_13221[31 : 0];
  assign _zz_1014 = 1'b1;
  assign _zz_3455 = _zz_13222;
  assign _zz_3456 = _zz_13230;
  assign _zz_1015 = 1'b1;
  assign _zz_3457 = _zz_13238;
  assign _zz_3458 = _zz_13246;
  assign _zz_1018 = ($signed(_zz_13254) * $signed(data_mid_27_real));
  assign _zz_3459 = _zz_13255;
  assign _zz_1016 = _zz_13258[31 : 0];
  assign _zz_3460 = _zz_13259;
  assign _zz_1017 = _zz_13262[31 : 0];
  assign _zz_1019 = 1'b1;
  assign _zz_3461 = _zz_13263;
  assign _zz_3462 = _zz_13271;
  assign _zz_1020 = 1'b1;
  assign _zz_3463 = _zz_13279;
  assign _zz_3464 = _zz_13287;
  assign _zz_1023 = ($signed(_zz_13295) * $signed(data_mid_28_real));
  assign _zz_3465 = _zz_13296;
  assign _zz_1021 = _zz_13299[31 : 0];
  assign _zz_3466 = _zz_13300;
  assign _zz_1022 = _zz_13303[31 : 0];
  assign _zz_1024 = 1'b1;
  assign _zz_3467 = _zz_13304;
  assign _zz_3468 = _zz_13312;
  assign _zz_1025 = 1'b1;
  assign _zz_3469 = _zz_13320;
  assign _zz_3470 = _zz_13328;
  assign _zz_1028 = ($signed(_zz_13336) * $signed(data_mid_29_real));
  assign _zz_3471 = _zz_13337;
  assign _zz_1026 = _zz_13340[31 : 0];
  assign _zz_3472 = _zz_13341;
  assign _zz_1027 = _zz_13344[31 : 0];
  assign _zz_1029 = 1'b1;
  assign _zz_3473 = _zz_13345;
  assign _zz_3474 = _zz_13353;
  assign _zz_1030 = 1'b1;
  assign _zz_3475 = _zz_13361;
  assign _zz_3476 = _zz_13369;
  assign _zz_1033 = ($signed(_zz_13377) * $signed(data_mid_30_real));
  assign _zz_3477 = _zz_13378;
  assign _zz_1031 = _zz_13381[31 : 0];
  assign _zz_3478 = _zz_13382;
  assign _zz_1032 = _zz_13385[31 : 0];
  assign _zz_1034 = 1'b1;
  assign _zz_3479 = _zz_13386;
  assign _zz_3480 = _zz_13394;
  assign _zz_1035 = 1'b1;
  assign _zz_3481 = _zz_13402;
  assign _zz_3482 = _zz_13410;
  assign _zz_1038 = ($signed(_zz_13418) * $signed(data_mid_31_real));
  assign _zz_3483 = _zz_13419;
  assign _zz_1036 = _zz_13422[31 : 0];
  assign _zz_3484 = _zz_13423;
  assign _zz_1037 = _zz_13426[31 : 0];
  assign _zz_1039 = 1'b1;
  assign _zz_3485 = _zz_13427;
  assign _zz_3486 = _zz_13435;
  assign _zz_1040 = 1'b1;
  assign _zz_3487 = _zz_13443;
  assign _zz_3488 = _zz_13451;
  assign _zz_1043 = ($signed(_zz_13459) * $signed(data_mid_40_real));
  assign _zz_3489 = _zz_13460;
  assign _zz_1041 = _zz_13463[31 : 0];
  assign _zz_3490 = _zz_13464;
  assign _zz_1042 = _zz_13467[31 : 0];
  assign _zz_1044 = 1'b1;
  assign _zz_3491 = _zz_13468;
  assign _zz_3492 = _zz_13476;
  assign _zz_1045 = 1'b1;
  assign _zz_3493 = _zz_13484;
  assign _zz_3494 = _zz_13492;
  assign _zz_1048 = ($signed(_zz_13500) * $signed(data_mid_41_real));
  assign _zz_3495 = _zz_13501;
  assign _zz_1046 = _zz_13504[31 : 0];
  assign _zz_3496 = _zz_13505;
  assign _zz_1047 = _zz_13508[31 : 0];
  assign _zz_1049 = 1'b1;
  assign _zz_3497 = _zz_13509;
  assign _zz_3498 = _zz_13517;
  assign _zz_1050 = 1'b1;
  assign _zz_3499 = _zz_13525;
  assign _zz_3500 = _zz_13533;
  assign _zz_1053 = ($signed(_zz_13541) * $signed(data_mid_42_real));
  assign _zz_3501 = _zz_13542;
  assign _zz_1051 = _zz_13545[31 : 0];
  assign _zz_3502 = _zz_13546;
  assign _zz_1052 = _zz_13549[31 : 0];
  assign _zz_1054 = 1'b1;
  assign _zz_3503 = _zz_13550;
  assign _zz_3504 = _zz_13558;
  assign _zz_1055 = 1'b1;
  assign _zz_3505 = _zz_13566;
  assign _zz_3506 = _zz_13574;
  assign _zz_1058 = ($signed(_zz_13582) * $signed(data_mid_43_real));
  assign _zz_3507 = _zz_13583;
  assign _zz_1056 = _zz_13586[31 : 0];
  assign _zz_3508 = _zz_13587;
  assign _zz_1057 = _zz_13590[31 : 0];
  assign _zz_1059 = 1'b1;
  assign _zz_3509 = _zz_13591;
  assign _zz_3510 = _zz_13599;
  assign _zz_1060 = 1'b1;
  assign _zz_3511 = _zz_13607;
  assign _zz_3512 = _zz_13615;
  assign _zz_1063 = ($signed(_zz_13623) * $signed(data_mid_44_real));
  assign _zz_3513 = _zz_13624;
  assign _zz_1061 = _zz_13627[31 : 0];
  assign _zz_3514 = _zz_13628;
  assign _zz_1062 = _zz_13631[31 : 0];
  assign _zz_1064 = 1'b1;
  assign _zz_3515 = _zz_13632;
  assign _zz_3516 = _zz_13640;
  assign _zz_1065 = 1'b1;
  assign _zz_3517 = _zz_13648;
  assign _zz_3518 = _zz_13656;
  assign _zz_1068 = ($signed(_zz_13664) * $signed(data_mid_45_real));
  assign _zz_3519 = _zz_13665;
  assign _zz_1066 = _zz_13668[31 : 0];
  assign _zz_3520 = _zz_13669;
  assign _zz_1067 = _zz_13672[31 : 0];
  assign _zz_1069 = 1'b1;
  assign _zz_3521 = _zz_13673;
  assign _zz_3522 = _zz_13681;
  assign _zz_1070 = 1'b1;
  assign _zz_3523 = _zz_13689;
  assign _zz_3524 = _zz_13697;
  assign _zz_1073 = ($signed(_zz_13705) * $signed(data_mid_46_real));
  assign _zz_3525 = _zz_13706;
  assign _zz_1071 = _zz_13709[31 : 0];
  assign _zz_3526 = _zz_13710;
  assign _zz_1072 = _zz_13713[31 : 0];
  assign _zz_1074 = 1'b1;
  assign _zz_3527 = _zz_13714;
  assign _zz_3528 = _zz_13722;
  assign _zz_1075 = 1'b1;
  assign _zz_3529 = _zz_13730;
  assign _zz_3530 = _zz_13738;
  assign _zz_1078 = ($signed(_zz_13746) * $signed(data_mid_47_real));
  assign _zz_3531 = _zz_13747;
  assign _zz_1076 = _zz_13750[31 : 0];
  assign _zz_3532 = _zz_13751;
  assign _zz_1077 = _zz_13754[31 : 0];
  assign _zz_1079 = 1'b1;
  assign _zz_3533 = _zz_13755;
  assign _zz_3534 = _zz_13763;
  assign _zz_1080 = 1'b1;
  assign _zz_3535 = _zz_13771;
  assign _zz_3536 = _zz_13779;
  assign _zz_1083 = ($signed(_zz_13787) * $signed(data_mid_56_real));
  assign _zz_3537 = _zz_13788;
  assign _zz_1081 = _zz_13791[31 : 0];
  assign _zz_3538 = _zz_13792;
  assign _zz_1082 = _zz_13795[31 : 0];
  assign _zz_1084 = 1'b1;
  assign _zz_3539 = _zz_13796;
  assign _zz_3540 = _zz_13804;
  assign _zz_1085 = 1'b1;
  assign _zz_3541 = _zz_13812;
  assign _zz_3542 = _zz_13820;
  assign _zz_1088 = ($signed(_zz_13828) * $signed(data_mid_57_real));
  assign _zz_3543 = _zz_13829;
  assign _zz_1086 = _zz_13832[31 : 0];
  assign _zz_3544 = _zz_13833;
  assign _zz_1087 = _zz_13836[31 : 0];
  assign _zz_1089 = 1'b1;
  assign _zz_3545 = _zz_13837;
  assign _zz_3546 = _zz_13845;
  assign _zz_1090 = 1'b1;
  assign _zz_3547 = _zz_13853;
  assign _zz_3548 = _zz_13861;
  assign _zz_1093 = ($signed(_zz_13869) * $signed(data_mid_58_real));
  assign _zz_3549 = _zz_13870;
  assign _zz_1091 = _zz_13873[31 : 0];
  assign _zz_3550 = _zz_13874;
  assign _zz_1092 = _zz_13877[31 : 0];
  assign _zz_1094 = 1'b1;
  assign _zz_3551 = _zz_13878;
  assign _zz_3552 = _zz_13886;
  assign _zz_1095 = 1'b1;
  assign _zz_3553 = _zz_13894;
  assign _zz_3554 = _zz_13902;
  assign _zz_1098 = ($signed(_zz_13910) * $signed(data_mid_59_real));
  assign _zz_3555 = _zz_13911;
  assign _zz_1096 = _zz_13914[31 : 0];
  assign _zz_3556 = _zz_13915;
  assign _zz_1097 = _zz_13918[31 : 0];
  assign _zz_1099 = 1'b1;
  assign _zz_3557 = _zz_13919;
  assign _zz_3558 = _zz_13927;
  assign _zz_1100 = 1'b1;
  assign _zz_3559 = _zz_13935;
  assign _zz_3560 = _zz_13943;
  assign _zz_1103 = ($signed(_zz_13951) * $signed(data_mid_60_real));
  assign _zz_3561 = _zz_13952;
  assign _zz_1101 = _zz_13955[31 : 0];
  assign _zz_3562 = _zz_13956;
  assign _zz_1102 = _zz_13959[31 : 0];
  assign _zz_1104 = 1'b1;
  assign _zz_3563 = _zz_13960;
  assign _zz_3564 = _zz_13968;
  assign _zz_1105 = 1'b1;
  assign _zz_3565 = _zz_13976;
  assign _zz_3566 = _zz_13984;
  assign _zz_1108 = ($signed(_zz_13992) * $signed(data_mid_61_real));
  assign _zz_3567 = _zz_13993;
  assign _zz_1106 = _zz_13996[31 : 0];
  assign _zz_3568 = _zz_13997;
  assign _zz_1107 = _zz_14000[31 : 0];
  assign _zz_1109 = 1'b1;
  assign _zz_3569 = _zz_14001;
  assign _zz_3570 = _zz_14009;
  assign _zz_1110 = 1'b1;
  assign _zz_3571 = _zz_14017;
  assign _zz_3572 = _zz_14025;
  assign _zz_1113 = ($signed(_zz_14033) * $signed(data_mid_62_real));
  assign _zz_3573 = _zz_14034;
  assign _zz_1111 = _zz_14037[31 : 0];
  assign _zz_3574 = _zz_14038;
  assign _zz_1112 = _zz_14041[31 : 0];
  assign _zz_1114 = 1'b1;
  assign _zz_3575 = _zz_14042;
  assign _zz_3576 = _zz_14050;
  assign _zz_1115 = 1'b1;
  assign _zz_3577 = _zz_14058;
  assign _zz_3578 = _zz_14066;
  assign _zz_1118 = ($signed(_zz_14074) * $signed(data_mid_63_real));
  assign _zz_3579 = _zz_14075;
  assign _zz_1116 = _zz_14078[31 : 0];
  assign _zz_3580 = _zz_14079;
  assign _zz_1117 = _zz_14082[31 : 0];
  assign _zz_1119 = 1'b1;
  assign _zz_3581 = _zz_14083;
  assign _zz_3582 = _zz_14091;
  assign _zz_1120 = 1'b1;
  assign _zz_3583 = _zz_14099;
  assign _zz_3584 = _zz_14107;
  assign _zz_1123 = ($signed(_zz_14115) * $signed(data_mid_72_real));
  assign _zz_3585 = _zz_14116;
  assign _zz_1121 = _zz_14119[31 : 0];
  assign _zz_3586 = _zz_14120;
  assign _zz_1122 = _zz_14123[31 : 0];
  assign _zz_1124 = 1'b1;
  assign _zz_3587 = _zz_14124;
  assign _zz_3588 = _zz_14132;
  assign _zz_1125 = 1'b1;
  assign _zz_3589 = _zz_14140;
  assign _zz_3590 = _zz_14148;
  assign _zz_1128 = ($signed(_zz_14156) * $signed(data_mid_73_real));
  assign _zz_3591 = _zz_14157;
  assign _zz_1126 = _zz_14160[31 : 0];
  assign _zz_3592 = _zz_14161;
  assign _zz_1127 = _zz_14164[31 : 0];
  assign _zz_1129 = 1'b1;
  assign _zz_3593 = _zz_14165;
  assign _zz_3594 = _zz_14173;
  assign _zz_1130 = 1'b1;
  assign _zz_3595 = _zz_14181;
  assign _zz_3596 = _zz_14189;
  assign _zz_1133 = ($signed(_zz_14197) * $signed(data_mid_74_real));
  assign _zz_3597 = _zz_14198;
  assign _zz_1131 = _zz_14201[31 : 0];
  assign _zz_3598 = _zz_14202;
  assign _zz_1132 = _zz_14205[31 : 0];
  assign _zz_1134 = 1'b1;
  assign _zz_3599 = _zz_14206;
  assign _zz_3600 = _zz_14214;
  assign _zz_1135 = 1'b1;
  assign _zz_3601 = _zz_14222;
  assign _zz_3602 = _zz_14230;
  assign _zz_1138 = ($signed(_zz_14238) * $signed(data_mid_75_real));
  assign _zz_3603 = _zz_14239;
  assign _zz_1136 = _zz_14242[31 : 0];
  assign _zz_3604 = _zz_14243;
  assign _zz_1137 = _zz_14246[31 : 0];
  assign _zz_1139 = 1'b1;
  assign _zz_3605 = _zz_14247;
  assign _zz_3606 = _zz_14255;
  assign _zz_1140 = 1'b1;
  assign _zz_3607 = _zz_14263;
  assign _zz_3608 = _zz_14271;
  assign _zz_1143 = ($signed(_zz_14279) * $signed(data_mid_76_real));
  assign _zz_3609 = _zz_14280;
  assign _zz_1141 = _zz_14283[31 : 0];
  assign _zz_3610 = _zz_14284;
  assign _zz_1142 = _zz_14287[31 : 0];
  assign _zz_1144 = 1'b1;
  assign _zz_3611 = _zz_14288;
  assign _zz_3612 = _zz_14296;
  assign _zz_1145 = 1'b1;
  assign _zz_3613 = _zz_14304;
  assign _zz_3614 = _zz_14312;
  assign _zz_1148 = ($signed(_zz_14320) * $signed(data_mid_77_real));
  assign _zz_3615 = _zz_14321;
  assign _zz_1146 = _zz_14324[31 : 0];
  assign _zz_3616 = _zz_14325;
  assign _zz_1147 = _zz_14328[31 : 0];
  assign _zz_1149 = 1'b1;
  assign _zz_3617 = _zz_14329;
  assign _zz_3618 = _zz_14337;
  assign _zz_1150 = 1'b1;
  assign _zz_3619 = _zz_14345;
  assign _zz_3620 = _zz_14353;
  assign _zz_1153 = ($signed(_zz_14361) * $signed(data_mid_78_real));
  assign _zz_3621 = _zz_14362;
  assign _zz_1151 = _zz_14365[31 : 0];
  assign _zz_3622 = _zz_14366;
  assign _zz_1152 = _zz_14369[31 : 0];
  assign _zz_1154 = 1'b1;
  assign _zz_3623 = _zz_14370;
  assign _zz_3624 = _zz_14378;
  assign _zz_1155 = 1'b1;
  assign _zz_3625 = _zz_14386;
  assign _zz_3626 = _zz_14394;
  assign _zz_1158 = ($signed(_zz_14402) * $signed(data_mid_79_real));
  assign _zz_3627 = _zz_14403;
  assign _zz_1156 = _zz_14406[31 : 0];
  assign _zz_3628 = _zz_14407;
  assign _zz_1157 = _zz_14410[31 : 0];
  assign _zz_1159 = 1'b1;
  assign _zz_3629 = _zz_14411;
  assign _zz_3630 = _zz_14419;
  assign _zz_1160 = 1'b1;
  assign _zz_3631 = _zz_14427;
  assign _zz_3632 = _zz_14435;
  assign _zz_1163 = ($signed(_zz_14443) * $signed(data_mid_88_real));
  assign _zz_3633 = _zz_14444;
  assign _zz_1161 = _zz_14447[31 : 0];
  assign _zz_3634 = _zz_14448;
  assign _zz_1162 = _zz_14451[31 : 0];
  assign _zz_1164 = 1'b1;
  assign _zz_3635 = _zz_14452;
  assign _zz_3636 = _zz_14460;
  assign _zz_1165 = 1'b1;
  assign _zz_3637 = _zz_14468;
  assign _zz_3638 = _zz_14476;
  assign _zz_1168 = ($signed(_zz_14484) * $signed(data_mid_89_real));
  assign _zz_3639 = _zz_14485;
  assign _zz_1166 = _zz_14488[31 : 0];
  assign _zz_3640 = _zz_14489;
  assign _zz_1167 = _zz_14492[31 : 0];
  assign _zz_1169 = 1'b1;
  assign _zz_3641 = _zz_14493;
  assign _zz_3642 = _zz_14501;
  assign _zz_1170 = 1'b1;
  assign _zz_3643 = _zz_14509;
  assign _zz_3644 = _zz_14517;
  assign _zz_1173 = ($signed(_zz_14525) * $signed(data_mid_90_real));
  assign _zz_3645 = _zz_14526;
  assign _zz_1171 = _zz_14529[31 : 0];
  assign _zz_3646 = _zz_14530;
  assign _zz_1172 = _zz_14533[31 : 0];
  assign _zz_1174 = 1'b1;
  assign _zz_3647 = _zz_14534;
  assign _zz_3648 = _zz_14542;
  assign _zz_1175 = 1'b1;
  assign _zz_3649 = _zz_14550;
  assign _zz_3650 = _zz_14558;
  assign _zz_1178 = ($signed(_zz_14566) * $signed(data_mid_91_real));
  assign _zz_3651 = _zz_14567;
  assign _zz_1176 = _zz_14570[31 : 0];
  assign _zz_3652 = _zz_14571;
  assign _zz_1177 = _zz_14574[31 : 0];
  assign _zz_1179 = 1'b1;
  assign _zz_3653 = _zz_14575;
  assign _zz_3654 = _zz_14583;
  assign _zz_1180 = 1'b1;
  assign _zz_3655 = _zz_14591;
  assign _zz_3656 = _zz_14599;
  assign _zz_1183 = ($signed(_zz_14607) * $signed(data_mid_92_real));
  assign _zz_3657 = _zz_14608;
  assign _zz_1181 = _zz_14611[31 : 0];
  assign _zz_3658 = _zz_14612;
  assign _zz_1182 = _zz_14615[31 : 0];
  assign _zz_1184 = 1'b1;
  assign _zz_3659 = _zz_14616;
  assign _zz_3660 = _zz_14624;
  assign _zz_1185 = 1'b1;
  assign _zz_3661 = _zz_14632;
  assign _zz_3662 = _zz_14640;
  assign _zz_1188 = ($signed(_zz_14648) * $signed(data_mid_93_real));
  assign _zz_3663 = _zz_14649;
  assign _zz_1186 = _zz_14652[31 : 0];
  assign _zz_3664 = _zz_14653;
  assign _zz_1187 = _zz_14656[31 : 0];
  assign _zz_1189 = 1'b1;
  assign _zz_3665 = _zz_14657;
  assign _zz_3666 = _zz_14665;
  assign _zz_1190 = 1'b1;
  assign _zz_3667 = _zz_14673;
  assign _zz_3668 = _zz_14681;
  assign _zz_1193 = ($signed(_zz_14689) * $signed(data_mid_94_real));
  assign _zz_3669 = _zz_14690;
  assign _zz_1191 = _zz_14693[31 : 0];
  assign _zz_3670 = _zz_14694;
  assign _zz_1192 = _zz_14697[31 : 0];
  assign _zz_1194 = 1'b1;
  assign _zz_3671 = _zz_14698;
  assign _zz_3672 = _zz_14706;
  assign _zz_1195 = 1'b1;
  assign _zz_3673 = _zz_14714;
  assign _zz_3674 = _zz_14722;
  assign _zz_1198 = ($signed(_zz_14730) * $signed(data_mid_95_real));
  assign _zz_3675 = _zz_14731;
  assign _zz_1196 = _zz_14734[31 : 0];
  assign _zz_3676 = _zz_14735;
  assign _zz_1197 = _zz_14738[31 : 0];
  assign _zz_1199 = 1'b1;
  assign _zz_3677 = _zz_14739;
  assign _zz_3678 = _zz_14747;
  assign _zz_1200 = 1'b1;
  assign _zz_3679 = _zz_14755;
  assign _zz_3680 = _zz_14763;
  assign _zz_1203 = ($signed(_zz_14771) * $signed(data_mid_104_real));
  assign _zz_3681 = _zz_14772;
  assign _zz_1201 = _zz_14775[31 : 0];
  assign _zz_3682 = _zz_14776;
  assign _zz_1202 = _zz_14779[31 : 0];
  assign _zz_1204 = 1'b1;
  assign _zz_3683 = _zz_14780;
  assign _zz_3684 = _zz_14788;
  assign _zz_1205 = 1'b1;
  assign _zz_3685 = _zz_14796;
  assign _zz_3686 = _zz_14804;
  assign _zz_1208 = ($signed(_zz_14812) * $signed(data_mid_105_real));
  assign _zz_3687 = _zz_14813;
  assign _zz_1206 = _zz_14816[31 : 0];
  assign _zz_3688 = _zz_14817;
  assign _zz_1207 = _zz_14820[31 : 0];
  assign _zz_1209 = 1'b1;
  assign _zz_3689 = _zz_14821;
  assign _zz_3690 = _zz_14829;
  assign _zz_1210 = 1'b1;
  assign _zz_3691 = _zz_14837;
  assign _zz_3692 = _zz_14845;
  assign _zz_1213 = ($signed(_zz_14853) * $signed(data_mid_106_real));
  assign _zz_3693 = _zz_14854;
  assign _zz_1211 = _zz_14857[31 : 0];
  assign _zz_3694 = _zz_14858;
  assign _zz_1212 = _zz_14861[31 : 0];
  assign _zz_1214 = 1'b1;
  assign _zz_3695 = _zz_14862;
  assign _zz_3696 = _zz_14870;
  assign _zz_1215 = 1'b1;
  assign _zz_3697 = _zz_14878;
  assign _zz_3698 = _zz_14886;
  assign _zz_1218 = ($signed(_zz_14894) * $signed(data_mid_107_real));
  assign _zz_3699 = _zz_14895;
  assign _zz_1216 = _zz_14898[31 : 0];
  assign _zz_3700 = _zz_14899;
  assign _zz_1217 = _zz_14902[31 : 0];
  assign _zz_1219 = 1'b1;
  assign _zz_3701 = _zz_14903;
  assign _zz_3702 = _zz_14911;
  assign _zz_1220 = 1'b1;
  assign _zz_3703 = _zz_14919;
  assign _zz_3704 = _zz_14927;
  assign _zz_1223 = ($signed(_zz_14935) * $signed(data_mid_108_real));
  assign _zz_3705 = _zz_14936;
  assign _zz_1221 = _zz_14939[31 : 0];
  assign _zz_3706 = _zz_14940;
  assign _zz_1222 = _zz_14943[31 : 0];
  assign _zz_1224 = 1'b1;
  assign _zz_3707 = _zz_14944;
  assign _zz_3708 = _zz_14952;
  assign _zz_1225 = 1'b1;
  assign _zz_3709 = _zz_14960;
  assign _zz_3710 = _zz_14968;
  assign _zz_1228 = ($signed(_zz_14976) * $signed(data_mid_109_real));
  assign _zz_3711 = _zz_14977;
  assign _zz_1226 = _zz_14980[31 : 0];
  assign _zz_3712 = _zz_14981;
  assign _zz_1227 = _zz_14984[31 : 0];
  assign _zz_1229 = 1'b1;
  assign _zz_3713 = _zz_14985;
  assign _zz_3714 = _zz_14993;
  assign _zz_1230 = 1'b1;
  assign _zz_3715 = _zz_15001;
  assign _zz_3716 = _zz_15009;
  assign _zz_1233 = ($signed(_zz_15017) * $signed(data_mid_110_real));
  assign _zz_3717 = _zz_15018;
  assign _zz_1231 = _zz_15021[31 : 0];
  assign _zz_3718 = _zz_15022;
  assign _zz_1232 = _zz_15025[31 : 0];
  assign _zz_1234 = 1'b1;
  assign _zz_3719 = _zz_15026;
  assign _zz_3720 = _zz_15034;
  assign _zz_1235 = 1'b1;
  assign _zz_3721 = _zz_15042;
  assign _zz_3722 = _zz_15050;
  assign _zz_1238 = ($signed(_zz_15058) * $signed(data_mid_111_real));
  assign _zz_3723 = _zz_15059;
  assign _zz_1236 = _zz_15062[31 : 0];
  assign _zz_3724 = _zz_15063;
  assign _zz_1237 = _zz_15066[31 : 0];
  assign _zz_1239 = 1'b1;
  assign _zz_3725 = _zz_15067;
  assign _zz_3726 = _zz_15075;
  assign _zz_1240 = 1'b1;
  assign _zz_3727 = _zz_15083;
  assign _zz_3728 = _zz_15091;
  assign _zz_1243 = ($signed(_zz_15099) * $signed(data_mid_120_real));
  assign _zz_3729 = _zz_15100;
  assign _zz_1241 = _zz_15103[31 : 0];
  assign _zz_3730 = _zz_15104;
  assign _zz_1242 = _zz_15107[31 : 0];
  assign _zz_1244 = 1'b1;
  assign _zz_3731 = _zz_15108;
  assign _zz_3732 = _zz_15116;
  assign _zz_1245 = 1'b1;
  assign _zz_3733 = _zz_15124;
  assign _zz_3734 = _zz_15132;
  assign _zz_1248 = ($signed(_zz_15140) * $signed(data_mid_121_real));
  assign _zz_3735 = _zz_15141;
  assign _zz_1246 = _zz_15144[31 : 0];
  assign _zz_3736 = _zz_15145;
  assign _zz_1247 = _zz_15148[31 : 0];
  assign _zz_1249 = 1'b1;
  assign _zz_3737 = _zz_15149;
  assign _zz_3738 = _zz_15157;
  assign _zz_1250 = 1'b1;
  assign _zz_3739 = _zz_15165;
  assign _zz_3740 = _zz_15173;
  assign _zz_1253 = ($signed(_zz_15181) * $signed(data_mid_122_real));
  assign _zz_3741 = _zz_15182;
  assign _zz_1251 = _zz_15185[31 : 0];
  assign _zz_3742 = _zz_15186;
  assign _zz_1252 = _zz_15189[31 : 0];
  assign _zz_1254 = 1'b1;
  assign _zz_3743 = _zz_15190;
  assign _zz_3744 = _zz_15198;
  assign _zz_1255 = 1'b1;
  assign _zz_3745 = _zz_15206;
  assign _zz_3746 = _zz_15214;
  assign _zz_1258 = ($signed(_zz_15222) * $signed(data_mid_123_real));
  assign _zz_3747 = _zz_15223;
  assign _zz_1256 = _zz_15226[31 : 0];
  assign _zz_3748 = _zz_15227;
  assign _zz_1257 = _zz_15230[31 : 0];
  assign _zz_1259 = 1'b1;
  assign _zz_3749 = _zz_15231;
  assign _zz_3750 = _zz_15239;
  assign _zz_1260 = 1'b1;
  assign _zz_3751 = _zz_15247;
  assign _zz_3752 = _zz_15255;
  assign _zz_1263 = ($signed(_zz_15263) * $signed(data_mid_124_real));
  assign _zz_3753 = _zz_15264;
  assign _zz_1261 = _zz_15267[31 : 0];
  assign _zz_3754 = _zz_15268;
  assign _zz_1262 = _zz_15271[31 : 0];
  assign _zz_1264 = 1'b1;
  assign _zz_3755 = _zz_15272;
  assign _zz_3756 = _zz_15280;
  assign _zz_1265 = 1'b1;
  assign _zz_3757 = _zz_15288;
  assign _zz_3758 = _zz_15296;
  assign _zz_1268 = ($signed(_zz_15304) * $signed(data_mid_125_real));
  assign _zz_3759 = _zz_15305;
  assign _zz_1266 = _zz_15308[31 : 0];
  assign _zz_3760 = _zz_15309;
  assign _zz_1267 = _zz_15312[31 : 0];
  assign _zz_1269 = 1'b1;
  assign _zz_3761 = _zz_15313;
  assign _zz_3762 = _zz_15321;
  assign _zz_1270 = 1'b1;
  assign _zz_3763 = _zz_15329;
  assign _zz_3764 = _zz_15337;
  assign _zz_1273 = ($signed(_zz_15345) * $signed(data_mid_126_real));
  assign _zz_3765 = _zz_15346;
  assign _zz_1271 = _zz_15349[31 : 0];
  assign _zz_3766 = _zz_15350;
  assign _zz_1272 = _zz_15353[31 : 0];
  assign _zz_1274 = 1'b1;
  assign _zz_3767 = _zz_15354;
  assign _zz_3768 = _zz_15362;
  assign _zz_1275 = 1'b1;
  assign _zz_3769 = _zz_15370;
  assign _zz_3770 = _zz_15378;
  assign _zz_1278 = ($signed(_zz_15386) * $signed(data_mid_127_real));
  assign _zz_3771 = _zz_15387;
  assign _zz_1276 = _zz_15390[31 : 0];
  assign _zz_3772 = _zz_15391;
  assign _zz_1277 = _zz_15394[31 : 0];
  assign _zz_1279 = 1'b1;
  assign _zz_3773 = _zz_15395;
  assign _zz_3774 = _zz_15403;
  assign _zz_1280 = 1'b1;
  assign _zz_3775 = _zz_15411;
  assign _zz_3776 = _zz_15419;
  assign _zz_1283 = ($signed(_zz_15427) * $signed(data_mid_16_real));
  assign _zz_3777 = _zz_15428;
  assign _zz_1281 = _zz_15431[31 : 0];
  assign _zz_3778 = _zz_15432;
  assign _zz_1282 = _zz_15435[31 : 0];
  assign _zz_1284 = 1'b1;
  assign _zz_3779 = _zz_15436;
  assign _zz_3780 = _zz_15444;
  assign _zz_1285 = 1'b1;
  assign _zz_3781 = _zz_15452;
  assign _zz_3782 = _zz_15460;
  assign _zz_1288 = ($signed(_zz_15468) * $signed(data_mid_17_real));
  assign _zz_3783 = _zz_15469;
  assign _zz_1286 = _zz_15472[31 : 0];
  assign _zz_3784 = _zz_15473;
  assign _zz_1287 = _zz_15476[31 : 0];
  assign _zz_1289 = 1'b1;
  assign _zz_3785 = _zz_15477;
  assign _zz_3786 = _zz_15485;
  assign _zz_1290 = 1'b1;
  assign _zz_3787 = _zz_15493;
  assign _zz_3788 = _zz_15501;
  assign _zz_1293 = ($signed(_zz_15509) * $signed(data_mid_18_real));
  assign _zz_3789 = _zz_15510;
  assign _zz_1291 = _zz_15513[31 : 0];
  assign _zz_3790 = _zz_15514;
  assign _zz_1292 = _zz_15517[31 : 0];
  assign _zz_1294 = 1'b1;
  assign _zz_3791 = _zz_15518;
  assign _zz_3792 = _zz_15526;
  assign _zz_1295 = 1'b1;
  assign _zz_3793 = _zz_15534;
  assign _zz_3794 = _zz_15542;
  assign _zz_1298 = ($signed(_zz_15550) * $signed(data_mid_19_real));
  assign _zz_3795 = _zz_15551;
  assign _zz_1296 = _zz_15554[31 : 0];
  assign _zz_3796 = _zz_15555;
  assign _zz_1297 = _zz_15558[31 : 0];
  assign _zz_1299 = 1'b1;
  assign _zz_3797 = _zz_15559;
  assign _zz_3798 = _zz_15567;
  assign _zz_1300 = 1'b1;
  assign _zz_3799 = _zz_15575;
  assign _zz_3800 = _zz_15583;
  assign _zz_1303 = ($signed(_zz_15591) * $signed(data_mid_20_real));
  assign _zz_3801 = _zz_15592;
  assign _zz_1301 = _zz_15595[31 : 0];
  assign _zz_3802 = _zz_15596;
  assign _zz_1302 = _zz_15599[31 : 0];
  assign _zz_1304 = 1'b1;
  assign _zz_3803 = _zz_15600;
  assign _zz_3804 = _zz_15608;
  assign _zz_1305 = 1'b1;
  assign _zz_3805 = _zz_15616;
  assign _zz_3806 = _zz_15624;
  assign _zz_1308 = ($signed(_zz_15632) * $signed(data_mid_21_real));
  assign _zz_3807 = _zz_15633;
  assign _zz_1306 = _zz_15636[31 : 0];
  assign _zz_3808 = _zz_15637;
  assign _zz_1307 = _zz_15640[31 : 0];
  assign _zz_1309 = 1'b1;
  assign _zz_3809 = _zz_15641;
  assign _zz_3810 = _zz_15649;
  assign _zz_1310 = 1'b1;
  assign _zz_3811 = _zz_15657;
  assign _zz_3812 = _zz_15665;
  assign _zz_1313 = ($signed(_zz_15673) * $signed(data_mid_22_real));
  assign _zz_3813 = _zz_15674;
  assign _zz_1311 = _zz_15677[31 : 0];
  assign _zz_3814 = _zz_15678;
  assign _zz_1312 = _zz_15681[31 : 0];
  assign _zz_1314 = 1'b1;
  assign _zz_3815 = _zz_15682;
  assign _zz_3816 = _zz_15690;
  assign _zz_1315 = 1'b1;
  assign _zz_3817 = _zz_15698;
  assign _zz_3818 = _zz_15706;
  assign _zz_1318 = ($signed(_zz_15714) * $signed(data_mid_23_real));
  assign _zz_3819 = _zz_15715;
  assign _zz_1316 = _zz_15718[31 : 0];
  assign _zz_3820 = _zz_15719;
  assign _zz_1317 = _zz_15722[31 : 0];
  assign _zz_1319 = 1'b1;
  assign _zz_3821 = _zz_15723;
  assign _zz_3822 = _zz_15731;
  assign _zz_1320 = 1'b1;
  assign _zz_3823 = _zz_15739;
  assign _zz_3824 = _zz_15747;
  assign _zz_1323 = ($signed(_zz_15755) * $signed(data_mid_24_real));
  assign _zz_3825 = _zz_15756;
  assign _zz_1321 = _zz_15759[31 : 0];
  assign _zz_3826 = _zz_15760;
  assign _zz_1322 = _zz_15763[31 : 0];
  assign _zz_1324 = 1'b1;
  assign _zz_3827 = _zz_15764;
  assign _zz_3828 = _zz_15772;
  assign _zz_1325 = 1'b1;
  assign _zz_3829 = _zz_15780;
  assign _zz_3830 = _zz_15788;
  assign _zz_1328 = ($signed(_zz_15796) * $signed(data_mid_25_real));
  assign _zz_3831 = _zz_15797;
  assign _zz_1326 = _zz_15800[31 : 0];
  assign _zz_3832 = _zz_15801;
  assign _zz_1327 = _zz_15804[31 : 0];
  assign _zz_1329 = 1'b1;
  assign _zz_3833 = _zz_15805;
  assign _zz_3834 = _zz_15813;
  assign _zz_1330 = 1'b1;
  assign _zz_3835 = _zz_15821;
  assign _zz_3836 = _zz_15829;
  assign _zz_1333 = ($signed(_zz_15837) * $signed(data_mid_26_real));
  assign _zz_3837 = _zz_15838;
  assign _zz_1331 = _zz_15841[31 : 0];
  assign _zz_3838 = _zz_15842;
  assign _zz_1332 = _zz_15845[31 : 0];
  assign _zz_1334 = 1'b1;
  assign _zz_3839 = _zz_15846;
  assign _zz_3840 = _zz_15854;
  assign _zz_1335 = 1'b1;
  assign _zz_3841 = _zz_15862;
  assign _zz_3842 = _zz_15870;
  assign _zz_1338 = ($signed(_zz_15878) * $signed(data_mid_27_real));
  assign _zz_3843 = _zz_15879;
  assign _zz_1336 = _zz_15882[31 : 0];
  assign _zz_3844 = _zz_15883;
  assign _zz_1337 = _zz_15886[31 : 0];
  assign _zz_1339 = 1'b1;
  assign _zz_3845 = _zz_15887;
  assign _zz_3846 = _zz_15895;
  assign _zz_1340 = 1'b1;
  assign _zz_3847 = _zz_15903;
  assign _zz_3848 = _zz_15911;
  assign _zz_1343 = ($signed(_zz_15919) * $signed(data_mid_28_real));
  assign _zz_3849 = _zz_15920;
  assign _zz_1341 = _zz_15923[31 : 0];
  assign _zz_3850 = _zz_15924;
  assign _zz_1342 = _zz_15927[31 : 0];
  assign _zz_1344 = 1'b1;
  assign _zz_3851 = _zz_15928;
  assign _zz_3852 = _zz_15936;
  assign _zz_1345 = 1'b1;
  assign _zz_3853 = _zz_15944;
  assign _zz_3854 = _zz_15952;
  assign _zz_1348 = ($signed(_zz_15960) * $signed(data_mid_29_real));
  assign _zz_3855 = _zz_15961;
  assign _zz_1346 = _zz_15964[31 : 0];
  assign _zz_3856 = _zz_15965;
  assign _zz_1347 = _zz_15968[31 : 0];
  assign _zz_1349 = 1'b1;
  assign _zz_3857 = _zz_15969;
  assign _zz_3858 = _zz_15977;
  assign _zz_1350 = 1'b1;
  assign _zz_3859 = _zz_15985;
  assign _zz_3860 = _zz_15993;
  assign _zz_1353 = ($signed(_zz_16001) * $signed(data_mid_30_real));
  assign _zz_3861 = _zz_16002;
  assign _zz_1351 = _zz_16005[31 : 0];
  assign _zz_3862 = _zz_16006;
  assign _zz_1352 = _zz_16009[31 : 0];
  assign _zz_1354 = 1'b1;
  assign _zz_3863 = _zz_16010;
  assign _zz_3864 = _zz_16018;
  assign _zz_1355 = 1'b1;
  assign _zz_3865 = _zz_16026;
  assign _zz_3866 = _zz_16034;
  assign _zz_1358 = ($signed(_zz_16042) * $signed(data_mid_31_real));
  assign _zz_3867 = _zz_16043;
  assign _zz_1356 = _zz_16046[31 : 0];
  assign _zz_3868 = _zz_16047;
  assign _zz_1357 = _zz_16050[31 : 0];
  assign _zz_1359 = 1'b1;
  assign _zz_3869 = _zz_16051;
  assign _zz_3870 = _zz_16059;
  assign _zz_1360 = 1'b1;
  assign _zz_3871 = _zz_16067;
  assign _zz_3872 = _zz_16075;
  assign _zz_1363 = ($signed(_zz_16083) * $signed(data_mid_48_real));
  assign _zz_3873 = _zz_16084;
  assign _zz_1361 = _zz_16087[31 : 0];
  assign _zz_3874 = _zz_16088;
  assign _zz_1362 = _zz_16091[31 : 0];
  assign _zz_1364 = 1'b1;
  assign _zz_3875 = _zz_16092;
  assign _zz_3876 = _zz_16100;
  assign _zz_1365 = 1'b1;
  assign _zz_3877 = _zz_16108;
  assign _zz_3878 = _zz_16116;
  assign _zz_1368 = ($signed(_zz_16124) * $signed(data_mid_49_real));
  assign _zz_3879 = _zz_16125;
  assign _zz_1366 = _zz_16128[31 : 0];
  assign _zz_3880 = _zz_16129;
  assign _zz_1367 = _zz_16132[31 : 0];
  assign _zz_1369 = 1'b1;
  assign _zz_3881 = _zz_16133;
  assign _zz_3882 = _zz_16141;
  assign _zz_1370 = 1'b1;
  assign _zz_3883 = _zz_16149;
  assign _zz_3884 = _zz_16157;
  assign _zz_1373 = ($signed(_zz_16165) * $signed(data_mid_50_real));
  assign _zz_3885 = _zz_16166;
  assign _zz_1371 = _zz_16169[31 : 0];
  assign _zz_3886 = _zz_16170;
  assign _zz_1372 = _zz_16173[31 : 0];
  assign _zz_1374 = 1'b1;
  assign _zz_3887 = _zz_16174;
  assign _zz_3888 = _zz_16182;
  assign _zz_1375 = 1'b1;
  assign _zz_3889 = _zz_16190;
  assign _zz_3890 = _zz_16198;
  assign _zz_1378 = ($signed(_zz_16206) * $signed(data_mid_51_real));
  assign _zz_3891 = _zz_16207;
  assign _zz_1376 = _zz_16210[31 : 0];
  assign _zz_3892 = _zz_16211;
  assign _zz_1377 = _zz_16214[31 : 0];
  assign _zz_1379 = 1'b1;
  assign _zz_3893 = _zz_16215;
  assign _zz_3894 = _zz_16223;
  assign _zz_1380 = 1'b1;
  assign _zz_3895 = _zz_16231;
  assign _zz_3896 = _zz_16239;
  assign _zz_1383 = ($signed(_zz_16247) * $signed(data_mid_52_real));
  assign _zz_3897 = _zz_16248;
  assign _zz_1381 = _zz_16251[31 : 0];
  assign _zz_3898 = _zz_16252;
  assign _zz_1382 = _zz_16255[31 : 0];
  assign _zz_1384 = 1'b1;
  assign _zz_3899 = _zz_16256;
  assign _zz_3900 = _zz_16264;
  assign _zz_1385 = 1'b1;
  assign _zz_3901 = _zz_16272;
  assign _zz_3902 = _zz_16280;
  assign _zz_1388 = ($signed(_zz_16288) * $signed(data_mid_53_real));
  assign _zz_3903 = _zz_16289;
  assign _zz_1386 = _zz_16292[31 : 0];
  assign _zz_3904 = _zz_16293;
  assign _zz_1387 = _zz_16296[31 : 0];
  assign _zz_1389 = 1'b1;
  assign _zz_3905 = _zz_16297;
  assign _zz_3906 = _zz_16305;
  assign _zz_1390 = 1'b1;
  assign _zz_3907 = _zz_16313;
  assign _zz_3908 = _zz_16321;
  assign _zz_1393 = ($signed(_zz_16329) * $signed(data_mid_54_real));
  assign _zz_3909 = _zz_16330;
  assign _zz_1391 = _zz_16333[31 : 0];
  assign _zz_3910 = _zz_16334;
  assign _zz_1392 = _zz_16337[31 : 0];
  assign _zz_1394 = 1'b1;
  assign _zz_3911 = _zz_16338;
  assign _zz_3912 = _zz_16346;
  assign _zz_1395 = 1'b1;
  assign _zz_3913 = _zz_16354;
  assign _zz_3914 = _zz_16362;
  assign _zz_1398 = ($signed(_zz_16370) * $signed(data_mid_55_real));
  assign _zz_3915 = _zz_16371;
  assign _zz_1396 = _zz_16374[31 : 0];
  assign _zz_3916 = _zz_16375;
  assign _zz_1397 = _zz_16378[31 : 0];
  assign _zz_1399 = 1'b1;
  assign _zz_3917 = _zz_16379;
  assign _zz_3918 = _zz_16387;
  assign _zz_1400 = 1'b1;
  assign _zz_3919 = _zz_16395;
  assign _zz_3920 = _zz_16403;
  assign _zz_1403 = ($signed(_zz_16411) * $signed(data_mid_56_real));
  assign _zz_3921 = _zz_16412;
  assign _zz_1401 = _zz_16415[31 : 0];
  assign _zz_3922 = _zz_16416;
  assign _zz_1402 = _zz_16419[31 : 0];
  assign _zz_1404 = 1'b1;
  assign _zz_3923 = _zz_16420;
  assign _zz_3924 = _zz_16428;
  assign _zz_1405 = 1'b1;
  assign _zz_3925 = _zz_16436;
  assign _zz_3926 = _zz_16444;
  assign _zz_1408 = ($signed(_zz_16452) * $signed(data_mid_57_real));
  assign _zz_3927 = _zz_16453;
  assign _zz_1406 = _zz_16456[31 : 0];
  assign _zz_3928 = _zz_16457;
  assign _zz_1407 = _zz_16460[31 : 0];
  assign _zz_1409 = 1'b1;
  assign _zz_3929 = _zz_16461;
  assign _zz_3930 = _zz_16469;
  assign _zz_1410 = 1'b1;
  assign _zz_3931 = _zz_16477;
  assign _zz_3932 = _zz_16485;
  assign _zz_1413 = ($signed(_zz_16493) * $signed(data_mid_58_real));
  assign _zz_3933 = _zz_16494;
  assign _zz_1411 = _zz_16497[31 : 0];
  assign _zz_3934 = _zz_16498;
  assign _zz_1412 = _zz_16501[31 : 0];
  assign _zz_1414 = 1'b1;
  assign _zz_3935 = _zz_16502;
  assign _zz_3936 = _zz_16510;
  assign _zz_1415 = 1'b1;
  assign _zz_3937 = _zz_16518;
  assign _zz_3938 = _zz_16526;
  assign _zz_1418 = ($signed(_zz_16534) * $signed(data_mid_59_real));
  assign _zz_3939 = _zz_16535;
  assign _zz_1416 = _zz_16538[31 : 0];
  assign _zz_3940 = _zz_16539;
  assign _zz_1417 = _zz_16542[31 : 0];
  assign _zz_1419 = 1'b1;
  assign _zz_3941 = _zz_16543;
  assign _zz_3942 = _zz_16551;
  assign _zz_1420 = 1'b1;
  assign _zz_3943 = _zz_16559;
  assign _zz_3944 = _zz_16567;
  assign _zz_1423 = ($signed(_zz_16575) * $signed(data_mid_60_real));
  assign _zz_3945 = _zz_16576;
  assign _zz_1421 = _zz_16579[31 : 0];
  assign _zz_3946 = _zz_16580;
  assign _zz_1422 = _zz_16583[31 : 0];
  assign _zz_1424 = 1'b1;
  assign _zz_3947 = _zz_16584;
  assign _zz_3948 = _zz_16592;
  assign _zz_1425 = 1'b1;
  assign _zz_3949 = _zz_16600;
  assign _zz_3950 = _zz_16608;
  assign _zz_1428 = ($signed(_zz_16616) * $signed(data_mid_61_real));
  assign _zz_3951 = _zz_16617;
  assign _zz_1426 = _zz_16620[31 : 0];
  assign _zz_3952 = _zz_16621;
  assign _zz_1427 = _zz_16624[31 : 0];
  assign _zz_1429 = 1'b1;
  assign _zz_3953 = _zz_16625;
  assign _zz_3954 = _zz_16633;
  assign _zz_1430 = 1'b1;
  assign _zz_3955 = _zz_16641;
  assign _zz_3956 = _zz_16649;
  assign _zz_1433 = ($signed(_zz_16657) * $signed(data_mid_62_real));
  assign _zz_3957 = _zz_16658;
  assign _zz_1431 = _zz_16661[31 : 0];
  assign _zz_3958 = _zz_16662;
  assign _zz_1432 = _zz_16665[31 : 0];
  assign _zz_1434 = 1'b1;
  assign _zz_3959 = _zz_16666;
  assign _zz_3960 = _zz_16674;
  assign _zz_1435 = 1'b1;
  assign _zz_3961 = _zz_16682;
  assign _zz_3962 = _zz_16690;
  assign _zz_1438 = ($signed(_zz_16698) * $signed(data_mid_63_real));
  assign _zz_3963 = _zz_16699;
  assign _zz_1436 = _zz_16702[31 : 0];
  assign _zz_3964 = _zz_16703;
  assign _zz_1437 = _zz_16706[31 : 0];
  assign _zz_1439 = 1'b1;
  assign _zz_3965 = _zz_16707;
  assign _zz_3966 = _zz_16715;
  assign _zz_1440 = 1'b1;
  assign _zz_3967 = _zz_16723;
  assign _zz_3968 = _zz_16731;
  assign _zz_1443 = ($signed(_zz_16739) * $signed(data_mid_80_real));
  assign _zz_3969 = _zz_16740;
  assign _zz_1441 = _zz_16743[31 : 0];
  assign _zz_3970 = _zz_16744;
  assign _zz_1442 = _zz_16747[31 : 0];
  assign _zz_1444 = 1'b1;
  assign _zz_3971 = _zz_16748;
  assign _zz_3972 = _zz_16756;
  assign _zz_1445 = 1'b1;
  assign _zz_3973 = _zz_16764;
  assign _zz_3974 = _zz_16772;
  assign _zz_1448 = ($signed(_zz_16780) * $signed(data_mid_81_real));
  assign _zz_3975 = _zz_16781;
  assign _zz_1446 = _zz_16784[31 : 0];
  assign _zz_3976 = _zz_16785;
  assign _zz_1447 = _zz_16788[31 : 0];
  assign _zz_1449 = 1'b1;
  assign _zz_3977 = _zz_16789;
  assign _zz_3978 = _zz_16797;
  assign _zz_1450 = 1'b1;
  assign _zz_3979 = _zz_16805;
  assign _zz_3980 = _zz_16813;
  assign _zz_1453 = ($signed(_zz_16821) * $signed(data_mid_82_real));
  assign _zz_3981 = _zz_16822;
  assign _zz_1451 = _zz_16825[31 : 0];
  assign _zz_3982 = _zz_16826;
  assign _zz_1452 = _zz_16829[31 : 0];
  assign _zz_1454 = 1'b1;
  assign _zz_3983 = _zz_16830;
  assign _zz_3984 = _zz_16838;
  assign _zz_1455 = 1'b1;
  assign _zz_3985 = _zz_16846;
  assign _zz_3986 = _zz_16854;
  assign _zz_1458 = ($signed(_zz_16862) * $signed(data_mid_83_real));
  assign _zz_3987 = _zz_16863;
  assign _zz_1456 = _zz_16866[31 : 0];
  assign _zz_3988 = _zz_16867;
  assign _zz_1457 = _zz_16870[31 : 0];
  assign _zz_1459 = 1'b1;
  assign _zz_3989 = _zz_16871;
  assign _zz_3990 = _zz_16879;
  assign _zz_1460 = 1'b1;
  assign _zz_3991 = _zz_16887;
  assign _zz_3992 = _zz_16895;
  assign _zz_1463 = ($signed(_zz_16903) * $signed(data_mid_84_real));
  assign _zz_3993 = _zz_16904;
  assign _zz_1461 = _zz_16907[31 : 0];
  assign _zz_3994 = _zz_16908;
  assign _zz_1462 = _zz_16911[31 : 0];
  assign _zz_1464 = 1'b1;
  assign _zz_3995 = _zz_16912;
  assign _zz_3996 = _zz_16920;
  assign _zz_1465 = 1'b1;
  assign _zz_3997 = _zz_16928;
  assign _zz_3998 = _zz_16936;
  assign _zz_1468 = ($signed(_zz_16944) * $signed(data_mid_85_real));
  assign _zz_3999 = _zz_16945;
  assign _zz_1466 = _zz_16948[31 : 0];
  assign _zz_4000 = _zz_16949;
  assign _zz_1467 = _zz_16952[31 : 0];
  assign _zz_1469 = 1'b1;
  assign _zz_4001 = _zz_16953;
  assign _zz_4002 = _zz_16961;
  assign _zz_1470 = 1'b1;
  assign _zz_4003 = _zz_16969;
  assign _zz_4004 = _zz_16977;
  assign _zz_1473 = ($signed(_zz_16985) * $signed(data_mid_86_real));
  assign _zz_4005 = _zz_16986;
  assign _zz_1471 = _zz_16989[31 : 0];
  assign _zz_4006 = _zz_16990;
  assign _zz_1472 = _zz_16993[31 : 0];
  assign _zz_1474 = 1'b1;
  assign _zz_4007 = _zz_16994;
  assign _zz_4008 = _zz_17002;
  assign _zz_1475 = 1'b1;
  assign _zz_4009 = _zz_17010;
  assign _zz_4010 = _zz_17018;
  assign _zz_1478 = ($signed(_zz_17026) * $signed(data_mid_87_real));
  assign _zz_4011 = _zz_17027;
  assign _zz_1476 = _zz_17030[31 : 0];
  assign _zz_4012 = _zz_17031;
  assign _zz_1477 = _zz_17034[31 : 0];
  assign _zz_1479 = 1'b1;
  assign _zz_4013 = _zz_17035;
  assign _zz_4014 = _zz_17043;
  assign _zz_1480 = 1'b1;
  assign _zz_4015 = _zz_17051;
  assign _zz_4016 = _zz_17059;
  assign _zz_1483 = ($signed(_zz_17067) * $signed(data_mid_88_real));
  assign _zz_4017 = _zz_17068;
  assign _zz_1481 = _zz_17071[31 : 0];
  assign _zz_4018 = _zz_17072;
  assign _zz_1482 = _zz_17075[31 : 0];
  assign _zz_1484 = 1'b1;
  assign _zz_4019 = _zz_17076;
  assign _zz_4020 = _zz_17084;
  assign _zz_1485 = 1'b1;
  assign _zz_4021 = _zz_17092;
  assign _zz_4022 = _zz_17100;
  assign _zz_1488 = ($signed(_zz_17108) * $signed(data_mid_89_real));
  assign _zz_4023 = _zz_17109;
  assign _zz_1486 = _zz_17112[31 : 0];
  assign _zz_4024 = _zz_17113;
  assign _zz_1487 = _zz_17116[31 : 0];
  assign _zz_1489 = 1'b1;
  assign _zz_4025 = _zz_17117;
  assign _zz_4026 = _zz_17125;
  assign _zz_1490 = 1'b1;
  assign _zz_4027 = _zz_17133;
  assign _zz_4028 = _zz_17141;
  assign _zz_1493 = ($signed(_zz_17149) * $signed(data_mid_90_real));
  assign _zz_4029 = _zz_17150;
  assign _zz_1491 = _zz_17153[31 : 0];
  assign _zz_4030 = _zz_17154;
  assign _zz_1492 = _zz_17157[31 : 0];
  assign _zz_1494 = 1'b1;
  assign _zz_4031 = _zz_17158;
  assign _zz_4032 = _zz_17166;
  assign _zz_1495 = 1'b1;
  assign _zz_4033 = _zz_17174;
  assign _zz_4034 = _zz_17182;
  assign _zz_1498 = ($signed(_zz_17190) * $signed(data_mid_91_real));
  assign _zz_4035 = _zz_17191;
  assign _zz_1496 = _zz_17194[31 : 0];
  assign _zz_4036 = _zz_17195;
  assign _zz_1497 = _zz_17198[31 : 0];
  assign _zz_1499 = 1'b1;
  assign _zz_4037 = _zz_17199;
  assign _zz_4038 = _zz_17207;
  assign _zz_1500 = 1'b1;
  assign _zz_4039 = _zz_17215;
  assign _zz_4040 = _zz_17223;
  assign _zz_1503 = ($signed(_zz_17231) * $signed(data_mid_92_real));
  assign _zz_4041 = _zz_17232;
  assign _zz_1501 = _zz_17235[31 : 0];
  assign _zz_4042 = _zz_17236;
  assign _zz_1502 = _zz_17239[31 : 0];
  assign _zz_1504 = 1'b1;
  assign _zz_4043 = _zz_17240;
  assign _zz_4044 = _zz_17248;
  assign _zz_1505 = 1'b1;
  assign _zz_4045 = _zz_17256;
  assign _zz_4046 = _zz_17264;
  assign _zz_1508 = ($signed(_zz_17272) * $signed(data_mid_93_real));
  assign _zz_4047 = _zz_17273;
  assign _zz_1506 = _zz_17276[31 : 0];
  assign _zz_4048 = _zz_17277;
  assign _zz_1507 = _zz_17280[31 : 0];
  assign _zz_1509 = 1'b1;
  assign _zz_4049 = _zz_17281;
  assign _zz_4050 = _zz_17289;
  assign _zz_1510 = 1'b1;
  assign _zz_4051 = _zz_17297;
  assign _zz_4052 = _zz_17305;
  assign _zz_1513 = ($signed(_zz_17313) * $signed(data_mid_94_real));
  assign _zz_4053 = _zz_17314;
  assign _zz_1511 = _zz_17317[31 : 0];
  assign _zz_4054 = _zz_17318;
  assign _zz_1512 = _zz_17321[31 : 0];
  assign _zz_1514 = 1'b1;
  assign _zz_4055 = _zz_17322;
  assign _zz_4056 = _zz_17330;
  assign _zz_1515 = 1'b1;
  assign _zz_4057 = _zz_17338;
  assign _zz_4058 = _zz_17346;
  assign _zz_1518 = ($signed(_zz_17354) * $signed(data_mid_95_real));
  assign _zz_4059 = _zz_17355;
  assign _zz_1516 = _zz_17358[31 : 0];
  assign _zz_4060 = _zz_17359;
  assign _zz_1517 = _zz_17362[31 : 0];
  assign _zz_1519 = 1'b1;
  assign _zz_4061 = _zz_17363;
  assign _zz_4062 = _zz_17371;
  assign _zz_1520 = 1'b1;
  assign _zz_4063 = _zz_17379;
  assign _zz_4064 = _zz_17387;
  assign _zz_1523 = ($signed(_zz_17395) * $signed(data_mid_112_real));
  assign _zz_4065 = _zz_17396;
  assign _zz_1521 = _zz_17399[31 : 0];
  assign _zz_4066 = _zz_17400;
  assign _zz_1522 = _zz_17403[31 : 0];
  assign _zz_1524 = 1'b1;
  assign _zz_4067 = _zz_17404;
  assign _zz_4068 = _zz_17412;
  assign _zz_1525 = 1'b1;
  assign _zz_4069 = _zz_17420;
  assign _zz_4070 = _zz_17428;
  assign _zz_1528 = ($signed(_zz_17436) * $signed(data_mid_113_real));
  assign _zz_4071 = _zz_17437;
  assign _zz_1526 = _zz_17440[31 : 0];
  assign _zz_4072 = _zz_17441;
  assign _zz_1527 = _zz_17444[31 : 0];
  assign _zz_1529 = 1'b1;
  assign _zz_4073 = _zz_17445;
  assign _zz_4074 = _zz_17453;
  assign _zz_1530 = 1'b1;
  assign _zz_4075 = _zz_17461;
  assign _zz_4076 = _zz_17469;
  assign _zz_1533 = ($signed(_zz_17477) * $signed(data_mid_114_real));
  assign _zz_4077 = _zz_17478;
  assign _zz_1531 = _zz_17481[31 : 0];
  assign _zz_4078 = _zz_17482;
  assign _zz_1532 = _zz_17485[31 : 0];
  assign _zz_1534 = 1'b1;
  assign _zz_4079 = _zz_17486;
  assign _zz_4080 = _zz_17494;
  assign _zz_1535 = 1'b1;
  assign _zz_4081 = _zz_17502;
  assign _zz_4082 = _zz_17510;
  assign _zz_1538 = ($signed(_zz_17518) * $signed(data_mid_115_real));
  assign _zz_4083 = _zz_17519;
  assign _zz_1536 = _zz_17522[31 : 0];
  assign _zz_4084 = _zz_17523;
  assign _zz_1537 = _zz_17526[31 : 0];
  assign _zz_1539 = 1'b1;
  assign _zz_4085 = _zz_17527;
  assign _zz_4086 = _zz_17535;
  assign _zz_1540 = 1'b1;
  assign _zz_4087 = _zz_17543;
  assign _zz_4088 = _zz_17551;
  assign _zz_1543 = ($signed(_zz_17559) * $signed(data_mid_116_real));
  assign _zz_4089 = _zz_17560;
  assign _zz_1541 = _zz_17563[31 : 0];
  assign _zz_4090 = _zz_17564;
  assign _zz_1542 = _zz_17567[31 : 0];
  assign _zz_1544 = 1'b1;
  assign _zz_4091 = _zz_17568;
  assign _zz_4092 = _zz_17576;
  assign _zz_1545 = 1'b1;
  assign _zz_4093 = _zz_17584;
  assign _zz_4094 = _zz_17592;
  assign _zz_1548 = ($signed(_zz_17600) * $signed(data_mid_117_real));
  assign _zz_4095 = _zz_17601;
  assign _zz_1546 = _zz_17604[31 : 0];
  assign _zz_4096 = _zz_17605;
  assign _zz_1547 = _zz_17608[31 : 0];
  assign _zz_1549 = 1'b1;
  assign _zz_4097 = _zz_17609;
  assign _zz_4098 = _zz_17617;
  assign _zz_1550 = 1'b1;
  assign _zz_4099 = _zz_17625;
  assign _zz_4100 = _zz_17633;
  assign _zz_1553 = ($signed(_zz_17641) * $signed(data_mid_118_real));
  assign _zz_4101 = _zz_17642;
  assign _zz_1551 = _zz_17645[31 : 0];
  assign _zz_4102 = _zz_17646;
  assign _zz_1552 = _zz_17649[31 : 0];
  assign _zz_1554 = 1'b1;
  assign _zz_4103 = _zz_17650;
  assign _zz_4104 = _zz_17658;
  assign _zz_1555 = 1'b1;
  assign _zz_4105 = _zz_17666;
  assign _zz_4106 = _zz_17674;
  assign _zz_1558 = ($signed(_zz_17682) * $signed(data_mid_119_real));
  assign _zz_4107 = _zz_17683;
  assign _zz_1556 = _zz_17686[31 : 0];
  assign _zz_4108 = _zz_17687;
  assign _zz_1557 = _zz_17690[31 : 0];
  assign _zz_1559 = 1'b1;
  assign _zz_4109 = _zz_17691;
  assign _zz_4110 = _zz_17699;
  assign _zz_1560 = 1'b1;
  assign _zz_4111 = _zz_17707;
  assign _zz_4112 = _zz_17715;
  assign _zz_1563 = ($signed(_zz_17723) * $signed(data_mid_120_real));
  assign _zz_4113 = _zz_17724;
  assign _zz_1561 = _zz_17727[31 : 0];
  assign _zz_4114 = _zz_17728;
  assign _zz_1562 = _zz_17731[31 : 0];
  assign _zz_1564 = 1'b1;
  assign _zz_4115 = _zz_17732;
  assign _zz_4116 = _zz_17740;
  assign _zz_1565 = 1'b1;
  assign _zz_4117 = _zz_17748;
  assign _zz_4118 = _zz_17756;
  assign _zz_1568 = ($signed(_zz_17764) * $signed(data_mid_121_real));
  assign _zz_4119 = _zz_17765;
  assign _zz_1566 = _zz_17768[31 : 0];
  assign _zz_4120 = _zz_17769;
  assign _zz_1567 = _zz_17772[31 : 0];
  assign _zz_1569 = 1'b1;
  assign _zz_4121 = _zz_17773;
  assign _zz_4122 = _zz_17781;
  assign _zz_1570 = 1'b1;
  assign _zz_4123 = _zz_17789;
  assign _zz_4124 = _zz_17797;
  assign _zz_1573 = ($signed(_zz_17805) * $signed(data_mid_122_real));
  assign _zz_4125 = _zz_17806;
  assign _zz_1571 = _zz_17809[31 : 0];
  assign _zz_4126 = _zz_17810;
  assign _zz_1572 = _zz_17813[31 : 0];
  assign _zz_1574 = 1'b1;
  assign _zz_4127 = _zz_17814;
  assign _zz_4128 = _zz_17822;
  assign _zz_1575 = 1'b1;
  assign _zz_4129 = _zz_17830;
  assign _zz_4130 = _zz_17838;
  assign _zz_1578 = ($signed(_zz_17846) * $signed(data_mid_123_real));
  assign _zz_4131 = _zz_17847;
  assign _zz_1576 = _zz_17850[31 : 0];
  assign _zz_4132 = _zz_17851;
  assign _zz_1577 = _zz_17854[31 : 0];
  assign _zz_1579 = 1'b1;
  assign _zz_4133 = _zz_17855;
  assign _zz_4134 = _zz_17863;
  assign _zz_1580 = 1'b1;
  assign _zz_4135 = _zz_17871;
  assign _zz_4136 = _zz_17879;
  assign _zz_1583 = ($signed(_zz_17887) * $signed(data_mid_124_real));
  assign _zz_4137 = _zz_17888;
  assign _zz_1581 = _zz_17891[31 : 0];
  assign _zz_4138 = _zz_17892;
  assign _zz_1582 = _zz_17895[31 : 0];
  assign _zz_1584 = 1'b1;
  assign _zz_4139 = _zz_17896;
  assign _zz_4140 = _zz_17904;
  assign _zz_1585 = 1'b1;
  assign _zz_4141 = _zz_17912;
  assign _zz_4142 = _zz_17920;
  assign _zz_1588 = ($signed(_zz_17928) * $signed(data_mid_125_real));
  assign _zz_4143 = _zz_17929;
  assign _zz_1586 = _zz_17932[31 : 0];
  assign _zz_4144 = _zz_17933;
  assign _zz_1587 = _zz_17936[31 : 0];
  assign _zz_1589 = 1'b1;
  assign _zz_4145 = _zz_17937;
  assign _zz_4146 = _zz_17945;
  assign _zz_1590 = 1'b1;
  assign _zz_4147 = _zz_17953;
  assign _zz_4148 = _zz_17961;
  assign _zz_1593 = ($signed(_zz_17969) * $signed(data_mid_126_real));
  assign _zz_4149 = _zz_17970;
  assign _zz_1591 = _zz_17973[31 : 0];
  assign _zz_4150 = _zz_17974;
  assign _zz_1592 = _zz_17977[31 : 0];
  assign _zz_1594 = 1'b1;
  assign _zz_4151 = _zz_17978;
  assign _zz_4152 = _zz_17986;
  assign _zz_1595 = 1'b1;
  assign _zz_4153 = _zz_17994;
  assign _zz_4154 = _zz_18002;
  assign _zz_1598 = ($signed(_zz_18010) * $signed(data_mid_127_real));
  assign _zz_4155 = _zz_18011;
  assign _zz_1596 = _zz_18014[31 : 0];
  assign _zz_4156 = _zz_18015;
  assign _zz_1597 = _zz_18018[31 : 0];
  assign _zz_1599 = 1'b1;
  assign _zz_4157 = _zz_18019;
  assign _zz_4158 = _zz_18027;
  assign _zz_1600 = 1'b1;
  assign _zz_4159 = _zz_18035;
  assign _zz_4160 = _zz_18043;
  assign _zz_1603 = ($signed(_zz_18051) * $signed(data_mid_32_real));
  assign _zz_4161 = _zz_18052;
  assign _zz_1601 = _zz_18055[31 : 0];
  assign _zz_4162 = _zz_18056;
  assign _zz_1602 = _zz_18059[31 : 0];
  assign _zz_1604 = 1'b1;
  assign _zz_4163 = _zz_18060;
  assign _zz_4164 = _zz_18068;
  assign _zz_1605 = 1'b1;
  assign _zz_4165 = _zz_18076;
  assign _zz_4166 = _zz_18084;
  assign _zz_1608 = ($signed(_zz_18092) * $signed(data_mid_33_real));
  assign _zz_4167 = _zz_18093;
  assign _zz_1606 = _zz_18096[31 : 0];
  assign _zz_4168 = _zz_18097;
  assign _zz_1607 = _zz_18100[31 : 0];
  assign _zz_1609 = 1'b1;
  assign _zz_4169 = _zz_18101;
  assign _zz_4170 = _zz_18109;
  assign _zz_1610 = 1'b1;
  assign _zz_4171 = _zz_18117;
  assign _zz_4172 = _zz_18125;
  assign _zz_1613 = ($signed(_zz_18133) * $signed(data_mid_34_real));
  assign _zz_4173 = _zz_18134;
  assign _zz_1611 = _zz_18137[31 : 0];
  assign _zz_4174 = _zz_18138;
  assign _zz_1612 = _zz_18141[31 : 0];
  assign _zz_1614 = 1'b1;
  assign _zz_4175 = _zz_18142;
  assign _zz_4176 = _zz_18150;
  assign _zz_1615 = 1'b1;
  assign _zz_4177 = _zz_18158;
  assign _zz_4178 = _zz_18166;
  assign _zz_1618 = ($signed(_zz_18174) * $signed(data_mid_35_real));
  assign _zz_4179 = _zz_18175;
  assign _zz_1616 = _zz_18178[31 : 0];
  assign _zz_4180 = _zz_18179;
  assign _zz_1617 = _zz_18182[31 : 0];
  assign _zz_1619 = 1'b1;
  assign _zz_4181 = _zz_18183;
  assign _zz_4182 = _zz_18191;
  assign _zz_1620 = 1'b1;
  assign _zz_4183 = _zz_18199;
  assign _zz_4184 = _zz_18207;
  assign _zz_1623 = ($signed(_zz_18215) * $signed(data_mid_36_real));
  assign _zz_4185 = _zz_18216;
  assign _zz_1621 = _zz_18219[31 : 0];
  assign _zz_4186 = _zz_18220;
  assign _zz_1622 = _zz_18223[31 : 0];
  assign _zz_1624 = 1'b1;
  assign _zz_4187 = _zz_18224;
  assign _zz_4188 = _zz_18232;
  assign _zz_1625 = 1'b1;
  assign _zz_4189 = _zz_18240;
  assign _zz_4190 = _zz_18248;
  assign _zz_1628 = ($signed(_zz_18256) * $signed(data_mid_37_real));
  assign _zz_4191 = _zz_18257;
  assign _zz_1626 = _zz_18260[31 : 0];
  assign _zz_4192 = _zz_18261;
  assign _zz_1627 = _zz_18264[31 : 0];
  assign _zz_1629 = 1'b1;
  assign _zz_4193 = _zz_18265;
  assign _zz_4194 = _zz_18273;
  assign _zz_1630 = 1'b1;
  assign _zz_4195 = _zz_18281;
  assign _zz_4196 = _zz_18289;
  assign _zz_1633 = ($signed(_zz_18297) * $signed(data_mid_38_real));
  assign _zz_4197 = _zz_18298;
  assign _zz_1631 = _zz_18301[31 : 0];
  assign _zz_4198 = _zz_18302;
  assign _zz_1632 = _zz_18305[31 : 0];
  assign _zz_1634 = 1'b1;
  assign _zz_4199 = _zz_18306;
  assign _zz_4200 = _zz_18314;
  assign _zz_1635 = 1'b1;
  assign _zz_4201 = _zz_18322;
  assign _zz_4202 = _zz_18330;
  assign _zz_1638 = ($signed(_zz_18338) * $signed(data_mid_39_real));
  assign _zz_4203 = _zz_18339;
  assign _zz_1636 = _zz_18342[31 : 0];
  assign _zz_4204 = _zz_18343;
  assign _zz_1637 = _zz_18346[31 : 0];
  assign _zz_1639 = 1'b1;
  assign _zz_4205 = _zz_18347;
  assign _zz_4206 = _zz_18355;
  assign _zz_1640 = 1'b1;
  assign _zz_4207 = _zz_18363;
  assign _zz_4208 = _zz_18371;
  assign _zz_1643 = ($signed(_zz_18379) * $signed(data_mid_40_real));
  assign _zz_4209 = _zz_18380;
  assign _zz_1641 = _zz_18383[31 : 0];
  assign _zz_4210 = _zz_18384;
  assign _zz_1642 = _zz_18387[31 : 0];
  assign _zz_1644 = 1'b1;
  assign _zz_4211 = _zz_18388;
  assign _zz_4212 = _zz_18396;
  assign _zz_1645 = 1'b1;
  assign _zz_4213 = _zz_18404;
  assign _zz_4214 = _zz_18412;
  assign _zz_1648 = ($signed(_zz_18420) * $signed(data_mid_41_real));
  assign _zz_4215 = _zz_18421;
  assign _zz_1646 = _zz_18424[31 : 0];
  assign _zz_4216 = _zz_18425;
  assign _zz_1647 = _zz_18428[31 : 0];
  assign _zz_1649 = 1'b1;
  assign _zz_4217 = _zz_18429;
  assign _zz_4218 = _zz_18437;
  assign _zz_1650 = 1'b1;
  assign _zz_4219 = _zz_18445;
  assign _zz_4220 = _zz_18453;
  assign _zz_1653 = ($signed(_zz_18461) * $signed(data_mid_42_real));
  assign _zz_4221 = _zz_18462;
  assign _zz_1651 = _zz_18465[31 : 0];
  assign _zz_4222 = _zz_18466;
  assign _zz_1652 = _zz_18469[31 : 0];
  assign _zz_1654 = 1'b1;
  assign _zz_4223 = _zz_18470;
  assign _zz_4224 = _zz_18478;
  assign _zz_1655 = 1'b1;
  assign _zz_4225 = _zz_18486;
  assign _zz_4226 = _zz_18494;
  assign _zz_1658 = ($signed(_zz_18502) * $signed(data_mid_43_real));
  assign _zz_4227 = _zz_18503;
  assign _zz_1656 = _zz_18506[31 : 0];
  assign _zz_4228 = _zz_18507;
  assign _zz_1657 = _zz_18510[31 : 0];
  assign _zz_1659 = 1'b1;
  assign _zz_4229 = _zz_18511;
  assign _zz_4230 = _zz_18519;
  assign _zz_1660 = 1'b1;
  assign _zz_4231 = _zz_18527;
  assign _zz_4232 = _zz_18535;
  assign _zz_1663 = ($signed(_zz_18543) * $signed(data_mid_44_real));
  assign _zz_4233 = _zz_18544;
  assign _zz_1661 = _zz_18547[31 : 0];
  assign _zz_4234 = _zz_18548;
  assign _zz_1662 = _zz_18551[31 : 0];
  assign _zz_1664 = 1'b1;
  assign _zz_4235 = _zz_18552;
  assign _zz_4236 = _zz_18560;
  assign _zz_1665 = 1'b1;
  assign _zz_4237 = _zz_18568;
  assign _zz_4238 = _zz_18576;
  assign _zz_1668 = ($signed(_zz_18584) * $signed(data_mid_45_real));
  assign _zz_4239 = _zz_18585;
  assign _zz_1666 = _zz_18588[31 : 0];
  assign _zz_4240 = _zz_18589;
  assign _zz_1667 = _zz_18592[31 : 0];
  assign _zz_1669 = 1'b1;
  assign _zz_4241 = _zz_18593;
  assign _zz_4242 = _zz_18601;
  assign _zz_1670 = 1'b1;
  assign _zz_4243 = _zz_18609;
  assign _zz_4244 = _zz_18617;
  assign _zz_1673 = ($signed(_zz_18625) * $signed(data_mid_46_real));
  assign _zz_4245 = _zz_18626;
  assign _zz_1671 = _zz_18629[31 : 0];
  assign _zz_4246 = _zz_18630;
  assign _zz_1672 = _zz_18633[31 : 0];
  assign _zz_1674 = 1'b1;
  assign _zz_4247 = _zz_18634;
  assign _zz_4248 = _zz_18642;
  assign _zz_1675 = 1'b1;
  assign _zz_4249 = _zz_18650;
  assign _zz_4250 = _zz_18658;
  assign _zz_1678 = ($signed(_zz_18666) * $signed(data_mid_47_real));
  assign _zz_4251 = _zz_18667;
  assign _zz_1676 = _zz_18670[31 : 0];
  assign _zz_4252 = _zz_18671;
  assign _zz_1677 = _zz_18674[31 : 0];
  assign _zz_1679 = 1'b1;
  assign _zz_4253 = _zz_18675;
  assign _zz_4254 = _zz_18683;
  assign _zz_1680 = 1'b1;
  assign _zz_4255 = _zz_18691;
  assign _zz_4256 = _zz_18699;
  assign _zz_1683 = ($signed(_zz_18707) * $signed(data_mid_48_real));
  assign _zz_4257 = _zz_18708;
  assign _zz_1681 = _zz_18711[31 : 0];
  assign _zz_4258 = _zz_18712;
  assign _zz_1682 = _zz_18715[31 : 0];
  assign _zz_1684 = 1'b1;
  assign _zz_4259 = _zz_18716;
  assign _zz_4260 = _zz_18724;
  assign _zz_1685 = 1'b1;
  assign _zz_4261 = _zz_18732;
  assign _zz_4262 = _zz_18740;
  assign _zz_1688 = ($signed(_zz_18748) * $signed(data_mid_49_real));
  assign _zz_4263 = _zz_18749;
  assign _zz_1686 = _zz_18752[31 : 0];
  assign _zz_4264 = _zz_18753;
  assign _zz_1687 = _zz_18756[31 : 0];
  assign _zz_1689 = 1'b1;
  assign _zz_4265 = _zz_18757;
  assign _zz_4266 = _zz_18765;
  assign _zz_1690 = 1'b1;
  assign _zz_4267 = _zz_18773;
  assign _zz_4268 = _zz_18781;
  assign _zz_1693 = ($signed(_zz_18789) * $signed(data_mid_50_real));
  assign _zz_4269 = _zz_18790;
  assign _zz_1691 = _zz_18793[31 : 0];
  assign _zz_4270 = _zz_18794;
  assign _zz_1692 = _zz_18797[31 : 0];
  assign _zz_1694 = 1'b1;
  assign _zz_4271 = _zz_18798;
  assign _zz_4272 = _zz_18806;
  assign _zz_1695 = 1'b1;
  assign _zz_4273 = _zz_18814;
  assign _zz_4274 = _zz_18822;
  assign _zz_1698 = ($signed(_zz_18830) * $signed(data_mid_51_real));
  assign _zz_4275 = _zz_18831;
  assign _zz_1696 = _zz_18834[31 : 0];
  assign _zz_4276 = _zz_18835;
  assign _zz_1697 = _zz_18838[31 : 0];
  assign _zz_1699 = 1'b1;
  assign _zz_4277 = _zz_18839;
  assign _zz_4278 = _zz_18847;
  assign _zz_1700 = 1'b1;
  assign _zz_4279 = _zz_18855;
  assign _zz_4280 = _zz_18863;
  assign _zz_1703 = ($signed(_zz_18871) * $signed(data_mid_52_real));
  assign _zz_4281 = _zz_18872;
  assign _zz_1701 = _zz_18875[31 : 0];
  assign _zz_4282 = _zz_18876;
  assign _zz_1702 = _zz_18879[31 : 0];
  assign _zz_1704 = 1'b1;
  assign _zz_4283 = _zz_18880;
  assign _zz_4284 = _zz_18888;
  assign _zz_1705 = 1'b1;
  assign _zz_4285 = _zz_18896;
  assign _zz_4286 = _zz_18904;
  assign _zz_1708 = ($signed(_zz_18912) * $signed(data_mid_53_real));
  assign _zz_4287 = _zz_18913;
  assign _zz_1706 = _zz_18916[31 : 0];
  assign _zz_4288 = _zz_18917;
  assign _zz_1707 = _zz_18920[31 : 0];
  assign _zz_1709 = 1'b1;
  assign _zz_4289 = _zz_18921;
  assign _zz_4290 = _zz_18929;
  assign _zz_1710 = 1'b1;
  assign _zz_4291 = _zz_18937;
  assign _zz_4292 = _zz_18945;
  assign _zz_1713 = ($signed(_zz_18953) * $signed(data_mid_54_real));
  assign _zz_4293 = _zz_18954;
  assign _zz_1711 = _zz_18957[31 : 0];
  assign _zz_4294 = _zz_18958;
  assign _zz_1712 = _zz_18961[31 : 0];
  assign _zz_1714 = 1'b1;
  assign _zz_4295 = _zz_18962;
  assign _zz_4296 = _zz_18970;
  assign _zz_1715 = 1'b1;
  assign _zz_4297 = _zz_18978;
  assign _zz_4298 = _zz_18986;
  assign _zz_1718 = ($signed(_zz_18994) * $signed(data_mid_55_real));
  assign _zz_4299 = _zz_18995;
  assign _zz_1716 = _zz_18998[31 : 0];
  assign _zz_4300 = _zz_18999;
  assign _zz_1717 = _zz_19002[31 : 0];
  assign _zz_1719 = 1'b1;
  assign _zz_4301 = _zz_19003;
  assign _zz_4302 = _zz_19011;
  assign _zz_1720 = 1'b1;
  assign _zz_4303 = _zz_19019;
  assign _zz_4304 = _zz_19027;
  assign _zz_1723 = ($signed(_zz_19035) * $signed(data_mid_56_real));
  assign _zz_4305 = _zz_19036;
  assign _zz_1721 = _zz_19039[31 : 0];
  assign _zz_4306 = _zz_19040;
  assign _zz_1722 = _zz_19043[31 : 0];
  assign _zz_1724 = 1'b1;
  assign _zz_4307 = _zz_19044;
  assign _zz_4308 = _zz_19052;
  assign _zz_1725 = 1'b1;
  assign _zz_4309 = _zz_19060;
  assign _zz_4310 = _zz_19068;
  assign _zz_1728 = ($signed(_zz_19076) * $signed(data_mid_57_real));
  assign _zz_4311 = _zz_19077;
  assign _zz_1726 = _zz_19080[31 : 0];
  assign _zz_4312 = _zz_19081;
  assign _zz_1727 = _zz_19084[31 : 0];
  assign _zz_1729 = 1'b1;
  assign _zz_4313 = _zz_19085;
  assign _zz_4314 = _zz_19093;
  assign _zz_1730 = 1'b1;
  assign _zz_4315 = _zz_19101;
  assign _zz_4316 = _zz_19109;
  assign _zz_1733 = ($signed(_zz_19117) * $signed(data_mid_58_real));
  assign _zz_4317 = _zz_19118;
  assign _zz_1731 = _zz_19121[31 : 0];
  assign _zz_4318 = _zz_19122;
  assign _zz_1732 = _zz_19125[31 : 0];
  assign _zz_1734 = 1'b1;
  assign _zz_4319 = _zz_19126;
  assign _zz_4320 = _zz_19134;
  assign _zz_1735 = 1'b1;
  assign _zz_4321 = _zz_19142;
  assign _zz_4322 = _zz_19150;
  assign _zz_1738 = ($signed(_zz_19158) * $signed(data_mid_59_real));
  assign _zz_4323 = _zz_19159;
  assign _zz_1736 = _zz_19162[31 : 0];
  assign _zz_4324 = _zz_19163;
  assign _zz_1737 = _zz_19166[31 : 0];
  assign _zz_1739 = 1'b1;
  assign _zz_4325 = _zz_19167;
  assign _zz_4326 = _zz_19175;
  assign _zz_1740 = 1'b1;
  assign _zz_4327 = _zz_19183;
  assign _zz_4328 = _zz_19191;
  assign _zz_1743 = ($signed(_zz_19199) * $signed(data_mid_60_real));
  assign _zz_4329 = _zz_19200;
  assign _zz_1741 = _zz_19203[31 : 0];
  assign _zz_4330 = _zz_19204;
  assign _zz_1742 = _zz_19207[31 : 0];
  assign _zz_1744 = 1'b1;
  assign _zz_4331 = _zz_19208;
  assign _zz_4332 = _zz_19216;
  assign _zz_1745 = 1'b1;
  assign _zz_4333 = _zz_19224;
  assign _zz_4334 = _zz_19232;
  assign _zz_1748 = ($signed(_zz_19240) * $signed(data_mid_61_real));
  assign _zz_4335 = _zz_19241;
  assign _zz_1746 = _zz_19244[31 : 0];
  assign _zz_4336 = _zz_19245;
  assign _zz_1747 = _zz_19248[31 : 0];
  assign _zz_1749 = 1'b1;
  assign _zz_4337 = _zz_19249;
  assign _zz_4338 = _zz_19257;
  assign _zz_1750 = 1'b1;
  assign _zz_4339 = _zz_19265;
  assign _zz_4340 = _zz_19273;
  assign _zz_1753 = ($signed(_zz_19281) * $signed(data_mid_62_real));
  assign _zz_4341 = _zz_19282;
  assign _zz_1751 = _zz_19285[31 : 0];
  assign _zz_4342 = _zz_19286;
  assign _zz_1752 = _zz_19289[31 : 0];
  assign _zz_1754 = 1'b1;
  assign _zz_4343 = _zz_19290;
  assign _zz_4344 = _zz_19298;
  assign _zz_1755 = 1'b1;
  assign _zz_4345 = _zz_19306;
  assign _zz_4346 = _zz_19314;
  assign _zz_1758 = ($signed(_zz_19322) * $signed(data_mid_63_real));
  assign _zz_4347 = _zz_19323;
  assign _zz_1756 = _zz_19326[31 : 0];
  assign _zz_4348 = _zz_19327;
  assign _zz_1757 = _zz_19330[31 : 0];
  assign _zz_1759 = 1'b1;
  assign _zz_4349 = _zz_19331;
  assign _zz_4350 = _zz_19339;
  assign _zz_1760 = 1'b1;
  assign _zz_4351 = _zz_19347;
  assign _zz_4352 = _zz_19355;
  assign _zz_1763 = ($signed(_zz_19363) * $signed(data_mid_96_real));
  assign _zz_4353 = _zz_19364;
  assign _zz_1761 = _zz_19367[31 : 0];
  assign _zz_4354 = _zz_19368;
  assign _zz_1762 = _zz_19371[31 : 0];
  assign _zz_1764 = 1'b1;
  assign _zz_4355 = _zz_19372;
  assign _zz_4356 = _zz_19380;
  assign _zz_1765 = 1'b1;
  assign _zz_4357 = _zz_19388;
  assign _zz_4358 = _zz_19396;
  assign _zz_1768 = ($signed(_zz_19404) * $signed(data_mid_97_real));
  assign _zz_4359 = _zz_19405;
  assign _zz_1766 = _zz_19408[31 : 0];
  assign _zz_4360 = _zz_19409;
  assign _zz_1767 = _zz_19412[31 : 0];
  assign _zz_1769 = 1'b1;
  assign _zz_4361 = _zz_19413;
  assign _zz_4362 = _zz_19421;
  assign _zz_1770 = 1'b1;
  assign _zz_4363 = _zz_19429;
  assign _zz_4364 = _zz_19437;
  assign _zz_1773 = ($signed(_zz_19445) * $signed(data_mid_98_real));
  assign _zz_4365 = _zz_19446;
  assign _zz_1771 = _zz_19449[31 : 0];
  assign _zz_4366 = _zz_19450;
  assign _zz_1772 = _zz_19453[31 : 0];
  assign _zz_1774 = 1'b1;
  assign _zz_4367 = _zz_19454;
  assign _zz_4368 = _zz_19462;
  assign _zz_1775 = 1'b1;
  assign _zz_4369 = _zz_19470;
  assign _zz_4370 = _zz_19478;
  assign _zz_1778 = ($signed(_zz_19486) * $signed(data_mid_99_real));
  assign _zz_4371 = _zz_19487;
  assign _zz_1776 = _zz_19490[31 : 0];
  assign _zz_4372 = _zz_19491;
  assign _zz_1777 = _zz_19494[31 : 0];
  assign _zz_1779 = 1'b1;
  assign _zz_4373 = _zz_19495;
  assign _zz_4374 = _zz_19503;
  assign _zz_1780 = 1'b1;
  assign _zz_4375 = _zz_19511;
  assign _zz_4376 = _zz_19519;
  assign _zz_1783 = ($signed(_zz_19527) * $signed(data_mid_100_real));
  assign _zz_4377 = _zz_19528;
  assign _zz_1781 = _zz_19531[31 : 0];
  assign _zz_4378 = _zz_19532;
  assign _zz_1782 = _zz_19535[31 : 0];
  assign _zz_1784 = 1'b1;
  assign _zz_4379 = _zz_19536;
  assign _zz_4380 = _zz_19544;
  assign _zz_1785 = 1'b1;
  assign _zz_4381 = _zz_19552;
  assign _zz_4382 = _zz_19560;
  assign _zz_1788 = ($signed(_zz_19568) * $signed(data_mid_101_real));
  assign _zz_4383 = _zz_19569;
  assign _zz_1786 = _zz_19572[31 : 0];
  assign _zz_4384 = _zz_19573;
  assign _zz_1787 = _zz_19576[31 : 0];
  assign _zz_1789 = 1'b1;
  assign _zz_4385 = _zz_19577;
  assign _zz_4386 = _zz_19585;
  assign _zz_1790 = 1'b1;
  assign _zz_4387 = _zz_19593;
  assign _zz_4388 = _zz_19601;
  assign _zz_1793 = ($signed(_zz_19609) * $signed(data_mid_102_real));
  assign _zz_4389 = _zz_19610;
  assign _zz_1791 = _zz_19613[31 : 0];
  assign _zz_4390 = _zz_19614;
  assign _zz_1792 = _zz_19617[31 : 0];
  assign _zz_1794 = 1'b1;
  assign _zz_4391 = _zz_19618;
  assign _zz_4392 = _zz_19626;
  assign _zz_1795 = 1'b1;
  assign _zz_4393 = _zz_19634;
  assign _zz_4394 = _zz_19642;
  assign _zz_1798 = ($signed(_zz_19650) * $signed(data_mid_103_real));
  assign _zz_4395 = _zz_19651;
  assign _zz_1796 = _zz_19654[31 : 0];
  assign _zz_4396 = _zz_19655;
  assign _zz_1797 = _zz_19658[31 : 0];
  assign _zz_1799 = 1'b1;
  assign _zz_4397 = _zz_19659;
  assign _zz_4398 = _zz_19667;
  assign _zz_1800 = 1'b1;
  assign _zz_4399 = _zz_19675;
  assign _zz_4400 = _zz_19683;
  assign _zz_1803 = ($signed(_zz_19691) * $signed(data_mid_104_real));
  assign _zz_4401 = _zz_19692;
  assign _zz_1801 = _zz_19695[31 : 0];
  assign _zz_4402 = _zz_19696;
  assign _zz_1802 = _zz_19699[31 : 0];
  assign _zz_1804 = 1'b1;
  assign _zz_4403 = _zz_19700;
  assign _zz_4404 = _zz_19708;
  assign _zz_1805 = 1'b1;
  assign _zz_4405 = _zz_19716;
  assign _zz_4406 = _zz_19724;
  assign _zz_1808 = ($signed(_zz_19732) * $signed(data_mid_105_real));
  assign _zz_4407 = _zz_19733;
  assign _zz_1806 = _zz_19736[31 : 0];
  assign _zz_4408 = _zz_19737;
  assign _zz_1807 = _zz_19740[31 : 0];
  assign _zz_1809 = 1'b1;
  assign _zz_4409 = _zz_19741;
  assign _zz_4410 = _zz_19749;
  assign _zz_1810 = 1'b1;
  assign _zz_4411 = _zz_19757;
  assign _zz_4412 = _zz_19765;
  assign _zz_1813 = ($signed(_zz_19773) * $signed(data_mid_106_real));
  assign _zz_4413 = _zz_19774;
  assign _zz_1811 = _zz_19777[31 : 0];
  assign _zz_4414 = _zz_19778;
  assign _zz_1812 = _zz_19781[31 : 0];
  assign _zz_1814 = 1'b1;
  assign _zz_4415 = _zz_19782;
  assign _zz_4416 = _zz_19790;
  assign _zz_1815 = 1'b1;
  assign _zz_4417 = _zz_19798;
  assign _zz_4418 = _zz_19806;
  assign _zz_1818 = ($signed(_zz_19814) * $signed(data_mid_107_real));
  assign _zz_4419 = _zz_19815;
  assign _zz_1816 = _zz_19818[31 : 0];
  assign _zz_4420 = _zz_19819;
  assign _zz_1817 = _zz_19822[31 : 0];
  assign _zz_1819 = 1'b1;
  assign _zz_4421 = _zz_19823;
  assign _zz_4422 = _zz_19831;
  assign _zz_1820 = 1'b1;
  assign _zz_4423 = _zz_19839;
  assign _zz_4424 = _zz_19847;
  assign _zz_1823 = ($signed(_zz_19855) * $signed(data_mid_108_real));
  assign _zz_4425 = _zz_19856;
  assign _zz_1821 = _zz_19859[31 : 0];
  assign _zz_4426 = _zz_19860;
  assign _zz_1822 = _zz_19863[31 : 0];
  assign _zz_1824 = 1'b1;
  assign _zz_4427 = _zz_19864;
  assign _zz_4428 = _zz_19872;
  assign _zz_1825 = 1'b1;
  assign _zz_4429 = _zz_19880;
  assign _zz_4430 = _zz_19888;
  assign _zz_1828 = ($signed(_zz_19896) * $signed(data_mid_109_real));
  assign _zz_4431 = _zz_19897;
  assign _zz_1826 = _zz_19900[31 : 0];
  assign _zz_4432 = _zz_19901;
  assign _zz_1827 = _zz_19904[31 : 0];
  assign _zz_1829 = 1'b1;
  assign _zz_4433 = _zz_19905;
  assign _zz_4434 = _zz_19913;
  assign _zz_1830 = 1'b1;
  assign _zz_4435 = _zz_19921;
  assign _zz_4436 = _zz_19929;
  assign _zz_1833 = ($signed(_zz_19937) * $signed(data_mid_110_real));
  assign _zz_4437 = _zz_19938;
  assign _zz_1831 = _zz_19941[31 : 0];
  assign _zz_4438 = _zz_19942;
  assign _zz_1832 = _zz_19945[31 : 0];
  assign _zz_1834 = 1'b1;
  assign _zz_4439 = _zz_19946;
  assign _zz_4440 = _zz_19954;
  assign _zz_1835 = 1'b1;
  assign _zz_4441 = _zz_19962;
  assign _zz_4442 = _zz_19970;
  assign _zz_1838 = ($signed(_zz_19978) * $signed(data_mid_111_real));
  assign _zz_4443 = _zz_19979;
  assign _zz_1836 = _zz_19982[31 : 0];
  assign _zz_4444 = _zz_19983;
  assign _zz_1837 = _zz_19986[31 : 0];
  assign _zz_1839 = 1'b1;
  assign _zz_4445 = _zz_19987;
  assign _zz_4446 = _zz_19995;
  assign _zz_1840 = 1'b1;
  assign _zz_4447 = _zz_20003;
  assign _zz_4448 = _zz_20011;
  assign _zz_1843 = ($signed(_zz_20019) * $signed(data_mid_112_real));
  assign _zz_4449 = _zz_20020;
  assign _zz_1841 = _zz_20023[31 : 0];
  assign _zz_4450 = _zz_20024;
  assign _zz_1842 = _zz_20027[31 : 0];
  assign _zz_1844 = 1'b1;
  assign _zz_4451 = _zz_20028;
  assign _zz_4452 = _zz_20036;
  assign _zz_1845 = 1'b1;
  assign _zz_4453 = _zz_20044;
  assign _zz_4454 = _zz_20052;
  assign _zz_1848 = ($signed(_zz_20060) * $signed(data_mid_113_real));
  assign _zz_4455 = _zz_20061;
  assign _zz_1846 = _zz_20064[31 : 0];
  assign _zz_4456 = _zz_20065;
  assign _zz_1847 = _zz_20068[31 : 0];
  assign _zz_1849 = 1'b1;
  assign _zz_4457 = _zz_20069;
  assign _zz_4458 = _zz_20077;
  assign _zz_1850 = 1'b1;
  assign _zz_4459 = _zz_20085;
  assign _zz_4460 = _zz_20093;
  assign _zz_1853 = ($signed(_zz_20101) * $signed(data_mid_114_real));
  assign _zz_4461 = _zz_20102;
  assign _zz_1851 = _zz_20105[31 : 0];
  assign _zz_4462 = _zz_20106;
  assign _zz_1852 = _zz_20109[31 : 0];
  assign _zz_1854 = 1'b1;
  assign _zz_4463 = _zz_20110;
  assign _zz_4464 = _zz_20118;
  assign _zz_1855 = 1'b1;
  assign _zz_4465 = _zz_20126;
  assign _zz_4466 = _zz_20134;
  assign _zz_1858 = ($signed(_zz_20142) * $signed(data_mid_115_real));
  assign _zz_4467 = _zz_20143;
  assign _zz_1856 = _zz_20146[31 : 0];
  assign _zz_4468 = _zz_20147;
  assign _zz_1857 = _zz_20150[31 : 0];
  assign _zz_1859 = 1'b1;
  assign _zz_4469 = _zz_20151;
  assign _zz_4470 = _zz_20159;
  assign _zz_1860 = 1'b1;
  assign _zz_4471 = _zz_20167;
  assign _zz_4472 = _zz_20175;
  assign _zz_1863 = ($signed(_zz_20183) * $signed(data_mid_116_real));
  assign _zz_4473 = _zz_20184;
  assign _zz_1861 = _zz_20187[31 : 0];
  assign _zz_4474 = _zz_20188;
  assign _zz_1862 = _zz_20191[31 : 0];
  assign _zz_1864 = 1'b1;
  assign _zz_4475 = _zz_20192;
  assign _zz_4476 = _zz_20200;
  assign _zz_1865 = 1'b1;
  assign _zz_4477 = _zz_20208;
  assign _zz_4478 = _zz_20216;
  assign _zz_1868 = ($signed(_zz_20224) * $signed(data_mid_117_real));
  assign _zz_4479 = _zz_20225;
  assign _zz_1866 = _zz_20228[31 : 0];
  assign _zz_4480 = _zz_20229;
  assign _zz_1867 = _zz_20232[31 : 0];
  assign _zz_1869 = 1'b1;
  assign _zz_4481 = _zz_20233;
  assign _zz_4482 = _zz_20241;
  assign _zz_1870 = 1'b1;
  assign _zz_4483 = _zz_20249;
  assign _zz_4484 = _zz_20257;
  assign _zz_1873 = ($signed(_zz_20265) * $signed(data_mid_118_real));
  assign _zz_4485 = _zz_20266;
  assign _zz_1871 = _zz_20269[31 : 0];
  assign _zz_4486 = _zz_20270;
  assign _zz_1872 = _zz_20273[31 : 0];
  assign _zz_1874 = 1'b1;
  assign _zz_4487 = _zz_20274;
  assign _zz_4488 = _zz_20282;
  assign _zz_1875 = 1'b1;
  assign _zz_4489 = _zz_20290;
  assign _zz_4490 = _zz_20298;
  assign _zz_1878 = ($signed(_zz_20306) * $signed(data_mid_119_real));
  assign _zz_4491 = _zz_20307;
  assign _zz_1876 = _zz_20310[31 : 0];
  assign _zz_4492 = _zz_20311;
  assign _zz_1877 = _zz_20314[31 : 0];
  assign _zz_1879 = 1'b1;
  assign _zz_4493 = _zz_20315;
  assign _zz_4494 = _zz_20323;
  assign _zz_1880 = 1'b1;
  assign _zz_4495 = _zz_20331;
  assign _zz_4496 = _zz_20339;
  assign _zz_1883 = ($signed(_zz_20347) * $signed(data_mid_120_real));
  assign _zz_4497 = _zz_20348;
  assign _zz_1881 = _zz_20351[31 : 0];
  assign _zz_4498 = _zz_20352;
  assign _zz_1882 = _zz_20355[31 : 0];
  assign _zz_1884 = 1'b1;
  assign _zz_4499 = _zz_20356;
  assign _zz_4500 = _zz_20364;
  assign _zz_1885 = 1'b1;
  assign _zz_4501 = _zz_20372;
  assign _zz_4502 = _zz_20380;
  assign _zz_1888 = ($signed(_zz_20388) * $signed(data_mid_121_real));
  assign _zz_4503 = _zz_20389;
  assign _zz_1886 = _zz_20392[31 : 0];
  assign _zz_4504 = _zz_20393;
  assign _zz_1887 = _zz_20396[31 : 0];
  assign _zz_1889 = 1'b1;
  assign _zz_4505 = _zz_20397;
  assign _zz_4506 = _zz_20405;
  assign _zz_1890 = 1'b1;
  assign _zz_4507 = _zz_20413;
  assign _zz_4508 = _zz_20421;
  assign _zz_1893 = ($signed(_zz_20429) * $signed(data_mid_122_real));
  assign _zz_4509 = _zz_20430;
  assign _zz_1891 = _zz_20433[31 : 0];
  assign _zz_4510 = _zz_20434;
  assign _zz_1892 = _zz_20437[31 : 0];
  assign _zz_1894 = 1'b1;
  assign _zz_4511 = _zz_20438;
  assign _zz_4512 = _zz_20446;
  assign _zz_1895 = 1'b1;
  assign _zz_4513 = _zz_20454;
  assign _zz_4514 = _zz_20462;
  assign _zz_1898 = ($signed(_zz_20470) * $signed(data_mid_123_real));
  assign _zz_4515 = _zz_20471;
  assign _zz_1896 = _zz_20474[31 : 0];
  assign _zz_4516 = _zz_20475;
  assign _zz_1897 = _zz_20478[31 : 0];
  assign _zz_1899 = 1'b1;
  assign _zz_4517 = _zz_20479;
  assign _zz_4518 = _zz_20487;
  assign _zz_1900 = 1'b1;
  assign _zz_4519 = _zz_20495;
  assign _zz_4520 = _zz_20503;
  assign _zz_1903 = ($signed(_zz_20511) * $signed(data_mid_124_real));
  assign _zz_4521 = _zz_20512;
  assign _zz_1901 = _zz_20515[31 : 0];
  assign _zz_4522 = _zz_20516;
  assign _zz_1902 = _zz_20519[31 : 0];
  assign _zz_1904 = 1'b1;
  assign _zz_4523 = _zz_20520;
  assign _zz_4524 = _zz_20528;
  assign _zz_1905 = 1'b1;
  assign _zz_4525 = _zz_20536;
  assign _zz_4526 = _zz_20544;
  assign _zz_1908 = ($signed(_zz_20552) * $signed(data_mid_125_real));
  assign _zz_4527 = _zz_20553;
  assign _zz_1906 = _zz_20556[31 : 0];
  assign _zz_4528 = _zz_20557;
  assign _zz_1907 = _zz_20560[31 : 0];
  assign _zz_1909 = 1'b1;
  assign _zz_4529 = _zz_20561;
  assign _zz_4530 = _zz_20569;
  assign _zz_1910 = 1'b1;
  assign _zz_4531 = _zz_20577;
  assign _zz_4532 = _zz_20585;
  assign _zz_1913 = ($signed(_zz_20593) * $signed(data_mid_126_real));
  assign _zz_4533 = _zz_20594;
  assign _zz_1911 = _zz_20597[31 : 0];
  assign _zz_4534 = _zz_20598;
  assign _zz_1912 = _zz_20601[31 : 0];
  assign _zz_1914 = 1'b1;
  assign _zz_4535 = _zz_20602;
  assign _zz_4536 = _zz_20610;
  assign _zz_1915 = 1'b1;
  assign _zz_4537 = _zz_20618;
  assign _zz_4538 = _zz_20626;
  assign _zz_1918 = ($signed(_zz_20634) * $signed(data_mid_127_real));
  assign _zz_4539 = _zz_20635;
  assign _zz_1916 = _zz_20638[31 : 0];
  assign _zz_4540 = _zz_20639;
  assign _zz_1917 = _zz_20642[31 : 0];
  assign _zz_1919 = 1'b1;
  assign _zz_4541 = _zz_20643;
  assign _zz_4542 = _zz_20651;
  assign _zz_1920 = 1'b1;
  assign _zz_4543 = _zz_20659;
  assign _zz_4544 = _zz_20667;
  assign _zz_1923 = ($signed(_zz_20675) * $signed(data_mid_64_real));
  assign _zz_4545 = _zz_20676;
  assign _zz_1921 = _zz_20679[31 : 0];
  assign _zz_4546 = _zz_20680;
  assign _zz_1922 = _zz_20683[31 : 0];
  assign _zz_1924 = 1'b1;
  assign _zz_4547 = _zz_20684;
  assign _zz_4548 = _zz_20692;
  assign _zz_1925 = 1'b1;
  assign _zz_4549 = _zz_20700;
  assign _zz_4550 = _zz_20708;
  assign _zz_1928 = ($signed(_zz_20716) * $signed(data_mid_65_real));
  assign _zz_4551 = _zz_20717;
  assign _zz_1926 = _zz_20720[31 : 0];
  assign _zz_4552 = _zz_20721;
  assign _zz_1927 = _zz_20724[31 : 0];
  assign _zz_1929 = 1'b1;
  assign _zz_4553 = _zz_20725;
  assign _zz_4554 = _zz_20733;
  assign _zz_1930 = 1'b1;
  assign _zz_4555 = _zz_20741;
  assign _zz_4556 = _zz_20749;
  assign _zz_1933 = ($signed(_zz_20757) * $signed(data_mid_66_real));
  assign _zz_4557 = _zz_20758;
  assign _zz_1931 = _zz_20761[31 : 0];
  assign _zz_4558 = _zz_20762;
  assign _zz_1932 = _zz_20765[31 : 0];
  assign _zz_1934 = 1'b1;
  assign _zz_4559 = _zz_20766;
  assign _zz_4560 = _zz_20774;
  assign _zz_1935 = 1'b1;
  assign _zz_4561 = _zz_20782;
  assign _zz_4562 = _zz_20790;
  assign _zz_1938 = ($signed(_zz_20798) * $signed(data_mid_67_real));
  assign _zz_4563 = _zz_20799;
  assign _zz_1936 = _zz_20802[31 : 0];
  assign _zz_4564 = _zz_20803;
  assign _zz_1937 = _zz_20806[31 : 0];
  assign _zz_1939 = 1'b1;
  assign _zz_4565 = _zz_20807;
  assign _zz_4566 = _zz_20815;
  assign _zz_1940 = 1'b1;
  assign _zz_4567 = _zz_20823;
  assign _zz_4568 = _zz_20831;
  assign _zz_1943 = ($signed(_zz_20839) * $signed(data_mid_68_real));
  assign _zz_4569 = _zz_20840;
  assign _zz_1941 = _zz_20843[31 : 0];
  assign _zz_4570 = _zz_20844;
  assign _zz_1942 = _zz_20847[31 : 0];
  assign _zz_1944 = 1'b1;
  assign _zz_4571 = _zz_20848;
  assign _zz_4572 = _zz_20856;
  assign _zz_1945 = 1'b1;
  assign _zz_4573 = _zz_20864;
  assign _zz_4574 = _zz_20872;
  assign _zz_1948 = ($signed(_zz_20880) * $signed(data_mid_69_real));
  assign _zz_4575 = _zz_20881;
  assign _zz_1946 = _zz_20884[31 : 0];
  assign _zz_4576 = _zz_20885;
  assign _zz_1947 = _zz_20888[31 : 0];
  assign _zz_1949 = 1'b1;
  assign _zz_4577 = _zz_20889;
  assign _zz_4578 = _zz_20897;
  assign _zz_1950 = 1'b1;
  assign _zz_4579 = _zz_20905;
  assign _zz_4580 = _zz_20913;
  assign _zz_1953 = ($signed(_zz_20921) * $signed(data_mid_70_real));
  assign _zz_4581 = _zz_20922;
  assign _zz_1951 = _zz_20925[31 : 0];
  assign _zz_4582 = _zz_20926;
  assign _zz_1952 = _zz_20929[31 : 0];
  assign _zz_1954 = 1'b1;
  assign _zz_4583 = _zz_20930;
  assign _zz_4584 = _zz_20938;
  assign _zz_1955 = 1'b1;
  assign _zz_4585 = _zz_20946;
  assign _zz_4586 = _zz_20954;
  assign _zz_1958 = ($signed(_zz_20962) * $signed(data_mid_71_real));
  assign _zz_4587 = _zz_20963;
  assign _zz_1956 = _zz_20966[31 : 0];
  assign _zz_4588 = _zz_20967;
  assign _zz_1957 = _zz_20970[31 : 0];
  assign _zz_1959 = 1'b1;
  assign _zz_4589 = _zz_20971;
  assign _zz_4590 = _zz_20979;
  assign _zz_1960 = 1'b1;
  assign _zz_4591 = _zz_20987;
  assign _zz_4592 = _zz_20995;
  assign _zz_1963 = ($signed(_zz_21003) * $signed(data_mid_72_real));
  assign _zz_4593 = _zz_21004;
  assign _zz_1961 = _zz_21007[31 : 0];
  assign _zz_4594 = _zz_21008;
  assign _zz_1962 = _zz_21011[31 : 0];
  assign _zz_1964 = 1'b1;
  assign _zz_4595 = _zz_21012;
  assign _zz_4596 = _zz_21020;
  assign _zz_1965 = 1'b1;
  assign _zz_4597 = _zz_21028;
  assign _zz_4598 = _zz_21036;
  assign _zz_1968 = ($signed(_zz_21044) * $signed(data_mid_73_real));
  assign _zz_4599 = _zz_21045;
  assign _zz_1966 = _zz_21048[31 : 0];
  assign _zz_4600 = _zz_21049;
  assign _zz_1967 = _zz_21052[31 : 0];
  assign _zz_1969 = 1'b1;
  assign _zz_4601 = _zz_21053;
  assign _zz_4602 = _zz_21061;
  assign _zz_1970 = 1'b1;
  assign _zz_4603 = _zz_21069;
  assign _zz_4604 = _zz_21077;
  assign _zz_1973 = ($signed(_zz_21085) * $signed(data_mid_74_real));
  assign _zz_4605 = _zz_21086;
  assign _zz_1971 = _zz_21089[31 : 0];
  assign _zz_4606 = _zz_21090;
  assign _zz_1972 = _zz_21093[31 : 0];
  assign _zz_1974 = 1'b1;
  assign _zz_4607 = _zz_21094;
  assign _zz_4608 = _zz_21102;
  assign _zz_1975 = 1'b1;
  assign _zz_4609 = _zz_21110;
  assign _zz_4610 = _zz_21118;
  assign _zz_1978 = ($signed(_zz_21126) * $signed(data_mid_75_real));
  assign _zz_4611 = _zz_21127;
  assign _zz_1976 = _zz_21130[31 : 0];
  assign _zz_4612 = _zz_21131;
  assign _zz_1977 = _zz_21134[31 : 0];
  assign _zz_1979 = 1'b1;
  assign _zz_4613 = _zz_21135;
  assign _zz_4614 = _zz_21143;
  assign _zz_1980 = 1'b1;
  assign _zz_4615 = _zz_21151;
  assign _zz_4616 = _zz_21159;
  assign _zz_1983 = ($signed(_zz_21167) * $signed(data_mid_76_real));
  assign _zz_4617 = _zz_21168;
  assign _zz_1981 = _zz_21171[31 : 0];
  assign _zz_4618 = _zz_21172;
  assign _zz_1982 = _zz_21175[31 : 0];
  assign _zz_1984 = 1'b1;
  assign _zz_4619 = _zz_21176;
  assign _zz_4620 = _zz_21184;
  assign _zz_1985 = 1'b1;
  assign _zz_4621 = _zz_21192;
  assign _zz_4622 = _zz_21200;
  assign _zz_1988 = ($signed(_zz_21208) * $signed(data_mid_77_real));
  assign _zz_4623 = _zz_21209;
  assign _zz_1986 = _zz_21212[31 : 0];
  assign _zz_4624 = _zz_21213;
  assign _zz_1987 = _zz_21216[31 : 0];
  assign _zz_1989 = 1'b1;
  assign _zz_4625 = _zz_21217;
  assign _zz_4626 = _zz_21225;
  assign _zz_1990 = 1'b1;
  assign _zz_4627 = _zz_21233;
  assign _zz_4628 = _zz_21241;
  assign _zz_1993 = ($signed(_zz_21249) * $signed(data_mid_78_real));
  assign _zz_4629 = _zz_21250;
  assign _zz_1991 = _zz_21253[31 : 0];
  assign _zz_4630 = _zz_21254;
  assign _zz_1992 = _zz_21257[31 : 0];
  assign _zz_1994 = 1'b1;
  assign _zz_4631 = _zz_21258;
  assign _zz_4632 = _zz_21266;
  assign _zz_1995 = 1'b1;
  assign _zz_4633 = _zz_21274;
  assign _zz_4634 = _zz_21282;
  assign _zz_1998 = ($signed(_zz_21290) * $signed(data_mid_79_real));
  assign _zz_4635 = _zz_21291;
  assign _zz_1996 = _zz_21294[31 : 0];
  assign _zz_4636 = _zz_21295;
  assign _zz_1997 = _zz_21298[31 : 0];
  assign _zz_1999 = 1'b1;
  assign _zz_4637 = _zz_21299;
  assign _zz_4638 = _zz_21307;
  assign _zz_2000 = 1'b1;
  assign _zz_4639 = _zz_21315;
  assign _zz_4640 = _zz_21323;
  assign _zz_2003 = ($signed(_zz_21331) * $signed(data_mid_80_real));
  assign _zz_4641 = _zz_21332;
  assign _zz_2001 = _zz_21335[31 : 0];
  assign _zz_4642 = _zz_21336;
  assign _zz_2002 = _zz_21339[31 : 0];
  assign _zz_2004 = 1'b1;
  assign _zz_4643 = _zz_21340;
  assign _zz_4644 = _zz_21348;
  assign _zz_2005 = 1'b1;
  assign _zz_4645 = _zz_21356;
  assign _zz_4646 = _zz_21364;
  assign _zz_2008 = ($signed(_zz_21372) * $signed(data_mid_81_real));
  assign _zz_4647 = _zz_21373;
  assign _zz_2006 = _zz_21376[31 : 0];
  assign _zz_4648 = _zz_21377;
  assign _zz_2007 = _zz_21380[31 : 0];
  assign _zz_2009 = 1'b1;
  assign _zz_4649 = _zz_21381;
  assign _zz_4650 = _zz_21389;
  assign _zz_2010 = 1'b1;
  assign _zz_4651 = _zz_21397;
  assign _zz_4652 = _zz_21405;
  assign _zz_2013 = ($signed(_zz_21413) * $signed(data_mid_82_real));
  assign _zz_4653 = _zz_21414;
  assign _zz_2011 = _zz_21417[31 : 0];
  assign _zz_4654 = _zz_21418;
  assign _zz_2012 = _zz_21421[31 : 0];
  assign _zz_2014 = 1'b1;
  assign _zz_4655 = _zz_21422;
  assign _zz_4656 = _zz_21430;
  assign _zz_2015 = 1'b1;
  assign _zz_4657 = _zz_21438;
  assign _zz_4658 = _zz_21446;
  assign _zz_2018 = ($signed(_zz_21454) * $signed(data_mid_83_real));
  assign _zz_4659 = _zz_21455;
  assign _zz_2016 = _zz_21458[31 : 0];
  assign _zz_4660 = _zz_21459;
  assign _zz_2017 = _zz_21462[31 : 0];
  assign _zz_2019 = 1'b1;
  assign _zz_4661 = _zz_21463;
  assign _zz_4662 = _zz_21471;
  assign _zz_2020 = 1'b1;
  assign _zz_4663 = _zz_21479;
  assign _zz_4664 = _zz_21487;
  assign _zz_2023 = ($signed(_zz_21495) * $signed(data_mid_84_real));
  assign _zz_4665 = _zz_21496;
  assign _zz_2021 = _zz_21499[31 : 0];
  assign _zz_4666 = _zz_21500;
  assign _zz_2022 = _zz_21503[31 : 0];
  assign _zz_2024 = 1'b1;
  assign _zz_4667 = _zz_21504;
  assign _zz_4668 = _zz_21512;
  assign _zz_2025 = 1'b1;
  assign _zz_4669 = _zz_21520;
  assign _zz_4670 = _zz_21528;
  assign _zz_2028 = ($signed(_zz_21536) * $signed(data_mid_85_real));
  assign _zz_4671 = _zz_21537;
  assign _zz_2026 = _zz_21540[31 : 0];
  assign _zz_4672 = _zz_21541;
  assign _zz_2027 = _zz_21544[31 : 0];
  assign _zz_2029 = 1'b1;
  assign _zz_4673 = _zz_21545;
  assign _zz_4674 = _zz_21553;
  assign _zz_2030 = 1'b1;
  assign _zz_4675 = _zz_21561;
  assign _zz_4676 = _zz_21569;
  assign _zz_2033 = ($signed(_zz_21577) * $signed(data_mid_86_real));
  assign _zz_4677 = _zz_21578;
  assign _zz_2031 = _zz_21581[31 : 0];
  assign _zz_4678 = _zz_21582;
  assign _zz_2032 = _zz_21585[31 : 0];
  assign _zz_2034 = 1'b1;
  assign _zz_4679 = _zz_21586;
  assign _zz_4680 = _zz_21594;
  assign _zz_2035 = 1'b1;
  assign _zz_4681 = _zz_21602;
  assign _zz_4682 = _zz_21610;
  assign _zz_2038 = ($signed(_zz_21618) * $signed(data_mid_87_real));
  assign _zz_4683 = _zz_21619;
  assign _zz_2036 = _zz_21622[31 : 0];
  assign _zz_4684 = _zz_21623;
  assign _zz_2037 = _zz_21626[31 : 0];
  assign _zz_2039 = 1'b1;
  assign _zz_4685 = _zz_21627;
  assign _zz_4686 = _zz_21635;
  assign _zz_2040 = 1'b1;
  assign _zz_4687 = _zz_21643;
  assign _zz_4688 = _zz_21651;
  assign _zz_2043 = ($signed(_zz_21659) * $signed(data_mid_88_real));
  assign _zz_4689 = _zz_21660;
  assign _zz_2041 = _zz_21663[31 : 0];
  assign _zz_4690 = _zz_21664;
  assign _zz_2042 = _zz_21667[31 : 0];
  assign _zz_2044 = 1'b1;
  assign _zz_4691 = _zz_21668;
  assign _zz_4692 = _zz_21676;
  assign _zz_2045 = 1'b1;
  assign _zz_4693 = _zz_21684;
  assign _zz_4694 = _zz_21692;
  assign _zz_2048 = ($signed(_zz_21700) * $signed(data_mid_89_real));
  assign _zz_4695 = _zz_21701;
  assign _zz_2046 = _zz_21704[31 : 0];
  assign _zz_4696 = _zz_21705;
  assign _zz_2047 = _zz_21708[31 : 0];
  assign _zz_2049 = 1'b1;
  assign _zz_4697 = _zz_21709;
  assign _zz_4698 = _zz_21717;
  assign _zz_2050 = 1'b1;
  assign _zz_4699 = _zz_21725;
  assign _zz_4700 = _zz_21733;
  assign _zz_2053 = ($signed(_zz_21741) * $signed(data_mid_90_real));
  assign _zz_4701 = _zz_21742;
  assign _zz_2051 = _zz_21745[31 : 0];
  assign _zz_4702 = _zz_21746;
  assign _zz_2052 = _zz_21749[31 : 0];
  assign _zz_2054 = 1'b1;
  assign _zz_4703 = _zz_21750;
  assign _zz_4704 = _zz_21758;
  assign _zz_2055 = 1'b1;
  assign _zz_4705 = _zz_21766;
  assign _zz_4706 = _zz_21774;
  assign _zz_2058 = ($signed(_zz_21782) * $signed(data_mid_91_real));
  assign _zz_4707 = _zz_21783;
  assign _zz_2056 = _zz_21786[31 : 0];
  assign _zz_4708 = _zz_21787;
  assign _zz_2057 = _zz_21790[31 : 0];
  assign _zz_2059 = 1'b1;
  assign _zz_4709 = _zz_21791;
  assign _zz_4710 = _zz_21799;
  assign _zz_2060 = 1'b1;
  assign _zz_4711 = _zz_21807;
  assign _zz_4712 = _zz_21815;
  assign _zz_2063 = ($signed(_zz_21823) * $signed(data_mid_92_real));
  assign _zz_4713 = _zz_21824;
  assign _zz_2061 = _zz_21827[31 : 0];
  assign _zz_4714 = _zz_21828;
  assign _zz_2062 = _zz_21831[31 : 0];
  assign _zz_2064 = 1'b1;
  assign _zz_4715 = _zz_21832;
  assign _zz_4716 = _zz_21840;
  assign _zz_2065 = 1'b1;
  assign _zz_4717 = _zz_21848;
  assign _zz_4718 = _zz_21856;
  assign _zz_2068 = ($signed(_zz_21864) * $signed(data_mid_93_real));
  assign _zz_4719 = _zz_21865;
  assign _zz_2066 = _zz_21868[31 : 0];
  assign _zz_4720 = _zz_21869;
  assign _zz_2067 = _zz_21872[31 : 0];
  assign _zz_2069 = 1'b1;
  assign _zz_4721 = _zz_21873;
  assign _zz_4722 = _zz_21881;
  assign _zz_2070 = 1'b1;
  assign _zz_4723 = _zz_21889;
  assign _zz_4724 = _zz_21897;
  assign _zz_2073 = ($signed(_zz_21905) * $signed(data_mid_94_real));
  assign _zz_4725 = _zz_21906;
  assign _zz_2071 = _zz_21909[31 : 0];
  assign _zz_4726 = _zz_21910;
  assign _zz_2072 = _zz_21913[31 : 0];
  assign _zz_2074 = 1'b1;
  assign _zz_4727 = _zz_21914;
  assign _zz_4728 = _zz_21922;
  assign _zz_2075 = 1'b1;
  assign _zz_4729 = _zz_21930;
  assign _zz_4730 = _zz_21938;
  assign _zz_2078 = ($signed(_zz_21946) * $signed(data_mid_95_real));
  assign _zz_4731 = _zz_21947;
  assign _zz_2076 = _zz_21950[31 : 0];
  assign _zz_4732 = _zz_21951;
  assign _zz_2077 = _zz_21954[31 : 0];
  assign _zz_2079 = 1'b1;
  assign _zz_4733 = _zz_21955;
  assign _zz_4734 = _zz_21963;
  assign _zz_2080 = 1'b1;
  assign _zz_4735 = _zz_21971;
  assign _zz_4736 = _zz_21979;
  assign _zz_2083 = ($signed(_zz_21987) * $signed(data_mid_96_real));
  assign _zz_4737 = _zz_21988;
  assign _zz_2081 = _zz_21991[31 : 0];
  assign _zz_4738 = _zz_21992;
  assign _zz_2082 = _zz_21995[31 : 0];
  assign _zz_2084 = 1'b1;
  assign _zz_4739 = _zz_21996;
  assign _zz_4740 = _zz_22004;
  assign _zz_2085 = 1'b1;
  assign _zz_4741 = _zz_22012;
  assign _zz_4742 = _zz_22020;
  assign _zz_2088 = ($signed(_zz_22028) * $signed(data_mid_97_real));
  assign _zz_4743 = _zz_22029;
  assign _zz_2086 = _zz_22032[31 : 0];
  assign _zz_4744 = _zz_22033;
  assign _zz_2087 = _zz_22036[31 : 0];
  assign _zz_2089 = 1'b1;
  assign _zz_4745 = _zz_22037;
  assign _zz_4746 = _zz_22045;
  assign _zz_2090 = 1'b1;
  assign _zz_4747 = _zz_22053;
  assign _zz_4748 = _zz_22061;
  assign _zz_2093 = ($signed(_zz_22069) * $signed(data_mid_98_real));
  assign _zz_4749 = _zz_22070;
  assign _zz_2091 = _zz_22073[31 : 0];
  assign _zz_4750 = _zz_22074;
  assign _zz_2092 = _zz_22077[31 : 0];
  assign _zz_2094 = 1'b1;
  assign _zz_4751 = _zz_22078;
  assign _zz_4752 = _zz_22086;
  assign _zz_2095 = 1'b1;
  assign _zz_4753 = _zz_22094;
  assign _zz_4754 = _zz_22102;
  assign _zz_2098 = ($signed(_zz_22110) * $signed(data_mid_99_real));
  assign _zz_4755 = _zz_22111;
  assign _zz_2096 = _zz_22114[31 : 0];
  assign _zz_4756 = _zz_22115;
  assign _zz_2097 = _zz_22118[31 : 0];
  assign _zz_2099 = 1'b1;
  assign _zz_4757 = _zz_22119;
  assign _zz_4758 = _zz_22127;
  assign _zz_2100 = 1'b1;
  assign _zz_4759 = _zz_22135;
  assign _zz_4760 = _zz_22143;
  assign _zz_2103 = ($signed(_zz_22151) * $signed(data_mid_100_real));
  assign _zz_4761 = _zz_22152;
  assign _zz_2101 = _zz_22155[31 : 0];
  assign _zz_4762 = _zz_22156;
  assign _zz_2102 = _zz_22159[31 : 0];
  assign _zz_2104 = 1'b1;
  assign _zz_4763 = _zz_22160;
  assign _zz_4764 = _zz_22168;
  assign _zz_2105 = 1'b1;
  assign _zz_4765 = _zz_22176;
  assign _zz_4766 = _zz_22184;
  assign _zz_2108 = ($signed(_zz_22192) * $signed(data_mid_101_real));
  assign _zz_4767 = _zz_22193;
  assign _zz_2106 = _zz_22196[31 : 0];
  assign _zz_4768 = _zz_22197;
  assign _zz_2107 = _zz_22200[31 : 0];
  assign _zz_2109 = 1'b1;
  assign _zz_4769 = _zz_22201;
  assign _zz_4770 = _zz_22209;
  assign _zz_2110 = 1'b1;
  assign _zz_4771 = _zz_22217;
  assign _zz_4772 = _zz_22225;
  assign _zz_2113 = ($signed(_zz_22233) * $signed(data_mid_102_real));
  assign _zz_4773 = _zz_22234;
  assign _zz_2111 = _zz_22237[31 : 0];
  assign _zz_4774 = _zz_22238;
  assign _zz_2112 = _zz_22241[31 : 0];
  assign _zz_2114 = 1'b1;
  assign _zz_4775 = _zz_22242;
  assign _zz_4776 = _zz_22250;
  assign _zz_2115 = 1'b1;
  assign _zz_4777 = _zz_22258;
  assign _zz_4778 = _zz_22266;
  assign _zz_2118 = ($signed(_zz_22274) * $signed(data_mid_103_real));
  assign _zz_4779 = _zz_22275;
  assign _zz_2116 = _zz_22278[31 : 0];
  assign _zz_4780 = _zz_22279;
  assign _zz_2117 = _zz_22282[31 : 0];
  assign _zz_2119 = 1'b1;
  assign _zz_4781 = _zz_22283;
  assign _zz_4782 = _zz_22291;
  assign _zz_2120 = 1'b1;
  assign _zz_4783 = _zz_22299;
  assign _zz_4784 = _zz_22307;
  assign _zz_2123 = ($signed(_zz_22315) * $signed(data_mid_104_real));
  assign _zz_4785 = _zz_22316;
  assign _zz_2121 = _zz_22319[31 : 0];
  assign _zz_4786 = _zz_22320;
  assign _zz_2122 = _zz_22323[31 : 0];
  assign _zz_2124 = 1'b1;
  assign _zz_4787 = _zz_22324;
  assign _zz_4788 = _zz_22332;
  assign _zz_2125 = 1'b1;
  assign _zz_4789 = _zz_22340;
  assign _zz_4790 = _zz_22348;
  assign _zz_2128 = ($signed(_zz_22356) * $signed(data_mid_105_real));
  assign _zz_4791 = _zz_22357;
  assign _zz_2126 = _zz_22360[31 : 0];
  assign _zz_4792 = _zz_22361;
  assign _zz_2127 = _zz_22364[31 : 0];
  assign _zz_2129 = 1'b1;
  assign _zz_4793 = _zz_22365;
  assign _zz_4794 = _zz_22373;
  assign _zz_2130 = 1'b1;
  assign _zz_4795 = _zz_22381;
  assign _zz_4796 = _zz_22389;
  assign _zz_2133 = ($signed(_zz_22397) * $signed(data_mid_106_real));
  assign _zz_4797 = _zz_22398;
  assign _zz_2131 = _zz_22401[31 : 0];
  assign _zz_4798 = _zz_22402;
  assign _zz_2132 = _zz_22405[31 : 0];
  assign _zz_2134 = 1'b1;
  assign _zz_4799 = _zz_22406;
  assign _zz_4800 = _zz_22414;
  assign _zz_2135 = 1'b1;
  assign _zz_4801 = _zz_22422;
  assign _zz_4802 = _zz_22430;
  assign _zz_2138 = ($signed(_zz_22438) * $signed(data_mid_107_real));
  assign _zz_4803 = _zz_22439;
  assign _zz_2136 = _zz_22442[31 : 0];
  assign _zz_4804 = _zz_22443;
  assign _zz_2137 = _zz_22446[31 : 0];
  assign _zz_2139 = 1'b1;
  assign _zz_4805 = _zz_22447;
  assign _zz_4806 = _zz_22455;
  assign _zz_2140 = 1'b1;
  assign _zz_4807 = _zz_22463;
  assign _zz_4808 = _zz_22471;
  assign _zz_2143 = ($signed(_zz_22479) * $signed(data_mid_108_real));
  assign _zz_4809 = _zz_22480;
  assign _zz_2141 = _zz_22483[31 : 0];
  assign _zz_4810 = _zz_22484;
  assign _zz_2142 = _zz_22487[31 : 0];
  assign _zz_2144 = 1'b1;
  assign _zz_4811 = _zz_22488;
  assign _zz_4812 = _zz_22496;
  assign _zz_2145 = 1'b1;
  assign _zz_4813 = _zz_22504;
  assign _zz_4814 = _zz_22512;
  assign _zz_2148 = ($signed(_zz_22520) * $signed(data_mid_109_real));
  assign _zz_4815 = _zz_22521;
  assign _zz_2146 = _zz_22524[31 : 0];
  assign _zz_4816 = _zz_22525;
  assign _zz_2147 = _zz_22528[31 : 0];
  assign _zz_2149 = 1'b1;
  assign _zz_4817 = _zz_22529;
  assign _zz_4818 = _zz_22537;
  assign _zz_2150 = 1'b1;
  assign _zz_4819 = _zz_22545;
  assign _zz_4820 = _zz_22553;
  assign _zz_2153 = ($signed(_zz_22561) * $signed(data_mid_110_real));
  assign _zz_4821 = _zz_22562;
  assign _zz_2151 = _zz_22565[31 : 0];
  assign _zz_4822 = _zz_22566;
  assign _zz_2152 = _zz_22569[31 : 0];
  assign _zz_2154 = 1'b1;
  assign _zz_4823 = _zz_22570;
  assign _zz_4824 = _zz_22578;
  assign _zz_2155 = 1'b1;
  assign _zz_4825 = _zz_22586;
  assign _zz_4826 = _zz_22594;
  assign _zz_2158 = ($signed(_zz_22602) * $signed(data_mid_111_real));
  assign _zz_4827 = _zz_22603;
  assign _zz_2156 = _zz_22606[31 : 0];
  assign _zz_4828 = _zz_22607;
  assign _zz_2157 = _zz_22610[31 : 0];
  assign _zz_2159 = 1'b1;
  assign _zz_4829 = _zz_22611;
  assign _zz_4830 = _zz_22619;
  assign _zz_2160 = 1'b1;
  assign _zz_4831 = _zz_22627;
  assign _zz_4832 = _zz_22635;
  assign _zz_2163 = ($signed(_zz_22643) * $signed(data_mid_112_real));
  assign _zz_4833 = _zz_22644;
  assign _zz_2161 = _zz_22647[31 : 0];
  assign _zz_4834 = _zz_22648;
  assign _zz_2162 = _zz_22651[31 : 0];
  assign _zz_2164 = 1'b1;
  assign _zz_4835 = _zz_22652;
  assign _zz_4836 = _zz_22660;
  assign _zz_2165 = 1'b1;
  assign _zz_4837 = _zz_22668;
  assign _zz_4838 = _zz_22676;
  assign _zz_2168 = ($signed(_zz_22684) * $signed(data_mid_113_real));
  assign _zz_4839 = _zz_22685;
  assign _zz_2166 = _zz_22688[31 : 0];
  assign _zz_4840 = _zz_22689;
  assign _zz_2167 = _zz_22692[31 : 0];
  assign _zz_2169 = 1'b1;
  assign _zz_4841 = _zz_22693;
  assign _zz_4842 = _zz_22701;
  assign _zz_2170 = 1'b1;
  assign _zz_4843 = _zz_22709;
  assign _zz_4844 = _zz_22717;
  assign _zz_2173 = ($signed(_zz_22725) * $signed(data_mid_114_real));
  assign _zz_4845 = _zz_22726;
  assign _zz_2171 = _zz_22729[31 : 0];
  assign _zz_4846 = _zz_22730;
  assign _zz_2172 = _zz_22733[31 : 0];
  assign _zz_2174 = 1'b1;
  assign _zz_4847 = _zz_22734;
  assign _zz_4848 = _zz_22742;
  assign _zz_2175 = 1'b1;
  assign _zz_4849 = _zz_22750;
  assign _zz_4850 = _zz_22758;
  assign _zz_2178 = ($signed(_zz_22766) * $signed(data_mid_115_real));
  assign _zz_4851 = _zz_22767;
  assign _zz_2176 = _zz_22770[31 : 0];
  assign _zz_4852 = _zz_22771;
  assign _zz_2177 = _zz_22774[31 : 0];
  assign _zz_2179 = 1'b1;
  assign _zz_4853 = _zz_22775;
  assign _zz_4854 = _zz_22783;
  assign _zz_2180 = 1'b1;
  assign _zz_4855 = _zz_22791;
  assign _zz_4856 = _zz_22799;
  assign _zz_2183 = ($signed(_zz_22807) * $signed(data_mid_116_real));
  assign _zz_4857 = _zz_22808;
  assign _zz_2181 = _zz_22811[31 : 0];
  assign _zz_4858 = _zz_22812;
  assign _zz_2182 = _zz_22815[31 : 0];
  assign _zz_2184 = 1'b1;
  assign _zz_4859 = _zz_22816;
  assign _zz_4860 = _zz_22824;
  assign _zz_2185 = 1'b1;
  assign _zz_4861 = _zz_22832;
  assign _zz_4862 = _zz_22840;
  assign _zz_2188 = ($signed(_zz_22848) * $signed(data_mid_117_real));
  assign _zz_4863 = _zz_22849;
  assign _zz_2186 = _zz_22852[31 : 0];
  assign _zz_4864 = _zz_22853;
  assign _zz_2187 = _zz_22856[31 : 0];
  assign _zz_2189 = 1'b1;
  assign _zz_4865 = _zz_22857;
  assign _zz_4866 = _zz_22865;
  assign _zz_2190 = 1'b1;
  assign _zz_4867 = _zz_22873;
  assign _zz_4868 = _zz_22881;
  assign _zz_2193 = ($signed(_zz_22889) * $signed(data_mid_118_real));
  assign _zz_4869 = _zz_22890;
  assign _zz_2191 = _zz_22893[31 : 0];
  assign _zz_4870 = _zz_22894;
  assign _zz_2192 = _zz_22897[31 : 0];
  assign _zz_2194 = 1'b1;
  assign _zz_4871 = _zz_22898;
  assign _zz_4872 = _zz_22906;
  assign _zz_2195 = 1'b1;
  assign _zz_4873 = _zz_22914;
  assign _zz_4874 = _zz_22922;
  assign _zz_2198 = ($signed(_zz_22930) * $signed(data_mid_119_real));
  assign _zz_4875 = _zz_22931;
  assign _zz_2196 = _zz_22934[31 : 0];
  assign _zz_4876 = _zz_22935;
  assign _zz_2197 = _zz_22938[31 : 0];
  assign _zz_2199 = 1'b1;
  assign _zz_4877 = _zz_22939;
  assign _zz_4878 = _zz_22947;
  assign _zz_2200 = 1'b1;
  assign _zz_4879 = _zz_22955;
  assign _zz_4880 = _zz_22963;
  assign _zz_2203 = ($signed(_zz_22971) * $signed(data_mid_120_real));
  assign _zz_4881 = _zz_22972;
  assign _zz_2201 = _zz_22975[31 : 0];
  assign _zz_4882 = _zz_22976;
  assign _zz_2202 = _zz_22979[31 : 0];
  assign _zz_2204 = 1'b1;
  assign _zz_4883 = _zz_22980;
  assign _zz_4884 = _zz_22988;
  assign _zz_2205 = 1'b1;
  assign _zz_4885 = _zz_22996;
  assign _zz_4886 = _zz_23004;
  assign _zz_2208 = ($signed(_zz_23012) * $signed(data_mid_121_real));
  assign _zz_4887 = _zz_23013;
  assign _zz_2206 = _zz_23016[31 : 0];
  assign _zz_4888 = _zz_23017;
  assign _zz_2207 = _zz_23020[31 : 0];
  assign _zz_2209 = 1'b1;
  assign _zz_4889 = _zz_23021;
  assign _zz_4890 = _zz_23029;
  assign _zz_2210 = 1'b1;
  assign _zz_4891 = _zz_23037;
  assign _zz_4892 = _zz_23045;
  assign _zz_2213 = ($signed(_zz_23053) * $signed(data_mid_122_real));
  assign _zz_4893 = _zz_23054;
  assign _zz_2211 = _zz_23057[31 : 0];
  assign _zz_4894 = _zz_23058;
  assign _zz_2212 = _zz_23061[31 : 0];
  assign _zz_2214 = 1'b1;
  assign _zz_4895 = _zz_23062;
  assign _zz_4896 = _zz_23070;
  assign _zz_2215 = 1'b1;
  assign _zz_4897 = _zz_23078;
  assign _zz_4898 = _zz_23086;
  assign _zz_2218 = ($signed(_zz_23094) * $signed(data_mid_123_real));
  assign _zz_4899 = _zz_23095;
  assign _zz_2216 = _zz_23098[31 : 0];
  assign _zz_4900 = _zz_23099;
  assign _zz_2217 = _zz_23102[31 : 0];
  assign _zz_2219 = 1'b1;
  assign _zz_4901 = _zz_23103;
  assign _zz_4902 = _zz_23111;
  assign _zz_2220 = 1'b1;
  assign _zz_4903 = _zz_23119;
  assign _zz_4904 = _zz_23127;
  assign _zz_2223 = ($signed(_zz_23135) * $signed(data_mid_124_real));
  assign _zz_4905 = _zz_23136;
  assign _zz_2221 = _zz_23139[31 : 0];
  assign _zz_4906 = _zz_23140;
  assign _zz_2222 = _zz_23143[31 : 0];
  assign _zz_2224 = 1'b1;
  assign _zz_4907 = _zz_23144;
  assign _zz_4908 = _zz_23152;
  assign _zz_2225 = 1'b1;
  assign _zz_4909 = _zz_23160;
  assign _zz_4910 = _zz_23168;
  assign _zz_2228 = ($signed(_zz_23176) * $signed(data_mid_125_real));
  assign _zz_4911 = _zz_23177;
  assign _zz_2226 = _zz_23180[31 : 0];
  assign _zz_4912 = _zz_23181;
  assign _zz_2227 = _zz_23184[31 : 0];
  assign _zz_2229 = 1'b1;
  assign _zz_4913 = _zz_23185;
  assign _zz_4914 = _zz_23193;
  assign _zz_2230 = 1'b1;
  assign _zz_4915 = _zz_23201;
  assign _zz_4916 = _zz_23209;
  assign _zz_2233 = ($signed(_zz_23217) * $signed(data_mid_126_real));
  assign _zz_4917 = _zz_23218;
  assign _zz_2231 = _zz_23221[31 : 0];
  assign _zz_4918 = _zz_23222;
  assign _zz_2232 = _zz_23225[31 : 0];
  assign _zz_2234 = 1'b1;
  assign _zz_4919 = _zz_23226;
  assign _zz_4920 = _zz_23234;
  assign _zz_2235 = 1'b1;
  assign _zz_4921 = _zz_23242;
  assign _zz_4922 = _zz_23250;
  assign _zz_2238 = ($signed(_zz_23258) * $signed(data_mid_127_real));
  assign _zz_4923 = _zz_23259;
  assign _zz_2236 = _zz_23262[31 : 0];
  assign _zz_4924 = _zz_23263;
  assign _zz_2237 = _zz_23266[31 : 0];
  assign _zz_2239 = 1'b1;
  assign _zz_4925 = _zz_23267;
  assign _zz_4926 = _zz_23275;
  assign _zz_2240 = 1'b1;
  assign _zz_4927 = _zz_23283;
  assign _zz_4928 = _zz_23291;
  assign sdata_out_valid = current_level_willOverflow_regNext;
  assign sdata_out_payload_0_real = data_mid_0_real;
  assign sdata_out_payload_0_imag = data_mid_0_imag;
  assign sdata_out_payload_1_real = data_mid_1_real;
  assign sdata_out_payload_1_imag = data_mid_1_imag;
  assign sdata_out_payload_2_real = data_mid_2_real;
  assign sdata_out_payload_2_imag = data_mid_2_imag;
  assign sdata_out_payload_3_real = data_mid_3_real;
  assign sdata_out_payload_3_imag = data_mid_3_imag;
  assign sdata_out_payload_4_real = data_mid_4_real;
  assign sdata_out_payload_4_imag = data_mid_4_imag;
  assign sdata_out_payload_5_real = data_mid_5_real;
  assign sdata_out_payload_5_imag = data_mid_5_imag;
  assign sdata_out_payload_6_real = data_mid_6_real;
  assign sdata_out_payload_6_imag = data_mid_6_imag;
  assign sdata_out_payload_7_real = data_mid_7_real;
  assign sdata_out_payload_7_imag = data_mid_7_imag;
  assign sdata_out_payload_8_real = data_mid_8_real;
  assign sdata_out_payload_8_imag = data_mid_8_imag;
  assign sdata_out_payload_9_real = data_mid_9_real;
  assign sdata_out_payload_9_imag = data_mid_9_imag;
  assign sdata_out_payload_10_real = data_mid_10_real;
  assign sdata_out_payload_10_imag = data_mid_10_imag;
  assign sdata_out_payload_11_real = data_mid_11_real;
  assign sdata_out_payload_11_imag = data_mid_11_imag;
  assign sdata_out_payload_12_real = data_mid_12_real;
  assign sdata_out_payload_12_imag = data_mid_12_imag;
  assign sdata_out_payload_13_real = data_mid_13_real;
  assign sdata_out_payload_13_imag = data_mid_13_imag;
  assign sdata_out_payload_14_real = data_mid_14_real;
  assign sdata_out_payload_14_imag = data_mid_14_imag;
  assign sdata_out_payload_15_real = data_mid_15_real;
  assign sdata_out_payload_15_imag = data_mid_15_imag;
  assign sdata_out_payload_16_real = data_mid_16_real;
  assign sdata_out_payload_16_imag = data_mid_16_imag;
  assign sdata_out_payload_17_real = data_mid_17_real;
  assign sdata_out_payload_17_imag = data_mid_17_imag;
  assign sdata_out_payload_18_real = data_mid_18_real;
  assign sdata_out_payload_18_imag = data_mid_18_imag;
  assign sdata_out_payload_19_real = data_mid_19_real;
  assign sdata_out_payload_19_imag = data_mid_19_imag;
  assign sdata_out_payload_20_real = data_mid_20_real;
  assign sdata_out_payload_20_imag = data_mid_20_imag;
  assign sdata_out_payload_21_real = data_mid_21_real;
  assign sdata_out_payload_21_imag = data_mid_21_imag;
  assign sdata_out_payload_22_real = data_mid_22_real;
  assign sdata_out_payload_22_imag = data_mid_22_imag;
  assign sdata_out_payload_23_real = data_mid_23_real;
  assign sdata_out_payload_23_imag = data_mid_23_imag;
  assign sdata_out_payload_24_real = data_mid_24_real;
  assign sdata_out_payload_24_imag = data_mid_24_imag;
  assign sdata_out_payload_25_real = data_mid_25_real;
  assign sdata_out_payload_25_imag = data_mid_25_imag;
  assign sdata_out_payload_26_real = data_mid_26_real;
  assign sdata_out_payload_26_imag = data_mid_26_imag;
  assign sdata_out_payload_27_real = data_mid_27_real;
  assign sdata_out_payload_27_imag = data_mid_27_imag;
  assign sdata_out_payload_28_real = data_mid_28_real;
  assign sdata_out_payload_28_imag = data_mid_28_imag;
  assign sdata_out_payload_29_real = data_mid_29_real;
  assign sdata_out_payload_29_imag = data_mid_29_imag;
  assign sdata_out_payload_30_real = data_mid_30_real;
  assign sdata_out_payload_30_imag = data_mid_30_imag;
  assign sdata_out_payload_31_real = data_mid_31_real;
  assign sdata_out_payload_31_imag = data_mid_31_imag;
  assign sdata_out_payload_32_real = data_mid_32_real;
  assign sdata_out_payload_32_imag = data_mid_32_imag;
  assign sdata_out_payload_33_real = data_mid_33_real;
  assign sdata_out_payload_33_imag = data_mid_33_imag;
  assign sdata_out_payload_34_real = data_mid_34_real;
  assign sdata_out_payload_34_imag = data_mid_34_imag;
  assign sdata_out_payload_35_real = data_mid_35_real;
  assign sdata_out_payload_35_imag = data_mid_35_imag;
  assign sdata_out_payload_36_real = data_mid_36_real;
  assign sdata_out_payload_36_imag = data_mid_36_imag;
  assign sdata_out_payload_37_real = data_mid_37_real;
  assign sdata_out_payload_37_imag = data_mid_37_imag;
  assign sdata_out_payload_38_real = data_mid_38_real;
  assign sdata_out_payload_38_imag = data_mid_38_imag;
  assign sdata_out_payload_39_real = data_mid_39_real;
  assign sdata_out_payload_39_imag = data_mid_39_imag;
  assign sdata_out_payload_40_real = data_mid_40_real;
  assign sdata_out_payload_40_imag = data_mid_40_imag;
  assign sdata_out_payload_41_real = data_mid_41_real;
  assign sdata_out_payload_41_imag = data_mid_41_imag;
  assign sdata_out_payload_42_real = data_mid_42_real;
  assign sdata_out_payload_42_imag = data_mid_42_imag;
  assign sdata_out_payload_43_real = data_mid_43_real;
  assign sdata_out_payload_43_imag = data_mid_43_imag;
  assign sdata_out_payload_44_real = data_mid_44_real;
  assign sdata_out_payload_44_imag = data_mid_44_imag;
  assign sdata_out_payload_45_real = data_mid_45_real;
  assign sdata_out_payload_45_imag = data_mid_45_imag;
  assign sdata_out_payload_46_real = data_mid_46_real;
  assign sdata_out_payload_46_imag = data_mid_46_imag;
  assign sdata_out_payload_47_real = data_mid_47_real;
  assign sdata_out_payload_47_imag = data_mid_47_imag;
  assign sdata_out_payload_48_real = data_mid_48_real;
  assign sdata_out_payload_48_imag = data_mid_48_imag;
  assign sdata_out_payload_49_real = data_mid_49_real;
  assign sdata_out_payload_49_imag = data_mid_49_imag;
  assign sdata_out_payload_50_real = data_mid_50_real;
  assign sdata_out_payload_50_imag = data_mid_50_imag;
  assign sdata_out_payload_51_real = data_mid_51_real;
  assign sdata_out_payload_51_imag = data_mid_51_imag;
  assign sdata_out_payload_52_real = data_mid_52_real;
  assign sdata_out_payload_52_imag = data_mid_52_imag;
  assign sdata_out_payload_53_real = data_mid_53_real;
  assign sdata_out_payload_53_imag = data_mid_53_imag;
  assign sdata_out_payload_54_real = data_mid_54_real;
  assign sdata_out_payload_54_imag = data_mid_54_imag;
  assign sdata_out_payload_55_real = data_mid_55_real;
  assign sdata_out_payload_55_imag = data_mid_55_imag;
  assign sdata_out_payload_56_real = data_mid_56_real;
  assign sdata_out_payload_56_imag = data_mid_56_imag;
  assign sdata_out_payload_57_real = data_mid_57_real;
  assign sdata_out_payload_57_imag = data_mid_57_imag;
  assign sdata_out_payload_58_real = data_mid_58_real;
  assign sdata_out_payload_58_imag = data_mid_58_imag;
  assign sdata_out_payload_59_real = data_mid_59_real;
  assign sdata_out_payload_59_imag = data_mid_59_imag;
  assign sdata_out_payload_60_real = data_mid_60_real;
  assign sdata_out_payload_60_imag = data_mid_60_imag;
  assign sdata_out_payload_61_real = data_mid_61_real;
  assign sdata_out_payload_61_imag = data_mid_61_imag;
  assign sdata_out_payload_62_real = data_mid_62_real;
  assign sdata_out_payload_62_imag = data_mid_62_imag;
  assign sdata_out_payload_63_real = data_mid_63_real;
  assign sdata_out_payload_63_imag = data_mid_63_imag;
  assign sdata_out_payload_64_real = data_mid_64_real;
  assign sdata_out_payload_64_imag = data_mid_64_imag;
  assign sdata_out_payload_65_real = data_mid_65_real;
  assign sdata_out_payload_65_imag = data_mid_65_imag;
  assign sdata_out_payload_66_real = data_mid_66_real;
  assign sdata_out_payload_66_imag = data_mid_66_imag;
  assign sdata_out_payload_67_real = data_mid_67_real;
  assign sdata_out_payload_67_imag = data_mid_67_imag;
  assign sdata_out_payload_68_real = data_mid_68_real;
  assign sdata_out_payload_68_imag = data_mid_68_imag;
  assign sdata_out_payload_69_real = data_mid_69_real;
  assign sdata_out_payload_69_imag = data_mid_69_imag;
  assign sdata_out_payload_70_real = data_mid_70_real;
  assign sdata_out_payload_70_imag = data_mid_70_imag;
  assign sdata_out_payload_71_real = data_mid_71_real;
  assign sdata_out_payload_71_imag = data_mid_71_imag;
  assign sdata_out_payload_72_real = data_mid_72_real;
  assign sdata_out_payload_72_imag = data_mid_72_imag;
  assign sdata_out_payload_73_real = data_mid_73_real;
  assign sdata_out_payload_73_imag = data_mid_73_imag;
  assign sdata_out_payload_74_real = data_mid_74_real;
  assign sdata_out_payload_74_imag = data_mid_74_imag;
  assign sdata_out_payload_75_real = data_mid_75_real;
  assign sdata_out_payload_75_imag = data_mid_75_imag;
  assign sdata_out_payload_76_real = data_mid_76_real;
  assign sdata_out_payload_76_imag = data_mid_76_imag;
  assign sdata_out_payload_77_real = data_mid_77_real;
  assign sdata_out_payload_77_imag = data_mid_77_imag;
  assign sdata_out_payload_78_real = data_mid_78_real;
  assign sdata_out_payload_78_imag = data_mid_78_imag;
  assign sdata_out_payload_79_real = data_mid_79_real;
  assign sdata_out_payload_79_imag = data_mid_79_imag;
  assign sdata_out_payload_80_real = data_mid_80_real;
  assign sdata_out_payload_80_imag = data_mid_80_imag;
  assign sdata_out_payload_81_real = data_mid_81_real;
  assign sdata_out_payload_81_imag = data_mid_81_imag;
  assign sdata_out_payload_82_real = data_mid_82_real;
  assign sdata_out_payload_82_imag = data_mid_82_imag;
  assign sdata_out_payload_83_real = data_mid_83_real;
  assign sdata_out_payload_83_imag = data_mid_83_imag;
  assign sdata_out_payload_84_real = data_mid_84_real;
  assign sdata_out_payload_84_imag = data_mid_84_imag;
  assign sdata_out_payload_85_real = data_mid_85_real;
  assign sdata_out_payload_85_imag = data_mid_85_imag;
  assign sdata_out_payload_86_real = data_mid_86_real;
  assign sdata_out_payload_86_imag = data_mid_86_imag;
  assign sdata_out_payload_87_real = data_mid_87_real;
  assign sdata_out_payload_87_imag = data_mid_87_imag;
  assign sdata_out_payload_88_real = data_mid_88_real;
  assign sdata_out_payload_88_imag = data_mid_88_imag;
  assign sdata_out_payload_89_real = data_mid_89_real;
  assign sdata_out_payload_89_imag = data_mid_89_imag;
  assign sdata_out_payload_90_real = data_mid_90_real;
  assign sdata_out_payload_90_imag = data_mid_90_imag;
  assign sdata_out_payload_91_real = data_mid_91_real;
  assign sdata_out_payload_91_imag = data_mid_91_imag;
  assign sdata_out_payload_92_real = data_mid_92_real;
  assign sdata_out_payload_92_imag = data_mid_92_imag;
  assign sdata_out_payload_93_real = data_mid_93_real;
  assign sdata_out_payload_93_imag = data_mid_93_imag;
  assign sdata_out_payload_94_real = data_mid_94_real;
  assign sdata_out_payload_94_imag = data_mid_94_imag;
  assign sdata_out_payload_95_real = data_mid_95_real;
  assign sdata_out_payload_95_imag = data_mid_95_imag;
  assign sdata_out_payload_96_real = data_mid_96_real;
  assign sdata_out_payload_96_imag = data_mid_96_imag;
  assign sdata_out_payload_97_real = data_mid_97_real;
  assign sdata_out_payload_97_imag = data_mid_97_imag;
  assign sdata_out_payload_98_real = data_mid_98_real;
  assign sdata_out_payload_98_imag = data_mid_98_imag;
  assign sdata_out_payload_99_real = data_mid_99_real;
  assign sdata_out_payload_99_imag = data_mid_99_imag;
  assign sdata_out_payload_100_real = data_mid_100_real;
  assign sdata_out_payload_100_imag = data_mid_100_imag;
  assign sdata_out_payload_101_real = data_mid_101_real;
  assign sdata_out_payload_101_imag = data_mid_101_imag;
  assign sdata_out_payload_102_real = data_mid_102_real;
  assign sdata_out_payload_102_imag = data_mid_102_imag;
  assign sdata_out_payload_103_real = data_mid_103_real;
  assign sdata_out_payload_103_imag = data_mid_103_imag;
  assign sdata_out_payload_104_real = data_mid_104_real;
  assign sdata_out_payload_104_imag = data_mid_104_imag;
  assign sdata_out_payload_105_real = data_mid_105_real;
  assign sdata_out_payload_105_imag = data_mid_105_imag;
  assign sdata_out_payload_106_real = data_mid_106_real;
  assign sdata_out_payload_106_imag = data_mid_106_imag;
  assign sdata_out_payload_107_real = data_mid_107_real;
  assign sdata_out_payload_107_imag = data_mid_107_imag;
  assign sdata_out_payload_108_real = data_mid_108_real;
  assign sdata_out_payload_108_imag = data_mid_108_imag;
  assign sdata_out_payload_109_real = data_mid_109_real;
  assign sdata_out_payload_109_imag = data_mid_109_imag;
  assign sdata_out_payload_110_real = data_mid_110_real;
  assign sdata_out_payload_110_imag = data_mid_110_imag;
  assign sdata_out_payload_111_real = data_mid_111_real;
  assign sdata_out_payload_111_imag = data_mid_111_imag;
  assign sdata_out_payload_112_real = data_mid_112_real;
  assign sdata_out_payload_112_imag = data_mid_112_imag;
  assign sdata_out_payload_113_real = data_mid_113_real;
  assign sdata_out_payload_113_imag = data_mid_113_imag;
  assign sdata_out_payload_114_real = data_mid_114_real;
  assign sdata_out_payload_114_imag = data_mid_114_imag;
  assign sdata_out_payload_115_real = data_mid_115_real;
  assign sdata_out_payload_115_imag = data_mid_115_imag;
  assign sdata_out_payload_116_real = data_mid_116_real;
  assign sdata_out_payload_116_imag = data_mid_116_imag;
  assign sdata_out_payload_117_real = data_mid_117_real;
  assign sdata_out_payload_117_imag = data_mid_117_imag;
  assign sdata_out_payload_118_real = data_mid_118_real;
  assign sdata_out_payload_118_imag = data_mid_118_imag;
  assign sdata_out_payload_119_real = data_mid_119_real;
  assign sdata_out_payload_119_imag = data_mid_119_imag;
  assign sdata_out_payload_120_real = data_mid_120_real;
  assign sdata_out_payload_120_imag = data_mid_120_imag;
  assign sdata_out_payload_121_real = data_mid_121_real;
  assign sdata_out_payload_121_imag = data_mid_121_imag;
  assign sdata_out_payload_122_real = data_mid_122_real;
  assign sdata_out_payload_122_imag = data_mid_122_imag;
  assign sdata_out_payload_123_real = data_mid_123_real;
  assign sdata_out_payload_123_imag = data_mid_123_imag;
  assign sdata_out_payload_124_real = data_mid_124_real;
  assign sdata_out_payload_124_imag = data_mid_124_imag;
  assign sdata_out_payload_125_real = data_mid_125_real;
  assign sdata_out_payload_125_imag = data_mid_125_imag;
  assign sdata_out_payload_126_real = data_mid_126_real;
  assign sdata_out_payload_126_imag = data_mid_126_imag;
  assign sdata_out_payload_127_real = data_mid_127_real;
  assign sdata_out_payload_127_imag = data_mid_127_imag;
  always @ (posedge clk) begin
    if(io_data_in_valid)begin
      data_in_0_real <= io_data_in_payload_0_real;
      data_in_0_imag <= io_data_in_payload_0_imag;
      data_in_1_real <= io_data_in_payload_1_real;
      data_in_1_imag <= io_data_in_payload_1_imag;
      data_in_2_real <= io_data_in_payload_2_real;
      data_in_2_imag <= io_data_in_payload_2_imag;
      data_in_3_real <= io_data_in_payload_3_real;
      data_in_3_imag <= io_data_in_payload_3_imag;
      data_in_4_real <= io_data_in_payload_4_real;
      data_in_4_imag <= io_data_in_payload_4_imag;
      data_in_5_real <= io_data_in_payload_5_real;
      data_in_5_imag <= io_data_in_payload_5_imag;
      data_in_6_real <= io_data_in_payload_6_real;
      data_in_6_imag <= io_data_in_payload_6_imag;
      data_in_7_real <= io_data_in_payload_7_real;
      data_in_7_imag <= io_data_in_payload_7_imag;
      data_in_8_real <= io_data_in_payload_8_real;
      data_in_8_imag <= io_data_in_payload_8_imag;
      data_in_9_real <= io_data_in_payload_9_real;
      data_in_9_imag <= io_data_in_payload_9_imag;
      data_in_10_real <= io_data_in_payload_10_real;
      data_in_10_imag <= io_data_in_payload_10_imag;
      data_in_11_real <= io_data_in_payload_11_real;
      data_in_11_imag <= io_data_in_payload_11_imag;
      data_in_12_real <= io_data_in_payload_12_real;
      data_in_12_imag <= io_data_in_payload_12_imag;
      data_in_13_real <= io_data_in_payload_13_real;
      data_in_13_imag <= io_data_in_payload_13_imag;
      data_in_14_real <= io_data_in_payload_14_real;
      data_in_14_imag <= io_data_in_payload_14_imag;
      data_in_15_real <= io_data_in_payload_15_real;
      data_in_15_imag <= io_data_in_payload_15_imag;
      data_in_16_real <= io_data_in_payload_16_real;
      data_in_16_imag <= io_data_in_payload_16_imag;
      data_in_17_real <= io_data_in_payload_17_real;
      data_in_17_imag <= io_data_in_payload_17_imag;
      data_in_18_real <= io_data_in_payload_18_real;
      data_in_18_imag <= io_data_in_payload_18_imag;
      data_in_19_real <= io_data_in_payload_19_real;
      data_in_19_imag <= io_data_in_payload_19_imag;
      data_in_20_real <= io_data_in_payload_20_real;
      data_in_20_imag <= io_data_in_payload_20_imag;
      data_in_21_real <= io_data_in_payload_21_real;
      data_in_21_imag <= io_data_in_payload_21_imag;
      data_in_22_real <= io_data_in_payload_22_real;
      data_in_22_imag <= io_data_in_payload_22_imag;
      data_in_23_real <= io_data_in_payload_23_real;
      data_in_23_imag <= io_data_in_payload_23_imag;
      data_in_24_real <= io_data_in_payload_24_real;
      data_in_24_imag <= io_data_in_payload_24_imag;
      data_in_25_real <= io_data_in_payload_25_real;
      data_in_25_imag <= io_data_in_payload_25_imag;
      data_in_26_real <= io_data_in_payload_26_real;
      data_in_26_imag <= io_data_in_payload_26_imag;
      data_in_27_real <= io_data_in_payload_27_real;
      data_in_27_imag <= io_data_in_payload_27_imag;
      data_in_28_real <= io_data_in_payload_28_real;
      data_in_28_imag <= io_data_in_payload_28_imag;
      data_in_29_real <= io_data_in_payload_29_real;
      data_in_29_imag <= io_data_in_payload_29_imag;
      data_in_30_real <= io_data_in_payload_30_real;
      data_in_30_imag <= io_data_in_payload_30_imag;
      data_in_31_real <= io_data_in_payload_31_real;
      data_in_31_imag <= io_data_in_payload_31_imag;
      data_in_32_real <= io_data_in_payload_32_real;
      data_in_32_imag <= io_data_in_payload_32_imag;
      data_in_33_real <= io_data_in_payload_33_real;
      data_in_33_imag <= io_data_in_payload_33_imag;
      data_in_34_real <= io_data_in_payload_34_real;
      data_in_34_imag <= io_data_in_payload_34_imag;
      data_in_35_real <= io_data_in_payload_35_real;
      data_in_35_imag <= io_data_in_payload_35_imag;
      data_in_36_real <= io_data_in_payload_36_real;
      data_in_36_imag <= io_data_in_payload_36_imag;
      data_in_37_real <= io_data_in_payload_37_real;
      data_in_37_imag <= io_data_in_payload_37_imag;
      data_in_38_real <= io_data_in_payload_38_real;
      data_in_38_imag <= io_data_in_payload_38_imag;
      data_in_39_real <= io_data_in_payload_39_real;
      data_in_39_imag <= io_data_in_payload_39_imag;
      data_in_40_real <= io_data_in_payload_40_real;
      data_in_40_imag <= io_data_in_payload_40_imag;
      data_in_41_real <= io_data_in_payload_41_real;
      data_in_41_imag <= io_data_in_payload_41_imag;
      data_in_42_real <= io_data_in_payload_42_real;
      data_in_42_imag <= io_data_in_payload_42_imag;
      data_in_43_real <= io_data_in_payload_43_real;
      data_in_43_imag <= io_data_in_payload_43_imag;
      data_in_44_real <= io_data_in_payload_44_real;
      data_in_44_imag <= io_data_in_payload_44_imag;
      data_in_45_real <= io_data_in_payload_45_real;
      data_in_45_imag <= io_data_in_payload_45_imag;
      data_in_46_real <= io_data_in_payload_46_real;
      data_in_46_imag <= io_data_in_payload_46_imag;
      data_in_47_real <= io_data_in_payload_47_real;
      data_in_47_imag <= io_data_in_payload_47_imag;
      data_in_48_real <= io_data_in_payload_48_real;
      data_in_48_imag <= io_data_in_payload_48_imag;
      data_in_49_real <= io_data_in_payload_49_real;
      data_in_49_imag <= io_data_in_payload_49_imag;
      data_in_50_real <= io_data_in_payload_50_real;
      data_in_50_imag <= io_data_in_payload_50_imag;
      data_in_51_real <= io_data_in_payload_51_real;
      data_in_51_imag <= io_data_in_payload_51_imag;
      data_in_52_real <= io_data_in_payload_52_real;
      data_in_52_imag <= io_data_in_payload_52_imag;
      data_in_53_real <= io_data_in_payload_53_real;
      data_in_53_imag <= io_data_in_payload_53_imag;
      data_in_54_real <= io_data_in_payload_54_real;
      data_in_54_imag <= io_data_in_payload_54_imag;
      data_in_55_real <= io_data_in_payload_55_real;
      data_in_55_imag <= io_data_in_payload_55_imag;
      data_in_56_real <= io_data_in_payload_56_real;
      data_in_56_imag <= io_data_in_payload_56_imag;
      data_in_57_real <= io_data_in_payload_57_real;
      data_in_57_imag <= io_data_in_payload_57_imag;
      data_in_58_real <= io_data_in_payload_58_real;
      data_in_58_imag <= io_data_in_payload_58_imag;
      data_in_59_real <= io_data_in_payload_59_real;
      data_in_59_imag <= io_data_in_payload_59_imag;
      data_in_60_real <= io_data_in_payload_60_real;
      data_in_60_imag <= io_data_in_payload_60_imag;
      data_in_61_real <= io_data_in_payload_61_real;
      data_in_61_imag <= io_data_in_payload_61_imag;
      data_in_62_real <= io_data_in_payload_62_real;
      data_in_62_imag <= io_data_in_payload_62_imag;
      data_in_63_real <= io_data_in_payload_63_real;
      data_in_63_imag <= io_data_in_payload_63_imag;
      data_in_64_real <= io_data_in_payload_64_real;
      data_in_64_imag <= io_data_in_payload_64_imag;
      data_in_65_real <= io_data_in_payload_65_real;
      data_in_65_imag <= io_data_in_payload_65_imag;
      data_in_66_real <= io_data_in_payload_66_real;
      data_in_66_imag <= io_data_in_payload_66_imag;
      data_in_67_real <= io_data_in_payload_67_real;
      data_in_67_imag <= io_data_in_payload_67_imag;
      data_in_68_real <= io_data_in_payload_68_real;
      data_in_68_imag <= io_data_in_payload_68_imag;
      data_in_69_real <= io_data_in_payload_69_real;
      data_in_69_imag <= io_data_in_payload_69_imag;
      data_in_70_real <= io_data_in_payload_70_real;
      data_in_70_imag <= io_data_in_payload_70_imag;
      data_in_71_real <= io_data_in_payload_71_real;
      data_in_71_imag <= io_data_in_payload_71_imag;
      data_in_72_real <= io_data_in_payload_72_real;
      data_in_72_imag <= io_data_in_payload_72_imag;
      data_in_73_real <= io_data_in_payload_73_real;
      data_in_73_imag <= io_data_in_payload_73_imag;
      data_in_74_real <= io_data_in_payload_74_real;
      data_in_74_imag <= io_data_in_payload_74_imag;
      data_in_75_real <= io_data_in_payload_75_real;
      data_in_75_imag <= io_data_in_payload_75_imag;
      data_in_76_real <= io_data_in_payload_76_real;
      data_in_76_imag <= io_data_in_payload_76_imag;
      data_in_77_real <= io_data_in_payload_77_real;
      data_in_77_imag <= io_data_in_payload_77_imag;
      data_in_78_real <= io_data_in_payload_78_real;
      data_in_78_imag <= io_data_in_payload_78_imag;
      data_in_79_real <= io_data_in_payload_79_real;
      data_in_79_imag <= io_data_in_payload_79_imag;
      data_in_80_real <= io_data_in_payload_80_real;
      data_in_80_imag <= io_data_in_payload_80_imag;
      data_in_81_real <= io_data_in_payload_81_real;
      data_in_81_imag <= io_data_in_payload_81_imag;
      data_in_82_real <= io_data_in_payload_82_real;
      data_in_82_imag <= io_data_in_payload_82_imag;
      data_in_83_real <= io_data_in_payload_83_real;
      data_in_83_imag <= io_data_in_payload_83_imag;
      data_in_84_real <= io_data_in_payload_84_real;
      data_in_84_imag <= io_data_in_payload_84_imag;
      data_in_85_real <= io_data_in_payload_85_real;
      data_in_85_imag <= io_data_in_payload_85_imag;
      data_in_86_real <= io_data_in_payload_86_real;
      data_in_86_imag <= io_data_in_payload_86_imag;
      data_in_87_real <= io_data_in_payload_87_real;
      data_in_87_imag <= io_data_in_payload_87_imag;
      data_in_88_real <= io_data_in_payload_88_real;
      data_in_88_imag <= io_data_in_payload_88_imag;
      data_in_89_real <= io_data_in_payload_89_real;
      data_in_89_imag <= io_data_in_payload_89_imag;
      data_in_90_real <= io_data_in_payload_90_real;
      data_in_90_imag <= io_data_in_payload_90_imag;
      data_in_91_real <= io_data_in_payload_91_real;
      data_in_91_imag <= io_data_in_payload_91_imag;
      data_in_92_real <= io_data_in_payload_92_real;
      data_in_92_imag <= io_data_in_payload_92_imag;
      data_in_93_real <= io_data_in_payload_93_real;
      data_in_93_imag <= io_data_in_payload_93_imag;
      data_in_94_real <= io_data_in_payload_94_real;
      data_in_94_imag <= io_data_in_payload_94_imag;
      data_in_95_real <= io_data_in_payload_95_real;
      data_in_95_imag <= io_data_in_payload_95_imag;
      data_in_96_real <= io_data_in_payload_96_real;
      data_in_96_imag <= io_data_in_payload_96_imag;
      data_in_97_real <= io_data_in_payload_97_real;
      data_in_97_imag <= io_data_in_payload_97_imag;
      data_in_98_real <= io_data_in_payload_98_real;
      data_in_98_imag <= io_data_in_payload_98_imag;
      data_in_99_real <= io_data_in_payload_99_real;
      data_in_99_imag <= io_data_in_payload_99_imag;
      data_in_100_real <= io_data_in_payload_100_real;
      data_in_100_imag <= io_data_in_payload_100_imag;
      data_in_101_real <= io_data_in_payload_101_real;
      data_in_101_imag <= io_data_in_payload_101_imag;
      data_in_102_real <= io_data_in_payload_102_real;
      data_in_102_imag <= io_data_in_payload_102_imag;
      data_in_103_real <= io_data_in_payload_103_real;
      data_in_103_imag <= io_data_in_payload_103_imag;
      data_in_104_real <= io_data_in_payload_104_real;
      data_in_104_imag <= io_data_in_payload_104_imag;
      data_in_105_real <= io_data_in_payload_105_real;
      data_in_105_imag <= io_data_in_payload_105_imag;
      data_in_106_real <= io_data_in_payload_106_real;
      data_in_106_imag <= io_data_in_payload_106_imag;
      data_in_107_real <= io_data_in_payload_107_real;
      data_in_107_imag <= io_data_in_payload_107_imag;
      data_in_108_real <= io_data_in_payload_108_real;
      data_in_108_imag <= io_data_in_payload_108_imag;
      data_in_109_real <= io_data_in_payload_109_real;
      data_in_109_imag <= io_data_in_payload_109_imag;
      data_in_110_real <= io_data_in_payload_110_real;
      data_in_110_imag <= io_data_in_payload_110_imag;
      data_in_111_real <= io_data_in_payload_111_real;
      data_in_111_imag <= io_data_in_payload_111_imag;
      data_in_112_real <= io_data_in_payload_112_real;
      data_in_112_imag <= io_data_in_payload_112_imag;
      data_in_113_real <= io_data_in_payload_113_real;
      data_in_113_imag <= io_data_in_payload_113_imag;
      data_in_114_real <= io_data_in_payload_114_real;
      data_in_114_imag <= io_data_in_payload_114_imag;
      data_in_115_real <= io_data_in_payload_115_real;
      data_in_115_imag <= io_data_in_payload_115_imag;
      data_in_116_real <= io_data_in_payload_116_real;
      data_in_116_imag <= io_data_in_payload_116_imag;
      data_in_117_real <= io_data_in_payload_117_real;
      data_in_117_imag <= io_data_in_payload_117_imag;
      data_in_118_real <= io_data_in_payload_118_real;
      data_in_118_imag <= io_data_in_payload_118_imag;
      data_in_119_real <= io_data_in_payload_119_real;
      data_in_119_imag <= io_data_in_payload_119_imag;
      data_in_120_real <= io_data_in_payload_120_real;
      data_in_120_imag <= io_data_in_payload_120_imag;
      data_in_121_real <= io_data_in_payload_121_real;
      data_in_121_imag <= io_data_in_payload_121_imag;
      data_in_122_real <= io_data_in_payload_122_real;
      data_in_122_imag <= io_data_in_payload_122_imag;
      data_in_123_real <= io_data_in_payload_123_real;
      data_in_123_imag <= io_data_in_payload_123_imag;
      data_in_124_real <= io_data_in_payload_124_real;
      data_in_124_imag <= io_data_in_payload_124_imag;
      data_in_125_real <= io_data_in_payload_125_real;
      data_in_125_imag <= io_data_in_payload_125_imag;
      data_in_126_real <= io_data_in_payload_126_real;
      data_in_126_imag <= io_data_in_payload_126_imag;
      data_in_127_real <= io_data_in_payload_127_real;
      data_in_127_imag <= io_data_in_payload_127_imag;
    end
    if((current_level_value == 3'b000))begin
      data_mid_0_real <= data_reorder_0_real;
      data_mid_0_imag <= data_reorder_0_imag;
      data_mid_1_real <= data_reorder_1_real;
      data_mid_1_imag <= data_reorder_1_imag;
      data_mid_2_real <= data_reorder_2_real;
      data_mid_2_imag <= data_reorder_2_imag;
      data_mid_3_real <= data_reorder_3_real;
      data_mid_3_imag <= data_reorder_3_imag;
      data_mid_4_real <= data_reorder_4_real;
      data_mid_4_imag <= data_reorder_4_imag;
      data_mid_5_real <= data_reorder_5_real;
      data_mid_5_imag <= data_reorder_5_imag;
      data_mid_6_real <= data_reorder_6_real;
      data_mid_6_imag <= data_reorder_6_imag;
      data_mid_7_real <= data_reorder_7_real;
      data_mid_7_imag <= data_reorder_7_imag;
      data_mid_8_real <= data_reorder_8_real;
      data_mid_8_imag <= data_reorder_8_imag;
      data_mid_9_real <= data_reorder_9_real;
      data_mid_9_imag <= data_reorder_9_imag;
      data_mid_10_real <= data_reorder_10_real;
      data_mid_10_imag <= data_reorder_10_imag;
      data_mid_11_real <= data_reorder_11_real;
      data_mid_11_imag <= data_reorder_11_imag;
      data_mid_12_real <= data_reorder_12_real;
      data_mid_12_imag <= data_reorder_12_imag;
      data_mid_13_real <= data_reorder_13_real;
      data_mid_13_imag <= data_reorder_13_imag;
      data_mid_14_real <= data_reorder_14_real;
      data_mid_14_imag <= data_reorder_14_imag;
      data_mid_15_real <= data_reorder_15_real;
      data_mid_15_imag <= data_reorder_15_imag;
      data_mid_16_real <= data_reorder_16_real;
      data_mid_16_imag <= data_reorder_16_imag;
      data_mid_17_real <= data_reorder_17_real;
      data_mid_17_imag <= data_reorder_17_imag;
      data_mid_18_real <= data_reorder_18_real;
      data_mid_18_imag <= data_reorder_18_imag;
      data_mid_19_real <= data_reorder_19_real;
      data_mid_19_imag <= data_reorder_19_imag;
      data_mid_20_real <= data_reorder_20_real;
      data_mid_20_imag <= data_reorder_20_imag;
      data_mid_21_real <= data_reorder_21_real;
      data_mid_21_imag <= data_reorder_21_imag;
      data_mid_22_real <= data_reorder_22_real;
      data_mid_22_imag <= data_reorder_22_imag;
      data_mid_23_real <= data_reorder_23_real;
      data_mid_23_imag <= data_reorder_23_imag;
      data_mid_24_real <= data_reorder_24_real;
      data_mid_24_imag <= data_reorder_24_imag;
      data_mid_25_real <= data_reorder_25_real;
      data_mid_25_imag <= data_reorder_25_imag;
      data_mid_26_real <= data_reorder_26_real;
      data_mid_26_imag <= data_reorder_26_imag;
      data_mid_27_real <= data_reorder_27_real;
      data_mid_27_imag <= data_reorder_27_imag;
      data_mid_28_real <= data_reorder_28_real;
      data_mid_28_imag <= data_reorder_28_imag;
      data_mid_29_real <= data_reorder_29_real;
      data_mid_29_imag <= data_reorder_29_imag;
      data_mid_30_real <= data_reorder_30_real;
      data_mid_30_imag <= data_reorder_30_imag;
      data_mid_31_real <= data_reorder_31_real;
      data_mid_31_imag <= data_reorder_31_imag;
      data_mid_32_real <= data_reorder_32_real;
      data_mid_32_imag <= data_reorder_32_imag;
      data_mid_33_real <= data_reorder_33_real;
      data_mid_33_imag <= data_reorder_33_imag;
      data_mid_34_real <= data_reorder_34_real;
      data_mid_34_imag <= data_reorder_34_imag;
      data_mid_35_real <= data_reorder_35_real;
      data_mid_35_imag <= data_reorder_35_imag;
      data_mid_36_real <= data_reorder_36_real;
      data_mid_36_imag <= data_reorder_36_imag;
      data_mid_37_real <= data_reorder_37_real;
      data_mid_37_imag <= data_reorder_37_imag;
      data_mid_38_real <= data_reorder_38_real;
      data_mid_38_imag <= data_reorder_38_imag;
      data_mid_39_real <= data_reorder_39_real;
      data_mid_39_imag <= data_reorder_39_imag;
      data_mid_40_real <= data_reorder_40_real;
      data_mid_40_imag <= data_reorder_40_imag;
      data_mid_41_real <= data_reorder_41_real;
      data_mid_41_imag <= data_reorder_41_imag;
      data_mid_42_real <= data_reorder_42_real;
      data_mid_42_imag <= data_reorder_42_imag;
      data_mid_43_real <= data_reorder_43_real;
      data_mid_43_imag <= data_reorder_43_imag;
      data_mid_44_real <= data_reorder_44_real;
      data_mid_44_imag <= data_reorder_44_imag;
      data_mid_45_real <= data_reorder_45_real;
      data_mid_45_imag <= data_reorder_45_imag;
      data_mid_46_real <= data_reorder_46_real;
      data_mid_46_imag <= data_reorder_46_imag;
      data_mid_47_real <= data_reorder_47_real;
      data_mid_47_imag <= data_reorder_47_imag;
      data_mid_48_real <= data_reorder_48_real;
      data_mid_48_imag <= data_reorder_48_imag;
      data_mid_49_real <= data_reorder_49_real;
      data_mid_49_imag <= data_reorder_49_imag;
      data_mid_50_real <= data_reorder_50_real;
      data_mid_50_imag <= data_reorder_50_imag;
      data_mid_51_real <= data_reorder_51_real;
      data_mid_51_imag <= data_reorder_51_imag;
      data_mid_52_real <= data_reorder_52_real;
      data_mid_52_imag <= data_reorder_52_imag;
      data_mid_53_real <= data_reorder_53_real;
      data_mid_53_imag <= data_reorder_53_imag;
      data_mid_54_real <= data_reorder_54_real;
      data_mid_54_imag <= data_reorder_54_imag;
      data_mid_55_real <= data_reorder_55_real;
      data_mid_55_imag <= data_reorder_55_imag;
      data_mid_56_real <= data_reorder_56_real;
      data_mid_56_imag <= data_reorder_56_imag;
      data_mid_57_real <= data_reorder_57_real;
      data_mid_57_imag <= data_reorder_57_imag;
      data_mid_58_real <= data_reorder_58_real;
      data_mid_58_imag <= data_reorder_58_imag;
      data_mid_59_real <= data_reorder_59_real;
      data_mid_59_imag <= data_reorder_59_imag;
      data_mid_60_real <= data_reorder_60_real;
      data_mid_60_imag <= data_reorder_60_imag;
      data_mid_61_real <= data_reorder_61_real;
      data_mid_61_imag <= data_reorder_61_imag;
      data_mid_62_real <= data_reorder_62_real;
      data_mid_62_imag <= data_reorder_62_imag;
      data_mid_63_real <= data_reorder_63_real;
      data_mid_63_imag <= data_reorder_63_imag;
      data_mid_64_real <= data_reorder_64_real;
      data_mid_64_imag <= data_reorder_64_imag;
      data_mid_65_real <= data_reorder_65_real;
      data_mid_65_imag <= data_reorder_65_imag;
      data_mid_66_real <= data_reorder_66_real;
      data_mid_66_imag <= data_reorder_66_imag;
      data_mid_67_real <= data_reorder_67_real;
      data_mid_67_imag <= data_reorder_67_imag;
      data_mid_68_real <= data_reorder_68_real;
      data_mid_68_imag <= data_reorder_68_imag;
      data_mid_69_real <= data_reorder_69_real;
      data_mid_69_imag <= data_reorder_69_imag;
      data_mid_70_real <= data_reorder_70_real;
      data_mid_70_imag <= data_reorder_70_imag;
      data_mid_71_real <= data_reorder_71_real;
      data_mid_71_imag <= data_reorder_71_imag;
      data_mid_72_real <= data_reorder_72_real;
      data_mid_72_imag <= data_reorder_72_imag;
      data_mid_73_real <= data_reorder_73_real;
      data_mid_73_imag <= data_reorder_73_imag;
      data_mid_74_real <= data_reorder_74_real;
      data_mid_74_imag <= data_reorder_74_imag;
      data_mid_75_real <= data_reorder_75_real;
      data_mid_75_imag <= data_reorder_75_imag;
      data_mid_76_real <= data_reorder_76_real;
      data_mid_76_imag <= data_reorder_76_imag;
      data_mid_77_real <= data_reorder_77_real;
      data_mid_77_imag <= data_reorder_77_imag;
      data_mid_78_real <= data_reorder_78_real;
      data_mid_78_imag <= data_reorder_78_imag;
      data_mid_79_real <= data_reorder_79_real;
      data_mid_79_imag <= data_reorder_79_imag;
      data_mid_80_real <= data_reorder_80_real;
      data_mid_80_imag <= data_reorder_80_imag;
      data_mid_81_real <= data_reorder_81_real;
      data_mid_81_imag <= data_reorder_81_imag;
      data_mid_82_real <= data_reorder_82_real;
      data_mid_82_imag <= data_reorder_82_imag;
      data_mid_83_real <= data_reorder_83_real;
      data_mid_83_imag <= data_reorder_83_imag;
      data_mid_84_real <= data_reorder_84_real;
      data_mid_84_imag <= data_reorder_84_imag;
      data_mid_85_real <= data_reorder_85_real;
      data_mid_85_imag <= data_reorder_85_imag;
      data_mid_86_real <= data_reorder_86_real;
      data_mid_86_imag <= data_reorder_86_imag;
      data_mid_87_real <= data_reorder_87_real;
      data_mid_87_imag <= data_reorder_87_imag;
      data_mid_88_real <= data_reorder_88_real;
      data_mid_88_imag <= data_reorder_88_imag;
      data_mid_89_real <= data_reorder_89_real;
      data_mid_89_imag <= data_reorder_89_imag;
      data_mid_90_real <= data_reorder_90_real;
      data_mid_90_imag <= data_reorder_90_imag;
      data_mid_91_real <= data_reorder_91_real;
      data_mid_91_imag <= data_reorder_91_imag;
      data_mid_92_real <= data_reorder_92_real;
      data_mid_92_imag <= data_reorder_92_imag;
      data_mid_93_real <= data_reorder_93_real;
      data_mid_93_imag <= data_reorder_93_imag;
      data_mid_94_real <= data_reorder_94_real;
      data_mid_94_imag <= data_reorder_94_imag;
      data_mid_95_real <= data_reorder_95_real;
      data_mid_95_imag <= data_reorder_95_imag;
      data_mid_96_real <= data_reorder_96_real;
      data_mid_96_imag <= data_reorder_96_imag;
      data_mid_97_real <= data_reorder_97_real;
      data_mid_97_imag <= data_reorder_97_imag;
      data_mid_98_real <= data_reorder_98_real;
      data_mid_98_imag <= data_reorder_98_imag;
      data_mid_99_real <= data_reorder_99_real;
      data_mid_99_imag <= data_reorder_99_imag;
      data_mid_100_real <= data_reorder_100_real;
      data_mid_100_imag <= data_reorder_100_imag;
      data_mid_101_real <= data_reorder_101_real;
      data_mid_101_imag <= data_reorder_101_imag;
      data_mid_102_real <= data_reorder_102_real;
      data_mid_102_imag <= data_reorder_102_imag;
      data_mid_103_real <= data_reorder_103_real;
      data_mid_103_imag <= data_reorder_103_imag;
      data_mid_104_real <= data_reorder_104_real;
      data_mid_104_imag <= data_reorder_104_imag;
      data_mid_105_real <= data_reorder_105_real;
      data_mid_105_imag <= data_reorder_105_imag;
      data_mid_106_real <= data_reorder_106_real;
      data_mid_106_imag <= data_reorder_106_imag;
      data_mid_107_real <= data_reorder_107_real;
      data_mid_107_imag <= data_reorder_107_imag;
      data_mid_108_real <= data_reorder_108_real;
      data_mid_108_imag <= data_reorder_108_imag;
      data_mid_109_real <= data_reorder_109_real;
      data_mid_109_imag <= data_reorder_109_imag;
      data_mid_110_real <= data_reorder_110_real;
      data_mid_110_imag <= data_reorder_110_imag;
      data_mid_111_real <= data_reorder_111_real;
      data_mid_111_imag <= data_reorder_111_imag;
      data_mid_112_real <= data_reorder_112_real;
      data_mid_112_imag <= data_reorder_112_imag;
      data_mid_113_real <= data_reorder_113_real;
      data_mid_113_imag <= data_reorder_113_imag;
      data_mid_114_real <= data_reorder_114_real;
      data_mid_114_imag <= data_reorder_114_imag;
      data_mid_115_real <= data_reorder_115_real;
      data_mid_115_imag <= data_reorder_115_imag;
      data_mid_116_real <= data_reorder_116_real;
      data_mid_116_imag <= data_reorder_116_imag;
      data_mid_117_real <= data_reorder_117_real;
      data_mid_117_imag <= data_reorder_117_imag;
      data_mid_118_real <= data_reorder_118_real;
      data_mid_118_imag <= data_reorder_118_imag;
      data_mid_119_real <= data_reorder_119_real;
      data_mid_119_imag <= data_reorder_119_imag;
      data_mid_120_real <= data_reorder_120_real;
      data_mid_120_imag <= data_reorder_120_imag;
      data_mid_121_real <= data_reorder_121_real;
      data_mid_121_imag <= data_reorder_121_imag;
      data_mid_122_real <= data_reorder_122_real;
      data_mid_122_imag <= data_reorder_122_imag;
      data_mid_123_real <= data_reorder_123_real;
      data_mid_123_imag <= data_reorder_123_imag;
      data_mid_124_real <= data_reorder_124_real;
      data_mid_124_imag <= data_reorder_124_imag;
      data_mid_125_real <= data_reorder_125_real;
      data_mid_125_imag <= data_reorder_125_imag;
      data_mid_126_real <= data_reorder_126_real;
      data_mid_126_imag <= data_reorder_126_imag;
      data_mid_127_real <= data_reorder_127_real;
      data_mid_127_imag <= data_reorder_127_imag;
    end else begin
      if((current_level_value == 3'b001))begin
        data_mid_1_real <= _zz_4947[15 : 0];
        data_mid_1_imag <= _zz_4955[15 : 0];
        data_mid_0_real <= _zz_4963[15 : 0];
        data_mid_0_imag <= _zz_4971[15 : 0];
      end
      if((current_level_value == 3'b001))begin
        data_mid_3_real <= _zz_4988[15 : 0];
        data_mid_3_imag <= _zz_4996[15 : 0];
        data_mid_2_real <= _zz_5004[15 : 0];
        data_mid_2_imag <= _zz_5012[15 : 0];
      end
      if((current_level_value == 3'b001))begin
        data_mid_5_real <= _zz_5029[15 : 0];
        data_mid_5_imag <= _zz_5037[15 : 0];
        data_mid_4_real <= _zz_5045[15 : 0];
        data_mid_4_imag <= _zz_5053[15 : 0];
      end
      if((current_level_value == 3'b001))begin
        data_mid_7_real <= _zz_5070[15 : 0];
        data_mid_7_imag <= _zz_5078[15 : 0];
        data_mid_6_real <= _zz_5086[15 : 0];
        data_mid_6_imag <= _zz_5094[15 : 0];
      end
      if((current_level_value == 3'b001))begin
        data_mid_9_real <= _zz_5111[15 : 0];
        data_mid_9_imag <= _zz_5119[15 : 0];
        data_mid_8_real <= _zz_5127[15 : 0];
        data_mid_8_imag <= _zz_5135[15 : 0];
      end
      if((current_level_value == 3'b001))begin
        data_mid_11_real <= _zz_5152[15 : 0];
        data_mid_11_imag <= _zz_5160[15 : 0];
        data_mid_10_real <= _zz_5168[15 : 0];
        data_mid_10_imag <= _zz_5176[15 : 0];
      end
      if((current_level_value == 3'b001))begin
        data_mid_13_real <= _zz_5193[15 : 0];
        data_mid_13_imag <= _zz_5201[15 : 0];
        data_mid_12_real <= _zz_5209[15 : 0];
        data_mid_12_imag <= _zz_5217[15 : 0];
      end
      if((current_level_value == 3'b001))begin
        data_mid_15_real <= _zz_5234[15 : 0];
        data_mid_15_imag <= _zz_5242[15 : 0];
        data_mid_14_real <= _zz_5250[15 : 0];
        data_mid_14_imag <= _zz_5258[15 : 0];
      end
      if((current_level_value == 3'b001))begin
        data_mid_17_real <= _zz_5275[15 : 0];
        data_mid_17_imag <= _zz_5283[15 : 0];
        data_mid_16_real <= _zz_5291[15 : 0];
        data_mid_16_imag <= _zz_5299[15 : 0];
      end
      if((current_level_value == 3'b001))begin
        data_mid_19_real <= _zz_5316[15 : 0];
        data_mid_19_imag <= _zz_5324[15 : 0];
        data_mid_18_real <= _zz_5332[15 : 0];
        data_mid_18_imag <= _zz_5340[15 : 0];
      end
      if((current_level_value == 3'b001))begin
        data_mid_21_real <= _zz_5357[15 : 0];
        data_mid_21_imag <= _zz_5365[15 : 0];
        data_mid_20_real <= _zz_5373[15 : 0];
        data_mid_20_imag <= _zz_5381[15 : 0];
      end
      if((current_level_value == 3'b001))begin
        data_mid_23_real <= _zz_5398[15 : 0];
        data_mid_23_imag <= _zz_5406[15 : 0];
        data_mid_22_real <= _zz_5414[15 : 0];
        data_mid_22_imag <= _zz_5422[15 : 0];
      end
      if((current_level_value == 3'b001))begin
        data_mid_25_real <= _zz_5439[15 : 0];
        data_mid_25_imag <= _zz_5447[15 : 0];
        data_mid_24_real <= _zz_5455[15 : 0];
        data_mid_24_imag <= _zz_5463[15 : 0];
      end
      if((current_level_value == 3'b001))begin
        data_mid_27_real <= _zz_5480[15 : 0];
        data_mid_27_imag <= _zz_5488[15 : 0];
        data_mid_26_real <= _zz_5496[15 : 0];
        data_mid_26_imag <= _zz_5504[15 : 0];
      end
      if((current_level_value == 3'b001))begin
        data_mid_29_real <= _zz_5521[15 : 0];
        data_mid_29_imag <= _zz_5529[15 : 0];
        data_mid_28_real <= _zz_5537[15 : 0];
        data_mid_28_imag <= _zz_5545[15 : 0];
      end
      if((current_level_value == 3'b001))begin
        data_mid_31_real <= _zz_5562[15 : 0];
        data_mid_31_imag <= _zz_5570[15 : 0];
        data_mid_30_real <= _zz_5578[15 : 0];
        data_mid_30_imag <= _zz_5586[15 : 0];
      end
      if((current_level_value == 3'b001))begin
        data_mid_33_real <= _zz_5603[15 : 0];
        data_mid_33_imag <= _zz_5611[15 : 0];
        data_mid_32_real <= _zz_5619[15 : 0];
        data_mid_32_imag <= _zz_5627[15 : 0];
      end
      if((current_level_value == 3'b001))begin
        data_mid_35_real <= _zz_5644[15 : 0];
        data_mid_35_imag <= _zz_5652[15 : 0];
        data_mid_34_real <= _zz_5660[15 : 0];
        data_mid_34_imag <= _zz_5668[15 : 0];
      end
      if((current_level_value == 3'b001))begin
        data_mid_37_real <= _zz_5685[15 : 0];
        data_mid_37_imag <= _zz_5693[15 : 0];
        data_mid_36_real <= _zz_5701[15 : 0];
        data_mid_36_imag <= _zz_5709[15 : 0];
      end
      if((current_level_value == 3'b001))begin
        data_mid_39_real <= _zz_5726[15 : 0];
        data_mid_39_imag <= _zz_5734[15 : 0];
        data_mid_38_real <= _zz_5742[15 : 0];
        data_mid_38_imag <= _zz_5750[15 : 0];
      end
      if((current_level_value == 3'b001))begin
        data_mid_41_real <= _zz_5767[15 : 0];
        data_mid_41_imag <= _zz_5775[15 : 0];
        data_mid_40_real <= _zz_5783[15 : 0];
        data_mid_40_imag <= _zz_5791[15 : 0];
      end
      if((current_level_value == 3'b001))begin
        data_mid_43_real <= _zz_5808[15 : 0];
        data_mid_43_imag <= _zz_5816[15 : 0];
        data_mid_42_real <= _zz_5824[15 : 0];
        data_mid_42_imag <= _zz_5832[15 : 0];
      end
      if((current_level_value == 3'b001))begin
        data_mid_45_real <= _zz_5849[15 : 0];
        data_mid_45_imag <= _zz_5857[15 : 0];
        data_mid_44_real <= _zz_5865[15 : 0];
        data_mid_44_imag <= _zz_5873[15 : 0];
      end
      if((current_level_value == 3'b001))begin
        data_mid_47_real <= _zz_5890[15 : 0];
        data_mid_47_imag <= _zz_5898[15 : 0];
        data_mid_46_real <= _zz_5906[15 : 0];
        data_mid_46_imag <= _zz_5914[15 : 0];
      end
      if((current_level_value == 3'b001))begin
        data_mid_49_real <= _zz_5931[15 : 0];
        data_mid_49_imag <= _zz_5939[15 : 0];
        data_mid_48_real <= _zz_5947[15 : 0];
        data_mid_48_imag <= _zz_5955[15 : 0];
      end
      if((current_level_value == 3'b001))begin
        data_mid_51_real <= _zz_5972[15 : 0];
        data_mid_51_imag <= _zz_5980[15 : 0];
        data_mid_50_real <= _zz_5988[15 : 0];
        data_mid_50_imag <= _zz_5996[15 : 0];
      end
      if((current_level_value == 3'b001))begin
        data_mid_53_real <= _zz_6013[15 : 0];
        data_mid_53_imag <= _zz_6021[15 : 0];
        data_mid_52_real <= _zz_6029[15 : 0];
        data_mid_52_imag <= _zz_6037[15 : 0];
      end
      if((current_level_value == 3'b001))begin
        data_mid_55_real <= _zz_6054[15 : 0];
        data_mid_55_imag <= _zz_6062[15 : 0];
        data_mid_54_real <= _zz_6070[15 : 0];
        data_mid_54_imag <= _zz_6078[15 : 0];
      end
      if((current_level_value == 3'b001))begin
        data_mid_57_real <= _zz_6095[15 : 0];
        data_mid_57_imag <= _zz_6103[15 : 0];
        data_mid_56_real <= _zz_6111[15 : 0];
        data_mid_56_imag <= _zz_6119[15 : 0];
      end
      if((current_level_value == 3'b001))begin
        data_mid_59_real <= _zz_6136[15 : 0];
        data_mid_59_imag <= _zz_6144[15 : 0];
        data_mid_58_real <= _zz_6152[15 : 0];
        data_mid_58_imag <= _zz_6160[15 : 0];
      end
      if((current_level_value == 3'b001))begin
        data_mid_61_real <= _zz_6177[15 : 0];
        data_mid_61_imag <= _zz_6185[15 : 0];
        data_mid_60_real <= _zz_6193[15 : 0];
        data_mid_60_imag <= _zz_6201[15 : 0];
      end
      if((current_level_value == 3'b001))begin
        data_mid_63_real <= _zz_6218[15 : 0];
        data_mid_63_imag <= _zz_6226[15 : 0];
        data_mid_62_real <= _zz_6234[15 : 0];
        data_mid_62_imag <= _zz_6242[15 : 0];
      end
      if((current_level_value == 3'b001))begin
        data_mid_65_real <= _zz_6259[15 : 0];
        data_mid_65_imag <= _zz_6267[15 : 0];
        data_mid_64_real <= _zz_6275[15 : 0];
        data_mid_64_imag <= _zz_6283[15 : 0];
      end
      if((current_level_value == 3'b001))begin
        data_mid_67_real <= _zz_6300[15 : 0];
        data_mid_67_imag <= _zz_6308[15 : 0];
        data_mid_66_real <= _zz_6316[15 : 0];
        data_mid_66_imag <= _zz_6324[15 : 0];
      end
      if((current_level_value == 3'b001))begin
        data_mid_69_real <= _zz_6341[15 : 0];
        data_mid_69_imag <= _zz_6349[15 : 0];
        data_mid_68_real <= _zz_6357[15 : 0];
        data_mid_68_imag <= _zz_6365[15 : 0];
      end
      if((current_level_value == 3'b001))begin
        data_mid_71_real <= _zz_6382[15 : 0];
        data_mid_71_imag <= _zz_6390[15 : 0];
        data_mid_70_real <= _zz_6398[15 : 0];
        data_mid_70_imag <= _zz_6406[15 : 0];
      end
      if((current_level_value == 3'b001))begin
        data_mid_73_real <= _zz_6423[15 : 0];
        data_mid_73_imag <= _zz_6431[15 : 0];
        data_mid_72_real <= _zz_6439[15 : 0];
        data_mid_72_imag <= _zz_6447[15 : 0];
      end
      if((current_level_value == 3'b001))begin
        data_mid_75_real <= _zz_6464[15 : 0];
        data_mid_75_imag <= _zz_6472[15 : 0];
        data_mid_74_real <= _zz_6480[15 : 0];
        data_mid_74_imag <= _zz_6488[15 : 0];
      end
      if((current_level_value == 3'b001))begin
        data_mid_77_real <= _zz_6505[15 : 0];
        data_mid_77_imag <= _zz_6513[15 : 0];
        data_mid_76_real <= _zz_6521[15 : 0];
        data_mid_76_imag <= _zz_6529[15 : 0];
      end
      if((current_level_value == 3'b001))begin
        data_mid_79_real <= _zz_6546[15 : 0];
        data_mid_79_imag <= _zz_6554[15 : 0];
        data_mid_78_real <= _zz_6562[15 : 0];
        data_mid_78_imag <= _zz_6570[15 : 0];
      end
      if((current_level_value == 3'b001))begin
        data_mid_81_real <= _zz_6587[15 : 0];
        data_mid_81_imag <= _zz_6595[15 : 0];
        data_mid_80_real <= _zz_6603[15 : 0];
        data_mid_80_imag <= _zz_6611[15 : 0];
      end
      if((current_level_value == 3'b001))begin
        data_mid_83_real <= _zz_6628[15 : 0];
        data_mid_83_imag <= _zz_6636[15 : 0];
        data_mid_82_real <= _zz_6644[15 : 0];
        data_mid_82_imag <= _zz_6652[15 : 0];
      end
      if((current_level_value == 3'b001))begin
        data_mid_85_real <= _zz_6669[15 : 0];
        data_mid_85_imag <= _zz_6677[15 : 0];
        data_mid_84_real <= _zz_6685[15 : 0];
        data_mid_84_imag <= _zz_6693[15 : 0];
      end
      if((current_level_value == 3'b001))begin
        data_mid_87_real <= _zz_6710[15 : 0];
        data_mid_87_imag <= _zz_6718[15 : 0];
        data_mid_86_real <= _zz_6726[15 : 0];
        data_mid_86_imag <= _zz_6734[15 : 0];
      end
      if((current_level_value == 3'b001))begin
        data_mid_89_real <= _zz_6751[15 : 0];
        data_mid_89_imag <= _zz_6759[15 : 0];
        data_mid_88_real <= _zz_6767[15 : 0];
        data_mid_88_imag <= _zz_6775[15 : 0];
      end
      if((current_level_value == 3'b001))begin
        data_mid_91_real <= _zz_6792[15 : 0];
        data_mid_91_imag <= _zz_6800[15 : 0];
        data_mid_90_real <= _zz_6808[15 : 0];
        data_mid_90_imag <= _zz_6816[15 : 0];
      end
      if((current_level_value == 3'b001))begin
        data_mid_93_real <= _zz_6833[15 : 0];
        data_mid_93_imag <= _zz_6841[15 : 0];
        data_mid_92_real <= _zz_6849[15 : 0];
        data_mid_92_imag <= _zz_6857[15 : 0];
      end
      if((current_level_value == 3'b001))begin
        data_mid_95_real <= _zz_6874[15 : 0];
        data_mid_95_imag <= _zz_6882[15 : 0];
        data_mid_94_real <= _zz_6890[15 : 0];
        data_mid_94_imag <= _zz_6898[15 : 0];
      end
      if((current_level_value == 3'b001))begin
        data_mid_97_real <= _zz_6915[15 : 0];
        data_mid_97_imag <= _zz_6923[15 : 0];
        data_mid_96_real <= _zz_6931[15 : 0];
        data_mid_96_imag <= _zz_6939[15 : 0];
      end
      if((current_level_value == 3'b001))begin
        data_mid_99_real <= _zz_6956[15 : 0];
        data_mid_99_imag <= _zz_6964[15 : 0];
        data_mid_98_real <= _zz_6972[15 : 0];
        data_mid_98_imag <= _zz_6980[15 : 0];
      end
      if((current_level_value == 3'b001))begin
        data_mid_101_real <= _zz_6997[15 : 0];
        data_mid_101_imag <= _zz_7005[15 : 0];
        data_mid_100_real <= _zz_7013[15 : 0];
        data_mid_100_imag <= _zz_7021[15 : 0];
      end
      if((current_level_value == 3'b001))begin
        data_mid_103_real <= _zz_7038[15 : 0];
        data_mid_103_imag <= _zz_7046[15 : 0];
        data_mid_102_real <= _zz_7054[15 : 0];
        data_mid_102_imag <= _zz_7062[15 : 0];
      end
      if((current_level_value == 3'b001))begin
        data_mid_105_real <= _zz_7079[15 : 0];
        data_mid_105_imag <= _zz_7087[15 : 0];
        data_mid_104_real <= _zz_7095[15 : 0];
        data_mid_104_imag <= _zz_7103[15 : 0];
      end
      if((current_level_value == 3'b001))begin
        data_mid_107_real <= _zz_7120[15 : 0];
        data_mid_107_imag <= _zz_7128[15 : 0];
        data_mid_106_real <= _zz_7136[15 : 0];
        data_mid_106_imag <= _zz_7144[15 : 0];
      end
      if((current_level_value == 3'b001))begin
        data_mid_109_real <= _zz_7161[15 : 0];
        data_mid_109_imag <= _zz_7169[15 : 0];
        data_mid_108_real <= _zz_7177[15 : 0];
        data_mid_108_imag <= _zz_7185[15 : 0];
      end
      if((current_level_value == 3'b001))begin
        data_mid_111_real <= _zz_7202[15 : 0];
        data_mid_111_imag <= _zz_7210[15 : 0];
        data_mid_110_real <= _zz_7218[15 : 0];
        data_mid_110_imag <= _zz_7226[15 : 0];
      end
      if((current_level_value == 3'b001))begin
        data_mid_113_real <= _zz_7243[15 : 0];
        data_mid_113_imag <= _zz_7251[15 : 0];
        data_mid_112_real <= _zz_7259[15 : 0];
        data_mid_112_imag <= _zz_7267[15 : 0];
      end
      if((current_level_value == 3'b001))begin
        data_mid_115_real <= _zz_7284[15 : 0];
        data_mid_115_imag <= _zz_7292[15 : 0];
        data_mid_114_real <= _zz_7300[15 : 0];
        data_mid_114_imag <= _zz_7308[15 : 0];
      end
      if((current_level_value == 3'b001))begin
        data_mid_117_real <= _zz_7325[15 : 0];
        data_mid_117_imag <= _zz_7333[15 : 0];
        data_mid_116_real <= _zz_7341[15 : 0];
        data_mid_116_imag <= _zz_7349[15 : 0];
      end
      if((current_level_value == 3'b001))begin
        data_mid_119_real <= _zz_7366[15 : 0];
        data_mid_119_imag <= _zz_7374[15 : 0];
        data_mid_118_real <= _zz_7382[15 : 0];
        data_mid_118_imag <= _zz_7390[15 : 0];
      end
      if((current_level_value == 3'b001))begin
        data_mid_121_real <= _zz_7407[15 : 0];
        data_mid_121_imag <= _zz_7415[15 : 0];
        data_mid_120_real <= _zz_7423[15 : 0];
        data_mid_120_imag <= _zz_7431[15 : 0];
      end
      if((current_level_value == 3'b001))begin
        data_mid_123_real <= _zz_7448[15 : 0];
        data_mid_123_imag <= _zz_7456[15 : 0];
        data_mid_122_real <= _zz_7464[15 : 0];
        data_mid_122_imag <= _zz_7472[15 : 0];
      end
      if((current_level_value == 3'b001))begin
        data_mid_125_real <= _zz_7489[15 : 0];
        data_mid_125_imag <= _zz_7497[15 : 0];
        data_mid_124_real <= _zz_7505[15 : 0];
        data_mid_124_imag <= _zz_7513[15 : 0];
      end
      if((current_level_value == 3'b001))begin
        data_mid_127_real <= _zz_7530[15 : 0];
        data_mid_127_imag <= _zz_7538[15 : 0];
        data_mid_126_real <= _zz_7546[15 : 0];
        data_mid_126_imag <= _zz_7554[15 : 0];
      end
      if((current_level_value == 3'b010))begin
        data_mid_2_real <= _zz_7571[15 : 0];
        data_mid_2_imag <= _zz_7579[15 : 0];
        data_mid_0_real <= _zz_7587[15 : 0];
        data_mid_0_imag <= _zz_7595[15 : 0];
      end
      if((current_level_value == 3'b010))begin
        data_mid_3_real <= _zz_7612[15 : 0];
        data_mid_3_imag <= _zz_7620[15 : 0];
        data_mid_1_real <= _zz_7628[15 : 0];
        data_mid_1_imag <= _zz_7636[15 : 0];
      end
      if((current_level_value == 3'b010))begin
        data_mid_6_real <= _zz_7653[15 : 0];
        data_mid_6_imag <= _zz_7661[15 : 0];
        data_mid_4_real <= _zz_7669[15 : 0];
        data_mid_4_imag <= _zz_7677[15 : 0];
      end
      if((current_level_value == 3'b010))begin
        data_mid_7_real <= _zz_7694[15 : 0];
        data_mid_7_imag <= _zz_7702[15 : 0];
        data_mid_5_real <= _zz_7710[15 : 0];
        data_mid_5_imag <= _zz_7718[15 : 0];
      end
      if((current_level_value == 3'b010))begin
        data_mid_10_real <= _zz_7735[15 : 0];
        data_mid_10_imag <= _zz_7743[15 : 0];
        data_mid_8_real <= _zz_7751[15 : 0];
        data_mid_8_imag <= _zz_7759[15 : 0];
      end
      if((current_level_value == 3'b010))begin
        data_mid_11_real <= _zz_7776[15 : 0];
        data_mid_11_imag <= _zz_7784[15 : 0];
        data_mid_9_real <= _zz_7792[15 : 0];
        data_mid_9_imag <= _zz_7800[15 : 0];
      end
      if((current_level_value == 3'b010))begin
        data_mid_14_real <= _zz_7817[15 : 0];
        data_mid_14_imag <= _zz_7825[15 : 0];
        data_mid_12_real <= _zz_7833[15 : 0];
        data_mid_12_imag <= _zz_7841[15 : 0];
      end
      if((current_level_value == 3'b010))begin
        data_mid_15_real <= _zz_7858[15 : 0];
        data_mid_15_imag <= _zz_7866[15 : 0];
        data_mid_13_real <= _zz_7874[15 : 0];
        data_mid_13_imag <= _zz_7882[15 : 0];
      end
      if((current_level_value == 3'b010))begin
        data_mid_18_real <= _zz_7899[15 : 0];
        data_mid_18_imag <= _zz_7907[15 : 0];
        data_mid_16_real <= _zz_7915[15 : 0];
        data_mid_16_imag <= _zz_7923[15 : 0];
      end
      if((current_level_value == 3'b010))begin
        data_mid_19_real <= _zz_7940[15 : 0];
        data_mid_19_imag <= _zz_7948[15 : 0];
        data_mid_17_real <= _zz_7956[15 : 0];
        data_mid_17_imag <= _zz_7964[15 : 0];
      end
      if((current_level_value == 3'b010))begin
        data_mid_22_real <= _zz_7981[15 : 0];
        data_mid_22_imag <= _zz_7989[15 : 0];
        data_mid_20_real <= _zz_7997[15 : 0];
        data_mid_20_imag <= _zz_8005[15 : 0];
      end
      if((current_level_value == 3'b010))begin
        data_mid_23_real <= _zz_8022[15 : 0];
        data_mid_23_imag <= _zz_8030[15 : 0];
        data_mid_21_real <= _zz_8038[15 : 0];
        data_mid_21_imag <= _zz_8046[15 : 0];
      end
      if((current_level_value == 3'b010))begin
        data_mid_26_real <= _zz_8063[15 : 0];
        data_mid_26_imag <= _zz_8071[15 : 0];
        data_mid_24_real <= _zz_8079[15 : 0];
        data_mid_24_imag <= _zz_8087[15 : 0];
      end
      if((current_level_value == 3'b010))begin
        data_mid_27_real <= _zz_8104[15 : 0];
        data_mid_27_imag <= _zz_8112[15 : 0];
        data_mid_25_real <= _zz_8120[15 : 0];
        data_mid_25_imag <= _zz_8128[15 : 0];
      end
      if((current_level_value == 3'b010))begin
        data_mid_30_real <= _zz_8145[15 : 0];
        data_mid_30_imag <= _zz_8153[15 : 0];
        data_mid_28_real <= _zz_8161[15 : 0];
        data_mid_28_imag <= _zz_8169[15 : 0];
      end
      if((current_level_value == 3'b010))begin
        data_mid_31_real <= _zz_8186[15 : 0];
        data_mid_31_imag <= _zz_8194[15 : 0];
        data_mid_29_real <= _zz_8202[15 : 0];
        data_mid_29_imag <= _zz_8210[15 : 0];
      end
      if((current_level_value == 3'b010))begin
        data_mid_34_real <= _zz_8227[15 : 0];
        data_mid_34_imag <= _zz_8235[15 : 0];
        data_mid_32_real <= _zz_8243[15 : 0];
        data_mid_32_imag <= _zz_8251[15 : 0];
      end
      if((current_level_value == 3'b010))begin
        data_mid_35_real <= _zz_8268[15 : 0];
        data_mid_35_imag <= _zz_8276[15 : 0];
        data_mid_33_real <= _zz_8284[15 : 0];
        data_mid_33_imag <= _zz_8292[15 : 0];
      end
      if((current_level_value == 3'b010))begin
        data_mid_38_real <= _zz_8309[15 : 0];
        data_mid_38_imag <= _zz_8317[15 : 0];
        data_mid_36_real <= _zz_8325[15 : 0];
        data_mid_36_imag <= _zz_8333[15 : 0];
      end
      if((current_level_value == 3'b010))begin
        data_mid_39_real <= _zz_8350[15 : 0];
        data_mid_39_imag <= _zz_8358[15 : 0];
        data_mid_37_real <= _zz_8366[15 : 0];
        data_mid_37_imag <= _zz_8374[15 : 0];
      end
      if((current_level_value == 3'b010))begin
        data_mid_42_real <= _zz_8391[15 : 0];
        data_mid_42_imag <= _zz_8399[15 : 0];
        data_mid_40_real <= _zz_8407[15 : 0];
        data_mid_40_imag <= _zz_8415[15 : 0];
      end
      if((current_level_value == 3'b010))begin
        data_mid_43_real <= _zz_8432[15 : 0];
        data_mid_43_imag <= _zz_8440[15 : 0];
        data_mid_41_real <= _zz_8448[15 : 0];
        data_mid_41_imag <= _zz_8456[15 : 0];
      end
      if((current_level_value == 3'b010))begin
        data_mid_46_real <= _zz_8473[15 : 0];
        data_mid_46_imag <= _zz_8481[15 : 0];
        data_mid_44_real <= _zz_8489[15 : 0];
        data_mid_44_imag <= _zz_8497[15 : 0];
      end
      if((current_level_value == 3'b010))begin
        data_mid_47_real <= _zz_8514[15 : 0];
        data_mid_47_imag <= _zz_8522[15 : 0];
        data_mid_45_real <= _zz_8530[15 : 0];
        data_mid_45_imag <= _zz_8538[15 : 0];
      end
      if((current_level_value == 3'b010))begin
        data_mid_50_real <= _zz_8555[15 : 0];
        data_mid_50_imag <= _zz_8563[15 : 0];
        data_mid_48_real <= _zz_8571[15 : 0];
        data_mid_48_imag <= _zz_8579[15 : 0];
      end
      if((current_level_value == 3'b010))begin
        data_mid_51_real <= _zz_8596[15 : 0];
        data_mid_51_imag <= _zz_8604[15 : 0];
        data_mid_49_real <= _zz_8612[15 : 0];
        data_mid_49_imag <= _zz_8620[15 : 0];
      end
      if((current_level_value == 3'b010))begin
        data_mid_54_real <= _zz_8637[15 : 0];
        data_mid_54_imag <= _zz_8645[15 : 0];
        data_mid_52_real <= _zz_8653[15 : 0];
        data_mid_52_imag <= _zz_8661[15 : 0];
      end
      if((current_level_value == 3'b010))begin
        data_mid_55_real <= _zz_8678[15 : 0];
        data_mid_55_imag <= _zz_8686[15 : 0];
        data_mid_53_real <= _zz_8694[15 : 0];
        data_mid_53_imag <= _zz_8702[15 : 0];
      end
      if((current_level_value == 3'b010))begin
        data_mid_58_real <= _zz_8719[15 : 0];
        data_mid_58_imag <= _zz_8727[15 : 0];
        data_mid_56_real <= _zz_8735[15 : 0];
        data_mid_56_imag <= _zz_8743[15 : 0];
      end
      if((current_level_value == 3'b010))begin
        data_mid_59_real <= _zz_8760[15 : 0];
        data_mid_59_imag <= _zz_8768[15 : 0];
        data_mid_57_real <= _zz_8776[15 : 0];
        data_mid_57_imag <= _zz_8784[15 : 0];
      end
      if((current_level_value == 3'b010))begin
        data_mid_62_real <= _zz_8801[15 : 0];
        data_mid_62_imag <= _zz_8809[15 : 0];
        data_mid_60_real <= _zz_8817[15 : 0];
        data_mid_60_imag <= _zz_8825[15 : 0];
      end
      if((current_level_value == 3'b010))begin
        data_mid_63_real <= _zz_8842[15 : 0];
        data_mid_63_imag <= _zz_8850[15 : 0];
        data_mid_61_real <= _zz_8858[15 : 0];
        data_mid_61_imag <= _zz_8866[15 : 0];
      end
      if((current_level_value == 3'b010))begin
        data_mid_66_real <= _zz_8883[15 : 0];
        data_mid_66_imag <= _zz_8891[15 : 0];
        data_mid_64_real <= _zz_8899[15 : 0];
        data_mid_64_imag <= _zz_8907[15 : 0];
      end
      if((current_level_value == 3'b010))begin
        data_mid_67_real <= _zz_8924[15 : 0];
        data_mid_67_imag <= _zz_8932[15 : 0];
        data_mid_65_real <= _zz_8940[15 : 0];
        data_mid_65_imag <= _zz_8948[15 : 0];
      end
      if((current_level_value == 3'b010))begin
        data_mid_70_real <= _zz_8965[15 : 0];
        data_mid_70_imag <= _zz_8973[15 : 0];
        data_mid_68_real <= _zz_8981[15 : 0];
        data_mid_68_imag <= _zz_8989[15 : 0];
      end
      if((current_level_value == 3'b010))begin
        data_mid_71_real <= _zz_9006[15 : 0];
        data_mid_71_imag <= _zz_9014[15 : 0];
        data_mid_69_real <= _zz_9022[15 : 0];
        data_mid_69_imag <= _zz_9030[15 : 0];
      end
      if((current_level_value == 3'b010))begin
        data_mid_74_real <= _zz_9047[15 : 0];
        data_mid_74_imag <= _zz_9055[15 : 0];
        data_mid_72_real <= _zz_9063[15 : 0];
        data_mid_72_imag <= _zz_9071[15 : 0];
      end
      if((current_level_value == 3'b010))begin
        data_mid_75_real <= _zz_9088[15 : 0];
        data_mid_75_imag <= _zz_9096[15 : 0];
        data_mid_73_real <= _zz_9104[15 : 0];
        data_mid_73_imag <= _zz_9112[15 : 0];
      end
      if((current_level_value == 3'b010))begin
        data_mid_78_real <= _zz_9129[15 : 0];
        data_mid_78_imag <= _zz_9137[15 : 0];
        data_mid_76_real <= _zz_9145[15 : 0];
        data_mid_76_imag <= _zz_9153[15 : 0];
      end
      if((current_level_value == 3'b010))begin
        data_mid_79_real <= _zz_9170[15 : 0];
        data_mid_79_imag <= _zz_9178[15 : 0];
        data_mid_77_real <= _zz_9186[15 : 0];
        data_mid_77_imag <= _zz_9194[15 : 0];
      end
      if((current_level_value == 3'b010))begin
        data_mid_82_real <= _zz_9211[15 : 0];
        data_mid_82_imag <= _zz_9219[15 : 0];
        data_mid_80_real <= _zz_9227[15 : 0];
        data_mid_80_imag <= _zz_9235[15 : 0];
      end
      if((current_level_value == 3'b010))begin
        data_mid_83_real <= _zz_9252[15 : 0];
        data_mid_83_imag <= _zz_9260[15 : 0];
        data_mid_81_real <= _zz_9268[15 : 0];
        data_mid_81_imag <= _zz_9276[15 : 0];
      end
      if((current_level_value == 3'b010))begin
        data_mid_86_real <= _zz_9293[15 : 0];
        data_mid_86_imag <= _zz_9301[15 : 0];
        data_mid_84_real <= _zz_9309[15 : 0];
        data_mid_84_imag <= _zz_9317[15 : 0];
      end
      if((current_level_value == 3'b010))begin
        data_mid_87_real <= _zz_9334[15 : 0];
        data_mid_87_imag <= _zz_9342[15 : 0];
        data_mid_85_real <= _zz_9350[15 : 0];
        data_mid_85_imag <= _zz_9358[15 : 0];
      end
      if((current_level_value == 3'b010))begin
        data_mid_90_real <= _zz_9375[15 : 0];
        data_mid_90_imag <= _zz_9383[15 : 0];
        data_mid_88_real <= _zz_9391[15 : 0];
        data_mid_88_imag <= _zz_9399[15 : 0];
      end
      if((current_level_value == 3'b010))begin
        data_mid_91_real <= _zz_9416[15 : 0];
        data_mid_91_imag <= _zz_9424[15 : 0];
        data_mid_89_real <= _zz_9432[15 : 0];
        data_mid_89_imag <= _zz_9440[15 : 0];
      end
      if((current_level_value == 3'b010))begin
        data_mid_94_real <= _zz_9457[15 : 0];
        data_mid_94_imag <= _zz_9465[15 : 0];
        data_mid_92_real <= _zz_9473[15 : 0];
        data_mid_92_imag <= _zz_9481[15 : 0];
      end
      if((current_level_value == 3'b010))begin
        data_mid_95_real <= _zz_9498[15 : 0];
        data_mid_95_imag <= _zz_9506[15 : 0];
        data_mid_93_real <= _zz_9514[15 : 0];
        data_mid_93_imag <= _zz_9522[15 : 0];
      end
      if((current_level_value == 3'b010))begin
        data_mid_98_real <= _zz_9539[15 : 0];
        data_mid_98_imag <= _zz_9547[15 : 0];
        data_mid_96_real <= _zz_9555[15 : 0];
        data_mid_96_imag <= _zz_9563[15 : 0];
      end
      if((current_level_value == 3'b010))begin
        data_mid_99_real <= _zz_9580[15 : 0];
        data_mid_99_imag <= _zz_9588[15 : 0];
        data_mid_97_real <= _zz_9596[15 : 0];
        data_mid_97_imag <= _zz_9604[15 : 0];
      end
      if((current_level_value == 3'b010))begin
        data_mid_102_real <= _zz_9621[15 : 0];
        data_mid_102_imag <= _zz_9629[15 : 0];
        data_mid_100_real <= _zz_9637[15 : 0];
        data_mid_100_imag <= _zz_9645[15 : 0];
      end
      if((current_level_value == 3'b010))begin
        data_mid_103_real <= _zz_9662[15 : 0];
        data_mid_103_imag <= _zz_9670[15 : 0];
        data_mid_101_real <= _zz_9678[15 : 0];
        data_mid_101_imag <= _zz_9686[15 : 0];
      end
      if((current_level_value == 3'b010))begin
        data_mid_106_real <= _zz_9703[15 : 0];
        data_mid_106_imag <= _zz_9711[15 : 0];
        data_mid_104_real <= _zz_9719[15 : 0];
        data_mid_104_imag <= _zz_9727[15 : 0];
      end
      if((current_level_value == 3'b010))begin
        data_mid_107_real <= _zz_9744[15 : 0];
        data_mid_107_imag <= _zz_9752[15 : 0];
        data_mid_105_real <= _zz_9760[15 : 0];
        data_mid_105_imag <= _zz_9768[15 : 0];
      end
      if((current_level_value == 3'b010))begin
        data_mid_110_real <= _zz_9785[15 : 0];
        data_mid_110_imag <= _zz_9793[15 : 0];
        data_mid_108_real <= _zz_9801[15 : 0];
        data_mid_108_imag <= _zz_9809[15 : 0];
      end
      if((current_level_value == 3'b010))begin
        data_mid_111_real <= _zz_9826[15 : 0];
        data_mid_111_imag <= _zz_9834[15 : 0];
        data_mid_109_real <= _zz_9842[15 : 0];
        data_mid_109_imag <= _zz_9850[15 : 0];
      end
      if((current_level_value == 3'b010))begin
        data_mid_114_real <= _zz_9867[15 : 0];
        data_mid_114_imag <= _zz_9875[15 : 0];
        data_mid_112_real <= _zz_9883[15 : 0];
        data_mid_112_imag <= _zz_9891[15 : 0];
      end
      if((current_level_value == 3'b010))begin
        data_mid_115_real <= _zz_9908[15 : 0];
        data_mid_115_imag <= _zz_9916[15 : 0];
        data_mid_113_real <= _zz_9924[15 : 0];
        data_mid_113_imag <= _zz_9932[15 : 0];
      end
      if((current_level_value == 3'b010))begin
        data_mid_118_real <= _zz_9949[15 : 0];
        data_mid_118_imag <= _zz_9957[15 : 0];
        data_mid_116_real <= _zz_9965[15 : 0];
        data_mid_116_imag <= _zz_9973[15 : 0];
      end
      if((current_level_value == 3'b010))begin
        data_mid_119_real <= _zz_9990[15 : 0];
        data_mid_119_imag <= _zz_9998[15 : 0];
        data_mid_117_real <= _zz_10006[15 : 0];
        data_mid_117_imag <= _zz_10014[15 : 0];
      end
      if((current_level_value == 3'b010))begin
        data_mid_122_real <= _zz_10031[15 : 0];
        data_mid_122_imag <= _zz_10039[15 : 0];
        data_mid_120_real <= _zz_10047[15 : 0];
        data_mid_120_imag <= _zz_10055[15 : 0];
      end
      if((current_level_value == 3'b010))begin
        data_mid_123_real <= _zz_10072[15 : 0];
        data_mid_123_imag <= _zz_10080[15 : 0];
        data_mid_121_real <= _zz_10088[15 : 0];
        data_mid_121_imag <= _zz_10096[15 : 0];
      end
      if((current_level_value == 3'b010))begin
        data_mid_126_real <= _zz_10113[15 : 0];
        data_mid_126_imag <= _zz_10121[15 : 0];
        data_mid_124_real <= _zz_10129[15 : 0];
        data_mid_124_imag <= _zz_10137[15 : 0];
      end
      if((current_level_value == 3'b010))begin
        data_mid_127_real <= _zz_10154[15 : 0];
        data_mid_127_imag <= _zz_10162[15 : 0];
        data_mid_125_real <= _zz_10170[15 : 0];
        data_mid_125_imag <= _zz_10178[15 : 0];
      end
      if((current_level_value == 3'b011))begin
        data_mid_4_real <= _zz_10195[15 : 0];
        data_mid_4_imag <= _zz_10203[15 : 0];
        data_mid_0_real <= _zz_10211[15 : 0];
        data_mid_0_imag <= _zz_10219[15 : 0];
      end
      if((current_level_value == 3'b011))begin
        data_mid_5_real <= _zz_10236[15 : 0];
        data_mid_5_imag <= _zz_10244[15 : 0];
        data_mid_1_real <= _zz_10252[15 : 0];
        data_mid_1_imag <= _zz_10260[15 : 0];
      end
      if((current_level_value == 3'b011))begin
        data_mid_6_real <= _zz_10277[15 : 0];
        data_mid_6_imag <= _zz_10285[15 : 0];
        data_mid_2_real <= _zz_10293[15 : 0];
        data_mid_2_imag <= _zz_10301[15 : 0];
      end
      if((current_level_value == 3'b011))begin
        data_mid_7_real <= _zz_10318[15 : 0];
        data_mid_7_imag <= _zz_10326[15 : 0];
        data_mid_3_real <= _zz_10334[15 : 0];
        data_mid_3_imag <= _zz_10342[15 : 0];
      end
      if((current_level_value == 3'b011))begin
        data_mid_12_real <= _zz_10359[15 : 0];
        data_mid_12_imag <= _zz_10367[15 : 0];
        data_mid_8_real <= _zz_10375[15 : 0];
        data_mid_8_imag <= _zz_10383[15 : 0];
      end
      if((current_level_value == 3'b011))begin
        data_mid_13_real <= _zz_10400[15 : 0];
        data_mid_13_imag <= _zz_10408[15 : 0];
        data_mid_9_real <= _zz_10416[15 : 0];
        data_mid_9_imag <= _zz_10424[15 : 0];
      end
      if((current_level_value == 3'b011))begin
        data_mid_14_real <= _zz_10441[15 : 0];
        data_mid_14_imag <= _zz_10449[15 : 0];
        data_mid_10_real <= _zz_10457[15 : 0];
        data_mid_10_imag <= _zz_10465[15 : 0];
      end
      if((current_level_value == 3'b011))begin
        data_mid_15_real <= _zz_10482[15 : 0];
        data_mid_15_imag <= _zz_10490[15 : 0];
        data_mid_11_real <= _zz_10498[15 : 0];
        data_mid_11_imag <= _zz_10506[15 : 0];
      end
      if((current_level_value == 3'b011))begin
        data_mid_20_real <= _zz_10523[15 : 0];
        data_mid_20_imag <= _zz_10531[15 : 0];
        data_mid_16_real <= _zz_10539[15 : 0];
        data_mid_16_imag <= _zz_10547[15 : 0];
      end
      if((current_level_value == 3'b011))begin
        data_mid_21_real <= _zz_10564[15 : 0];
        data_mid_21_imag <= _zz_10572[15 : 0];
        data_mid_17_real <= _zz_10580[15 : 0];
        data_mid_17_imag <= _zz_10588[15 : 0];
      end
      if((current_level_value == 3'b011))begin
        data_mid_22_real <= _zz_10605[15 : 0];
        data_mid_22_imag <= _zz_10613[15 : 0];
        data_mid_18_real <= _zz_10621[15 : 0];
        data_mid_18_imag <= _zz_10629[15 : 0];
      end
      if((current_level_value == 3'b011))begin
        data_mid_23_real <= _zz_10646[15 : 0];
        data_mid_23_imag <= _zz_10654[15 : 0];
        data_mid_19_real <= _zz_10662[15 : 0];
        data_mid_19_imag <= _zz_10670[15 : 0];
      end
      if((current_level_value == 3'b011))begin
        data_mid_28_real <= _zz_10687[15 : 0];
        data_mid_28_imag <= _zz_10695[15 : 0];
        data_mid_24_real <= _zz_10703[15 : 0];
        data_mid_24_imag <= _zz_10711[15 : 0];
      end
      if((current_level_value == 3'b011))begin
        data_mid_29_real <= _zz_10728[15 : 0];
        data_mid_29_imag <= _zz_10736[15 : 0];
        data_mid_25_real <= _zz_10744[15 : 0];
        data_mid_25_imag <= _zz_10752[15 : 0];
      end
      if((current_level_value == 3'b011))begin
        data_mid_30_real <= _zz_10769[15 : 0];
        data_mid_30_imag <= _zz_10777[15 : 0];
        data_mid_26_real <= _zz_10785[15 : 0];
        data_mid_26_imag <= _zz_10793[15 : 0];
      end
      if((current_level_value == 3'b011))begin
        data_mid_31_real <= _zz_10810[15 : 0];
        data_mid_31_imag <= _zz_10818[15 : 0];
        data_mid_27_real <= _zz_10826[15 : 0];
        data_mid_27_imag <= _zz_10834[15 : 0];
      end
      if((current_level_value == 3'b011))begin
        data_mid_36_real <= _zz_10851[15 : 0];
        data_mid_36_imag <= _zz_10859[15 : 0];
        data_mid_32_real <= _zz_10867[15 : 0];
        data_mid_32_imag <= _zz_10875[15 : 0];
      end
      if((current_level_value == 3'b011))begin
        data_mid_37_real <= _zz_10892[15 : 0];
        data_mid_37_imag <= _zz_10900[15 : 0];
        data_mid_33_real <= _zz_10908[15 : 0];
        data_mid_33_imag <= _zz_10916[15 : 0];
      end
      if((current_level_value == 3'b011))begin
        data_mid_38_real <= _zz_10933[15 : 0];
        data_mid_38_imag <= _zz_10941[15 : 0];
        data_mid_34_real <= _zz_10949[15 : 0];
        data_mid_34_imag <= _zz_10957[15 : 0];
      end
      if((current_level_value == 3'b011))begin
        data_mid_39_real <= _zz_10974[15 : 0];
        data_mid_39_imag <= _zz_10982[15 : 0];
        data_mid_35_real <= _zz_10990[15 : 0];
        data_mid_35_imag <= _zz_10998[15 : 0];
      end
      if((current_level_value == 3'b011))begin
        data_mid_44_real <= _zz_11015[15 : 0];
        data_mid_44_imag <= _zz_11023[15 : 0];
        data_mid_40_real <= _zz_11031[15 : 0];
        data_mid_40_imag <= _zz_11039[15 : 0];
      end
      if((current_level_value == 3'b011))begin
        data_mid_45_real <= _zz_11056[15 : 0];
        data_mid_45_imag <= _zz_11064[15 : 0];
        data_mid_41_real <= _zz_11072[15 : 0];
        data_mid_41_imag <= _zz_11080[15 : 0];
      end
      if((current_level_value == 3'b011))begin
        data_mid_46_real <= _zz_11097[15 : 0];
        data_mid_46_imag <= _zz_11105[15 : 0];
        data_mid_42_real <= _zz_11113[15 : 0];
        data_mid_42_imag <= _zz_11121[15 : 0];
      end
      if((current_level_value == 3'b011))begin
        data_mid_47_real <= _zz_11138[15 : 0];
        data_mid_47_imag <= _zz_11146[15 : 0];
        data_mid_43_real <= _zz_11154[15 : 0];
        data_mid_43_imag <= _zz_11162[15 : 0];
      end
      if((current_level_value == 3'b011))begin
        data_mid_52_real <= _zz_11179[15 : 0];
        data_mid_52_imag <= _zz_11187[15 : 0];
        data_mid_48_real <= _zz_11195[15 : 0];
        data_mid_48_imag <= _zz_11203[15 : 0];
      end
      if((current_level_value == 3'b011))begin
        data_mid_53_real <= _zz_11220[15 : 0];
        data_mid_53_imag <= _zz_11228[15 : 0];
        data_mid_49_real <= _zz_11236[15 : 0];
        data_mid_49_imag <= _zz_11244[15 : 0];
      end
      if((current_level_value == 3'b011))begin
        data_mid_54_real <= _zz_11261[15 : 0];
        data_mid_54_imag <= _zz_11269[15 : 0];
        data_mid_50_real <= _zz_11277[15 : 0];
        data_mid_50_imag <= _zz_11285[15 : 0];
      end
      if((current_level_value == 3'b011))begin
        data_mid_55_real <= _zz_11302[15 : 0];
        data_mid_55_imag <= _zz_11310[15 : 0];
        data_mid_51_real <= _zz_11318[15 : 0];
        data_mid_51_imag <= _zz_11326[15 : 0];
      end
      if((current_level_value == 3'b011))begin
        data_mid_60_real <= _zz_11343[15 : 0];
        data_mid_60_imag <= _zz_11351[15 : 0];
        data_mid_56_real <= _zz_11359[15 : 0];
        data_mid_56_imag <= _zz_11367[15 : 0];
      end
      if((current_level_value == 3'b011))begin
        data_mid_61_real <= _zz_11384[15 : 0];
        data_mid_61_imag <= _zz_11392[15 : 0];
        data_mid_57_real <= _zz_11400[15 : 0];
        data_mid_57_imag <= _zz_11408[15 : 0];
      end
      if((current_level_value == 3'b011))begin
        data_mid_62_real <= _zz_11425[15 : 0];
        data_mid_62_imag <= _zz_11433[15 : 0];
        data_mid_58_real <= _zz_11441[15 : 0];
        data_mid_58_imag <= _zz_11449[15 : 0];
      end
      if((current_level_value == 3'b011))begin
        data_mid_63_real <= _zz_11466[15 : 0];
        data_mid_63_imag <= _zz_11474[15 : 0];
        data_mid_59_real <= _zz_11482[15 : 0];
        data_mid_59_imag <= _zz_11490[15 : 0];
      end
      if((current_level_value == 3'b011))begin
        data_mid_68_real <= _zz_11507[15 : 0];
        data_mid_68_imag <= _zz_11515[15 : 0];
        data_mid_64_real <= _zz_11523[15 : 0];
        data_mid_64_imag <= _zz_11531[15 : 0];
      end
      if((current_level_value == 3'b011))begin
        data_mid_69_real <= _zz_11548[15 : 0];
        data_mid_69_imag <= _zz_11556[15 : 0];
        data_mid_65_real <= _zz_11564[15 : 0];
        data_mid_65_imag <= _zz_11572[15 : 0];
      end
      if((current_level_value == 3'b011))begin
        data_mid_70_real <= _zz_11589[15 : 0];
        data_mid_70_imag <= _zz_11597[15 : 0];
        data_mid_66_real <= _zz_11605[15 : 0];
        data_mid_66_imag <= _zz_11613[15 : 0];
      end
      if((current_level_value == 3'b011))begin
        data_mid_71_real <= _zz_11630[15 : 0];
        data_mid_71_imag <= _zz_11638[15 : 0];
        data_mid_67_real <= _zz_11646[15 : 0];
        data_mid_67_imag <= _zz_11654[15 : 0];
      end
      if((current_level_value == 3'b011))begin
        data_mid_76_real <= _zz_11671[15 : 0];
        data_mid_76_imag <= _zz_11679[15 : 0];
        data_mid_72_real <= _zz_11687[15 : 0];
        data_mid_72_imag <= _zz_11695[15 : 0];
      end
      if((current_level_value == 3'b011))begin
        data_mid_77_real <= _zz_11712[15 : 0];
        data_mid_77_imag <= _zz_11720[15 : 0];
        data_mid_73_real <= _zz_11728[15 : 0];
        data_mid_73_imag <= _zz_11736[15 : 0];
      end
      if((current_level_value == 3'b011))begin
        data_mid_78_real <= _zz_11753[15 : 0];
        data_mid_78_imag <= _zz_11761[15 : 0];
        data_mid_74_real <= _zz_11769[15 : 0];
        data_mid_74_imag <= _zz_11777[15 : 0];
      end
      if((current_level_value == 3'b011))begin
        data_mid_79_real <= _zz_11794[15 : 0];
        data_mid_79_imag <= _zz_11802[15 : 0];
        data_mid_75_real <= _zz_11810[15 : 0];
        data_mid_75_imag <= _zz_11818[15 : 0];
      end
      if((current_level_value == 3'b011))begin
        data_mid_84_real <= _zz_11835[15 : 0];
        data_mid_84_imag <= _zz_11843[15 : 0];
        data_mid_80_real <= _zz_11851[15 : 0];
        data_mid_80_imag <= _zz_11859[15 : 0];
      end
      if((current_level_value == 3'b011))begin
        data_mid_85_real <= _zz_11876[15 : 0];
        data_mid_85_imag <= _zz_11884[15 : 0];
        data_mid_81_real <= _zz_11892[15 : 0];
        data_mid_81_imag <= _zz_11900[15 : 0];
      end
      if((current_level_value == 3'b011))begin
        data_mid_86_real <= _zz_11917[15 : 0];
        data_mid_86_imag <= _zz_11925[15 : 0];
        data_mid_82_real <= _zz_11933[15 : 0];
        data_mid_82_imag <= _zz_11941[15 : 0];
      end
      if((current_level_value == 3'b011))begin
        data_mid_87_real <= _zz_11958[15 : 0];
        data_mid_87_imag <= _zz_11966[15 : 0];
        data_mid_83_real <= _zz_11974[15 : 0];
        data_mid_83_imag <= _zz_11982[15 : 0];
      end
      if((current_level_value == 3'b011))begin
        data_mid_92_real <= _zz_11999[15 : 0];
        data_mid_92_imag <= _zz_12007[15 : 0];
        data_mid_88_real <= _zz_12015[15 : 0];
        data_mid_88_imag <= _zz_12023[15 : 0];
      end
      if((current_level_value == 3'b011))begin
        data_mid_93_real <= _zz_12040[15 : 0];
        data_mid_93_imag <= _zz_12048[15 : 0];
        data_mid_89_real <= _zz_12056[15 : 0];
        data_mid_89_imag <= _zz_12064[15 : 0];
      end
      if((current_level_value == 3'b011))begin
        data_mid_94_real <= _zz_12081[15 : 0];
        data_mid_94_imag <= _zz_12089[15 : 0];
        data_mid_90_real <= _zz_12097[15 : 0];
        data_mid_90_imag <= _zz_12105[15 : 0];
      end
      if((current_level_value == 3'b011))begin
        data_mid_95_real <= _zz_12122[15 : 0];
        data_mid_95_imag <= _zz_12130[15 : 0];
        data_mid_91_real <= _zz_12138[15 : 0];
        data_mid_91_imag <= _zz_12146[15 : 0];
      end
      if((current_level_value == 3'b011))begin
        data_mid_100_real <= _zz_12163[15 : 0];
        data_mid_100_imag <= _zz_12171[15 : 0];
        data_mid_96_real <= _zz_12179[15 : 0];
        data_mid_96_imag <= _zz_12187[15 : 0];
      end
      if((current_level_value == 3'b011))begin
        data_mid_101_real <= _zz_12204[15 : 0];
        data_mid_101_imag <= _zz_12212[15 : 0];
        data_mid_97_real <= _zz_12220[15 : 0];
        data_mid_97_imag <= _zz_12228[15 : 0];
      end
      if((current_level_value == 3'b011))begin
        data_mid_102_real <= _zz_12245[15 : 0];
        data_mid_102_imag <= _zz_12253[15 : 0];
        data_mid_98_real <= _zz_12261[15 : 0];
        data_mid_98_imag <= _zz_12269[15 : 0];
      end
      if((current_level_value == 3'b011))begin
        data_mid_103_real <= _zz_12286[15 : 0];
        data_mid_103_imag <= _zz_12294[15 : 0];
        data_mid_99_real <= _zz_12302[15 : 0];
        data_mid_99_imag <= _zz_12310[15 : 0];
      end
      if((current_level_value == 3'b011))begin
        data_mid_108_real <= _zz_12327[15 : 0];
        data_mid_108_imag <= _zz_12335[15 : 0];
        data_mid_104_real <= _zz_12343[15 : 0];
        data_mid_104_imag <= _zz_12351[15 : 0];
      end
      if((current_level_value == 3'b011))begin
        data_mid_109_real <= _zz_12368[15 : 0];
        data_mid_109_imag <= _zz_12376[15 : 0];
        data_mid_105_real <= _zz_12384[15 : 0];
        data_mid_105_imag <= _zz_12392[15 : 0];
      end
      if((current_level_value == 3'b011))begin
        data_mid_110_real <= _zz_12409[15 : 0];
        data_mid_110_imag <= _zz_12417[15 : 0];
        data_mid_106_real <= _zz_12425[15 : 0];
        data_mid_106_imag <= _zz_12433[15 : 0];
      end
      if((current_level_value == 3'b011))begin
        data_mid_111_real <= _zz_12450[15 : 0];
        data_mid_111_imag <= _zz_12458[15 : 0];
        data_mid_107_real <= _zz_12466[15 : 0];
        data_mid_107_imag <= _zz_12474[15 : 0];
      end
      if((current_level_value == 3'b011))begin
        data_mid_116_real <= _zz_12491[15 : 0];
        data_mid_116_imag <= _zz_12499[15 : 0];
        data_mid_112_real <= _zz_12507[15 : 0];
        data_mid_112_imag <= _zz_12515[15 : 0];
      end
      if((current_level_value == 3'b011))begin
        data_mid_117_real <= _zz_12532[15 : 0];
        data_mid_117_imag <= _zz_12540[15 : 0];
        data_mid_113_real <= _zz_12548[15 : 0];
        data_mid_113_imag <= _zz_12556[15 : 0];
      end
      if((current_level_value == 3'b011))begin
        data_mid_118_real <= _zz_12573[15 : 0];
        data_mid_118_imag <= _zz_12581[15 : 0];
        data_mid_114_real <= _zz_12589[15 : 0];
        data_mid_114_imag <= _zz_12597[15 : 0];
      end
      if((current_level_value == 3'b011))begin
        data_mid_119_real <= _zz_12614[15 : 0];
        data_mid_119_imag <= _zz_12622[15 : 0];
        data_mid_115_real <= _zz_12630[15 : 0];
        data_mid_115_imag <= _zz_12638[15 : 0];
      end
      if((current_level_value == 3'b011))begin
        data_mid_124_real <= _zz_12655[15 : 0];
        data_mid_124_imag <= _zz_12663[15 : 0];
        data_mid_120_real <= _zz_12671[15 : 0];
        data_mid_120_imag <= _zz_12679[15 : 0];
      end
      if((current_level_value == 3'b011))begin
        data_mid_125_real <= _zz_12696[15 : 0];
        data_mid_125_imag <= _zz_12704[15 : 0];
        data_mid_121_real <= _zz_12712[15 : 0];
        data_mid_121_imag <= _zz_12720[15 : 0];
      end
      if((current_level_value == 3'b011))begin
        data_mid_126_real <= _zz_12737[15 : 0];
        data_mid_126_imag <= _zz_12745[15 : 0];
        data_mid_122_real <= _zz_12753[15 : 0];
        data_mid_122_imag <= _zz_12761[15 : 0];
      end
      if((current_level_value == 3'b011))begin
        data_mid_127_real <= _zz_12778[15 : 0];
        data_mid_127_imag <= _zz_12786[15 : 0];
        data_mid_123_real <= _zz_12794[15 : 0];
        data_mid_123_imag <= _zz_12802[15 : 0];
      end
      if((current_level_value == 3'b100))begin
        data_mid_8_real <= _zz_12819[15 : 0];
        data_mid_8_imag <= _zz_12827[15 : 0];
        data_mid_0_real <= _zz_12835[15 : 0];
        data_mid_0_imag <= _zz_12843[15 : 0];
      end
      if((current_level_value == 3'b100))begin
        data_mid_9_real <= _zz_12860[15 : 0];
        data_mid_9_imag <= _zz_12868[15 : 0];
        data_mid_1_real <= _zz_12876[15 : 0];
        data_mid_1_imag <= _zz_12884[15 : 0];
      end
      if((current_level_value == 3'b100))begin
        data_mid_10_real <= _zz_12901[15 : 0];
        data_mid_10_imag <= _zz_12909[15 : 0];
        data_mid_2_real <= _zz_12917[15 : 0];
        data_mid_2_imag <= _zz_12925[15 : 0];
      end
      if((current_level_value == 3'b100))begin
        data_mid_11_real <= _zz_12942[15 : 0];
        data_mid_11_imag <= _zz_12950[15 : 0];
        data_mid_3_real <= _zz_12958[15 : 0];
        data_mid_3_imag <= _zz_12966[15 : 0];
      end
      if((current_level_value == 3'b100))begin
        data_mid_12_real <= _zz_12983[15 : 0];
        data_mid_12_imag <= _zz_12991[15 : 0];
        data_mid_4_real <= _zz_12999[15 : 0];
        data_mid_4_imag <= _zz_13007[15 : 0];
      end
      if((current_level_value == 3'b100))begin
        data_mid_13_real <= _zz_13024[15 : 0];
        data_mid_13_imag <= _zz_13032[15 : 0];
        data_mid_5_real <= _zz_13040[15 : 0];
        data_mid_5_imag <= _zz_13048[15 : 0];
      end
      if((current_level_value == 3'b100))begin
        data_mid_14_real <= _zz_13065[15 : 0];
        data_mid_14_imag <= _zz_13073[15 : 0];
        data_mid_6_real <= _zz_13081[15 : 0];
        data_mid_6_imag <= _zz_13089[15 : 0];
      end
      if((current_level_value == 3'b100))begin
        data_mid_15_real <= _zz_13106[15 : 0];
        data_mid_15_imag <= _zz_13114[15 : 0];
        data_mid_7_real <= _zz_13122[15 : 0];
        data_mid_7_imag <= _zz_13130[15 : 0];
      end
      if((current_level_value == 3'b100))begin
        data_mid_24_real <= _zz_13147[15 : 0];
        data_mid_24_imag <= _zz_13155[15 : 0];
        data_mid_16_real <= _zz_13163[15 : 0];
        data_mid_16_imag <= _zz_13171[15 : 0];
      end
      if((current_level_value == 3'b100))begin
        data_mid_25_real <= _zz_13188[15 : 0];
        data_mid_25_imag <= _zz_13196[15 : 0];
        data_mid_17_real <= _zz_13204[15 : 0];
        data_mid_17_imag <= _zz_13212[15 : 0];
      end
      if((current_level_value == 3'b100))begin
        data_mid_26_real <= _zz_13229[15 : 0];
        data_mid_26_imag <= _zz_13237[15 : 0];
        data_mid_18_real <= _zz_13245[15 : 0];
        data_mid_18_imag <= _zz_13253[15 : 0];
      end
      if((current_level_value == 3'b100))begin
        data_mid_27_real <= _zz_13270[15 : 0];
        data_mid_27_imag <= _zz_13278[15 : 0];
        data_mid_19_real <= _zz_13286[15 : 0];
        data_mid_19_imag <= _zz_13294[15 : 0];
      end
      if((current_level_value == 3'b100))begin
        data_mid_28_real <= _zz_13311[15 : 0];
        data_mid_28_imag <= _zz_13319[15 : 0];
        data_mid_20_real <= _zz_13327[15 : 0];
        data_mid_20_imag <= _zz_13335[15 : 0];
      end
      if((current_level_value == 3'b100))begin
        data_mid_29_real <= _zz_13352[15 : 0];
        data_mid_29_imag <= _zz_13360[15 : 0];
        data_mid_21_real <= _zz_13368[15 : 0];
        data_mid_21_imag <= _zz_13376[15 : 0];
      end
      if((current_level_value == 3'b100))begin
        data_mid_30_real <= _zz_13393[15 : 0];
        data_mid_30_imag <= _zz_13401[15 : 0];
        data_mid_22_real <= _zz_13409[15 : 0];
        data_mid_22_imag <= _zz_13417[15 : 0];
      end
      if((current_level_value == 3'b100))begin
        data_mid_31_real <= _zz_13434[15 : 0];
        data_mid_31_imag <= _zz_13442[15 : 0];
        data_mid_23_real <= _zz_13450[15 : 0];
        data_mid_23_imag <= _zz_13458[15 : 0];
      end
      if((current_level_value == 3'b100))begin
        data_mid_40_real <= _zz_13475[15 : 0];
        data_mid_40_imag <= _zz_13483[15 : 0];
        data_mid_32_real <= _zz_13491[15 : 0];
        data_mid_32_imag <= _zz_13499[15 : 0];
      end
      if((current_level_value == 3'b100))begin
        data_mid_41_real <= _zz_13516[15 : 0];
        data_mid_41_imag <= _zz_13524[15 : 0];
        data_mid_33_real <= _zz_13532[15 : 0];
        data_mid_33_imag <= _zz_13540[15 : 0];
      end
      if((current_level_value == 3'b100))begin
        data_mid_42_real <= _zz_13557[15 : 0];
        data_mid_42_imag <= _zz_13565[15 : 0];
        data_mid_34_real <= _zz_13573[15 : 0];
        data_mid_34_imag <= _zz_13581[15 : 0];
      end
      if((current_level_value == 3'b100))begin
        data_mid_43_real <= _zz_13598[15 : 0];
        data_mid_43_imag <= _zz_13606[15 : 0];
        data_mid_35_real <= _zz_13614[15 : 0];
        data_mid_35_imag <= _zz_13622[15 : 0];
      end
      if((current_level_value == 3'b100))begin
        data_mid_44_real <= _zz_13639[15 : 0];
        data_mid_44_imag <= _zz_13647[15 : 0];
        data_mid_36_real <= _zz_13655[15 : 0];
        data_mid_36_imag <= _zz_13663[15 : 0];
      end
      if((current_level_value == 3'b100))begin
        data_mid_45_real <= _zz_13680[15 : 0];
        data_mid_45_imag <= _zz_13688[15 : 0];
        data_mid_37_real <= _zz_13696[15 : 0];
        data_mid_37_imag <= _zz_13704[15 : 0];
      end
      if((current_level_value == 3'b100))begin
        data_mid_46_real <= _zz_13721[15 : 0];
        data_mid_46_imag <= _zz_13729[15 : 0];
        data_mid_38_real <= _zz_13737[15 : 0];
        data_mid_38_imag <= _zz_13745[15 : 0];
      end
      if((current_level_value == 3'b100))begin
        data_mid_47_real <= _zz_13762[15 : 0];
        data_mid_47_imag <= _zz_13770[15 : 0];
        data_mid_39_real <= _zz_13778[15 : 0];
        data_mid_39_imag <= _zz_13786[15 : 0];
      end
      if((current_level_value == 3'b100))begin
        data_mid_56_real <= _zz_13803[15 : 0];
        data_mid_56_imag <= _zz_13811[15 : 0];
        data_mid_48_real <= _zz_13819[15 : 0];
        data_mid_48_imag <= _zz_13827[15 : 0];
      end
      if((current_level_value == 3'b100))begin
        data_mid_57_real <= _zz_13844[15 : 0];
        data_mid_57_imag <= _zz_13852[15 : 0];
        data_mid_49_real <= _zz_13860[15 : 0];
        data_mid_49_imag <= _zz_13868[15 : 0];
      end
      if((current_level_value == 3'b100))begin
        data_mid_58_real <= _zz_13885[15 : 0];
        data_mid_58_imag <= _zz_13893[15 : 0];
        data_mid_50_real <= _zz_13901[15 : 0];
        data_mid_50_imag <= _zz_13909[15 : 0];
      end
      if((current_level_value == 3'b100))begin
        data_mid_59_real <= _zz_13926[15 : 0];
        data_mid_59_imag <= _zz_13934[15 : 0];
        data_mid_51_real <= _zz_13942[15 : 0];
        data_mid_51_imag <= _zz_13950[15 : 0];
      end
      if((current_level_value == 3'b100))begin
        data_mid_60_real <= _zz_13967[15 : 0];
        data_mid_60_imag <= _zz_13975[15 : 0];
        data_mid_52_real <= _zz_13983[15 : 0];
        data_mid_52_imag <= _zz_13991[15 : 0];
      end
      if((current_level_value == 3'b100))begin
        data_mid_61_real <= _zz_14008[15 : 0];
        data_mid_61_imag <= _zz_14016[15 : 0];
        data_mid_53_real <= _zz_14024[15 : 0];
        data_mid_53_imag <= _zz_14032[15 : 0];
      end
      if((current_level_value == 3'b100))begin
        data_mid_62_real <= _zz_14049[15 : 0];
        data_mid_62_imag <= _zz_14057[15 : 0];
        data_mid_54_real <= _zz_14065[15 : 0];
        data_mid_54_imag <= _zz_14073[15 : 0];
      end
      if((current_level_value == 3'b100))begin
        data_mid_63_real <= _zz_14090[15 : 0];
        data_mid_63_imag <= _zz_14098[15 : 0];
        data_mid_55_real <= _zz_14106[15 : 0];
        data_mid_55_imag <= _zz_14114[15 : 0];
      end
      if((current_level_value == 3'b100))begin
        data_mid_72_real <= _zz_14131[15 : 0];
        data_mid_72_imag <= _zz_14139[15 : 0];
        data_mid_64_real <= _zz_14147[15 : 0];
        data_mid_64_imag <= _zz_14155[15 : 0];
      end
      if((current_level_value == 3'b100))begin
        data_mid_73_real <= _zz_14172[15 : 0];
        data_mid_73_imag <= _zz_14180[15 : 0];
        data_mid_65_real <= _zz_14188[15 : 0];
        data_mid_65_imag <= _zz_14196[15 : 0];
      end
      if((current_level_value == 3'b100))begin
        data_mid_74_real <= _zz_14213[15 : 0];
        data_mid_74_imag <= _zz_14221[15 : 0];
        data_mid_66_real <= _zz_14229[15 : 0];
        data_mid_66_imag <= _zz_14237[15 : 0];
      end
      if((current_level_value == 3'b100))begin
        data_mid_75_real <= _zz_14254[15 : 0];
        data_mid_75_imag <= _zz_14262[15 : 0];
        data_mid_67_real <= _zz_14270[15 : 0];
        data_mid_67_imag <= _zz_14278[15 : 0];
      end
      if((current_level_value == 3'b100))begin
        data_mid_76_real <= _zz_14295[15 : 0];
        data_mid_76_imag <= _zz_14303[15 : 0];
        data_mid_68_real <= _zz_14311[15 : 0];
        data_mid_68_imag <= _zz_14319[15 : 0];
      end
      if((current_level_value == 3'b100))begin
        data_mid_77_real <= _zz_14336[15 : 0];
        data_mid_77_imag <= _zz_14344[15 : 0];
        data_mid_69_real <= _zz_14352[15 : 0];
        data_mid_69_imag <= _zz_14360[15 : 0];
      end
      if((current_level_value == 3'b100))begin
        data_mid_78_real <= _zz_14377[15 : 0];
        data_mid_78_imag <= _zz_14385[15 : 0];
        data_mid_70_real <= _zz_14393[15 : 0];
        data_mid_70_imag <= _zz_14401[15 : 0];
      end
      if((current_level_value == 3'b100))begin
        data_mid_79_real <= _zz_14418[15 : 0];
        data_mid_79_imag <= _zz_14426[15 : 0];
        data_mid_71_real <= _zz_14434[15 : 0];
        data_mid_71_imag <= _zz_14442[15 : 0];
      end
      if((current_level_value == 3'b100))begin
        data_mid_88_real <= _zz_14459[15 : 0];
        data_mid_88_imag <= _zz_14467[15 : 0];
        data_mid_80_real <= _zz_14475[15 : 0];
        data_mid_80_imag <= _zz_14483[15 : 0];
      end
      if((current_level_value == 3'b100))begin
        data_mid_89_real <= _zz_14500[15 : 0];
        data_mid_89_imag <= _zz_14508[15 : 0];
        data_mid_81_real <= _zz_14516[15 : 0];
        data_mid_81_imag <= _zz_14524[15 : 0];
      end
      if((current_level_value == 3'b100))begin
        data_mid_90_real <= _zz_14541[15 : 0];
        data_mid_90_imag <= _zz_14549[15 : 0];
        data_mid_82_real <= _zz_14557[15 : 0];
        data_mid_82_imag <= _zz_14565[15 : 0];
      end
      if((current_level_value == 3'b100))begin
        data_mid_91_real <= _zz_14582[15 : 0];
        data_mid_91_imag <= _zz_14590[15 : 0];
        data_mid_83_real <= _zz_14598[15 : 0];
        data_mid_83_imag <= _zz_14606[15 : 0];
      end
      if((current_level_value == 3'b100))begin
        data_mid_92_real <= _zz_14623[15 : 0];
        data_mid_92_imag <= _zz_14631[15 : 0];
        data_mid_84_real <= _zz_14639[15 : 0];
        data_mid_84_imag <= _zz_14647[15 : 0];
      end
      if((current_level_value == 3'b100))begin
        data_mid_93_real <= _zz_14664[15 : 0];
        data_mid_93_imag <= _zz_14672[15 : 0];
        data_mid_85_real <= _zz_14680[15 : 0];
        data_mid_85_imag <= _zz_14688[15 : 0];
      end
      if((current_level_value == 3'b100))begin
        data_mid_94_real <= _zz_14705[15 : 0];
        data_mid_94_imag <= _zz_14713[15 : 0];
        data_mid_86_real <= _zz_14721[15 : 0];
        data_mid_86_imag <= _zz_14729[15 : 0];
      end
      if((current_level_value == 3'b100))begin
        data_mid_95_real <= _zz_14746[15 : 0];
        data_mid_95_imag <= _zz_14754[15 : 0];
        data_mid_87_real <= _zz_14762[15 : 0];
        data_mid_87_imag <= _zz_14770[15 : 0];
      end
      if((current_level_value == 3'b100))begin
        data_mid_104_real <= _zz_14787[15 : 0];
        data_mid_104_imag <= _zz_14795[15 : 0];
        data_mid_96_real <= _zz_14803[15 : 0];
        data_mid_96_imag <= _zz_14811[15 : 0];
      end
      if((current_level_value == 3'b100))begin
        data_mid_105_real <= _zz_14828[15 : 0];
        data_mid_105_imag <= _zz_14836[15 : 0];
        data_mid_97_real <= _zz_14844[15 : 0];
        data_mid_97_imag <= _zz_14852[15 : 0];
      end
      if((current_level_value == 3'b100))begin
        data_mid_106_real <= _zz_14869[15 : 0];
        data_mid_106_imag <= _zz_14877[15 : 0];
        data_mid_98_real <= _zz_14885[15 : 0];
        data_mid_98_imag <= _zz_14893[15 : 0];
      end
      if((current_level_value == 3'b100))begin
        data_mid_107_real <= _zz_14910[15 : 0];
        data_mid_107_imag <= _zz_14918[15 : 0];
        data_mid_99_real <= _zz_14926[15 : 0];
        data_mid_99_imag <= _zz_14934[15 : 0];
      end
      if((current_level_value == 3'b100))begin
        data_mid_108_real <= _zz_14951[15 : 0];
        data_mid_108_imag <= _zz_14959[15 : 0];
        data_mid_100_real <= _zz_14967[15 : 0];
        data_mid_100_imag <= _zz_14975[15 : 0];
      end
      if((current_level_value == 3'b100))begin
        data_mid_109_real <= _zz_14992[15 : 0];
        data_mid_109_imag <= _zz_15000[15 : 0];
        data_mid_101_real <= _zz_15008[15 : 0];
        data_mid_101_imag <= _zz_15016[15 : 0];
      end
      if((current_level_value == 3'b100))begin
        data_mid_110_real <= _zz_15033[15 : 0];
        data_mid_110_imag <= _zz_15041[15 : 0];
        data_mid_102_real <= _zz_15049[15 : 0];
        data_mid_102_imag <= _zz_15057[15 : 0];
      end
      if((current_level_value == 3'b100))begin
        data_mid_111_real <= _zz_15074[15 : 0];
        data_mid_111_imag <= _zz_15082[15 : 0];
        data_mid_103_real <= _zz_15090[15 : 0];
        data_mid_103_imag <= _zz_15098[15 : 0];
      end
      if((current_level_value == 3'b100))begin
        data_mid_120_real <= _zz_15115[15 : 0];
        data_mid_120_imag <= _zz_15123[15 : 0];
        data_mid_112_real <= _zz_15131[15 : 0];
        data_mid_112_imag <= _zz_15139[15 : 0];
      end
      if((current_level_value == 3'b100))begin
        data_mid_121_real <= _zz_15156[15 : 0];
        data_mid_121_imag <= _zz_15164[15 : 0];
        data_mid_113_real <= _zz_15172[15 : 0];
        data_mid_113_imag <= _zz_15180[15 : 0];
      end
      if((current_level_value == 3'b100))begin
        data_mid_122_real <= _zz_15197[15 : 0];
        data_mid_122_imag <= _zz_15205[15 : 0];
        data_mid_114_real <= _zz_15213[15 : 0];
        data_mid_114_imag <= _zz_15221[15 : 0];
      end
      if((current_level_value == 3'b100))begin
        data_mid_123_real <= _zz_15238[15 : 0];
        data_mid_123_imag <= _zz_15246[15 : 0];
        data_mid_115_real <= _zz_15254[15 : 0];
        data_mid_115_imag <= _zz_15262[15 : 0];
      end
      if((current_level_value == 3'b100))begin
        data_mid_124_real <= _zz_15279[15 : 0];
        data_mid_124_imag <= _zz_15287[15 : 0];
        data_mid_116_real <= _zz_15295[15 : 0];
        data_mid_116_imag <= _zz_15303[15 : 0];
      end
      if((current_level_value == 3'b100))begin
        data_mid_125_real <= _zz_15320[15 : 0];
        data_mid_125_imag <= _zz_15328[15 : 0];
        data_mid_117_real <= _zz_15336[15 : 0];
        data_mid_117_imag <= _zz_15344[15 : 0];
      end
      if((current_level_value == 3'b100))begin
        data_mid_126_real <= _zz_15361[15 : 0];
        data_mid_126_imag <= _zz_15369[15 : 0];
        data_mid_118_real <= _zz_15377[15 : 0];
        data_mid_118_imag <= _zz_15385[15 : 0];
      end
      if((current_level_value == 3'b100))begin
        data_mid_127_real <= _zz_15402[15 : 0];
        data_mid_127_imag <= _zz_15410[15 : 0];
        data_mid_119_real <= _zz_15418[15 : 0];
        data_mid_119_imag <= _zz_15426[15 : 0];
      end
      if((current_level_value == 3'b101))begin
        data_mid_16_real <= _zz_15443[15 : 0];
        data_mid_16_imag <= _zz_15451[15 : 0];
        data_mid_0_real <= _zz_15459[15 : 0];
        data_mid_0_imag <= _zz_15467[15 : 0];
      end
      if((current_level_value == 3'b101))begin
        data_mid_17_real <= _zz_15484[15 : 0];
        data_mid_17_imag <= _zz_15492[15 : 0];
        data_mid_1_real <= _zz_15500[15 : 0];
        data_mid_1_imag <= _zz_15508[15 : 0];
      end
      if((current_level_value == 3'b101))begin
        data_mid_18_real <= _zz_15525[15 : 0];
        data_mid_18_imag <= _zz_15533[15 : 0];
        data_mid_2_real <= _zz_15541[15 : 0];
        data_mid_2_imag <= _zz_15549[15 : 0];
      end
      if((current_level_value == 3'b101))begin
        data_mid_19_real <= _zz_15566[15 : 0];
        data_mid_19_imag <= _zz_15574[15 : 0];
        data_mid_3_real <= _zz_15582[15 : 0];
        data_mid_3_imag <= _zz_15590[15 : 0];
      end
      if((current_level_value == 3'b101))begin
        data_mid_20_real <= _zz_15607[15 : 0];
        data_mid_20_imag <= _zz_15615[15 : 0];
        data_mid_4_real <= _zz_15623[15 : 0];
        data_mid_4_imag <= _zz_15631[15 : 0];
      end
      if((current_level_value == 3'b101))begin
        data_mid_21_real <= _zz_15648[15 : 0];
        data_mid_21_imag <= _zz_15656[15 : 0];
        data_mid_5_real <= _zz_15664[15 : 0];
        data_mid_5_imag <= _zz_15672[15 : 0];
      end
      if((current_level_value == 3'b101))begin
        data_mid_22_real <= _zz_15689[15 : 0];
        data_mid_22_imag <= _zz_15697[15 : 0];
        data_mid_6_real <= _zz_15705[15 : 0];
        data_mid_6_imag <= _zz_15713[15 : 0];
      end
      if((current_level_value == 3'b101))begin
        data_mid_23_real <= _zz_15730[15 : 0];
        data_mid_23_imag <= _zz_15738[15 : 0];
        data_mid_7_real <= _zz_15746[15 : 0];
        data_mid_7_imag <= _zz_15754[15 : 0];
      end
      if((current_level_value == 3'b101))begin
        data_mid_24_real <= _zz_15771[15 : 0];
        data_mid_24_imag <= _zz_15779[15 : 0];
        data_mid_8_real <= _zz_15787[15 : 0];
        data_mid_8_imag <= _zz_15795[15 : 0];
      end
      if((current_level_value == 3'b101))begin
        data_mid_25_real <= _zz_15812[15 : 0];
        data_mid_25_imag <= _zz_15820[15 : 0];
        data_mid_9_real <= _zz_15828[15 : 0];
        data_mid_9_imag <= _zz_15836[15 : 0];
      end
      if((current_level_value == 3'b101))begin
        data_mid_26_real <= _zz_15853[15 : 0];
        data_mid_26_imag <= _zz_15861[15 : 0];
        data_mid_10_real <= _zz_15869[15 : 0];
        data_mid_10_imag <= _zz_15877[15 : 0];
      end
      if((current_level_value == 3'b101))begin
        data_mid_27_real <= _zz_15894[15 : 0];
        data_mid_27_imag <= _zz_15902[15 : 0];
        data_mid_11_real <= _zz_15910[15 : 0];
        data_mid_11_imag <= _zz_15918[15 : 0];
      end
      if((current_level_value == 3'b101))begin
        data_mid_28_real <= _zz_15935[15 : 0];
        data_mid_28_imag <= _zz_15943[15 : 0];
        data_mid_12_real <= _zz_15951[15 : 0];
        data_mid_12_imag <= _zz_15959[15 : 0];
      end
      if((current_level_value == 3'b101))begin
        data_mid_29_real <= _zz_15976[15 : 0];
        data_mid_29_imag <= _zz_15984[15 : 0];
        data_mid_13_real <= _zz_15992[15 : 0];
        data_mid_13_imag <= _zz_16000[15 : 0];
      end
      if((current_level_value == 3'b101))begin
        data_mid_30_real <= _zz_16017[15 : 0];
        data_mid_30_imag <= _zz_16025[15 : 0];
        data_mid_14_real <= _zz_16033[15 : 0];
        data_mid_14_imag <= _zz_16041[15 : 0];
      end
      if((current_level_value == 3'b101))begin
        data_mid_31_real <= _zz_16058[15 : 0];
        data_mid_31_imag <= _zz_16066[15 : 0];
        data_mid_15_real <= _zz_16074[15 : 0];
        data_mid_15_imag <= _zz_16082[15 : 0];
      end
      if((current_level_value == 3'b101))begin
        data_mid_48_real <= _zz_16099[15 : 0];
        data_mid_48_imag <= _zz_16107[15 : 0];
        data_mid_32_real <= _zz_16115[15 : 0];
        data_mid_32_imag <= _zz_16123[15 : 0];
      end
      if((current_level_value == 3'b101))begin
        data_mid_49_real <= _zz_16140[15 : 0];
        data_mid_49_imag <= _zz_16148[15 : 0];
        data_mid_33_real <= _zz_16156[15 : 0];
        data_mid_33_imag <= _zz_16164[15 : 0];
      end
      if((current_level_value == 3'b101))begin
        data_mid_50_real <= _zz_16181[15 : 0];
        data_mid_50_imag <= _zz_16189[15 : 0];
        data_mid_34_real <= _zz_16197[15 : 0];
        data_mid_34_imag <= _zz_16205[15 : 0];
      end
      if((current_level_value == 3'b101))begin
        data_mid_51_real <= _zz_16222[15 : 0];
        data_mid_51_imag <= _zz_16230[15 : 0];
        data_mid_35_real <= _zz_16238[15 : 0];
        data_mid_35_imag <= _zz_16246[15 : 0];
      end
      if((current_level_value == 3'b101))begin
        data_mid_52_real <= _zz_16263[15 : 0];
        data_mid_52_imag <= _zz_16271[15 : 0];
        data_mid_36_real <= _zz_16279[15 : 0];
        data_mid_36_imag <= _zz_16287[15 : 0];
      end
      if((current_level_value == 3'b101))begin
        data_mid_53_real <= _zz_16304[15 : 0];
        data_mid_53_imag <= _zz_16312[15 : 0];
        data_mid_37_real <= _zz_16320[15 : 0];
        data_mid_37_imag <= _zz_16328[15 : 0];
      end
      if((current_level_value == 3'b101))begin
        data_mid_54_real <= _zz_16345[15 : 0];
        data_mid_54_imag <= _zz_16353[15 : 0];
        data_mid_38_real <= _zz_16361[15 : 0];
        data_mid_38_imag <= _zz_16369[15 : 0];
      end
      if((current_level_value == 3'b101))begin
        data_mid_55_real <= _zz_16386[15 : 0];
        data_mid_55_imag <= _zz_16394[15 : 0];
        data_mid_39_real <= _zz_16402[15 : 0];
        data_mid_39_imag <= _zz_16410[15 : 0];
      end
      if((current_level_value == 3'b101))begin
        data_mid_56_real <= _zz_16427[15 : 0];
        data_mid_56_imag <= _zz_16435[15 : 0];
        data_mid_40_real <= _zz_16443[15 : 0];
        data_mid_40_imag <= _zz_16451[15 : 0];
      end
      if((current_level_value == 3'b101))begin
        data_mid_57_real <= _zz_16468[15 : 0];
        data_mid_57_imag <= _zz_16476[15 : 0];
        data_mid_41_real <= _zz_16484[15 : 0];
        data_mid_41_imag <= _zz_16492[15 : 0];
      end
      if((current_level_value == 3'b101))begin
        data_mid_58_real <= _zz_16509[15 : 0];
        data_mid_58_imag <= _zz_16517[15 : 0];
        data_mid_42_real <= _zz_16525[15 : 0];
        data_mid_42_imag <= _zz_16533[15 : 0];
      end
      if((current_level_value == 3'b101))begin
        data_mid_59_real <= _zz_16550[15 : 0];
        data_mid_59_imag <= _zz_16558[15 : 0];
        data_mid_43_real <= _zz_16566[15 : 0];
        data_mid_43_imag <= _zz_16574[15 : 0];
      end
      if((current_level_value == 3'b101))begin
        data_mid_60_real <= _zz_16591[15 : 0];
        data_mid_60_imag <= _zz_16599[15 : 0];
        data_mid_44_real <= _zz_16607[15 : 0];
        data_mid_44_imag <= _zz_16615[15 : 0];
      end
      if((current_level_value == 3'b101))begin
        data_mid_61_real <= _zz_16632[15 : 0];
        data_mid_61_imag <= _zz_16640[15 : 0];
        data_mid_45_real <= _zz_16648[15 : 0];
        data_mid_45_imag <= _zz_16656[15 : 0];
      end
      if((current_level_value == 3'b101))begin
        data_mid_62_real <= _zz_16673[15 : 0];
        data_mid_62_imag <= _zz_16681[15 : 0];
        data_mid_46_real <= _zz_16689[15 : 0];
        data_mid_46_imag <= _zz_16697[15 : 0];
      end
      if((current_level_value == 3'b101))begin
        data_mid_63_real <= _zz_16714[15 : 0];
        data_mid_63_imag <= _zz_16722[15 : 0];
        data_mid_47_real <= _zz_16730[15 : 0];
        data_mid_47_imag <= _zz_16738[15 : 0];
      end
      if((current_level_value == 3'b101))begin
        data_mid_80_real <= _zz_16755[15 : 0];
        data_mid_80_imag <= _zz_16763[15 : 0];
        data_mid_64_real <= _zz_16771[15 : 0];
        data_mid_64_imag <= _zz_16779[15 : 0];
      end
      if((current_level_value == 3'b101))begin
        data_mid_81_real <= _zz_16796[15 : 0];
        data_mid_81_imag <= _zz_16804[15 : 0];
        data_mid_65_real <= _zz_16812[15 : 0];
        data_mid_65_imag <= _zz_16820[15 : 0];
      end
      if((current_level_value == 3'b101))begin
        data_mid_82_real <= _zz_16837[15 : 0];
        data_mid_82_imag <= _zz_16845[15 : 0];
        data_mid_66_real <= _zz_16853[15 : 0];
        data_mid_66_imag <= _zz_16861[15 : 0];
      end
      if((current_level_value == 3'b101))begin
        data_mid_83_real <= _zz_16878[15 : 0];
        data_mid_83_imag <= _zz_16886[15 : 0];
        data_mid_67_real <= _zz_16894[15 : 0];
        data_mid_67_imag <= _zz_16902[15 : 0];
      end
      if((current_level_value == 3'b101))begin
        data_mid_84_real <= _zz_16919[15 : 0];
        data_mid_84_imag <= _zz_16927[15 : 0];
        data_mid_68_real <= _zz_16935[15 : 0];
        data_mid_68_imag <= _zz_16943[15 : 0];
      end
      if((current_level_value == 3'b101))begin
        data_mid_85_real <= _zz_16960[15 : 0];
        data_mid_85_imag <= _zz_16968[15 : 0];
        data_mid_69_real <= _zz_16976[15 : 0];
        data_mid_69_imag <= _zz_16984[15 : 0];
      end
      if((current_level_value == 3'b101))begin
        data_mid_86_real <= _zz_17001[15 : 0];
        data_mid_86_imag <= _zz_17009[15 : 0];
        data_mid_70_real <= _zz_17017[15 : 0];
        data_mid_70_imag <= _zz_17025[15 : 0];
      end
      if((current_level_value == 3'b101))begin
        data_mid_87_real <= _zz_17042[15 : 0];
        data_mid_87_imag <= _zz_17050[15 : 0];
        data_mid_71_real <= _zz_17058[15 : 0];
        data_mid_71_imag <= _zz_17066[15 : 0];
      end
      if((current_level_value == 3'b101))begin
        data_mid_88_real <= _zz_17083[15 : 0];
        data_mid_88_imag <= _zz_17091[15 : 0];
        data_mid_72_real <= _zz_17099[15 : 0];
        data_mid_72_imag <= _zz_17107[15 : 0];
      end
      if((current_level_value == 3'b101))begin
        data_mid_89_real <= _zz_17124[15 : 0];
        data_mid_89_imag <= _zz_17132[15 : 0];
        data_mid_73_real <= _zz_17140[15 : 0];
        data_mid_73_imag <= _zz_17148[15 : 0];
      end
      if((current_level_value == 3'b101))begin
        data_mid_90_real <= _zz_17165[15 : 0];
        data_mid_90_imag <= _zz_17173[15 : 0];
        data_mid_74_real <= _zz_17181[15 : 0];
        data_mid_74_imag <= _zz_17189[15 : 0];
      end
      if((current_level_value == 3'b101))begin
        data_mid_91_real <= _zz_17206[15 : 0];
        data_mid_91_imag <= _zz_17214[15 : 0];
        data_mid_75_real <= _zz_17222[15 : 0];
        data_mid_75_imag <= _zz_17230[15 : 0];
      end
      if((current_level_value == 3'b101))begin
        data_mid_92_real <= _zz_17247[15 : 0];
        data_mid_92_imag <= _zz_17255[15 : 0];
        data_mid_76_real <= _zz_17263[15 : 0];
        data_mid_76_imag <= _zz_17271[15 : 0];
      end
      if((current_level_value == 3'b101))begin
        data_mid_93_real <= _zz_17288[15 : 0];
        data_mid_93_imag <= _zz_17296[15 : 0];
        data_mid_77_real <= _zz_17304[15 : 0];
        data_mid_77_imag <= _zz_17312[15 : 0];
      end
      if((current_level_value == 3'b101))begin
        data_mid_94_real <= _zz_17329[15 : 0];
        data_mid_94_imag <= _zz_17337[15 : 0];
        data_mid_78_real <= _zz_17345[15 : 0];
        data_mid_78_imag <= _zz_17353[15 : 0];
      end
      if((current_level_value == 3'b101))begin
        data_mid_95_real <= _zz_17370[15 : 0];
        data_mid_95_imag <= _zz_17378[15 : 0];
        data_mid_79_real <= _zz_17386[15 : 0];
        data_mid_79_imag <= _zz_17394[15 : 0];
      end
      if((current_level_value == 3'b101))begin
        data_mid_112_real <= _zz_17411[15 : 0];
        data_mid_112_imag <= _zz_17419[15 : 0];
        data_mid_96_real <= _zz_17427[15 : 0];
        data_mid_96_imag <= _zz_17435[15 : 0];
      end
      if((current_level_value == 3'b101))begin
        data_mid_113_real <= _zz_17452[15 : 0];
        data_mid_113_imag <= _zz_17460[15 : 0];
        data_mid_97_real <= _zz_17468[15 : 0];
        data_mid_97_imag <= _zz_17476[15 : 0];
      end
      if((current_level_value == 3'b101))begin
        data_mid_114_real <= _zz_17493[15 : 0];
        data_mid_114_imag <= _zz_17501[15 : 0];
        data_mid_98_real <= _zz_17509[15 : 0];
        data_mid_98_imag <= _zz_17517[15 : 0];
      end
      if((current_level_value == 3'b101))begin
        data_mid_115_real <= _zz_17534[15 : 0];
        data_mid_115_imag <= _zz_17542[15 : 0];
        data_mid_99_real <= _zz_17550[15 : 0];
        data_mid_99_imag <= _zz_17558[15 : 0];
      end
      if((current_level_value == 3'b101))begin
        data_mid_116_real <= _zz_17575[15 : 0];
        data_mid_116_imag <= _zz_17583[15 : 0];
        data_mid_100_real <= _zz_17591[15 : 0];
        data_mid_100_imag <= _zz_17599[15 : 0];
      end
      if((current_level_value == 3'b101))begin
        data_mid_117_real <= _zz_17616[15 : 0];
        data_mid_117_imag <= _zz_17624[15 : 0];
        data_mid_101_real <= _zz_17632[15 : 0];
        data_mid_101_imag <= _zz_17640[15 : 0];
      end
      if((current_level_value == 3'b101))begin
        data_mid_118_real <= _zz_17657[15 : 0];
        data_mid_118_imag <= _zz_17665[15 : 0];
        data_mid_102_real <= _zz_17673[15 : 0];
        data_mid_102_imag <= _zz_17681[15 : 0];
      end
      if((current_level_value == 3'b101))begin
        data_mid_119_real <= _zz_17698[15 : 0];
        data_mid_119_imag <= _zz_17706[15 : 0];
        data_mid_103_real <= _zz_17714[15 : 0];
        data_mid_103_imag <= _zz_17722[15 : 0];
      end
      if((current_level_value == 3'b101))begin
        data_mid_120_real <= _zz_17739[15 : 0];
        data_mid_120_imag <= _zz_17747[15 : 0];
        data_mid_104_real <= _zz_17755[15 : 0];
        data_mid_104_imag <= _zz_17763[15 : 0];
      end
      if((current_level_value == 3'b101))begin
        data_mid_121_real <= _zz_17780[15 : 0];
        data_mid_121_imag <= _zz_17788[15 : 0];
        data_mid_105_real <= _zz_17796[15 : 0];
        data_mid_105_imag <= _zz_17804[15 : 0];
      end
      if((current_level_value == 3'b101))begin
        data_mid_122_real <= _zz_17821[15 : 0];
        data_mid_122_imag <= _zz_17829[15 : 0];
        data_mid_106_real <= _zz_17837[15 : 0];
        data_mid_106_imag <= _zz_17845[15 : 0];
      end
      if((current_level_value == 3'b101))begin
        data_mid_123_real <= _zz_17862[15 : 0];
        data_mid_123_imag <= _zz_17870[15 : 0];
        data_mid_107_real <= _zz_17878[15 : 0];
        data_mid_107_imag <= _zz_17886[15 : 0];
      end
      if((current_level_value == 3'b101))begin
        data_mid_124_real <= _zz_17903[15 : 0];
        data_mid_124_imag <= _zz_17911[15 : 0];
        data_mid_108_real <= _zz_17919[15 : 0];
        data_mid_108_imag <= _zz_17927[15 : 0];
      end
      if((current_level_value == 3'b101))begin
        data_mid_125_real <= _zz_17944[15 : 0];
        data_mid_125_imag <= _zz_17952[15 : 0];
        data_mid_109_real <= _zz_17960[15 : 0];
        data_mid_109_imag <= _zz_17968[15 : 0];
      end
      if((current_level_value == 3'b101))begin
        data_mid_126_real <= _zz_17985[15 : 0];
        data_mid_126_imag <= _zz_17993[15 : 0];
        data_mid_110_real <= _zz_18001[15 : 0];
        data_mid_110_imag <= _zz_18009[15 : 0];
      end
      if((current_level_value == 3'b101))begin
        data_mid_127_real <= _zz_18026[15 : 0];
        data_mid_127_imag <= _zz_18034[15 : 0];
        data_mid_111_real <= _zz_18042[15 : 0];
        data_mid_111_imag <= _zz_18050[15 : 0];
      end
      if((current_level_value == 3'b110))begin
        data_mid_32_real <= _zz_18067[15 : 0];
        data_mid_32_imag <= _zz_18075[15 : 0];
        data_mid_0_real <= _zz_18083[15 : 0];
        data_mid_0_imag <= _zz_18091[15 : 0];
      end
      if((current_level_value == 3'b110))begin
        data_mid_33_real <= _zz_18108[15 : 0];
        data_mid_33_imag <= _zz_18116[15 : 0];
        data_mid_1_real <= _zz_18124[15 : 0];
        data_mid_1_imag <= _zz_18132[15 : 0];
      end
      if((current_level_value == 3'b110))begin
        data_mid_34_real <= _zz_18149[15 : 0];
        data_mid_34_imag <= _zz_18157[15 : 0];
        data_mid_2_real <= _zz_18165[15 : 0];
        data_mid_2_imag <= _zz_18173[15 : 0];
      end
      if((current_level_value == 3'b110))begin
        data_mid_35_real <= _zz_18190[15 : 0];
        data_mid_35_imag <= _zz_18198[15 : 0];
        data_mid_3_real <= _zz_18206[15 : 0];
        data_mid_3_imag <= _zz_18214[15 : 0];
      end
      if((current_level_value == 3'b110))begin
        data_mid_36_real <= _zz_18231[15 : 0];
        data_mid_36_imag <= _zz_18239[15 : 0];
        data_mid_4_real <= _zz_18247[15 : 0];
        data_mid_4_imag <= _zz_18255[15 : 0];
      end
      if((current_level_value == 3'b110))begin
        data_mid_37_real <= _zz_18272[15 : 0];
        data_mid_37_imag <= _zz_18280[15 : 0];
        data_mid_5_real <= _zz_18288[15 : 0];
        data_mid_5_imag <= _zz_18296[15 : 0];
      end
      if((current_level_value == 3'b110))begin
        data_mid_38_real <= _zz_18313[15 : 0];
        data_mid_38_imag <= _zz_18321[15 : 0];
        data_mid_6_real <= _zz_18329[15 : 0];
        data_mid_6_imag <= _zz_18337[15 : 0];
      end
      if((current_level_value == 3'b110))begin
        data_mid_39_real <= _zz_18354[15 : 0];
        data_mid_39_imag <= _zz_18362[15 : 0];
        data_mid_7_real <= _zz_18370[15 : 0];
        data_mid_7_imag <= _zz_18378[15 : 0];
      end
      if((current_level_value == 3'b110))begin
        data_mid_40_real <= _zz_18395[15 : 0];
        data_mid_40_imag <= _zz_18403[15 : 0];
        data_mid_8_real <= _zz_18411[15 : 0];
        data_mid_8_imag <= _zz_18419[15 : 0];
      end
      if((current_level_value == 3'b110))begin
        data_mid_41_real <= _zz_18436[15 : 0];
        data_mid_41_imag <= _zz_18444[15 : 0];
        data_mid_9_real <= _zz_18452[15 : 0];
        data_mid_9_imag <= _zz_18460[15 : 0];
      end
      if((current_level_value == 3'b110))begin
        data_mid_42_real <= _zz_18477[15 : 0];
        data_mid_42_imag <= _zz_18485[15 : 0];
        data_mid_10_real <= _zz_18493[15 : 0];
        data_mid_10_imag <= _zz_18501[15 : 0];
      end
      if((current_level_value == 3'b110))begin
        data_mid_43_real <= _zz_18518[15 : 0];
        data_mid_43_imag <= _zz_18526[15 : 0];
        data_mid_11_real <= _zz_18534[15 : 0];
        data_mid_11_imag <= _zz_18542[15 : 0];
      end
      if((current_level_value == 3'b110))begin
        data_mid_44_real <= _zz_18559[15 : 0];
        data_mid_44_imag <= _zz_18567[15 : 0];
        data_mid_12_real <= _zz_18575[15 : 0];
        data_mid_12_imag <= _zz_18583[15 : 0];
      end
      if((current_level_value == 3'b110))begin
        data_mid_45_real <= _zz_18600[15 : 0];
        data_mid_45_imag <= _zz_18608[15 : 0];
        data_mid_13_real <= _zz_18616[15 : 0];
        data_mid_13_imag <= _zz_18624[15 : 0];
      end
      if((current_level_value == 3'b110))begin
        data_mid_46_real <= _zz_18641[15 : 0];
        data_mid_46_imag <= _zz_18649[15 : 0];
        data_mid_14_real <= _zz_18657[15 : 0];
        data_mid_14_imag <= _zz_18665[15 : 0];
      end
      if((current_level_value == 3'b110))begin
        data_mid_47_real <= _zz_18682[15 : 0];
        data_mid_47_imag <= _zz_18690[15 : 0];
        data_mid_15_real <= _zz_18698[15 : 0];
        data_mid_15_imag <= _zz_18706[15 : 0];
      end
      if((current_level_value == 3'b110))begin
        data_mid_48_real <= _zz_18723[15 : 0];
        data_mid_48_imag <= _zz_18731[15 : 0];
        data_mid_16_real <= _zz_18739[15 : 0];
        data_mid_16_imag <= _zz_18747[15 : 0];
      end
      if((current_level_value == 3'b110))begin
        data_mid_49_real <= _zz_18764[15 : 0];
        data_mid_49_imag <= _zz_18772[15 : 0];
        data_mid_17_real <= _zz_18780[15 : 0];
        data_mid_17_imag <= _zz_18788[15 : 0];
      end
      if((current_level_value == 3'b110))begin
        data_mid_50_real <= _zz_18805[15 : 0];
        data_mid_50_imag <= _zz_18813[15 : 0];
        data_mid_18_real <= _zz_18821[15 : 0];
        data_mid_18_imag <= _zz_18829[15 : 0];
      end
      if((current_level_value == 3'b110))begin
        data_mid_51_real <= _zz_18846[15 : 0];
        data_mid_51_imag <= _zz_18854[15 : 0];
        data_mid_19_real <= _zz_18862[15 : 0];
        data_mid_19_imag <= _zz_18870[15 : 0];
      end
      if((current_level_value == 3'b110))begin
        data_mid_52_real <= _zz_18887[15 : 0];
        data_mid_52_imag <= _zz_18895[15 : 0];
        data_mid_20_real <= _zz_18903[15 : 0];
        data_mid_20_imag <= _zz_18911[15 : 0];
      end
      if((current_level_value == 3'b110))begin
        data_mid_53_real <= _zz_18928[15 : 0];
        data_mid_53_imag <= _zz_18936[15 : 0];
        data_mid_21_real <= _zz_18944[15 : 0];
        data_mid_21_imag <= _zz_18952[15 : 0];
      end
      if((current_level_value == 3'b110))begin
        data_mid_54_real <= _zz_18969[15 : 0];
        data_mid_54_imag <= _zz_18977[15 : 0];
        data_mid_22_real <= _zz_18985[15 : 0];
        data_mid_22_imag <= _zz_18993[15 : 0];
      end
      if((current_level_value == 3'b110))begin
        data_mid_55_real <= _zz_19010[15 : 0];
        data_mid_55_imag <= _zz_19018[15 : 0];
        data_mid_23_real <= _zz_19026[15 : 0];
        data_mid_23_imag <= _zz_19034[15 : 0];
      end
      if((current_level_value == 3'b110))begin
        data_mid_56_real <= _zz_19051[15 : 0];
        data_mid_56_imag <= _zz_19059[15 : 0];
        data_mid_24_real <= _zz_19067[15 : 0];
        data_mid_24_imag <= _zz_19075[15 : 0];
      end
      if((current_level_value == 3'b110))begin
        data_mid_57_real <= _zz_19092[15 : 0];
        data_mid_57_imag <= _zz_19100[15 : 0];
        data_mid_25_real <= _zz_19108[15 : 0];
        data_mid_25_imag <= _zz_19116[15 : 0];
      end
      if((current_level_value == 3'b110))begin
        data_mid_58_real <= _zz_19133[15 : 0];
        data_mid_58_imag <= _zz_19141[15 : 0];
        data_mid_26_real <= _zz_19149[15 : 0];
        data_mid_26_imag <= _zz_19157[15 : 0];
      end
      if((current_level_value == 3'b110))begin
        data_mid_59_real <= _zz_19174[15 : 0];
        data_mid_59_imag <= _zz_19182[15 : 0];
        data_mid_27_real <= _zz_19190[15 : 0];
        data_mid_27_imag <= _zz_19198[15 : 0];
      end
      if((current_level_value == 3'b110))begin
        data_mid_60_real <= _zz_19215[15 : 0];
        data_mid_60_imag <= _zz_19223[15 : 0];
        data_mid_28_real <= _zz_19231[15 : 0];
        data_mid_28_imag <= _zz_19239[15 : 0];
      end
      if((current_level_value == 3'b110))begin
        data_mid_61_real <= _zz_19256[15 : 0];
        data_mid_61_imag <= _zz_19264[15 : 0];
        data_mid_29_real <= _zz_19272[15 : 0];
        data_mid_29_imag <= _zz_19280[15 : 0];
      end
      if((current_level_value == 3'b110))begin
        data_mid_62_real <= _zz_19297[15 : 0];
        data_mid_62_imag <= _zz_19305[15 : 0];
        data_mid_30_real <= _zz_19313[15 : 0];
        data_mid_30_imag <= _zz_19321[15 : 0];
      end
      if((current_level_value == 3'b110))begin
        data_mid_63_real <= _zz_19338[15 : 0];
        data_mid_63_imag <= _zz_19346[15 : 0];
        data_mid_31_real <= _zz_19354[15 : 0];
        data_mid_31_imag <= _zz_19362[15 : 0];
      end
      if((current_level_value == 3'b110))begin
        data_mid_96_real <= _zz_19379[15 : 0];
        data_mid_96_imag <= _zz_19387[15 : 0];
        data_mid_64_real <= _zz_19395[15 : 0];
        data_mid_64_imag <= _zz_19403[15 : 0];
      end
      if((current_level_value == 3'b110))begin
        data_mid_97_real <= _zz_19420[15 : 0];
        data_mid_97_imag <= _zz_19428[15 : 0];
        data_mid_65_real <= _zz_19436[15 : 0];
        data_mid_65_imag <= _zz_19444[15 : 0];
      end
      if((current_level_value == 3'b110))begin
        data_mid_98_real <= _zz_19461[15 : 0];
        data_mid_98_imag <= _zz_19469[15 : 0];
        data_mid_66_real <= _zz_19477[15 : 0];
        data_mid_66_imag <= _zz_19485[15 : 0];
      end
      if((current_level_value == 3'b110))begin
        data_mid_99_real <= _zz_19502[15 : 0];
        data_mid_99_imag <= _zz_19510[15 : 0];
        data_mid_67_real <= _zz_19518[15 : 0];
        data_mid_67_imag <= _zz_19526[15 : 0];
      end
      if((current_level_value == 3'b110))begin
        data_mid_100_real <= _zz_19543[15 : 0];
        data_mid_100_imag <= _zz_19551[15 : 0];
        data_mid_68_real <= _zz_19559[15 : 0];
        data_mid_68_imag <= _zz_19567[15 : 0];
      end
      if((current_level_value == 3'b110))begin
        data_mid_101_real <= _zz_19584[15 : 0];
        data_mid_101_imag <= _zz_19592[15 : 0];
        data_mid_69_real <= _zz_19600[15 : 0];
        data_mid_69_imag <= _zz_19608[15 : 0];
      end
      if((current_level_value == 3'b110))begin
        data_mid_102_real <= _zz_19625[15 : 0];
        data_mid_102_imag <= _zz_19633[15 : 0];
        data_mid_70_real <= _zz_19641[15 : 0];
        data_mid_70_imag <= _zz_19649[15 : 0];
      end
      if((current_level_value == 3'b110))begin
        data_mid_103_real <= _zz_19666[15 : 0];
        data_mid_103_imag <= _zz_19674[15 : 0];
        data_mid_71_real <= _zz_19682[15 : 0];
        data_mid_71_imag <= _zz_19690[15 : 0];
      end
      if((current_level_value == 3'b110))begin
        data_mid_104_real <= _zz_19707[15 : 0];
        data_mid_104_imag <= _zz_19715[15 : 0];
        data_mid_72_real <= _zz_19723[15 : 0];
        data_mid_72_imag <= _zz_19731[15 : 0];
      end
      if((current_level_value == 3'b110))begin
        data_mid_105_real <= _zz_19748[15 : 0];
        data_mid_105_imag <= _zz_19756[15 : 0];
        data_mid_73_real <= _zz_19764[15 : 0];
        data_mid_73_imag <= _zz_19772[15 : 0];
      end
      if((current_level_value == 3'b110))begin
        data_mid_106_real <= _zz_19789[15 : 0];
        data_mid_106_imag <= _zz_19797[15 : 0];
        data_mid_74_real <= _zz_19805[15 : 0];
        data_mid_74_imag <= _zz_19813[15 : 0];
      end
      if((current_level_value == 3'b110))begin
        data_mid_107_real <= _zz_19830[15 : 0];
        data_mid_107_imag <= _zz_19838[15 : 0];
        data_mid_75_real <= _zz_19846[15 : 0];
        data_mid_75_imag <= _zz_19854[15 : 0];
      end
      if((current_level_value == 3'b110))begin
        data_mid_108_real <= _zz_19871[15 : 0];
        data_mid_108_imag <= _zz_19879[15 : 0];
        data_mid_76_real <= _zz_19887[15 : 0];
        data_mid_76_imag <= _zz_19895[15 : 0];
      end
      if((current_level_value == 3'b110))begin
        data_mid_109_real <= _zz_19912[15 : 0];
        data_mid_109_imag <= _zz_19920[15 : 0];
        data_mid_77_real <= _zz_19928[15 : 0];
        data_mid_77_imag <= _zz_19936[15 : 0];
      end
      if((current_level_value == 3'b110))begin
        data_mid_110_real <= _zz_19953[15 : 0];
        data_mid_110_imag <= _zz_19961[15 : 0];
        data_mid_78_real <= _zz_19969[15 : 0];
        data_mid_78_imag <= _zz_19977[15 : 0];
      end
      if((current_level_value == 3'b110))begin
        data_mid_111_real <= _zz_19994[15 : 0];
        data_mid_111_imag <= _zz_20002[15 : 0];
        data_mid_79_real <= _zz_20010[15 : 0];
        data_mid_79_imag <= _zz_20018[15 : 0];
      end
      if((current_level_value == 3'b110))begin
        data_mid_112_real <= _zz_20035[15 : 0];
        data_mid_112_imag <= _zz_20043[15 : 0];
        data_mid_80_real <= _zz_20051[15 : 0];
        data_mid_80_imag <= _zz_20059[15 : 0];
      end
      if((current_level_value == 3'b110))begin
        data_mid_113_real <= _zz_20076[15 : 0];
        data_mid_113_imag <= _zz_20084[15 : 0];
        data_mid_81_real <= _zz_20092[15 : 0];
        data_mid_81_imag <= _zz_20100[15 : 0];
      end
      if((current_level_value == 3'b110))begin
        data_mid_114_real <= _zz_20117[15 : 0];
        data_mid_114_imag <= _zz_20125[15 : 0];
        data_mid_82_real <= _zz_20133[15 : 0];
        data_mid_82_imag <= _zz_20141[15 : 0];
      end
      if((current_level_value == 3'b110))begin
        data_mid_115_real <= _zz_20158[15 : 0];
        data_mid_115_imag <= _zz_20166[15 : 0];
        data_mid_83_real <= _zz_20174[15 : 0];
        data_mid_83_imag <= _zz_20182[15 : 0];
      end
      if((current_level_value == 3'b110))begin
        data_mid_116_real <= _zz_20199[15 : 0];
        data_mid_116_imag <= _zz_20207[15 : 0];
        data_mid_84_real <= _zz_20215[15 : 0];
        data_mid_84_imag <= _zz_20223[15 : 0];
      end
      if((current_level_value == 3'b110))begin
        data_mid_117_real <= _zz_20240[15 : 0];
        data_mid_117_imag <= _zz_20248[15 : 0];
        data_mid_85_real <= _zz_20256[15 : 0];
        data_mid_85_imag <= _zz_20264[15 : 0];
      end
      if((current_level_value == 3'b110))begin
        data_mid_118_real <= _zz_20281[15 : 0];
        data_mid_118_imag <= _zz_20289[15 : 0];
        data_mid_86_real <= _zz_20297[15 : 0];
        data_mid_86_imag <= _zz_20305[15 : 0];
      end
      if((current_level_value == 3'b110))begin
        data_mid_119_real <= _zz_20322[15 : 0];
        data_mid_119_imag <= _zz_20330[15 : 0];
        data_mid_87_real <= _zz_20338[15 : 0];
        data_mid_87_imag <= _zz_20346[15 : 0];
      end
      if((current_level_value == 3'b110))begin
        data_mid_120_real <= _zz_20363[15 : 0];
        data_mid_120_imag <= _zz_20371[15 : 0];
        data_mid_88_real <= _zz_20379[15 : 0];
        data_mid_88_imag <= _zz_20387[15 : 0];
      end
      if((current_level_value == 3'b110))begin
        data_mid_121_real <= _zz_20404[15 : 0];
        data_mid_121_imag <= _zz_20412[15 : 0];
        data_mid_89_real <= _zz_20420[15 : 0];
        data_mid_89_imag <= _zz_20428[15 : 0];
      end
      if((current_level_value == 3'b110))begin
        data_mid_122_real <= _zz_20445[15 : 0];
        data_mid_122_imag <= _zz_20453[15 : 0];
        data_mid_90_real <= _zz_20461[15 : 0];
        data_mid_90_imag <= _zz_20469[15 : 0];
      end
      if((current_level_value == 3'b110))begin
        data_mid_123_real <= _zz_20486[15 : 0];
        data_mid_123_imag <= _zz_20494[15 : 0];
        data_mid_91_real <= _zz_20502[15 : 0];
        data_mid_91_imag <= _zz_20510[15 : 0];
      end
      if((current_level_value == 3'b110))begin
        data_mid_124_real <= _zz_20527[15 : 0];
        data_mid_124_imag <= _zz_20535[15 : 0];
        data_mid_92_real <= _zz_20543[15 : 0];
        data_mid_92_imag <= _zz_20551[15 : 0];
      end
      if((current_level_value == 3'b110))begin
        data_mid_125_real <= _zz_20568[15 : 0];
        data_mid_125_imag <= _zz_20576[15 : 0];
        data_mid_93_real <= _zz_20584[15 : 0];
        data_mid_93_imag <= _zz_20592[15 : 0];
      end
      if((current_level_value == 3'b110))begin
        data_mid_126_real <= _zz_20609[15 : 0];
        data_mid_126_imag <= _zz_20617[15 : 0];
        data_mid_94_real <= _zz_20625[15 : 0];
        data_mid_94_imag <= _zz_20633[15 : 0];
      end
      if((current_level_value == 3'b110))begin
        data_mid_127_real <= _zz_20650[15 : 0];
        data_mid_127_imag <= _zz_20658[15 : 0];
        data_mid_95_real <= _zz_20666[15 : 0];
        data_mid_95_imag <= _zz_20674[15 : 0];
      end
      if((current_level_value == 3'b111))begin
        data_mid_64_real <= _zz_20691[15 : 0];
        data_mid_64_imag <= _zz_20699[15 : 0];
        data_mid_0_real <= _zz_20707[15 : 0];
        data_mid_0_imag <= _zz_20715[15 : 0];
      end
      if((current_level_value == 3'b111))begin
        data_mid_65_real <= _zz_20732[15 : 0];
        data_mid_65_imag <= _zz_20740[15 : 0];
        data_mid_1_real <= _zz_20748[15 : 0];
        data_mid_1_imag <= _zz_20756[15 : 0];
      end
      if((current_level_value == 3'b111))begin
        data_mid_66_real <= _zz_20773[15 : 0];
        data_mid_66_imag <= _zz_20781[15 : 0];
        data_mid_2_real <= _zz_20789[15 : 0];
        data_mid_2_imag <= _zz_20797[15 : 0];
      end
      if((current_level_value == 3'b111))begin
        data_mid_67_real <= _zz_20814[15 : 0];
        data_mid_67_imag <= _zz_20822[15 : 0];
        data_mid_3_real <= _zz_20830[15 : 0];
        data_mid_3_imag <= _zz_20838[15 : 0];
      end
      if((current_level_value == 3'b111))begin
        data_mid_68_real <= _zz_20855[15 : 0];
        data_mid_68_imag <= _zz_20863[15 : 0];
        data_mid_4_real <= _zz_20871[15 : 0];
        data_mid_4_imag <= _zz_20879[15 : 0];
      end
      if((current_level_value == 3'b111))begin
        data_mid_69_real <= _zz_20896[15 : 0];
        data_mid_69_imag <= _zz_20904[15 : 0];
        data_mid_5_real <= _zz_20912[15 : 0];
        data_mid_5_imag <= _zz_20920[15 : 0];
      end
      if((current_level_value == 3'b111))begin
        data_mid_70_real <= _zz_20937[15 : 0];
        data_mid_70_imag <= _zz_20945[15 : 0];
        data_mid_6_real <= _zz_20953[15 : 0];
        data_mid_6_imag <= _zz_20961[15 : 0];
      end
      if((current_level_value == 3'b111))begin
        data_mid_71_real <= _zz_20978[15 : 0];
        data_mid_71_imag <= _zz_20986[15 : 0];
        data_mid_7_real <= _zz_20994[15 : 0];
        data_mid_7_imag <= _zz_21002[15 : 0];
      end
      if((current_level_value == 3'b111))begin
        data_mid_72_real <= _zz_21019[15 : 0];
        data_mid_72_imag <= _zz_21027[15 : 0];
        data_mid_8_real <= _zz_21035[15 : 0];
        data_mid_8_imag <= _zz_21043[15 : 0];
      end
      if((current_level_value == 3'b111))begin
        data_mid_73_real <= _zz_21060[15 : 0];
        data_mid_73_imag <= _zz_21068[15 : 0];
        data_mid_9_real <= _zz_21076[15 : 0];
        data_mid_9_imag <= _zz_21084[15 : 0];
      end
      if((current_level_value == 3'b111))begin
        data_mid_74_real <= _zz_21101[15 : 0];
        data_mid_74_imag <= _zz_21109[15 : 0];
        data_mid_10_real <= _zz_21117[15 : 0];
        data_mid_10_imag <= _zz_21125[15 : 0];
      end
      if((current_level_value == 3'b111))begin
        data_mid_75_real <= _zz_21142[15 : 0];
        data_mid_75_imag <= _zz_21150[15 : 0];
        data_mid_11_real <= _zz_21158[15 : 0];
        data_mid_11_imag <= _zz_21166[15 : 0];
      end
      if((current_level_value == 3'b111))begin
        data_mid_76_real <= _zz_21183[15 : 0];
        data_mid_76_imag <= _zz_21191[15 : 0];
        data_mid_12_real <= _zz_21199[15 : 0];
        data_mid_12_imag <= _zz_21207[15 : 0];
      end
      if((current_level_value == 3'b111))begin
        data_mid_77_real <= _zz_21224[15 : 0];
        data_mid_77_imag <= _zz_21232[15 : 0];
        data_mid_13_real <= _zz_21240[15 : 0];
        data_mid_13_imag <= _zz_21248[15 : 0];
      end
      if((current_level_value == 3'b111))begin
        data_mid_78_real <= _zz_21265[15 : 0];
        data_mid_78_imag <= _zz_21273[15 : 0];
        data_mid_14_real <= _zz_21281[15 : 0];
        data_mid_14_imag <= _zz_21289[15 : 0];
      end
      if((current_level_value == 3'b111))begin
        data_mid_79_real <= _zz_21306[15 : 0];
        data_mid_79_imag <= _zz_21314[15 : 0];
        data_mid_15_real <= _zz_21322[15 : 0];
        data_mid_15_imag <= _zz_21330[15 : 0];
      end
      if((current_level_value == 3'b111))begin
        data_mid_80_real <= _zz_21347[15 : 0];
        data_mid_80_imag <= _zz_21355[15 : 0];
        data_mid_16_real <= _zz_21363[15 : 0];
        data_mid_16_imag <= _zz_21371[15 : 0];
      end
      if((current_level_value == 3'b111))begin
        data_mid_81_real <= _zz_21388[15 : 0];
        data_mid_81_imag <= _zz_21396[15 : 0];
        data_mid_17_real <= _zz_21404[15 : 0];
        data_mid_17_imag <= _zz_21412[15 : 0];
      end
      if((current_level_value == 3'b111))begin
        data_mid_82_real <= _zz_21429[15 : 0];
        data_mid_82_imag <= _zz_21437[15 : 0];
        data_mid_18_real <= _zz_21445[15 : 0];
        data_mid_18_imag <= _zz_21453[15 : 0];
      end
      if((current_level_value == 3'b111))begin
        data_mid_83_real <= _zz_21470[15 : 0];
        data_mid_83_imag <= _zz_21478[15 : 0];
        data_mid_19_real <= _zz_21486[15 : 0];
        data_mid_19_imag <= _zz_21494[15 : 0];
      end
      if((current_level_value == 3'b111))begin
        data_mid_84_real <= _zz_21511[15 : 0];
        data_mid_84_imag <= _zz_21519[15 : 0];
        data_mid_20_real <= _zz_21527[15 : 0];
        data_mid_20_imag <= _zz_21535[15 : 0];
      end
      if((current_level_value == 3'b111))begin
        data_mid_85_real <= _zz_21552[15 : 0];
        data_mid_85_imag <= _zz_21560[15 : 0];
        data_mid_21_real <= _zz_21568[15 : 0];
        data_mid_21_imag <= _zz_21576[15 : 0];
      end
      if((current_level_value == 3'b111))begin
        data_mid_86_real <= _zz_21593[15 : 0];
        data_mid_86_imag <= _zz_21601[15 : 0];
        data_mid_22_real <= _zz_21609[15 : 0];
        data_mid_22_imag <= _zz_21617[15 : 0];
      end
      if((current_level_value == 3'b111))begin
        data_mid_87_real <= _zz_21634[15 : 0];
        data_mid_87_imag <= _zz_21642[15 : 0];
        data_mid_23_real <= _zz_21650[15 : 0];
        data_mid_23_imag <= _zz_21658[15 : 0];
      end
      if((current_level_value == 3'b111))begin
        data_mid_88_real <= _zz_21675[15 : 0];
        data_mid_88_imag <= _zz_21683[15 : 0];
        data_mid_24_real <= _zz_21691[15 : 0];
        data_mid_24_imag <= _zz_21699[15 : 0];
      end
      if((current_level_value == 3'b111))begin
        data_mid_89_real <= _zz_21716[15 : 0];
        data_mid_89_imag <= _zz_21724[15 : 0];
        data_mid_25_real <= _zz_21732[15 : 0];
        data_mid_25_imag <= _zz_21740[15 : 0];
      end
      if((current_level_value == 3'b111))begin
        data_mid_90_real <= _zz_21757[15 : 0];
        data_mid_90_imag <= _zz_21765[15 : 0];
        data_mid_26_real <= _zz_21773[15 : 0];
        data_mid_26_imag <= _zz_21781[15 : 0];
      end
      if((current_level_value == 3'b111))begin
        data_mid_91_real <= _zz_21798[15 : 0];
        data_mid_91_imag <= _zz_21806[15 : 0];
        data_mid_27_real <= _zz_21814[15 : 0];
        data_mid_27_imag <= _zz_21822[15 : 0];
      end
      if((current_level_value == 3'b111))begin
        data_mid_92_real <= _zz_21839[15 : 0];
        data_mid_92_imag <= _zz_21847[15 : 0];
        data_mid_28_real <= _zz_21855[15 : 0];
        data_mid_28_imag <= _zz_21863[15 : 0];
      end
      if((current_level_value == 3'b111))begin
        data_mid_93_real <= _zz_21880[15 : 0];
        data_mid_93_imag <= _zz_21888[15 : 0];
        data_mid_29_real <= _zz_21896[15 : 0];
        data_mid_29_imag <= _zz_21904[15 : 0];
      end
      if((current_level_value == 3'b111))begin
        data_mid_94_real <= _zz_21921[15 : 0];
        data_mid_94_imag <= _zz_21929[15 : 0];
        data_mid_30_real <= _zz_21937[15 : 0];
        data_mid_30_imag <= _zz_21945[15 : 0];
      end
      if((current_level_value == 3'b111))begin
        data_mid_95_real <= _zz_21962[15 : 0];
        data_mid_95_imag <= _zz_21970[15 : 0];
        data_mid_31_real <= _zz_21978[15 : 0];
        data_mid_31_imag <= _zz_21986[15 : 0];
      end
      if((current_level_value == 3'b111))begin
        data_mid_96_real <= _zz_22003[15 : 0];
        data_mid_96_imag <= _zz_22011[15 : 0];
        data_mid_32_real <= _zz_22019[15 : 0];
        data_mid_32_imag <= _zz_22027[15 : 0];
      end
      if((current_level_value == 3'b111))begin
        data_mid_97_real <= _zz_22044[15 : 0];
        data_mid_97_imag <= _zz_22052[15 : 0];
        data_mid_33_real <= _zz_22060[15 : 0];
        data_mid_33_imag <= _zz_22068[15 : 0];
      end
      if((current_level_value == 3'b111))begin
        data_mid_98_real <= _zz_22085[15 : 0];
        data_mid_98_imag <= _zz_22093[15 : 0];
        data_mid_34_real <= _zz_22101[15 : 0];
        data_mid_34_imag <= _zz_22109[15 : 0];
      end
      if((current_level_value == 3'b111))begin
        data_mid_99_real <= _zz_22126[15 : 0];
        data_mid_99_imag <= _zz_22134[15 : 0];
        data_mid_35_real <= _zz_22142[15 : 0];
        data_mid_35_imag <= _zz_22150[15 : 0];
      end
      if((current_level_value == 3'b111))begin
        data_mid_100_real <= _zz_22167[15 : 0];
        data_mid_100_imag <= _zz_22175[15 : 0];
        data_mid_36_real <= _zz_22183[15 : 0];
        data_mid_36_imag <= _zz_22191[15 : 0];
      end
      if((current_level_value == 3'b111))begin
        data_mid_101_real <= _zz_22208[15 : 0];
        data_mid_101_imag <= _zz_22216[15 : 0];
        data_mid_37_real <= _zz_22224[15 : 0];
        data_mid_37_imag <= _zz_22232[15 : 0];
      end
      if((current_level_value == 3'b111))begin
        data_mid_102_real <= _zz_22249[15 : 0];
        data_mid_102_imag <= _zz_22257[15 : 0];
        data_mid_38_real <= _zz_22265[15 : 0];
        data_mid_38_imag <= _zz_22273[15 : 0];
      end
      if((current_level_value == 3'b111))begin
        data_mid_103_real <= _zz_22290[15 : 0];
        data_mid_103_imag <= _zz_22298[15 : 0];
        data_mid_39_real <= _zz_22306[15 : 0];
        data_mid_39_imag <= _zz_22314[15 : 0];
      end
      if((current_level_value == 3'b111))begin
        data_mid_104_real <= _zz_22331[15 : 0];
        data_mid_104_imag <= _zz_22339[15 : 0];
        data_mid_40_real <= _zz_22347[15 : 0];
        data_mid_40_imag <= _zz_22355[15 : 0];
      end
      if((current_level_value == 3'b111))begin
        data_mid_105_real <= _zz_22372[15 : 0];
        data_mid_105_imag <= _zz_22380[15 : 0];
        data_mid_41_real <= _zz_22388[15 : 0];
        data_mid_41_imag <= _zz_22396[15 : 0];
      end
      if((current_level_value == 3'b111))begin
        data_mid_106_real <= _zz_22413[15 : 0];
        data_mid_106_imag <= _zz_22421[15 : 0];
        data_mid_42_real <= _zz_22429[15 : 0];
        data_mid_42_imag <= _zz_22437[15 : 0];
      end
      if((current_level_value == 3'b111))begin
        data_mid_107_real <= _zz_22454[15 : 0];
        data_mid_107_imag <= _zz_22462[15 : 0];
        data_mid_43_real <= _zz_22470[15 : 0];
        data_mid_43_imag <= _zz_22478[15 : 0];
      end
      if((current_level_value == 3'b111))begin
        data_mid_108_real <= _zz_22495[15 : 0];
        data_mid_108_imag <= _zz_22503[15 : 0];
        data_mid_44_real <= _zz_22511[15 : 0];
        data_mid_44_imag <= _zz_22519[15 : 0];
      end
      if((current_level_value == 3'b111))begin
        data_mid_109_real <= _zz_22536[15 : 0];
        data_mid_109_imag <= _zz_22544[15 : 0];
        data_mid_45_real <= _zz_22552[15 : 0];
        data_mid_45_imag <= _zz_22560[15 : 0];
      end
      if((current_level_value == 3'b111))begin
        data_mid_110_real <= _zz_22577[15 : 0];
        data_mid_110_imag <= _zz_22585[15 : 0];
        data_mid_46_real <= _zz_22593[15 : 0];
        data_mid_46_imag <= _zz_22601[15 : 0];
      end
      if((current_level_value == 3'b111))begin
        data_mid_111_real <= _zz_22618[15 : 0];
        data_mid_111_imag <= _zz_22626[15 : 0];
        data_mid_47_real <= _zz_22634[15 : 0];
        data_mid_47_imag <= _zz_22642[15 : 0];
      end
      if((current_level_value == 3'b111))begin
        data_mid_112_real <= _zz_22659[15 : 0];
        data_mid_112_imag <= _zz_22667[15 : 0];
        data_mid_48_real <= _zz_22675[15 : 0];
        data_mid_48_imag <= _zz_22683[15 : 0];
      end
      if((current_level_value == 3'b111))begin
        data_mid_113_real <= _zz_22700[15 : 0];
        data_mid_113_imag <= _zz_22708[15 : 0];
        data_mid_49_real <= _zz_22716[15 : 0];
        data_mid_49_imag <= _zz_22724[15 : 0];
      end
      if((current_level_value == 3'b111))begin
        data_mid_114_real <= _zz_22741[15 : 0];
        data_mid_114_imag <= _zz_22749[15 : 0];
        data_mid_50_real <= _zz_22757[15 : 0];
        data_mid_50_imag <= _zz_22765[15 : 0];
      end
      if((current_level_value == 3'b111))begin
        data_mid_115_real <= _zz_22782[15 : 0];
        data_mid_115_imag <= _zz_22790[15 : 0];
        data_mid_51_real <= _zz_22798[15 : 0];
        data_mid_51_imag <= _zz_22806[15 : 0];
      end
      if((current_level_value == 3'b111))begin
        data_mid_116_real <= _zz_22823[15 : 0];
        data_mid_116_imag <= _zz_22831[15 : 0];
        data_mid_52_real <= _zz_22839[15 : 0];
        data_mid_52_imag <= _zz_22847[15 : 0];
      end
      if((current_level_value == 3'b111))begin
        data_mid_117_real <= _zz_22864[15 : 0];
        data_mid_117_imag <= _zz_22872[15 : 0];
        data_mid_53_real <= _zz_22880[15 : 0];
        data_mid_53_imag <= _zz_22888[15 : 0];
      end
      if((current_level_value == 3'b111))begin
        data_mid_118_real <= _zz_22905[15 : 0];
        data_mid_118_imag <= _zz_22913[15 : 0];
        data_mid_54_real <= _zz_22921[15 : 0];
        data_mid_54_imag <= _zz_22929[15 : 0];
      end
      if((current_level_value == 3'b111))begin
        data_mid_119_real <= _zz_22946[15 : 0];
        data_mid_119_imag <= _zz_22954[15 : 0];
        data_mid_55_real <= _zz_22962[15 : 0];
        data_mid_55_imag <= _zz_22970[15 : 0];
      end
      if((current_level_value == 3'b111))begin
        data_mid_120_real <= _zz_22987[15 : 0];
        data_mid_120_imag <= _zz_22995[15 : 0];
        data_mid_56_real <= _zz_23003[15 : 0];
        data_mid_56_imag <= _zz_23011[15 : 0];
      end
      if((current_level_value == 3'b111))begin
        data_mid_121_real <= _zz_23028[15 : 0];
        data_mid_121_imag <= _zz_23036[15 : 0];
        data_mid_57_real <= _zz_23044[15 : 0];
        data_mid_57_imag <= _zz_23052[15 : 0];
      end
      if((current_level_value == 3'b111))begin
        data_mid_122_real <= _zz_23069[15 : 0];
        data_mid_122_imag <= _zz_23077[15 : 0];
        data_mid_58_real <= _zz_23085[15 : 0];
        data_mid_58_imag <= _zz_23093[15 : 0];
      end
      if((current_level_value == 3'b111))begin
        data_mid_123_real <= _zz_23110[15 : 0];
        data_mid_123_imag <= _zz_23118[15 : 0];
        data_mid_59_real <= _zz_23126[15 : 0];
        data_mid_59_imag <= _zz_23134[15 : 0];
      end
      if((current_level_value == 3'b111))begin
        data_mid_124_real <= _zz_23151[15 : 0];
        data_mid_124_imag <= _zz_23159[15 : 0];
        data_mid_60_real <= _zz_23167[15 : 0];
        data_mid_60_imag <= _zz_23175[15 : 0];
      end
      if((current_level_value == 3'b111))begin
        data_mid_125_real <= _zz_23192[15 : 0];
        data_mid_125_imag <= _zz_23200[15 : 0];
        data_mid_61_real <= _zz_23208[15 : 0];
        data_mid_61_imag <= _zz_23216[15 : 0];
      end
      if((current_level_value == 3'b111))begin
        data_mid_126_real <= _zz_23233[15 : 0];
        data_mid_126_imag <= _zz_23241[15 : 0];
        data_mid_62_real <= _zz_23249[15 : 0];
        data_mid_62_imag <= _zz_23257[15 : 0];
      end
      if((current_level_value == 3'b111))begin
        data_mid_127_real <= _zz_23274[15 : 0];
        data_mid_127_imag <= _zz_23282[15 : 0];
        data_mid_63_real <= _zz_23290[15 : 0];
        data_mid_63_imag <= _zz_23298[15 : 0];
      end
    end
  end

  always @ (posedge clk or posedge reset) begin
    if (reset) begin
      io_data_in_valid_regNext <= 1'b0;
      current_level_value <= 3'b000;
      null_cond_period_minus_1 <= 1'b0;
      current_level_willOverflow_regNext <= 1'b0;
    end else begin
      io_data_in_valid_regNext <= io_data_in_valid;
      current_level_value <= current_level_valueNext;
      if(io_data_in_valid_regNext)begin
        null_cond_period_minus_1 <= 1'b1;
      end else begin
        if(current_level_willOverflow)begin
          null_cond_period_minus_1 <= 1'b0;
        end
      end
      current_level_willOverflow_regNext <= current_level_willOverflow;
    end
  end


endmodule

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

module SInt32fixTo23_8_ROUNDTOINF (
  input      [31:0]   din,
  output     [15:0]   dout
);
  wire       [32:0]   _zz_9;
  wire       [32:0]   _zz_10;
  wire       [7:0]    _zz_11;
  wire       [24:0]   _zz_12;
  wire       [24:0]   _zz_13;
  wire       [32:0]   _zz_14;
  wire       [32:0]   _zz_15;
  wire       [32:0]   _zz_16;
  wire       [9:0]    _zz_17;
  wire       [8:0]    _zz_18;
  reg        [24:0]   _zz_1;
  wire       [31:0]   _zz_2;
  wire       [31:0]   _zz_3;
  wire       [31:0]   _zz_4;
  wire       [32:0]   _zz_5;
  wire       [31:0]   _zz_6;
  reg        [24:0]   _zz_7;
  reg        [15:0]   _zz_8;

  assign _zz_9 = {_zz_4[31],_zz_4};
  assign _zz_10 = {_zz_3[31],_zz_3};
  assign _zz_11 = _zz_5[7 : 0];
  assign _zz_12 = _zz_5[32 : 8];
  assign _zz_13 = 25'h0000001;
  assign _zz_14 = ($signed(_zz_15) + $signed(_zz_16));
  assign _zz_15 = {_zz_6[31],_zz_6};
  assign _zz_16 = {_zz_2[31],_zz_2};
  assign _zz_17 = _zz_1[24 : 15];
  assign _zz_18 = _zz_1[23 : 15];
  assign _zz_2 = {{24'h0,1'b1},7'h0};
  assign _zz_3 = {25'h1ffffff,7'h0};
  assign _zz_4 = din[31 : 0];
  assign _zz_5 = ($signed(_zz_9) + $signed(_zz_10));
  assign _zz_6 = din[31 : 0];
  always @ (*) begin
    if((_zz_11 != 8'h0))begin
      _zz_7 = ($signed(_zz_12) + $signed(_zz_13));
    end else begin
      _zz_7 = _zz_5[32 : 8];
    end
  end

  always @ (*) begin
    if(_zz_5[32])begin
      _zz_1 = _zz_7;
    end else begin
      _zz_1 = (_zz_14 >>> 8);
    end
  end

  always @ (*) begin
    if(_zz_1[24])begin
      if((! (_zz_17 == 10'h3ff)))begin
        _zz_8 = 16'h8000;
      end else begin
        _zz_8 = _zz_1[15 : 0];
      end
    end else begin
      if((_zz_18 != 9'h0))begin
        _zz_8 = 16'h7fff;
      end else begin
        _zz_8 = _zz_1[15 : 0];
      end
    end
  end

  assign dout = _zz_8;

endmodule

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

module SInt32fixTo31_0_ROUNDTOINF (
  input      [31:0]   din,
  output     [31:0]   dout
);

  assign dout = din;

endmodule
