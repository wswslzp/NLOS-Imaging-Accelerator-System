// Generator : SpinalHDL v1.4.1    git head : d1b4746673438bc5f242515335278fa39a666c38
// Component : CoefGenArray
// Git hash  : 2a34fe18f42a28946060dbf37f9913e1060dc674



module CoefGenArray (
  input               io_wave_front_valid,
  input      [15:0]   io_wave_front_payload_0_0,
  input               io_distance_valid,
  input      [15:0]   io_distance_payload_0_0,
  input               io_timeshift_valid,
  input      [15:0]   io_timeshift_payload_0_0_real,
  input      [15:0]   io_timeshift_payload_0_0_imag,
  output              io_coef_valid,
  output     [15:0]   io_coef_payload_0_0_0_real,
  output     [15:0]   io_coef_payload_0_0_0_imag,
  input               clk,
  input               reset
);
  wire       [15:0]   coefGenCore_1_io_coef_real;
  wire       [15:0]   coefGenCore_1_io_coef_imag;
  reg        [15:0]   wave_front_0_0;
  reg        [15:0]   distance_0_0;
  reg        [15:0]   timeshift_0_0_real;
  reg        [15:0]   timeshift_0_0_imag;
  reg                 _zz_1;
  reg                 _zz_2;
  reg                 _zz_3;
  reg                 _zz_4;
  reg                 _zz_5;
  reg                 _zz_6;

  CoefGenCore coefGenCore_1 (
    .io_wave              (wave_front_0_0[15:0]              ), //i
    .io_distance          (distance_0_0[15:0]                ), //i
    .io_timeshift_real    (timeshift_0_0_real[15:0]          ), //i
    .io_timeshift_imag    (timeshift_0_0_imag[15:0]          ), //i
    .io_coef_real         (coefGenCore_1_io_coef_real[15:0]  ), //o
    .io_coef_imag         (coefGenCore_1_io_coef_imag[15:0]  ), //o
    .clk                  (clk                               ), //i
    .reset                (reset                             )  //i
  );
  assign io_coef_payload_0_0_0_real = coefGenCore_1_io_coef_real;
  assign io_coef_payload_0_0_0_imag = coefGenCore_1_io_coef_imag;
  assign io_coef_valid = _zz_6;
  always @ (posedge clk) begin
    if(io_wave_front_valid)begin
      wave_front_0_0 <= io_wave_front_payload_0_0;
    end
    if(io_distance_valid)begin
      distance_0_0 <= io_distance_payload_0_0;
    end
    if(io_timeshift_valid)begin
      timeshift_0_0_real <= io_timeshift_payload_0_0_real;
      timeshift_0_0_imag <= io_timeshift_payload_0_0_imag;
    end
    _zz_1 <= ((io_wave_front_valid && io_distance_valid) && io_timeshift_valid);
    _zz_2 <= _zz_1;
    _zz_3 <= _zz_2;
    _zz_4 <= _zz_3;
    _zz_5 <= _zz_4;
    _zz_6 <= _zz_5;
  end


endmodule

module CoefGenCore (
  input      [15:0]   io_wave,
  input      [15:0]   io_distance,
  input      [15:0]   io_timeshift_real,
  input      [15:0]   io_timeshift_imag,
  output     [15:0]   io_coef_real,
  output     [15:0]   io_coef_imag,
  input               clk,
  input               reset
);
  wire       [15:0]   _zz_413;
  wire       [15:0]   _zz_414;
  wire       [7:0]    _zz_415;
  wire       [7:0]    _zz_416;
  wire       [7:0]    _zz_417;
  wire       [7:0]    _zz_418;
  wire       [15:0]   _zz_419;
  wire       [15:0]   _zz_420;
  wire       [15:0]   _zz_421;
  wire       [15:0]   _zz_422;
  wire       [7:0]    _zz_423;
  wire       [15:0]   _zz_424;
  wire       [15:0]   _zz_425;
  wire       [15:0]   _zz_426;
  wire       [7:0]    _zz_427;
  wire       [15:0]   _zz_428;
  wire       [15:0]   _zz_429;
  wire       [15:0]   _zz_430;
  wire       [15:0]   _zz_431;
  wire       [15:0]   _zz_432;
  wire       [15:0]   _zz_433;
  wire       [15:0]   _zz_434;
  wire       [31:0]   _zz_435;
  wire       [31:0]   _zz_436;
  wire       [31:0]   _zz_437;
  wire       [31:0]   _zz_438;
  wire       [15:0]   _zz_439;
  wire       [31:0]   _zz_440;
  wire       [31:0]   _zz_441;
  wire       [31:0]   _zz_442;
  wire       [15:0]   _zz_443;
  wire       [31:0]   _zz_444;
  wire       [31:0]   _zz_445;
  wire       [31:0]   _zz_446;
  reg        [15:0]   _zz_447;
  reg        [15:0]   _zz_448;
  reg        [15:0]   _zz_449;
  reg        [15:0]   _zz_450;
  reg        [15:0]   _zz_451;
  reg        [15:0]   _zz_452;
  wire       [7:0]    fixTo_dout;
  wire       [7:0]    fixTo_1_dout;
  wire       [7:0]    fixTo_2_dout;
  wire       [7:0]    divUnit_1_c;
  wire       [7:0]    divUnit_2_c;
  wire       [15:0]   fixTo_3_dout;
  wire       [15:0]   fixTo_4_dout;
  wire       [15:0]   mulUnit_1_c;
  wire       [15:0]   fixTo_5_dout;
  wire       [15:0]   fixTo_6_dout;
  wire       [15:0]   fixTo_7_dout;
  wire       [15:0]   mulUnit_2_c;
  wire       [15:0]   fixTo_8_dout;
  wire       [15:0]   fixTo_9_dout;
  wire       [15:0]   fixTo_10_dout;
  wire       [15:0]   mulUnit_3_c;
  wire       [15:0]   fixTo_11_dout;
  wire       [15:0]   fixTo_12_dout;
  wire       [15:0]   fixTo_13_dout;
  wire       [15:0]   divUnit_3_c;
  wire       [15:0]   divUnit_4_c;
  wire       [31:0]   fixTo_14_dout;
  wire       [31:0]   fixTo_15_dout;
  wire       [31:0]   mulUnit_4_c;
  wire       [31:0]   fixTo_16_dout;
  wire       [31:0]   fixTo_17_dout;
  wire       [31:0]   fixTo_18_dout;
  wire       [31:0]   mulUnit_5_c;
  wire       [31:0]   fixTo_19_dout;
  wire       [31:0]   fixTo_20_dout;
  wire       [31:0]   fixTo_21_dout;
  wire       [31:0]   mulUnit_6_c;
  wire       [31:0]   fixTo_22_dout;
  wire       [15:0]   fixTo_23_dout;
  wire       [15:0]   fixTo_24_dout;
  wire                _zz_453;
  wire                _zz_454;
  wire       [7:0]    _zz_455;
  wire       [7:0]    _zz_456;
  wire       [15:0]   _zz_457;
  wire       [7:0]    _zz_458;
  wire       [15:0]   _zz_459;
  wire       [7:0]    _zz_460;
  wire       [15:0]   _zz_461;
  wire       [7:0]    _zz_462;
  wire       [15:0]   _zz_463;
  wire       [7:0]    _zz_464;
  wire       [15:0]   _zz_465;
  wire       [7:0]    _zz_466;
  wire       [15:0]   _zz_467;
  wire       [7:0]    _zz_468;
  wire       [15:0]   _zz_469;
  wire       [7:0]    _zz_470;
  wire       [15:0]   _zz_471;
  wire       [7:0]    _zz_472;
  wire       [15:0]   _zz_473;
  wire       [7:0]    _zz_474;
  wire       [15:0]   _zz_475;
  wire       [7:0]    _zz_476;
  wire       [15:0]   _zz_477;
  wire       [7:0]    _zz_478;
  wire       [15:0]   _zz_479;
  wire       [7:0]    _zz_480;
  wire       [15:0]   _zz_481;
  wire       [7:0]    _zz_482;
  wire       [15:0]   _zz_483;
  wire       [7:0]    _zz_484;
  wire       [15:0]   _zz_485;
  wire       [7:0]    _zz_486;
  wire       [15:0]   _zz_487;
  wire       [7:0]    _zz_488;
  wire       [15:0]   _zz_489;
  wire       [7:0]    _zz_490;
  wire       [15:0]   _zz_491;
  wire       [7:0]    _zz_492;
  wire       [15:0]   _zz_493;
  wire       [7:0]    _zz_494;
  wire       [15:0]   _zz_495;
  wire       [7:0]    _zz_496;
  wire       [15:0]   _zz_497;
  wire       [7:0]    _zz_498;
  wire       [15:0]   _zz_499;
  wire       [7:0]    _zz_500;
  wire       [15:0]   _zz_501;
  wire       [7:0]    _zz_502;
  wire       [15:0]   _zz_503;
  wire       [7:0]    _zz_504;
  wire       [15:0]   _zz_505;
  wire       [7:0]    _zz_506;
  wire       [15:0]   _zz_507;
  wire       [7:0]    _zz_508;
  wire       [15:0]   _zz_509;
  wire       [7:0]    _zz_510;
  wire       [15:0]   _zz_511;
  wire       [7:0]    _zz_512;
  wire       [15:0]   _zz_513;
  wire       [7:0]    _zz_514;
  wire       [15:0]   _zz_515;
  wire       [7:0]    _zz_516;
  wire       [15:0]   _zz_517;
  wire       [7:0]    _zz_518;
  wire       [15:0]   _zz_519;
  wire       [7:0]    _zz_520;
  wire       [15:0]   _zz_521;
  wire       [7:0]    _zz_522;
  wire       [15:0]   _zz_523;
  wire       [7:0]    _zz_524;
  wire       [15:0]   _zz_525;
  wire       [7:0]    _zz_526;
  wire       [15:0]   _zz_527;
  wire       [7:0]    _zz_528;
  wire       [15:0]   _zz_529;
  wire       [7:0]    _zz_530;
  wire       [15:0]   _zz_531;
  wire       [7:0]    _zz_532;
  wire       [15:0]   _zz_533;
  wire       [7:0]    _zz_534;
  wire       [15:0]   _zz_535;
  wire       [7:0]    _zz_536;
  wire       [15:0]   _zz_537;
  wire       [7:0]    _zz_538;
  wire       [15:0]   _zz_539;
  wire       [7:0]    _zz_540;
  wire       [15:0]   _zz_541;
  wire       [7:0]    _zz_542;
  wire       [15:0]   _zz_543;
  wire       [7:0]    _zz_544;
  wire       [15:0]   _zz_545;
  wire       [7:0]    _zz_546;
  wire       [15:0]   _zz_547;
  wire       [7:0]    _zz_548;
  wire       [15:0]   _zz_549;
  wire       [7:0]    _zz_550;
  wire       [15:0]   _zz_551;
  wire       [7:0]    _zz_552;
  wire       [15:0]   _zz_553;
  wire       [7:0]    _zz_554;
  wire       [15:0]   _zz_555;
  wire       [7:0]    _zz_556;
  wire       [15:0]   _zz_557;
  wire       [7:0]    _zz_558;
  wire       [15:0]   _zz_559;
  wire       [7:0]    _zz_560;
  wire       [15:0]   _zz_561;
  wire       [7:0]    _zz_562;
  wire       [15:0]   _zz_563;
  wire       [7:0]    _zz_564;
  wire       [15:0]   _zz_565;
  wire       [7:0]    _zz_566;
  wire       [15:0]   _zz_567;
  wire       [7:0]    _zz_568;
  wire       [15:0]   _zz_569;
  wire       [7:0]    _zz_570;
  wire       [15:0]   _zz_571;
  wire       [7:0]    _zz_572;
  wire       [15:0]   _zz_573;
  wire       [7:0]    _zz_574;
  wire       [15:0]   _zz_575;
  wire       [7:0]    _zz_576;
  wire       [15:0]   _zz_577;
  wire       [7:0]    _zz_578;
  wire       [15:0]   _zz_579;
  wire       [7:0]    _zz_580;
  wire       [15:0]   _zz_581;
  wire       [7:0]    _zz_582;
  wire       [15:0]   _zz_583;
  wire       [7:0]    _zz_584;
  wire       [15:0]   _zz_585;
  wire       [7:0]    _zz_586;
  wire       [15:0]   _zz_587;
  wire       [7:0]    _zz_588;
  wire       [15:0]   _zz_589;
  wire       [7:0]    _zz_590;
  wire       [15:0]   _zz_591;
  wire       [7:0]    _zz_592;
  wire       [15:0]   _zz_593;
  wire       [7:0]    _zz_594;
  wire       [15:0]   _zz_595;
  wire       [7:0]    _zz_596;
  wire       [15:0]   _zz_597;
  wire       [7:0]    _zz_598;
  wire       [15:0]   _zz_599;
  wire       [7:0]    _zz_600;
  wire       [15:0]   _zz_601;
  wire       [7:0]    _zz_602;
  wire       [15:0]   _zz_603;
  wire       [7:0]    _zz_604;
  wire       [15:0]   _zz_605;
  wire       [7:0]    _zz_606;
  wire       [15:0]   _zz_607;
  wire       [7:0]    _zz_608;
  wire       [15:0]   _zz_609;
  wire       [7:0]    _zz_610;
  wire       [15:0]   _zz_611;
  wire       [7:0]    _zz_612;
  wire       [15:0]   _zz_613;
  wire       [7:0]    _zz_614;
  wire       [15:0]   _zz_615;
  wire       [7:0]    _zz_616;
  wire       [15:0]   _zz_617;
  wire       [7:0]    _zz_618;
  wire       [15:0]   _zz_619;
  wire       [7:0]    _zz_620;
  wire       [15:0]   _zz_621;
  wire       [7:0]    _zz_622;
  wire       [15:0]   _zz_623;
  wire       [7:0]    _zz_624;
  wire       [15:0]   _zz_625;
  wire       [7:0]    _zz_626;
  wire       [15:0]   _zz_627;
  wire       [7:0]    _zz_628;
  wire       [15:0]   _zz_629;
  wire       [7:0]    _zz_630;
  wire       [15:0]   _zz_631;
  wire       [7:0]    _zz_632;
  wire       [15:0]   _zz_633;
  wire       [7:0]    _zz_634;
  wire       [15:0]   _zz_635;
  wire       [7:0]    _zz_636;
  wire       [15:0]   _zz_637;
  wire       [7:0]    _zz_638;
  wire       [15:0]   _zz_639;
  wire       [7:0]    _zz_640;
  wire       [15:0]   _zz_641;
  wire       [7:0]    _zz_642;
  wire       [15:0]   _zz_643;
  wire       [7:0]    _zz_644;
  wire       [15:0]   _zz_645;
  wire       [7:0]    _zz_646;
  wire       [15:0]   _zz_647;
  wire       [7:0]    _zz_648;
  wire       [15:0]   _zz_649;
  wire       [7:0]    _zz_650;
  wire       [15:0]   _zz_651;
  wire       [7:0]    _zz_652;
  wire       [15:0]   _zz_653;
  wire       [7:0]    _zz_654;
  wire       [15:0]   _zz_655;
  wire       [7:0]    _zz_656;
  wire       [15:0]   _zz_657;
  wire       [7:0]    _zz_658;
  wire       [15:0]   _zz_659;
  wire       [7:0]    _zz_660;
  wire       [15:0]   _zz_661;
  wire       [7:0]    _zz_662;
  wire       [15:0]   _zz_663;
  wire       [7:0]    _zz_664;
  wire       [15:0]   _zz_665;
  wire       [7:0]    _zz_666;
  wire       [15:0]   _zz_667;
  wire       [7:0]    _zz_668;
  wire       [15:0]   _zz_669;
  wire       [7:0]    _zz_670;
  wire       [15:0]   _zz_671;
  wire       [7:0]    _zz_672;
  wire       [15:0]   _zz_673;
  wire       [7:0]    _zz_674;
  wire       [15:0]   _zz_675;
  wire       [7:0]    _zz_676;
  wire       [15:0]   _zz_677;
  wire       [7:0]    _zz_678;
  wire       [15:0]   _zz_679;
  wire       [7:0]    _zz_680;
  wire       [15:0]   _zz_681;
  wire       [7:0]    _zz_682;
  wire       [15:0]   _zz_683;
  wire       [7:0]    _zz_684;
  wire       [15:0]   _zz_685;
  wire       [7:0]    _zz_686;
  wire       [15:0]   _zz_687;
  wire       [7:0]    _zz_688;
  wire       [15:0]   _zz_689;
  wire       [7:0]    _zz_690;
  wire       [15:0]   _zz_691;
  wire       [7:0]    _zz_692;
  wire       [15:0]   _zz_693;
  wire       [7:0]    _zz_694;
  wire       [15:0]   _zz_695;
  wire       [7:0]    _zz_696;
  wire       [15:0]   _zz_697;
  wire       [7:0]    _zz_698;
  wire       [15:0]   _zz_699;
  wire       [7:0]    _zz_700;
  wire       [15:0]   _zz_701;
  wire       [7:0]    _zz_702;
  wire       [15:0]   _zz_703;
  wire       [7:0]    _zz_704;
  wire       [15:0]   _zz_705;
  wire       [7:0]    _zz_706;
  wire       [15:0]   _zz_707;
  wire       [7:0]    _zz_708;
  wire       [15:0]   _zz_709;
  wire       [7:0]    _zz_710;
  wire       [15:0]   _zz_711;
  wire       [1:0]    _zz_712;
  wire       [0:0]    _zz_713;
  wire       [1:0]    _zz_714;
  wire       [0:0]    _zz_715;
  wire       [1:0]    _zz_716;
  wire       [2:0]    _zz_717;
  wire       [1:0]    _zz_718;
  wire       [2:0]    _zz_719;
  wire       [1:0]    _zz_720;
  wire       [1:0]    _zz_721;
  wire       [0:0]    _zz_722;
  wire       [1:0]    _zz_723;
  wire       [0:0]    _zz_724;
  wire       [1:0]    _zz_725;
  wire       [1:0]    _zz_726;
  wire       [2:0]    _zz_727;
  wire       [1:0]    _zz_728;
  wire       [3:0]    _zz_729;
  wire       [2:0]    _zz_730;
  wire       [3:0]    _zz_731;
  wire       [2:0]    _zz_732;
  wire       [1:0]    _zz_733;
  wire       [0:0]    _zz_734;
  wire       [1:0]    _zz_735;
  wire       [0:0]    _zz_736;
  wire       [1:0]    _zz_737;
  wire       [2:0]    _zz_738;
  wire       [1:0]    _zz_739;
  wire       [2:0]    _zz_740;
  wire       [1:0]    _zz_741;
  wire       [1:0]    _zz_742;
  wire       [0:0]    _zz_743;
  wire       [1:0]    _zz_744;
  wire       [0:0]    _zz_745;
  wire       [1:0]    _zz_746;
  wire       [1:0]    _zz_747;
  wire       [2:0]    _zz_748;
  wire       [1:0]    _zz_749;
  wire       [2:0]    _zz_750;
  wire       [3:0]    _zz_751;
  wire       [2:0]    _zz_752;
  wire       [4:0]    _zz_753;
  wire       [3:0]    _zz_754;
  wire       [4:0]    _zz_755;
  wire       [3:0]    _zz_756;
  wire       [1:0]    _zz_757;
  wire       [0:0]    _zz_758;
  wire       [1:0]    _zz_759;
  wire       [0:0]    _zz_760;
  wire       [1:0]    _zz_761;
  wire       [2:0]    _zz_762;
  wire       [1:0]    _zz_763;
  wire       [2:0]    _zz_764;
  wire       [1:0]    _zz_765;
  wire       [1:0]    _zz_766;
  wire       [0:0]    _zz_767;
  wire       [1:0]    _zz_768;
  wire       [0:0]    _zz_769;
  wire       [1:0]    _zz_770;
  wire       [1:0]    _zz_771;
  wire       [2:0]    _zz_772;
  wire       [1:0]    _zz_773;
  wire       [3:0]    _zz_774;
  wire       [2:0]    _zz_775;
  wire       [3:0]    _zz_776;
  wire       [2:0]    _zz_777;
  wire       [1:0]    _zz_778;
  wire       [0:0]    _zz_779;
  wire       [1:0]    _zz_780;
  wire       [0:0]    _zz_781;
  wire       [1:0]    _zz_782;
  wire       [2:0]    _zz_783;
  wire       [1:0]    _zz_784;
  wire       [2:0]    _zz_785;
  wire       [1:0]    _zz_786;
  wire       [1:0]    _zz_787;
  wire       [0:0]    _zz_788;
  wire       [1:0]    _zz_789;
  wire       [0:0]    _zz_790;
  wire       [1:0]    _zz_791;
  wire       [1:0]    _zz_792;
  wire       [2:0]    _zz_793;
  wire       [1:0]    _zz_794;
  wire       [2:0]    _zz_795;
  wire       [3:0]    _zz_796;
  wire       [2:0]    _zz_797;
  wire       [3:0]    _zz_798;
  wire       [4:0]    _zz_799;
  wire       [3:0]    _zz_800;
  wire       [5:0]    _zz_801;
  wire       [4:0]    _zz_802;
  wire       [5:0]    _zz_803;
  wire       [4:0]    _zz_804;
  wire       [1:0]    _zz_805;
  wire       [0:0]    _zz_806;
  wire       [1:0]    _zz_807;
  wire       [0:0]    _zz_808;
  wire       [1:0]    _zz_809;
  wire       [2:0]    _zz_810;
  wire       [1:0]    _zz_811;
  wire       [2:0]    _zz_812;
  wire       [1:0]    _zz_813;
  wire       [1:0]    _zz_814;
  wire       [0:0]    _zz_815;
  wire       [1:0]    _zz_816;
  wire       [0:0]    _zz_817;
  wire       [1:0]    _zz_818;
  wire       [1:0]    _zz_819;
  wire       [2:0]    _zz_820;
  wire       [1:0]    _zz_821;
  wire       [3:0]    _zz_822;
  wire       [2:0]    _zz_823;
  wire       [3:0]    _zz_824;
  wire       [2:0]    _zz_825;
  wire       [1:0]    _zz_826;
  wire       [0:0]    _zz_827;
  wire       [1:0]    _zz_828;
  wire       [0:0]    _zz_829;
  wire       [1:0]    _zz_830;
  wire       [2:0]    _zz_831;
  wire       [1:0]    _zz_832;
  wire       [2:0]    _zz_833;
  wire       [1:0]    _zz_834;
  wire       [1:0]    _zz_835;
  wire       [0:0]    _zz_836;
  wire       [1:0]    _zz_837;
  wire       [0:0]    _zz_838;
  wire       [1:0]    _zz_839;
  wire       [1:0]    _zz_840;
  wire       [2:0]    _zz_841;
  wire       [1:0]    _zz_842;
  wire       [2:0]    _zz_843;
  wire       [3:0]    _zz_844;
  wire       [2:0]    _zz_845;
  wire       [4:0]    _zz_846;
  wire       [3:0]    _zz_847;
  wire       [4:0]    _zz_848;
  wire       [3:0]    _zz_849;
  wire       [1:0]    _zz_850;
  wire       [0:0]    _zz_851;
  wire       [1:0]    _zz_852;
  wire       [0:0]    _zz_853;
  wire       [1:0]    _zz_854;
  wire       [2:0]    _zz_855;
  wire       [1:0]    _zz_856;
  wire       [2:0]    _zz_857;
  wire       [1:0]    _zz_858;
  wire       [1:0]    _zz_859;
  wire       [0:0]    _zz_860;
  wire       [1:0]    _zz_861;
  wire       [0:0]    _zz_862;
  wire       [1:0]    _zz_863;
  wire       [1:0]    _zz_864;
  wire       [2:0]    _zz_865;
  wire       [1:0]    _zz_866;
  wire       [3:0]    _zz_867;
  wire       [2:0]    _zz_868;
  wire       [3:0]    _zz_869;
  wire       [2:0]    _zz_870;
  wire       [1:0]    _zz_871;
  wire       [0:0]    _zz_872;
  wire       [1:0]    _zz_873;
  wire       [0:0]    _zz_874;
  wire       [1:0]    _zz_875;
  wire       [2:0]    _zz_876;
  wire       [1:0]    _zz_877;
  wire       [2:0]    _zz_878;
  wire       [1:0]    _zz_879;
  wire       [1:0]    _zz_880;
  wire       [0:0]    _zz_881;
  wire       [1:0]    _zz_882;
  wire       [0:0]    _zz_883;
  wire       [1:0]    _zz_884;
  wire       [1:0]    _zz_885;
  wire       [2:0]    _zz_886;
  wire       [1:0]    _zz_887;
  wire       [2:0]    _zz_888;
  wire       [3:0]    _zz_889;
  wire       [2:0]    _zz_890;
  wire       [3:0]    _zz_891;
  wire       [4:0]    _zz_892;
  wire       [3:0]    _zz_893;
  wire       [4:0]    _zz_894;
  wire       [5:0]    _zz_895;
  wire       [4:0]    _zz_896;
  wire       [6:0]    _zz_897;
  wire       [5:0]    _zz_898;
  wire       [6:0]    _zz_899;
  wire       [5:0]    _zz_900;
  wire       [1:0]    _zz_901;
  wire       [0:0]    _zz_902;
  wire       [1:0]    _zz_903;
  wire       [0:0]    _zz_904;
  wire       [1:0]    _zz_905;
  wire       [2:0]    _zz_906;
  wire       [1:0]    _zz_907;
  wire       [2:0]    _zz_908;
  wire       [1:0]    _zz_909;
  wire       [1:0]    _zz_910;
  wire       [0:0]    _zz_911;
  wire       [1:0]    _zz_912;
  wire       [0:0]    _zz_913;
  wire       [1:0]    _zz_914;
  wire       [1:0]    _zz_915;
  wire       [2:0]    _zz_916;
  wire       [1:0]    _zz_917;
  wire       [3:0]    _zz_918;
  wire       [2:0]    _zz_919;
  wire       [3:0]    _zz_920;
  wire       [2:0]    _zz_921;
  wire       [1:0]    _zz_922;
  wire       [0:0]    _zz_923;
  wire       [1:0]    _zz_924;
  wire       [0:0]    _zz_925;
  wire       [1:0]    _zz_926;
  wire       [2:0]    _zz_927;
  wire       [1:0]    _zz_928;
  wire       [2:0]    _zz_929;
  wire       [1:0]    _zz_930;
  wire       [1:0]    _zz_931;
  wire       [0:0]    _zz_932;
  wire       [1:0]    _zz_933;
  wire       [0:0]    _zz_934;
  wire       [1:0]    _zz_935;
  wire       [1:0]    _zz_936;
  wire       [2:0]    _zz_937;
  wire       [1:0]    _zz_938;
  wire       [2:0]    _zz_939;
  wire       [3:0]    _zz_940;
  wire       [2:0]    _zz_941;
  wire       [4:0]    _zz_942;
  wire       [3:0]    _zz_943;
  wire       [4:0]    _zz_944;
  wire       [3:0]    _zz_945;
  wire       [1:0]    _zz_946;
  wire       [0:0]    _zz_947;
  wire       [1:0]    _zz_948;
  wire       [0:0]    _zz_949;
  wire       [1:0]    _zz_950;
  wire       [2:0]    _zz_951;
  wire       [1:0]    _zz_952;
  wire       [2:0]    _zz_953;
  wire       [1:0]    _zz_954;
  wire       [1:0]    _zz_955;
  wire       [0:0]    _zz_956;
  wire       [1:0]    _zz_957;
  wire       [0:0]    _zz_958;
  wire       [1:0]    _zz_959;
  wire       [1:0]    _zz_960;
  wire       [2:0]    _zz_961;
  wire       [1:0]    _zz_962;
  wire       [3:0]    _zz_963;
  wire       [2:0]    _zz_964;
  wire       [3:0]    _zz_965;
  wire       [2:0]    _zz_966;
  wire       [1:0]    _zz_967;
  wire       [0:0]    _zz_968;
  wire       [1:0]    _zz_969;
  wire       [0:0]    _zz_970;
  wire       [1:0]    _zz_971;
  wire       [2:0]    _zz_972;
  wire       [1:0]    _zz_973;
  wire       [2:0]    _zz_974;
  wire       [1:0]    _zz_975;
  wire       [1:0]    _zz_976;
  wire       [0:0]    _zz_977;
  wire       [1:0]    _zz_978;
  wire       [0:0]    _zz_979;
  wire       [1:0]    _zz_980;
  wire       [1:0]    _zz_981;
  wire       [2:0]    _zz_982;
  wire       [1:0]    _zz_983;
  wire       [2:0]    _zz_984;
  wire       [3:0]    _zz_985;
  wire       [2:0]    _zz_986;
  wire       [3:0]    _zz_987;
  wire       [4:0]    _zz_988;
  wire       [3:0]    _zz_989;
  wire       [5:0]    _zz_990;
  wire       [4:0]    _zz_991;
  wire       [5:0]    _zz_992;
  wire       [4:0]    _zz_993;
  wire       [1:0]    _zz_994;
  wire       [0:0]    _zz_995;
  wire       [1:0]    _zz_996;
  wire       [0:0]    _zz_997;
  wire       [1:0]    _zz_998;
  wire       [2:0]    _zz_999;
  wire       [1:0]    _zz_1000;
  wire       [2:0]    _zz_1001;
  wire       [1:0]    _zz_1002;
  wire       [1:0]    _zz_1003;
  wire       [0:0]    _zz_1004;
  wire       [1:0]    _zz_1005;
  wire       [0:0]    _zz_1006;
  wire       [1:0]    _zz_1007;
  wire       [1:0]    _zz_1008;
  wire       [2:0]    _zz_1009;
  wire       [1:0]    _zz_1010;
  wire       [3:0]    _zz_1011;
  wire       [2:0]    _zz_1012;
  wire       [3:0]    _zz_1013;
  wire       [2:0]    _zz_1014;
  wire       [1:0]    _zz_1015;
  wire       [0:0]    _zz_1016;
  wire       [1:0]    _zz_1017;
  wire       [0:0]    _zz_1018;
  wire       [1:0]    _zz_1019;
  wire       [2:0]    _zz_1020;
  wire       [1:0]    _zz_1021;
  wire       [2:0]    _zz_1022;
  wire       [1:0]    _zz_1023;
  wire       [1:0]    _zz_1024;
  wire       [0:0]    _zz_1025;
  wire       [1:0]    _zz_1026;
  wire       [0:0]    _zz_1027;
  wire       [1:0]    _zz_1028;
  wire       [1:0]    _zz_1029;
  wire       [2:0]    _zz_1030;
  wire       [1:0]    _zz_1031;
  wire       [2:0]    _zz_1032;
  wire       [3:0]    _zz_1033;
  wire       [2:0]    _zz_1034;
  wire       [4:0]    _zz_1035;
  wire       [3:0]    _zz_1036;
  wire       [4:0]    _zz_1037;
  wire       [3:0]    _zz_1038;
  wire       [1:0]    _zz_1039;
  wire       [0:0]    _zz_1040;
  wire       [1:0]    _zz_1041;
  wire       [0:0]    _zz_1042;
  wire       [1:0]    _zz_1043;
  wire       [2:0]    _zz_1044;
  wire       [1:0]    _zz_1045;
  wire       [2:0]    _zz_1046;
  wire       [1:0]    _zz_1047;
  wire       [1:0]    _zz_1048;
  wire       [0:0]    _zz_1049;
  wire       [1:0]    _zz_1050;
  wire       [0:0]    _zz_1051;
  wire       [1:0]    _zz_1052;
  wire       [1:0]    _zz_1053;
  wire       [2:0]    _zz_1054;
  wire       [1:0]    _zz_1055;
  wire       [3:0]    _zz_1056;
  wire       [2:0]    _zz_1057;
  wire       [3:0]    _zz_1058;
  wire       [2:0]    _zz_1059;
  wire       [1:0]    _zz_1060;
  wire       [0:0]    _zz_1061;
  wire       [1:0]    _zz_1062;
  wire       [0:0]    _zz_1063;
  wire       [1:0]    _zz_1064;
  wire       [2:0]    _zz_1065;
  wire       [1:0]    _zz_1066;
  wire       [2:0]    _zz_1067;
  wire       [1:0]    _zz_1068;
  wire       [1:0]    _zz_1069;
  wire       [0:0]    _zz_1070;
  wire       [1:0]    _zz_1071;
  wire       [0:0]    _zz_1072;
  wire       [1:0]    _zz_1073;
  wire       [1:0]    _zz_1074;
  wire       [2:0]    _zz_1075;
  wire       [1:0]    _zz_1076;
  wire       [2:0]    _zz_1077;
  wire       [3:0]    _zz_1078;
  wire       [2:0]    _zz_1079;
  wire       [3:0]    _zz_1080;
  wire       [4:0]    _zz_1081;
  wire       [3:0]    _zz_1082;
  wire       [4:0]    _zz_1083;
  wire       [5:0]    _zz_1084;
  wire       [4:0]    _zz_1085;
  wire       [5:0]    _zz_1086;
  wire       [6:0]    _zz_1087;
  wire       [5:0]    _zz_1088;
  wire       [7:0]    _zz_1089;
  wire       [6:0]    _zz_1090;
  wire       [7:0]    _zz_1091;
  wire       [6:0]    _zz_1092;
  wire       [1:0]    _zz_1093;
  wire       [0:0]    _zz_1094;
  wire       [1:0]    _zz_1095;
  wire       [0:0]    _zz_1096;
  wire       [1:0]    _zz_1097;
  wire       [2:0]    _zz_1098;
  wire       [1:0]    _zz_1099;
  wire       [2:0]    _zz_1100;
  wire       [1:0]    _zz_1101;
  wire       [1:0]    _zz_1102;
  wire       [0:0]    _zz_1103;
  wire       [1:0]    _zz_1104;
  wire       [0:0]    _zz_1105;
  wire       [1:0]    _zz_1106;
  wire       [1:0]    _zz_1107;
  wire       [2:0]    _zz_1108;
  wire       [1:0]    _zz_1109;
  wire       [3:0]    _zz_1110;
  wire       [2:0]    _zz_1111;
  wire       [3:0]    _zz_1112;
  wire       [2:0]    _zz_1113;
  wire       [1:0]    _zz_1114;
  wire       [0:0]    _zz_1115;
  wire       [1:0]    _zz_1116;
  wire       [0:0]    _zz_1117;
  wire       [1:0]    _zz_1118;
  wire       [2:0]    _zz_1119;
  wire       [1:0]    _zz_1120;
  wire       [2:0]    _zz_1121;
  wire       [1:0]    _zz_1122;
  wire       [1:0]    _zz_1123;
  wire       [0:0]    _zz_1124;
  wire       [1:0]    _zz_1125;
  wire       [0:0]    _zz_1126;
  wire       [1:0]    _zz_1127;
  wire       [1:0]    _zz_1128;
  wire       [2:0]    _zz_1129;
  wire       [1:0]    _zz_1130;
  wire       [2:0]    _zz_1131;
  wire       [3:0]    _zz_1132;
  wire       [2:0]    _zz_1133;
  wire       [4:0]    _zz_1134;
  wire       [3:0]    _zz_1135;
  wire       [4:0]    _zz_1136;
  wire       [3:0]    _zz_1137;
  wire       [1:0]    _zz_1138;
  wire       [0:0]    _zz_1139;
  wire       [1:0]    _zz_1140;
  wire       [0:0]    _zz_1141;
  wire       [1:0]    _zz_1142;
  wire       [2:0]    _zz_1143;
  wire       [1:0]    _zz_1144;
  wire       [2:0]    _zz_1145;
  wire       [1:0]    _zz_1146;
  wire       [1:0]    _zz_1147;
  wire       [0:0]    _zz_1148;
  wire       [1:0]    _zz_1149;
  wire       [0:0]    _zz_1150;
  wire       [1:0]    _zz_1151;
  wire       [1:0]    _zz_1152;
  wire       [2:0]    _zz_1153;
  wire       [1:0]    _zz_1154;
  wire       [3:0]    _zz_1155;
  wire       [2:0]    _zz_1156;
  wire       [3:0]    _zz_1157;
  wire       [2:0]    _zz_1158;
  wire       [1:0]    _zz_1159;
  wire       [0:0]    _zz_1160;
  wire       [1:0]    _zz_1161;
  wire       [0:0]    _zz_1162;
  wire       [1:0]    _zz_1163;
  wire       [2:0]    _zz_1164;
  wire       [1:0]    _zz_1165;
  wire       [2:0]    _zz_1166;
  wire       [1:0]    _zz_1167;
  wire       [1:0]    _zz_1168;
  wire       [0:0]    _zz_1169;
  wire       [1:0]    _zz_1170;
  wire       [0:0]    _zz_1171;
  wire       [1:0]    _zz_1172;
  wire       [1:0]    _zz_1173;
  wire       [2:0]    _zz_1174;
  wire       [1:0]    _zz_1175;
  wire       [2:0]    _zz_1176;
  wire       [3:0]    _zz_1177;
  wire       [2:0]    _zz_1178;
  wire       [3:0]    _zz_1179;
  wire       [4:0]    _zz_1180;
  wire       [3:0]    _zz_1181;
  wire       [5:0]    _zz_1182;
  wire       [4:0]    _zz_1183;
  wire       [5:0]    _zz_1184;
  wire       [4:0]    _zz_1185;
  wire       [1:0]    _zz_1186;
  wire       [0:0]    _zz_1187;
  wire       [1:0]    _zz_1188;
  wire       [0:0]    _zz_1189;
  wire       [1:0]    _zz_1190;
  wire       [2:0]    _zz_1191;
  wire       [1:0]    _zz_1192;
  wire       [2:0]    _zz_1193;
  wire       [1:0]    _zz_1194;
  wire       [1:0]    _zz_1195;
  wire       [0:0]    _zz_1196;
  wire       [1:0]    _zz_1197;
  wire       [0:0]    _zz_1198;
  wire       [1:0]    _zz_1199;
  wire       [1:0]    _zz_1200;
  wire       [2:0]    _zz_1201;
  wire       [1:0]    _zz_1202;
  wire       [3:0]    _zz_1203;
  wire       [2:0]    _zz_1204;
  wire       [3:0]    _zz_1205;
  wire       [2:0]    _zz_1206;
  wire       [1:0]    _zz_1207;
  wire       [0:0]    _zz_1208;
  wire       [1:0]    _zz_1209;
  wire       [0:0]    _zz_1210;
  wire       [1:0]    _zz_1211;
  wire       [2:0]    _zz_1212;
  wire       [1:0]    _zz_1213;
  wire       [2:0]    _zz_1214;
  wire       [1:0]    _zz_1215;
  wire       [1:0]    _zz_1216;
  wire       [0:0]    _zz_1217;
  wire       [1:0]    _zz_1218;
  wire       [0:0]    _zz_1219;
  wire       [1:0]    _zz_1220;
  wire       [1:0]    _zz_1221;
  wire       [2:0]    _zz_1222;
  wire       [1:0]    _zz_1223;
  wire       [2:0]    _zz_1224;
  wire       [3:0]    _zz_1225;
  wire       [2:0]    _zz_1226;
  wire       [4:0]    _zz_1227;
  wire       [3:0]    _zz_1228;
  wire       [4:0]    _zz_1229;
  wire       [3:0]    _zz_1230;
  wire       [1:0]    _zz_1231;
  wire       [0:0]    _zz_1232;
  wire       [1:0]    _zz_1233;
  wire       [0:0]    _zz_1234;
  wire       [1:0]    _zz_1235;
  wire       [2:0]    _zz_1236;
  wire       [1:0]    _zz_1237;
  wire       [2:0]    _zz_1238;
  wire       [1:0]    _zz_1239;
  wire       [1:0]    _zz_1240;
  wire       [0:0]    _zz_1241;
  wire       [1:0]    _zz_1242;
  wire       [0:0]    _zz_1243;
  wire       [1:0]    _zz_1244;
  wire       [1:0]    _zz_1245;
  wire       [2:0]    _zz_1246;
  wire       [1:0]    _zz_1247;
  wire       [3:0]    _zz_1248;
  wire       [2:0]    _zz_1249;
  wire       [3:0]    _zz_1250;
  wire       [2:0]    _zz_1251;
  wire       [1:0]    _zz_1252;
  wire       [0:0]    _zz_1253;
  wire       [1:0]    _zz_1254;
  wire       [0:0]    _zz_1255;
  wire       [1:0]    _zz_1256;
  wire       [2:0]    _zz_1257;
  wire       [1:0]    _zz_1258;
  wire       [2:0]    _zz_1259;
  wire       [1:0]    _zz_1260;
  wire       [1:0]    _zz_1261;
  wire       [0:0]    _zz_1262;
  wire       [1:0]    _zz_1263;
  wire       [0:0]    _zz_1264;
  wire       [1:0]    _zz_1265;
  wire       [1:0]    _zz_1266;
  wire       [2:0]    _zz_1267;
  wire       [1:0]    _zz_1268;
  wire       [2:0]    _zz_1269;
  wire       [3:0]    _zz_1270;
  wire       [2:0]    _zz_1271;
  wire       [3:0]    _zz_1272;
  wire       [4:0]    _zz_1273;
  wire       [3:0]    _zz_1274;
  wire       [4:0]    _zz_1275;
  wire       [5:0]    _zz_1276;
  wire       [4:0]    _zz_1277;
  wire       [6:0]    _zz_1278;
  wire       [5:0]    _zz_1279;
  wire       [6:0]    _zz_1280;
  wire       [5:0]    _zz_1281;
  wire       [1:0]    _zz_1282;
  wire       [0:0]    _zz_1283;
  wire       [1:0]    _zz_1284;
  wire       [0:0]    _zz_1285;
  wire       [1:0]    _zz_1286;
  wire       [2:0]    _zz_1287;
  wire       [1:0]    _zz_1288;
  wire       [2:0]    _zz_1289;
  wire       [1:0]    _zz_1290;
  wire       [1:0]    _zz_1291;
  wire       [0:0]    _zz_1292;
  wire       [1:0]    _zz_1293;
  wire       [0:0]    _zz_1294;
  wire       [1:0]    _zz_1295;
  wire       [1:0]    _zz_1296;
  wire       [2:0]    _zz_1297;
  wire       [1:0]    _zz_1298;
  wire       [3:0]    _zz_1299;
  wire       [2:0]    _zz_1300;
  wire       [3:0]    _zz_1301;
  wire       [2:0]    _zz_1302;
  wire       [1:0]    _zz_1303;
  wire       [0:0]    _zz_1304;
  wire       [1:0]    _zz_1305;
  wire       [0:0]    _zz_1306;
  wire       [1:0]    _zz_1307;
  wire       [2:0]    _zz_1308;
  wire       [1:0]    _zz_1309;
  wire       [2:0]    _zz_1310;
  wire       [1:0]    _zz_1311;
  wire       [1:0]    _zz_1312;
  wire       [0:0]    _zz_1313;
  wire       [1:0]    _zz_1314;
  wire       [0:0]    _zz_1315;
  wire       [1:0]    _zz_1316;
  wire       [1:0]    _zz_1317;
  wire       [2:0]    _zz_1318;
  wire       [1:0]    _zz_1319;
  wire       [2:0]    _zz_1320;
  wire       [3:0]    _zz_1321;
  wire       [2:0]    _zz_1322;
  wire       [4:0]    _zz_1323;
  wire       [3:0]    _zz_1324;
  wire       [4:0]    _zz_1325;
  wire       [3:0]    _zz_1326;
  wire       [1:0]    _zz_1327;
  wire       [0:0]    _zz_1328;
  wire       [1:0]    _zz_1329;
  wire       [0:0]    _zz_1330;
  wire       [1:0]    _zz_1331;
  wire       [2:0]    _zz_1332;
  wire       [1:0]    _zz_1333;
  wire       [2:0]    _zz_1334;
  wire       [1:0]    _zz_1335;
  wire       [1:0]    _zz_1336;
  wire       [0:0]    _zz_1337;
  wire       [1:0]    _zz_1338;
  wire       [0:0]    _zz_1339;
  wire       [1:0]    _zz_1340;
  wire       [1:0]    _zz_1341;
  wire       [2:0]    _zz_1342;
  wire       [1:0]    _zz_1343;
  wire       [3:0]    _zz_1344;
  wire       [2:0]    _zz_1345;
  wire       [3:0]    _zz_1346;
  wire       [2:0]    _zz_1347;
  wire       [1:0]    _zz_1348;
  wire       [0:0]    _zz_1349;
  wire       [1:0]    _zz_1350;
  wire       [0:0]    _zz_1351;
  wire       [1:0]    _zz_1352;
  wire       [2:0]    _zz_1353;
  wire       [1:0]    _zz_1354;
  wire       [2:0]    _zz_1355;
  wire       [1:0]    _zz_1356;
  wire       [1:0]    _zz_1357;
  wire       [0:0]    _zz_1358;
  wire       [1:0]    _zz_1359;
  wire       [0:0]    _zz_1360;
  wire       [1:0]    _zz_1361;
  wire       [1:0]    _zz_1362;
  wire       [2:0]    _zz_1363;
  wire       [1:0]    _zz_1364;
  wire       [2:0]    _zz_1365;
  wire       [3:0]    _zz_1366;
  wire       [2:0]    _zz_1367;
  wire       [3:0]    _zz_1368;
  wire       [4:0]    _zz_1369;
  wire       [3:0]    _zz_1370;
  wire       [5:0]    _zz_1371;
  wire       [4:0]    _zz_1372;
  wire       [5:0]    _zz_1373;
  wire       [4:0]    _zz_1374;
  wire       [1:0]    _zz_1375;
  wire       [0:0]    _zz_1376;
  wire       [1:0]    _zz_1377;
  wire       [0:0]    _zz_1378;
  wire       [1:0]    _zz_1379;
  wire       [2:0]    _zz_1380;
  wire       [1:0]    _zz_1381;
  wire       [2:0]    _zz_1382;
  wire       [1:0]    _zz_1383;
  wire       [1:0]    _zz_1384;
  wire       [0:0]    _zz_1385;
  wire       [1:0]    _zz_1386;
  wire       [0:0]    _zz_1387;
  wire       [1:0]    _zz_1388;
  wire       [1:0]    _zz_1389;
  wire       [2:0]    _zz_1390;
  wire       [1:0]    _zz_1391;
  wire       [3:0]    _zz_1392;
  wire       [2:0]    _zz_1393;
  wire       [3:0]    _zz_1394;
  wire       [2:0]    _zz_1395;
  wire       [1:0]    _zz_1396;
  wire       [0:0]    _zz_1397;
  wire       [1:0]    _zz_1398;
  wire       [0:0]    _zz_1399;
  wire       [1:0]    _zz_1400;
  wire       [2:0]    _zz_1401;
  wire       [1:0]    _zz_1402;
  wire       [2:0]    _zz_1403;
  wire       [1:0]    _zz_1404;
  wire       [1:0]    _zz_1405;
  wire       [0:0]    _zz_1406;
  wire       [1:0]    _zz_1407;
  wire       [0:0]    _zz_1408;
  wire       [1:0]    _zz_1409;
  wire       [1:0]    _zz_1410;
  wire       [2:0]    _zz_1411;
  wire       [1:0]    _zz_1412;
  wire       [2:0]    _zz_1413;
  wire       [3:0]    _zz_1414;
  wire       [2:0]    _zz_1415;
  wire       [4:0]    _zz_1416;
  wire       [3:0]    _zz_1417;
  wire       [4:0]    _zz_1418;
  wire       [3:0]    _zz_1419;
  wire       [1:0]    _zz_1420;
  wire       [0:0]    _zz_1421;
  wire       [1:0]    _zz_1422;
  wire       [0:0]    _zz_1423;
  wire       [1:0]    _zz_1424;
  wire       [2:0]    _zz_1425;
  wire       [1:0]    _zz_1426;
  wire       [2:0]    _zz_1427;
  wire       [1:0]    _zz_1428;
  wire       [1:0]    _zz_1429;
  wire       [0:0]    _zz_1430;
  wire       [1:0]    _zz_1431;
  wire       [0:0]    _zz_1432;
  wire       [1:0]    _zz_1433;
  wire       [1:0]    _zz_1434;
  wire       [2:0]    _zz_1435;
  wire       [1:0]    _zz_1436;
  wire       [3:0]    _zz_1437;
  wire       [2:0]    _zz_1438;
  wire       [3:0]    _zz_1439;
  wire       [2:0]    _zz_1440;
  wire       [1:0]    _zz_1441;
  wire       [0:0]    _zz_1442;
  wire       [1:0]    _zz_1443;
  wire       [0:0]    _zz_1444;
  wire       [1:0]    _zz_1445;
  wire       [2:0]    _zz_1446;
  wire       [1:0]    _zz_1447;
  wire       [2:0]    _zz_1448;
  wire       [1:0]    _zz_1449;
  wire       [1:0]    _zz_1450;
  wire       [0:0]    _zz_1451;
  wire       [1:0]    _zz_1452;
  wire       [0:0]    _zz_1453;
  wire       [1:0]    _zz_1454;
  wire       [1:0]    _zz_1455;
  wire       [2:0]    _zz_1456;
  wire       [1:0]    _zz_1457;
  wire       [2:0]    _zz_1458;
  wire       [3:0]    _zz_1459;
  wire       [2:0]    _zz_1460;
  wire       [3:0]    _zz_1461;
  wire       [4:0]    _zz_1462;
  wire       [3:0]    _zz_1463;
  wire       [4:0]    _zz_1464;
  wire       [5:0]    _zz_1465;
  wire       [4:0]    _zz_1466;
  wire       [5:0]    _zz_1467;
  wire       [6:0]    _zz_1468;
  wire       [5:0]    _zz_1469;
  wire       [6:0]    _zz_1470;
  wire       [7:0]    _zz_1471;
  wire       [6:0]    _zz_1472;
  wire       [7:0]    _zz_1473;
  wire       [7:0]    _zz_1474;
  wire       [15:0]   _zz_1475;
  wire       [7:0]    _zz_1476;
  wire       [15:0]   _zz_1477;
  wire       [7:0]    _zz_1478;
  wire       [7:0]    _zz_1479;
  wire       [7:0]    _zz_1480;
  wire       [7:0]    _zz_1481;
  wire       [7:0]    _zz_1482;
  wire       [7:0]    _zz_1483;
  wire       [15:0]   _zz_1484;
  wire       [15:0]   _zz_1485;
  wire       [15:0]   _zz_1486;
  wire       [15:0]   _zz_1487;
  wire       [15:0]   _zz_1488;
  wire       [15:0]   _zz_1489;
  wire       [15:0]   _zz_1490;
  wire       [15:0]   _zz_1491;
  wire       [15:0]   _zz_1492;
  wire       [15:0]   _zz_1493;
  wire       [15:0]   _zz_1494;
  wire       [15:0]   _zz_1495;
  wire       [15:0]   _zz_1496;
  wire       [23:0]   _zz_1497;
  wire       [31:0]   _zz_1498;
  wire       [15:0]   _zz_1499;
  wire       [15:0]   _zz_1500;
  wire       [15:0]   _zz_1501;
  wire       [23:0]   _zz_1502;
  wire       [31:0]   _zz_1503;
  wire       [23:0]   _zz_1504;
  wire       [31:0]   _zz_1505;
  wire       [15:0]   _zz_1506;
  wire       [15:0]   _zz_1507;
  wire       [15:0]   _zz_1508;
  wire       [23:0]   _zz_1509;
  wire       [31:0]   _zz_1510;
  wire       [23:0]   _zz_1511;
  wire       [23:0]   _zz_1512;
  wire       [23:0]   _zz_1513;
  wire       [23:0]   _zz_1514;
  wire       [15:0]   _zz_1515;
  wire       [15:0]   _zz_1516;
  wire       [15:0]   _zz_1517;
  wire       [15:0]   _zz_1518;
  wire       [23:0]   _zz_1519;
  wire       [15:0]   _zz_1520;
  wire       [23:0]   _zz_1521;
  wire       [15:0]   _zz_1522;
  wire       [31:0]   _zz_1523;
  wire       [31:0]   _zz_1524;
  wire       [31:0]   _zz_1525;
  wire       [31:0]   _zz_1526;
  wire       [31:0]   _zz_1527;
  wire       [31:0]   _zz_1528;
  wire       [31:0]   _zz_1529;
  wire       [31:0]   _zz_1530;
  wire       [31:0]   _zz_1531;
  wire       [31:0]   _zz_1532;
  wire       [31:0]   _zz_1533;
  wire       [31:0]   _zz_1534;
  wire       [31:0]   _zz_1535;
  wire       [47:0]   _zz_1536;
  wire       [31:0]   _zz_1537;
  wire       [31:0]   _zz_1538;
  wire       [31:0]   _zz_1539;
  wire       [47:0]   _zz_1540;
  wire       [31:0]   _zz_1541;
  wire       [31:0]   _zz_1542;
  wire       [31:0]   _zz_1543;
  wire       [15:0]   _zz_1544;
  wire       [15:0]   _zz_1545;
  wire       [15:0]   func_table_0_real;
  wire       [15:0]   func_table_0_imag;
  wire       [15:0]   func_table_1_real;
  wire       [15:0]   func_table_1_imag;
  wire       [15:0]   func_table_2_real;
  wire       [15:0]   func_table_2_imag;
  wire       [15:0]   func_table_3_real;
  wire       [15:0]   func_table_3_imag;
  wire       [15:0]   func_table_4_real;
  wire       [15:0]   func_table_4_imag;
  wire       [15:0]   func_table_5_real;
  wire       [15:0]   func_table_5_imag;
  wire       [15:0]   func_table_6_real;
  wire       [15:0]   func_table_6_imag;
  wire       [15:0]   func_table_7_real;
  wire       [15:0]   func_table_7_imag;
  wire       [15:0]   func_table_8_real;
  wire       [15:0]   func_table_8_imag;
  wire       [15:0]   func_table_9_real;
  wire       [15:0]   func_table_9_imag;
  wire       [15:0]   func_table_10_real;
  wire       [15:0]   func_table_10_imag;
  wire       [15:0]   func_table_11_real;
  wire       [15:0]   func_table_11_imag;
  wire       [15:0]   func_table_12_real;
  wire       [15:0]   func_table_12_imag;
  wire       [15:0]   func_table_13_real;
  wire       [15:0]   func_table_13_imag;
  wire       [15:0]   func_table_14_real;
  wire       [15:0]   func_table_14_imag;
  wire       [15:0]   func_table_15_real;
  wire       [15:0]   func_table_15_imag;
  wire       [15:0]   func_table_16_real;
  wire       [15:0]   func_table_16_imag;
  wire       [15:0]   func_table_17_real;
  wire       [15:0]   func_table_17_imag;
  wire       [15:0]   func_table_18_real;
  wire       [15:0]   func_table_18_imag;
  wire       [15:0]   func_table_19_real;
  wire       [15:0]   func_table_19_imag;
  wire       [15:0]   func_table_20_real;
  wire       [15:0]   func_table_20_imag;
  wire       [15:0]   func_table_21_real;
  wire       [15:0]   func_table_21_imag;
  wire       [15:0]   func_table_22_real;
  wire       [15:0]   func_table_22_imag;
  wire       [15:0]   func_table_23_real;
  wire       [15:0]   func_table_23_imag;
  wire       [15:0]   func_table_24_real;
  wire       [15:0]   func_table_24_imag;
  wire       [15:0]   func_table_25_real;
  wire       [15:0]   func_table_25_imag;
  wire       [15:0]   func_table_26_real;
  wire       [15:0]   func_table_26_imag;
  wire       [15:0]   func_table_27_real;
  wire       [15:0]   func_table_27_imag;
  wire       [15:0]   func_table_28_real;
  wire       [15:0]   func_table_28_imag;
  wire       [15:0]   func_table_29_real;
  wire       [15:0]   func_table_29_imag;
  wire       [15:0]   func_table_30_real;
  wire       [15:0]   func_table_30_imag;
  wire       [15:0]   func_table_31_real;
  wire       [15:0]   func_table_31_imag;
  wire       [15:0]   func_table_32_real;
  wire       [15:0]   func_table_32_imag;
  wire       [15:0]   func_table_33_real;
  wire       [15:0]   func_table_33_imag;
  wire       [15:0]   func_table_34_real;
  wire       [15:0]   func_table_34_imag;
  wire       [15:0]   func_table_35_real;
  wire       [15:0]   func_table_35_imag;
  wire       [15:0]   func_table_36_real;
  wire       [15:0]   func_table_36_imag;
  wire       [15:0]   func_table_37_real;
  wire       [15:0]   func_table_37_imag;
  wire       [15:0]   func_table_38_real;
  wire       [15:0]   func_table_38_imag;
  wire       [15:0]   func_table_39_real;
  wire       [15:0]   func_table_39_imag;
  wire       [15:0]   func_table_40_real;
  wire       [15:0]   func_table_40_imag;
  wire       [15:0]   func_table_41_real;
  wire       [15:0]   func_table_41_imag;
  wire       [15:0]   func_table_42_real;
  wire       [15:0]   func_table_42_imag;
  wire       [15:0]   func_table_43_real;
  wire       [15:0]   func_table_43_imag;
  wire       [15:0]   func_table_44_real;
  wire       [15:0]   func_table_44_imag;
  wire       [15:0]   func_table_45_real;
  wire       [15:0]   func_table_45_imag;
  wire       [15:0]   func_table_46_real;
  wire       [15:0]   func_table_46_imag;
  wire       [15:0]   func_table_47_real;
  wire       [15:0]   func_table_47_imag;
  wire       [15:0]   func_table_48_real;
  wire       [15:0]   func_table_48_imag;
  wire       [15:0]   func_table_49_real;
  wire       [15:0]   func_table_49_imag;
  wire       [15:0]   func_table_50_real;
  wire       [15:0]   func_table_50_imag;
  wire       [15:0]   func_table_51_real;
  wire       [15:0]   func_table_51_imag;
  wire       [15:0]   func_table_52_real;
  wire       [15:0]   func_table_52_imag;
  wire       [15:0]   func_table_53_real;
  wire       [15:0]   func_table_53_imag;
  wire       [15:0]   func_table_54_real;
  wire       [15:0]   func_table_54_imag;
  wire       [15:0]   func_table_55_real;
  wire       [15:0]   func_table_55_imag;
  wire       [15:0]   func_table_56_real;
  wire       [15:0]   func_table_56_imag;
  wire       [15:0]   func_table_57_real;
  wire       [15:0]   func_table_57_imag;
  wire       [15:0]   func_table_58_real;
  wire       [15:0]   func_table_58_imag;
  wire       [15:0]   func_table_59_real;
  wire       [15:0]   func_table_59_imag;
  wire       [15:0]   func_table_60_real;
  wire       [15:0]   func_table_60_imag;
  wire       [15:0]   func_table_61_real;
  wire       [15:0]   func_table_61_imag;
  wire       [15:0]   func_table_62_real;
  wire       [15:0]   func_table_62_imag;
  wire       [15:0]   func_table_63_real;
  wire       [15:0]   func_table_63_imag;
  wire       [15:0]   func_table_64_real;
  wire       [15:0]   func_table_64_imag;
  wire       [15:0]   func_table_65_real;
  wire       [15:0]   func_table_65_imag;
  wire       [15:0]   func_table_66_real;
  wire       [15:0]   func_table_66_imag;
  wire       [15:0]   func_table_67_real;
  wire       [15:0]   func_table_67_imag;
  wire       [15:0]   func_table_68_real;
  wire       [15:0]   func_table_68_imag;
  wire       [15:0]   func_table_69_real;
  wire       [15:0]   func_table_69_imag;
  wire       [15:0]   func_table_70_real;
  wire       [15:0]   func_table_70_imag;
  wire       [15:0]   func_table_71_real;
  wire       [15:0]   func_table_71_imag;
  wire       [15:0]   func_table_72_real;
  wire       [15:0]   func_table_72_imag;
  wire       [15:0]   func_table_73_real;
  wire       [15:0]   func_table_73_imag;
  wire       [15:0]   func_table_74_real;
  wire       [15:0]   func_table_74_imag;
  wire       [15:0]   func_table_75_real;
  wire       [15:0]   func_table_75_imag;
  wire       [15:0]   func_table_76_real;
  wire       [15:0]   func_table_76_imag;
  wire       [15:0]   func_table_77_real;
  wire       [15:0]   func_table_77_imag;
  wire       [15:0]   func_table_78_real;
  wire       [15:0]   func_table_78_imag;
  wire       [15:0]   func_table_79_real;
  wire       [15:0]   func_table_79_imag;
  wire       [15:0]   func_table_80_real;
  wire       [15:0]   func_table_80_imag;
  wire       [15:0]   func_table_81_real;
  wire       [15:0]   func_table_81_imag;
  wire       [15:0]   func_table_82_real;
  wire       [15:0]   func_table_82_imag;
  wire       [15:0]   func_table_83_real;
  wire       [15:0]   func_table_83_imag;
  wire       [15:0]   func_table_84_real;
  wire       [15:0]   func_table_84_imag;
  wire       [15:0]   func_table_85_real;
  wire       [15:0]   func_table_85_imag;
  wire       [15:0]   func_table_86_real;
  wire       [15:0]   func_table_86_imag;
  wire       [15:0]   func_table_87_real;
  wire       [15:0]   func_table_87_imag;
  wire       [15:0]   func_table_88_real;
  wire       [15:0]   func_table_88_imag;
  wire       [15:0]   func_table_89_real;
  wire       [15:0]   func_table_89_imag;
  wire       [15:0]   func_table_90_real;
  wire       [15:0]   func_table_90_imag;
  wire       [15:0]   func_table_91_real;
  wire       [15:0]   func_table_91_imag;
  wire       [15:0]   func_table_92_real;
  wire       [15:0]   func_table_92_imag;
  wire       [15:0]   func_table_93_real;
  wire       [15:0]   func_table_93_imag;
  wire       [15:0]   func_table_94_real;
  wire       [15:0]   func_table_94_imag;
  wire       [15:0]   func_table_95_real;
  wire       [15:0]   func_table_95_imag;
  wire       [15:0]   func_table_96_real;
  wire       [15:0]   func_table_96_imag;
  wire       [15:0]   func_table_97_real;
  wire       [15:0]   func_table_97_imag;
  wire       [15:0]   func_table_98_real;
  wire       [15:0]   func_table_98_imag;
  wire       [15:0]   func_table_99_real;
  wire       [15:0]   func_table_99_imag;
  wire       [15:0]   func_table_100_real;
  wire       [15:0]   func_table_100_imag;
  wire       [15:0]   func_table_101_real;
  wire       [15:0]   func_table_101_imag;
  wire       [15:0]   func_table_102_real;
  wire       [15:0]   func_table_102_imag;
  wire       [15:0]   func_table_103_real;
  wire       [15:0]   func_table_103_imag;
  wire       [15:0]   func_table_104_real;
  wire       [15:0]   func_table_104_imag;
  wire       [15:0]   func_table_105_real;
  wire       [15:0]   func_table_105_imag;
  wire       [15:0]   func_table_106_real;
  wire       [15:0]   func_table_106_imag;
  wire       [15:0]   func_table_107_real;
  wire       [15:0]   func_table_107_imag;
  wire       [15:0]   func_table_108_real;
  wire       [15:0]   func_table_108_imag;
  wire       [15:0]   func_table_109_real;
  wire       [15:0]   func_table_109_imag;
  wire       [15:0]   func_table_110_real;
  wire       [15:0]   func_table_110_imag;
  wire       [15:0]   func_table_111_real;
  wire       [15:0]   func_table_111_imag;
  wire       [15:0]   func_table_112_real;
  wire       [15:0]   func_table_112_imag;
  wire       [15:0]   func_table_113_real;
  wire       [15:0]   func_table_113_imag;
  wire       [15:0]   func_table_114_real;
  wire       [15:0]   func_table_114_imag;
  wire       [15:0]   func_table_115_real;
  wire       [15:0]   func_table_115_imag;
  wire       [15:0]   func_table_116_real;
  wire       [15:0]   func_table_116_imag;
  wire       [15:0]   func_table_117_real;
  wire       [15:0]   func_table_117_imag;
  wire       [15:0]   func_table_118_real;
  wire       [15:0]   func_table_118_imag;
  wire       [15:0]   func_table_119_real;
  wire       [15:0]   func_table_119_imag;
  wire       [15:0]   func_table_120_real;
  wire       [15:0]   func_table_120_imag;
  wire       [15:0]   func_table_121_real;
  wire       [15:0]   func_table_121_imag;
  wire       [15:0]   func_table_122_real;
  wire       [15:0]   func_table_122_imag;
  wire       [15:0]   func_table_123_real;
  wire       [15:0]   func_table_123_imag;
  wire       [15:0]   func_table_124_real;
  wire       [15:0]   func_table_124_imag;
  wire       [15:0]   func_table_125_real;
  wire       [15:0]   func_table_125_imag;
  wire       [15:0]   func_table_126_real;
  wire       [15:0]   func_table_126_imag;
  wire       [15:0]   func_table_127_real;
  wire       [15:0]   func_table_127_imag;
  reg        [15:0]   wave;
  reg        [15:0]   distance;
  wire       [15:0]   timeshift_real;
  wire       [15:0]   timeshift_imag;
  reg        [15:0]   io_timeshift_regNext_real;
  reg        [15:0]   io_timeshift_regNext_imag;
  reg        [15:0]   _zz_1;
  reg        [15:0]   _zz_2;
  reg        [15:0]   _zz_3;
  reg        [15:0]   _zz_4;
  reg        [15:0]   _zz_5;
  reg        [15:0]   _zz_6;
  reg        [15:0]   _zz_7;
  reg        [15:0]   _zz_8;
  reg        [31:0]   _zz_9;
  wire       [7:0]    wd_prod;
  wire       [15:0]   indx_table_0;
  wire       [15:0]   indx_table_1;
  wire       [15:0]   indx_table_2;
  wire       [15:0]   indx_table_3;
  wire       [15:0]   indx_table_4;
  wire       [15:0]   indx_table_5;
  wire       [15:0]   indx_table_6;
  wire       [15:0]   indx_table_7;
  wire       [15:0]   indx_table_8;
  wire       [15:0]   indx_table_9;
  wire       [15:0]   indx_table_10;
  wire       [15:0]   indx_table_11;
  wire       [15:0]   indx_table_12;
  wire       [15:0]   indx_table_13;
  wire       [15:0]   indx_table_14;
  wire       [15:0]   indx_table_15;
  wire       [15:0]   indx_table_16;
  wire       [15:0]   indx_table_17;
  wire       [15:0]   indx_table_18;
  wire       [15:0]   indx_table_19;
  wire       [15:0]   indx_table_20;
  wire       [15:0]   indx_table_21;
  wire       [15:0]   indx_table_22;
  wire       [15:0]   indx_table_23;
  wire       [15:0]   indx_table_24;
  wire       [15:0]   indx_table_25;
  wire       [15:0]   indx_table_26;
  wire       [15:0]   indx_table_27;
  wire       [15:0]   indx_table_28;
  wire       [15:0]   indx_table_29;
  wire       [15:0]   indx_table_30;
  wire       [15:0]   indx_table_31;
  wire       [15:0]   indx_table_32;
  wire       [15:0]   indx_table_33;
  wire       [15:0]   indx_table_34;
  wire       [15:0]   indx_table_35;
  wire       [15:0]   indx_table_36;
  wire       [15:0]   indx_table_37;
  wire       [15:0]   indx_table_38;
  wire       [15:0]   indx_table_39;
  wire       [15:0]   indx_table_40;
  wire       [15:0]   indx_table_41;
  wire       [15:0]   indx_table_42;
  wire       [15:0]   indx_table_43;
  wire       [15:0]   indx_table_44;
  wire       [15:0]   indx_table_45;
  wire       [15:0]   indx_table_46;
  wire       [15:0]   indx_table_47;
  wire       [15:0]   indx_table_48;
  wire       [15:0]   indx_table_49;
  wire       [15:0]   indx_table_50;
  wire       [15:0]   indx_table_51;
  wire       [15:0]   indx_table_52;
  wire       [15:0]   indx_table_53;
  wire       [15:0]   indx_table_54;
  wire       [15:0]   indx_table_55;
  wire       [15:0]   indx_table_56;
  wire       [15:0]   indx_table_57;
  wire       [15:0]   indx_table_58;
  wire       [15:0]   indx_table_59;
  wire       [15:0]   indx_table_60;
  wire       [15:0]   indx_table_61;
  wire       [15:0]   indx_table_62;
  wire       [15:0]   indx_table_63;
  wire       [15:0]   indx_table_64;
  wire       [15:0]   indx_table_65;
  wire       [15:0]   indx_table_66;
  wire       [15:0]   indx_table_67;
  wire       [15:0]   indx_table_68;
  wire       [15:0]   indx_table_69;
  wire       [15:0]   indx_table_70;
  wire       [15:0]   indx_table_71;
  wire       [15:0]   indx_table_72;
  wire       [15:0]   indx_table_73;
  wire       [15:0]   indx_table_74;
  wire       [15:0]   indx_table_75;
  wire       [15:0]   indx_table_76;
  wire       [15:0]   indx_table_77;
  wire       [15:0]   indx_table_78;
  wire       [15:0]   indx_table_79;
  wire       [15:0]   indx_table_80;
  wire       [15:0]   indx_table_81;
  wire       [15:0]   indx_table_82;
  wire       [15:0]   indx_table_83;
  wire       [15:0]   indx_table_84;
  wire       [15:0]   indx_table_85;
  wire       [15:0]   indx_table_86;
  wire       [15:0]   indx_table_87;
  wire       [15:0]   indx_table_88;
  wire       [15:0]   indx_table_89;
  wire       [15:0]   indx_table_90;
  wire       [15:0]   indx_table_91;
  wire       [15:0]   indx_table_92;
  wire       [15:0]   indx_table_93;
  wire       [15:0]   indx_table_94;
  wire       [15:0]   indx_table_95;
  wire       [15:0]   indx_table_96;
  wire       [15:0]   indx_table_97;
  wire       [15:0]   indx_table_98;
  wire       [15:0]   indx_table_99;
  wire       [15:0]   indx_table_100;
  wire       [15:0]   indx_table_101;
  wire       [15:0]   indx_table_102;
  wire       [15:0]   indx_table_103;
  wire       [15:0]   indx_table_104;
  wire       [15:0]   indx_table_105;
  wire       [15:0]   indx_table_106;
  wire       [15:0]   indx_table_107;
  wire       [15:0]   indx_table_108;
  wire       [15:0]   indx_table_109;
  wire       [15:0]   indx_table_110;
  wire       [15:0]   indx_table_111;
  wire       [15:0]   indx_table_112;
  wire       [15:0]   indx_table_113;
  wire       [15:0]   indx_table_114;
  wire       [15:0]   indx_table_115;
  wire       [15:0]   indx_table_116;
  wire       [15:0]   indx_table_117;
  wire       [15:0]   indx_table_118;
  wire       [15:0]   indx_table_119;
  wire       [15:0]   indx_table_120;
  wire       [15:0]   indx_table_121;
  wire       [15:0]   indx_table_122;
  wire       [15:0]   indx_table_123;
  wire       [15:0]   indx_table_124;
  wire       [15:0]   indx_table_125;
  wire       [15:0]   indx_table_126;
  wire       [15:0]   indx_table_127;
  wire                idx_comp_0;
  wire                idx_comp_1;
  wire                idx_comp_2;
  wire                idx_comp_3;
  wire                idx_comp_4;
  wire                idx_comp_5;
  wire                idx_comp_6;
  wire                idx_comp_7;
  wire                idx_comp_8;
  wire                idx_comp_9;
  wire                idx_comp_10;
  wire                idx_comp_11;
  wire                idx_comp_12;
  wire                idx_comp_13;
  wire                idx_comp_14;
  wire                idx_comp_15;
  wire                idx_comp_16;
  wire                idx_comp_17;
  wire                idx_comp_18;
  wire                idx_comp_19;
  wire                idx_comp_20;
  wire                idx_comp_21;
  wire                idx_comp_22;
  wire                idx_comp_23;
  wire                idx_comp_24;
  wire                idx_comp_25;
  wire                idx_comp_26;
  wire                idx_comp_27;
  wire                idx_comp_28;
  wire                idx_comp_29;
  wire                idx_comp_30;
  wire                idx_comp_31;
  wire                idx_comp_32;
  wire                idx_comp_33;
  wire                idx_comp_34;
  wire                idx_comp_35;
  wire                idx_comp_36;
  wire                idx_comp_37;
  wire                idx_comp_38;
  wire                idx_comp_39;
  wire                idx_comp_40;
  wire                idx_comp_41;
  wire                idx_comp_42;
  wire                idx_comp_43;
  wire                idx_comp_44;
  wire                idx_comp_45;
  wire                idx_comp_46;
  wire                idx_comp_47;
  wire                idx_comp_48;
  wire                idx_comp_49;
  wire                idx_comp_50;
  wire                idx_comp_51;
  wire                idx_comp_52;
  wire                idx_comp_53;
  wire                idx_comp_54;
  wire                idx_comp_55;
  wire                idx_comp_56;
  wire                idx_comp_57;
  wire                idx_comp_58;
  wire                idx_comp_59;
  wire                idx_comp_60;
  wire                idx_comp_61;
  wire                idx_comp_62;
  wire                idx_comp_63;
  wire                idx_comp_64;
  wire                idx_comp_65;
  wire                idx_comp_66;
  wire                idx_comp_67;
  wire                idx_comp_68;
  wire                idx_comp_69;
  wire                idx_comp_70;
  wire                idx_comp_71;
  wire                idx_comp_72;
  wire                idx_comp_73;
  wire                idx_comp_74;
  wire                idx_comp_75;
  wire                idx_comp_76;
  wire                idx_comp_77;
  wire                idx_comp_78;
  wire                idx_comp_79;
  wire                idx_comp_80;
  wire                idx_comp_81;
  wire                idx_comp_82;
  wire                idx_comp_83;
  wire                idx_comp_84;
  wire                idx_comp_85;
  wire                idx_comp_86;
  wire                idx_comp_87;
  wire                idx_comp_88;
  wire                idx_comp_89;
  wire                idx_comp_90;
  wire                idx_comp_91;
  wire                idx_comp_92;
  wire                idx_comp_93;
  wire                idx_comp_94;
  wire                idx_comp_95;
  wire                idx_comp_96;
  wire                idx_comp_97;
  wire                idx_comp_98;
  wire                idx_comp_99;
  wire                idx_comp_100;
  wire                idx_comp_101;
  wire                idx_comp_102;
  wire                idx_comp_103;
  wire                idx_comp_104;
  wire                idx_comp_105;
  wire                idx_comp_106;
  wire                idx_comp_107;
  wire                idx_comp_108;
  wire                idx_comp_109;
  wire                idx_comp_110;
  wire                idx_comp_111;
  wire                idx_comp_112;
  wire                idx_comp_113;
  wire                idx_comp_114;
  wire                idx_comp_115;
  wire                idx_comp_116;
  wire                idx_comp_117;
  wire                idx_comp_118;
  wire                idx_comp_119;
  wire                idx_comp_120;
  wire                idx_comp_121;
  wire                idx_comp_122;
  wire                idx_comp_123;
  wire                idx_comp_124;
  wire                idx_comp_125;
  wire                idx_comp_126;
  wire                idx_comp_127;
  reg        [127:0]  _zz_10;
  wire       [127:0]  _zz_11;
  wire       [7:0]    all_zeros;
  wire       [7:0]    all_left_zeros;
  wire       [7:0]    whole_bit_count;
  wire       [7:0]    left_bit_count;
  wire       [63:0]   _zz_12;
  wire       [6:0]    all_zeros_1;
  wire       [6:0]    all_left_zeros_1;
  wire       [6:0]    whole_bit_count_1;
  wire       [6:0]    left_bit_count_1;
  wire       [31:0]   _zz_13;
  wire       [5:0]    all_zeros_2;
  wire       [5:0]    all_left_zeros_2;
  wire       [5:0]    whole_bit_count_2;
  wire       [5:0]    left_bit_count_2;
  wire       [15:0]   _zz_14;
  wire       [4:0]    all_zeros_3;
  wire       [4:0]    all_left_zeros_3;
  wire       [4:0]    whole_bit_count_3;
  wire       [4:0]    left_bit_count_3;
  wire       [7:0]    _zz_15;
  wire       [3:0]    all_zeros_4;
  wire       [3:0]    all_left_zeros_4;
  wire       [3:0]    whole_bit_count_4;
  wire       [3:0]    left_bit_count_4;
  wire       [3:0]    _zz_16;
  wire       [2:0]    all_zeros_5;
  wire       [2:0]    all_left_zeros_5;
  wire       [2:0]    whole_bit_count_5;
  wire       [2:0]    left_bit_count_5;
  wire       [1:0]    _zz_17;
  wire       [1:0]    all_zeros_6;
  wire       [1:0]    all_left_zeros_6;
  wire       [1:0]    whole_bit_count_6;
  wire       [1:0]    left_bit_count_6;
  wire       [0:0]    _zz_18;
  wire       [0:0]    _zz_19;
  wire       [0:0]    all_zeros_7;
  wire       [0:0]    all_left_zeros_7;
  wire       [1:0]    left_all_zeros_count;
  wire       [0:0]    _zz_20;
  wire       [0:0]    _zz_21;
  wire       [0:0]    all_zeros_8;
  wire       [0:0]    all_left_zeros_8;
  wire       [1:0]    left_non_all_zeros_count;
  wire       [1:0]    non_zeros_lzc;
  wire       [2:0]    left_all_zeros_count_1;
  wire       [1:0]    _zz_22;
  wire       [1:0]    all_zeros_9;
  wire       [1:0]    all_left_zeros_9;
  wire       [1:0]    whole_bit_count_7;
  wire       [1:0]    left_bit_count_7;
  wire       [0:0]    _zz_23;
  wire       [0:0]    _zz_24;
  wire       [0:0]    all_zeros_10;
  wire       [0:0]    all_left_zeros_10;
  wire       [1:0]    left_all_zeros_count_2;
  wire       [0:0]    _zz_25;
  wire       [0:0]    _zz_26;
  wire       [0:0]    all_zeros_11;
  wire       [0:0]    all_left_zeros_11;
  wire       [1:0]    left_non_all_zeros_count_1;
  wire       [1:0]    non_zeros_lzc_1;
  wire       [2:0]    left_non_all_zeros_count_2;
  wire       [2:0]    non_zeros_lzc_2;
  wire       [3:0]    left_all_zeros_count_3;
  wire       [3:0]    _zz_27;
  wire       [2:0]    all_zeros_12;
  wire       [2:0]    all_left_zeros_12;
  wire       [2:0]    whole_bit_count_8;
  wire       [2:0]    left_bit_count_8;
  wire       [1:0]    _zz_28;
  wire       [1:0]    all_zeros_13;
  wire       [1:0]    all_left_zeros_13;
  wire       [1:0]    whole_bit_count_9;
  wire       [1:0]    left_bit_count_9;
  wire       [0:0]    _zz_29;
  wire       [0:0]    _zz_30;
  wire       [0:0]    all_zeros_14;
  wire       [0:0]    all_left_zeros_14;
  wire       [1:0]    left_all_zeros_count_4;
  wire       [0:0]    _zz_31;
  wire       [0:0]    _zz_32;
  wire       [0:0]    all_zeros_15;
  wire       [0:0]    all_left_zeros_15;
  wire       [1:0]    left_non_all_zeros_count_3;
  wire       [1:0]    non_zeros_lzc_3;
  wire       [2:0]    left_all_zeros_count_5;
  wire       [1:0]    _zz_33;
  wire       [1:0]    all_zeros_16;
  wire       [1:0]    all_left_zeros_16;
  wire       [1:0]    whole_bit_count_10;
  wire       [1:0]    left_bit_count_10;
  wire       [0:0]    _zz_34;
  wire       [0:0]    _zz_35;
  wire       [0:0]    all_zeros_17;
  wire       [0:0]    all_left_zeros_17;
  wire       [1:0]    left_all_zeros_count_6;
  wire       [0:0]    _zz_36;
  wire       [0:0]    _zz_37;
  wire       [0:0]    all_zeros_18;
  wire       [0:0]    all_left_zeros_18;
  wire       [1:0]    left_non_all_zeros_count_4;
  wire       [1:0]    non_zeros_lzc_4;
  wire       [2:0]    left_non_all_zeros_count_5;
  wire       [2:0]    non_zeros_lzc_5;
  wire       [3:0]    left_non_all_zeros_count_6;
  wire       [3:0]    non_zeros_lzc_6;
  wire       [4:0]    left_all_zeros_count_7;
  wire       [7:0]    _zz_38;
  wire       [3:0]    all_zeros_19;
  wire       [3:0]    all_left_zeros_19;
  wire       [3:0]    whole_bit_count_11;
  wire       [3:0]    left_bit_count_11;
  wire       [3:0]    _zz_39;
  wire       [2:0]    all_zeros_20;
  wire       [2:0]    all_left_zeros_20;
  wire       [2:0]    whole_bit_count_12;
  wire       [2:0]    left_bit_count_12;
  wire       [1:0]    _zz_40;
  wire       [1:0]    all_zeros_21;
  wire       [1:0]    all_left_zeros_21;
  wire       [1:0]    whole_bit_count_13;
  wire       [1:0]    left_bit_count_13;
  wire       [0:0]    _zz_41;
  wire       [0:0]    _zz_42;
  wire       [0:0]    all_zeros_22;
  wire       [0:0]    all_left_zeros_22;
  wire       [1:0]    left_all_zeros_count_8;
  wire       [0:0]    _zz_43;
  wire       [0:0]    _zz_44;
  wire       [0:0]    all_zeros_23;
  wire       [0:0]    all_left_zeros_23;
  wire       [1:0]    left_non_all_zeros_count_7;
  wire       [1:0]    non_zeros_lzc_7;
  wire       [2:0]    left_all_zeros_count_9;
  wire       [1:0]    _zz_45;
  wire       [1:0]    all_zeros_24;
  wire       [1:0]    all_left_zeros_24;
  wire       [1:0]    whole_bit_count_14;
  wire       [1:0]    left_bit_count_14;
  wire       [0:0]    _zz_46;
  wire       [0:0]    _zz_47;
  wire       [0:0]    all_zeros_25;
  wire       [0:0]    all_left_zeros_25;
  wire       [1:0]    left_all_zeros_count_10;
  wire       [0:0]    _zz_48;
  wire       [0:0]    _zz_49;
  wire       [0:0]    all_zeros_26;
  wire       [0:0]    all_left_zeros_26;
  wire       [1:0]    left_non_all_zeros_count_8;
  wire       [1:0]    non_zeros_lzc_8;
  wire       [2:0]    left_non_all_zeros_count_9;
  wire       [2:0]    non_zeros_lzc_9;
  wire       [3:0]    left_all_zeros_count_11;
  wire       [3:0]    _zz_50;
  wire       [2:0]    all_zeros_27;
  wire       [2:0]    all_left_zeros_27;
  wire       [2:0]    whole_bit_count_15;
  wire       [2:0]    left_bit_count_15;
  wire       [1:0]    _zz_51;
  wire       [1:0]    all_zeros_28;
  wire       [1:0]    all_left_zeros_28;
  wire       [1:0]    whole_bit_count_16;
  wire       [1:0]    left_bit_count_16;
  wire       [0:0]    _zz_52;
  wire       [0:0]    _zz_53;
  wire       [0:0]    all_zeros_29;
  wire       [0:0]    all_left_zeros_29;
  wire       [1:0]    left_all_zeros_count_12;
  wire       [0:0]    _zz_54;
  wire       [0:0]    _zz_55;
  wire       [0:0]    all_zeros_30;
  wire       [0:0]    all_left_zeros_30;
  wire       [1:0]    left_non_all_zeros_count_10;
  wire       [1:0]    non_zeros_lzc_10;
  wire       [2:0]    left_all_zeros_count_13;
  wire       [1:0]    _zz_56;
  wire       [1:0]    all_zeros_31;
  wire       [1:0]    all_left_zeros_31;
  wire       [1:0]    whole_bit_count_17;
  wire       [1:0]    left_bit_count_17;
  wire       [0:0]    _zz_57;
  wire       [0:0]    _zz_58;
  wire       [0:0]    all_zeros_32;
  wire       [0:0]    all_left_zeros_32;
  wire       [1:0]    left_all_zeros_count_14;
  wire       [0:0]    _zz_59;
  wire       [0:0]    _zz_60;
  wire       [0:0]    all_zeros_33;
  wire       [0:0]    all_left_zeros_33;
  wire       [1:0]    left_non_all_zeros_count_11;
  wire       [1:0]    non_zeros_lzc_11;
  wire       [2:0]    left_non_all_zeros_count_12;
  wire       [2:0]    non_zeros_lzc_12;
  wire       [3:0]    left_non_all_zeros_count_13;
  wire       [3:0]    non_zeros_lzc_13;
  wire       [4:0]    left_non_all_zeros_count_14;
  wire       [4:0]    non_zeros_lzc_14;
  wire       [5:0]    left_all_zeros_count_15;
  wire       [15:0]   _zz_61;
  wire       [4:0]    all_zeros_34;
  wire       [4:0]    all_left_zeros_34;
  wire       [4:0]    whole_bit_count_18;
  wire       [4:0]    left_bit_count_18;
  wire       [7:0]    _zz_62;
  wire       [3:0]    all_zeros_35;
  wire       [3:0]    all_left_zeros_35;
  wire       [3:0]    whole_bit_count_19;
  wire       [3:0]    left_bit_count_19;
  wire       [3:0]    _zz_63;
  wire       [2:0]    all_zeros_36;
  wire       [2:0]    all_left_zeros_36;
  wire       [2:0]    whole_bit_count_20;
  wire       [2:0]    left_bit_count_20;
  wire       [1:0]    _zz_64;
  wire       [1:0]    all_zeros_37;
  wire       [1:0]    all_left_zeros_37;
  wire       [1:0]    whole_bit_count_21;
  wire       [1:0]    left_bit_count_21;
  wire       [0:0]    _zz_65;
  wire       [0:0]    _zz_66;
  wire       [0:0]    all_zeros_38;
  wire       [0:0]    all_left_zeros_38;
  wire       [1:0]    left_all_zeros_count_16;
  wire       [0:0]    _zz_67;
  wire       [0:0]    _zz_68;
  wire       [0:0]    all_zeros_39;
  wire       [0:0]    all_left_zeros_39;
  wire       [1:0]    left_non_all_zeros_count_15;
  wire       [1:0]    non_zeros_lzc_15;
  wire       [2:0]    left_all_zeros_count_17;
  wire       [1:0]    _zz_69;
  wire       [1:0]    all_zeros_40;
  wire       [1:0]    all_left_zeros_40;
  wire       [1:0]    whole_bit_count_22;
  wire       [1:0]    left_bit_count_22;
  wire       [0:0]    _zz_70;
  wire       [0:0]    _zz_71;
  wire       [0:0]    all_zeros_41;
  wire       [0:0]    all_left_zeros_41;
  wire       [1:0]    left_all_zeros_count_18;
  wire       [0:0]    _zz_72;
  wire       [0:0]    _zz_73;
  wire       [0:0]    all_zeros_42;
  wire       [0:0]    all_left_zeros_42;
  wire       [1:0]    left_non_all_zeros_count_16;
  wire       [1:0]    non_zeros_lzc_16;
  wire       [2:0]    left_non_all_zeros_count_17;
  wire       [2:0]    non_zeros_lzc_17;
  wire       [3:0]    left_all_zeros_count_19;
  wire       [3:0]    _zz_74;
  wire       [2:0]    all_zeros_43;
  wire       [2:0]    all_left_zeros_43;
  wire       [2:0]    whole_bit_count_23;
  wire       [2:0]    left_bit_count_23;
  wire       [1:0]    _zz_75;
  wire       [1:0]    all_zeros_44;
  wire       [1:0]    all_left_zeros_44;
  wire       [1:0]    whole_bit_count_24;
  wire       [1:0]    left_bit_count_24;
  wire       [0:0]    _zz_76;
  wire       [0:0]    _zz_77;
  wire       [0:0]    all_zeros_45;
  wire       [0:0]    all_left_zeros_45;
  wire       [1:0]    left_all_zeros_count_20;
  wire       [0:0]    _zz_78;
  wire       [0:0]    _zz_79;
  wire       [0:0]    all_zeros_46;
  wire       [0:0]    all_left_zeros_46;
  wire       [1:0]    left_non_all_zeros_count_18;
  wire       [1:0]    non_zeros_lzc_18;
  wire       [2:0]    left_all_zeros_count_21;
  wire       [1:0]    _zz_80;
  wire       [1:0]    all_zeros_47;
  wire       [1:0]    all_left_zeros_47;
  wire       [1:0]    whole_bit_count_25;
  wire       [1:0]    left_bit_count_25;
  wire       [0:0]    _zz_81;
  wire       [0:0]    _zz_82;
  wire       [0:0]    all_zeros_48;
  wire       [0:0]    all_left_zeros_48;
  wire       [1:0]    left_all_zeros_count_22;
  wire       [0:0]    _zz_83;
  wire       [0:0]    _zz_84;
  wire       [0:0]    all_zeros_49;
  wire       [0:0]    all_left_zeros_49;
  wire       [1:0]    left_non_all_zeros_count_19;
  wire       [1:0]    non_zeros_lzc_19;
  wire       [2:0]    left_non_all_zeros_count_20;
  wire       [2:0]    non_zeros_lzc_20;
  wire       [3:0]    left_non_all_zeros_count_21;
  wire       [3:0]    non_zeros_lzc_21;
  wire       [4:0]    left_all_zeros_count_23;
  wire       [7:0]    _zz_85;
  wire       [3:0]    all_zeros_50;
  wire       [3:0]    all_left_zeros_50;
  wire       [3:0]    whole_bit_count_26;
  wire       [3:0]    left_bit_count_26;
  wire       [3:0]    _zz_86;
  wire       [2:0]    all_zeros_51;
  wire       [2:0]    all_left_zeros_51;
  wire       [2:0]    whole_bit_count_27;
  wire       [2:0]    left_bit_count_27;
  wire       [1:0]    _zz_87;
  wire       [1:0]    all_zeros_52;
  wire       [1:0]    all_left_zeros_52;
  wire       [1:0]    whole_bit_count_28;
  wire       [1:0]    left_bit_count_28;
  wire       [0:0]    _zz_88;
  wire       [0:0]    _zz_89;
  wire       [0:0]    all_zeros_53;
  wire       [0:0]    all_left_zeros_53;
  wire       [1:0]    left_all_zeros_count_24;
  wire       [0:0]    _zz_90;
  wire       [0:0]    _zz_91;
  wire       [0:0]    all_zeros_54;
  wire       [0:0]    all_left_zeros_54;
  wire       [1:0]    left_non_all_zeros_count_22;
  wire       [1:0]    non_zeros_lzc_22;
  wire       [2:0]    left_all_zeros_count_25;
  wire       [1:0]    _zz_92;
  wire       [1:0]    all_zeros_55;
  wire       [1:0]    all_left_zeros_55;
  wire       [1:0]    whole_bit_count_29;
  wire       [1:0]    left_bit_count_29;
  wire       [0:0]    _zz_93;
  wire       [0:0]    _zz_94;
  wire       [0:0]    all_zeros_56;
  wire       [0:0]    all_left_zeros_56;
  wire       [1:0]    left_all_zeros_count_26;
  wire       [0:0]    _zz_95;
  wire       [0:0]    _zz_96;
  wire       [0:0]    all_zeros_57;
  wire       [0:0]    all_left_zeros_57;
  wire       [1:0]    left_non_all_zeros_count_23;
  wire       [1:0]    non_zeros_lzc_23;
  wire       [2:0]    left_non_all_zeros_count_24;
  wire       [2:0]    non_zeros_lzc_24;
  wire       [3:0]    left_all_zeros_count_27;
  wire       [3:0]    _zz_97;
  wire       [2:0]    all_zeros_58;
  wire       [2:0]    all_left_zeros_58;
  wire       [2:0]    whole_bit_count_30;
  wire       [2:0]    left_bit_count_30;
  wire       [1:0]    _zz_98;
  wire       [1:0]    all_zeros_59;
  wire       [1:0]    all_left_zeros_59;
  wire       [1:0]    whole_bit_count_31;
  wire       [1:0]    left_bit_count_31;
  wire       [0:0]    _zz_99;
  wire       [0:0]    _zz_100;
  wire       [0:0]    all_zeros_60;
  wire       [0:0]    all_left_zeros_60;
  wire       [1:0]    left_all_zeros_count_28;
  wire       [0:0]    _zz_101;
  wire       [0:0]    _zz_102;
  wire       [0:0]    all_zeros_61;
  wire       [0:0]    all_left_zeros_61;
  wire       [1:0]    left_non_all_zeros_count_25;
  wire       [1:0]    non_zeros_lzc_25;
  wire       [2:0]    left_all_zeros_count_29;
  wire       [1:0]    _zz_103;
  wire       [1:0]    all_zeros_62;
  wire       [1:0]    all_left_zeros_62;
  wire       [1:0]    whole_bit_count_32;
  wire       [1:0]    left_bit_count_32;
  wire       [0:0]    _zz_104;
  wire       [0:0]    _zz_105;
  wire       [0:0]    all_zeros_63;
  wire       [0:0]    all_left_zeros_63;
  wire       [1:0]    left_all_zeros_count_30;
  wire       [0:0]    _zz_106;
  wire       [0:0]    _zz_107;
  wire       [0:0]    all_zeros_64;
  wire       [0:0]    all_left_zeros_64;
  wire       [1:0]    left_non_all_zeros_count_26;
  wire       [1:0]    non_zeros_lzc_26;
  wire       [2:0]    left_non_all_zeros_count_27;
  wire       [2:0]    non_zeros_lzc_27;
  wire       [3:0]    left_non_all_zeros_count_28;
  wire       [3:0]    non_zeros_lzc_28;
  wire       [4:0]    left_non_all_zeros_count_29;
  wire       [4:0]    non_zeros_lzc_29;
  wire       [5:0]    left_non_all_zeros_count_30;
  wire       [5:0]    non_zeros_lzc_30;
  wire       [6:0]    left_all_zeros_count_31;
  wire       [31:0]   _zz_108;
  wire       [5:0]    all_zeros_65;
  wire       [5:0]    all_left_zeros_65;
  wire       [5:0]    whole_bit_count_33;
  wire       [5:0]    left_bit_count_33;
  wire       [15:0]   _zz_109;
  wire       [4:0]    all_zeros_66;
  wire       [4:0]    all_left_zeros_66;
  wire       [4:0]    whole_bit_count_34;
  wire       [4:0]    left_bit_count_34;
  wire       [7:0]    _zz_110;
  wire       [3:0]    all_zeros_67;
  wire       [3:0]    all_left_zeros_67;
  wire       [3:0]    whole_bit_count_35;
  wire       [3:0]    left_bit_count_35;
  wire       [3:0]    _zz_111;
  wire       [2:0]    all_zeros_68;
  wire       [2:0]    all_left_zeros_68;
  wire       [2:0]    whole_bit_count_36;
  wire       [2:0]    left_bit_count_36;
  wire       [1:0]    _zz_112;
  wire       [1:0]    all_zeros_69;
  wire       [1:0]    all_left_zeros_69;
  wire       [1:0]    whole_bit_count_37;
  wire       [1:0]    left_bit_count_37;
  wire       [0:0]    _zz_113;
  wire       [0:0]    _zz_114;
  wire       [0:0]    all_zeros_70;
  wire       [0:0]    all_left_zeros_70;
  wire       [1:0]    left_all_zeros_count_32;
  wire       [0:0]    _zz_115;
  wire       [0:0]    _zz_116;
  wire       [0:0]    all_zeros_71;
  wire       [0:0]    all_left_zeros_71;
  wire       [1:0]    left_non_all_zeros_count_31;
  wire       [1:0]    non_zeros_lzc_31;
  wire       [2:0]    left_all_zeros_count_33;
  wire       [1:0]    _zz_117;
  wire       [1:0]    all_zeros_72;
  wire       [1:0]    all_left_zeros_72;
  wire       [1:0]    whole_bit_count_38;
  wire       [1:0]    left_bit_count_38;
  wire       [0:0]    _zz_118;
  wire       [0:0]    _zz_119;
  wire       [0:0]    all_zeros_73;
  wire       [0:0]    all_left_zeros_73;
  wire       [1:0]    left_all_zeros_count_34;
  wire       [0:0]    _zz_120;
  wire       [0:0]    _zz_121;
  wire       [0:0]    all_zeros_74;
  wire       [0:0]    all_left_zeros_74;
  wire       [1:0]    left_non_all_zeros_count_32;
  wire       [1:0]    non_zeros_lzc_32;
  wire       [2:0]    left_non_all_zeros_count_33;
  wire       [2:0]    non_zeros_lzc_33;
  wire       [3:0]    left_all_zeros_count_35;
  wire       [3:0]    _zz_122;
  wire       [2:0]    all_zeros_75;
  wire       [2:0]    all_left_zeros_75;
  wire       [2:0]    whole_bit_count_39;
  wire       [2:0]    left_bit_count_39;
  wire       [1:0]    _zz_123;
  wire       [1:0]    all_zeros_76;
  wire       [1:0]    all_left_zeros_76;
  wire       [1:0]    whole_bit_count_40;
  wire       [1:0]    left_bit_count_40;
  wire       [0:0]    _zz_124;
  wire       [0:0]    _zz_125;
  wire       [0:0]    all_zeros_77;
  wire       [0:0]    all_left_zeros_77;
  wire       [1:0]    left_all_zeros_count_36;
  wire       [0:0]    _zz_126;
  wire       [0:0]    _zz_127;
  wire       [0:0]    all_zeros_78;
  wire       [0:0]    all_left_zeros_78;
  wire       [1:0]    left_non_all_zeros_count_34;
  wire       [1:0]    non_zeros_lzc_34;
  wire       [2:0]    left_all_zeros_count_37;
  wire       [1:0]    _zz_128;
  wire       [1:0]    all_zeros_79;
  wire       [1:0]    all_left_zeros_79;
  wire       [1:0]    whole_bit_count_41;
  wire       [1:0]    left_bit_count_41;
  wire       [0:0]    _zz_129;
  wire       [0:0]    _zz_130;
  wire       [0:0]    all_zeros_80;
  wire       [0:0]    all_left_zeros_80;
  wire       [1:0]    left_all_zeros_count_38;
  wire       [0:0]    _zz_131;
  wire       [0:0]    _zz_132;
  wire       [0:0]    all_zeros_81;
  wire       [0:0]    all_left_zeros_81;
  wire       [1:0]    left_non_all_zeros_count_35;
  wire       [1:0]    non_zeros_lzc_35;
  wire       [2:0]    left_non_all_zeros_count_36;
  wire       [2:0]    non_zeros_lzc_36;
  wire       [3:0]    left_non_all_zeros_count_37;
  wire       [3:0]    non_zeros_lzc_37;
  wire       [4:0]    left_all_zeros_count_39;
  wire       [7:0]    _zz_133;
  wire       [3:0]    all_zeros_82;
  wire       [3:0]    all_left_zeros_82;
  wire       [3:0]    whole_bit_count_42;
  wire       [3:0]    left_bit_count_42;
  wire       [3:0]    _zz_134;
  wire       [2:0]    all_zeros_83;
  wire       [2:0]    all_left_zeros_83;
  wire       [2:0]    whole_bit_count_43;
  wire       [2:0]    left_bit_count_43;
  wire       [1:0]    _zz_135;
  wire       [1:0]    all_zeros_84;
  wire       [1:0]    all_left_zeros_84;
  wire       [1:0]    whole_bit_count_44;
  wire       [1:0]    left_bit_count_44;
  wire       [0:0]    _zz_136;
  wire       [0:0]    _zz_137;
  wire       [0:0]    all_zeros_85;
  wire       [0:0]    all_left_zeros_85;
  wire       [1:0]    left_all_zeros_count_40;
  wire       [0:0]    _zz_138;
  wire       [0:0]    _zz_139;
  wire       [0:0]    all_zeros_86;
  wire       [0:0]    all_left_zeros_86;
  wire       [1:0]    left_non_all_zeros_count_38;
  wire       [1:0]    non_zeros_lzc_38;
  wire       [2:0]    left_all_zeros_count_41;
  wire       [1:0]    _zz_140;
  wire       [1:0]    all_zeros_87;
  wire       [1:0]    all_left_zeros_87;
  wire       [1:0]    whole_bit_count_45;
  wire       [1:0]    left_bit_count_45;
  wire       [0:0]    _zz_141;
  wire       [0:0]    _zz_142;
  wire       [0:0]    all_zeros_88;
  wire       [0:0]    all_left_zeros_88;
  wire       [1:0]    left_all_zeros_count_42;
  wire       [0:0]    _zz_143;
  wire       [0:0]    _zz_144;
  wire       [0:0]    all_zeros_89;
  wire       [0:0]    all_left_zeros_89;
  wire       [1:0]    left_non_all_zeros_count_39;
  wire       [1:0]    non_zeros_lzc_39;
  wire       [2:0]    left_non_all_zeros_count_40;
  wire       [2:0]    non_zeros_lzc_40;
  wire       [3:0]    left_all_zeros_count_43;
  wire       [3:0]    _zz_145;
  wire       [2:0]    all_zeros_90;
  wire       [2:0]    all_left_zeros_90;
  wire       [2:0]    whole_bit_count_46;
  wire       [2:0]    left_bit_count_46;
  wire       [1:0]    _zz_146;
  wire       [1:0]    all_zeros_91;
  wire       [1:0]    all_left_zeros_91;
  wire       [1:0]    whole_bit_count_47;
  wire       [1:0]    left_bit_count_47;
  wire       [0:0]    _zz_147;
  wire       [0:0]    _zz_148;
  wire       [0:0]    all_zeros_92;
  wire       [0:0]    all_left_zeros_92;
  wire       [1:0]    left_all_zeros_count_44;
  wire       [0:0]    _zz_149;
  wire       [0:0]    _zz_150;
  wire       [0:0]    all_zeros_93;
  wire       [0:0]    all_left_zeros_93;
  wire       [1:0]    left_non_all_zeros_count_41;
  wire       [1:0]    non_zeros_lzc_41;
  wire       [2:0]    left_all_zeros_count_45;
  wire       [1:0]    _zz_151;
  wire       [1:0]    all_zeros_94;
  wire       [1:0]    all_left_zeros_94;
  wire       [1:0]    whole_bit_count_48;
  wire       [1:0]    left_bit_count_48;
  wire       [0:0]    _zz_152;
  wire       [0:0]    _zz_153;
  wire       [0:0]    all_zeros_95;
  wire       [0:0]    all_left_zeros_95;
  wire       [1:0]    left_all_zeros_count_46;
  wire       [0:0]    _zz_154;
  wire       [0:0]    _zz_155;
  wire       [0:0]    all_zeros_96;
  wire       [0:0]    all_left_zeros_96;
  wire       [1:0]    left_non_all_zeros_count_42;
  wire       [1:0]    non_zeros_lzc_42;
  wire       [2:0]    left_non_all_zeros_count_43;
  wire       [2:0]    non_zeros_lzc_43;
  wire       [3:0]    left_non_all_zeros_count_44;
  wire       [3:0]    non_zeros_lzc_44;
  wire       [4:0]    left_non_all_zeros_count_45;
  wire       [4:0]    non_zeros_lzc_45;
  wire       [5:0]    left_all_zeros_count_47;
  wire       [15:0]   _zz_156;
  wire       [4:0]    all_zeros_97;
  wire       [4:0]    all_left_zeros_97;
  wire       [4:0]    whole_bit_count_49;
  wire       [4:0]    left_bit_count_49;
  wire       [7:0]    _zz_157;
  wire       [3:0]    all_zeros_98;
  wire       [3:0]    all_left_zeros_98;
  wire       [3:0]    whole_bit_count_50;
  wire       [3:0]    left_bit_count_50;
  wire       [3:0]    _zz_158;
  wire       [2:0]    all_zeros_99;
  wire       [2:0]    all_left_zeros_99;
  wire       [2:0]    whole_bit_count_51;
  wire       [2:0]    left_bit_count_51;
  wire       [1:0]    _zz_159;
  wire       [1:0]    all_zeros_100;
  wire       [1:0]    all_left_zeros_100;
  wire       [1:0]    whole_bit_count_52;
  wire       [1:0]    left_bit_count_52;
  wire       [0:0]    _zz_160;
  wire       [0:0]    _zz_161;
  wire       [0:0]    all_zeros_101;
  wire       [0:0]    all_left_zeros_101;
  wire       [1:0]    left_all_zeros_count_48;
  wire       [0:0]    _zz_162;
  wire       [0:0]    _zz_163;
  wire       [0:0]    all_zeros_102;
  wire       [0:0]    all_left_zeros_102;
  wire       [1:0]    left_non_all_zeros_count_46;
  wire       [1:0]    non_zeros_lzc_46;
  wire       [2:0]    left_all_zeros_count_49;
  wire       [1:0]    _zz_164;
  wire       [1:0]    all_zeros_103;
  wire       [1:0]    all_left_zeros_103;
  wire       [1:0]    whole_bit_count_53;
  wire       [1:0]    left_bit_count_53;
  wire       [0:0]    _zz_165;
  wire       [0:0]    _zz_166;
  wire       [0:0]    all_zeros_104;
  wire       [0:0]    all_left_zeros_104;
  wire       [1:0]    left_all_zeros_count_50;
  wire       [0:0]    _zz_167;
  wire       [0:0]    _zz_168;
  wire       [0:0]    all_zeros_105;
  wire       [0:0]    all_left_zeros_105;
  wire       [1:0]    left_non_all_zeros_count_47;
  wire       [1:0]    non_zeros_lzc_47;
  wire       [2:0]    left_non_all_zeros_count_48;
  wire       [2:0]    non_zeros_lzc_48;
  wire       [3:0]    left_all_zeros_count_51;
  wire       [3:0]    _zz_169;
  wire       [2:0]    all_zeros_106;
  wire       [2:0]    all_left_zeros_106;
  wire       [2:0]    whole_bit_count_54;
  wire       [2:0]    left_bit_count_54;
  wire       [1:0]    _zz_170;
  wire       [1:0]    all_zeros_107;
  wire       [1:0]    all_left_zeros_107;
  wire       [1:0]    whole_bit_count_55;
  wire       [1:0]    left_bit_count_55;
  wire       [0:0]    _zz_171;
  wire       [0:0]    _zz_172;
  wire       [0:0]    all_zeros_108;
  wire       [0:0]    all_left_zeros_108;
  wire       [1:0]    left_all_zeros_count_52;
  wire       [0:0]    _zz_173;
  wire       [0:0]    _zz_174;
  wire       [0:0]    all_zeros_109;
  wire       [0:0]    all_left_zeros_109;
  wire       [1:0]    left_non_all_zeros_count_49;
  wire       [1:0]    non_zeros_lzc_49;
  wire       [2:0]    left_all_zeros_count_53;
  wire       [1:0]    _zz_175;
  wire       [1:0]    all_zeros_110;
  wire       [1:0]    all_left_zeros_110;
  wire       [1:0]    whole_bit_count_56;
  wire       [1:0]    left_bit_count_56;
  wire       [0:0]    _zz_176;
  wire       [0:0]    _zz_177;
  wire       [0:0]    all_zeros_111;
  wire       [0:0]    all_left_zeros_111;
  wire       [1:0]    left_all_zeros_count_54;
  wire       [0:0]    _zz_178;
  wire       [0:0]    _zz_179;
  wire       [0:0]    all_zeros_112;
  wire       [0:0]    all_left_zeros_112;
  wire       [1:0]    left_non_all_zeros_count_50;
  wire       [1:0]    non_zeros_lzc_50;
  wire       [2:0]    left_non_all_zeros_count_51;
  wire       [2:0]    non_zeros_lzc_51;
  wire       [3:0]    left_non_all_zeros_count_52;
  wire       [3:0]    non_zeros_lzc_52;
  wire       [4:0]    left_all_zeros_count_55;
  wire       [7:0]    _zz_180;
  wire       [3:0]    all_zeros_113;
  wire       [3:0]    all_left_zeros_113;
  wire       [3:0]    whole_bit_count_57;
  wire       [3:0]    left_bit_count_57;
  wire       [3:0]    _zz_181;
  wire       [2:0]    all_zeros_114;
  wire       [2:0]    all_left_zeros_114;
  wire       [2:0]    whole_bit_count_58;
  wire       [2:0]    left_bit_count_58;
  wire       [1:0]    _zz_182;
  wire       [1:0]    all_zeros_115;
  wire       [1:0]    all_left_zeros_115;
  wire       [1:0]    whole_bit_count_59;
  wire       [1:0]    left_bit_count_59;
  wire       [0:0]    _zz_183;
  wire       [0:0]    _zz_184;
  wire       [0:0]    all_zeros_116;
  wire       [0:0]    all_left_zeros_116;
  wire       [1:0]    left_all_zeros_count_56;
  wire       [0:0]    _zz_185;
  wire       [0:0]    _zz_186;
  wire       [0:0]    all_zeros_117;
  wire       [0:0]    all_left_zeros_117;
  wire       [1:0]    left_non_all_zeros_count_53;
  wire       [1:0]    non_zeros_lzc_53;
  wire       [2:0]    left_all_zeros_count_57;
  wire       [1:0]    _zz_187;
  wire       [1:0]    all_zeros_118;
  wire       [1:0]    all_left_zeros_118;
  wire       [1:0]    whole_bit_count_60;
  wire       [1:0]    left_bit_count_60;
  wire       [0:0]    _zz_188;
  wire       [0:0]    _zz_189;
  wire       [0:0]    all_zeros_119;
  wire       [0:0]    all_left_zeros_119;
  wire       [1:0]    left_all_zeros_count_58;
  wire       [0:0]    _zz_190;
  wire       [0:0]    _zz_191;
  wire       [0:0]    all_zeros_120;
  wire       [0:0]    all_left_zeros_120;
  wire       [1:0]    left_non_all_zeros_count_54;
  wire       [1:0]    non_zeros_lzc_54;
  wire       [2:0]    left_non_all_zeros_count_55;
  wire       [2:0]    non_zeros_lzc_55;
  wire       [3:0]    left_all_zeros_count_59;
  wire       [3:0]    _zz_192;
  wire       [2:0]    all_zeros_121;
  wire       [2:0]    all_left_zeros_121;
  wire       [2:0]    whole_bit_count_61;
  wire       [2:0]    left_bit_count_61;
  wire       [1:0]    _zz_193;
  wire       [1:0]    all_zeros_122;
  wire       [1:0]    all_left_zeros_122;
  wire       [1:0]    whole_bit_count_62;
  wire       [1:0]    left_bit_count_62;
  wire       [0:0]    _zz_194;
  wire       [0:0]    _zz_195;
  wire       [0:0]    all_zeros_123;
  wire       [0:0]    all_left_zeros_123;
  wire       [1:0]    left_all_zeros_count_60;
  wire       [0:0]    _zz_196;
  wire       [0:0]    _zz_197;
  wire       [0:0]    all_zeros_124;
  wire       [0:0]    all_left_zeros_124;
  wire       [1:0]    left_non_all_zeros_count_56;
  wire       [1:0]    non_zeros_lzc_56;
  wire       [2:0]    left_all_zeros_count_61;
  wire       [1:0]    _zz_198;
  wire       [1:0]    all_zeros_125;
  wire       [1:0]    all_left_zeros_125;
  wire       [1:0]    whole_bit_count_63;
  wire       [1:0]    left_bit_count_63;
  wire       [0:0]    _zz_199;
  wire       [0:0]    _zz_200;
  wire       [0:0]    all_zeros_126;
  wire       [0:0]    all_left_zeros_126;
  wire       [1:0]    left_all_zeros_count_62;
  wire       [0:0]    _zz_201;
  wire       [0:0]    _zz_202;
  wire       [0:0]    all_zeros_127;
  wire       [0:0]    all_left_zeros_127;
  wire       [1:0]    left_non_all_zeros_count_57;
  wire       [1:0]    non_zeros_lzc_57;
  wire       [2:0]    left_non_all_zeros_count_58;
  wire       [2:0]    non_zeros_lzc_58;
  wire       [3:0]    left_non_all_zeros_count_59;
  wire       [3:0]    non_zeros_lzc_59;
  wire       [4:0]    left_non_all_zeros_count_60;
  wire       [4:0]    non_zeros_lzc_60;
  wire       [5:0]    left_non_all_zeros_count_61;
  wire       [5:0]    non_zeros_lzc_61;
  wire       [6:0]    left_non_all_zeros_count_62;
  wire       [6:0]    non_zeros_lzc_62;
  wire       [7:0]    left_all_zeros_count_63;
  wire       [63:0]   _zz_203;
  wire       [6:0]    all_zeros_128;
  wire       [6:0]    all_left_zeros_128;
  wire       [6:0]    whole_bit_count_64;
  wire       [6:0]    left_bit_count_64;
  wire       [31:0]   _zz_204;
  wire       [5:0]    all_zeros_129;
  wire       [5:0]    all_left_zeros_129;
  wire       [5:0]    whole_bit_count_65;
  wire       [5:0]    left_bit_count_65;
  wire       [15:0]   _zz_205;
  wire       [4:0]    all_zeros_130;
  wire       [4:0]    all_left_zeros_130;
  wire       [4:0]    whole_bit_count_66;
  wire       [4:0]    left_bit_count_66;
  wire       [7:0]    _zz_206;
  wire       [3:0]    all_zeros_131;
  wire       [3:0]    all_left_zeros_131;
  wire       [3:0]    whole_bit_count_67;
  wire       [3:0]    left_bit_count_67;
  wire       [3:0]    _zz_207;
  wire       [2:0]    all_zeros_132;
  wire       [2:0]    all_left_zeros_132;
  wire       [2:0]    whole_bit_count_68;
  wire       [2:0]    left_bit_count_68;
  wire       [1:0]    _zz_208;
  wire       [1:0]    all_zeros_133;
  wire       [1:0]    all_left_zeros_133;
  wire       [1:0]    whole_bit_count_69;
  wire       [1:0]    left_bit_count_69;
  wire       [0:0]    _zz_209;
  wire       [0:0]    _zz_210;
  wire       [0:0]    all_zeros_134;
  wire       [0:0]    all_left_zeros_134;
  wire       [1:0]    left_all_zeros_count_64;
  wire       [0:0]    _zz_211;
  wire       [0:0]    _zz_212;
  wire       [0:0]    all_zeros_135;
  wire       [0:0]    all_left_zeros_135;
  wire       [1:0]    left_non_all_zeros_count_63;
  wire       [1:0]    non_zeros_lzc_63;
  wire       [2:0]    left_all_zeros_count_65;
  wire       [1:0]    _zz_213;
  wire       [1:0]    all_zeros_136;
  wire       [1:0]    all_left_zeros_136;
  wire       [1:0]    whole_bit_count_70;
  wire       [1:0]    left_bit_count_70;
  wire       [0:0]    _zz_214;
  wire       [0:0]    _zz_215;
  wire       [0:0]    all_zeros_137;
  wire       [0:0]    all_left_zeros_137;
  wire       [1:0]    left_all_zeros_count_66;
  wire       [0:0]    _zz_216;
  wire       [0:0]    _zz_217;
  wire       [0:0]    all_zeros_138;
  wire       [0:0]    all_left_zeros_138;
  wire       [1:0]    left_non_all_zeros_count_64;
  wire       [1:0]    non_zeros_lzc_64;
  wire       [2:0]    left_non_all_zeros_count_65;
  wire       [2:0]    non_zeros_lzc_65;
  wire       [3:0]    left_all_zeros_count_67;
  wire       [3:0]    _zz_218;
  wire       [2:0]    all_zeros_139;
  wire       [2:0]    all_left_zeros_139;
  wire       [2:0]    whole_bit_count_71;
  wire       [2:0]    left_bit_count_71;
  wire       [1:0]    _zz_219;
  wire       [1:0]    all_zeros_140;
  wire       [1:0]    all_left_zeros_140;
  wire       [1:0]    whole_bit_count_72;
  wire       [1:0]    left_bit_count_72;
  wire       [0:0]    _zz_220;
  wire       [0:0]    _zz_221;
  wire       [0:0]    all_zeros_141;
  wire       [0:0]    all_left_zeros_141;
  wire       [1:0]    left_all_zeros_count_68;
  wire       [0:0]    _zz_222;
  wire       [0:0]    _zz_223;
  wire       [0:0]    all_zeros_142;
  wire       [0:0]    all_left_zeros_142;
  wire       [1:0]    left_non_all_zeros_count_66;
  wire       [1:0]    non_zeros_lzc_66;
  wire       [2:0]    left_all_zeros_count_69;
  wire       [1:0]    _zz_224;
  wire       [1:0]    all_zeros_143;
  wire       [1:0]    all_left_zeros_143;
  wire       [1:0]    whole_bit_count_73;
  wire       [1:0]    left_bit_count_73;
  wire       [0:0]    _zz_225;
  wire       [0:0]    _zz_226;
  wire       [0:0]    all_zeros_144;
  wire       [0:0]    all_left_zeros_144;
  wire       [1:0]    left_all_zeros_count_70;
  wire       [0:0]    _zz_227;
  wire       [0:0]    _zz_228;
  wire       [0:0]    all_zeros_145;
  wire       [0:0]    all_left_zeros_145;
  wire       [1:0]    left_non_all_zeros_count_67;
  wire       [1:0]    non_zeros_lzc_67;
  wire       [2:0]    left_non_all_zeros_count_68;
  wire       [2:0]    non_zeros_lzc_68;
  wire       [3:0]    left_non_all_zeros_count_69;
  wire       [3:0]    non_zeros_lzc_69;
  wire       [4:0]    left_all_zeros_count_71;
  wire       [7:0]    _zz_229;
  wire       [3:0]    all_zeros_146;
  wire       [3:0]    all_left_zeros_146;
  wire       [3:0]    whole_bit_count_74;
  wire       [3:0]    left_bit_count_74;
  wire       [3:0]    _zz_230;
  wire       [2:0]    all_zeros_147;
  wire       [2:0]    all_left_zeros_147;
  wire       [2:0]    whole_bit_count_75;
  wire       [2:0]    left_bit_count_75;
  wire       [1:0]    _zz_231;
  wire       [1:0]    all_zeros_148;
  wire       [1:0]    all_left_zeros_148;
  wire       [1:0]    whole_bit_count_76;
  wire       [1:0]    left_bit_count_76;
  wire       [0:0]    _zz_232;
  wire       [0:0]    _zz_233;
  wire       [0:0]    all_zeros_149;
  wire       [0:0]    all_left_zeros_149;
  wire       [1:0]    left_all_zeros_count_72;
  wire       [0:0]    _zz_234;
  wire       [0:0]    _zz_235;
  wire       [0:0]    all_zeros_150;
  wire       [0:0]    all_left_zeros_150;
  wire       [1:0]    left_non_all_zeros_count_70;
  wire       [1:0]    non_zeros_lzc_70;
  wire       [2:0]    left_all_zeros_count_73;
  wire       [1:0]    _zz_236;
  wire       [1:0]    all_zeros_151;
  wire       [1:0]    all_left_zeros_151;
  wire       [1:0]    whole_bit_count_77;
  wire       [1:0]    left_bit_count_77;
  wire       [0:0]    _zz_237;
  wire       [0:0]    _zz_238;
  wire       [0:0]    all_zeros_152;
  wire       [0:0]    all_left_zeros_152;
  wire       [1:0]    left_all_zeros_count_74;
  wire       [0:0]    _zz_239;
  wire       [0:0]    _zz_240;
  wire       [0:0]    all_zeros_153;
  wire       [0:0]    all_left_zeros_153;
  wire       [1:0]    left_non_all_zeros_count_71;
  wire       [1:0]    non_zeros_lzc_71;
  wire       [2:0]    left_non_all_zeros_count_72;
  wire       [2:0]    non_zeros_lzc_72;
  wire       [3:0]    left_all_zeros_count_75;
  wire       [3:0]    _zz_241;
  wire       [2:0]    all_zeros_154;
  wire       [2:0]    all_left_zeros_154;
  wire       [2:0]    whole_bit_count_78;
  wire       [2:0]    left_bit_count_78;
  wire       [1:0]    _zz_242;
  wire       [1:0]    all_zeros_155;
  wire       [1:0]    all_left_zeros_155;
  wire       [1:0]    whole_bit_count_79;
  wire       [1:0]    left_bit_count_79;
  wire       [0:0]    _zz_243;
  wire       [0:0]    _zz_244;
  wire       [0:0]    all_zeros_156;
  wire       [0:0]    all_left_zeros_156;
  wire       [1:0]    left_all_zeros_count_76;
  wire       [0:0]    _zz_245;
  wire       [0:0]    _zz_246;
  wire       [0:0]    all_zeros_157;
  wire       [0:0]    all_left_zeros_157;
  wire       [1:0]    left_non_all_zeros_count_73;
  wire       [1:0]    non_zeros_lzc_73;
  wire       [2:0]    left_all_zeros_count_77;
  wire       [1:0]    _zz_247;
  wire       [1:0]    all_zeros_158;
  wire       [1:0]    all_left_zeros_158;
  wire       [1:0]    whole_bit_count_80;
  wire       [1:0]    left_bit_count_80;
  wire       [0:0]    _zz_248;
  wire       [0:0]    _zz_249;
  wire       [0:0]    all_zeros_159;
  wire       [0:0]    all_left_zeros_159;
  wire       [1:0]    left_all_zeros_count_78;
  wire       [0:0]    _zz_250;
  wire       [0:0]    _zz_251;
  wire       [0:0]    all_zeros_160;
  wire       [0:0]    all_left_zeros_160;
  wire       [1:0]    left_non_all_zeros_count_74;
  wire       [1:0]    non_zeros_lzc_74;
  wire       [2:0]    left_non_all_zeros_count_75;
  wire       [2:0]    non_zeros_lzc_75;
  wire       [3:0]    left_non_all_zeros_count_76;
  wire       [3:0]    non_zeros_lzc_76;
  wire       [4:0]    left_non_all_zeros_count_77;
  wire       [4:0]    non_zeros_lzc_77;
  wire       [5:0]    left_all_zeros_count_79;
  wire       [15:0]   _zz_252;
  wire       [4:0]    all_zeros_161;
  wire       [4:0]    all_left_zeros_161;
  wire       [4:0]    whole_bit_count_81;
  wire       [4:0]    left_bit_count_81;
  wire       [7:0]    _zz_253;
  wire       [3:0]    all_zeros_162;
  wire       [3:0]    all_left_zeros_162;
  wire       [3:0]    whole_bit_count_82;
  wire       [3:0]    left_bit_count_82;
  wire       [3:0]    _zz_254;
  wire       [2:0]    all_zeros_163;
  wire       [2:0]    all_left_zeros_163;
  wire       [2:0]    whole_bit_count_83;
  wire       [2:0]    left_bit_count_83;
  wire       [1:0]    _zz_255;
  wire       [1:0]    all_zeros_164;
  wire       [1:0]    all_left_zeros_164;
  wire       [1:0]    whole_bit_count_84;
  wire       [1:0]    left_bit_count_84;
  wire       [0:0]    _zz_256;
  wire       [0:0]    _zz_257;
  wire       [0:0]    all_zeros_165;
  wire       [0:0]    all_left_zeros_165;
  wire       [1:0]    left_all_zeros_count_80;
  wire       [0:0]    _zz_258;
  wire       [0:0]    _zz_259;
  wire       [0:0]    all_zeros_166;
  wire       [0:0]    all_left_zeros_166;
  wire       [1:0]    left_non_all_zeros_count_78;
  wire       [1:0]    non_zeros_lzc_78;
  wire       [2:0]    left_all_zeros_count_81;
  wire       [1:0]    _zz_260;
  wire       [1:0]    all_zeros_167;
  wire       [1:0]    all_left_zeros_167;
  wire       [1:0]    whole_bit_count_85;
  wire       [1:0]    left_bit_count_85;
  wire       [0:0]    _zz_261;
  wire       [0:0]    _zz_262;
  wire       [0:0]    all_zeros_168;
  wire       [0:0]    all_left_zeros_168;
  wire       [1:0]    left_all_zeros_count_82;
  wire       [0:0]    _zz_263;
  wire       [0:0]    _zz_264;
  wire       [0:0]    all_zeros_169;
  wire       [0:0]    all_left_zeros_169;
  wire       [1:0]    left_non_all_zeros_count_79;
  wire       [1:0]    non_zeros_lzc_79;
  wire       [2:0]    left_non_all_zeros_count_80;
  wire       [2:0]    non_zeros_lzc_80;
  wire       [3:0]    left_all_zeros_count_83;
  wire       [3:0]    _zz_265;
  wire       [2:0]    all_zeros_170;
  wire       [2:0]    all_left_zeros_170;
  wire       [2:0]    whole_bit_count_86;
  wire       [2:0]    left_bit_count_86;
  wire       [1:0]    _zz_266;
  wire       [1:0]    all_zeros_171;
  wire       [1:0]    all_left_zeros_171;
  wire       [1:0]    whole_bit_count_87;
  wire       [1:0]    left_bit_count_87;
  wire       [0:0]    _zz_267;
  wire       [0:0]    _zz_268;
  wire       [0:0]    all_zeros_172;
  wire       [0:0]    all_left_zeros_172;
  wire       [1:0]    left_all_zeros_count_84;
  wire       [0:0]    _zz_269;
  wire       [0:0]    _zz_270;
  wire       [0:0]    all_zeros_173;
  wire       [0:0]    all_left_zeros_173;
  wire       [1:0]    left_non_all_zeros_count_81;
  wire       [1:0]    non_zeros_lzc_81;
  wire       [2:0]    left_all_zeros_count_85;
  wire       [1:0]    _zz_271;
  wire       [1:0]    all_zeros_174;
  wire       [1:0]    all_left_zeros_174;
  wire       [1:0]    whole_bit_count_88;
  wire       [1:0]    left_bit_count_88;
  wire       [0:0]    _zz_272;
  wire       [0:0]    _zz_273;
  wire       [0:0]    all_zeros_175;
  wire       [0:0]    all_left_zeros_175;
  wire       [1:0]    left_all_zeros_count_86;
  wire       [0:0]    _zz_274;
  wire       [0:0]    _zz_275;
  wire       [0:0]    all_zeros_176;
  wire       [0:0]    all_left_zeros_176;
  wire       [1:0]    left_non_all_zeros_count_82;
  wire       [1:0]    non_zeros_lzc_82;
  wire       [2:0]    left_non_all_zeros_count_83;
  wire       [2:0]    non_zeros_lzc_83;
  wire       [3:0]    left_non_all_zeros_count_84;
  wire       [3:0]    non_zeros_lzc_84;
  wire       [4:0]    left_all_zeros_count_87;
  wire       [7:0]    _zz_276;
  wire       [3:0]    all_zeros_177;
  wire       [3:0]    all_left_zeros_177;
  wire       [3:0]    whole_bit_count_89;
  wire       [3:0]    left_bit_count_89;
  wire       [3:0]    _zz_277;
  wire       [2:0]    all_zeros_178;
  wire       [2:0]    all_left_zeros_178;
  wire       [2:0]    whole_bit_count_90;
  wire       [2:0]    left_bit_count_90;
  wire       [1:0]    _zz_278;
  wire       [1:0]    all_zeros_179;
  wire       [1:0]    all_left_zeros_179;
  wire       [1:0]    whole_bit_count_91;
  wire       [1:0]    left_bit_count_91;
  wire       [0:0]    _zz_279;
  wire       [0:0]    _zz_280;
  wire       [0:0]    all_zeros_180;
  wire       [0:0]    all_left_zeros_180;
  wire       [1:0]    left_all_zeros_count_88;
  wire       [0:0]    _zz_281;
  wire       [0:0]    _zz_282;
  wire       [0:0]    all_zeros_181;
  wire       [0:0]    all_left_zeros_181;
  wire       [1:0]    left_non_all_zeros_count_85;
  wire       [1:0]    non_zeros_lzc_85;
  wire       [2:0]    left_all_zeros_count_89;
  wire       [1:0]    _zz_283;
  wire       [1:0]    all_zeros_182;
  wire       [1:0]    all_left_zeros_182;
  wire       [1:0]    whole_bit_count_92;
  wire       [1:0]    left_bit_count_92;
  wire       [0:0]    _zz_284;
  wire       [0:0]    _zz_285;
  wire       [0:0]    all_zeros_183;
  wire       [0:0]    all_left_zeros_183;
  wire       [1:0]    left_all_zeros_count_90;
  wire       [0:0]    _zz_286;
  wire       [0:0]    _zz_287;
  wire       [0:0]    all_zeros_184;
  wire       [0:0]    all_left_zeros_184;
  wire       [1:0]    left_non_all_zeros_count_86;
  wire       [1:0]    non_zeros_lzc_86;
  wire       [2:0]    left_non_all_zeros_count_87;
  wire       [2:0]    non_zeros_lzc_87;
  wire       [3:0]    left_all_zeros_count_91;
  wire       [3:0]    _zz_288;
  wire       [2:0]    all_zeros_185;
  wire       [2:0]    all_left_zeros_185;
  wire       [2:0]    whole_bit_count_93;
  wire       [2:0]    left_bit_count_93;
  wire       [1:0]    _zz_289;
  wire       [1:0]    all_zeros_186;
  wire       [1:0]    all_left_zeros_186;
  wire       [1:0]    whole_bit_count_94;
  wire       [1:0]    left_bit_count_94;
  wire       [0:0]    _zz_290;
  wire       [0:0]    _zz_291;
  wire       [0:0]    all_zeros_187;
  wire       [0:0]    all_left_zeros_187;
  wire       [1:0]    left_all_zeros_count_92;
  wire       [0:0]    _zz_292;
  wire       [0:0]    _zz_293;
  wire       [0:0]    all_zeros_188;
  wire       [0:0]    all_left_zeros_188;
  wire       [1:0]    left_non_all_zeros_count_88;
  wire       [1:0]    non_zeros_lzc_88;
  wire       [2:0]    left_all_zeros_count_93;
  wire       [1:0]    _zz_294;
  wire       [1:0]    all_zeros_189;
  wire       [1:0]    all_left_zeros_189;
  wire       [1:0]    whole_bit_count_95;
  wire       [1:0]    left_bit_count_95;
  wire       [0:0]    _zz_295;
  wire       [0:0]    _zz_296;
  wire       [0:0]    all_zeros_190;
  wire       [0:0]    all_left_zeros_190;
  wire       [1:0]    left_all_zeros_count_94;
  wire       [0:0]    _zz_297;
  wire       [0:0]    _zz_298;
  wire       [0:0]    all_zeros_191;
  wire       [0:0]    all_left_zeros_191;
  wire       [1:0]    left_non_all_zeros_count_89;
  wire       [1:0]    non_zeros_lzc_89;
  wire       [2:0]    left_non_all_zeros_count_90;
  wire       [2:0]    non_zeros_lzc_90;
  wire       [3:0]    left_non_all_zeros_count_91;
  wire       [3:0]    non_zeros_lzc_91;
  wire       [4:0]    left_non_all_zeros_count_92;
  wire       [4:0]    non_zeros_lzc_92;
  wire       [5:0]    left_non_all_zeros_count_93;
  wire       [5:0]    non_zeros_lzc_93;
  wire       [6:0]    left_all_zeros_count_95;
  wire       [31:0]   _zz_299;
  wire       [5:0]    all_zeros_192;
  wire       [5:0]    all_left_zeros_192;
  wire       [5:0]    whole_bit_count_96;
  wire       [5:0]    left_bit_count_96;
  wire       [15:0]   _zz_300;
  wire       [4:0]    all_zeros_193;
  wire       [4:0]    all_left_zeros_193;
  wire       [4:0]    whole_bit_count_97;
  wire       [4:0]    left_bit_count_97;
  wire       [7:0]    _zz_301;
  wire       [3:0]    all_zeros_194;
  wire       [3:0]    all_left_zeros_194;
  wire       [3:0]    whole_bit_count_98;
  wire       [3:0]    left_bit_count_98;
  wire       [3:0]    _zz_302;
  wire       [2:0]    all_zeros_195;
  wire       [2:0]    all_left_zeros_195;
  wire       [2:0]    whole_bit_count_99;
  wire       [2:0]    left_bit_count_99;
  wire       [1:0]    _zz_303;
  wire       [1:0]    all_zeros_196;
  wire       [1:0]    all_left_zeros_196;
  wire       [1:0]    whole_bit_count_100;
  wire       [1:0]    left_bit_count_100;
  wire       [0:0]    _zz_304;
  wire       [0:0]    _zz_305;
  wire       [0:0]    all_zeros_197;
  wire       [0:0]    all_left_zeros_197;
  wire       [1:0]    left_all_zeros_count_96;
  wire       [0:0]    _zz_306;
  wire       [0:0]    _zz_307;
  wire       [0:0]    all_zeros_198;
  wire       [0:0]    all_left_zeros_198;
  wire       [1:0]    left_non_all_zeros_count_94;
  wire       [1:0]    non_zeros_lzc_94;
  wire       [2:0]    left_all_zeros_count_97;
  wire       [1:0]    _zz_308;
  wire       [1:0]    all_zeros_199;
  wire       [1:0]    all_left_zeros_199;
  wire       [1:0]    whole_bit_count_101;
  wire       [1:0]    left_bit_count_101;
  wire       [0:0]    _zz_309;
  wire       [0:0]    _zz_310;
  wire       [0:0]    all_zeros_200;
  wire       [0:0]    all_left_zeros_200;
  wire       [1:0]    left_all_zeros_count_98;
  wire       [0:0]    _zz_311;
  wire       [0:0]    _zz_312;
  wire       [0:0]    all_zeros_201;
  wire       [0:0]    all_left_zeros_201;
  wire       [1:0]    left_non_all_zeros_count_95;
  wire       [1:0]    non_zeros_lzc_95;
  wire       [2:0]    left_non_all_zeros_count_96;
  wire       [2:0]    non_zeros_lzc_96;
  wire       [3:0]    left_all_zeros_count_99;
  wire       [3:0]    _zz_313;
  wire       [2:0]    all_zeros_202;
  wire       [2:0]    all_left_zeros_202;
  wire       [2:0]    whole_bit_count_102;
  wire       [2:0]    left_bit_count_102;
  wire       [1:0]    _zz_314;
  wire       [1:0]    all_zeros_203;
  wire       [1:0]    all_left_zeros_203;
  wire       [1:0]    whole_bit_count_103;
  wire       [1:0]    left_bit_count_103;
  wire       [0:0]    _zz_315;
  wire       [0:0]    _zz_316;
  wire       [0:0]    all_zeros_204;
  wire       [0:0]    all_left_zeros_204;
  wire       [1:0]    left_all_zeros_count_100;
  wire       [0:0]    _zz_317;
  wire       [0:0]    _zz_318;
  wire       [0:0]    all_zeros_205;
  wire       [0:0]    all_left_zeros_205;
  wire       [1:0]    left_non_all_zeros_count_97;
  wire       [1:0]    non_zeros_lzc_97;
  wire       [2:0]    left_all_zeros_count_101;
  wire       [1:0]    _zz_319;
  wire       [1:0]    all_zeros_206;
  wire       [1:0]    all_left_zeros_206;
  wire       [1:0]    whole_bit_count_104;
  wire       [1:0]    left_bit_count_104;
  wire       [0:0]    _zz_320;
  wire       [0:0]    _zz_321;
  wire       [0:0]    all_zeros_207;
  wire       [0:0]    all_left_zeros_207;
  wire       [1:0]    left_all_zeros_count_102;
  wire       [0:0]    _zz_322;
  wire       [0:0]    _zz_323;
  wire       [0:0]    all_zeros_208;
  wire       [0:0]    all_left_zeros_208;
  wire       [1:0]    left_non_all_zeros_count_98;
  wire       [1:0]    non_zeros_lzc_98;
  wire       [2:0]    left_non_all_zeros_count_99;
  wire       [2:0]    non_zeros_lzc_99;
  wire       [3:0]    left_non_all_zeros_count_100;
  wire       [3:0]    non_zeros_lzc_100;
  wire       [4:0]    left_all_zeros_count_103;
  wire       [7:0]    _zz_324;
  wire       [3:0]    all_zeros_209;
  wire       [3:0]    all_left_zeros_209;
  wire       [3:0]    whole_bit_count_105;
  wire       [3:0]    left_bit_count_105;
  wire       [3:0]    _zz_325;
  wire       [2:0]    all_zeros_210;
  wire       [2:0]    all_left_zeros_210;
  wire       [2:0]    whole_bit_count_106;
  wire       [2:0]    left_bit_count_106;
  wire       [1:0]    _zz_326;
  wire       [1:0]    all_zeros_211;
  wire       [1:0]    all_left_zeros_211;
  wire       [1:0]    whole_bit_count_107;
  wire       [1:0]    left_bit_count_107;
  wire       [0:0]    _zz_327;
  wire       [0:0]    _zz_328;
  wire       [0:0]    all_zeros_212;
  wire       [0:0]    all_left_zeros_212;
  wire       [1:0]    left_all_zeros_count_104;
  wire       [0:0]    _zz_329;
  wire       [0:0]    _zz_330;
  wire       [0:0]    all_zeros_213;
  wire       [0:0]    all_left_zeros_213;
  wire       [1:0]    left_non_all_zeros_count_101;
  wire       [1:0]    non_zeros_lzc_101;
  wire       [2:0]    left_all_zeros_count_105;
  wire       [1:0]    _zz_331;
  wire       [1:0]    all_zeros_214;
  wire       [1:0]    all_left_zeros_214;
  wire       [1:0]    whole_bit_count_108;
  wire       [1:0]    left_bit_count_108;
  wire       [0:0]    _zz_332;
  wire       [0:0]    _zz_333;
  wire       [0:0]    all_zeros_215;
  wire       [0:0]    all_left_zeros_215;
  wire       [1:0]    left_all_zeros_count_106;
  wire       [0:0]    _zz_334;
  wire       [0:0]    _zz_335;
  wire       [0:0]    all_zeros_216;
  wire       [0:0]    all_left_zeros_216;
  wire       [1:0]    left_non_all_zeros_count_102;
  wire       [1:0]    non_zeros_lzc_102;
  wire       [2:0]    left_non_all_zeros_count_103;
  wire       [2:0]    non_zeros_lzc_103;
  wire       [3:0]    left_all_zeros_count_107;
  wire       [3:0]    _zz_336;
  wire       [2:0]    all_zeros_217;
  wire       [2:0]    all_left_zeros_217;
  wire       [2:0]    whole_bit_count_109;
  wire       [2:0]    left_bit_count_109;
  wire       [1:0]    _zz_337;
  wire       [1:0]    all_zeros_218;
  wire       [1:0]    all_left_zeros_218;
  wire       [1:0]    whole_bit_count_110;
  wire       [1:0]    left_bit_count_110;
  wire       [0:0]    _zz_338;
  wire       [0:0]    _zz_339;
  wire       [0:0]    all_zeros_219;
  wire       [0:0]    all_left_zeros_219;
  wire       [1:0]    left_all_zeros_count_108;
  wire       [0:0]    _zz_340;
  wire       [0:0]    _zz_341;
  wire       [0:0]    all_zeros_220;
  wire       [0:0]    all_left_zeros_220;
  wire       [1:0]    left_non_all_zeros_count_104;
  wire       [1:0]    non_zeros_lzc_104;
  wire       [2:0]    left_all_zeros_count_109;
  wire       [1:0]    _zz_342;
  wire       [1:0]    all_zeros_221;
  wire       [1:0]    all_left_zeros_221;
  wire       [1:0]    whole_bit_count_111;
  wire       [1:0]    left_bit_count_111;
  wire       [0:0]    _zz_343;
  wire       [0:0]    _zz_344;
  wire       [0:0]    all_zeros_222;
  wire       [0:0]    all_left_zeros_222;
  wire       [1:0]    left_all_zeros_count_110;
  wire       [0:0]    _zz_345;
  wire       [0:0]    _zz_346;
  wire       [0:0]    all_zeros_223;
  wire       [0:0]    all_left_zeros_223;
  wire       [1:0]    left_non_all_zeros_count_105;
  wire       [1:0]    non_zeros_lzc_105;
  wire       [2:0]    left_non_all_zeros_count_106;
  wire       [2:0]    non_zeros_lzc_106;
  wire       [3:0]    left_non_all_zeros_count_107;
  wire       [3:0]    non_zeros_lzc_107;
  wire       [4:0]    left_non_all_zeros_count_108;
  wire       [4:0]    non_zeros_lzc_108;
  wire       [5:0]    left_all_zeros_count_111;
  wire       [15:0]   _zz_347;
  wire       [4:0]    all_zeros_224;
  wire       [4:0]    all_left_zeros_224;
  wire       [4:0]    whole_bit_count_112;
  wire       [4:0]    left_bit_count_112;
  wire       [7:0]    _zz_348;
  wire       [3:0]    all_zeros_225;
  wire       [3:0]    all_left_zeros_225;
  wire       [3:0]    whole_bit_count_113;
  wire       [3:0]    left_bit_count_113;
  wire       [3:0]    _zz_349;
  wire       [2:0]    all_zeros_226;
  wire       [2:0]    all_left_zeros_226;
  wire       [2:0]    whole_bit_count_114;
  wire       [2:0]    left_bit_count_114;
  wire       [1:0]    _zz_350;
  wire       [1:0]    all_zeros_227;
  wire       [1:0]    all_left_zeros_227;
  wire       [1:0]    whole_bit_count_115;
  wire       [1:0]    left_bit_count_115;
  wire       [0:0]    _zz_351;
  wire       [0:0]    _zz_352;
  wire       [0:0]    all_zeros_228;
  wire       [0:0]    all_left_zeros_228;
  wire       [1:0]    left_all_zeros_count_112;
  wire       [0:0]    _zz_353;
  wire       [0:0]    _zz_354;
  wire       [0:0]    all_zeros_229;
  wire       [0:0]    all_left_zeros_229;
  wire       [1:0]    left_non_all_zeros_count_109;
  wire       [1:0]    non_zeros_lzc_109;
  wire       [2:0]    left_all_zeros_count_113;
  wire       [1:0]    _zz_355;
  wire       [1:0]    all_zeros_230;
  wire       [1:0]    all_left_zeros_230;
  wire       [1:0]    whole_bit_count_116;
  wire       [1:0]    left_bit_count_116;
  wire       [0:0]    _zz_356;
  wire       [0:0]    _zz_357;
  wire       [0:0]    all_zeros_231;
  wire       [0:0]    all_left_zeros_231;
  wire       [1:0]    left_all_zeros_count_114;
  wire       [0:0]    _zz_358;
  wire       [0:0]    _zz_359;
  wire       [0:0]    all_zeros_232;
  wire       [0:0]    all_left_zeros_232;
  wire       [1:0]    left_non_all_zeros_count_110;
  wire       [1:0]    non_zeros_lzc_110;
  wire       [2:0]    left_non_all_zeros_count_111;
  wire       [2:0]    non_zeros_lzc_111;
  wire       [3:0]    left_all_zeros_count_115;
  wire       [3:0]    _zz_360;
  wire       [2:0]    all_zeros_233;
  wire       [2:0]    all_left_zeros_233;
  wire       [2:0]    whole_bit_count_117;
  wire       [2:0]    left_bit_count_117;
  wire       [1:0]    _zz_361;
  wire       [1:0]    all_zeros_234;
  wire       [1:0]    all_left_zeros_234;
  wire       [1:0]    whole_bit_count_118;
  wire       [1:0]    left_bit_count_118;
  wire       [0:0]    _zz_362;
  wire       [0:0]    _zz_363;
  wire       [0:0]    all_zeros_235;
  wire       [0:0]    all_left_zeros_235;
  wire       [1:0]    left_all_zeros_count_116;
  wire       [0:0]    _zz_364;
  wire       [0:0]    _zz_365;
  wire       [0:0]    all_zeros_236;
  wire       [0:0]    all_left_zeros_236;
  wire       [1:0]    left_non_all_zeros_count_112;
  wire       [1:0]    non_zeros_lzc_112;
  wire       [2:0]    left_all_zeros_count_117;
  wire       [1:0]    _zz_366;
  wire       [1:0]    all_zeros_237;
  wire       [1:0]    all_left_zeros_237;
  wire       [1:0]    whole_bit_count_119;
  wire       [1:0]    left_bit_count_119;
  wire       [0:0]    _zz_367;
  wire       [0:0]    _zz_368;
  wire       [0:0]    all_zeros_238;
  wire       [0:0]    all_left_zeros_238;
  wire       [1:0]    left_all_zeros_count_118;
  wire       [0:0]    _zz_369;
  wire       [0:0]    _zz_370;
  wire       [0:0]    all_zeros_239;
  wire       [0:0]    all_left_zeros_239;
  wire       [1:0]    left_non_all_zeros_count_113;
  wire       [1:0]    non_zeros_lzc_113;
  wire       [2:0]    left_non_all_zeros_count_114;
  wire       [2:0]    non_zeros_lzc_114;
  wire       [3:0]    left_non_all_zeros_count_115;
  wire       [3:0]    non_zeros_lzc_115;
  wire       [4:0]    left_all_zeros_count_119;
  wire       [7:0]    _zz_371;
  wire       [3:0]    all_zeros_240;
  wire       [3:0]    all_left_zeros_240;
  wire       [3:0]    whole_bit_count_120;
  wire       [3:0]    left_bit_count_120;
  wire       [3:0]    _zz_372;
  wire       [2:0]    all_zeros_241;
  wire       [2:0]    all_left_zeros_241;
  wire       [2:0]    whole_bit_count_121;
  wire       [2:0]    left_bit_count_121;
  wire       [1:0]    _zz_373;
  wire       [1:0]    all_zeros_242;
  wire       [1:0]    all_left_zeros_242;
  wire       [1:0]    whole_bit_count_122;
  wire       [1:0]    left_bit_count_122;
  wire       [0:0]    _zz_374;
  wire       [0:0]    _zz_375;
  wire       [0:0]    all_zeros_243;
  wire       [0:0]    all_left_zeros_243;
  wire       [1:0]    left_all_zeros_count_120;
  wire       [0:0]    _zz_376;
  wire       [0:0]    _zz_377;
  wire       [0:0]    all_zeros_244;
  wire       [0:0]    all_left_zeros_244;
  wire       [1:0]    left_non_all_zeros_count_116;
  wire       [1:0]    non_zeros_lzc_116;
  wire       [2:0]    left_all_zeros_count_121;
  wire       [1:0]    _zz_378;
  wire       [1:0]    all_zeros_245;
  wire       [1:0]    all_left_zeros_245;
  wire       [1:0]    whole_bit_count_123;
  wire       [1:0]    left_bit_count_123;
  wire       [0:0]    _zz_379;
  wire       [0:0]    _zz_380;
  wire       [0:0]    all_zeros_246;
  wire       [0:0]    all_left_zeros_246;
  wire       [1:0]    left_all_zeros_count_122;
  wire       [0:0]    _zz_381;
  wire       [0:0]    _zz_382;
  wire       [0:0]    all_zeros_247;
  wire       [0:0]    all_left_zeros_247;
  wire       [1:0]    left_non_all_zeros_count_117;
  wire       [1:0]    non_zeros_lzc_117;
  wire       [2:0]    left_non_all_zeros_count_118;
  wire       [2:0]    non_zeros_lzc_118;
  wire       [3:0]    left_all_zeros_count_123;
  wire       [3:0]    _zz_383;
  wire       [2:0]    all_zeros_248;
  wire       [2:0]    all_left_zeros_248;
  wire       [2:0]    whole_bit_count_124;
  wire       [2:0]    left_bit_count_124;
  wire       [1:0]    _zz_384;
  wire       [1:0]    all_zeros_249;
  wire       [1:0]    all_left_zeros_249;
  wire       [1:0]    whole_bit_count_125;
  wire       [1:0]    left_bit_count_125;
  wire       [0:0]    _zz_385;
  wire       [0:0]    _zz_386;
  wire       [0:0]    all_zeros_250;
  wire       [0:0]    all_left_zeros_250;
  wire       [1:0]    left_all_zeros_count_124;
  wire       [0:0]    _zz_387;
  wire       [0:0]    _zz_388;
  wire       [0:0]    all_zeros_251;
  wire       [0:0]    all_left_zeros_251;
  wire       [1:0]    left_non_all_zeros_count_119;
  wire       [1:0]    non_zeros_lzc_119;
  wire       [2:0]    left_all_zeros_count_125;
  wire       [1:0]    _zz_389;
  wire       [1:0]    all_zeros_252;
  wire       [1:0]    all_left_zeros_252;
  wire       [1:0]    whole_bit_count_126;
  wire       [1:0]    left_bit_count_126;
  wire       [0:0]    _zz_390;
  wire       [0:0]    _zz_391;
  wire       [0:0]    all_zeros_253;
  wire       [0:0]    all_left_zeros_253;
  wire       [1:0]    left_all_zeros_count_126;
  wire       [0:0]    _zz_392;
  wire       [0:0]    _zz_393;
  wire       [0:0]    all_zeros_254;
  wire       [0:0]    all_left_zeros_254;
  wire       [1:0]    left_non_all_zeros_count_120;
  wire       [1:0]    non_zeros_lzc_120;
  wire       [2:0]    left_non_all_zeros_count_121;
  wire       [2:0]    non_zeros_lzc_121;
  wire       [3:0]    left_non_all_zeros_count_122;
  wire       [3:0]    non_zeros_lzc_122;
  wire       [4:0]    left_non_all_zeros_count_123;
  wire       [4:0]    non_zeros_lzc_123;
  wire       [5:0]    left_non_all_zeros_count_124;
  wire       [5:0]    non_zeros_lzc_124;
  wire       [6:0]    left_non_all_zeros_count_125;
  wire       [6:0]    non_zeros_lzc_125;
  wire       [7:0]    left_non_all_zeros_count_126;
  wire       [7:0]    non_zeros_lzc_126;
  reg        [7:0]    _zz_394;
  wire       [6:0]    lzc;
  reg        [31:0]   exp_wd_prod_real;
  reg        [31:0]   exp_wd_prod_imag;
  wire       [6:0]    _zz_395;
  wire       [7:0]    _zz_396;
  wire       [15:0]   _zz_397;
  wire       [15:0]   _zz_398;
  wire       [7:0]    _zz_399;
  wire       [15:0]   _zz_400;
  wire       [15:0]   _zz_401;
  wire       [7:0]    _zz_402;
  wire       [7:0]    _zz_403;
  wire       [15:0]   _zz_404;
  reg        [31:0]   _zz_405;
  reg        [31:0]   _zz_406;
  reg        [15:0]   func_table_0_regNext_real;
  reg        [15:0]   func_table_0_regNext_imag;
  reg        [15:0]   func_table_127_regNext_real;
  reg        [15:0]   func_table_127_regNext_imag;
  wire       [15:0]   _zz_407;
  reg        [15:0]   wave_regNext;
  reg        [15:0]   _zz_408;
  reg        [15:0]   _zz_409;
  reg        [31:0]   exp_wd_prod_divw_real;
  reg        [31:0]   exp_wd_prod_divw_imag;
  wire       [31:0]   _zz_410;
  reg        [63:0]   _zz_411;
  reg        [63:0]   _zz_412;

  assign _zz_453 = ((lzc != 7'h0) && (_zz_1474 < 8'h80));
  assign _zz_454 = (lzc == 7'h0);
  assign _zz_455 = fixTo_dout;
  assign _zz_456 = wd_prod;
  assign _zz_457 = {8'd0, _zz_456};
  assign _zz_458 = wd_prod;
  assign _zz_459 = {8'd0, _zz_458};
  assign _zz_460 = wd_prod;
  assign _zz_461 = {8'd0, _zz_460};
  assign _zz_462 = wd_prod;
  assign _zz_463 = {8'd0, _zz_462};
  assign _zz_464 = wd_prod;
  assign _zz_465 = {8'd0, _zz_464};
  assign _zz_466 = wd_prod;
  assign _zz_467 = {8'd0, _zz_466};
  assign _zz_468 = wd_prod;
  assign _zz_469 = {8'd0, _zz_468};
  assign _zz_470 = wd_prod;
  assign _zz_471 = {8'd0, _zz_470};
  assign _zz_472 = wd_prod;
  assign _zz_473 = {8'd0, _zz_472};
  assign _zz_474 = wd_prod;
  assign _zz_475 = {8'd0, _zz_474};
  assign _zz_476 = wd_prod;
  assign _zz_477 = {8'd0, _zz_476};
  assign _zz_478 = wd_prod;
  assign _zz_479 = {8'd0, _zz_478};
  assign _zz_480 = wd_prod;
  assign _zz_481 = {8'd0, _zz_480};
  assign _zz_482 = wd_prod;
  assign _zz_483 = {8'd0, _zz_482};
  assign _zz_484 = wd_prod;
  assign _zz_485 = {8'd0, _zz_484};
  assign _zz_486 = wd_prod;
  assign _zz_487 = {8'd0, _zz_486};
  assign _zz_488 = wd_prod;
  assign _zz_489 = {8'd0, _zz_488};
  assign _zz_490 = wd_prod;
  assign _zz_491 = {8'd0, _zz_490};
  assign _zz_492 = wd_prod;
  assign _zz_493 = {8'd0, _zz_492};
  assign _zz_494 = wd_prod;
  assign _zz_495 = {8'd0, _zz_494};
  assign _zz_496 = wd_prod;
  assign _zz_497 = {8'd0, _zz_496};
  assign _zz_498 = wd_prod;
  assign _zz_499 = {8'd0, _zz_498};
  assign _zz_500 = wd_prod;
  assign _zz_501 = {8'd0, _zz_500};
  assign _zz_502 = wd_prod;
  assign _zz_503 = {8'd0, _zz_502};
  assign _zz_504 = wd_prod;
  assign _zz_505 = {8'd0, _zz_504};
  assign _zz_506 = wd_prod;
  assign _zz_507 = {8'd0, _zz_506};
  assign _zz_508 = wd_prod;
  assign _zz_509 = {8'd0, _zz_508};
  assign _zz_510 = wd_prod;
  assign _zz_511 = {8'd0, _zz_510};
  assign _zz_512 = wd_prod;
  assign _zz_513 = {8'd0, _zz_512};
  assign _zz_514 = wd_prod;
  assign _zz_515 = {8'd0, _zz_514};
  assign _zz_516 = wd_prod;
  assign _zz_517 = {8'd0, _zz_516};
  assign _zz_518 = wd_prod;
  assign _zz_519 = {8'd0, _zz_518};
  assign _zz_520 = wd_prod;
  assign _zz_521 = {8'd0, _zz_520};
  assign _zz_522 = wd_prod;
  assign _zz_523 = {8'd0, _zz_522};
  assign _zz_524 = wd_prod;
  assign _zz_525 = {8'd0, _zz_524};
  assign _zz_526 = wd_prod;
  assign _zz_527 = {8'd0, _zz_526};
  assign _zz_528 = wd_prod;
  assign _zz_529 = {8'd0, _zz_528};
  assign _zz_530 = wd_prod;
  assign _zz_531 = {8'd0, _zz_530};
  assign _zz_532 = wd_prod;
  assign _zz_533 = {8'd0, _zz_532};
  assign _zz_534 = wd_prod;
  assign _zz_535 = {8'd0, _zz_534};
  assign _zz_536 = wd_prod;
  assign _zz_537 = {8'd0, _zz_536};
  assign _zz_538 = wd_prod;
  assign _zz_539 = {8'd0, _zz_538};
  assign _zz_540 = wd_prod;
  assign _zz_541 = {8'd0, _zz_540};
  assign _zz_542 = wd_prod;
  assign _zz_543 = {8'd0, _zz_542};
  assign _zz_544 = wd_prod;
  assign _zz_545 = {8'd0, _zz_544};
  assign _zz_546 = wd_prod;
  assign _zz_547 = {8'd0, _zz_546};
  assign _zz_548 = wd_prod;
  assign _zz_549 = {8'd0, _zz_548};
  assign _zz_550 = wd_prod;
  assign _zz_551 = {8'd0, _zz_550};
  assign _zz_552 = wd_prod;
  assign _zz_553 = {8'd0, _zz_552};
  assign _zz_554 = wd_prod;
  assign _zz_555 = {8'd0, _zz_554};
  assign _zz_556 = wd_prod;
  assign _zz_557 = {8'd0, _zz_556};
  assign _zz_558 = wd_prod;
  assign _zz_559 = {8'd0, _zz_558};
  assign _zz_560 = wd_prod;
  assign _zz_561 = {8'd0, _zz_560};
  assign _zz_562 = wd_prod;
  assign _zz_563 = {8'd0, _zz_562};
  assign _zz_564 = wd_prod;
  assign _zz_565 = {8'd0, _zz_564};
  assign _zz_566 = wd_prod;
  assign _zz_567 = {8'd0, _zz_566};
  assign _zz_568 = wd_prod;
  assign _zz_569 = {8'd0, _zz_568};
  assign _zz_570 = wd_prod;
  assign _zz_571 = {8'd0, _zz_570};
  assign _zz_572 = wd_prod;
  assign _zz_573 = {8'd0, _zz_572};
  assign _zz_574 = wd_prod;
  assign _zz_575 = {8'd0, _zz_574};
  assign _zz_576 = wd_prod;
  assign _zz_577 = {8'd0, _zz_576};
  assign _zz_578 = wd_prod;
  assign _zz_579 = {8'd0, _zz_578};
  assign _zz_580 = wd_prod;
  assign _zz_581 = {8'd0, _zz_580};
  assign _zz_582 = wd_prod;
  assign _zz_583 = {8'd0, _zz_582};
  assign _zz_584 = wd_prod;
  assign _zz_585 = {8'd0, _zz_584};
  assign _zz_586 = wd_prod;
  assign _zz_587 = {8'd0, _zz_586};
  assign _zz_588 = wd_prod;
  assign _zz_589 = {8'd0, _zz_588};
  assign _zz_590 = wd_prod;
  assign _zz_591 = {8'd0, _zz_590};
  assign _zz_592 = wd_prod;
  assign _zz_593 = {8'd0, _zz_592};
  assign _zz_594 = wd_prod;
  assign _zz_595 = {8'd0, _zz_594};
  assign _zz_596 = wd_prod;
  assign _zz_597 = {8'd0, _zz_596};
  assign _zz_598 = wd_prod;
  assign _zz_599 = {8'd0, _zz_598};
  assign _zz_600 = wd_prod;
  assign _zz_601 = {8'd0, _zz_600};
  assign _zz_602 = wd_prod;
  assign _zz_603 = {8'd0, _zz_602};
  assign _zz_604 = wd_prod;
  assign _zz_605 = {8'd0, _zz_604};
  assign _zz_606 = wd_prod;
  assign _zz_607 = {8'd0, _zz_606};
  assign _zz_608 = wd_prod;
  assign _zz_609 = {8'd0, _zz_608};
  assign _zz_610 = wd_prod;
  assign _zz_611 = {8'd0, _zz_610};
  assign _zz_612 = wd_prod;
  assign _zz_613 = {8'd0, _zz_612};
  assign _zz_614 = wd_prod;
  assign _zz_615 = {8'd0, _zz_614};
  assign _zz_616 = wd_prod;
  assign _zz_617 = {8'd0, _zz_616};
  assign _zz_618 = wd_prod;
  assign _zz_619 = {8'd0, _zz_618};
  assign _zz_620 = wd_prod;
  assign _zz_621 = {8'd0, _zz_620};
  assign _zz_622 = wd_prod;
  assign _zz_623 = {8'd0, _zz_622};
  assign _zz_624 = wd_prod;
  assign _zz_625 = {8'd0, _zz_624};
  assign _zz_626 = wd_prod;
  assign _zz_627 = {8'd0, _zz_626};
  assign _zz_628 = wd_prod;
  assign _zz_629 = {8'd0, _zz_628};
  assign _zz_630 = wd_prod;
  assign _zz_631 = {8'd0, _zz_630};
  assign _zz_632 = wd_prod;
  assign _zz_633 = {8'd0, _zz_632};
  assign _zz_634 = wd_prod;
  assign _zz_635 = {8'd0, _zz_634};
  assign _zz_636 = wd_prod;
  assign _zz_637 = {8'd0, _zz_636};
  assign _zz_638 = wd_prod;
  assign _zz_639 = {8'd0, _zz_638};
  assign _zz_640 = wd_prod;
  assign _zz_641 = {8'd0, _zz_640};
  assign _zz_642 = wd_prod;
  assign _zz_643 = {8'd0, _zz_642};
  assign _zz_644 = wd_prod;
  assign _zz_645 = {8'd0, _zz_644};
  assign _zz_646 = wd_prod;
  assign _zz_647 = {8'd0, _zz_646};
  assign _zz_648 = wd_prod;
  assign _zz_649 = {8'd0, _zz_648};
  assign _zz_650 = wd_prod;
  assign _zz_651 = {8'd0, _zz_650};
  assign _zz_652 = wd_prod;
  assign _zz_653 = {8'd0, _zz_652};
  assign _zz_654 = wd_prod;
  assign _zz_655 = {8'd0, _zz_654};
  assign _zz_656 = wd_prod;
  assign _zz_657 = {8'd0, _zz_656};
  assign _zz_658 = wd_prod;
  assign _zz_659 = {8'd0, _zz_658};
  assign _zz_660 = wd_prod;
  assign _zz_661 = {8'd0, _zz_660};
  assign _zz_662 = wd_prod;
  assign _zz_663 = {8'd0, _zz_662};
  assign _zz_664 = wd_prod;
  assign _zz_665 = {8'd0, _zz_664};
  assign _zz_666 = wd_prod;
  assign _zz_667 = {8'd0, _zz_666};
  assign _zz_668 = wd_prod;
  assign _zz_669 = {8'd0, _zz_668};
  assign _zz_670 = wd_prod;
  assign _zz_671 = {8'd0, _zz_670};
  assign _zz_672 = wd_prod;
  assign _zz_673 = {8'd0, _zz_672};
  assign _zz_674 = wd_prod;
  assign _zz_675 = {8'd0, _zz_674};
  assign _zz_676 = wd_prod;
  assign _zz_677 = {8'd0, _zz_676};
  assign _zz_678 = wd_prod;
  assign _zz_679 = {8'd0, _zz_678};
  assign _zz_680 = wd_prod;
  assign _zz_681 = {8'd0, _zz_680};
  assign _zz_682 = wd_prod;
  assign _zz_683 = {8'd0, _zz_682};
  assign _zz_684 = wd_prod;
  assign _zz_685 = {8'd0, _zz_684};
  assign _zz_686 = wd_prod;
  assign _zz_687 = {8'd0, _zz_686};
  assign _zz_688 = wd_prod;
  assign _zz_689 = {8'd0, _zz_688};
  assign _zz_690 = wd_prod;
  assign _zz_691 = {8'd0, _zz_690};
  assign _zz_692 = wd_prod;
  assign _zz_693 = {8'd0, _zz_692};
  assign _zz_694 = wd_prod;
  assign _zz_695 = {8'd0, _zz_694};
  assign _zz_696 = wd_prod;
  assign _zz_697 = {8'd0, _zz_696};
  assign _zz_698 = wd_prod;
  assign _zz_699 = {8'd0, _zz_698};
  assign _zz_700 = wd_prod;
  assign _zz_701 = {8'd0, _zz_700};
  assign _zz_702 = wd_prod;
  assign _zz_703 = {8'd0, _zz_702};
  assign _zz_704 = wd_prod;
  assign _zz_705 = {8'd0, _zz_704};
  assign _zz_706 = wd_prod;
  assign _zz_707 = {8'd0, _zz_706};
  assign _zz_708 = wd_prod;
  assign _zz_709 = {8'd0, _zz_708};
  assign _zz_710 = wd_prod;
  assign _zz_711 = {8'd0, _zz_710};
  assign _zz_712 = (left_bit_count_6 + _zz_714);
  assign _zz_713 = _zz_18[0];
  assign _zz_714 = {1'd0, _zz_713};
  assign _zz_715 = _zz_20[0];
  assign _zz_716 = {1'd0, _zz_715};
  assign _zz_717 = (left_bit_count_5 + _zz_719);
  assign _zz_718 = ((all_zeros_6 & _zz_720) & non_zeros_lzc);
  assign _zz_719 = {1'd0, _zz_718};
  assign _zz_720 = (whole_bit_count_6 + (~ all_zeros_6));
  assign _zz_721 = (left_bit_count_7 + _zz_723);
  assign _zz_722 = _zz_23[0];
  assign _zz_723 = {1'd0, _zz_722};
  assign _zz_724 = _zz_25[0];
  assign _zz_725 = {1'd0, _zz_724};
  assign _zz_726 = ((all_zeros_9 & _zz_728) & non_zeros_lzc_1);
  assign _zz_727 = {1'd0, _zz_726};
  assign _zz_728 = (whole_bit_count_7 + (~ all_zeros_9));
  assign _zz_729 = (left_bit_count_4 + _zz_731);
  assign _zz_730 = ((all_zeros_5 & _zz_732) & non_zeros_lzc_2);
  assign _zz_731 = {1'd0, _zz_730};
  assign _zz_732 = (whole_bit_count_5 + (~ all_zeros_5));
  assign _zz_733 = (left_bit_count_9 + _zz_735);
  assign _zz_734 = _zz_29[0];
  assign _zz_735 = {1'd0, _zz_734};
  assign _zz_736 = _zz_31[0];
  assign _zz_737 = {1'd0, _zz_736};
  assign _zz_738 = (left_bit_count_8 + _zz_740);
  assign _zz_739 = ((all_zeros_13 & _zz_741) & non_zeros_lzc_3);
  assign _zz_740 = {1'd0, _zz_739};
  assign _zz_741 = (whole_bit_count_9 + (~ all_zeros_13));
  assign _zz_742 = (left_bit_count_10 + _zz_744);
  assign _zz_743 = _zz_34[0];
  assign _zz_744 = {1'd0, _zz_743};
  assign _zz_745 = _zz_36[0];
  assign _zz_746 = {1'd0, _zz_745};
  assign _zz_747 = ((all_zeros_16 & _zz_749) & non_zeros_lzc_4);
  assign _zz_748 = {1'd0, _zz_747};
  assign _zz_749 = (whole_bit_count_10 + (~ all_zeros_16));
  assign _zz_750 = ((all_zeros_12 & _zz_752) & non_zeros_lzc_5);
  assign _zz_751 = {1'd0, _zz_750};
  assign _zz_752 = (whole_bit_count_8 + (~ all_zeros_12));
  assign _zz_753 = (left_bit_count_3 + _zz_755);
  assign _zz_754 = ((all_zeros_4 & _zz_756) & non_zeros_lzc_6);
  assign _zz_755 = {1'd0, _zz_754};
  assign _zz_756 = (whole_bit_count_4 + (~ all_zeros_4));
  assign _zz_757 = (left_bit_count_13 + _zz_759);
  assign _zz_758 = _zz_41[0];
  assign _zz_759 = {1'd0, _zz_758};
  assign _zz_760 = _zz_43[0];
  assign _zz_761 = {1'd0, _zz_760};
  assign _zz_762 = (left_bit_count_12 + _zz_764);
  assign _zz_763 = ((all_zeros_21 & _zz_765) & non_zeros_lzc_7);
  assign _zz_764 = {1'd0, _zz_763};
  assign _zz_765 = (whole_bit_count_13 + (~ all_zeros_21));
  assign _zz_766 = (left_bit_count_14 + _zz_768);
  assign _zz_767 = _zz_46[0];
  assign _zz_768 = {1'd0, _zz_767};
  assign _zz_769 = _zz_48[0];
  assign _zz_770 = {1'd0, _zz_769};
  assign _zz_771 = ((all_zeros_24 & _zz_773) & non_zeros_lzc_8);
  assign _zz_772 = {1'd0, _zz_771};
  assign _zz_773 = (whole_bit_count_14 + (~ all_zeros_24));
  assign _zz_774 = (left_bit_count_11 + _zz_776);
  assign _zz_775 = ((all_zeros_20 & _zz_777) & non_zeros_lzc_9);
  assign _zz_776 = {1'd0, _zz_775};
  assign _zz_777 = (whole_bit_count_12 + (~ all_zeros_20));
  assign _zz_778 = (left_bit_count_16 + _zz_780);
  assign _zz_779 = _zz_52[0];
  assign _zz_780 = {1'd0, _zz_779};
  assign _zz_781 = _zz_54[0];
  assign _zz_782 = {1'd0, _zz_781};
  assign _zz_783 = (left_bit_count_15 + _zz_785);
  assign _zz_784 = ((all_zeros_28 & _zz_786) & non_zeros_lzc_10);
  assign _zz_785 = {1'd0, _zz_784};
  assign _zz_786 = (whole_bit_count_16 + (~ all_zeros_28));
  assign _zz_787 = (left_bit_count_17 + _zz_789);
  assign _zz_788 = _zz_57[0];
  assign _zz_789 = {1'd0, _zz_788};
  assign _zz_790 = _zz_59[0];
  assign _zz_791 = {1'd0, _zz_790};
  assign _zz_792 = ((all_zeros_31 & _zz_794) & non_zeros_lzc_11);
  assign _zz_793 = {1'd0, _zz_792};
  assign _zz_794 = (whole_bit_count_17 + (~ all_zeros_31));
  assign _zz_795 = ((all_zeros_27 & _zz_797) & non_zeros_lzc_12);
  assign _zz_796 = {1'd0, _zz_795};
  assign _zz_797 = (whole_bit_count_15 + (~ all_zeros_27));
  assign _zz_798 = ((all_zeros_19 & _zz_800) & non_zeros_lzc_13);
  assign _zz_799 = {1'd0, _zz_798};
  assign _zz_800 = (whole_bit_count_11 + (~ all_zeros_19));
  assign _zz_801 = (left_bit_count_2 + _zz_803);
  assign _zz_802 = ((all_zeros_3 & _zz_804) & non_zeros_lzc_14);
  assign _zz_803 = {1'd0, _zz_802};
  assign _zz_804 = (whole_bit_count_3 + (~ all_zeros_3));
  assign _zz_805 = (left_bit_count_21 + _zz_807);
  assign _zz_806 = _zz_65[0];
  assign _zz_807 = {1'd0, _zz_806};
  assign _zz_808 = _zz_67[0];
  assign _zz_809 = {1'd0, _zz_808};
  assign _zz_810 = (left_bit_count_20 + _zz_812);
  assign _zz_811 = ((all_zeros_37 & _zz_813) & non_zeros_lzc_15);
  assign _zz_812 = {1'd0, _zz_811};
  assign _zz_813 = (whole_bit_count_21 + (~ all_zeros_37));
  assign _zz_814 = (left_bit_count_22 + _zz_816);
  assign _zz_815 = _zz_70[0];
  assign _zz_816 = {1'd0, _zz_815};
  assign _zz_817 = _zz_72[0];
  assign _zz_818 = {1'd0, _zz_817};
  assign _zz_819 = ((all_zeros_40 & _zz_821) & non_zeros_lzc_16);
  assign _zz_820 = {1'd0, _zz_819};
  assign _zz_821 = (whole_bit_count_22 + (~ all_zeros_40));
  assign _zz_822 = (left_bit_count_19 + _zz_824);
  assign _zz_823 = ((all_zeros_36 & _zz_825) & non_zeros_lzc_17);
  assign _zz_824 = {1'd0, _zz_823};
  assign _zz_825 = (whole_bit_count_20 + (~ all_zeros_36));
  assign _zz_826 = (left_bit_count_24 + _zz_828);
  assign _zz_827 = _zz_76[0];
  assign _zz_828 = {1'd0, _zz_827};
  assign _zz_829 = _zz_78[0];
  assign _zz_830 = {1'd0, _zz_829};
  assign _zz_831 = (left_bit_count_23 + _zz_833);
  assign _zz_832 = ((all_zeros_44 & _zz_834) & non_zeros_lzc_18);
  assign _zz_833 = {1'd0, _zz_832};
  assign _zz_834 = (whole_bit_count_24 + (~ all_zeros_44));
  assign _zz_835 = (left_bit_count_25 + _zz_837);
  assign _zz_836 = _zz_81[0];
  assign _zz_837 = {1'd0, _zz_836};
  assign _zz_838 = _zz_83[0];
  assign _zz_839 = {1'd0, _zz_838};
  assign _zz_840 = ((all_zeros_47 & _zz_842) & non_zeros_lzc_19);
  assign _zz_841 = {1'd0, _zz_840};
  assign _zz_842 = (whole_bit_count_25 + (~ all_zeros_47));
  assign _zz_843 = ((all_zeros_43 & _zz_845) & non_zeros_lzc_20);
  assign _zz_844 = {1'd0, _zz_843};
  assign _zz_845 = (whole_bit_count_23 + (~ all_zeros_43));
  assign _zz_846 = (left_bit_count_18 + _zz_848);
  assign _zz_847 = ((all_zeros_35 & _zz_849) & non_zeros_lzc_21);
  assign _zz_848 = {1'd0, _zz_847};
  assign _zz_849 = (whole_bit_count_19 + (~ all_zeros_35));
  assign _zz_850 = (left_bit_count_28 + _zz_852);
  assign _zz_851 = _zz_88[0];
  assign _zz_852 = {1'd0, _zz_851};
  assign _zz_853 = _zz_90[0];
  assign _zz_854 = {1'd0, _zz_853};
  assign _zz_855 = (left_bit_count_27 + _zz_857);
  assign _zz_856 = ((all_zeros_52 & _zz_858) & non_zeros_lzc_22);
  assign _zz_857 = {1'd0, _zz_856};
  assign _zz_858 = (whole_bit_count_28 + (~ all_zeros_52));
  assign _zz_859 = (left_bit_count_29 + _zz_861);
  assign _zz_860 = _zz_93[0];
  assign _zz_861 = {1'd0, _zz_860};
  assign _zz_862 = _zz_95[0];
  assign _zz_863 = {1'd0, _zz_862};
  assign _zz_864 = ((all_zeros_55 & _zz_866) & non_zeros_lzc_23);
  assign _zz_865 = {1'd0, _zz_864};
  assign _zz_866 = (whole_bit_count_29 + (~ all_zeros_55));
  assign _zz_867 = (left_bit_count_26 + _zz_869);
  assign _zz_868 = ((all_zeros_51 & _zz_870) & non_zeros_lzc_24);
  assign _zz_869 = {1'd0, _zz_868};
  assign _zz_870 = (whole_bit_count_27 + (~ all_zeros_51));
  assign _zz_871 = (left_bit_count_31 + _zz_873);
  assign _zz_872 = _zz_99[0];
  assign _zz_873 = {1'd0, _zz_872};
  assign _zz_874 = _zz_101[0];
  assign _zz_875 = {1'd0, _zz_874};
  assign _zz_876 = (left_bit_count_30 + _zz_878);
  assign _zz_877 = ((all_zeros_59 & _zz_879) & non_zeros_lzc_25);
  assign _zz_878 = {1'd0, _zz_877};
  assign _zz_879 = (whole_bit_count_31 + (~ all_zeros_59));
  assign _zz_880 = (left_bit_count_32 + _zz_882);
  assign _zz_881 = _zz_104[0];
  assign _zz_882 = {1'd0, _zz_881};
  assign _zz_883 = _zz_106[0];
  assign _zz_884 = {1'd0, _zz_883};
  assign _zz_885 = ((all_zeros_62 & _zz_887) & non_zeros_lzc_26);
  assign _zz_886 = {1'd0, _zz_885};
  assign _zz_887 = (whole_bit_count_32 + (~ all_zeros_62));
  assign _zz_888 = ((all_zeros_58 & _zz_890) & non_zeros_lzc_27);
  assign _zz_889 = {1'd0, _zz_888};
  assign _zz_890 = (whole_bit_count_30 + (~ all_zeros_58));
  assign _zz_891 = ((all_zeros_50 & _zz_893) & non_zeros_lzc_28);
  assign _zz_892 = {1'd0, _zz_891};
  assign _zz_893 = (whole_bit_count_26 + (~ all_zeros_50));
  assign _zz_894 = ((all_zeros_34 & _zz_896) & non_zeros_lzc_29);
  assign _zz_895 = {1'd0, _zz_894};
  assign _zz_896 = (whole_bit_count_18 + (~ all_zeros_34));
  assign _zz_897 = (left_bit_count_1 + _zz_899);
  assign _zz_898 = ((all_zeros_2 & _zz_900) & non_zeros_lzc_30);
  assign _zz_899 = {1'd0, _zz_898};
  assign _zz_900 = (whole_bit_count_2 + (~ all_zeros_2));
  assign _zz_901 = (left_bit_count_37 + _zz_903);
  assign _zz_902 = _zz_113[0];
  assign _zz_903 = {1'd0, _zz_902};
  assign _zz_904 = _zz_115[0];
  assign _zz_905 = {1'd0, _zz_904};
  assign _zz_906 = (left_bit_count_36 + _zz_908);
  assign _zz_907 = ((all_zeros_69 & _zz_909) & non_zeros_lzc_31);
  assign _zz_908 = {1'd0, _zz_907};
  assign _zz_909 = (whole_bit_count_37 + (~ all_zeros_69));
  assign _zz_910 = (left_bit_count_38 + _zz_912);
  assign _zz_911 = _zz_118[0];
  assign _zz_912 = {1'd0, _zz_911};
  assign _zz_913 = _zz_120[0];
  assign _zz_914 = {1'd0, _zz_913};
  assign _zz_915 = ((all_zeros_72 & _zz_917) & non_zeros_lzc_32);
  assign _zz_916 = {1'd0, _zz_915};
  assign _zz_917 = (whole_bit_count_38 + (~ all_zeros_72));
  assign _zz_918 = (left_bit_count_35 + _zz_920);
  assign _zz_919 = ((all_zeros_68 & _zz_921) & non_zeros_lzc_33);
  assign _zz_920 = {1'd0, _zz_919};
  assign _zz_921 = (whole_bit_count_36 + (~ all_zeros_68));
  assign _zz_922 = (left_bit_count_40 + _zz_924);
  assign _zz_923 = _zz_124[0];
  assign _zz_924 = {1'd0, _zz_923};
  assign _zz_925 = _zz_126[0];
  assign _zz_926 = {1'd0, _zz_925};
  assign _zz_927 = (left_bit_count_39 + _zz_929);
  assign _zz_928 = ((all_zeros_76 & _zz_930) & non_zeros_lzc_34);
  assign _zz_929 = {1'd0, _zz_928};
  assign _zz_930 = (whole_bit_count_40 + (~ all_zeros_76));
  assign _zz_931 = (left_bit_count_41 + _zz_933);
  assign _zz_932 = _zz_129[0];
  assign _zz_933 = {1'd0, _zz_932};
  assign _zz_934 = _zz_131[0];
  assign _zz_935 = {1'd0, _zz_934};
  assign _zz_936 = ((all_zeros_79 & _zz_938) & non_zeros_lzc_35);
  assign _zz_937 = {1'd0, _zz_936};
  assign _zz_938 = (whole_bit_count_41 + (~ all_zeros_79));
  assign _zz_939 = ((all_zeros_75 & _zz_941) & non_zeros_lzc_36);
  assign _zz_940 = {1'd0, _zz_939};
  assign _zz_941 = (whole_bit_count_39 + (~ all_zeros_75));
  assign _zz_942 = (left_bit_count_34 + _zz_944);
  assign _zz_943 = ((all_zeros_67 & _zz_945) & non_zeros_lzc_37);
  assign _zz_944 = {1'd0, _zz_943};
  assign _zz_945 = (whole_bit_count_35 + (~ all_zeros_67));
  assign _zz_946 = (left_bit_count_44 + _zz_948);
  assign _zz_947 = _zz_136[0];
  assign _zz_948 = {1'd0, _zz_947};
  assign _zz_949 = _zz_138[0];
  assign _zz_950 = {1'd0, _zz_949};
  assign _zz_951 = (left_bit_count_43 + _zz_953);
  assign _zz_952 = ((all_zeros_84 & _zz_954) & non_zeros_lzc_38);
  assign _zz_953 = {1'd0, _zz_952};
  assign _zz_954 = (whole_bit_count_44 + (~ all_zeros_84));
  assign _zz_955 = (left_bit_count_45 + _zz_957);
  assign _zz_956 = _zz_141[0];
  assign _zz_957 = {1'd0, _zz_956};
  assign _zz_958 = _zz_143[0];
  assign _zz_959 = {1'd0, _zz_958};
  assign _zz_960 = ((all_zeros_87 & _zz_962) & non_zeros_lzc_39);
  assign _zz_961 = {1'd0, _zz_960};
  assign _zz_962 = (whole_bit_count_45 + (~ all_zeros_87));
  assign _zz_963 = (left_bit_count_42 + _zz_965);
  assign _zz_964 = ((all_zeros_83 & _zz_966) & non_zeros_lzc_40);
  assign _zz_965 = {1'd0, _zz_964};
  assign _zz_966 = (whole_bit_count_43 + (~ all_zeros_83));
  assign _zz_967 = (left_bit_count_47 + _zz_969);
  assign _zz_968 = _zz_147[0];
  assign _zz_969 = {1'd0, _zz_968};
  assign _zz_970 = _zz_149[0];
  assign _zz_971 = {1'd0, _zz_970};
  assign _zz_972 = (left_bit_count_46 + _zz_974);
  assign _zz_973 = ((all_zeros_91 & _zz_975) & non_zeros_lzc_41);
  assign _zz_974 = {1'd0, _zz_973};
  assign _zz_975 = (whole_bit_count_47 + (~ all_zeros_91));
  assign _zz_976 = (left_bit_count_48 + _zz_978);
  assign _zz_977 = _zz_152[0];
  assign _zz_978 = {1'd0, _zz_977};
  assign _zz_979 = _zz_154[0];
  assign _zz_980 = {1'd0, _zz_979};
  assign _zz_981 = ((all_zeros_94 & _zz_983) & non_zeros_lzc_42);
  assign _zz_982 = {1'd0, _zz_981};
  assign _zz_983 = (whole_bit_count_48 + (~ all_zeros_94));
  assign _zz_984 = ((all_zeros_90 & _zz_986) & non_zeros_lzc_43);
  assign _zz_985 = {1'd0, _zz_984};
  assign _zz_986 = (whole_bit_count_46 + (~ all_zeros_90));
  assign _zz_987 = ((all_zeros_82 & _zz_989) & non_zeros_lzc_44);
  assign _zz_988 = {1'd0, _zz_987};
  assign _zz_989 = (whole_bit_count_42 + (~ all_zeros_82));
  assign _zz_990 = (left_bit_count_33 + _zz_992);
  assign _zz_991 = ((all_zeros_66 & _zz_993) & non_zeros_lzc_45);
  assign _zz_992 = {1'd0, _zz_991};
  assign _zz_993 = (whole_bit_count_34 + (~ all_zeros_66));
  assign _zz_994 = (left_bit_count_52 + _zz_996);
  assign _zz_995 = _zz_160[0];
  assign _zz_996 = {1'd0, _zz_995};
  assign _zz_997 = _zz_162[0];
  assign _zz_998 = {1'd0, _zz_997};
  assign _zz_999 = (left_bit_count_51 + _zz_1001);
  assign _zz_1000 = ((all_zeros_100 & _zz_1002) & non_zeros_lzc_46);
  assign _zz_1001 = {1'd0, _zz_1000};
  assign _zz_1002 = (whole_bit_count_52 + (~ all_zeros_100));
  assign _zz_1003 = (left_bit_count_53 + _zz_1005);
  assign _zz_1004 = _zz_165[0];
  assign _zz_1005 = {1'd0, _zz_1004};
  assign _zz_1006 = _zz_167[0];
  assign _zz_1007 = {1'd0, _zz_1006};
  assign _zz_1008 = ((all_zeros_103 & _zz_1010) & non_zeros_lzc_47);
  assign _zz_1009 = {1'd0, _zz_1008};
  assign _zz_1010 = (whole_bit_count_53 + (~ all_zeros_103));
  assign _zz_1011 = (left_bit_count_50 + _zz_1013);
  assign _zz_1012 = ((all_zeros_99 & _zz_1014) & non_zeros_lzc_48);
  assign _zz_1013 = {1'd0, _zz_1012};
  assign _zz_1014 = (whole_bit_count_51 + (~ all_zeros_99));
  assign _zz_1015 = (left_bit_count_55 + _zz_1017);
  assign _zz_1016 = _zz_171[0];
  assign _zz_1017 = {1'd0, _zz_1016};
  assign _zz_1018 = _zz_173[0];
  assign _zz_1019 = {1'd0, _zz_1018};
  assign _zz_1020 = (left_bit_count_54 + _zz_1022);
  assign _zz_1021 = ((all_zeros_107 & _zz_1023) & non_zeros_lzc_49);
  assign _zz_1022 = {1'd0, _zz_1021};
  assign _zz_1023 = (whole_bit_count_55 + (~ all_zeros_107));
  assign _zz_1024 = (left_bit_count_56 + _zz_1026);
  assign _zz_1025 = _zz_176[0];
  assign _zz_1026 = {1'd0, _zz_1025};
  assign _zz_1027 = _zz_178[0];
  assign _zz_1028 = {1'd0, _zz_1027};
  assign _zz_1029 = ((all_zeros_110 & _zz_1031) & non_zeros_lzc_50);
  assign _zz_1030 = {1'd0, _zz_1029};
  assign _zz_1031 = (whole_bit_count_56 + (~ all_zeros_110));
  assign _zz_1032 = ((all_zeros_106 & _zz_1034) & non_zeros_lzc_51);
  assign _zz_1033 = {1'd0, _zz_1032};
  assign _zz_1034 = (whole_bit_count_54 + (~ all_zeros_106));
  assign _zz_1035 = (left_bit_count_49 + _zz_1037);
  assign _zz_1036 = ((all_zeros_98 & _zz_1038) & non_zeros_lzc_52);
  assign _zz_1037 = {1'd0, _zz_1036};
  assign _zz_1038 = (whole_bit_count_50 + (~ all_zeros_98));
  assign _zz_1039 = (left_bit_count_59 + _zz_1041);
  assign _zz_1040 = _zz_183[0];
  assign _zz_1041 = {1'd0, _zz_1040};
  assign _zz_1042 = _zz_185[0];
  assign _zz_1043 = {1'd0, _zz_1042};
  assign _zz_1044 = (left_bit_count_58 + _zz_1046);
  assign _zz_1045 = ((all_zeros_115 & _zz_1047) & non_zeros_lzc_53);
  assign _zz_1046 = {1'd0, _zz_1045};
  assign _zz_1047 = (whole_bit_count_59 + (~ all_zeros_115));
  assign _zz_1048 = (left_bit_count_60 + _zz_1050);
  assign _zz_1049 = _zz_188[0];
  assign _zz_1050 = {1'd0, _zz_1049};
  assign _zz_1051 = _zz_190[0];
  assign _zz_1052 = {1'd0, _zz_1051};
  assign _zz_1053 = ((all_zeros_118 & _zz_1055) & non_zeros_lzc_54);
  assign _zz_1054 = {1'd0, _zz_1053};
  assign _zz_1055 = (whole_bit_count_60 + (~ all_zeros_118));
  assign _zz_1056 = (left_bit_count_57 + _zz_1058);
  assign _zz_1057 = ((all_zeros_114 & _zz_1059) & non_zeros_lzc_55);
  assign _zz_1058 = {1'd0, _zz_1057};
  assign _zz_1059 = (whole_bit_count_58 + (~ all_zeros_114));
  assign _zz_1060 = (left_bit_count_62 + _zz_1062);
  assign _zz_1061 = _zz_194[0];
  assign _zz_1062 = {1'd0, _zz_1061};
  assign _zz_1063 = _zz_196[0];
  assign _zz_1064 = {1'd0, _zz_1063};
  assign _zz_1065 = (left_bit_count_61 + _zz_1067);
  assign _zz_1066 = ((all_zeros_122 & _zz_1068) & non_zeros_lzc_56);
  assign _zz_1067 = {1'd0, _zz_1066};
  assign _zz_1068 = (whole_bit_count_62 + (~ all_zeros_122));
  assign _zz_1069 = (left_bit_count_63 + _zz_1071);
  assign _zz_1070 = _zz_199[0];
  assign _zz_1071 = {1'd0, _zz_1070};
  assign _zz_1072 = _zz_201[0];
  assign _zz_1073 = {1'd0, _zz_1072};
  assign _zz_1074 = ((all_zeros_125 & _zz_1076) & non_zeros_lzc_57);
  assign _zz_1075 = {1'd0, _zz_1074};
  assign _zz_1076 = (whole_bit_count_63 + (~ all_zeros_125));
  assign _zz_1077 = ((all_zeros_121 & _zz_1079) & non_zeros_lzc_58);
  assign _zz_1078 = {1'd0, _zz_1077};
  assign _zz_1079 = (whole_bit_count_61 + (~ all_zeros_121));
  assign _zz_1080 = ((all_zeros_113 & _zz_1082) & non_zeros_lzc_59);
  assign _zz_1081 = {1'd0, _zz_1080};
  assign _zz_1082 = (whole_bit_count_57 + (~ all_zeros_113));
  assign _zz_1083 = ((all_zeros_97 & _zz_1085) & non_zeros_lzc_60);
  assign _zz_1084 = {1'd0, _zz_1083};
  assign _zz_1085 = (whole_bit_count_49 + (~ all_zeros_97));
  assign _zz_1086 = ((all_zeros_65 & _zz_1088) & non_zeros_lzc_61);
  assign _zz_1087 = {1'd0, _zz_1086};
  assign _zz_1088 = (whole_bit_count_33 + (~ all_zeros_65));
  assign _zz_1089 = (left_bit_count + _zz_1091);
  assign _zz_1090 = ((all_zeros_1 & _zz_1092) & non_zeros_lzc_62);
  assign _zz_1091 = {1'd0, _zz_1090};
  assign _zz_1092 = (whole_bit_count_1 + (~ all_zeros_1));
  assign _zz_1093 = (left_bit_count_69 + _zz_1095);
  assign _zz_1094 = _zz_209[0];
  assign _zz_1095 = {1'd0, _zz_1094};
  assign _zz_1096 = _zz_211[0];
  assign _zz_1097 = {1'd0, _zz_1096};
  assign _zz_1098 = (left_bit_count_68 + _zz_1100);
  assign _zz_1099 = ((all_zeros_133 & _zz_1101) & non_zeros_lzc_63);
  assign _zz_1100 = {1'd0, _zz_1099};
  assign _zz_1101 = (whole_bit_count_69 + (~ all_zeros_133));
  assign _zz_1102 = (left_bit_count_70 + _zz_1104);
  assign _zz_1103 = _zz_214[0];
  assign _zz_1104 = {1'd0, _zz_1103};
  assign _zz_1105 = _zz_216[0];
  assign _zz_1106 = {1'd0, _zz_1105};
  assign _zz_1107 = ((all_zeros_136 & _zz_1109) & non_zeros_lzc_64);
  assign _zz_1108 = {1'd0, _zz_1107};
  assign _zz_1109 = (whole_bit_count_70 + (~ all_zeros_136));
  assign _zz_1110 = (left_bit_count_67 + _zz_1112);
  assign _zz_1111 = ((all_zeros_132 & _zz_1113) & non_zeros_lzc_65);
  assign _zz_1112 = {1'd0, _zz_1111};
  assign _zz_1113 = (whole_bit_count_68 + (~ all_zeros_132));
  assign _zz_1114 = (left_bit_count_72 + _zz_1116);
  assign _zz_1115 = _zz_220[0];
  assign _zz_1116 = {1'd0, _zz_1115};
  assign _zz_1117 = _zz_222[0];
  assign _zz_1118 = {1'd0, _zz_1117};
  assign _zz_1119 = (left_bit_count_71 + _zz_1121);
  assign _zz_1120 = ((all_zeros_140 & _zz_1122) & non_zeros_lzc_66);
  assign _zz_1121 = {1'd0, _zz_1120};
  assign _zz_1122 = (whole_bit_count_72 + (~ all_zeros_140));
  assign _zz_1123 = (left_bit_count_73 + _zz_1125);
  assign _zz_1124 = _zz_225[0];
  assign _zz_1125 = {1'd0, _zz_1124};
  assign _zz_1126 = _zz_227[0];
  assign _zz_1127 = {1'd0, _zz_1126};
  assign _zz_1128 = ((all_zeros_143 & _zz_1130) & non_zeros_lzc_67);
  assign _zz_1129 = {1'd0, _zz_1128};
  assign _zz_1130 = (whole_bit_count_73 + (~ all_zeros_143));
  assign _zz_1131 = ((all_zeros_139 & _zz_1133) & non_zeros_lzc_68);
  assign _zz_1132 = {1'd0, _zz_1131};
  assign _zz_1133 = (whole_bit_count_71 + (~ all_zeros_139));
  assign _zz_1134 = (left_bit_count_66 + _zz_1136);
  assign _zz_1135 = ((all_zeros_131 & _zz_1137) & non_zeros_lzc_69);
  assign _zz_1136 = {1'd0, _zz_1135};
  assign _zz_1137 = (whole_bit_count_67 + (~ all_zeros_131));
  assign _zz_1138 = (left_bit_count_76 + _zz_1140);
  assign _zz_1139 = _zz_232[0];
  assign _zz_1140 = {1'd0, _zz_1139};
  assign _zz_1141 = _zz_234[0];
  assign _zz_1142 = {1'd0, _zz_1141};
  assign _zz_1143 = (left_bit_count_75 + _zz_1145);
  assign _zz_1144 = ((all_zeros_148 & _zz_1146) & non_zeros_lzc_70);
  assign _zz_1145 = {1'd0, _zz_1144};
  assign _zz_1146 = (whole_bit_count_76 + (~ all_zeros_148));
  assign _zz_1147 = (left_bit_count_77 + _zz_1149);
  assign _zz_1148 = _zz_237[0];
  assign _zz_1149 = {1'd0, _zz_1148};
  assign _zz_1150 = _zz_239[0];
  assign _zz_1151 = {1'd0, _zz_1150};
  assign _zz_1152 = ((all_zeros_151 & _zz_1154) & non_zeros_lzc_71);
  assign _zz_1153 = {1'd0, _zz_1152};
  assign _zz_1154 = (whole_bit_count_77 + (~ all_zeros_151));
  assign _zz_1155 = (left_bit_count_74 + _zz_1157);
  assign _zz_1156 = ((all_zeros_147 & _zz_1158) & non_zeros_lzc_72);
  assign _zz_1157 = {1'd0, _zz_1156};
  assign _zz_1158 = (whole_bit_count_75 + (~ all_zeros_147));
  assign _zz_1159 = (left_bit_count_79 + _zz_1161);
  assign _zz_1160 = _zz_243[0];
  assign _zz_1161 = {1'd0, _zz_1160};
  assign _zz_1162 = _zz_245[0];
  assign _zz_1163 = {1'd0, _zz_1162};
  assign _zz_1164 = (left_bit_count_78 + _zz_1166);
  assign _zz_1165 = ((all_zeros_155 & _zz_1167) & non_zeros_lzc_73);
  assign _zz_1166 = {1'd0, _zz_1165};
  assign _zz_1167 = (whole_bit_count_79 + (~ all_zeros_155));
  assign _zz_1168 = (left_bit_count_80 + _zz_1170);
  assign _zz_1169 = _zz_248[0];
  assign _zz_1170 = {1'd0, _zz_1169};
  assign _zz_1171 = _zz_250[0];
  assign _zz_1172 = {1'd0, _zz_1171};
  assign _zz_1173 = ((all_zeros_158 & _zz_1175) & non_zeros_lzc_74);
  assign _zz_1174 = {1'd0, _zz_1173};
  assign _zz_1175 = (whole_bit_count_80 + (~ all_zeros_158));
  assign _zz_1176 = ((all_zeros_154 & _zz_1178) & non_zeros_lzc_75);
  assign _zz_1177 = {1'd0, _zz_1176};
  assign _zz_1178 = (whole_bit_count_78 + (~ all_zeros_154));
  assign _zz_1179 = ((all_zeros_146 & _zz_1181) & non_zeros_lzc_76);
  assign _zz_1180 = {1'd0, _zz_1179};
  assign _zz_1181 = (whole_bit_count_74 + (~ all_zeros_146));
  assign _zz_1182 = (left_bit_count_65 + _zz_1184);
  assign _zz_1183 = ((all_zeros_130 & _zz_1185) & non_zeros_lzc_77);
  assign _zz_1184 = {1'd0, _zz_1183};
  assign _zz_1185 = (whole_bit_count_66 + (~ all_zeros_130));
  assign _zz_1186 = (left_bit_count_84 + _zz_1188);
  assign _zz_1187 = _zz_256[0];
  assign _zz_1188 = {1'd0, _zz_1187};
  assign _zz_1189 = _zz_258[0];
  assign _zz_1190 = {1'd0, _zz_1189};
  assign _zz_1191 = (left_bit_count_83 + _zz_1193);
  assign _zz_1192 = ((all_zeros_164 & _zz_1194) & non_zeros_lzc_78);
  assign _zz_1193 = {1'd0, _zz_1192};
  assign _zz_1194 = (whole_bit_count_84 + (~ all_zeros_164));
  assign _zz_1195 = (left_bit_count_85 + _zz_1197);
  assign _zz_1196 = _zz_261[0];
  assign _zz_1197 = {1'd0, _zz_1196};
  assign _zz_1198 = _zz_263[0];
  assign _zz_1199 = {1'd0, _zz_1198};
  assign _zz_1200 = ((all_zeros_167 & _zz_1202) & non_zeros_lzc_79);
  assign _zz_1201 = {1'd0, _zz_1200};
  assign _zz_1202 = (whole_bit_count_85 + (~ all_zeros_167));
  assign _zz_1203 = (left_bit_count_82 + _zz_1205);
  assign _zz_1204 = ((all_zeros_163 & _zz_1206) & non_zeros_lzc_80);
  assign _zz_1205 = {1'd0, _zz_1204};
  assign _zz_1206 = (whole_bit_count_83 + (~ all_zeros_163));
  assign _zz_1207 = (left_bit_count_87 + _zz_1209);
  assign _zz_1208 = _zz_267[0];
  assign _zz_1209 = {1'd0, _zz_1208};
  assign _zz_1210 = _zz_269[0];
  assign _zz_1211 = {1'd0, _zz_1210};
  assign _zz_1212 = (left_bit_count_86 + _zz_1214);
  assign _zz_1213 = ((all_zeros_171 & _zz_1215) & non_zeros_lzc_81);
  assign _zz_1214 = {1'd0, _zz_1213};
  assign _zz_1215 = (whole_bit_count_87 + (~ all_zeros_171));
  assign _zz_1216 = (left_bit_count_88 + _zz_1218);
  assign _zz_1217 = _zz_272[0];
  assign _zz_1218 = {1'd0, _zz_1217};
  assign _zz_1219 = _zz_274[0];
  assign _zz_1220 = {1'd0, _zz_1219};
  assign _zz_1221 = ((all_zeros_174 & _zz_1223) & non_zeros_lzc_82);
  assign _zz_1222 = {1'd0, _zz_1221};
  assign _zz_1223 = (whole_bit_count_88 + (~ all_zeros_174));
  assign _zz_1224 = ((all_zeros_170 & _zz_1226) & non_zeros_lzc_83);
  assign _zz_1225 = {1'd0, _zz_1224};
  assign _zz_1226 = (whole_bit_count_86 + (~ all_zeros_170));
  assign _zz_1227 = (left_bit_count_81 + _zz_1229);
  assign _zz_1228 = ((all_zeros_162 & _zz_1230) & non_zeros_lzc_84);
  assign _zz_1229 = {1'd0, _zz_1228};
  assign _zz_1230 = (whole_bit_count_82 + (~ all_zeros_162));
  assign _zz_1231 = (left_bit_count_91 + _zz_1233);
  assign _zz_1232 = _zz_279[0];
  assign _zz_1233 = {1'd0, _zz_1232};
  assign _zz_1234 = _zz_281[0];
  assign _zz_1235 = {1'd0, _zz_1234};
  assign _zz_1236 = (left_bit_count_90 + _zz_1238);
  assign _zz_1237 = ((all_zeros_179 & _zz_1239) & non_zeros_lzc_85);
  assign _zz_1238 = {1'd0, _zz_1237};
  assign _zz_1239 = (whole_bit_count_91 + (~ all_zeros_179));
  assign _zz_1240 = (left_bit_count_92 + _zz_1242);
  assign _zz_1241 = _zz_284[0];
  assign _zz_1242 = {1'd0, _zz_1241};
  assign _zz_1243 = _zz_286[0];
  assign _zz_1244 = {1'd0, _zz_1243};
  assign _zz_1245 = ((all_zeros_182 & _zz_1247) & non_zeros_lzc_86);
  assign _zz_1246 = {1'd0, _zz_1245};
  assign _zz_1247 = (whole_bit_count_92 + (~ all_zeros_182));
  assign _zz_1248 = (left_bit_count_89 + _zz_1250);
  assign _zz_1249 = ((all_zeros_178 & _zz_1251) & non_zeros_lzc_87);
  assign _zz_1250 = {1'd0, _zz_1249};
  assign _zz_1251 = (whole_bit_count_90 + (~ all_zeros_178));
  assign _zz_1252 = (left_bit_count_94 + _zz_1254);
  assign _zz_1253 = _zz_290[0];
  assign _zz_1254 = {1'd0, _zz_1253};
  assign _zz_1255 = _zz_292[0];
  assign _zz_1256 = {1'd0, _zz_1255};
  assign _zz_1257 = (left_bit_count_93 + _zz_1259);
  assign _zz_1258 = ((all_zeros_186 & _zz_1260) & non_zeros_lzc_88);
  assign _zz_1259 = {1'd0, _zz_1258};
  assign _zz_1260 = (whole_bit_count_94 + (~ all_zeros_186));
  assign _zz_1261 = (left_bit_count_95 + _zz_1263);
  assign _zz_1262 = _zz_295[0];
  assign _zz_1263 = {1'd0, _zz_1262};
  assign _zz_1264 = _zz_297[0];
  assign _zz_1265 = {1'd0, _zz_1264};
  assign _zz_1266 = ((all_zeros_189 & _zz_1268) & non_zeros_lzc_89);
  assign _zz_1267 = {1'd0, _zz_1266};
  assign _zz_1268 = (whole_bit_count_95 + (~ all_zeros_189));
  assign _zz_1269 = ((all_zeros_185 & _zz_1271) & non_zeros_lzc_90);
  assign _zz_1270 = {1'd0, _zz_1269};
  assign _zz_1271 = (whole_bit_count_93 + (~ all_zeros_185));
  assign _zz_1272 = ((all_zeros_177 & _zz_1274) & non_zeros_lzc_91);
  assign _zz_1273 = {1'd0, _zz_1272};
  assign _zz_1274 = (whole_bit_count_89 + (~ all_zeros_177));
  assign _zz_1275 = ((all_zeros_161 & _zz_1277) & non_zeros_lzc_92);
  assign _zz_1276 = {1'd0, _zz_1275};
  assign _zz_1277 = (whole_bit_count_81 + (~ all_zeros_161));
  assign _zz_1278 = (left_bit_count_64 + _zz_1280);
  assign _zz_1279 = ((all_zeros_129 & _zz_1281) & non_zeros_lzc_93);
  assign _zz_1280 = {1'd0, _zz_1279};
  assign _zz_1281 = (whole_bit_count_65 + (~ all_zeros_129));
  assign _zz_1282 = (left_bit_count_100 + _zz_1284);
  assign _zz_1283 = _zz_304[0];
  assign _zz_1284 = {1'd0, _zz_1283};
  assign _zz_1285 = _zz_306[0];
  assign _zz_1286 = {1'd0, _zz_1285};
  assign _zz_1287 = (left_bit_count_99 + _zz_1289);
  assign _zz_1288 = ((all_zeros_196 & _zz_1290) & non_zeros_lzc_94);
  assign _zz_1289 = {1'd0, _zz_1288};
  assign _zz_1290 = (whole_bit_count_100 + (~ all_zeros_196));
  assign _zz_1291 = (left_bit_count_101 + _zz_1293);
  assign _zz_1292 = _zz_309[0];
  assign _zz_1293 = {1'd0, _zz_1292};
  assign _zz_1294 = _zz_311[0];
  assign _zz_1295 = {1'd0, _zz_1294};
  assign _zz_1296 = ((all_zeros_199 & _zz_1298) & non_zeros_lzc_95);
  assign _zz_1297 = {1'd0, _zz_1296};
  assign _zz_1298 = (whole_bit_count_101 + (~ all_zeros_199));
  assign _zz_1299 = (left_bit_count_98 + _zz_1301);
  assign _zz_1300 = ((all_zeros_195 & _zz_1302) & non_zeros_lzc_96);
  assign _zz_1301 = {1'd0, _zz_1300};
  assign _zz_1302 = (whole_bit_count_99 + (~ all_zeros_195));
  assign _zz_1303 = (left_bit_count_103 + _zz_1305);
  assign _zz_1304 = _zz_315[0];
  assign _zz_1305 = {1'd0, _zz_1304};
  assign _zz_1306 = _zz_317[0];
  assign _zz_1307 = {1'd0, _zz_1306};
  assign _zz_1308 = (left_bit_count_102 + _zz_1310);
  assign _zz_1309 = ((all_zeros_203 & _zz_1311) & non_zeros_lzc_97);
  assign _zz_1310 = {1'd0, _zz_1309};
  assign _zz_1311 = (whole_bit_count_103 + (~ all_zeros_203));
  assign _zz_1312 = (left_bit_count_104 + _zz_1314);
  assign _zz_1313 = _zz_320[0];
  assign _zz_1314 = {1'd0, _zz_1313};
  assign _zz_1315 = _zz_322[0];
  assign _zz_1316 = {1'd0, _zz_1315};
  assign _zz_1317 = ((all_zeros_206 & _zz_1319) & non_zeros_lzc_98);
  assign _zz_1318 = {1'd0, _zz_1317};
  assign _zz_1319 = (whole_bit_count_104 + (~ all_zeros_206));
  assign _zz_1320 = ((all_zeros_202 & _zz_1322) & non_zeros_lzc_99);
  assign _zz_1321 = {1'd0, _zz_1320};
  assign _zz_1322 = (whole_bit_count_102 + (~ all_zeros_202));
  assign _zz_1323 = (left_bit_count_97 + _zz_1325);
  assign _zz_1324 = ((all_zeros_194 & _zz_1326) & non_zeros_lzc_100);
  assign _zz_1325 = {1'd0, _zz_1324};
  assign _zz_1326 = (whole_bit_count_98 + (~ all_zeros_194));
  assign _zz_1327 = (left_bit_count_107 + _zz_1329);
  assign _zz_1328 = _zz_327[0];
  assign _zz_1329 = {1'd0, _zz_1328};
  assign _zz_1330 = _zz_329[0];
  assign _zz_1331 = {1'd0, _zz_1330};
  assign _zz_1332 = (left_bit_count_106 + _zz_1334);
  assign _zz_1333 = ((all_zeros_211 & _zz_1335) & non_zeros_lzc_101);
  assign _zz_1334 = {1'd0, _zz_1333};
  assign _zz_1335 = (whole_bit_count_107 + (~ all_zeros_211));
  assign _zz_1336 = (left_bit_count_108 + _zz_1338);
  assign _zz_1337 = _zz_332[0];
  assign _zz_1338 = {1'd0, _zz_1337};
  assign _zz_1339 = _zz_334[0];
  assign _zz_1340 = {1'd0, _zz_1339};
  assign _zz_1341 = ((all_zeros_214 & _zz_1343) & non_zeros_lzc_102);
  assign _zz_1342 = {1'd0, _zz_1341};
  assign _zz_1343 = (whole_bit_count_108 + (~ all_zeros_214));
  assign _zz_1344 = (left_bit_count_105 + _zz_1346);
  assign _zz_1345 = ((all_zeros_210 & _zz_1347) & non_zeros_lzc_103);
  assign _zz_1346 = {1'd0, _zz_1345};
  assign _zz_1347 = (whole_bit_count_106 + (~ all_zeros_210));
  assign _zz_1348 = (left_bit_count_110 + _zz_1350);
  assign _zz_1349 = _zz_338[0];
  assign _zz_1350 = {1'd0, _zz_1349};
  assign _zz_1351 = _zz_340[0];
  assign _zz_1352 = {1'd0, _zz_1351};
  assign _zz_1353 = (left_bit_count_109 + _zz_1355);
  assign _zz_1354 = ((all_zeros_218 & _zz_1356) & non_zeros_lzc_104);
  assign _zz_1355 = {1'd0, _zz_1354};
  assign _zz_1356 = (whole_bit_count_110 + (~ all_zeros_218));
  assign _zz_1357 = (left_bit_count_111 + _zz_1359);
  assign _zz_1358 = _zz_343[0];
  assign _zz_1359 = {1'd0, _zz_1358};
  assign _zz_1360 = _zz_345[0];
  assign _zz_1361 = {1'd0, _zz_1360};
  assign _zz_1362 = ((all_zeros_221 & _zz_1364) & non_zeros_lzc_105);
  assign _zz_1363 = {1'd0, _zz_1362};
  assign _zz_1364 = (whole_bit_count_111 + (~ all_zeros_221));
  assign _zz_1365 = ((all_zeros_217 & _zz_1367) & non_zeros_lzc_106);
  assign _zz_1366 = {1'd0, _zz_1365};
  assign _zz_1367 = (whole_bit_count_109 + (~ all_zeros_217));
  assign _zz_1368 = ((all_zeros_209 & _zz_1370) & non_zeros_lzc_107);
  assign _zz_1369 = {1'd0, _zz_1368};
  assign _zz_1370 = (whole_bit_count_105 + (~ all_zeros_209));
  assign _zz_1371 = (left_bit_count_96 + _zz_1373);
  assign _zz_1372 = ((all_zeros_193 & _zz_1374) & non_zeros_lzc_108);
  assign _zz_1373 = {1'd0, _zz_1372};
  assign _zz_1374 = (whole_bit_count_97 + (~ all_zeros_193));
  assign _zz_1375 = (left_bit_count_115 + _zz_1377);
  assign _zz_1376 = _zz_351[0];
  assign _zz_1377 = {1'd0, _zz_1376};
  assign _zz_1378 = _zz_353[0];
  assign _zz_1379 = {1'd0, _zz_1378};
  assign _zz_1380 = (left_bit_count_114 + _zz_1382);
  assign _zz_1381 = ((all_zeros_227 & _zz_1383) & non_zeros_lzc_109);
  assign _zz_1382 = {1'd0, _zz_1381};
  assign _zz_1383 = (whole_bit_count_115 + (~ all_zeros_227));
  assign _zz_1384 = (left_bit_count_116 + _zz_1386);
  assign _zz_1385 = _zz_356[0];
  assign _zz_1386 = {1'd0, _zz_1385};
  assign _zz_1387 = _zz_358[0];
  assign _zz_1388 = {1'd0, _zz_1387};
  assign _zz_1389 = ((all_zeros_230 & _zz_1391) & non_zeros_lzc_110);
  assign _zz_1390 = {1'd0, _zz_1389};
  assign _zz_1391 = (whole_bit_count_116 + (~ all_zeros_230));
  assign _zz_1392 = (left_bit_count_113 + _zz_1394);
  assign _zz_1393 = ((all_zeros_226 & _zz_1395) & non_zeros_lzc_111);
  assign _zz_1394 = {1'd0, _zz_1393};
  assign _zz_1395 = (whole_bit_count_114 + (~ all_zeros_226));
  assign _zz_1396 = (left_bit_count_118 + _zz_1398);
  assign _zz_1397 = _zz_362[0];
  assign _zz_1398 = {1'd0, _zz_1397};
  assign _zz_1399 = _zz_364[0];
  assign _zz_1400 = {1'd0, _zz_1399};
  assign _zz_1401 = (left_bit_count_117 + _zz_1403);
  assign _zz_1402 = ((all_zeros_234 & _zz_1404) & non_zeros_lzc_112);
  assign _zz_1403 = {1'd0, _zz_1402};
  assign _zz_1404 = (whole_bit_count_118 + (~ all_zeros_234));
  assign _zz_1405 = (left_bit_count_119 + _zz_1407);
  assign _zz_1406 = _zz_367[0];
  assign _zz_1407 = {1'd0, _zz_1406};
  assign _zz_1408 = _zz_369[0];
  assign _zz_1409 = {1'd0, _zz_1408};
  assign _zz_1410 = ((all_zeros_237 & _zz_1412) & non_zeros_lzc_113);
  assign _zz_1411 = {1'd0, _zz_1410};
  assign _zz_1412 = (whole_bit_count_119 + (~ all_zeros_237));
  assign _zz_1413 = ((all_zeros_233 & _zz_1415) & non_zeros_lzc_114);
  assign _zz_1414 = {1'd0, _zz_1413};
  assign _zz_1415 = (whole_bit_count_117 + (~ all_zeros_233));
  assign _zz_1416 = (left_bit_count_112 + _zz_1418);
  assign _zz_1417 = ((all_zeros_225 & _zz_1419) & non_zeros_lzc_115);
  assign _zz_1418 = {1'd0, _zz_1417};
  assign _zz_1419 = (whole_bit_count_113 + (~ all_zeros_225));
  assign _zz_1420 = (left_bit_count_122 + _zz_1422);
  assign _zz_1421 = _zz_374[0];
  assign _zz_1422 = {1'd0, _zz_1421};
  assign _zz_1423 = _zz_376[0];
  assign _zz_1424 = {1'd0, _zz_1423};
  assign _zz_1425 = (left_bit_count_121 + _zz_1427);
  assign _zz_1426 = ((all_zeros_242 & _zz_1428) & non_zeros_lzc_116);
  assign _zz_1427 = {1'd0, _zz_1426};
  assign _zz_1428 = (whole_bit_count_122 + (~ all_zeros_242));
  assign _zz_1429 = (left_bit_count_123 + _zz_1431);
  assign _zz_1430 = _zz_379[0];
  assign _zz_1431 = {1'd0, _zz_1430};
  assign _zz_1432 = _zz_381[0];
  assign _zz_1433 = {1'd0, _zz_1432};
  assign _zz_1434 = ((all_zeros_245 & _zz_1436) & non_zeros_lzc_117);
  assign _zz_1435 = {1'd0, _zz_1434};
  assign _zz_1436 = (whole_bit_count_123 + (~ all_zeros_245));
  assign _zz_1437 = (left_bit_count_120 + _zz_1439);
  assign _zz_1438 = ((all_zeros_241 & _zz_1440) & non_zeros_lzc_118);
  assign _zz_1439 = {1'd0, _zz_1438};
  assign _zz_1440 = (whole_bit_count_121 + (~ all_zeros_241));
  assign _zz_1441 = (left_bit_count_125 + _zz_1443);
  assign _zz_1442 = _zz_385[0];
  assign _zz_1443 = {1'd0, _zz_1442};
  assign _zz_1444 = _zz_387[0];
  assign _zz_1445 = {1'd0, _zz_1444};
  assign _zz_1446 = (left_bit_count_124 + _zz_1448);
  assign _zz_1447 = ((all_zeros_249 & _zz_1449) & non_zeros_lzc_119);
  assign _zz_1448 = {1'd0, _zz_1447};
  assign _zz_1449 = (whole_bit_count_125 + (~ all_zeros_249));
  assign _zz_1450 = (left_bit_count_126 + _zz_1452);
  assign _zz_1451 = _zz_390[0];
  assign _zz_1452 = {1'd0, _zz_1451};
  assign _zz_1453 = _zz_392[0];
  assign _zz_1454 = {1'd0, _zz_1453};
  assign _zz_1455 = ((all_zeros_252 & _zz_1457) & non_zeros_lzc_120);
  assign _zz_1456 = {1'd0, _zz_1455};
  assign _zz_1457 = (whole_bit_count_126 + (~ all_zeros_252));
  assign _zz_1458 = ((all_zeros_248 & _zz_1460) & non_zeros_lzc_121);
  assign _zz_1459 = {1'd0, _zz_1458};
  assign _zz_1460 = (whole_bit_count_124 + (~ all_zeros_248));
  assign _zz_1461 = ((all_zeros_240 & _zz_1463) & non_zeros_lzc_122);
  assign _zz_1462 = {1'd0, _zz_1461};
  assign _zz_1463 = (whole_bit_count_120 + (~ all_zeros_240));
  assign _zz_1464 = ((all_zeros_224 & _zz_1466) & non_zeros_lzc_123);
  assign _zz_1465 = {1'd0, _zz_1464};
  assign _zz_1466 = (whole_bit_count_112 + (~ all_zeros_224));
  assign _zz_1467 = ((all_zeros_192 & _zz_1469) & non_zeros_lzc_124);
  assign _zz_1468 = {1'd0, _zz_1467};
  assign _zz_1469 = (whole_bit_count_96 + (~ all_zeros_192));
  assign _zz_1470 = ((all_zeros_128 & _zz_1472) & non_zeros_lzc_125);
  assign _zz_1471 = {1'd0, _zz_1470};
  assign _zz_1472 = (whole_bit_count_64 + (~ all_zeros_128));
  assign _zz_1473 = (whole_bit_count + (~ all_zeros));
  assign _zz_1474 = {1'd0, lzc};
  assign _zz_1475 = _zz_447;
  assign _zz_1476 = _zz_1477[7 : 0];
  assign _zz_1477 = _zz_450;
  assign _zz_1478 = _zz_1479[7 : 0];
  assign _zz_1479 = fixTo_1_dout;
  assign _zz_1480 = divUnit_1_c[7 : 0];
  assign _zz_1481 = _zz_1482[7 : 0];
  assign _zz_1482 = fixTo_2_dout;
  assign _zz_1483 = divUnit_2_c[7 : 0];
  assign _zz_1484 = _zz_1485[15 : 0];
  assign _zz_1485 = fixTo_3_dout;
  assign _zz_1486 = _zz_1487[15 : 0];
  assign _zz_1487 = fixTo_4_dout;
  assign _zz_1488 = fixTo_5_dout;
  assign _zz_1489 = _zz_1490[15 : 0];
  assign _zz_1490 = fixTo_6_dout;
  assign _zz_1491 = _zz_1492[15 : 0];
  assign _zz_1492 = fixTo_7_dout;
  assign _zz_1493 = _zz_1494[15 : 0];
  assign _zz_1494 = fixTo_9_dout;
  assign _zz_1495 = _zz_1496[15 : 0];
  assign _zz_1496 = fixTo_10_dout;
  assign _zz_1497 = ({8'd0,_zz_1499} <<< 8);
  assign _zz_1498 = {{8{_zz_1497[23]}}, _zz_1497};
  assign _zz_1499 = ($signed(_zz_404) - $signed(_zz_1500));
  assign _zz_1500 = _zz_1501[15 : 0];
  assign _zz_1501 = fixTo_11_dout;
  assign _zz_1502 = ({8'd0,_zz_397} <<< 8);
  assign _zz_1503 = {{8{_zz_1502[23]}}, _zz_1502};
  assign _zz_1504 = ({8'd0,_zz_1506} <<< 8);
  assign _zz_1505 = {{8{_zz_1504[23]}}, _zz_1504};
  assign _zz_1506 = ($signed(_zz_404) + $signed(_zz_1507));
  assign _zz_1507 = _zz_1508[15 : 0];
  assign _zz_1508 = fixTo_8_dout;
  assign _zz_1509 = ({8'd0,_zz_398} <<< 8);
  assign _zz_1510 = {{8{_zz_1509[23]}}, _zz_1509};
  assign _zz_1511 = ({8'd0,func_table_0_regNext_real} <<< 8);
  assign _zz_1512 = ({8'd0,func_table_0_regNext_imag} <<< 8);
  assign _zz_1513 = ({8'd0,func_table_127_regNext_real} <<< 8);
  assign _zz_1514 = ({8'd0,func_table_127_regNext_imag} <<< 8);
  assign _zz_1515 = _zz_1516[15 : 0];
  assign _zz_1516 = fixTo_12_dout;
  assign _zz_1517 = _zz_1518[15 : 0];
  assign _zz_1518 = fixTo_13_dout;
  assign _zz_1519 = ({8'd0,_zz_1520} <<< 8);
  assign _zz_1520 = divUnit_3_c[15 : 0];
  assign _zz_1521 = ({8'd0,_zz_1522} <<< 8);
  assign _zz_1522 = divUnit_4_c[15 : 0];
  assign _zz_1523 = _zz_1524[31 : 0];
  assign _zz_1524 = fixTo_14_dout;
  assign _zz_1525 = _zz_1526[31 : 0];
  assign _zz_1526 = fixTo_15_dout;
  assign _zz_1527 = fixTo_16_dout;
  assign _zz_1528 = _zz_1529[31 : 0];
  assign _zz_1529 = fixTo_17_dout;
  assign _zz_1530 = _zz_1531[31 : 0];
  assign _zz_1531 = fixTo_18_dout;
  assign _zz_1532 = _zz_1533[31 : 0];
  assign _zz_1533 = fixTo_20_dout;
  assign _zz_1534 = _zz_1535[31 : 0];
  assign _zz_1535 = fixTo_21_dout;
  assign _zz_1536 = ({16'd0,_zz_1537} <<< 16);
  assign _zz_1537 = ($signed(_zz_410) - $signed(_zz_1538));
  assign _zz_1538 = _zz_1539[31 : 0];
  assign _zz_1539 = fixTo_22_dout;
  assign _zz_1540 = ({16'd0,_zz_1541} <<< 16);
  assign _zz_1541 = ($signed(_zz_410) + $signed(_zz_1542));
  assign _zz_1542 = _zz_1543[31 : 0];
  assign _zz_1543 = fixTo_19_dout;
  assign _zz_1544 = fixTo_23_dout;
  assign _zz_1545 = fixTo_24_dout;
  SInt32fixTo15_8_ROUNDTOINF fixTo (
    .din     (_zz_9[31:0]      ), //i
    .dout    (fixTo_dout[7:0]  )  //o
  );
  SInt16fixTo7_0_ROUNDTOINF fixTo_1 (
    .din     (_zz_413[15:0]      ), //i
    .dout    (fixTo_1_dout[7:0]  )  //o
  );
  SInt16fixTo7_0_ROUNDTOINF fixTo_2 (
    .din     (_zz_414[15:0]      ), //i
    .dout    (fixTo_2_dout[7:0]  )  //o
  );
  DivUnit divUnit_1 (
    .a    (_zz_415[7:0]      ), //i
    .b    (_zz_416[7:0]      ), //i
    .c    (divUnit_1_c[7:0]  )  //o
  );
  DivUnit divUnit_2 (
    .a    (_zz_417[7:0]      ), //i
    .b    (_zz_418[7:0]      ), //i
    .c    (divUnit_2_c[7:0]  )  //o
  );
  SInt16fixTo15_0_ROUNDTOINF fixTo_3 (
    .din     (_zz_419[15:0]       ), //i
    .dout    (fixTo_3_dout[15:0]  )  //o
  );
  SInt8fixTo15_0_ROUNDTOINF fixTo_4 (
    .din     (_zz_402[7:0]        ), //i
    .dout    (fixTo_4_dout[15:0]  )  //o
  );
  MulUnit mulUnit_1 (
    .a    (_zz_420[15:0]      ), //i
    .b    (_zz_421[15:0]      ), //i
    .c    (mulUnit_1_c[15:0]  )  //o
  );
  SInt16fixTo15_0_ROUNDTOINF fixTo_5 (
    .din     (_zz_422[15:0]       ), //i
    .dout    (fixTo_5_dout[15:0]  )  //o
  );
  SInt8fixTo15_0_ROUNDTOINF fixTo_6 (
    .din     (_zz_423[7:0]        ), //i
    .dout    (fixTo_6_dout[15:0]  )  //o
  );
  SInt16fixTo15_0_ROUNDTOINF fixTo_7 (
    .din     (_zz_400[15:0]       ), //i
    .dout    (fixTo_7_dout[15:0]  )  //o
  );
  MulUnit mulUnit_2 (
    .a    (_zz_424[15:0]      ), //i
    .b    (_zz_425[15:0]      ), //i
    .c    (mulUnit_2_c[15:0]  )  //o
  );
  SInt16fixTo15_0_ROUNDTOINF fixTo_8 (
    .din     (_zz_426[15:0]       ), //i
    .dout    (fixTo_8_dout[15:0]  )  //o
  );
  SInt8fixTo15_0_ROUNDTOINF fixTo_9 (
    .din     (_zz_427[7:0]        ), //i
    .dout    (fixTo_9_dout[15:0]  )  //o
  );
  SInt16fixTo15_0_ROUNDTOINF fixTo_10 (
    .din     (_zz_401[15:0]        ), //i
    .dout    (fixTo_10_dout[15:0]  )  //o
  );
  MulUnit mulUnit_3 (
    .a    (_zz_428[15:0]      ), //i
    .b    (_zz_429[15:0]      ), //i
    .c    (mulUnit_3_c[15:0]  )  //o
  );
  SInt16fixTo15_0_ROUNDTOINF fixTo_11 (
    .din     (_zz_430[15:0]        ), //i
    .dout    (fixTo_11_dout[15:0]  )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_12 (
    .din     (exp_wd_prod_real[31:0]  ), //i
    .dout    (fixTo_12_dout[15:0]     )  //o
  );
  SInt32fixTo23_8_ROUNDTOINF fixTo_13 (
    .din     (exp_wd_prod_imag[31:0]  ), //i
    .dout    (fixTo_13_dout[15:0]     )  //o
  );
  DivUnit divUnit_3 (
    .a    (_zz_431[15:0]      ), //i
    .b    (_zz_432[15:0]      ), //i
    .c    (divUnit_3_c[15:0]  )  //o
  );
  DivUnit divUnit_4 (
    .a    (_zz_433[15:0]      ), //i
    .b    (_zz_434[15:0]      ), //i
    .c    (divUnit_4_c[15:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_14 (
    .din     (_zz_435[31:0]        ), //i
    .dout    (fixTo_14_dout[31:0]  )  //o
  );
  SInt16fixTo31_0_ROUNDTOINF fixTo_15 (
    .din     (timeshift_real[15:0]  ), //i
    .dout    (fixTo_15_dout[31:0]   )  //o
  );
  MulUnit mulUnit_4 (
    .a    (_zz_436[31:0]      ), //i
    .b    (_zz_437[31:0]      ), //i
    .c    (mulUnit_4_c[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_16 (
    .din     (_zz_438[31:0]        ), //i
    .dout    (fixTo_16_dout[31:0]  )  //o
  );
  SInt16fixTo31_0_ROUNDTOINF fixTo_17 (
    .din     (_zz_439[15:0]        ), //i
    .dout    (fixTo_17_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_18 (
    .din     (exp_wd_prod_divw_real[31:0]  ), //i
    .dout    (fixTo_18_dout[31:0]          )  //o
  );
  MulUnit mulUnit_5 (
    .a    (_zz_440[31:0]      ), //i
    .b    (_zz_441[31:0]      ), //i
    .c    (mulUnit_5_c[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_19 (
    .din     (_zz_442[31:0]        ), //i
    .dout    (fixTo_19_dout[31:0]  )  //o
  );
  SInt16fixTo31_0_ROUNDTOINF fixTo_20 (
    .din     (_zz_443[15:0]        ), //i
    .dout    (fixTo_20_dout[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_21 (
    .din     (exp_wd_prod_divw_imag[31:0]  ), //i
    .dout    (fixTo_21_dout[31:0]          )  //o
  );
  MulUnit mulUnit_6 (
    .a    (_zz_444[31:0]      ), //i
    .b    (_zz_445[31:0]      ), //i
    .c    (mulUnit_6_c[31:0]  )  //o
  );
  SInt32fixTo31_0_ROUNDTOINF fixTo_22 (
    .din     (_zz_446[31:0]        ), //i
    .dout    (fixTo_22_dout[31:0]  )  //o
  );
  SInt64fixTo39_24_ROUNDTOINF fixTo_23 (
    .din     (_zz_411[63:0]        ), //i
    .dout    (fixTo_23_dout[15:0]  )  //o
  );
  SInt64fixTo39_24_ROUNDTOINF fixTo_24 (
    .din     (_zz_412[63:0]        ), //i
    .dout    (fixTo_24_dout[15:0]  )  //o
  );
  always @(*) begin
    case(_zz_395)
      7'b0000000 : begin
        _zz_447 = indx_table_0;
        _zz_448 = func_table_0_real;
        _zz_449 = func_table_0_imag;
      end
      7'b0000001 : begin
        _zz_447 = indx_table_1;
        _zz_448 = func_table_1_real;
        _zz_449 = func_table_1_imag;
      end
      7'b0000010 : begin
        _zz_447 = indx_table_2;
        _zz_448 = func_table_2_real;
        _zz_449 = func_table_2_imag;
      end
      7'b0000011 : begin
        _zz_447 = indx_table_3;
        _zz_448 = func_table_3_real;
        _zz_449 = func_table_3_imag;
      end
      7'b0000100 : begin
        _zz_447 = indx_table_4;
        _zz_448 = func_table_4_real;
        _zz_449 = func_table_4_imag;
      end
      7'b0000101 : begin
        _zz_447 = indx_table_5;
        _zz_448 = func_table_5_real;
        _zz_449 = func_table_5_imag;
      end
      7'b0000110 : begin
        _zz_447 = indx_table_6;
        _zz_448 = func_table_6_real;
        _zz_449 = func_table_6_imag;
      end
      7'b0000111 : begin
        _zz_447 = indx_table_7;
        _zz_448 = func_table_7_real;
        _zz_449 = func_table_7_imag;
      end
      7'b0001000 : begin
        _zz_447 = indx_table_8;
        _zz_448 = func_table_8_real;
        _zz_449 = func_table_8_imag;
      end
      7'b0001001 : begin
        _zz_447 = indx_table_9;
        _zz_448 = func_table_9_real;
        _zz_449 = func_table_9_imag;
      end
      7'b0001010 : begin
        _zz_447 = indx_table_10;
        _zz_448 = func_table_10_real;
        _zz_449 = func_table_10_imag;
      end
      7'b0001011 : begin
        _zz_447 = indx_table_11;
        _zz_448 = func_table_11_real;
        _zz_449 = func_table_11_imag;
      end
      7'b0001100 : begin
        _zz_447 = indx_table_12;
        _zz_448 = func_table_12_real;
        _zz_449 = func_table_12_imag;
      end
      7'b0001101 : begin
        _zz_447 = indx_table_13;
        _zz_448 = func_table_13_real;
        _zz_449 = func_table_13_imag;
      end
      7'b0001110 : begin
        _zz_447 = indx_table_14;
        _zz_448 = func_table_14_real;
        _zz_449 = func_table_14_imag;
      end
      7'b0001111 : begin
        _zz_447 = indx_table_15;
        _zz_448 = func_table_15_real;
        _zz_449 = func_table_15_imag;
      end
      7'b0010000 : begin
        _zz_447 = indx_table_16;
        _zz_448 = func_table_16_real;
        _zz_449 = func_table_16_imag;
      end
      7'b0010001 : begin
        _zz_447 = indx_table_17;
        _zz_448 = func_table_17_real;
        _zz_449 = func_table_17_imag;
      end
      7'b0010010 : begin
        _zz_447 = indx_table_18;
        _zz_448 = func_table_18_real;
        _zz_449 = func_table_18_imag;
      end
      7'b0010011 : begin
        _zz_447 = indx_table_19;
        _zz_448 = func_table_19_real;
        _zz_449 = func_table_19_imag;
      end
      7'b0010100 : begin
        _zz_447 = indx_table_20;
        _zz_448 = func_table_20_real;
        _zz_449 = func_table_20_imag;
      end
      7'b0010101 : begin
        _zz_447 = indx_table_21;
        _zz_448 = func_table_21_real;
        _zz_449 = func_table_21_imag;
      end
      7'b0010110 : begin
        _zz_447 = indx_table_22;
        _zz_448 = func_table_22_real;
        _zz_449 = func_table_22_imag;
      end
      7'b0010111 : begin
        _zz_447 = indx_table_23;
        _zz_448 = func_table_23_real;
        _zz_449 = func_table_23_imag;
      end
      7'b0011000 : begin
        _zz_447 = indx_table_24;
        _zz_448 = func_table_24_real;
        _zz_449 = func_table_24_imag;
      end
      7'b0011001 : begin
        _zz_447 = indx_table_25;
        _zz_448 = func_table_25_real;
        _zz_449 = func_table_25_imag;
      end
      7'b0011010 : begin
        _zz_447 = indx_table_26;
        _zz_448 = func_table_26_real;
        _zz_449 = func_table_26_imag;
      end
      7'b0011011 : begin
        _zz_447 = indx_table_27;
        _zz_448 = func_table_27_real;
        _zz_449 = func_table_27_imag;
      end
      7'b0011100 : begin
        _zz_447 = indx_table_28;
        _zz_448 = func_table_28_real;
        _zz_449 = func_table_28_imag;
      end
      7'b0011101 : begin
        _zz_447 = indx_table_29;
        _zz_448 = func_table_29_real;
        _zz_449 = func_table_29_imag;
      end
      7'b0011110 : begin
        _zz_447 = indx_table_30;
        _zz_448 = func_table_30_real;
        _zz_449 = func_table_30_imag;
      end
      7'b0011111 : begin
        _zz_447 = indx_table_31;
        _zz_448 = func_table_31_real;
        _zz_449 = func_table_31_imag;
      end
      7'b0100000 : begin
        _zz_447 = indx_table_32;
        _zz_448 = func_table_32_real;
        _zz_449 = func_table_32_imag;
      end
      7'b0100001 : begin
        _zz_447 = indx_table_33;
        _zz_448 = func_table_33_real;
        _zz_449 = func_table_33_imag;
      end
      7'b0100010 : begin
        _zz_447 = indx_table_34;
        _zz_448 = func_table_34_real;
        _zz_449 = func_table_34_imag;
      end
      7'b0100011 : begin
        _zz_447 = indx_table_35;
        _zz_448 = func_table_35_real;
        _zz_449 = func_table_35_imag;
      end
      7'b0100100 : begin
        _zz_447 = indx_table_36;
        _zz_448 = func_table_36_real;
        _zz_449 = func_table_36_imag;
      end
      7'b0100101 : begin
        _zz_447 = indx_table_37;
        _zz_448 = func_table_37_real;
        _zz_449 = func_table_37_imag;
      end
      7'b0100110 : begin
        _zz_447 = indx_table_38;
        _zz_448 = func_table_38_real;
        _zz_449 = func_table_38_imag;
      end
      7'b0100111 : begin
        _zz_447 = indx_table_39;
        _zz_448 = func_table_39_real;
        _zz_449 = func_table_39_imag;
      end
      7'b0101000 : begin
        _zz_447 = indx_table_40;
        _zz_448 = func_table_40_real;
        _zz_449 = func_table_40_imag;
      end
      7'b0101001 : begin
        _zz_447 = indx_table_41;
        _zz_448 = func_table_41_real;
        _zz_449 = func_table_41_imag;
      end
      7'b0101010 : begin
        _zz_447 = indx_table_42;
        _zz_448 = func_table_42_real;
        _zz_449 = func_table_42_imag;
      end
      7'b0101011 : begin
        _zz_447 = indx_table_43;
        _zz_448 = func_table_43_real;
        _zz_449 = func_table_43_imag;
      end
      7'b0101100 : begin
        _zz_447 = indx_table_44;
        _zz_448 = func_table_44_real;
        _zz_449 = func_table_44_imag;
      end
      7'b0101101 : begin
        _zz_447 = indx_table_45;
        _zz_448 = func_table_45_real;
        _zz_449 = func_table_45_imag;
      end
      7'b0101110 : begin
        _zz_447 = indx_table_46;
        _zz_448 = func_table_46_real;
        _zz_449 = func_table_46_imag;
      end
      7'b0101111 : begin
        _zz_447 = indx_table_47;
        _zz_448 = func_table_47_real;
        _zz_449 = func_table_47_imag;
      end
      7'b0110000 : begin
        _zz_447 = indx_table_48;
        _zz_448 = func_table_48_real;
        _zz_449 = func_table_48_imag;
      end
      7'b0110001 : begin
        _zz_447 = indx_table_49;
        _zz_448 = func_table_49_real;
        _zz_449 = func_table_49_imag;
      end
      7'b0110010 : begin
        _zz_447 = indx_table_50;
        _zz_448 = func_table_50_real;
        _zz_449 = func_table_50_imag;
      end
      7'b0110011 : begin
        _zz_447 = indx_table_51;
        _zz_448 = func_table_51_real;
        _zz_449 = func_table_51_imag;
      end
      7'b0110100 : begin
        _zz_447 = indx_table_52;
        _zz_448 = func_table_52_real;
        _zz_449 = func_table_52_imag;
      end
      7'b0110101 : begin
        _zz_447 = indx_table_53;
        _zz_448 = func_table_53_real;
        _zz_449 = func_table_53_imag;
      end
      7'b0110110 : begin
        _zz_447 = indx_table_54;
        _zz_448 = func_table_54_real;
        _zz_449 = func_table_54_imag;
      end
      7'b0110111 : begin
        _zz_447 = indx_table_55;
        _zz_448 = func_table_55_real;
        _zz_449 = func_table_55_imag;
      end
      7'b0111000 : begin
        _zz_447 = indx_table_56;
        _zz_448 = func_table_56_real;
        _zz_449 = func_table_56_imag;
      end
      7'b0111001 : begin
        _zz_447 = indx_table_57;
        _zz_448 = func_table_57_real;
        _zz_449 = func_table_57_imag;
      end
      7'b0111010 : begin
        _zz_447 = indx_table_58;
        _zz_448 = func_table_58_real;
        _zz_449 = func_table_58_imag;
      end
      7'b0111011 : begin
        _zz_447 = indx_table_59;
        _zz_448 = func_table_59_real;
        _zz_449 = func_table_59_imag;
      end
      7'b0111100 : begin
        _zz_447 = indx_table_60;
        _zz_448 = func_table_60_real;
        _zz_449 = func_table_60_imag;
      end
      7'b0111101 : begin
        _zz_447 = indx_table_61;
        _zz_448 = func_table_61_real;
        _zz_449 = func_table_61_imag;
      end
      7'b0111110 : begin
        _zz_447 = indx_table_62;
        _zz_448 = func_table_62_real;
        _zz_449 = func_table_62_imag;
      end
      7'b0111111 : begin
        _zz_447 = indx_table_63;
        _zz_448 = func_table_63_real;
        _zz_449 = func_table_63_imag;
      end
      7'b1000000 : begin
        _zz_447 = indx_table_64;
        _zz_448 = func_table_64_real;
        _zz_449 = func_table_64_imag;
      end
      7'b1000001 : begin
        _zz_447 = indx_table_65;
        _zz_448 = func_table_65_real;
        _zz_449 = func_table_65_imag;
      end
      7'b1000010 : begin
        _zz_447 = indx_table_66;
        _zz_448 = func_table_66_real;
        _zz_449 = func_table_66_imag;
      end
      7'b1000011 : begin
        _zz_447 = indx_table_67;
        _zz_448 = func_table_67_real;
        _zz_449 = func_table_67_imag;
      end
      7'b1000100 : begin
        _zz_447 = indx_table_68;
        _zz_448 = func_table_68_real;
        _zz_449 = func_table_68_imag;
      end
      7'b1000101 : begin
        _zz_447 = indx_table_69;
        _zz_448 = func_table_69_real;
        _zz_449 = func_table_69_imag;
      end
      7'b1000110 : begin
        _zz_447 = indx_table_70;
        _zz_448 = func_table_70_real;
        _zz_449 = func_table_70_imag;
      end
      7'b1000111 : begin
        _zz_447 = indx_table_71;
        _zz_448 = func_table_71_real;
        _zz_449 = func_table_71_imag;
      end
      7'b1001000 : begin
        _zz_447 = indx_table_72;
        _zz_448 = func_table_72_real;
        _zz_449 = func_table_72_imag;
      end
      7'b1001001 : begin
        _zz_447 = indx_table_73;
        _zz_448 = func_table_73_real;
        _zz_449 = func_table_73_imag;
      end
      7'b1001010 : begin
        _zz_447 = indx_table_74;
        _zz_448 = func_table_74_real;
        _zz_449 = func_table_74_imag;
      end
      7'b1001011 : begin
        _zz_447 = indx_table_75;
        _zz_448 = func_table_75_real;
        _zz_449 = func_table_75_imag;
      end
      7'b1001100 : begin
        _zz_447 = indx_table_76;
        _zz_448 = func_table_76_real;
        _zz_449 = func_table_76_imag;
      end
      7'b1001101 : begin
        _zz_447 = indx_table_77;
        _zz_448 = func_table_77_real;
        _zz_449 = func_table_77_imag;
      end
      7'b1001110 : begin
        _zz_447 = indx_table_78;
        _zz_448 = func_table_78_real;
        _zz_449 = func_table_78_imag;
      end
      7'b1001111 : begin
        _zz_447 = indx_table_79;
        _zz_448 = func_table_79_real;
        _zz_449 = func_table_79_imag;
      end
      7'b1010000 : begin
        _zz_447 = indx_table_80;
        _zz_448 = func_table_80_real;
        _zz_449 = func_table_80_imag;
      end
      7'b1010001 : begin
        _zz_447 = indx_table_81;
        _zz_448 = func_table_81_real;
        _zz_449 = func_table_81_imag;
      end
      7'b1010010 : begin
        _zz_447 = indx_table_82;
        _zz_448 = func_table_82_real;
        _zz_449 = func_table_82_imag;
      end
      7'b1010011 : begin
        _zz_447 = indx_table_83;
        _zz_448 = func_table_83_real;
        _zz_449 = func_table_83_imag;
      end
      7'b1010100 : begin
        _zz_447 = indx_table_84;
        _zz_448 = func_table_84_real;
        _zz_449 = func_table_84_imag;
      end
      7'b1010101 : begin
        _zz_447 = indx_table_85;
        _zz_448 = func_table_85_real;
        _zz_449 = func_table_85_imag;
      end
      7'b1010110 : begin
        _zz_447 = indx_table_86;
        _zz_448 = func_table_86_real;
        _zz_449 = func_table_86_imag;
      end
      7'b1010111 : begin
        _zz_447 = indx_table_87;
        _zz_448 = func_table_87_real;
        _zz_449 = func_table_87_imag;
      end
      7'b1011000 : begin
        _zz_447 = indx_table_88;
        _zz_448 = func_table_88_real;
        _zz_449 = func_table_88_imag;
      end
      7'b1011001 : begin
        _zz_447 = indx_table_89;
        _zz_448 = func_table_89_real;
        _zz_449 = func_table_89_imag;
      end
      7'b1011010 : begin
        _zz_447 = indx_table_90;
        _zz_448 = func_table_90_real;
        _zz_449 = func_table_90_imag;
      end
      7'b1011011 : begin
        _zz_447 = indx_table_91;
        _zz_448 = func_table_91_real;
        _zz_449 = func_table_91_imag;
      end
      7'b1011100 : begin
        _zz_447 = indx_table_92;
        _zz_448 = func_table_92_real;
        _zz_449 = func_table_92_imag;
      end
      7'b1011101 : begin
        _zz_447 = indx_table_93;
        _zz_448 = func_table_93_real;
        _zz_449 = func_table_93_imag;
      end
      7'b1011110 : begin
        _zz_447 = indx_table_94;
        _zz_448 = func_table_94_real;
        _zz_449 = func_table_94_imag;
      end
      7'b1011111 : begin
        _zz_447 = indx_table_95;
        _zz_448 = func_table_95_real;
        _zz_449 = func_table_95_imag;
      end
      7'b1100000 : begin
        _zz_447 = indx_table_96;
        _zz_448 = func_table_96_real;
        _zz_449 = func_table_96_imag;
      end
      7'b1100001 : begin
        _zz_447 = indx_table_97;
        _zz_448 = func_table_97_real;
        _zz_449 = func_table_97_imag;
      end
      7'b1100010 : begin
        _zz_447 = indx_table_98;
        _zz_448 = func_table_98_real;
        _zz_449 = func_table_98_imag;
      end
      7'b1100011 : begin
        _zz_447 = indx_table_99;
        _zz_448 = func_table_99_real;
        _zz_449 = func_table_99_imag;
      end
      7'b1100100 : begin
        _zz_447 = indx_table_100;
        _zz_448 = func_table_100_real;
        _zz_449 = func_table_100_imag;
      end
      7'b1100101 : begin
        _zz_447 = indx_table_101;
        _zz_448 = func_table_101_real;
        _zz_449 = func_table_101_imag;
      end
      7'b1100110 : begin
        _zz_447 = indx_table_102;
        _zz_448 = func_table_102_real;
        _zz_449 = func_table_102_imag;
      end
      7'b1100111 : begin
        _zz_447 = indx_table_103;
        _zz_448 = func_table_103_real;
        _zz_449 = func_table_103_imag;
      end
      7'b1101000 : begin
        _zz_447 = indx_table_104;
        _zz_448 = func_table_104_real;
        _zz_449 = func_table_104_imag;
      end
      7'b1101001 : begin
        _zz_447 = indx_table_105;
        _zz_448 = func_table_105_real;
        _zz_449 = func_table_105_imag;
      end
      7'b1101010 : begin
        _zz_447 = indx_table_106;
        _zz_448 = func_table_106_real;
        _zz_449 = func_table_106_imag;
      end
      7'b1101011 : begin
        _zz_447 = indx_table_107;
        _zz_448 = func_table_107_real;
        _zz_449 = func_table_107_imag;
      end
      7'b1101100 : begin
        _zz_447 = indx_table_108;
        _zz_448 = func_table_108_real;
        _zz_449 = func_table_108_imag;
      end
      7'b1101101 : begin
        _zz_447 = indx_table_109;
        _zz_448 = func_table_109_real;
        _zz_449 = func_table_109_imag;
      end
      7'b1101110 : begin
        _zz_447 = indx_table_110;
        _zz_448 = func_table_110_real;
        _zz_449 = func_table_110_imag;
      end
      7'b1101111 : begin
        _zz_447 = indx_table_111;
        _zz_448 = func_table_111_real;
        _zz_449 = func_table_111_imag;
      end
      7'b1110000 : begin
        _zz_447 = indx_table_112;
        _zz_448 = func_table_112_real;
        _zz_449 = func_table_112_imag;
      end
      7'b1110001 : begin
        _zz_447 = indx_table_113;
        _zz_448 = func_table_113_real;
        _zz_449 = func_table_113_imag;
      end
      7'b1110010 : begin
        _zz_447 = indx_table_114;
        _zz_448 = func_table_114_real;
        _zz_449 = func_table_114_imag;
      end
      7'b1110011 : begin
        _zz_447 = indx_table_115;
        _zz_448 = func_table_115_real;
        _zz_449 = func_table_115_imag;
      end
      7'b1110100 : begin
        _zz_447 = indx_table_116;
        _zz_448 = func_table_116_real;
        _zz_449 = func_table_116_imag;
      end
      7'b1110101 : begin
        _zz_447 = indx_table_117;
        _zz_448 = func_table_117_real;
        _zz_449 = func_table_117_imag;
      end
      7'b1110110 : begin
        _zz_447 = indx_table_118;
        _zz_448 = func_table_118_real;
        _zz_449 = func_table_118_imag;
      end
      7'b1110111 : begin
        _zz_447 = indx_table_119;
        _zz_448 = func_table_119_real;
        _zz_449 = func_table_119_imag;
      end
      7'b1111000 : begin
        _zz_447 = indx_table_120;
        _zz_448 = func_table_120_real;
        _zz_449 = func_table_120_imag;
      end
      7'b1111001 : begin
        _zz_447 = indx_table_121;
        _zz_448 = func_table_121_real;
        _zz_449 = func_table_121_imag;
      end
      7'b1111010 : begin
        _zz_447 = indx_table_122;
        _zz_448 = func_table_122_real;
        _zz_449 = func_table_122_imag;
      end
      7'b1111011 : begin
        _zz_447 = indx_table_123;
        _zz_448 = func_table_123_real;
        _zz_449 = func_table_123_imag;
      end
      7'b1111100 : begin
        _zz_447 = indx_table_124;
        _zz_448 = func_table_124_real;
        _zz_449 = func_table_124_imag;
      end
      7'b1111101 : begin
        _zz_447 = indx_table_125;
        _zz_448 = func_table_125_real;
        _zz_449 = func_table_125_imag;
      end
      7'b1111110 : begin
        _zz_447 = indx_table_126;
        _zz_448 = func_table_126_real;
        _zz_449 = func_table_126_imag;
      end
      default : begin
        _zz_447 = indx_table_127;
        _zz_448 = func_table_127_real;
        _zz_449 = func_table_127_imag;
      end
    endcase
  end

  always @(*) begin
    case(lzc)
      7'b0000000 : begin
        _zz_450 = indx_table_0;
        _zz_451 = func_table_0_real;
        _zz_452 = func_table_0_imag;
      end
      7'b0000001 : begin
        _zz_450 = indx_table_1;
        _zz_451 = func_table_1_real;
        _zz_452 = func_table_1_imag;
      end
      7'b0000010 : begin
        _zz_450 = indx_table_2;
        _zz_451 = func_table_2_real;
        _zz_452 = func_table_2_imag;
      end
      7'b0000011 : begin
        _zz_450 = indx_table_3;
        _zz_451 = func_table_3_real;
        _zz_452 = func_table_3_imag;
      end
      7'b0000100 : begin
        _zz_450 = indx_table_4;
        _zz_451 = func_table_4_real;
        _zz_452 = func_table_4_imag;
      end
      7'b0000101 : begin
        _zz_450 = indx_table_5;
        _zz_451 = func_table_5_real;
        _zz_452 = func_table_5_imag;
      end
      7'b0000110 : begin
        _zz_450 = indx_table_6;
        _zz_451 = func_table_6_real;
        _zz_452 = func_table_6_imag;
      end
      7'b0000111 : begin
        _zz_450 = indx_table_7;
        _zz_451 = func_table_7_real;
        _zz_452 = func_table_7_imag;
      end
      7'b0001000 : begin
        _zz_450 = indx_table_8;
        _zz_451 = func_table_8_real;
        _zz_452 = func_table_8_imag;
      end
      7'b0001001 : begin
        _zz_450 = indx_table_9;
        _zz_451 = func_table_9_real;
        _zz_452 = func_table_9_imag;
      end
      7'b0001010 : begin
        _zz_450 = indx_table_10;
        _zz_451 = func_table_10_real;
        _zz_452 = func_table_10_imag;
      end
      7'b0001011 : begin
        _zz_450 = indx_table_11;
        _zz_451 = func_table_11_real;
        _zz_452 = func_table_11_imag;
      end
      7'b0001100 : begin
        _zz_450 = indx_table_12;
        _zz_451 = func_table_12_real;
        _zz_452 = func_table_12_imag;
      end
      7'b0001101 : begin
        _zz_450 = indx_table_13;
        _zz_451 = func_table_13_real;
        _zz_452 = func_table_13_imag;
      end
      7'b0001110 : begin
        _zz_450 = indx_table_14;
        _zz_451 = func_table_14_real;
        _zz_452 = func_table_14_imag;
      end
      7'b0001111 : begin
        _zz_450 = indx_table_15;
        _zz_451 = func_table_15_real;
        _zz_452 = func_table_15_imag;
      end
      7'b0010000 : begin
        _zz_450 = indx_table_16;
        _zz_451 = func_table_16_real;
        _zz_452 = func_table_16_imag;
      end
      7'b0010001 : begin
        _zz_450 = indx_table_17;
        _zz_451 = func_table_17_real;
        _zz_452 = func_table_17_imag;
      end
      7'b0010010 : begin
        _zz_450 = indx_table_18;
        _zz_451 = func_table_18_real;
        _zz_452 = func_table_18_imag;
      end
      7'b0010011 : begin
        _zz_450 = indx_table_19;
        _zz_451 = func_table_19_real;
        _zz_452 = func_table_19_imag;
      end
      7'b0010100 : begin
        _zz_450 = indx_table_20;
        _zz_451 = func_table_20_real;
        _zz_452 = func_table_20_imag;
      end
      7'b0010101 : begin
        _zz_450 = indx_table_21;
        _zz_451 = func_table_21_real;
        _zz_452 = func_table_21_imag;
      end
      7'b0010110 : begin
        _zz_450 = indx_table_22;
        _zz_451 = func_table_22_real;
        _zz_452 = func_table_22_imag;
      end
      7'b0010111 : begin
        _zz_450 = indx_table_23;
        _zz_451 = func_table_23_real;
        _zz_452 = func_table_23_imag;
      end
      7'b0011000 : begin
        _zz_450 = indx_table_24;
        _zz_451 = func_table_24_real;
        _zz_452 = func_table_24_imag;
      end
      7'b0011001 : begin
        _zz_450 = indx_table_25;
        _zz_451 = func_table_25_real;
        _zz_452 = func_table_25_imag;
      end
      7'b0011010 : begin
        _zz_450 = indx_table_26;
        _zz_451 = func_table_26_real;
        _zz_452 = func_table_26_imag;
      end
      7'b0011011 : begin
        _zz_450 = indx_table_27;
        _zz_451 = func_table_27_real;
        _zz_452 = func_table_27_imag;
      end
      7'b0011100 : begin
        _zz_450 = indx_table_28;
        _zz_451 = func_table_28_real;
        _zz_452 = func_table_28_imag;
      end
      7'b0011101 : begin
        _zz_450 = indx_table_29;
        _zz_451 = func_table_29_real;
        _zz_452 = func_table_29_imag;
      end
      7'b0011110 : begin
        _zz_450 = indx_table_30;
        _zz_451 = func_table_30_real;
        _zz_452 = func_table_30_imag;
      end
      7'b0011111 : begin
        _zz_450 = indx_table_31;
        _zz_451 = func_table_31_real;
        _zz_452 = func_table_31_imag;
      end
      7'b0100000 : begin
        _zz_450 = indx_table_32;
        _zz_451 = func_table_32_real;
        _zz_452 = func_table_32_imag;
      end
      7'b0100001 : begin
        _zz_450 = indx_table_33;
        _zz_451 = func_table_33_real;
        _zz_452 = func_table_33_imag;
      end
      7'b0100010 : begin
        _zz_450 = indx_table_34;
        _zz_451 = func_table_34_real;
        _zz_452 = func_table_34_imag;
      end
      7'b0100011 : begin
        _zz_450 = indx_table_35;
        _zz_451 = func_table_35_real;
        _zz_452 = func_table_35_imag;
      end
      7'b0100100 : begin
        _zz_450 = indx_table_36;
        _zz_451 = func_table_36_real;
        _zz_452 = func_table_36_imag;
      end
      7'b0100101 : begin
        _zz_450 = indx_table_37;
        _zz_451 = func_table_37_real;
        _zz_452 = func_table_37_imag;
      end
      7'b0100110 : begin
        _zz_450 = indx_table_38;
        _zz_451 = func_table_38_real;
        _zz_452 = func_table_38_imag;
      end
      7'b0100111 : begin
        _zz_450 = indx_table_39;
        _zz_451 = func_table_39_real;
        _zz_452 = func_table_39_imag;
      end
      7'b0101000 : begin
        _zz_450 = indx_table_40;
        _zz_451 = func_table_40_real;
        _zz_452 = func_table_40_imag;
      end
      7'b0101001 : begin
        _zz_450 = indx_table_41;
        _zz_451 = func_table_41_real;
        _zz_452 = func_table_41_imag;
      end
      7'b0101010 : begin
        _zz_450 = indx_table_42;
        _zz_451 = func_table_42_real;
        _zz_452 = func_table_42_imag;
      end
      7'b0101011 : begin
        _zz_450 = indx_table_43;
        _zz_451 = func_table_43_real;
        _zz_452 = func_table_43_imag;
      end
      7'b0101100 : begin
        _zz_450 = indx_table_44;
        _zz_451 = func_table_44_real;
        _zz_452 = func_table_44_imag;
      end
      7'b0101101 : begin
        _zz_450 = indx_table_45;
        _zz_451 = func_table_45_real;
        _zz_452 = func_table_45_imag;
      end
      7'b0101110 : begin
        _zz_450 = indx_table_46;
        _zz_451 = func_table_46_real;
        _zz_452 = func_table_46_imag;
      end
      7'b0101111 : begin
        _zz_450 = indx_table_47;
        _zz_451 = func_table_47_real;
        _zz_452 = func_table_47_imag;
      end
      7'b0110000 : begin
        _zz_450 = indx_table_48;
        _zz_451 = func_table_48_real;
        _zz_452 = func_table_48_imag;
      end
      7'b0110001 : begin
        _zz_450 = indx_table_49;
        _zz_451 = func_table_49_real;
        _zz_452 = func_table_49_imag;
      end
      7'b0110010 : begin
        _zz_450 = indx_table_50;
        _zz_451 = func_table_50_real;
        _zz_452 = func_table_50_imag;
      end
      7'b0110011 : begin
        _zz_450 = indx_table_51;
        _zz_451 = func_table_51_real;
        _zz_452 = func_table_51_imag;
      end
      7'b0110100 : begin
        _zz_450 = indx_table_52;
        _zz_451 = func_table_52_real;
        _zz_452 = func_table_52_imag;
      end
      7'b0110101 : begin
        _zz_450 = indx_table_53;
        _zz_451 = func_table_53_real;
        _zz_452 = func_table_53_imag;
      end
      7'b0110110 : begin
        _zz_450 = indx_table_54;
        _zz_451 = func_table_54_real;
        _zz_452 = func_table_54_imag;
      end
      7'b0110111 : begin
        _zz_450 = indx_table_55;
        _zz_451 = func_table_55_real;
        _zz_452 = func_table_55_imag;
      end
      7'b0111000 : begin
        _zz_450 = indx_table_56;
        _zz_451 = func_table_56_real;
        _zz_452 = func_table_56_imag;
      end
      7'b0111001 : begin
        _zz_450 = indx_table_57;
        _zz_451 = func_table_57_real;
        _zz_452 = func_table_57_imag;
      end
      7'b0111010 : begin
        _zz_450 = indx_table_58;
        _zz_451 = func_table_58_real;
        _zz_452 = func_table_58_imag;
      end
      7'b0111011 : begin
        _zz_450 = indx_table_59;
        _zz_451 = func_table_59_real;
        _zz_452 = func_table_59_imag;
      end
      7'b0111100 : begin
        _zz_450 = indx_table_60;
        _zz_451 = func_table_60_real;
        _zz_452 = func_table_60_imag;
      end
      7'b0111101 : begin
        _zz_450 = indx_table_61;
        _zz_451 = func_table_61_real;
        _zz_452 = func_table_61_imag;
      end
      7'b0111110 : begin
        _zz_450 = indx_table_62;
        _zz_451 = func_table_62_real;
        _zz_452 = func_table_62_imag;
      end
      7'b0111111 : begin
        _zz_450 = indx_table_63;
        _zz_451 = func_table_63_real;
        _zz_452 = func_table_63_imag;
      end
      7'b1000000 : begin
        _zz_450 = indx_table_64;
        _zz_451 = func_table_64_real;
        _zz_452 = func_table_64_imag;
      end
      7'b1000001 : begin
        _zz_450 = indx_table_65;
        _zz_451 = func_table_65_real;
        _zz_452 = func_table_65_imag;
      end
      7'b1000010 : begin
        _zz_450 = indx_table_66;
        _zz_451 = func_table_66_real;
        _zz_452 = func_table_66_imag;
      end
      7'b1000011 : begin
        _zz_450 = indx_table_67;
        _zz_451 = func_table_67_real;
        _zz_452 = func_table_67_imag;
      end
      7'b1000100 : begin
        _zz_450 = indx_table_68;
        _zz_451 = func_table_68_real;
        _zz_452 = func_table_68_imag;
      end
      7'b1000101 : begin
        _zz_450 = indx_table_69;
        _zz_451 = func_table_69_real;
        _zz_452 = func_table_69_imag;
      end
      7'b1000110 : begin
        _zz_450 = indx_table_70;
        _zz_451 = func_table_70_real;
        _zz_452 = func_table_70_imag;
      end
      7'b1000111 : begin
        _zz_450 = indx_table_71;
        _zz_451 = func_table_71_real;
        _zz_452 = func_table_71_imag;
      end
      7'b1001000 : begin
        _zz_450 = indx_table_72;
        _zz_451 = func_table_72_real;
        _zz_452 = func_table_72_imag;
      end
      7'b1001001 : begin
        _zz_450 = indx_table_73;
        _zz_451 = func_table_73_real;
        _zz_452 = func_table_73_imag;
      end
      7'b1001010 : begin
        _zz_450 = indx_table_74;
        _zz_451 = func_table_74_real;
        _zz_452 = func_table_74_imag;
      end
      7'b1001011 : begin
        _zz_450 = indx_table_75;
        _zz_451 = func_table_75_real;
        _zz_452 = func_table_75_imag;
      end
      7'b1001100 : begin
        _zz_450 = indx_table_76;
        _zz_451 = func_table_76_real;
        _zz_452 = func_table_76_imag;
      end
      7'b1001101 : begin
        _zz_450 = indx_table_77;
        _zz_451 = func_table_77_real;
        _zz_452 = func_table_77_imag;
      end
      7'b1001110 : begin
        _zz_450 = indx_table_78;
        _zz_451 = func_table_78_real;
        _zz_452 = func_table_78_imag;
      end
      7'b1001111 : begin
        _zz_450 = indx_table_79;
        _zz_451 = func_table_79_real;
        _zz_452 = func_table_79_imag;
      end
      7'b1010000 : begin
        _zz_450 = indx_table_80;
        _zz_451 = func_table_80_real;
        _zz_452 = func_table_80_imag;
      end
      7'b1010001 : begin
        _zz_450 = indx_table_81;
        _zz_451 = func_table_81_real;
        _zz_452 = func_table_81_imag;
      end
      7'b1010010 : begin
        _zz_450 = indx_table_82;
        _zz_451 = func_table_82_real;
        _zz_452 = func_table_82_imag;
      end
      7'b1010011 : begin
        _zz_450 = indx_table_83;
        _zz_451 = func_table_83_real;
        _zz_452 = func_table_83_imag;
      end
      7'b1010100 : begin
        _zz_450 = indx_table_84;
        _zz_451 = func_table_84_real;
        _zz_452 = func_table_84_imag;
      end
      7'b1010101 : begin
        _zz_450 = indx_table_85;
        _zz_451 = func_table_85_real;
        _zz_452 = func_table_85_imag;
      end
      7'b1010110 : begin
        _zz_450 = indx_table_86;
        _zz_451 = func_table_86_real;
        _zz_452 = func_table_86_imag;
      end
      7'b1010111 : begin
        _zz_450 = indx_table_87;
        _zz_451 = func_table_87_real;
        _zz_452 = func_table_87_imag;
      end
      7'b1011000 : begin
        _zz_450 = indx_table_88;
        _zz_451 = func_table_88_real;
        _zz_452 = func_table_88_imag;
      end
      7'b1011001 : begin
        _zz_450 = indx_table_89;
        _zz_451 = func_table_89_real;
        _zz_452 = func_table_89_imag;
      end
      7'b1011010 : begin
        _zz_450 = indx_table_90;
        _zz_451 = func_table_90_real;
        _zz_452 = func_table_90_imag;
      end
      7'b1011011 : begin
        _zz_450 = indx_table_91;
        _zz_451 = func_table_91_real;
        _zz_452 = func_table_91_imag;
      end
      7'b1011100 : begin
        _zz_450 = indx_table_92;
        _zz_451 = func_table_92_real;
        _zz_452 = func_table_92_imag;
      end
      7'b1011101 : begin
        _zz_450 = indx_table_93;
        _zz_451 = func_table_93_real;
        _zz_452 = func_table_93_imag;
      end
      7'b1011110 : begin
        _zz_450 = indx_table_94;
        _zz_451 = func_table_94_real;
        _zz_452 = func_table_94_imag;
      end
      7'b1011111 : begin
        _zz_450 = indx_table_95;
        _zz_451 = func_table_95_real;
        _zz_452 = func_table_95_imag;
      end
      7'b1100000 : begin
        _zz_450 = indx_table_96;
        _zz_451 = func_table_96_real;
        _zz_452 = func_table_96_imag;
      end
      7'b1100001 : begin
        _zz_450 = indx_table_97;
        _zz_451 = func_table_97_real;
        _zz_452 = func_table_97_imag;
      end
      7'b1100010 : begin
        _zz_450 = indx_table_98;
        _zz_451 = func_table_98_real;
        _zz_452 = func_table_98_imag;
      end
      7'b1100011 : begin
        _zz_450 = indx_table_99;
        _zz_451 = func_table_99_real;
        _zz_452 = func_table_99_imag;
      end
      7'b1100100 : begin
        _zz_450 = indx_table_100;
        _zz_451 = func_table_100_real;
        _zz_452 = func_table_100_imag;
      end
      7'b1100101 : begin
        _zz_450 = indx_table_101;
        _zz_451 = func_table_101_real;
        _zz_452 = func_table_101_imag;
      end
      7'b1100110 : begin
        _zz_450 = indx_table_102;
        _zz_451 = func_table_102_real;
        _zz_452 = func_table_102_imag;
      end
      7'b1100111 : begin
        _zz_450 = indx_table_103;
        _zz_451 = func_table_103_real;
        _zz_452 = func_table_103_imag;
      end
      7'b1101000 : begin
        _zz_450 = indx_table_104;
        _zz_451 = func_table_104_real;
        _zz_452 = func_table_104_imag;
      end
      7'b1101001 : begin
        _zz_450 = indx_table_105;
        _zz_451 = func_table_105_real;
        _zz_452 = func_table_105_imag;
      end
      7'b1101010 : begin
        _zz_450 = indx_table_106;
        _zz_451 = func_table_106_real;
        _zz_452 = func_table_106_imag;
      end
      7'b1101011 : begin
        _zz_450 = indx_table_107;
        _zz_451 = func_table_107_real;
        _zz_452 = func_table_107_imag;
      end
      7'b1101100 : begin
        _zz_450 = indx_table_108;
        _zz_451 = func_table_108_real;
        _zz_452 = func_table_108_imag;
      end
      7'b1101101 : begin
        _zz_450 = indx_table_109;
        _zz_451 = func_table_109_real;
        _zz_452 = func_table_109_imag;
      end
      7'b1101110 : begin
        _zz_450 = indx_table_110;
        _zz_451 = func_table_110_real;
        _zz_452 = func_table_110_imag;
      end
      7'b1101111 : begin
        _zz_450 = indx_table_111;
        _zz_451 = func_table_111_real;
        _zz_452 = func_table_111_imag;
      end
      7'b1110000 : begin
        _zz_450 = indx_table_112;
        _zz_451 = func_table_112_real;
        _zz_452 = func_table_112_imag;
      end
      7'b1110001 : begin
        _zz_450 = indx_table_113;
        _zz_451 = func_table_113_real;
        _zz_452 = func_table_113_imag;
      end
      7'b1110010 : begin
        _zz_450 = indx_table_114;
        _zz_451 = func_table_114_real;
        _zz_452 = func_table_114_imag;
      end
      7'b1110011 : begin
        _zz_450 = indx_table_115;
        _zz_451 = func_table_115_real;
        _zz_452 = func_table_115_imag;
      end
      7'b1110100 : begin
        _zz_450 = indx_table_116;
        _zz_451 = func_table_116_real;
        _zz_452 = func_table_116_imag;
      end
      7'b1110101 : begin
        _zz_450 = indx_table_117;
        _zz_451 = func_table_117_real;
        _zz_452 = func_table_117_imag;
      end
      7'b1110110 : begin
        _zz_450 = indx_table_118;
        _zz_451 = func_table_118_real;
        _zz_452 = func_table_118_imag;
      end
      7'b1110111 : begin
        _zz_450 = indx_table_119;
        _zz_451 = func_table_119_real;
        _zz_452 = func_table_119_imag;
      end
      7'b1111000 : begin
        _zz_450 = indx_table_120;
        _zz_451 = func_table_120_real;
        _zz_452 = func_table_120_imag;
      end
      7'b1111001 : begin
        _zz_450 = indx_table_121;
        _zz_451 = func_table_121_real;
        _zz_452 = func_table_121_imag;
      end
      7'b1111010 : begin
        _zz_450 = indx_table_122;
        _zz_451 = func_table_122_real;
        _zz_452 = func_table_122_imag;
      end
      7'b1111011 : begin
        _zz_450 = indx_table_123;
        _zz_451 = func_table_123_real;
        _zz_452 = func_table_123_imag;
      end
      7'b1111100 : begin
        _zz_450 = indx_table_124;
        _zz_451 = func_table_124_real;
        _zz_452 = func_table_124_imag;
      end
      7'b1111101 : begin
        _zz_450 = indx_table_125;
        _zz_451 = func_table_125_real;
        _zz_452 = func_table_125_imag;
      end
      7'b1111110 : begin
        _zz_450 = indx_table_126;
        _zz_451 = func_table_126_real;
        _zz_452 = func_table_126_imag;
      end
      default : begin
        _zz_450 = indx_table_127;
        _zz_451 = func_table_127_real;
        _zz_452 = func_table_127_imag;
      end
    endcase
  end

  assign func_table_0_real = 16'h00e1;
  assign func_table_0_imag = 16'h0078;
  assign func_table_1_real = 16'h008e;
  assign func_table_1_imag = 16'h00d4;
  assign func_table_2_real = 16'h0019;
  assign func_table_2_imag = 16'h00fe;
  assign func_table_3_real = 16'hff9f;
  assign func_table_3_imag = 16'h00ec;
  assign func_table_4_real = 16'hff3b;
  assign func_table_4_imag = 16'h00a2;
  assign func_table_5_real = 16'hff05;
  assign func_table_5_imag = 16'h0031;
  assign func_table_6_real = 16'hff0c;
  assign func_table_6_imag = 16'hffb6;
  assign func_table_7_real = 16'hff4b;
  assign func_table_7_imag = 16'hff4b;
  assign func_table_8_real = 16'hffb6;
  assign func_table_8_imag = 16'hff0c;
  assign func_table_9_real = 16'h0031;
  assign func_table_9_imag = 16'hff05;
  assign func_table_10_real = 16'h00a2;
  assign func_table_10_imag = 16'hff3b;
  assign func_table_11_real = 16'h00ec;
  assign func_table_11_imag = 16'hff9f;
  assign func_table_12_real = 16'h00fe;
  assign func_table_12_imag = 16'h0019;
  assign func_table_13_real = 16'h00d4;
  assign func_table_13_imag = 16'h008e;
  assign func_table_14_real = 16'h0078;
  assign func_table_14_imag = 16'h00e1;
  assign func_table_15_real = 16'h0;
  assign func_table_15_imag = 16'h0100;
  assign func_table_16_real = 16'hff88;
  assign func_table_16_imag = 16'h00e1;
  assign func_table_17_real = 16'hff2c;
  assign func_table_17_imag = 16'h008e;
  assign func_table_18_real = 16'hff02;
  assign func_table_18_imag = 16'h0019;
  assign func_table_19_real = 16'hff14;
  assign func_table_19_imag = 16'hff9f;
  assign func_table_20_real = 16'hff5e;
  assign func_table_20_imag = 16'hff3b;
  assign func_table_21_real = 16'hffcf;
  assign func_table_21_imag = 16'hff05;
  assign func_table_22_real = 16'h004a;
  assign func_table_22_imag = 16'hff0c;
  assign func_table_23_real = 16'h00b5;
  assign func_table_23_imag = 16'hff4b;
  assign func_table_24_real = 16'h00f4;
  assign func_table_24_imag = 16'hffb6;
  assign func_table_25_real = 16'h00fb;
  assign func_table_25_imag = 16'h0031;
  assign func_table_26_real = 16'h00c5;
  assign func_table_26_imag = 16'h00a2;
  assign func_table_27_real = 16'h0061;
  assign func_table_27_imag = 16'h00ec;
  assign func_table_28_real = 16'hffe7;
  assign func_table_28_imag = 16'h00fe;
  assign func_table_29_real = 16'hff72;
  assign func_table_29_imag = 16'h00d4;
  assign func_table_30_real = 16'hff1f;
  assign func_table_30_imag = 16'h0078;
  assign func_table_31_real = 16'hff00;
  assign func_table_31_imag = 16'h0;
  assign func_table_32_real = 16'hff1f;
  assign func_table_32_imag = 16'hff88;
  assign func_table_33_real = 16'hff72;
  assign func_table_33_imag = 16'hff2c;
  assign func_table_34_real = 16'hffe7;
  assign func_table_34_imag = 16'hff02;
  assign func_table_35_real = 16'h0061;
  assign func_table_35_imag = 16'hff14;
  assign func_table_36_real = 16'h00c5;
  assign func_table_36_imag = 16'hff5e;
  assign func_table_37_real = 16'h00fb;
  assign func_table_37_imag = 16'hffcf;
  assign func_table_38_real = 16'h00f4;
  assign func_table_38_imag = 16'h004a;
  assign func_table_39_real = 16'h00b5;
  assign func_table_39_imag = 16'h00b5;
  assign func_table_40_real = 16'h004a;
  assign func_table_40_imag = 16'h00f4;
  assign func_table_41_real = 16'hffcf;
  assign func_table_41_imag = 16'h00fb;
  assign func_table_42_real = 16'hff5e;
  assign func_table_42_imag = 16'h00c5;
  assign func_table_43_real = 16'hff14;
  assign func_table_43_imag = 16'h0061;
  assign func_table_44_real = 16'hff02;
  assign func_table_44_imag = 16'hffe7;
  assign func_table_45_real = 16'hff2c;
  assign func_table_45_imag = 16'hff72;
  assign func_table_46_real = 16'hff88;
  assign func_table_46_imag = 16'hff1f;
  assign func_table_47_real = 16'h0;
  assign func_table_47_imag = 16'hff00;
  assign func_table_48_real = 16'h0078;
  assign func_table_48_imag = 16'hff1f;
  assign func_table_49_real = 16'h00d4;
  assign func_table_49_imag = 16'hff72;
  assign func_table_50_real = 16'h00fe;
  assign func_table_50_imag = 16'hffe7;
  assign func_table_51_real = 16'h00ec;
  assign func_table_51_imag = 16'h0061;
  assign func_table_52_real = 16'h00a2;
  assign func_table_52_imag = 16'h00c5;
  assign func_table_53_real = 16'h0031;
  assign func_table_53_imag = 16'h00fb;
  assign func_table_54_real = 16'hffb6;
  assign func_table_54_imag = 16'h00f4;
  assign func_table_55_real = 16'hff4b;
  assign func_table_55_imag = 16'h00b5;
  assign func_table_56_real = 16'hff0c;
  assign func_table_56_imag = 16'h004a;
  assign func_table_57_real = 16'hff05;
  assign func_table_57_imag = 16'hffcf;
  assign func_table_58_real = 16'hff3b;
  assign func_table_58_imag = 16'hff5e;
  assign func_table_59_real = 16'hff9f;
  assign func_table_59_imag = 16'hff14;
  assign func_table_60_real = 16'h0019;
  assign func_table_60_imag = 16'hff02;
  assign func_table_61_real = 16'h008e;
  assign func_table_61_imag = 16'hff2c;
  assign func_table_62_real = 16'h00e1;
  assign func_table_62_imag = 16'hff88;
  assign func_table_63_real = 16'h0100;
  assign func_table_63_imag = 16'h0;
  assign func_table_64_real = 16'h00e1;
  assign func_table_64_imag = 16'h0078;
  assign func_table_65_real = 16'h008e;
  assign func_table_65_imag = 16'h00d4;
  assign func_table_66_real = 16'h0019;
  assign func_table_66_imag = 16'h00fe;
  assign func_table_67_real = 16'hff9f;
  assign func_table_67_imag = 16'h00ec;
  assign func_table_68_real = 16'hff3b;
  assign func_table_68_imag = 16'h00a2;
  assign func_table_69_real = 16'hff05;
  assign func_table_69_imag = 16'h0031;
  assign func_table_70_real = 16'hff0c;
  assign func_table_70_imag = 16'hffb6;
  assign func_table_71_real = 16'hff4b;
  assign func_table_71_imag = 16'hff4b;
  assign func_table_72_real = 16'hffb6;
  assign func_table_72_imag = 16'hff0c;
  assign func_table_73_real = 16'h0031;
  assign func_table_73_imag = 16'hff05;
  assign func_table_74_real = 16'h00a2;
  assign func_table_74_imag = 16'hff3b;
  assign func_table_75_real = 16'h00ec;
  assign func_table_75_imag = 16'hff9f;
  assign func_table_76_real = 16'h00fe;
  assign func_table_76_imag = 16'h0019;
  assign func_table_77_real = 16'h00d4;
  assign func_table_77_imag = 16'h008e;
  assign func_table_78_real = 16'h0078;
  assign func_table_78_imag = 16'h00e1;
  assign func_table_79_real = 16'h0;
  assign func_table_79_imag = 16'h0100;
  assign func_table_80_real = 16'hff88;
  assign func_table_80_imag = 16'h00e1;
  assign func_table_81_real = 16'hff2c;
  assign func_table_81_imag = 16'h008e;
  assign func_table_82_real = 16'hff02;
  assign func_table_82_imag = 16'h0019;
  assign func_table_83_real = 16'hff14;
  assign func_table_83_imag = 16'hff9f;
  assign func_table_84_real = 16'hff5e;
  assign func_table_84_imag = 16'hff3b;
  assign func_table_85_real = 16'hffcf;
  assign func_table_85_imag = 16'hff05;
  assign func_table_86_real = 16'h004a;
  assign func_table_86_imag = 16'hff0c;
  assign func_table_87_real = 16'h00b5;
  assign func_table_87_imag = 16'hff4b;
  assign func_table_88_real = 16'h00f4;
  assign func_table_88_imag = 16'hffb6;
  assign func_table_89_real = 16'h00fb;
  assign func_table_89_imag = 16'h0031;
  assign func_table_90_real = 16'h00c5;
  assign func_table_90_imag = 16'h00a2;
  assign func_table_91_real = 16'h0061;
  assign func_table_91_imag = 16'h00ec;
  assign func_table_92_real = 16'hffe7;
  assign func_table_92_imag = 16'h00fe;
  assign func_table_93_real = 16'hff72;
  assign func_table_93_imag = 16'h00d4;
  assign func_table_94_real = 16'hff1f;
  assign func_table_94_imag = 16'h0078;
  assign func_table_95_real = 16'hff00;
  assign func_table_95_imag = 16'h0;
  assign func_table_96_real = 16'hff1f;
  assign func_table_96_imag = 16'hff88;
  assign func_table_97_real = 16'hff72;
  assign func_table_97_imag = 16'hff2c;
  assign func_table_98_real = 16'hffe7;
  assign func_table_98_imag = 16'hff02;
  assign func_table_99_real = 16'h0061;
  assign func_table_99_imag = 16'hff14;
  assign func_table_100_real = 16'h00c5;
  assign func_table_100_imag = 16'hff5e;
  assign func_table_101_real = 16'h00fb;
  assign func_table_101_imag = 16'hffcf;
  assign func_table_102_real = 16'h00f4;
  assign func_table_102_imag = 16'h004a;
  assign func_table_103_real = 16'h00b5;
  assign func_table_103_imag = 16'h00b5;
  assign func_table_104_real = 16'h004a;
  assign func_table_104_imag = 16'h00f4;
  assign func_table_105_real = 16'hffcf;
  assign func_table_105_imag = 16'h00fb;
  assign func_table_106_real = 16'hff5e;
  assign func_table_106_imag = 16'h00c5;
  assign func_table_107_real = 16'hff14;
  assign func_table_107_imag = 16'h0061;
  assign func_table_108_real = 16'hff02;
  assign func_table_108_imag = 16'hffe7;
  assign func_table_109_real = 16'hff2c;
  assign func_table_109_imag = 16'hff72;
  assign func_table_110_real = 16'hff88;
  assign func_table_110_imag = 16'hff1f;
  assign func_table_111_real = 16'h0;
  assign func_table_111_imag = 16'hff00;
  assign func_table_112_real = 16'h0078;
  assign func_table_112_imag = 16'hff1f;
  assign func_table_113_real = 16'h00d4;
  assign func_table_113_imag = 16'hff72;
  assign func_table_114_real = 16'h00fe;
  assign func_table_114_imag = 16'hffe7;
  assign func_table_115_real = 16'h00ec;
  assign func_table_115_imag = 16'h0061;
  assign func_table_116_real = 16'h00a2;
  assign func_table_116_imag = 16'h00c5;
  assign func_table_117_real = 16'h0031;
  assign func_table_117_imag = 16'h00fb;
  assign func_table_118_real = 16'hffb6;
  assign func_table_118_imag = 16'h00f4;
  assign func_table_119_real = 16'hff4b;
  assign func_table_119_imag = 16'h00b5;
  assign func_table_120_real = 16'hff0c;
  assign func_table_120_imag = 16'h004a;
  assign func_table_121_real = 16'hff05;
  assign func_table_121_imag = 16'hffcf;
  assign func_table_122_real = 16'hff3b;
  assign func_table_122_imag = 16'hff5e;
  assign func_table_123_real = 16'hff9f;
  assign func_table_123_imag = 16'hff14;
  assign func_table_124_real = 16'h0019;
  assign func_table_124_imag = 16'hff02;
  assign func_table_125_real = 16'h008e;
  assign func_table_125_imag = 16'hff2c;
  assign func_table_126_real = 16'h00e1;
  assign func_table_126_imag = 16'hff88;
  assign func_table_127_real = 16'h0100;
  assign func_table_127_imag = 16'h0;
  assign timeshift_real = _zz_7;
  assign timeshift_imag = _zz_8;
  assign wd_prod = _zz_455[7 : 0];
  assign indx_table_0 = 16'h0;
  assign indx_table_1 = 16'h0200;
  assign indx_table_2 = 16'h0400;
  assign indx_table_3 = 16'h0600;
  assign indx_table_4 = 16'h0800;
  assign indx_table_5 = 16'h0a00;
  assign indx_table_6 = 16'h0c00;
  assign indx_table_7 = 16'h0e00;
  assign indx_table_8 = 16'h1000;
  assign indx_table_9 = 16'h1200;
  assign indx_table_10 = 16'h1400;
  assign indx_table_11 = 16'h1600;
  assign indx_table_12 = 16'h1800;
  assign indx_table_13 = 16'h1a00;
  assign indx_table_14 = 16'h1c00;
  assign indx_table_15 = 16'h1e00;
  assign indx_table_16 = 16'h2000;
  assign indx_table_17 = 16'h2200;
  assign indx_table_18 = 16'h2400;
  assign indx_table_19 = 16'h2600;
  assign indx_table_20 = 16'h2800;
  assign indx_table_21 = 16'h2a00;
  assign indx_table_22 = 16'h2c00;
  assign indx_table_23 = 16'h2e00;
  assign indx_table_24 = 16'h3000;
  assign indx_table_25 = 16'h3200;
  assign indx_table_26 = 16'h3400;
  assign indx_table_27 = 16'h3600;
  assign indx_table_28 = 16'h3800;
  assign indx_table_29 = 16'h3a00;
  assign indx_table_30 = 16'h3c00;
  assign indx_table_31 = 16'h3e00;
  assign indx_table_32 = 16'h4000;
  assign indx_table_33 = 16'h4200;
  assign indx_table_34 = 16'h4400;
  assign indx_table_35 = 16'h4600;
  assign indx_table_36 = 16'h4800;
  assign indx_table_37 = 16'h4a00;
  assign indx_table_38 = 16'h4c00;
  assign indx_table_39 = 16'h4e00;
  assign indx_table_40 = 16'h5000;
  assign indx_table_41 = 16'h5200;
  assign indx_table_42 = 16'h5400;
  assign indx_table_43 = 16'h5600;
  assign indx_table_44 = 16'h5800;
  assign indx_table_45 = 16'h5a00;
  assign indx_table_46 = 16'h5c00;
  assign indx_table_47 = 16'h5e00;
  assign indx_table_48 = 16'h6000;
  assign indx_table_49 = 16'h6200;
  assign indx_table_50 = 16'h6400;
  assign indx_table_51 = 16'h6600;
  assign indx_table_52 = 16'h6800;
  assign indx_table_53 = 16'h6a00;
  assign indx_table_54 = 16'h6c00;
  assign indx_table_55 = 16'h6e00;
  assign indx_table_56 = 16'h7000;
  assign indx_table_57 = 16'h7200;
  assign indx_table_58 = 16'h7400;
  assign indx_table_59 = 16'h7600;
  assign indx_table_60 = 16'h7800;
  assign indx_table_61 = 16'h7a00;
  assign indx_table_62 = 16'h7c00;
  assign indx_table_63 = 16'h7e00;
  assign indx_table_64 = 16'h8000;
  assign indx_table_65 = 16'h8200;
  assign indx_table_66 = 16'h8400;
  assign indx_table_67 = 16'h8600;
  assign indx_table_68 = 16'h8800;
  assign indx_table_69 = 16'h8a00;
  assign indx_table_70 = 16'h8c00;
  assign indx_table_71 = 16'h8e00;
  assign indx_table_72 = 16'h9000;
  assign indx_table_73 = 16'h9200;
  assign indx_table_74 = 16'h9400;
  assign indx_table_75 = 16'h9600;
  assign indx_table_76 = 16'h9800;
  assign indx_table_77 = 16'h9a00;
  assign indx_table_78 = 16'h9c00;
  assign indx_table_79 = 16'h9e00;
  assign indx_table_80 = 16'ha000;
  assign indx_table_81 = 16'ha200;
  assign indx_table_82 = 16'ha400;
  assign indx_table_83 = 16'ha600;
  assign indx_table_84 = 16'ha800;
  assign indx_table_85 = 16'haa00;
  assign indx_table_86 = 16'hac00;
  assign indx_table_87 = 16'hae00;
  assign indx_table_88 = 16'hb000;
  assign indx_table_89 = 16'hb200;
  assign indx_table_90 = 16'hb400;
  assign indx_table_91 = 16'hb600;
  assign indx_table_92 = 16'hb800;
  assign indx_table_93 = 16'hba00;
  assign indx_table_94 = 16'hbc00;
  assign indx_table_95 = 16'hbe00;
  assign indx_table_96 = 16'hc000;
  assign indx_table_97 = 16'hc200;
  assign indx_table_98 = 16'hc400;
  assign indx_table_99 = 16'hc600;
  assign indx_table_100 = 16'hc800;
  assign indx_table_101 = 16'hca00;
  assign indx_table_102 = 16'hcc00;
  assign indx_table_103 = 16'hce00;
  assign indx_table_104 = 16'hd000;
  assign indx_table_105 = 16'hd200;
  assign indx_table_106 = 16'hd400;
  assign indx_table_107 = 16'hd600;
  assign indx_table_108 = 16'hd800;
  assign indx_table_109 = 16'hda00;
  assign indx_table_110 = 16'hdc00;
  assign indx_table_111 = 16'hde00;
  assign indx_table_112 = 16'he000;
  assign indx_table_113 = 16'he200;
  assign indx_table_114 = 16'he400;
  assign indx_table_115 = 16'he600;
  assign indx_table_116 = 16'he800;
  assign indx_table_117 = 16'hea00;
  assign indx_table_118 = 16'hec00;
  assign indx_table_119 = 16'hee00;
  assign indx_table_120 = 16'hf000;
  assign indx_table_121 = 16'hf200;
  assign indx_table_122 = 16'hf400;
  assign indx_table_123 = 16'hf600;
  assign indx_table_124 = 16'hf800;
  assign indx_table_125 = 16'hfa00;
  assign indx_table_126 = 16'hfc00;
  assign indx_table_127 = 16'hfe00;
  assign idx_comp_0 = (_zz_457 < indx_table_0);
  assign idx_comp_1 = (_zz_459 < indx_table_1);
  assign idx_comp_2 = (_zz_461 < indx_table_2);
  assign idx_comp_3 = (_zz_463 < indx_table_3);
  assign idx_comp_4 = (_zz_465 < indx_table_4);
  assign idx_comp_5 = (_zz_467 < indx_table_5);
  assign idx_comp_6 = (_zz_469 < indx_table_6);
  assign idx_comp_7 = (_zz_471 < indx_table_7);
  assign idx_comp_8 = (_zz_473 < indx_table_8);
  assign idx_comp_9 = (_zz_475 < indx_table_9);
  assign idx_comp_10 = (_zz_477 < indx_table_10);
  assign idx_comp_11 = (_zz_479 < indx_table_11);
  assign idx_comp_12 = (_zz_481 < indx_table_12);
  assign idx_comp_13 = (_zz_483 < indx_table_13);
  assign idx_comp_14 = (_zz_485 < indx_table_14);
  assign idx_comp_15 = (_zz_487 < indx_table_15);
  assign idx_comp_16 = (_zz_489 < indx_table_16);
  assign idx_comp_17 = (_zz_491 < indx_table_17);
  assign idx_comp_18 = (_zz_493 < indx_table_18);
  assign idx_comp_19 = (_zz_495 < indx_table_19);
  assign idx_comp_20 = (_zz_497 < indx_table_20);
  assign idx_comp_21 = (_zz_499 < indx_table_21);
  assign idx_comp_22 = (_zz_501 < indx_table_22);
  assign idx_comp_23 = (_zz_503 < indx_table_23);
  assign idx_comp_24 = (_zz_505 < indx_table_24);
  assign idx_comp_25 = (_zz_507 < indx_table_25);
  assign idx_comp_26 = (_zz_509 < indx_table_26);
  assign idx_comp_27 = (_zz_511 < indx_table_27);
  assign idx_comp_28 = (_zz_513 < indx_table_28);
  assign idx_comp_29 = (_zz_515 < indx_table_29);
  assign idx_comp_30 = (_zz_517 < indx_table_30);
  assign idx_comp_31 = (_zz_519 < indx_table_31);
  assign idx_comp_32 = (_zz_521 < indx_table_32);
  assign idx_comp_33 = (_zz_523 < indx_table_33);
  assign idx_comp_34 = (_zz_525 < indx_table_34);
  assign idx_comp_35 = (_zz_527 < indx_table_35);
  assign idx_comp_36 = (_zz_529 < indx_table_36);
  assign idx_comp_37 = (_zz_531 < indx_table_37);
  assign idx_comp_38 = (_zz_533 < indx_table_38);
  assign idx_comp_39 = (_zz_535 < indx_table_39);
  assign idx_comp_40 = (_zz_537 < indx_table_40);
  assign idx_comp_41 = (_zz_539 < indx_table_41);
  assign idx_comp_42 = (_zz_541 < indx_table_42);
  assign idx_comp_43 = (_zz_543 < indx_table_43);
  assign idx_comp_44 = (_zz_545 < indx_table_44);
  assign idx_comp_45 = (_zz_547 < indx_table_45);
  assign idx_comp_46 = (_zz_549 < indx_table_46);
  assign idx_comp_47 = (_zz_551 < indx_table_47);
  assign idx_comp_48 = (_zz_553 < indx_table_48);
  assign idx_comp_49 = (_zz_555 < indx_table_49);
  assign idx_comp_50 = (_zz_557 < indx_table_50);
  assign idx_comp_51 = (_zz_559 < indx_table_51);
  assign idx_comp_52 = (_zz_561 < indx_table_52);
  assign idx_comp_53 = (_zz_563 < indx_table_53);
  assign idx_comp_54 = (_zz_565 < indx_table_54);
  assign idx_comp_55 = (_zz_567 < indx_table_55);
  assign idx_comp_56 = (_zz_569 < indx_table_56);
  assign idx_comp_57 = (_zz_571 < indx_table_57);
  assign idx_comp_58 = (_zz_573 < indx_table_58);
  assign idx_comp_59 = (_zz_575 < indx_table_59);
  assign idx_comp_60 = (_zz_577 < indx_table_60);
  assign idx_comp_61 = (_zz_579 < indx_table_61);
  assign idx_comp_62 = (_zz_581 < indx_table_62);
  assign idx_comp_63 = (_zz_583 < indx_table_63);
  assign idx_comp_64 = (_zz_585 < indx_table_64);
  assign idx_comp_65 = (_zz_587 < indx_table_65);
  assign idx_comp_66 = (_zz_589 < indx_table_66);
  assign idx_comp_67 = (_zz_591 < indx_table_67);
  assign idx_comp_68 = (_zz_593 < indx_table_68);
  assign idx_comp_69 = (_zz_595 < indx_table_69);
  assign idx_comp_70 = (_zz_597 < indx_table_70);
  assign idx_comp_71 = (_zz_599 < indx_table_71);
  assign idx_comp_72 = (_zz_601 < indx_table_72);
  assign idx_comp_73 = (_zz_603 < indx_table_73);
  assign idx_comp_74 = (_zz_605 < indx_table_74);
  assign idx_comp_75 = (_zz_607 < indx_table_75);
  assign idx_comp_76 = (_zz_609 < indx_table_76);
  assign idx_comp_77 = (_zz_611 < indx_table_77);
  assign idx_comp_78 = (_zz_613 < indx_table_78);
  assign idx_comp_79 = (_zz_615 < indx_table_79);
  assign idx_comp_80 = (_zz_617 < indx_table_80);
  assign idx_comp_81 = (_zz_619 < indx_table_81);
  assign idx_comp_82 = (_zz_621 < indx_table_82);
  assign idx_comp_83 = (_zz_623 < indx_table_83);
  assign idx_comp_84 = (_zz_625 < indx_table_84);
  assign idx_comp_85 = (_zz_627 < indx_table_85);
  assign idx_comp_86 = (_zz_629 < indx_table_86);
  assign idx_comp_87 = (_zz_631 < indx_table_87);
  assign idx_comp_88 = (_zz_633 < indx_table_88);
  assign idx_comp_89 = (_zz_635 < indx_table_89);
  assign idx_comp_90 = (_zz_637 < indx_table_90);
  assign idx_comp_91 = (_zz_639 < indx_table_91);
  assign idx_comp_92 = (_zz_641 < indx_table_92);
  assign idx_comp_93 = (_zz_643 < indx_table_93);
  assign idx_comp_94 = (_zz_645 < indx_table_94);
  assign idx_comp_95 = (_zz_647 < indx_table_95);
  assign idx_comp_96 = (_zz_649 < indx_table_96);
  assign idx_comp_97 = (_zz_651 < indx_table_97);
  assign idx_comp_98 = (_zz_653 < indx_table_98);
  assign idx_comp_99 = (_zz_655 < indx_table_99);
  assign idx_comp_100 = (_zz_657 < indx_table_100);
  assign idx_comp_101 = (_zz_659 < indx_table_101);
  assign idx_comp_102 = (_zz_661 < indx_table_102);
  assign idx_comp_103 = (_zz_663 < indx_table_103);
  assign idx_comp_104 = (_zz_665 < indx_table_104);
  assign idx_comp_105 = (_zz_667 < indx_table_105);
  assign idx_comp_106 = (_zz_669 < indx_table_106);
  assign idx_comp_107 = (_zz_671 < indx_table_107);
  assign idx_comp_108 = (_zz_673 < indx_table_108);
  assign idx_comp_109 = (_zz_675 < indx_table_109);
  assign idx_comp_110 = (_zz_677 < indx_table_110);
  assign idx_comp_111 = (_zz_679 < indx_table_111);
  assign idx_comp_112 = (_zz_681 < indx_table_112);
  assign idx_comp_113 = (_zz_683 < indx_table_113);
  assign idx_comp_114 = (_zz_685 < indx_table_114);
  assign idx_comp_115 = (_zz_687 < indx_table_115);
  assign idx_comp_116 = (_zz_689 < indx_table_116);
  assign idx_comp_117 = (_zz_691 < indx_table_117);
  assign idx_comp_118 = (_zz_693 < indx_table_118);
  assign idx_comp_119 = (_zz_695 < indx_table_119);
  assign idx_comp_120 = (_zz_697 < indx_table_120);
  assign idx_comp_121 = (_zz_699 < indx_table_121);
  assign idx_comp_122 = (_zz_701 < indx_table_122);
  assign idx_comp_123 = (_zz_703 < indx_table_123);
  assign idx_comp_124 = (_zz_705 < indx_table_124);
  assign idx_comp_125 = (_zz_707 < indx_table_125);
  assign idx_comp_126 = (_zz_709 < indx_table_126);
  assign idx_comp_127 = (_zz_711 < indx_table_127);
  always @ (*) begin
    _zz_10[0] = idx_comp_0;
    _zz_10[1] = idx_comp_1;
    _zz_10[2] = idx_comp_2;
    _zz_10[3] = idx_comp_3;
    _zz_10[4] = idx_comp_4;
    _zz_10[5] = idx_comp_5;
    _zz_10[6] = idx_comp_6;
    _zz_10[7] = idx_comp_7;
    _zz_10[8] = idx_comp_8;
    _zz_10[9] = idx_comp_9;
    _zz_10[10] = idx_comp_10;
    _zz_10[11] = idx_comp_11;
    _zz_10[12] = idx_comp_12;
    _zz_10[13] = idx_comp_13;
    _zz_10[14] = idx_comp_14;
    _zz_10[15] = idx_comp_15;
    _zz_10[16] = idx_comp_16;
    _zz_10[17] = idx_comp_17;
    _zz_10[18] = idx_comp_18;
    _zz_10[19] = idx_comp_19;
    _zz_10[20] = idx_comp_20;
    _zz_10[21] = idx_comp_21;
    _zz_10[22] = idx_comp_22;
    _zz_10[23] = idx_comp_23;
    _zz_10[24] = idx_comp_24;
    _zz_10[25] = idx_comp_25;
    _zz_10[26] = idx_comp_26;
    _zz_10[27] = idx_comp_27;
    _zz_10[28] = idx_comp_28;
    _zz_10[29] = idx_comp_29;
    _zz_10[30] = idx_comp_30;
    _zz_10[31] = idx_comp_31;
    _zz_10[32] = idx_comp_32;
    _zz_10[33] = idx_comp_33;
    _zz_10[34] = idx_comp_34;
    _zz_10[35] = idx_comp_35;
    _zz_10[36] = idx_comp_36;
    _zz_10[37] = idx_comp_37;
    _zz_10[38] = idx_comp_38;
    _zz_10[39] = idx_comp_39;
    _zz_10[40] = idx_comp_40;
    _zz_10[41] = idx_comp_41;
    _zz_10[42] = idx_comp_42;
    _zz_10[43] = idx_comp_43;
    _zz_10[44] = idx_comp_44;
    _zz_10[45] = idx_comp_45;
    _zz_10[46] = idx_comp_46;
    _zz_10[47] = idx_comp_47;
    _zz_10[48] = idx_comp_48;
    _zz_10[49] = idx_comp_49;
    _zz_10[50] = idx_comp_50;
    _zz_10[51] = idx_comp_51;
    _zz_10[52] = idx_comp_52;
    _zz_10[53] = idx_comp_53;
    _zz_10[54] = idx_comp_54;
    _zz_10[55] = idx_comp_55;
    _zz_10[56] = idx_comp_56;
    _zz_10[57] = idx_comp_57;
    _zz_10[58] = idx_comp_58;
    _zz_10[59] = idx_comp_59;
    _zz_10[60] = idx_comp_60;
    _zz_10[61] = idx_comp_61;
    _zz_10[62] = idx_comp_62;
    _zz_10[63] = idx_comp_63;
    _zz_10[64] = idx_comp_64;
    _zz_10[65] = idx_comp_65;
    _zz_10[66] = idx_comp_66;
    _zz_10[67] = idx_comp_67;
    _zz_10[68] = idx_comp_68;
    _zz_10[69] = idx_comp_69;
    _zz_10[70] = idx_comp_70;
    _zz_10[71] = idx_comp_71;
    _zz_10[72] = idx_comp_72;
    _zz_10[73] = idx_comp_73;
    _zz_10[74] = idx_comp_74;
    _zz_10[75] = idx_comp_75;
    _zz_10[76] = idx_comp_76;
    _zz_10[77] = idx_comp_77;
    _zz_10[78] = idx_comp_78;
    _zz_10[79] = idx_comp_79;
    _zz_10[80] = idx_comp_80;
    _zz_10[81] = idx_comp_81;
    _zz_10[82] = idx_comp_82;
    _zz_10[83] = idx_comp_83;
    _zz_10[84] = idx_comp_84;
    _zz_10[85] = idx_comp_85;
    _zz_10[86] = idx_comp_86;
    _zz_10[87] = idx_comp_87;
    _zz_10[88] = idx_comp_88;
    _zz_10[89] = idx_comp_89;
    _zz_10[90] = idx_comp_90;
    _zz_10[91] = idx_comp_91;
    _zz_10[92] = idx_comp_92;
    _zz_10[93] = idx_comp_93;
    _zz_10[94] = idx_comp_94;
    _zz_10[95] = idx_comp_95;
    _zz_10[96] = idx_comp_96;
    _zz_10[97] = idx_comp_97;
    _zz_10[98] = idx_comp_98;
    _zz_10[99] = idx_comp_99;
    _zz_10[100] = idx_comp_100;
    _zz_10[101] = idx_comp_101;
    _zz_10[102] = idx_comp_102;
    _zz_10[103] = idx_comp_103;
    _zz_10[104] = idx_comp_104;
    _zz_10[105] = idx_comp_105;
    _zz_10[106] = idx_comp_106;
    _zz_10[107] = idx_comp_107;
    _zz_10[108] = idx_comp_108;
    _zz_10[109] = idx_comp_109;
    _zz_10[110] = idx_comp_110;
    _zz_10[111] = idx_comp_111;
    _zz_10[112] = idx_comp_112;
    _zz_10[113] = idx_comp_113;
    _zz_10[114] = idx_comp_114;
    _zz_10[115] = idx_comp_115;
    _zz_10[116] = idx_comp_116;
    _zz_10[117] = idx_comp_117;
    _zz_10[118] = idx_comp_118;
    _zz_10[119] = idx_comp_119;
    _zz_10[120] = idx_comp_120;
    _zz_10[121] = idx_comp_121;
    _zz_10[122] = idx_comp_122;
    _zz_10[123] = idx_comp_123;
    _zz_10[124] = idx_comp_124;
    _zz_10[125] = idx_comp_125;
    _zz_10[126] = idx_comp_126;
    _zz_10[127] = idx_comp_127;
  end

  assign _zz_11 = _zz_10;
  assign all_zeros = ((! (_zz_11 != 128'h0)) ? 8'hff : 8'h0);
  assign all_left_zeros = ((! (_zz_11[127 : 64] != 64'h0)) ? 8'hff : 8'h0);
  assign whole_bit_count = 8'h80;
  assign left_bit_count = 8'h40;
  assign _zz_12 = _zz_11[63 : 0];
  assign all_zeros_1 = ((! (_zz_12 != 64'h0)) ? 7'h7f : 7'h0);
  assign all_left_zeros_1 = ((! (_zz_12[63 : 32] != 32'h0)) ? 7'h7f : 7'h0);
  assign whole_bit_count_1 = 7'h40;
  assign left_bit_count_1 = 7'h20;
  assign _zz_13 = _zz_12[31 : 0];
  assign all_zeros_2 = ((! (_zz_13 != 32'h0)) ? 6'h3f : 6'h0);
  assign all_left_zeros_2 = ((! (_zz_13[31 : 16] != 16'h0)) ? 6'h3f : 6'h0);
  assign whole_bit_count_2 = 6'h20;
  assign left_bit_count_2 = 6'h10;
  assign _zz_14 = _zz_13[15 : 0];
  assign all_zeros_3 = ((! (_zz_14 != 16'h0)) ? 5'h1f : 5'h0);
  assign all_left_zeros_3 = ((! (_zz_14[15 : 8] != 8'h0)) ? 5'h1f : 5'h0);
  assign whole_bit_count_3 = 5'h10;
  assign left_bit_count_3 = 5'h08;
  assign _zz_15 = _zz_14[7 : 0];
  assign all_zeros_4 = ((! (_zz_15 != 8'h0)) ? 4'b1111 : 4'b0000);
  assign all_left_zeros_4 = ((! (_zz_15[7 : 4] != 4'b0000)) ? 4'b1111 : 4'b0000);
  assign whole_bit_count_4 = 4'b1000;
  assign left_bit_count_4 = 4'b0100;
  assign _zz_16 = _zz_15[3 : 0];
  assign all_zeros_5 = ((! (_zz_16 != 4'b0000)) ? 3'b111 : 3'b000);
  assign all_left_zeros_5 = ((! (_zz_16[3 : 2] != 2'b00)) ? 3'b111 : 3'b000);
  assign whole_bit_count_5 = 3'b100;
  assign left_bit_count_5 = 3'b010;
  assign _zz_17 = _zz_16[1 : 0];
  assign all_zeros_6 = ((! (_zz_17 != 2'b00)) ? 2'b11 : 2'b00);
  assign all_left_zeros_6 = ((! (_zz_17[1 : 1] != 1'b0)) ? 2'b11 : 2'b00);
  assign whole_bit_count_6 = 2'b10;
  assign left_bit_count_6 = 2'b01;
  assign _zz_18 = _zz_17[0 : 0];
  assign _zz_19 = _zz_18;
  assign all_zeros_7 = ((! (_zz_19 != 1'b0)) ? 1'b1 : 1'b0);
  assign all_left_zeros_7 = ((! (_zz_19[0 : 0] != 1'b0)) ? 1'b1 : 1'b0);
  assign left_all_zeros_count = (all_left_zeros_6 & _zz_712);
  assign _zz_20 = _zz_17[1 : 1];
  assign _zz_21 = _zz_20;
  assign all_zeros_8 = ((! (_zz_21 != 1'b0)) ? 1'b1 : 1'b0);
  assign all_left_zeros_8 = ((! (_zz_21[0 : 0] != 1'b0)) ? 1'b1 : 1'b0);
  assign left_non_all_zeros_count = ((~ all_left_zeros_6) & _zz_716);
  assign non_zeros_lzc = (left_all_zeros_count + left_non_all_zeros_count);
  assign left_all_zeros_count_1 = (all_left_zeros_5 & _zz_717);
  assign _zz_22 = _zz_16[3 : 2];
  assign all_zeros_9 = ((! (_zz_22 != 2'b00)) ? 2'b11 : 2'b00);
  assign all_left_zeros_9 = ((! (_zz_22[1 : 1] != 1'b0)) ? 2'b11 : 2'b00);
  assign whole_bit_count_7 = 2'b10;
  assign left_bit_count_7 = 2'b01;
  assign _zz_23 = _zz_22[0 : 0];
  assign _zz_24 = _zz_23;
  assign all_zeros_10 = ((! (_zz_24 != 1'b0)) ? 1'b1 : 1'b0);
  assign all_left_zeros_10 = ((! (_zz_24[0 : 0] != 1'b0)) ? 1'b1 : 1'b0);
  assign left_all_zeros_count_2 = (all_left_zeros_9 & _zz_721);
  assign _zz_25 = _zz_22[1 : 1];
  assign _zz_26 = _zz_25;
  assign all_zeros_11 = ((! (_zz_26 != 1'b0)) ? 1'b1 : 1'b0);
  assign all_left_zeros_11 = ((! (_zz_26[0 : 0] != 1'b0)) ? 1'b1 : 1'b0);
  assign left_non_all_zeros_count_1 = ((~ all_left_zeros_9) & _zz_725);
  assign non_zeros_lzc_1 = (left_all_zeros_count_2 + left_non_all_zeros_count_1);
  assign left_non_all_zeros_count_2 = ((~ all_left_zeros_5) & _zz_727);
  assign non_zeros_lzc_2 = (left_all_zeros_count_1 + left_non_all_zeros_count_2);
  assign left_all_zeros_count_3 = (all_left_zeros_4 & _zz_729);
  assign _zz_27 = _zz_15[7 : 4];
  assign all_zeros_12 = ((! (_zz_27 != 4'b0000)) ? 3'b111 : 3'b000);
  assign all_left_zeros_12 = ((! (_zz_27[3 : 2] != 2'b00)) ? 3'b111 : 3'b000);
  assign whole_bit_count_8 = 3'b100;
  assign left_bit_count_8 = 3'b010;
  assign _zz_28 = _zz_27[1 : 0];
  assign all_zeros_13 = ((! (_zz_28 != 2'b00)) ? 2'b11 : 2'b00);
  assign all_left_zeros_13 = ((! (_zz_28[1 : 1] != 1'b0)) ? 2'b11 : 2'b00);
  assign whole_bit_count_9 = 2'b10;
  assign left_bit_count_9 = 2'b01;
  assign _zz_29 = _zz_28[0 : 0];
  assign _zz_30 = _zz_29;
  assign all_zeros_14 = ((! (_zz_30 != 1'b0)) ? 1'b1 : 1'b0);
  assign all_left_zeros_14 = ((! (_zz_30[0 : 0] != 1'b0)) ? 1'b1 : 1'b0);
  assign left_all_zeros_count_4 = (all_left_zeros_13 & _zz_733);
  assign _zz_31 = _zz_28[1 : 1];
  assign _zz_32 = _zz_31;
  assign all_zeros_15 = ((! (_zz_32 != 1'b0)) ? 1'b1 : 1'b0);
  assign all_left_zeros_15 = ((! (_zz_32[0 : 0] != 1'b0)) ? 1'b1 : 1'b0);
  assign left_non_all_zeros_count_3 = ((~ all_left_zeros_13) & _zz_737);
  assign non_zeros_lzc_3 = (left_all_zeros_count_4 + left_non_all_zeros_count_3);
  assign left_all_zeros_count_5 = (all_left_zeros_12 & _zz_738);
  assign _zz_33 = _zz_27[3 : 2];
  assign all_zeros_16 = ((! (_zz_33 != 2'b00)) ? 2'b11 : 2'b00);
  assign all_left_zeros_16 = ((! (_zz_33[1 : 1] != 1'b0)) ? 2'b11 : 2'b00);
  assign whole_bit_count_10 = 2'b10;
  assign left_bit_count_10 = 2'b01;
  assign _zz_34 = _zz_33[0 : 0];
  assign _zz_35 = _zz_34;
  assign all_zeros_17 = ((! (_zz_35 != 1'b0)) ? 1'b1 : 1'b0);
  assign all_left_zeros_17 = ((! (_zz_35[0 : 0] != 1'b0)) ? 1'b1 : 1'b0);
  assign left_all_zeros_count_6 = (all_left_zeros_16 & _zz_742);
  assign _zz_36 = _zz_33[1 : 1];
  assign _zz_37 = _zz_36;
  assign all_zeros_18 = ((! (_zz_37 != 1'b0)) ? 1'b1 : 1'b0);
  assign all_left_zeros_18 = ((! (_zz_37[0 : 0] != 1'b0)) ? 1'b1 : 1'b0);
  assign left_non_all_zeros_count_4 = ((~ all_left_zeros_16) & _zz_746);
  assign non_zeros_lzc_4 = (left_all_zeros_count_6 + left_non_all_zeros_count_4);
  assign left_non_all_zeros_count_5 = ((~ all_left_zeros_12) & _zz_748);
  assign non_zeros_lzc_5 = (left_all_zeros_count_5 + left_non_all_zeros_count_5);
  assign left_non_all_zeros_count_6 = ((~ all_left_zeros_4) & _zz_751);
  assign non_zeros_lzc_6 = (left_all_zeros_count_3 + left_non_all_zeros_count_6);
  assign left_all_zeros_count_7 = (all_left_zeros_3 & _zz_753);
  assign _zz_38 = _zz_14[15 : 8];
  assign all_zeros_19 = ((! (_zz_38 != 8'h0)) ? 4'b1111 : 4'b0000);
  assign all_left_zeros_19 = ((! (_zz_38[7 : 4] != 4'b0000)) ? 4'b1111 : 4'b0000);
  assign whole_bit_count_11 = 4'b1000;
  assign left_bit_count_11 = 4'b0100;
  assign _zz_39 = _zz_38[3 : 0];
  assign all_zeros_20 = ((! (_zz_39 != 4'b0000)) ? 3'b111 : 3'b000);
  assign all_left_zeros_20 = ((! (_zz_39[3 : 2] != 2'b00)) ? 3'b111 : 3'b000);
  assign whole_bit_count_12 = 3'b100;
  assign left_bit_count_12 = 3'b010;
  assign _zz_40 = _zz_39[1 : 0];
  assign all_zeros_21 = ((! (_zz_40 != 2'b00)) ? 2'b11 : 2'b00);
  assign all_left_zeros_21 = ((! (_zz_40[1 : 1] != 1'b0)) ? 2'b11 : 2'b00);
  assign whole_bit_count_13 = 2'b10;
  assign left_bit_count_13 = 2'b01;
  assign _zz_41 = _zz_40[0 : 0];
  assign _zz_42 = _zz_41;
  assign all_zeros_22 = ((! (_zz_42 != 1'b0)) ? 1'b1 : 1'b0);
  assign all_left_zeros_22 = ((! (_zz_42[0 : 0] != 1'b0)) ? 1'b1 : 1'b0);
  assign left_all_zeros_count_8 = (all_left_zeros_21 & _zz_757);
  assign _zz_43 = _zz_40[1 : 1];
  assign _zz_44 = _zz_43;
  assign all_zeros_23 = ((! (_zz_44 != 1'b0)) ? 1'b1 : 1'b0);
  assign all_left_zeros_23 = ((! (_zz_44[0 : 0] != 1'b0)) ? 1'b1 : 1'b0);
  assign left_non_all_zeros_count_7 = ((~ all_left_zeros_21) & _zz_761);
  assign non_zeros_lzc_7 = (left_all_zeros_count_8 + left_non_all_zeros_count_7);
  assign left_all_zeros_count_9 = (all_left_zeros_20 & _zz_762);
  assign _zz_45 = _zz_39[3 : 2];
  assign all_zeros_24 = ((! (_zz_45 != 2'b00)) ? 2'b11 : 2'b00);
  assign all_left_zeros_24 = ((! (_zz_45[1 : 1] != 1'b0)) ? 2'b11 : 2'b00);
  assign whole_bit_count_14 = 2'b10;
  assign left_bit_count_14 = 2'b01;
  assign _zz_46 = _zz_45[0 : 0];
  assign _zz_47 = _zz_46;
  assign all_zeros_25 = ((! (_zz_47 != 1'b0)) ? 1'b1 : 1'b0);
  assign all_left_zeros_25 = ((! (_zz_47[0 : 0] != 1'b0)) ? 1'b1 : 1'b0);
  assign left_all_zeros_count_10 = (all_left_zeros_24 & _zz_766);
  assign _zz_48 = _zz_45[1 : 1];
  assign _zz_49 = _zz_48;
  assign all_zeros_26 = ((! (_zz_49 != 1'b0)) ? 1'b1 : 1'b0);
  assign all_left_zeros_26 = ((! (_zz_49[0 : 0] != 1'b0)) ? 1'b1 : 1'b0);
  assign left_non_all_zeros_count_8 = ((~ all_left_zeros_24) & _zz_770);
  assign non_zeros_lzc_8 = (left_all_zeros_count_10 + left_non_all_zeros_count_8);
  assign left_non_all_zeros_count_9 = ((~ all_left_zeros_20) & _zz_772);
  assign non_zeros_lzc_9 = (left_all_zeros_count_9 + left_non_all_zeros_count_9);
  assign left_all_zeros_count_11 = (all_left_zeros_19 & _zz_774);
  assign _zz_50 = _zz_38[7 : 4];
  assign all_zeros_27 = ((! (_zz_50 != 4'b0000)) ? 3'b111 : 3'b000);
  assign all_left_zeros_27 = ((! (_zz_50[3 : 2] != 2'b00)) ? 3'b111 : 3'b000);
  assign whole_bit_count_15 = 3'b100;
  assign left_bit_count_15 = 3'b010;
  assign _zz_51 = _zz_50[1 : 0];
  assign all_zeros_28 = ((! (_zz_51 != 2'b00)) ? 2'b11 : 2'b00);
  assign all_left_zeros_28 = ((! (_zz_51[1 : 1] != 1'b0)) ? 2'b11 : 2'b00);
  assign whole_bit_count_16 = 2'b10;
  assign left_bit_count_16 = 2'b01;
  assign _zz_52 = _zz_51[0 : 0];
  assign _zz_53 = _zz_52;
  assign all_zeros_29 = ((! (_zz_53 != 1'b0)) ? 1'b1 : 1'b0);
  assign all_left_zeros_29 = ((! (_zz_53[0 : 0] != 1'b0)) ? 1'b1 : 1'b0);
  assign left_all_zeros_count_12 = (all_left_zeros_28 & _zz_778);
  assign _zz_54 = _zz_51[1 : 1];
  assign _zz_55 = _zz_54;
  assign all_zeros_30 = ((! (_zz_55 != 1'b0)) ? 1'b1 : 1'b0);
  assign all_left_zeros_30 = ((! (_zz_55[0 : 0] != 1'b0)) ? 1'b1 : 1'b0);
  assign left_non_all_zeros_count_10 = ((~ all_left_zeros_28) & _zz_782);
  assign non_zeros_lzc_10 = (left_all_zeros_count_12 + left_non_all_zeros_count_10);
  assign left_all_zeros_count_13 = (all_left_zeros_27 & _zz_783);
  assign _zz_56 = _zz_50[3 : 2];
  assign all_zeros_31 = ((! (_zz_56 != 2'b00)) ? 2'b11 : 2'b00);
  assign all_left_zeros_31 = ((! (_zz_56[1 : 1] != 1'b0)) ? 2'b11 : 2'b00);
  assign whole_bit_count_17 = 2'b10;
  assign left_bit_count_17 = 2'b01;
  assign _zz_57 = _zz_56[0 : 0];
  assign _zz_58 = _zz_57;
  assign all_zeros_32 = ((! (_zz_58 != 1'b0)) ? 1'b1 : 1'b0);
  assign all_left_zeros_32 = ((! (_zz_58[0 : 0] != 1'b0)) ? 1'b1 : 1'b0);
  assign left_all_zeros_count_14 = (all_left_zeros_31 & _zz_787);
  assign _zz_59 = _zz_56[1 : 1];
  assign _zz_60 = _zz_59;
  assign all_zeros_33 = ((! (_zz_60 != 1'b0)) ? 1'b1 : 1'b0);
  assign all_left_zeros_33 = ((! (_zz_60[0 : 0] != 1'b0)) ? 1'b1 : 1'b0);
  assign left_non_all_zeros_count_11 = ((~ all_left_zeros_31) & _zz_791);
  assign non_zeros_lzc_11 = (left_all_zeros_count_14 + left_non_all_zeros_count_11);
  assign left_non_all_zeros_count_12 = ((~ all_left_zeros_27) & _zz_793);
  assign non_zeros_lzc_12 = (left_all_zeros_count_13 + left_non_all_zeros_count_12);
  assign left_non_all_zeros_count_13 = ((~ all_left_zeros_19) & _zz_796);
  assign non_zeros_lzc_13 = (left_all_zeros_count_11 + left_non_all_zeros_count_13);
  assign left_non_all_zeros_count_14 = ((~ all_left_zeros_3) & _zz_799);
  assign non_zeros_lzc_14 = (left_all_zeros_count_7 + left_non_all_zeros_count_14);
  assign left_all_zeros_count_15 = (all_left_zeros_2 & _zz_801);
  assign _zz_61 = _zz_13[31 : 16];
  assign all_zeros_34 = ((! (_zz_61 != 16'h0)) ? 5'h1f : 5'h0);
  assign all_left_zeros_34 = ((! (_zz_61[15 : 8] != 8'h0)) ? 5'h1f : 5'h0);
  assign whole_bit_count_18 = 5'h10;
  assign left_bit_count_18 = 5'h08;
  assign _zz_62 = _zz_61[7 : 0];
  assign all_zeros_35 = ((! (_zz_62 != 8'h0)) ? 4'b1111 : 4'b0000);
  assign all_left_zeros_35 = ((! (_zz_62[7 : 4] != 4'b0000)) ? 4'b1111 : 4'b0000);
  assign whole_bit_count_19 = 4'b1000;
  assign left_bit_count_19 = 4'b0100;
  assign _zz_63 = _zz_62[3 : 0];
  assign all_zeros_36 = ((! (_zz_63 != 4'b0000)) ? 3'b111 : 3'b000);
  assign all_left_zeros_36 = ((! (_zz_63[3 : 2] != 2'b00)) ? 3'b111 : 3'b000);
  assign whole_bit_count_20 = 3'b100;
  assign left_bit_count_20 = 3'b010;
  assign _zz_64 = _zz_63[1 : 0];
  assign all_zeros_37 = ((! (_zz_64 != 2'b00)) ? 2'b11 : 2'b00);
  assign all_left_zeros_37 = ((! (_zz_64[1 : 1] != 1'b0)) ? 2'b11 : 2'b00);
  assign whole_bit_count_21 = 2'b10;
  assign left_bit_count_21 = 2'b01;
  assign _zz_65 = _zz_64[0 : 0];
  assign _zz_66 = _zz_65;
  assign all_zeros_38 = ((! (_zz_66 != 1'b0)) ? 1'b1 : 1'b0);
  assign all_left_zeros_38 = ((! (_zz_66[0 : 0] != 1'b0)) ? 1'b1 : 1'b0);
  assign left_all_zeros_count_16 = (all_left_zeros_37 & _zz_805);
  assign _zz_67 = _zz_64[1 : 1];
  assign _zz_68 = _zz_67;
  assign all_zeros_39 = ((! (_zz_68 != 1'b0)) ? 1'b1 : 1'b0);
  assign all_left_zeros_39 = ((! (_zz_68[0 : 0] != 1'b0)) ? 1'b1 : 1'b0);
  assign left_non_all_zeros_count_15 = ((~ all_left_zeros_37) & _zz_809);
  assign non_zeros_lzc_15 = (left_all_zeros_count_16 + left_non_all_zeros_count_15);
  assign left_all_zeros_count_17 = (all_left_zeros_36 & _zz_810);
  assign _zz_69 = _zz_63[3 : 2];
  assign all_zeros_40 = ((! (_zz_69 != 2'b00)) ? 2'b11 : 2'b00);
  assign all_left_zeros_40 = ((! (_zz_69[1 : 1] != 1'b0)) ? 2'b11 : 2'b00);
  assign whole_bit_count_22 = 2'b10;
  assign left_bit_count_22 = 2'b01;
  assign _zz_70 = _zz_69[0 : 0];
  assign _zz_71 = _zz_70;
  assign all_zeros_41 = ((! (_zz_71 != 1'b0)) ? 1'b1 : 1'b0);
  assign all_left_zeros_41 = ((! (_zz_71[0 : 0] != 1'b0)) ? 1'b1 : 1'b0);
  assign left_all_zeros_count_18 = (all_left_zeros_40 & _zz_814);
  assign _zz_72 = _zz_69[1 : 1];
  assign _zz_73 = _zz_72;
  assign all_zeros_42 = ((! (_zz_73 != 1'b0)) ? 1'b1 : 1'b0);
  assign all_left_zeros_42 = ((! (_zz_73[0 : 0] != 1'b0)) ? 1'b1 : 1'b0);
  assign left_non_all_zeros_count_16 = ((~ all_left_zeros_40) & _zz_818);
  assign non_zeros_lzc_16 = (left_all_zeros_count_18 + left_non_all_zeros_count_16);
  assign left_non_all_zeros_count_17 = ((~ all_left_zeros_36) & _zz_820);
  assign non_zeros_lzc_17 = (left_all_zeros_count_17 + left_non_all_zeros_count_17);
  assign left_all_zeros_count_19 = (all_left_zeros_35 & _zz_822);
  assign _zz_74 = _zz_62[7 : 4];
  assign all_zeros_43 = ((! (_zz_74 != 4'b0000)) ? 3'b111 : 3'b000);
  assign all_left_zeros_43 = ((! (_zz_74[3 : 2] != 2'b00)) ? 3'b111 : 3'b000);
  assign whole_bit_count_23 = 3'b100;
  assign left_bit_count_23 = 3'b010;
  assign _zz_75 = _zz_74[1 : 0];
  assign all_zeros_44 = ((! (_zz_75 != 2'b00)) ? 2'b11 : 2'b00);
  assign all_left_zeros_44 = ((! (_zz_75[1 : 1] != 1'b0)) ? 2'b11 : 2'b00);
  assign whole_bit_count_24 = 2'b10;
  assign left_bit_count_24 = 2'b01;
  assign _zz_76 = _zz_75[0 : 0];
  assign _zz_77 = _zz_76;
  assign all_zeros_45 = ((! (_zz_77 != 1'b0)) ? 1'b1 : 1'b0);
  assign all_left_zeros_45 = ((! (_zz_77[0 : 0] != 1'b0)) ? 1'b1 : 1'b0);
  assign left_all_zeros_count_20 = (all_left_zeros_44 & _zz_826);
  assign _zz_78 = _zz_75[1 : 1];
  assign _zz_79 = _zz_78;
  assign all_zeros_46 = ((! (_zz_79 != 1'b0)) ? 1'b1 : 1'b0);
  assign all_left_zeros_46 = ((! (_zz_79[0 : 0] != 1'b0)) ? 1'b1 : 1'b0);
  assign left_non_all_zeros_count_18 = ((~ all_left_zeros_44) & _zz_830);
  assign non_zeros_lzc_18 = (left_all_zeros_count_20 + left_non_all_zeros_count_18);
  assign left_all_zeros_count_21 = (all_left_zeros_43 & _zz_831);
  assign _zz_80 = _zz_74[3 : 2];
  assign all_zeros_47 = ((! (_zz_80 != 2'b00)) ? 2'b11 : 2'b00);
  assign all_left_zeros_47 = ((! (_zz_80[1 : 1] != 1'b0)) ? 2'b11 : 2'b00);
  assign whole_bit_count_25 = 2'b10;
  assign left_bit_count_25 = 2'b01;
  assign _zz_81 = _zz_80[0 : 0];
  assign _zz_82 = _zz_81;
  assign all_zeros_48 = ((! (_zz_82 != 1'b0)) ? 1'b1 : 1'b0);
  assign all_left_zeros_48 = ((! (_zz_82[0 : 0] != 1'b0)) ? 1'b1 : 1'b0);
  assign left_all_zeros_count_22 = (all_left_zeros_47 & _zz_835);
  assign _zz_83 = _zz_80[1 : 1];
  assign _zz_84 = _zz_83;
  assign all_zeros_49 = ((! (_zz_84 != 1'b0)) ? 1'b1 : 1'b0);
  assign all_left_zeros_49 = ((! (_zz_84[0 : 0] != 1'b0)) ? 1'b1 : 1'b0);
  assign left_non_all_zeros_count_19 = ((~ all_left_zeros_47) & _zz_839);
  assign non_zeros_lzc_19 = (left_all_zeros_count_22 + left_non_all_zeros_count_19);
  assign left_non_all_zeros_count_20 = ((~ all_left_zeros_43) & _zz_841);
  assign non_zeros_lzc_20 = (left_all_zeros_count_21 + left_non_all_zeros_count_20);
  assign left_non_all_zeros_count_21 = ((~ all_left_zeros_35) & _zz_844);
  assign non_zeros_lzc_21 = (left_all_zeros_count_19 + left_non_all_zeros_count_21);
  assign left_all_zeros_count_23 = (all_left_zeros_34 & _zz_846);
  assign _zz_85 = _zz_61[15 : 8];
  assign all_zeros_50 = ((! (_zz_85 != 8'h0)) ? 4'b1111 : 4'b0000);
  assign all_left_zeros_50 = ((! (_zz_85[7 : 4] != 4'b0000)) ? 4'b1111 : 4'b0000);
  assign whole_bit_count_26 = 4'b1000;
  assign left_bit_count_26 = 4'b0100;
  assign _zz_86 = _zz_85[3 : 0];
  assign all_zeros_51 = ((! (_zz_86 != 4'b0000)) ? 3'b111 : 3'b000);
  assign all_left_zeros_51 = ((! (_zz_86[3 : 2] != 2'b00)) ? 3'b111 : 3'b000);
  assign whole_bit_count_27 = 3'b100;
  assign left_bit_count_27 = 3'b010;
  assign _zz_87 = _zz_86[1 : 0];
  assign all_zeros_52 = ((! (_zz_87 != 2'b00)) ? 2'b11 : 2'b00);
  assign all_left_zeros_52 = ((! (_zz_87[1 : 1] != 1'b0)) ? 2'b11 : 2'b00);
  assign whole_bit_count_28 = 2'b10;
  assign left_bit_count_28 = 2'b01;
  assign _zz_88 = _zz_87[0 : 0];
  assign _zz_89 = _zz_88;
  assign all_zeros_53 = ((! (_zz_89 != 1'b0)) ? 1'b1 : 1'b0);
  assign all_left_zeros_53 = ((! (_zz_89[0 : 0] != 1'b0)) ? 1'b1 : 1'b0);
  assign left_all_zeros_count_24 = (all_left_zeros_52 & _zz_850);
  assign _zz_90 = _zz_87[1 : 1];
  assign _zz_91 = _zz_90;
  assign all_zeros_54 = ((! (_zz_91 != 1'b0)) ? 1'b1 : 1'b0);
  assign all_left_zeros_54 = ((! (_zz_91[0 : 0] != 1'b0)) ? 1'b1 : 1'b0);
  assign left_non_all_zeros_count_22 = ((~ all_left_zeros_52) & _zz_854);
  assign non_zeros_lzc_22 = (left_all_zeros_count_24 + left_non_all_zeros_count_22);
  assign left_all_zeros_count_25 = (all_left_zeros_51 & _zz_855);
  assign _zz_92 = _zz_86[3 : 2];
  assign all_zeros_55 = ((! (_zz_92 != 2'b00)) ? 2'b11 : 2'b00);
  assign all_left_zeros_55 = ((! (_zz_92[1 : 1] != 1'b0)) ? 2'b11 : 2'b00);
  assign whole_bit_count_29 = 2'b10;
  assign left_bit_count_29 = 2'b01;
  assign _zz_93 = _zz_92[0 : 0];
  assign _zz_94 = _zz_93;
  assign all_zeros_56 = ((! (_zz_94 != 1'b0)) ? 1'b1 : 1'b0);
  assign all_left_zeros_56 = ((! (_zz_94[0 : 0] != 1'b0)) ? 1'b1 : 1'b0);
  assign left_all_zeros_count_26 = (all_left_zeros_55 & _zz_859);
  assign _zz_95 = _zz_92[1 : 1];
  assign _zz_96 = _zz_95;
  assign all_zeros_57 = ((! (_zz_96 != 1'b0)) ? 1'b1 : 1'b0);
  assign all_left_zeros_57 = ((! (_zz_96[0 : 0] != 1'b0)) ? 1'b1 : 1'b0);
  assign left_non_all_zeros_count_23 = ((~ all_left_zeros_55) & _zz_863);
  assign non_zeros_lzc_23 = (left_all_zeros_count_26 + left_non_all_zeros_count_23);
  assign left_non_all_zeros_count_24 = ((~ all_left_zeros_51) & _zz_865);
  assign non_zeros_lzc_24 = (left_all_zeros_count_25 + left_non_all_zeros_count_24);
  assign left_all_zeros_count_27 = (all_left_zeros_50 & _zz_867);
  assign _zz_97 = _zz_85[7 : 4];
  assign all_zeros_58 = ((! (_zz_97 != 4'b0000)) ? 3'b111 : 3'b000);
  assign all_left_zeros_58 = ((! (_zz_97[3 : 2] != 2'b00)) ? 3'b111 : 3'b000);
  assign whole_bit_count_30 = 3'b100;
  assign left_bit_count_30 = 3'b010;
  assign _zz_98 = _zz_97[1 : 0];
  assign all_zeros_59 = ((! (_zz_98 != 2'b00)) ? 2'b11 : 2'b00);
  assign all_left_zeros_59 = ((! (_zz_98[1 : 1] != 1'b0)) ? 2'b11 : 2'b00);
  assign whole_bit_count_31 = 2'b10;
  assign left_bit_count_31 = 2'b01;
  assign _zz_99 = _zz_98[0 : 0];
  assign _zz_100 = _zz_99;
  assign all_zeros_60 = ((! (_zz_100 != 1'b0)) ? 1'b1 : 1'b0);
  assign all_left_zeros_60 = ((! (_zz_100[0 : 0] != 1'b0)) ? 1'b1 : 1'b0);
  assign left_all_zeros_count_28 = (all_left_zeros_59 & _zz_871);
  assign _zz_101 = _zz_98[1 : 1];
  assign _zz_102 = _zz_101;
  assign all_zeros_61 = ((! (_zz_102 != 1'b0)) ? 1'b1 : 1'b0);
  assign all_left_zeros_61 = ((! (_zz_102[0 : 0] != 1'b0)) ? 1'b1 : 1'b0);
  assign left_non_all_zeros_count_25 = ((~ all_left_zeros_59) & _zz_875);
  assign non_zeros_lzc_25 = (left_all_zeros_count_28 + left_non_all_zeros_count_25);
  assign left_all_zeros_count_29 = (all_left_zeros_58 & _zz_876);
  assign _zz_103 = _zz_97[3 : 2];
  assign all_zeros_62 = ((! (_zz_103 != 2'b00)) ? 2'b11 : 2'b00);
  assign all_left_zeros_62 = ((! (_zz_103[1 : 1] != 1'b0)) ? 2'b11 : 2'b00);
  assign whole_bit_count_32 = 2'b10;
  assign left_bit_count_32 = 2'b01;
  assign _zz_104 = _zz_103[0 : 0];
  assign _zz_105 = _zz_104;
  assign all_zeros_63 = ((! (_zz_105 != 1'b0)) ? 1'b1 : 1'b0);
  assign all_left_zeros_63 = ((! (_zz_105[0 : 0] != 1'b0)) ? 1'b1 : 1'b0);
  assign left_all_zeros_count_30 = (all_left_zeros_62 & _zz_880);
  assign _zz_106 = _zz_103[1 : 1];
  assign _zz_107 = _zz_106;
  assign all_zeros_64 = ((! (_zz_107 != 1'b0)) ? 1'b1 : 1'b0);
  assign all_left_zeros_64 = ((! (_zz_107[0 : 0] != 1'b0)) ? 1'b1 : 1'b0);
  assign left_non_all_zeros_count_26 = ((~ all_left_zeros_62) & _zz_884);
  assign non_zeros_lzc_26 = (left_all_zeros_count_30 + left_non_all_zeros_count_26);
  assign left_non_all_zeros_count_27 = ((~ all_left_zeros_58) & _zz_886);
  assign non_zeros_lzc_27 = (left_all_zeros_count_29 + left_non_all_zeros_count_27);
  assign left_non_all_zeros_count_28 = ((~ all_left_zeros_50) & _zz_889);
  assign non_zeros_lzc_28 = (left_all_zeros_count_27 + left_non_all_zeros_count_28);
  assign left_non_all_zeros_count_29 = ((~ all_left_zeros_34) & _zz_892);
  assign non_zeros_lzc_29 = (left_all_zeros_count_23 + left_non_all_zeros_count_29);
  assign left_non_all_zeros_count_30 = ((~ all_left_zeros_2) & _zz_895);
  assign non_zeros_lzc_30 = (left_all_zeros_count_15 + left_non_all_zeros_count_30);
  assign left_all_zeros_count_31 = (all_left_zeros_1 & _zz_897);
  assign _zz_108 = _zz_12[63 : 32];
  assign all_zeros_65 = ((! (_zz_108 != 32'h0)) ? 6'h3f : 6'h0);
  assign all_left_zeros_65 = ((! (_zz_108[31 : 16] != 16'h0)) ? 6'h3f : 6'h0);
  assign whole_bit_count_33 = 6'h20;
  assign left_bit_count_33 = 6'h10;
  assign _zz_109 = _zz_108[15 : 0];
  assign all_zeros_66 = ((! (_zz_109 != 16'h0)) ? 5'h1f : 5'h0);
  assign all_left_zeros_66 = ((! (_zz_109[15 : 8] != 8'h0)) ? 5'h1f : 5'h0);
  assign whole_bit_count_34 = 5'h10;
  assign left_bit_count_34 = 5'h08;
  assign _zz_110 = _zz_109[7 : 0];
  assign all_zeros_67 = ((! (_zz_110 != 8'h0)) ? 4'b1111 : 4'b0000);
  assign all_left_zeros_67 = ((! (_zz_110[7 : 4] != 4'b0000)) ? 4'b1111 : 4'b0000);
  assign whole_bit_count_35 = 4'b1000;
  assign left_bit_count_35 = 4'b0100;
  assign _zz_111 = _zz_110[3 : 0];
  assign all_zeros_68 = ((! (_zz_111 != 4'b0000)) ? 3'b111 : 3'b000);
  assign all_left_zeros_68 = ((! (_zz_111[3 : 2] != 2'b00)) ? 3'b111 : 3'b000);
  assign whole_bit_count_36 = 3'b100;
  assign left_bit_count_36 = 3'b010;
  assign _zz_112 = _zz_111[1 : 0];
  assign all_zeros_69 = ((! (_zz_112 != 2'b00)) ? 2'b11 : 2'b00);
  assign all_left_zeros_69 = ((! (_zz_112[1 : 1] != 1'b0)) ? 2'b11 : 2'b00);
  assign whole_bit_count_37 = 2'b10;
  assign left_bit_count_37 = 2'b01;
  assign _zz_113 = _zz_112[0 : 0];
  assign _zz_114 = _zz_113;
  assign all_zeros_70 = ((! (_zz_114 != 1'b0)) ? 1'b1 : 1'b0);
  assign all_left_zeros_70 = ((! (_zz_114[0 : 0] != 1'b0)) ? 1'b1 : 1'b0);
  assign left_all_zeros_count_32 = (all_left_zeros_69 & _zz_901);
  assign _zz_115 = _zz_112[1 : 1];
  assign _zz_116 = _zz_115;
  assign all_zeros_71 = ((! (_zz_116 != 1'b0)) ? 1'b1 : 1'b0);
  assign all_left_zeros_71 = ((! (_zz_116[0 : 0] != 1'b0)) ? 1'b1 : 1'b0);
  assign left_non_all_zeros_count_31 = ((~ all_left_zeros_69) & _zz_905);
  assign non_zeros_lzc_31 = (left_all_zeros_count_32 + left_non_all_zeros_count_31);
  assign left_all_zeros_count_33 = (all_left_zeros_68 & _zz_906);
  assign _zz_117 = _zz_111[3 : 2];
  assign all_zeros_72 = ((! (_zz_117 != 2'b00)) ? 2'b11 : 2'b00);
  assign all_left_zeros_72 = ((! (_zz_117[1 : 1] != 1'b0)) ? 2'b11 : 2'b00);
  assign whole_bit_count_38 = 2'b10;
  assign left_bit_count_38 = 2'b01;
  assign _zz_118 = _zz_117[0 : 0];
  assign _zz_119 = _zz_118;
  assign all_zeros_73 = ((! (_zz_119 != 1'b0)) ? 1'b1 : 1'b0);
  assign all_left_zeros_73 = ((! (_zz_119[0 : 0] != 1'b0)) ? 1'b1 : 1'b0);
  assign left_all_zeros_count_34 = (all_left_zeros_72 & _zz_910);
  assign _zz_120 = _zz_117[1 : 1];
  assign _zz_121 = _zz_120;
  assign all_zeros_74 = ((! (_zz_121 != 1'b0)) ? 1'b1 : 1'b0);
  assign all_left_zeros_74 = ((! (_zz_121[0 : 0] != 1'b0)) ? 1'b1 : 1'b0);
  assign left_non_all_zeros_count_32 = ((~ all_left_zeros_72) & _zz_914);
  assign non_zeros_lzc_32 = (left_all_zeros_count_34 + left_non_all_zeros_count_32);
  assign left_non_all_zeros_count_33 = ((~ all_left_zeros_68) & _zz_916);
  assign non_zeros_lzc_33 = (left_all_zeros_count_33 + left_non_all_zeros_count_33);
  assign left_all_zeros_count_35 = (all_left_zeros_67 & _zz_918);
  assign _zz_122 = _zz_110[7 : 4];
  assign all_zeros_75 = ((! (_zz_122 != 4'b0000)) ? 3'b111 : 3'b000);
  assign all_left_zeros_75 = ((! (_zz_122[3 : 2] != 2'b00)) ? 3'b111 : 3'b000);
  assign whole_bit_count_39 = 3'b100;
  assign left_bit_count_39 = 3'b010;
  assign _zz_123 = _zz_122[1 : 0];
  assign all_zeros_76 = ((! (_zz_123 != 2'b00)) ? 2'b11 : 2'b00);
  assign all_left_zeros_76 = ((! (_zz_123[1 : 1] != 1'b0)) ? 2'b11 : 2'b00);
  assign whole_bit_count_40 = 2'b10;
  assign left_bit_count_40 = 2'b01;
  assign _zz_124 = _zz_123[0 : 0];
  assign _zz_125 = _zz_124;
  assign all_zeros_77 = ((! (_zz_125 != 1'b0)) ? 1'b1 : 1'b0);
  assign all_left_zeros_77 = ((! (_zz_125[0 : 0] != 1'b0)) ? 1'b1 : 1'b0);
  assign left_all_zeros_count_36 = (all_left_zeros_76 & _zz_922);
  assign _zz_126 = _zz_123[1 : 1];
  assign _zz_127 = _zz_126;
  assign all_zeros_78 = ((! (_zz_127 != 1'b0)) ? 1'b1 : 1'b0);
  assign all_left_zeros_78 = ((! (_zz_127[0 : 0] != 1'b0)) ? 1'b1 : 1'b0);
  assign left_non_all_zeros_count_34 = ((~ all_left_zeros_76) & _zz_926);
  assign non_zeros_lzc_34 = (left_all_zeros_count_36 + left_non_all_zeros_count_34);
  assign left_all_zeros_count_37 = (all_left_zeros_75 & _zz_927);
  assign _zz_128 = _zz_122[3 : 2];
  assign all_zeros_79 = ((! (_zz_128 != 2'b00)) ? 2'b11 : 2'b00);
  assign all_left_zeros_79 = ((! (_zz_128[1 : 1] != 1'b0)) ? 2'b11 : 2'b00);
  assign whole_bit_count_41 = 2'b10;
  assign left_bit_count_41 = 2'b01;
  assign _zz_129 = _zz_128[0 : 0];
  assign _zz_130 = _zz_129;
  assign all_zeros_80 = ((! (_zz_130 != 1'b0)) ? 1'b1 : 1'b0);
  assign all_left_zeros_80 = ((! (_zz_130[0 : 0] != 1'b0)) ? 1'b1 : 1'b0);
  assign left_all_zeros_count_38 = (all_left_zeros_79 & _zz_931);
  assign _zz_131 = _zz_128[1 : 1];
  assign _zz_132 = _zz_131;
  assign all_zeros_81 = ((! (_zz_132 != 1'b0)) ? 1'b1 : 1'b0);
  assign all_left_zeros_81 = ((! (_zz_132[0 : 0] != 1'b0)) ? 1'b1 : 1'b0);
  assign left_non_all_zeros_count_35 = ((~ all_left_zeros_79) & _zz_935);
  assign non_zeros_lzc_35 = (left_all_zeros_count_38 + left_non_all_zeros_count_35);
  assign left_non_all_zeros_count_36 = ((~ all_left_zeros_75) & _zz_937);
  assign non_zeros_lzc_36 = (left_all_zeros_count_37 + left_non_all_zeros_count_36);
  assign left_non_all_zeros_count_37 = ((~ all_left_zeros_67) & _zz_940);
  assign non_zeros_lzc_37 = (left_all_zeros_count_35 + left_non_all_zeros_count_37);
  assign left_all_zeros_count_39 = (all_left_zeros_66 & _zz_942);
  assign _zz_133 = _zz_109[15 : 8];
  assign all_zeros_82 = ((! (_zz_133 != 8'h0)) ? 4'b1111 : 4'b0000);
  assign all_left_zeros_82 = ((! (_zz_133[7 : 4] != 4'b0000)) ? 4'b1111 : 4'b0000);
  assign whole_bit_count_42 = 4'b1000;
  assign left_bit_count_42 = 4'b0100;
  assign _zz_134 = _zz_133[3 : 0];
  assign all_zeros_83 = ((! (_zz_134 != 4'b0000)) ? 3'b111 : 3'b000);
  assign all_left_zeros_83 = ((! (_zz_134[3 : 2] != 2'b00)) ? 3'b111 : 3'b000);
  assign whole_bit_count_43 = 3'b100;
  assign left_bit_count_43 = 3'b010;
  assign _zz_135 = _zz_134[1 : 0];
  assign all_zeros_84 = ((! (_zz_135 != 2'b00)) ? 2'b11 : 2'b00);
  assign all_left_zeros_84 = ((! (_zz_135[1 : 1] != 1'b0)) ? 2'b11 : 2'b00);
  assign whole_bit_count_44 = 2'b10;
  assign left_bit_count_44 = 2'b01;
  assign _zz_136 = _zz_135[0 : 0];
  assign _zz_137 = _zz_136;
  assign all_zeros_85 = ((! (_zz_137 != 1'b0)) ? 1'b1 : 1'b0);
  assign all_left_zeros_85 = ((! (_zz_137[0 : 0] != 1'b0)) ? 1'b1 : 1'b0);
  assign left_all_zeros_count_40 = (all_left_zeros_84 & _zz_946);
  assign _zz_138 = _zz_135[1 : 1];
  assign _zz_139 = _zz_138;
  assign all_zeros_86 = ((! (_zz_139 != 1'b0)) ? 1'b1 : 1'b0);
  assign all_left_zeros_86 = ((! (_zz_139[0 : 0] != 1'b0)) ? 1'b1 : 1'b0);
  assign left_non_all_zeros_count_38 = ((~ all_left_zeros_84) & _zz_950);
  assign non_zeros_lzc_38 = (left_all_zeros_count_40 + left_non_all_zeros_count_38);
  assign left_all_zeros_count_41 = (all_left_zeros_83 & _zz_951);
  assign _zz_140 = _zz_134[3 : 2];
  assign all_zeros_87 = ((! (_zz_140 != 2'b00)) ? 2'b11 : 2'b00);
  assign all_left_zeros_87 = ((! (_zz_140[1 : 1] != 1'b0)) ? 2'b11 : 2'b00);
  assign whole_bit_count_45 = 2'b10;
  assign left_bit_count_45 = 2'b01;
  assign _zz_141 = _zz_140[0 : 0];
  assign _zz_142 = _zz_141;
  assign all_zeros_88 = ((! (_zz_142 != 1'b0)) ? 1'b1 : 1'b0);
  assign all_left_zeros_88 = ((! (_zz_142[0 : 0] != 1'b0)) ? 1'b1 : 1'b0);
  assign left_all_zeros_count_42 = (all_left_zeros_87 & _zz_955);
  assign _zz_143 = _zz_140[1 : 1];
  assign _zz_144 = _zz_143;
  assign all_zeros_89 = ((! (_zz_144 != 1'b0)) ? 1'b1 : 1'b0);
  assign all_left_zeros_89 = ((! (_zz_144[0 : 0] != 1'b0)) ? 1'b1 : 1'b0);
  assign left_non_all_zeros_count_39 = ((~ all_left_zeros_87) & _zz_959);
  assign non_zeros_lzc_39 = (left_all_zeros_count_42 + left_non_all_zeros_count_39);
  assign left_non_all_zeros_count_40 = ((~ all_left_zeros_83) & _zz_961);
  assign non_zeros_lzc_40 = (left_all_zeros_count_41 + left_non_all_zeros_count_40);
  assign left_all_zeros_count_43 = (all_left_zeros_82 & _zz_963);
  assign _zz_145 = _zz_133[7 : 4];
  assign all_zeros_90 = ((! (_zz_145 != 4'b0000)) ? 3'b111 : 3'b000);
  assign all_left_zeros_90 = ((! (_zz_145[3 : 2] != 2'b00)) ? 3'b111 : 3'b000);
  assign whole_bit_count_46 = 3'b100;
  assign left_bit_count_46 = 3'b010;
  assign _zz_146 = _zz_145[1 : 0];
  assign all_zeros_91 = ((! (_zz_146 != 2'b00)) ? 2'b11 : 2'b00);
  assign all_left_zeros_91 = ((! (_zz_146[1 : 1] != 1'b0)) ? 2'b11 : 2'b00);
  assign whole_bit_count_47 = 2'b10;
  assign left_bit_count_47 = 2'b01;
  assign _zz_147 = _zz_146[0 : 0];
  assign _zz_148 = _zz_147;
  assign all_zeros_92 = ((! (_zz_148 != 1'b0)) ? 1'b1 : 1'b0);
  assign all_left_zeros_92 = ((! (_zz_148[0 : 0] != 1'b0)) ? 1'b1 : 1'b0);
  assign left_all_zeros_count_44 = (all_left_zeros_91 & _zz_967);
  assign _zz_149 = _zz_146[1 : 1];
  assign _zz_150 = _zz_149;
  assign all_zeros_93 = ((! (_zz_150 != 1'b0)) ? 1'b1 : 1'b0);
  assign all_left_zeros_93 = ((! (_zz_150[0 : 0] != 1'b0)) ? 1'b1 : 1'b0);
  assign left_non_all_zeros_count_41 = ((~ all_left_zeros_91) & _zz_971);
  assign non_zeros_lzc_41 = (left_all_zeros_count_44 + left_non_all_zeros_count_41);
  assign left_all_zeros_count_45 = (all_left_zeros_90 & _zz_972);
  assign _zz_151 = _zz_145[3 : 2];
  assign all_zeros_94 = ((! (_zz_151 != 2'b00)) ? 2'b11 : 2'b00);
  assign all_left_zeros_94 = ((! (_zz_151[1 : 1] != 1'b0)) ? 2'b11 : 2'b00);
  assign whole_bit_count_48 = 2'b10;
  assign left_bit_count_48 = 2'b01;
  assign _zz_152 = _zz_151[0 : 0];
  assign _zz_153 = _zz_152;
  assign all_zeros_95 = ((! (_zz_153 != 1'b0)) ? 1'b1 : 1'b0);
  assign all_left_zeros_95 = ((! (_zz_153[0 : 0] != 1'b0)) ? 1'b1 : 1'b0);
  assign left_all_zeros_count_46 = (all_left_zeros_94 & _zz_976);
  assign _zz_154 = _zz_151[1 : 1];
  assign _zz_155 = _zz_154;
  assign all_zeros_96 = ((! (_zz_155 != 1'b0)) ? 1'b1 : 1'b0);
  assign all_left_zeros_96 = ((! (_zz_155[0 : 0] != 1'b0)) ? 1'b1 : 1'b0);
  assign left_non_all_zeros_count_42 = ((~ all_left_zeros_94) & _zz_980);
  assign non_zeros_lzc_42 = (left_all_zeros_count_46 + left_non_all_zeros_count_42);
  assign left_non_all_zeros_count_43 = ((~ all_left_zeros_90) & _zz_982);
  assign non_zeros_lzc_43 = (left_all_zeros_count_45 + left_non_all_zeros_count_43);
  assign left_non_all_zeros_count_44 = ((~ all_left_zeros_82) & _zz_985);
  assign non_zeros_lzc_44 = (left_all_zeros_count_43 + left_non_all_zeros_count_44);
  assign left_non_all_zeros_count_45 = ((~ all_left_zeros_66) & _zz_988);
  assign non_zeros_lzc_45 = (left_all_zeros_count_39 + left_non_all_zeros_count_45);
  assign left_all_zeros_count_47 = (all_left_zeros_65 & _zz_990);
  assign _zz_156 = _zz_108[31 : 16];
  assign all_zeros_97 = ((! (_zz_156 != 16'h0)) ? 5'h1f : 5'h0);
  assign all_left_zeros_97 = ((! (_zz_156[15 : 8] != 8'h0)) ? 5'h1f : 5'h0);
  assign whole_bit_count_49 = 5'h10;
  assign left_bit_count_49 = 5'h08;
  assign _zz_157 = _zz_156[7 : 0];
  assign all_zeros_98 = ((! (_zz_157 != 8'h0)) ? 4'b1111 : 4'b0000);
  assign all_left_zeros_98 = ((! (_zz_157[7 : 4] != 4'b0000)) ? 4'b1111 : 4'b0000);
  assign whole_bit_count_50 = 4'b1000;
  assign left_bit_count_50 = 4'b0100;
  assign _zz_158 = _zz_157[3 : 0];
  assign all_zeros_99 = ((! (_zz_158 != 4'b0000)) ? 3'b111 : 3'b000);
  assign all_left_zeros_99 = ((! (_zz_158[3 : 2] != 2'b00)) ? 3'b111 : 3'b000);
  assign whole_bit_count_51 = 3'b100;
  assign left_bit_count_51 = 3'b010;
  assign _zz_159 = _zz_158[1 : 0];
  assign all_zeros_100 = ((! (_zz_159 != 2'b00)) ? 2'b11 : 2'b00);
  assign all_left_zeros_100 = ((! (_zz_159[1 : 1] != 1'b0)) ? 2'b11 : 2'b00);
  assign whole_bit_count_52 = 2'b10;
  assign left_bit_count_52 = 2'b01;
  assign _zz_160 = _zz_159[0 : 0];
  assign _zz_161 = _zz_160;
  assign all_zeros_101 = ((! (_zz_161 != 1'b0)) ? 1'b1 : 1'b0);
  assign all_left_zeros_101 = ((! (_zz_161[0 : 0] != 1'b0)) ? 1'b1 : 1'b0);
  assign left_all_zeros_count_48 = (all_left_zeros_100 & _zz_994);
  assign _zz_162 = _zz_159[1 : 1];
  assign _zz_163 = _zz_162;
  assign all_zeros_102 = ((! (_zz_163 != 1'b0)) ? 1'b1 : 1'b0);
  assign all_left_zeros_102 = ((! (_zz_163[0 : 0] != 1'b0)) ? 1'b1 : 1'b0);
  assign left_non_all_zeros_count_46 = ((~ all_left_zeros_100) & _zz_998);
  assign non_zeros_lzc_46 = (left_all_zeros_count_48 + left_non_all_zeros_count_46);
  assign left_all_zeros_count_49 = (all_left_zeros_99 & _zz_999);
  assign _zz_164 = _zz_158[3 : 2];
  assign all_zeros_103 = ((! (_zz_164 != 2'b00)) ? 2'b11 : 2'b00);
  assign all_left_zeros_103 = ((! (_zz_164[1 : 1] != 1'b0)) ? 2'b11 : 2'b00);
  assign whole_bit_count_53 = 2'b10;
  assign left_bit_count_53 = 2'b01;
  assign _zz_165 = _zz_164[0 : 0];
  assign _zz_166 = _zz_165;
  assign all_zeros_104 = ((! (_zz_166 != 1'b0)) ? 1'b1 : 1'b0);
  assign all_left_zeros_104 = ((! (_zz_166[0 : 0] != 1'b0)) ? 1'b1 : 1'b0);
  assign left_all_zeros_count_50 = (all_left_zeros_103 & _zz_1003);
  assign _zz_167 = _zz_164[1 : 1];
  assign _zz_168 = _zz_167;
  assign all_zeros_105 = ((! (_zz_168 != 1'b0)) ? 1'b1 : 1'b0);
  assign all_left_zeros_105 = ((! (_zz_168[0 : 0] != 1'b0)) ? 1'b1 : 1'b0);
  assign left_non_all_zeros_count_47 = ((~ all_left_zeros_103) & _zz_1007);
  assign non_zeros_lzc_47 = (left_all_zeros_count_50 + left_non_all_zeros_count_47);
  assign left_non_all_zeros_count_48 = ((~ all_left_zeros_99) & _zz_1009);
  assign non_zeros_lzc_48 = (left_all_zeros_count_49 + left_non_all_zeros_count_48);
  assign left_all_zeros_count_51 = (all_left_zeros_98 & _zz_1011);
  assign _zz_169 = _zz_157[7 : 4];
  assign all_zeros_106 = ((! (_zz_169 != 4'b0000)) ? 3'b111 : 3'b000);
  assign all_left_zeros_106 = ((! (_zz_169[3 : 2] != 2'b00)) ? 3'b111 : 3'b000);
  assign whole_bit_count_54 = 3'b100;
  assign left_bit_count_54 = 3'b010;
  assign _zz_170 = _zz_169[1 : 0];
  assign all_zeros_107 = ((! (_zz_170 != 2'b00)) ? 2'b11 : 2'b00);
  assign all_left_zeros_107 = ((! (_zz_170[1 : 1] != 1'b0)) ? 2'b11 : 2'b00);
  assign whole_bit_count_55 = 2'b10;
  assign left_bit_count_55 = 2'b01;
  assign _zz_171 = _zz_170[0 : 0];
  assign _zz_172 = _zz_171;
  assign all_zeros_108 = ((! (_zz_172 != 1'b0)) ? 1'b1 : 1'b0);
  assign all_left_zeros_108 = ((! (_zz_172[0 : 0] != 1'b0)) ? 1'b1 : 1'b0);
  assign left_all_zeros_count_52 = (all_left_zeros_107 & _zz_1015);
  assign _zz_173 = _zz_170[1 : 1];
  assign _zz_174 = _zz_173;
  assign all_zeros_109 = ((! (_zz_174 != 1'b0)) ? 1'b1 : 1'b0);
  assign all_left_zeros_109 = ((! (_zz_174[0 : 0] != 1'b0)) ? 1'b1 : 1'b0);
  assign left_non_all_zeros_count_49 = ((~ all_left_zeros_107) & _zz_1019);
  assign non_zeros_lzc_49 = (left_all_zeros_count_52 + left_non_all_zeros_count_49);
  assign left_all_zeros_count_53 = (all_left_zeros_106 & _zz_1020);
  assign _zz_175 = _zz_169[3 : 2];
  assign all_zeros_110 = ((! (_zz_175 != 2'b00)) ? 2'b11 : 2'b00);
  assign all_left_zeros_110 = ((! (_zz_175[1 : 1] != 1'b0)) ? 2'b11 : 2'b00);
  assign whole_bit_count_56 = 2'b10;
  assign left_bit_count_56 = 2'b01;
  assign _zz_176 = _zz_175[0 : 0];
  assign _zz_177 = _zz_176;
  assign all_zeros_111 = ((! (_zz_177 != 1'b0)) ? 1'b1 : 1'b0);
  assign all_left_zeros_111 = ((! (_zz_177[0 : 0] != 1'b0)) ? 1'b1 : 1'b0);
  assign left_all_zeros_count_54 = (all_left_zeros_110 & _zz_1024);
  assign _zz_178 = _zz_175[1 : 1];
  assign _zz_179 = _zz_178;
  assign all_zeros_112 = ((! (_zz_179 != 1'b0)) ? 1'b1 : 1'b0);
  assign all_left_zeros_112 = ((! (_zz_179[0 : 0] != 1'b0)) ? 1'b1 : 1'b0);
  assign left_non_all_zeros_count_50 = ((~ all_left_zeros_110) & _zz_1028);
  assign non_zeros_lzc_50 = (left_all_zeros_count_54 + left_non_all_zeros_count_50);
  assign left_non_all_zeros_count_51 = ((~ all_left_zeros_106) & _zz_1030);
  assign non_zeros_lzc_51 = (left_all_zeros_count_53 + left_non_all_zeros_count_51);
  assign left_non_all_zeros_count_52 = ((~ all_left_zeros_98) & _zz_1033);
  assign non_zeros_lzc_52 = (left_all_zeros_count_51 + left_non_all_zeros_count_52);
  assign left_all_zeros_count_55 = (all_left_zeros_97 & _zz_1035);
  assign _zz_180 = _zz_156[15 : 8];
  assign all_zeros_113 = ((! (_zz_180 != 8'h0)) ? 4'b1111 : 4'b0000);
  assign all_left_zeros_113 = ((! (_zz_180[7 : 4] != 4'b0000)) ? 4'b1111 : 4'b0000);
  assign whole_bit_count_57 = 4'b1000;
  assign left_bit_count_57 = 4'b0100;
  assign _zz_181 = _zz_180[3 : 0];
  assign all_zeros_114 = ((! (_zz_181 != 4'b0000)) ? 3'b111 : 3'b000);
  assign all_left_zeros_114 = ((! (_zz_181[3 : 2] != 2'b00)) ? 3'b111 : 3'b000);
  assign whole_bit_count_58 = 3'b100;
  assign left_bit_count_58 = 3'b010;
  assign _zz_182 = _zz_181[1 : 0];
  assign all_zeros_115 = ((! (_zz_182 != 2'b00)) ? 2'b11 : 2'b00);
  assign all_left_zeros_115 = ((! (_zz_182[1 : 1] != 1'b0)) ? 2'b11 : 2'b00);
  assign whole_bit_count_59 = 2'b10;
  assign left_bit_count_59 = 2'b01;
  assign _zz_183 = _zz_182[0 : 0];
  assign _zz_184 = _zz_183;
  assign all_zeros_116 = ((! (_zz_184 != 1'b0)) ? 1'b1 : 1'b0);
  assign all_left_zeros_116 = ((! (_zz_184[0 : 0] != 1'b0)) ? 1'b1 : 1'b0);
  assign left_all_zeros_count_56 = (all_left_zeros_115 & _zz_1039);
  assign _zz_185 = _zz_182[1 : 1];
  assign _zz_186 = _zz_185;
  assign all_zeros_117 = ((! (_zz_186 != 1'b0)) ? 1'b1 : 1'b0);
  assign all_left_zeros_117 = ((! (_zz_186[0 : 0] != 1'b0)) ? 1'b1 : 1'b0);
  assign left_non_all_zeros_count_53 = ((~ all_left_zeros_115) & _zz_1043);
  assign non_zeros_lzc_53 = (left_all_zeros_count_56 + left_non_all_zeros_count_53);
  assign left_all_zeros_count_57 = (all_left_zeros_114 & _zz_1044);
  assign _zz_187 = _zz_181[3 : 2];
  assign all_zeros_118 = ((! (_zz_187 != 2'b00)) ? 2'b11 : 2'b00);
  assign all_left_zeros_118 = ((! (_zz_187[1 : 1] != 1'b0)) ? 2'b11 : 2'b00);
  assign whole_bit_count_60 = 2'b10;
  assign left_bit_count_60 = 2'b01;
  assign _zz_188 = _zz_187[0 : 0];
  assign _zz_189 = _zz_188;
  assign all_zeros_119 = ((! (_zz_189 != 1'b0)) ? 1'b1 : 1'b0);
  assign all_left_zeros_119 = ((! (_zz_189[0 : 0] != 1'b0)) ? 1'b1 : 1'b0);
  assign left_all_zeros_count_58 = (all_left_zeros_118 & _zz_1048);
  assign _zz_190 = _zz_187[1 : 1];
  assign _zz_191 = _zz_190;
  assign all_zeros_120 = ((! (_zz_191 != 1'b0)) ? 1'b1 : 1'b0);
  assign all_left_zeros_120 = ((! (_zz_191[0 : 0] != 1'b0)) ? 1'b1 : 1'b0);
  assign left_non_all_zeros_count_54 = ((~ all_left_zeros_118) & _zz_1052);
  assign non_zeros_lzc_54 = (left_all_zeros_count_58 + left_non_all_zeros_count_54);
  assign left_non_all_zeros_count_55 = ((~ all_left_zeros_114) & _zz_1054);
  assign non_zeros_lzc_55 = (left_all_zeros_count_57 + left_non_all_zeros_count_55);
  assign left_all_zeros_count_59 = (all_left_zeros_113 & _zz_1056);
  assign _zz_192 = _zz_180[7 : 4];
  assign all_zeros_121 = ((! (_zz_192 != 4'b0000)) ? 3'b111 : 3'b000);
  assign all_left_zeros_121 = ((! (_zz_192[3 : 2] != 2'b00)) ? 3'b111 : 3'b000);
  assign whole_bit_count_61 = 3'b100;
  assign left_bit_count_61 = 3'b010;
  assign _zz_193 = _zz_192[1 : 0];
  assign all_zeros_122 = ((! (_zz_193 != 2'b00)) ? 2'b11 : 2'b00);
  assign all_left_zeros_122 = ((! (_zz_193[1 : 1] != 1'b0)) ? 2'b11 : 2'b00);
  assign whole_bit_count_62 = 2'b10;
  assign left_bit_count_62 = 2'b01;
  assign _zz_194 = _zz_193[0 : 0];
  assign _zz_195 = _zz_194;
  assign all_zeros_123 = ((! (_zz_195 != 1'b0)) ? 1'b1 : 1'b0);
  assign all_left_zeros_123 = ((! (_zz_195[0 : 0] != 1'b0)) ? 1'b1 : 1'b0);
  assign left_all_zeros_count_60 = (all_left_zeros_122 & _zz_1060);
  assign _zz_196 = _zz_193[1 : 1];
  assign _zz_197 = _zz_196;
  assign all_zeros_124 = ((! (_zz_197 != 1'b0)) ? 1'b1 : 1'b0);
  assign all_left_zeros_124 = ((! (_zz_197[0 : 0] != 1'b0)) ? 1'b1 : 1'b0);
  assign left_non_all_zeros_count_56 = ((~ all_left_zeros_122) & _zz_1064);
  assign non_zeros_lzc_56 = (left_all_zeros_count_60 + left_non_all_zeros_count_56);
  assign left_all_zeros_count_61 = (all_left_zeros_121 & _zz_1065);
  assign _zz_198 = _zz_192[3 : 2];
  assign all_zeros_125 = ((! (_zz_198 != 2'b00)) ? 2'b11 : 2'b00);
  assign all_left_zeros_125 = ((! (_zz_198[1 : 1] != 1'b0)) ? 2'b11 : 2'b00);
  assign whole_bit_count_63 = 2'b10;
  assign left_bit_count_63 = 2'b01;
  assign _zz_199 = _zz_198[0 : 0];
  assign _zz_200 = _zz_199;
  assign all_zeros_126 = ((! (_zz_200 != 1'b0)) ? 1'b1 : 1'b0);
  assign all_left_zeros_126 = ((! (_zz_200[0 : 0] != 1'b0)) ? 1'b1 : 1'b0);
  assign left_all_zeros_count_62 = (all_left_zeros_125 & _zz_1069);
  assign _zz_201 = _zz_198[1 : 1];
  assign _zz_202 = _zz_201;
  assign all_zeros_127 = ((! (_zz_202 != 1'b0)) ? 1'b1 : 1'b0);
  assign all_left_zeros_127 = ((! (_zz_202[0 : 0] != 1'b0)) ? 1'b1 : 1'b0);
  assign left_non_all_zeros_count_57 = ((~ all_left_zeros_125) & _zz_1073);
  assign non_zeros_lzc_57 = (left_all_zeros_count_62 + left_non_all_zeros_count_57);
  assign left_non_all_zeros_count_58 = ((~ all_left_zeros_121) & _zz_1075);
  assign non_zeros_lzc_58 = (left_all_zeros_count_61 + left_non_all_zeros_count_58);
  assign left_non_all_zeros_count_59 = ((~ all_left_zeros_113) & _zz_1078);
  assign non_zeros_lzc_59 = (left_all_zeros_count_59 + left_non_all_zeros_count_59);
  assign left_non_all_zeros_count_60 = ((~ all_left_zeros_97) & _zz_1081);
  assign non_zeros_lzc_60 = (left_all_zeros_count_55 + left_non_all_zeros_count_60);
  assign left_non_all_zeros_count_61 = ((~ all_left_zeros_65) & _zz_1084);
  assign non_zeros_lzc_61 = (left_all_zeros_count_47 + left_non_all_zeros_count_61);
  assign left_non_all_zeros_count_62 = ((~ all_left_zeros_1) & _zz_1087);
  assign non_zeros_lzc_62 = (left_all_zeros_count_31 + left_non_all_zeros_count_62);
  assign left_all_zeros_count_63 = (all_left_zeros & _zz_1089);
  assign _zz_203 = _zz_11[127 : 64];
  assign all_zeros_128 = ((! (_zz_203 != 64'h0)) ? 7'h7f : 7'h0);
  assign all_left_zeros_128 = ((! (_zz_203[63 : 32] != 32'h0)) ? 7'h7f : 7'h0);
  assign whole_bit_count_64 = 7'h40;
  assign left_bit_count_64 = 7'h20;
  assign _zz_204 = _zz_203[31 : 0];
  assign all_zeros_129 = ((! (_zz_204 != 32'h0)) ? 6'h3f : 6'h0);
  assign all_left_zeros_129 = ((! (_zz_204[31 : 16] != 16'h0)) ? 6'h3f : 6'h0);
  assign whole_bit_count_65 = 6'h20;
  assign left_bit_count_65 = 6'h10;
  assign _zz_205 = _zz_204[15 : 0];
  assign all_zeros_130 = ((! (_zz_205 != 16'h0)) ? 5'h1f : 5'h0);
  assign all_left_zeros_130 = ((! (_zz_205[15 : 8] != 8'h0)) ? 5'h1f : 5'h0);
  assign whole_bit_count_66 = 5'h10;
  assign left_bit_count_66 = 5'h08;
  assign _zz_206 = _zz_205[7 : 0];
  assign all_zeros_131 = ((! (_zz_206 != 8'h0)) ? 4'b1111 : 4'b0000);
  assign all_left_zeros_131 = ((! (_zz_206[7 : 4] != 4'b0000)) ? 4'b1111 : 4'b0000);
  assign whole_bit_count_67 = 4'b1000;
  assign left_bit_count_67 = 4'b0100;
  assign _zz_207 = _zz_206[3 : 0];
  assign all_zeros_132 = ((! (_zz_207 != 4'b0000)) ? 3'b111 : 3'b000);
  assign all_left_zeros_132 = ((! (_zz_207[3 : 2] != 2'b00)) ? 3'b111 : 3'b000);
  assign whole_bit_count_68 = 3'b100;
  assign left_bit_count_68 = 3'b010;
  assign _zz_208 = _zz_207[1 : 0];
  assign all_zeros_133 = ((! (_zz_208 != 2'b00)) ? 2'b11 : 2'b00);
  assign all_left_zeros_133 = ((! (_zz_208[1 : 1] != 1'b0)) ? 2'b11 : 2'b00);
  assign whole_bit_count_69 = 2'b10;
  assign left_bit_count_69 = 2'b01;
  assign _zz_209 = _zz_208[0 : 0];
  assign _zz_210 = _zz_209;
  assign all_zeros_134 = ((! (_zz_210 != 1'b0)) ? 1'b1 : 1'b0);
  assign all_left_zeros_134 = ((! (_zz_210[0 : 0] != 1'b0)) ? 1'b1 : 1'b0);
  assign left_all_zeros_count_64 = (all_left_zeros_133 & _zz_1093);
  assign _zz_211 = _zz_208[1 : 1];
  assign _zz_212 = _zz_211;
  assign all_zeros_135 = ((! (_zz_212 != 1'b0)) ? 1'b1 : 1'b0);
  assign all_left_zeros_135 = ((! (_zz_212[0 : 0] != 1'b0)) ? 1'b1 : 1'b0);
  assign left_non_all_zeros_count_63 = ((~ all_left_zeros_133) & _zz_1097);
  assign non_zeros_lzc_63 = (left_all_zeros_count_64 + left_non_all_zeros_count_63);
  assign left_all_zeros_count_65 = (all_left_zeros_132 & _zz_1098);
  assign _zz_213 = _zz_207[3 : 2];
  assign all_zeros_136 = ((! (_zz_213 != 2'b00)) ? 2'b11 : 2'b00);
  assign all_left_zeros_136 = ((! (_zz_213[1 : 1] != 1'b0)) ? 2'b11 : 2'b00);
  assign whole_bit_count_70 = 2'b10;
  assign left_bit_count_70 = 2'b01;
  assign _zz_214 = _zz_213[0 : 0];
  assign _zz_215 = _zz_214;
  assign all_zeros_137 = ((! (_zz_215 != 1'b0)) ? 1'b1 : 1'b0);
  assign all_left_zeros_137 = ((! (_zz_215[0 : 0] != 1'b0)) ? 1'b1 : 1'b0);
  assign left_all_zeros_count_66 = (all_left_zeros_136 & _zz_1102);
  assign _zz_216 = _zz_213[1 : 1];
  assign _zz_217 = _zz_216;
  assign all_zeros_138 = ((! (_zz_217 != 1'b0)) ? 1'b1 : 1'b0);
  assign all_left_zeros_138 = ((! (_zz_217[0 : 0] != 1'b0)) ? 1'b1 : 1'b0);
  assign left_non_all_zeros_count_64 = ((~ all_left_zeros_136) & _zz_1106);
  assign non_zeros_lzc_64 = (left_all_zeros_count_66 + left_non_all_zeros_count_64);
  assign left_non_all_zeros_count_65 = ((~ all_left_zeros_132) & _zz_1108);
  assign non_zeros_lzc_65 = (left_all_zeros_count_65 + left_non_all_zeros_count_65);
  assign left_all_zeros_count_67 = (all_left_zeros_131 & _zz_1110);
  assign _zz_218 = _zz_206[7 : 4];
  assign all_zeros_139 = ((! (_zz_218 != 4'b0000)) ? 3'b111 : 3'b000);
  assign all_left_zeros_139 = ((! (_zz_218[3 : 2] != 2'b00)) ? 3'b111 : 3'b000);
  assign whole_bit_count_71 = 3'b100;
  assign left_bit_count_71 = 3'b010;
  assign _zz_219 = _zz_218[1 : 0];
  assign all_zeros_140 = ((! (_zz_219 != 2'b00)) ? 2'b11 : 2'b00);
  assign all_left_zeros_140 = ((! (_zz_219[1 : 1] != 1'b0)) ? 2'b11 : 2'b00);
  assign whole_bit_count_72 = 2'b10;
  assign left_bit_count_72 = 2'b01;
  assign _zz_220 = _zz_219[0 : 0];
  assign _zz_221 = _zz_220;
  assign all_zeros_141 = ((! (_zz_221 != 1'b0)) ? 1'b1 : 1'b0);
  assign all_left_zeros_141 = ((! (_zz_221[0 : 0] != 1'b0)) ? 1'b1 : 1'b0);
  assign left_all_zeros_count_68 = (all_left_zeros_140 & _zz_1114);
  assign _zz_222 = _zz_219[1 : 1];
  assign _zz_223 = _zz_222;
  assign all_zeros_142 = ((! (_zz_223 != 1'b0)) ? 1'b1 : 1'b0);
  assign all_left_zeros_142 = ((! (_zz_223[0 : 0] != 1'b0)) ? 1'b1 : 1'b0);
  assign left_non_all_zeros_count_66 = ((~ all_left_zeros_140) & _zz_1118);
  assign non_zeros_lzc_66 = (left_all_zeros_count_68 + left_non_all_zeros_count_66);
  assign left_all_zeros_count_69 = (all_left_zeros_139 & _zz_1119);
  assign _zz_224 = _zz_218[3 : 2];
  assign all_zeros_143 = ((! (_zz_224 != 2'b00)) ? 2'b11 : 2'b00);
  assign all_left_zeros_143 = ((! (_zz_224[1 : 1] != 1'b0)) ? 2'b11 : 2'b00);
  assign whole_bit_count_73 = 2'b10;
  assign left_bit_count_73 = 2'b01;
  assign _zz_225 = _zz_224[0 : 0];
  assign _zz_226 = _zz_225;
  assign all_zeros_144 = ((! (_zz_226 != 1'b0)) ? 1'b1 : 1'b0);
  assign all_left_zeros_144 = ((! (_zz_226[0 : 0] != 1'b0)) ? 1'b1 : 1'b0);
  assign left_all_zeros_count_70 = (all_left_zeros_143 & _zz_1123);
  assign _zz_227 = _zz_224[1 : 1];
  assign _zz_228 = _zz_227;
  assign all_zeros_145 = ((! (_zz_228 != 1'b0)) ? 1'b1 : 1'b0);
  assign all_left_zeros_145 = ((! (_zz_228[0 : 0] != 1'b0)) ? 1'b1 : 1'b0);
  assign left_non_all_zeros_count_67 = ((~ all_left_zeros_143) & _zz_1127);
  assign non_zeros_lzc_67 = (left_all_zeros_count_70 + left_non_all_zeros_count_67);
  assign left_non_all_zeros_count_68 = ((~ all_left_zeros_139) & _zz_1129);
  assign non_zeros_lzc_68 = (left_all_zeros_count_69 + left_non_all_zeros_count_68);
  assign left_non_all_zeros_count_69 = ((~ all_left_zeros_131) & _zz_1132);
  assign non_zeros_lzc_69 = (left_all_zeros_count_67 + left_non_all_zeros_count_69);
  assign left_all_zeros_count_71 = (all_left_zeros_130 & _zz_1134);
  assign _zz_229 = _zz_205[15 : 8];
  assign all_zeros_146 = ((! (_zz_229 != 8'h0)) ? 4'b1111 : 4'b0000);
  assign all_left_zeros_146 = ((! (_zz_229[7 : 4] != 4'b0000)) ? 4'b1111 : 4'b0000);
  assign whole_bit_count_74 = 4'b1000;
  assign left_bit_count_74 = 4'b0100;
  assign _zz_230 = _zz_229[3 : 0];
  assign all_zeros_147 = ((! (_zz_230 != 4'b0000)) ? 3'b111 : 3'b000);
  assign all_left_zeros_147 = ((! (_zz_230[3 : 2] != 2'b00)) ? 3'b111 : 3'b000);
  assign whole_bit_count_75 = 3'b100;
  assign left_bit_count_75 = 3'b010;
  assign _zz_231 = _zz_230[1 : 0];
  assign all_zeros_148 = ((! (_zz_231 != 2'b00)) ? 2'b11 : 2'b00);
  assign all_left_zeros_148 = ((! (_zz_231[1 : 1] != 1'b0)) ? 2'b11 : 2'b00);
  assign whole_bit_count_76 = 2'b10;
  assign left_bit_count_76 = 2'b01;
  assign _zz_232 = _zz_231[0 : 0];
  assign _zz_233 = _zz_232;
  assign all_zeros_149 = ((! (_zz_233 != 1'b0)) ? 1'b1 : 1'b0);
  assign all_left_zeros_149 = ((! (_zz_233[0 : 0] != 1'b0)) ? 1'b1 : 1'b0);
  assign left_all_zeros_count_72 = (all_left_zeros_148 & _zz_1138);
  assign _zz_234 = _zz_231[1 : 1];
  assign _zz_235 = _zz_234;
  assign all_zeros_150 = ((! (_zz_235 != 1'b0)) ? 1'b1 : 1'b0);
  assign all_left_zeros_150 = ((! (_zz_235[0 : 0] != 1'b0)) ? 1'b1 : 1'b0);
  assign left_non_all_zeros_count_70 = ((~ all_left_zeros_148) & _zz_1142);
  assign non_zeros_lzc_70 = (left_all_zeros_count_72 + left_non_all_zeros_count_70);
  assign left_all_zeros_count_73 = (all_left_zeros_147 & _zz_1143);
  assign _zz_236 = _zz_230[3 : 2];
  assign all_zeros_151 = ((! (_zz_236 != 2'b00)) ? 2'b11 : 2'b00);
  assign all_left_zeros_151 = ((! (_zz_236[1 : 1] != 1'b0)) ? 2'b11 : 2'b00);
  assign whole_bit_count_77 = 2'b10;
  assign left_bit_count_77 = 2'b01;
  assign _zz_237 = _zz_236[0 : 0];
  assign _zz_238 = _zz_237;
  assign all_zeros_152 = ((! (_zz_238 != 1'b0)) ? 1'b1 : 1'b0);
  assign all_left_zeros_152 = ((! (_zz_238[0 : 0] != 1'b0)) ? 1'b1 : 1'b0);
  assign left_all_zeros_count_74 = (all_left_zeros_151 & _zz_1147);
  assign _zz_239 = _zz_236[1 : 1];
  assign _zz_240 = _zz_239;
  assign all_zeros_153 = ((! (_zz_240 != 1'b0)) ? 1'b1 : 1'b0);
  assign all_left_zeros_153 = ((! (_zz_240[0 : 0] != 1'b0)) ? 1'b1 : 1'b0);
  assign left_non_all_zeros_count_71 = ((~ all_left_zeros_151) & _zz_1151);
  assign non_zeros_lzc_71 = (left_all_zeros_count_74 + left_non_all_zeros_count_71);
  assign left_non_all_zeros_count_72 = ((~ all_left_zeros_147) & _zz_1153);
  assign non_zeros_lzc_72 = (left_all_zeros_count_73 + left_non_all_zeros_count_72);
  assign left_all_zeros_count_75 = (all_left_zeros_146 & _zz_1155);
  assign _zz_241 = _zz_229[7 : 4];
  assign all_zeros_154 = ((! (_zz_241 != 4'b0000)) ? 3'b111 : 3'b000);
  assign all_left_zeros_154 = ((! (_zz_241[3 : 2] != 2'b00)) ? 3'b111 : 3'b000);
  assign whole_bit_count_78 = 3'b100;
  assign left_bit_count_78 = 3'b010;
  assign _zz_242 = _zz_241[1 : 0];
  assign all_zeros_155 = ((! (_zz_242 != 2'b00)) ? 2'b11 : 2'b00);
  assign all_left_zeros_155 = ((! (_zz_242[1 : 1] != 1'b0)) ? 2'b11 : 2'b00);
  assign whole_bit_count_79 = 2'b10;
  assign left_bit_count_79 = 2'b01;
  assign _zz_243 = _zz_242[0 : 0];
  assign _zz_244 = _zz_243;
  assign all_zeros_156 = ((! (_zz_244 != 1'b0)) ? 1'b1 : 1'b0);
  assign all_left_zeros_156 = ((! (_zz_244[0 : 0] != 1'b0)) ? 1'b1 : 1'b0);
  assign left_all_zeros_count_76 = (all_left_zeros_155 & _zz_1159);
  assign _zz_245 = _zz_242[1 : 1];
  assign _zz_246 = _zz_245;
  assign all_zeros_157 = ((! (_zz_246 != 1'b0)) ? 1'b1 : 1'b0);
  assign all_left_zeros_157 = ((! (_zz_246[0 : 0] != 1'b0)) ? 1'b1 : 1'b0);
  assign left_non_all_zeros_count_73 = ((~ all_left_zeros_155) & _zz_1163);
  assign non_zeros_lzc_73 = (left_all_zeros_count_76 + left_non_all_zeros_count_73);
  assign left_all_zeros_count_77 = (all_left_zeros_154 & _zz_1164);
  assign _zz_247 = _zz_241[3 : 2];
  assign all_zeros_158 = ((! (_zz_247 != 2'b00)) ? 2'b11 : 2'b00);
  assign all_left_zeros_158 = ((! (_zz_247[1 : 1] != 1'b0)) ? 2'b11 : 2'b00);
  assign whole_bit_count_80 = 2'b10;
  assign left_bit_count_80 = 2'b01;
  assign _zz_248 = _zz_247[0 : 0];
  assign _zz_249 = _zz_248;
  assign all_zeros_159 = ((! (_zz_249 != 1'b0)) ? 1'b1 : 1'b0);
  assign all_left_zeros_159 = ((! (_zz_249[0 : 0] != 1'b0)) ? 1'b1 : 1'b0);
  assign left_all_zeros_count_78 = (all_left_zeros_158 & _zz_1168);
  assign _zz_250 = _zz_247[1 : 1];
  assign _zz_251 = _zz_250;
  assign all_zeros_160 = ((! (_zz_251 != 1'b0)) ? 1'b1 : 1'b0);
  assign all_left_zeros_160 = ((! (_zz_251[0 : 0] != 1'b0)) ? 1'b1 : 1'b0);
  assign left_non_all_zeros_count_74 = ((~ all_left_zeros_158) & _zz_1172);
  assign non_zeros_lzc_74 = (left_all_zeros_count_78 + left_non_all_zeros_count_74);
  assign left_non_all_zeros_count_75 = ((~ all_left_zeros_154) & _zz_1174);
  assign non_zeros_lzc_75 = (left_all_zeros_count_77 + left_non_all_zeros_count_75);
  assign left_non_all_zeros_count_76 = ((~ all_left_zeros_146) & _zz_1177);
  assign non_zeros_lzc_76 = (left_all_zeros_count_75 + left_non_all_zeros_count_76);
  assign left_non_all_zeros_count_77 = ((~ all_left_zeros_130) & _zz_1180);
  assign non_zeros_lzc_77 = (left_all_zeros_count_71 + left_non_all_zeros_count_77);
  assign left_all_zeros_count_79 = (all_left_zeros_129 & _zz_1182);
  assign _zz_252 = _zz_204[31 : 16];
  assign all_zeros_161 = ((! (_zz_252 != 16'h0)) ? 5'h1f : 5'h0);
  assign all_left_zeros_161 = ((! (_zz_252[15 : 8] != 8'h0)) ? 5'h1f : 5'h0);
  assign whole_bit_count_81 = 5'h10;
  assign left_bit_count_81 = 5'h08;
  assign _zz_253 = _zz_252[7 : 0];
  assign all_zeros_162 = ((! (_zz_253 != 8'h0)) ? 4'b1111 : 4'b0000);
  assign all_left_zeros_162 = ((! (_zz_253[7 : 4] != 4'b0000)) ? 4'b1111 : 4'b0000);
  assign whole_bit_count_82 = 4'b1000;
  assign left_bit_count_82 = 4'b0100;
  assign _zz_254 = _zz_253[3 : 0];
  assign all_zeros_163 = ((! (_zz_254 != 4'b0000)) ? 3'b111 : 3'b000);
  assign all_left_zeros_163 = ((! (_zz_254[3 : 2] != 2'b00)) ? 3'b111 : 3'b000);
  assign whole_bit_count_83 = 3'b100;
  assign left_bit_count_83 = 3'b010;
  assign _zz_255 = _zz_254[1 : 0];
  assign all_zeros_164 = ((! (_zz_255 != 2'b00)) ? 2'b11 : 2'b00);
  assign all_left_zeros_164 = ((! (_zz_255[1 : 1] != 1'b0)) ? 2'b11 : 2'b00);
  assign whole_bit_count_84 = 2'b10;
  assign left_bit_count_84 = 2'b01;
  assign _zz_256 = _zz_255[0 : 0];
  assign _zz_257 = _zz_256;
  assign all_zeros_165 = ((! (_zz_257 != 1'b0)) ? 1'b1 : 1'b0);
  assign all_left_zeros_165 = ((! (_zz_257[0 : 0] != 1'b0)) ? 1'b1 : 1'b0);
  assign left_all_zeros_count_80 = (all_left_zeros_164 & _zz_1186);
  assign _zz_258 = _zz_255[1 : 1];
  assign _zz_259 = _zz_258;
  assign all_zeros_166 = ((! (_zz_259 != 1'b0)) ? 1'b1 : 1'b0);
  assign all_left_zeros_166 = ((! (_zz_259[0 : 0] != 1'b0)) ? 1'b1 : 1'b0);
  assign left_non_all_zeros_count_78 = ((~ all_left_zeros_164) & _zz_1190);
  assign non_zeros_lzc_78 = (left_all_zeros_count_80 + left_non_all_zeros_count_78);
  assign left_all_zeros_count_81 = (all_left_zeros_163 & _zz_1191);
  assign _zz_260 = _zz_254[3 : 2];
  assign all_zeros_167 = ((! (_zz_260 != 2'b00)) ? 2'b11 : 2'b00);
  assign all_left_zeros_167 = ((! (_zz_260[1 : 1] != 1'b0)) ? 2'b11 : 2'b00);
  assign whole_bit_count_85 = 2'b10;
  assign left_bit_count_85 = 2'b01;
  assign _zz_261 = _zz_260[0 : 0];
  assign _zz_262 = _zz_261;
  assign all_zeros_168 = ((! (_zz_262 != 1'b0)) ? 1'b1 : 1'b0);
  assign all_left_zeros_168 = ((! (_zz_262[0 : 0] != 1'b0)) ? 1'b1 : 1'b0);
  assign left_all_zeros_count_82 = (all_left_zeros_167 & _zz_1195);
  assign _zz_263 = _zz_260[1 : 1];
  assign _zz_264 = _zz_263;
  assign all_zeros_169 = ((! (_zz_264 != 1'b0)) ? 1'b1 : 1'b0);
  assign all_left_zeros_169 = ((! (_zz_264[0 : 0] != 1'b0)) ? 1'b1 : 1'b0);
  assign left_non_all_zeros_count_79 = ((~ all_left_zeros_167) & _zz_1199);
  assign non_zeros_lzc_79 = (left_all_zeros_count_82 + left_non_all_zeros_count_79);
  assign left_non_all_zeros_count_80 = ((~ all_left_zeros_163) & _zz_1201);
  assign non_zeros_lzc_80 = (left_all_zeros_count_81 + left_non_all_zeros_count_80);
  assign left_all_zeros_count_83 = (all_left_zeros_162 & _zz_1203);
  assign _zz_265 = _zz_253[7 : 4];
  assign all_zeros_170 = ((! (_zz_265 != 4'b0000)) ? 3'b111 : 3'b000);
  assign all_left_zeros_170 = ((! (_zz_265[3 : 2] != 2'b00)) ? 3'b111 : 3'b000);
  assign whole_bit_count_86 = 3'b100;
  assign left_bit_count_86 = 3'b010;
  assign _zz_266 = _zz_265[1 : 0];
  assign all_zeros_171 = ((! (_zz_266 != 2'b00)) ? 2'b11 : 2'b00);
  assign all_left_zeros_171 = ((! (_zz_266[1 : 1] != 1'b0)) ? 2'b11 : 2'b00);
  assign whole_bit_count_87 = 2'b10;
  assign left_bit_count_87 = 2'b01;
  assign _zz_267 = _zz_266[0 : 0];
  assign _zz_268 = _zz_267;
  assign all_zeros_172 = ((! (_zz_268 != 1'b0)) ? 1'b1 : 1'b0);
  assign all_left_zeros_172 = ((! (_zz_268[0 : 0] != 1'b0)) ? 1'b1 : 1'b0);
  assign left_all_zeros_count_84 = (all_left_zeros_171 & _zz_1207);
  assign _zz_269 = _zz_266[1 : 1];
  assign _zz_270 = _zz_269;
  assign all_zeros_173 = ((! (_zz_270 != 1'b0)) ? 1'b1 : 1'b0);
  assign all_left_zeros_173 = ((! (_zz_270[0 : 0] != 1'b0)) ? 1'b1 : 1'b0);
  assign left_non_all_zeros_count_81 = ((~ all_left_zeros_171) & _zz_1211);
  assign non_zeros_lzc_81 = (left_all_zeros_count_84 + left_non_all_zeros_count_81);
  assign left_all_zeros_count_85 = (all_left_zeros_170 & _zz_1212);
  assign _zz_271 = _zz_265[3 : 2];
  assign all_zeros_174 = ((! (_zz_271 != 2'b00)) ? 2'b11 : 2'b00);
  assign all_left_zeros_174 = ((! (_zz_271[1 : 1] != 1'b0)) ? 2'b11 : 2'b00);
  assign whole_bit_count_88 = 2'b10;
  assign left_bit_count_88 = 2'b01;
  assign _zz_272 = _zz_271[0 : 0];
  assign _zz_273 = _zz_272;
  assign all_zeros_175 = ((! (_zz_273 != 1'b0)) ? 1'b1 : 1'b0);
  assign all_left_zeros_175 = ((! (_zz_273[0 : 0] != 1'b0)) ? 1'b1 : 1'b0);
  assign left_all_zeros_count_86 = (all_left_zeros_174 & _zz_1216);
  assign _zz_274 = _zz_271[1 : 1];
  assign _zz_275 = _zz_274;
  assign all_zeros_176 = ((! (_zz_275 != 1'b0)) ? 1'b1 : 1'b0);
  assign all_left_zeros_176 = ((! (_zz_275[0 : 0] != 1'b0)) ? 1'b1 : 1'b0);
  assign left_non_all_zeros_count_82 = ((~ all_left_zeros_174) & _zz_1220);
  assign non_zeros_lzc_82 = (left_all_zeros_count_86 + left_non_all_zeros_count_82);
  assign left_non_all_zeros_count_83 = ((~ all_left_zeros_170) & _zz_1222);
  assign non_zeros_lzc_83 = (left_all_zeros_count_85 + left_non_all_zeros_count_83);
  assign left_non_all_zeros_count_84 = ((~ all_left_zeros_162) & _zz_1225);
  assign non_zeros_lzc_84 = (left_all_zeros_count_83 + left_non_all_zeros_count_84);
  assign left_all_zeros_count_87 = (all_left_zeros_161 & _zz_1227);
  assign _zz_276 = _zz_252[15 : 8];
  assign all_zeros_177 = ((! (_zz_276 != 8'h0)) ? 4'b1111 : 4'b0000);
  assign all_left_zeros_177 = ((! (_zz_276[7 : 4] != 4'b0000)) ? 4'b1111 : 4'b0000);
  assign whole_bit_count_89 = 4'b1000;
  assign left_bit_count_89 = 4'b0100;
  assign _zz_277 = _zz_276[3 : 0];
  assign all_zeros_178 = ((! (_zz_277 != 4'b0000)) ? 3'b111 : 3'b000);
  assign all_left_zeros_178 = ((! (_zz_277[3 : 2] != 2'b00)) ? 3'b111 : 3'b000);
  assign whole_bit_count_90 = 3'b100;
  assign left_bit_count_90 = 3'b010;
  assign _zz_278 = _zz_277[1 : 0];
  assign all_zeros_179 = ((! (_zz_278 != 2'b00)) ? 2'b11 : 2'b00);
  assign all_left_zeros_179 = ((! (_zz_278[1 : 1] != 1'b0)) ? 2'b11 : 2'b00);
  assign whole_bit_count_91 = 2'b10;
  assign left_bit_count_91 = 2'b01;
  assign _zz_279 = _zz_278[0 : 0];
  assign _zz_280 = _zz_279;
  assign all_zeros_180 = ((! (_zz_280 != 1'b0)) ? 1'b1 : 1'b0);
  assign all_left_zeros_180 = ((! (_zz_280[0 : 0] != 1'b0)) ? 1'b1 : 1'b0);
  assign left_all_zeros_count_88 = (all_left_zeros_179 & _zz_1231);
  assign _zz_281 = _zz_278[1 : 1];
  assign _zz_282 = _zz_281;
  assign all_zeros_181 = ((! (_zz_282 != 1'b0)) ? 1'b1 : 1'b0);
  assign all_left_zeros_181 = ((! (_zz_282[0 : 0] != 1'b0)) ? 1'b1 : 1'b0);
  assign left_non_all_zeros_count_85 = ((~ all_left_zeros_179) & _zz_1235);
  assign non_zeros_lzc_85 = (left_all_zeros_count_88 + left_non_all_zeros_count_85);
  assign left_all_zeros_count_89 = (all_left_zeros_178 & _zz_1236);
  assign _zz_283 = _zz_277[3 : 2];
  assign all_zeros_182 = ((! (_zz_283 != 2'b00)) ? 2'b11 : 2'b00);
  assign all_left_zeros_182 = ((! (_zz_283[1 : 1] != 1'b0)) ? 2'b11 : 2'b00);
  assign whole_bit_count_92 = 2'b10;
  assign left_bit_count_92 = 2'b01;
  assign _zz_284 = _zz_283[0 : 0];
  assign _zz_285 = _zz_284;
  assign all_zeros_183 = ((! (_zz_285 != 1'b0)) ? 1'b1 : 1'b0);
  assign all_left_zeros_183 = ((! (_zz_285[0 : 0] != 1'b0)) ? 1'b1 : 1'b0);
  assign left_all_zeros_count_90 = (all_left_zeros_182 & _zz_1240);
  assign _zz_286 = _zz_283[1 : 1];
  assign _zz_287 = _zz_286;
  assign all_zeros_184 = ((! (_zz_287 != 1'b0)) ? 1'b1 : 1'b0);
  assign all_left_zeros_184 = ((! (_zz_287[0 : 0] != 1'b0)) ? 1'b1 : 1'b0);
  assign left_non_all_zeros_count_86 = ((~ all_left_zeros_182) & _zz_1244);
  assign non_zeros_lzc_86 = (left_all_zeros_count_90 + left_non_all_zeros_count_86);
  assign left_non_all_zeros_count_87 = ((~ all_left_zeros_178) & _zz_1246);
  assign non_zeros_lzc_87 = (left_all_zeros_count_89 + left_non_all_zeros_count_87);
  assign left_all_zeros_count_91 = (all_left_zeros_177 & _zz_1248);
  assign _zz_288 = _zz_276[7 : 4];
  assign all_zeros_185 = ((! (_zz_288 != 4'b0000)) ? 3'b111 : 3'b000);
  assign all_left_zeros_185 = ((! (_zz_288[3 : 2] != 2'b00)) ? 3'b111 : 3'b000);
  assign whole_bit_count_93 = 3'b100;
  assign left_bit_count_93 = 3'b010;
  assign _zz_289 = _zz_288[1 : 0];
  assign all_zeros_186 = ((! (_zz_289 != 2'b00)) ? 2'b11 : 2'b00);
  assign all_left_zeros_186 = ((! (_zz_289[1 : 1] != 1'b0)) ? 2'b11 : 2'b00);
  assign whole_bit_count_94 = 2'b10;
  assign left_bit_count_94 = 2'b01;
  assign _zz_290 = _zz_289[0 : 0];
  assign _zz_291 = _zz_290;
  assign all_zeros_187 = ((! (_zz_291 != 1'b0)) ? 1'b1 : 1'b0);
  assign all_left_zeros_187 = ((! (_zz_291[0 : 0] != 1'b0)) ? 1'b1 : 1'b0);
  assign left_all_zeros_count_92 = (all_left_zeros_186 & _zz_1252);
  assign _zz_292 = _zz_289[1 : 1];
  assign _zz_293 = _zz_292;
  assign all_zeros_188 = ((! (_zz_293 != 1'b0)) ? 1'b1 : 1'b0);
  assign all_left_zeros_188 = ((! (_zz_293[0 : 0] != 1'b0)) ? 1'b1 : 1'b0);
  assign left_non_all_zeros_count_88 = ((~ all_left_zeros_186) & _zz_1256);
  assign non_zeros_lzc_88 = (left_all_zeros_count_92 + left_non_all_zeros_count_88);
  assign left_all_zeros_count_93 = (all_left_zeros_185 & _zz_1257);
  assign _zz_294 = _zz_288[3 : 2];
  assign all_zeros_189 = ((! (_zz_294 != 2'b00)) ? 2'b11 : 2'b00);
  assign all_left_zeros_189 = ((! (_zz_294[1 : 1] != 1'b0)) ? 2'b11 : 2'b00);
  assign whole_bit_count_95 = 2'b10;
  assign left_bit_count_95 = 2'b01;
  assign _zz_295 = _zz_294[0 : 0];
  assign _zz_296 = _zz_295;
  assign all_zeros_190 = ((! (_zz_296 != 1'b0)) ? 1'b1 : 1'b0);
  assign all_left_zeros_190 = ((! (_zz_296[0 : 0] != 1'b0)) ? 1'b1 : 1'b0);
  assign left_all_zeros_count_94 = (all_left_zeros_189 & _zz_1261);
  assign _zz_297 = _zz_294[1 : 1];
  assign _zz_298 = _zz_297;
  assign all_zeros_191 = ((! (_zz_298 != 1'b0)) ? 1'b1 : 1'b0);
  assign all_left_zeros_191 = ((! (_zz_298[0 : 0] != 1'b0)) ? 1'b1 : 1'b0);
  assign left_non_all_zeros_count_89 = ((~ all_left_zeros_189) & _zz_1265);
  assign non_zeros_lzc_89 = (left_all_zeros_count_94 + left_non_all_zeros_count_89);
  assign left_non_all_zeros_count_90 = ((~ all_left_zeros_185) & _zz_1267);
  assign non_zeros_lzc_90 = (left_all_zeros_count_93 + left_non_all_zeros_count_90);
  assign left_non_all_zeros_count_91 = ((~ all_left_zeros_177) & _zz_1270);
  assign non_zeros_lzc_91 = (left_all_zeros_count_91 + left_non_all_zeros_count_91);
  assign left_non_all_zeros_count_92 = ((~ all_left_zeros_161) & _zz_1273);
  assign non_zeros_lzc_92 = (left_all_zeros_count_87 + left_non_all_zeros_count_92);
  assign left_non_all_zeros_count_93 = ((~ all_left_zeros_129) & _zz_1276);
  assign non_zeros_lzc_93 = (left_all_zeros_count_79 + left_non_all_zeros_count_93);
  assign left_all_zeros_count_95 = (all_left_zeros_128 & _zz_1278);
  assign _zz_299 = _zz_203[63 : 32];
  assign all_zeros_192 = ((! (_zz_299 != 32'h0)) ? 6'h3f : 6'h0);
  assign all_left_zeros_192 = ((! (_zz_299[31 : 16] != 16'h0)) ? 6'h3f : 6'h0);
  assign whole_bit_count_96 = 6'h20;
  assign left_bit_count_96 = 6'h10;
  assign _zz_300 = _zz_299[15 : 0];
  assign all_zeros_193 = ((! (_zz_300 != 16'h0)) ? 5'h1f : 5'h0);
  assign all_left_zeros_193 = ((! (_zz_300[15 : 8] != 8'h0)) ? 5'h1f : 5'h0);
  assign whole_bit_count_97 = 5'h10;
  assign left_bit_count_97 = 5'h08;
  assign _zz_301 = _zz_300[7 : 0];
  assign all_zeros_194 = ((! (_zz_301 != 8'h0)) ? 4'b1111 : 4'b0000);
  assign all_left_zeros_194 = ((! (_zz_301[7 : 4] != 4'b0000)) ? 4'b1111 : 4'b0000);
  assign whole_bit_count_98 = 4'b1000;
  assign left_bit_count_98 = 4'b0100;
  assign _zz_302 = _zz_301[3 : 0];
  assign all_zeros_195 = ((! (_zz_302 != 4'b0000)) ? 3'b111 : 3'b000);
  assign all_left_zeros_195 = ((! (_zz_302[3 : 2] != 2'b00)) ? 3'b111 : 3'b000);
  assign whole_bit_count_99 = 3'b100;
  assign left_bit_count_99 = 3'b010;
  assign _zz_303 = _zz_302[1 : 0];
  assign all_zeros_196 = ((! (_zz_303 != 2'b00)) ? 2'b11 : 2'b00);
  assign all_left_zeros_196 = ((! (_zz_303[1 : 1] != 1'b0)) ? 2'b11 : 2'b00);
  assign whole_bit_count_100 = 2'b10;
  assign left_bit_count_100 = 2'b01;
  assign _zz_304 = _zz_303[0 : 0];
  assign _zz_305 = _zz_304;
  assign all_zeros_197 = ((! (_zz_305 != 1'b0)) ? 1'b1 : 1'b0);
  assign all_left_zeros_197 = ((! (_zz_305[0 : 0] != 1'b0)) ? 1'b1 : 1'b0);
  assign left_all_zeros_count_96 = (all_left_zeros_196 & _zz_1282);
  assign _zz_306 = _zz_303[1 : 1];
  assign _zz_307 = _zz_306;
  assign all_zeros_198 = ((! (_zz_307 != 1'b0)) ? 1'b1 : 1'b0);
  assign all_left_zeros_198 = ((! (_zz_307[0 : 0] != 1'b0)) ? 1'b1 : 1'b0);
  assign left_non_all_zeros_count_94 = ((~ all_left_zeros_196) & _zz_1286);
  assign non_zeros_lzc_94 = (left_all_zeros_count_96 + left_non_all_zeros_count_94);
  assign left_all_zeros_count_97 = (all_left_zeros_195 & _zz_1287);
  assign _zz_308 = _zz_302[3 : 2];
  assign all_zeros_199 = ((! (_zz_308 != 2'b00)) ? 2'b11 : 2'b00);
  assign all_left_zeros_199 = ((! (_zz_308[1 : 1] != 1'b0)) ? 2'b11 : 2'b00);
  assign whole_bit_count_101 = 2'b10;
  assign left_bit_count_101 = 2'b01;
  assign _zz_309 = _zz_308[0 : 0];
  assign _zz_310 = _zz_309;
  assign all_zeros_200 = ((! (_zz_310 != 1'b0)) ? 1'b1 : 1'b0);
  assign all_left_zeros_200 = ((! (_zz_310[0 : 0] != 1'b0)) ? 1'b1 : 1'b0);
  assign left_all_zeros_count_98 = (all_left_zeros_199 & _zz_1291);
  assign _zz_311 = _zz_308[1 : 1];
  assign _zz_312 = _zz_311;
  assign all_zeros_201 = ((! (_zz_312 != 1'b0)) ? 1'b1 : 1'b0);
  assign all_left_zeros_201 = ((! (_zz_312[0 : 0] != 1'b0)) ? 1'b1 : 1'b0);
  assign left_non_all_zeros_count_95 = ((~ all_left_zeros_199) & _zz_1295);
  assign non_zeros_lzc_95 = (left_all_zeros_count_98 + left_non_all_zeros_count_95);
  assign left_non_all_zeros_count_96 = ((~ all_left_zeros_195) & _zz_1297);
  assign non_zeros_lzc_96 = (left_all_zeros_count_97 + left_non_all_zeros_count_96);
  assign left_all_zeros_count_99 = (all_left_zeros_194 & _zz_1299);
  assign _zz_313 = _zz_301[7 : 4];
  assign all_zeros_202 = ((! (_zz_313 != 4'b0000)) ? 3'b111 : 3'b000);
  assign all_left_zeros_202 = ((! (_zz_313[3 : 2] != 2'b00)) ? 3'b111 : 3'b000);
  assign whole_bit_count_102 = 3'b100;
  assign left_bit_count_102 = 3'b010;
  assign _zz_314 = _zz_313[1 : 0];
  assign all_zeros_203 = ((! (_zz_314 != 2'b00)) ? 2'b11 : 2'b00);
  assign all_left_zeros_203 = ((! (_zz_314[1 : 1] != 1'b0)) ? 2'b11 : 2'b00);
  assign whole_bit_count_103 = 2'b10;
  assign left_bit_count_103 = 2'b01;
  assign _zz_315 = _zz_314[0 : 0];
  assign _zz_316 = _zz_315;
  assign all_zeros_204 = ((! (_zz_316 != 1'b0)) ? 1'b1 : 1'b0);
  assign all_left_zeros_204 = ((! (_zz_316[0 : 0] != 1'b0)) ? 1'b1 : 1'b0);
  assign left_all_zeros_count_100 = (all_left_zeros_203 & _zz_1303);
  assign _zz_317 = _zz_314[1 : 1];
  assign _zz_318 = _zz_317;
  assign all_zeros_205 = ((! (_zz_318 != 1'b0)) ? 1'b1 : 1'b0);
  assign all_left_zeros_205 = ((! (_zz_318[0 : 0] != 1'b0)) ? 1'b1 : 1'b0);
  assign left_non_all_zeros_count_97 = ((~ all_left_zeros_203) & _zz_1307);
  assign non_zeros_lzc_97 = (left_all_zeros_count_100 + left_non_all_zeros_count_97);
  assign left_all_zeros_count_101 = (all_left_zeros_202 & _zz_1308);
  assign _zz_319 = _zz_313[3 : 2];
  assign all_zeros_206 = ((! (_zz_319 != 2'b00)) ? 2'b11 : 2'b00);
  assign all_left_zeros_206 = ((! (_zz_319[1 : 1] != 1'b0)) ? 2'b11 : 2'b00);
  assign whole_bit_count_104 = 2'b10;
  assign left_bit_count_104 = 2'b01;
  assign _zz_320 = _zz_319[0 : 0];
  assign _zz_321 = _zz_320;
  assign all_zeros_207 = ((! (_zz_321 != 1'b0)) ? 1'b1 : 1'b0);
  assign all_left_zeros_207 = ((! (_zz_321[0 : 0] != 1'b0)) ? 1'b1 : 1'b0);
  assign left_all_zeros_count_102 = (all_left_zeros_206 & _zz_1312);
  assign _zz_322 = _zz_319[1 : 1];
  assign _zz_323 = _zz_322;
  assign all_zeros_208 = ((! (_zz_323 != 1'b0)) ? 1'b1 : 1'b0);
  assign all_left_zeros_208 = ((! (_zz_323[0 : 0] != 1'b0)) ? 1'b1 : 1'b0);
  assign left_non_all_zeros_count_98 = ((~ all_left_zeros_206) & _zz_1316);
  assign non_zeros_lzc_98 = (left_all_zeros_count_102 + left_non_all_zeros_count_98);
  assign left_non_all_zeros_count_99 = ((~ all_left_zeros_202) & _zz_1318);
  assign non_zeros_lzc_99 = (left_all_zeros_count_101 + left_non_all_zeros_count_99);
  assign left_non_all_zeros_count_100 = ((~ all_left_zeros_194) & _zz_1321);
  assign non_zeros_lzc_100 = (left_all_zeros_count_99 + left_non_all_zeros_count_100);
  assign left_all_zeros_count_103 = (all_left_zeros_193 & _zz_1323);
  assign _zz_324 = _zz_300[15 : 8];
  assign all_zeros_209 = ((! (_zz_324 != 8'h0)) ? 4'b1111 : 4'b0000);
  assign all_left_zeros_209 = ((! (_zz_324[7 : 4] != 4'b0000)) ? 4'b1111 : 4'b0000);
  assign whole_bit_count_105 = 4'b1000;
  assign left_bit_count_105 = 4'b0100;
  assign _zz_325 = _zz_324[3 : 0];
  assign all_zeros_210 = ((! (_zz_325 != 4'b0000)) ? 3'b111 : 3'b000);
  assign all_left_zeros_210 = ((! (_zz_325[3 : 2] != 2'b00)) ? 3'b111 : 3'b000);
  assign whole_bit_count_106 = 3'b100;
  assign left_bit_count_106 = 3'b010;
  assign _zz_326 = _zz_325[1 : 0];
  assign all_zeros_211 = ((! (_zz_326 != 2'b00)) ? 2'b11 : 2'b00);
  assign all_left_zeros_211 = ((! (_zz_326[1 : 1] != 1'b0)) ? 2'b11 : 2'b00);
  assign whole_bit_count_107 = 2'b10;
  assign left_bit_count_107 = 2'b01;
  assign _zz_327 = _zz_326[0 : 0];
  assign _zz_328 = _zz_327;
  assign all_zeros_212 = ((! (_zz_328 != 1'b0)) ? 1'b1 : 1'b0);
  assign all_left_zeros_212 = ((! (_zz_328[0 : 0] != 1'b0)) ? 1'b1 : 1'b0);
  assign left_all_zeros_count_104 = (all_left_zeros_211 & _zz_1327);
  assign _zz_329 = _zz_326[1 : 1];
  assign _zz_330 = _zz_329;
  assign all_zeros_213 = ((! (_zz_330 != 1'b0)) ? 1'b1 : 1'b0);
  assign all_left_zeros_213 = ((! (_zz_330[0 : 0] != 1'b0)) ? 1'b1 : 1'b0);
  assign left_non_all_zeros_count_101 = ((~ all_left_zeros_211) & _zz_1331);
  assign non_zeros_lzc_101 = (left_all_zeros_count_104 + left_non_all_zeros_count_101);
  assign left_all_zeros_count_105 = (all_left_zeros_210 & _zz_1332);
  assign _zz_331 = _zz_325[3 : 2];
  assign all_zeros_214 = ((! (_zz_331 != 2'b00)) ? 2'b11 : 2'b00);
  assign all_left_zeros_214 = ((! (_zz_331[1 : 1] != 1'b0)) ? 2'b11 : 2'b00);
  assign whole_bit_count_108 = 2'b10;
  assign left_bit_count_108 = 2'b01;
  assign _zz_332 = _zz_331[0 : 0];
  assign _zz_333 = _zz_332;
  assign all_zeros_215 = ((! (_zz_333 != 1'b0)) ? 1'b1 : 1'b0);
  assign all_left_zeros_215 = ((! (_zz_333[0 : 0] != 1'b0)) ? 1'b1 : 1'b0);
  assign left_all_zeros_count_106 = (all_left_zeros_214 & _zz_1336);
  assign _zz_334 = _zz_331[1 : 1];
  assign _zz_335 = _zz_334;
  assign all_zeros_216 = ((! (_zz_335 != 1'b0)) ? 1'b1 : 1'b0);
  assign all_left_zeros_216 = ((! (_zz_335[0 : 0] != 1'b0)) ? 1'b1 : 1'b0);
  assign left_non_all_zeros_count_102 = ((~ all_left_zeros_214) & _zz_1340);
  assign non_zeros_lzc_102 = (left_all_zeros_count_106 + left_non_all_zeros_count_102);
  assign left_non_all_zeros_count_103 = ((~ all_left_zeros_210) & _zz_1342);
  assign non_zeros_lzc_103 = (left_all_zeros_count_105 + left_non_all_zeros_count_103);
  assign left_all_zeros_count_107 = (all_left_zeros_209 & _zz_1344);
  assign _zz_336 = _zz_324[7 : 4];
  assign all_zeros_217 = ((! (_zz_336 != 4'b0000)) ? 3'b111 : 3'b000);
  assign all_left_zeros_217 = ((! (_zz_336[3 : 2] != 2'b00)) ? 3'b111 : 3'b000);
  assign whole_bit_count_109 = 3'b100;
  assign left_bit_count_109 = 3'b010;
  assign _zz_337 = _zz_336[1 : 0];
  assign all_zeros_218 = ((! (_zz_337 != 2'b00)) ? 2'b11 : 2'b00);
  assign all_left_zeros_218 = ((! (_zz_337[1 : 1] != 1'b0)) ? 2'b11 : 2'b00);
  assign whole_bit_count_110 = 2'b10;
  assign left_bit_count_110 = 2'b01;
  assign _zz_338 = _zz_337[0 : 0];
  assign _zz_339 = _zz_338;
  assign all_zeros_219 = ((! (_zz_339 != 1'b0)) ? 1'b1 : 1'b0);
  assign all_left_zeros_219 = ((! (_zz_339[0 : 0] != 1'b0)) ? 1'b1 : 1'b0);
  assign left_all_zeros_count_108 = (all_left_zeros_218 & _zz_1348);
  assign _zz_340 = _zz_337[1 : 1];
  assign _zz_341 = _zz_340;
  assign all_zeros_220 = ((! (_zz_341 != 1'b0)) ? 1'b1 : 1'b0);
  assign all_left_zeros_220 = ((! (_zz_341[0 : 0] != 1'b0)) ? 1'b1 : 1'b0);
  assign left_non_all_zeros_count_104 = ((~ all_left_zeros_218) & _zz_1352);
  assign non_zeros_lzc_104 = (left_all_zeros_count_108 + left_non_all_zeros_count_104);
  assign left_all_zeros_count_109 = (all_left_zeros_217 & _zz_1353);
  assign _zz_342 = _zz_336[3 : 2];
  assign all_zeros_221 = ((! (_zz_342 != 2'b00)) ? 2'b11 : 2'b00);
  assign all_left_zeros_221 = ((! (_zz_342[1 : 1] != 1'b0)) ? 2'b11 : 2'b00);
  assign whole_bit_count_111 = 2'b10;
  assign left_bit_count_111 = 2'b01;
  assign _zz_343 = _zz_342[0 : 0];
  assign _zz_344 = _zz_343;
  assign all_zeros_222 = ((! (_zz_344 != 1'b0)) ? 1'b1 : 1'b0);
  assign all_left_zeros_222 = ((! (_zz_344[0 : 0] != 1'b0)) ? 1'b1 : 1'b0);
  assign left_all_zeros_count_110 = (all_left_zeros_221 & _zz_1357);
  assign _zz_345 = _zz_342[1 : 1];
  assign _zz_346 = _zz_345;
  assign all_zeros_223 = ((! (_zz_346 != 1'b0)) ? 1'b1 : 1'b0);
  assign all_left_zeros_223 = ((! (_zz_346[0 : 0] != 1'b0)) ? 1'b1 : 1'b0);
  assign left_non_all_zeros_count_105 = ((~ all_left_zeros_221) & _zz_1361);
  assign non_zeros_lzc_105 = (left_all_zeros_count_110 + left_non_all_zeros_count_105);
  assign left_non_all_zeros_count_106 = ((~ all_left_zeros_217) & _zz_1363);
  assign non_zeros_lzc_106 = (left_all_zeros_count_109 + left_non_all_zeros_count_106);
  assign left_non_all_zeros_count_107 = ((~ all_left_zeros_209) & _zz_1366);
  assign non_zeros_lzc_107 = (left_all_zeros_count_107 + left_non_all_zeros_count_107);
  assign left_non_all_zeros_count_108 = ((~ all_left_zeros_193) & _zz_1369);
  assign non_zeros_lzc_108 = (left_all_zeros_count_103 + left_non_all_zeros_count_108);
  assign left_all_zeros_count_111 = (all_left_zeros_192 & _zz_1371);
  assign _zz_347 = _zz_299[31 : 16];
  assign all_zeros_224 = ((! (_zz_347 != 16'h0)) ? 5'h1f : 5'h0);
  assign all_left_zeros_224 = ((! (_zz_347[15 : 8] != 8'h0)) ? 5'h1f : 5'h0);
  assign whole_bit_count_112 = 5'h10;
  assign left_bit_count_112 = 5'h08;
  assign _zz_348 = _zz_347[7 : 0];
  assign all_zeros_225 = ((! (_zz_348 != 8'h0)) ? 4'b1111 : 4'b0000);
  assign all_left_zeros_225 = ((! (_zz_348[7 : 4] != 4'b0000)) ? 4'b1111 : 4'b0000);
  assign whole_bit_count_113 = 4'b1000;
  assign left_bit_count_113 = 4'b0100;
  assign _zz_349 = _zz_348[3 : 0];
  assign all_zeros_226 = ((! (_zz_349 != 4'b0000)) ? 3'b111 : 3'b000);
  assign all_left_zeros_226 = ((! (_zz_349[3 : 2] != 2'b00)) ? 3'b111 : 3'b000);
  assign whole_bit_count_114 = 3'b100;
  assign left_bit_count_114 = 3'b010;
  assign _zz_350 = _zz_349[1 : 0];
  assign all_zeros_227 = ((! (_zz_350 != 2'b00)) ? 2'b11 : 2'b00);
  assign all_left_zeros_227 = ((! (_zz_350[1 : 1] != 1'b0)) ? 2'b11 : 2'b00);
  assign whole_bit_count_115 = 2'b10;
  assign left_bit_count_115 = 2'b01;
  assign _zz_351 = _zz_350[0 : 0];
  assign _zz_352 = _zz_351;
  assign all_zeros_228 = ((! (_zz_352 != 1'b0)) ? 1'b1 : 1'b0);
  assign all_left_zeros_228 = ((! (_zz_352[0 : 0] != 1'b0)) ? 1'b1 : 1'b0);
  assign left_all_zeros_count_112 = (all_left_zeros_227 & _zz_1375);
  assign _zz_353 = _zz_350[1 : 1];
  assign _zz_354 = _zz_353;
  assign all_zeros_229 = ((! (_zz_354 != 1'b0)) ? 1'b1 : 1'b0);
  assign all_left_zeros_229 = ((! (_zz_354[0 : 0] != 1'b0)) ? 1'b1 : 1'b0);
  assign left_non_all_zeros_count_109 = ((~ all_left_zeros_227) & _zz_1379);
  assign non_zeros_lzc_109 = (left_all_zeros_count_112 + left_non_all_zeros_count_109);
  assign left_all_zeros_count_113 = (all_left_zeros_226 & _zz_1380);
  assign _zz_355 = _zz_349[3 : 2];
  assign all_zeros_230 = ((! (_zz_355 != 2'b00)) ? 2'b11 : 2'b00);
  assign all_left_zeros_230 = ((! (_zz_355[1 : 1] != 1'b0)) ? 2'b11 : 2'b00);
  assign whole_bit_count_116 = 2'b10;
  assign left_bit_count_116 = 2'b01;
  assign _zz_356 = _zz_355[0 : 0];
  assign _zz_357 = _zz_356;
  assign all_zeros_231 = ((! (_zz_357 != 1'b0)) ? 1'b1 : 1'b0);
  assign all_left_zeros_231 = ((! (_zz_357[0 : 0] != 1'b0)) ? 1'b1 : 1'b0);
  assign left_all_zeros_count_114 = (all_left_zeros_230 & _zz_1384);
  assign _zz_358 = _zz_355[1 : 1];
  assign _zz_359 = _zz_358;
  assign all_zeros_232 = ((! (_zz_359 != 1'b0)) ? 1'b1 : 1'b0);
  assign all_left_zeros_232 = ((! (_zz_359[0 : 0] != 1'b0)) ? 1'b1 : 1'b0);
  assign left_non_all_zeros_count_110 = ((~ all_left_zeros_230) & _zz_1388);
  assign non_zeros_lzc_110 = (left_all_zeros_count_114 + left_non_all_zeros_count_110);
  assign left_non_all_zeros_count_111 = ((~ all_left_zeros_226) & _zz_1390);
  assign non_zeros_lzc_111 = (left_all_zeros_count_113 + left_non_all_zeros_count_111);
  assign left_all_zeros_count_115 = (all_left_zeros_225 & _zz_1392);
  assign _zz_360 = _zz_348[7 : 4];
  assign all_zeros_233 = ((! (_zz_360 != 4'b0000)) ? 3'b111 : 3'b000);
  assign all_left_zeros_233 = ((! (_zz_360[3 : 2] != 2'b00)) ? 3'b111 : 3'b000);
  assign whole_bit_count_117 = 3'b100;
  assign left_bit_count_117 = 3'b010;
  assign _zz_361 = _zz_360[1 : 0];
  assign all_zeros_234 = ((! (_zz_361 != 2'b00)) ? 2'b11 : 2'b00);
  assign all_left_zeros_234 = ((! (_zz_361[1 : 1] != 1'b0)) ? 2'b11 : 2'b00);
  assign whole_bit_count_118 = 2'b10;
  assign left_bit_count_118 = 2'b01;
  assign _zz_362 = _zz_361[0 : 0];
  assign _zz_363 = _zz_362;
  assign all_zeros_235 = ((! (_zz_363 != 1'b0)) ? 1'b1 : 1'b0);
  assign all_left_zeros_235 = ((! (_zz_363[0 : 0] != 1'b0)) ? 1'b1 : 1'b0);
  assign left_all_zeros_count_116 = (all_left_zeros_234 & _zz_1396);
  assign _zz_364 = _zz_361[1 : 1];
  assign _zz_365 = _zz_364;
  assign all_zeros_236 = ((! (_zz_365 != 1'b0)) ? 1'b1 : 1'b0);
  assign all_left_zeros_236 = ((! (_zz_365[0 : 0] != 1'b0)) ? 1'b1 : 1'b0);
  assign left_non_all_zeros_count_112 = ((~ all_left_zeros_234) & _zz_1400);
  assign non_zeros_lzc_112 = (left_all_zeros_count_116 + left_non_all_zeros_count_112);
  assign left_all_zeros_count_117 = (all_left_zeros_233 & _zz_1401);
  assign _zz_366 = _zz_360[3 : 2];
  assign all_zeros_237 = ((! (_zz_366 != 2'b00)) ? 2'b11 : 2'b00);
  assign all_left_zeros_237 = ((! (_zz_366[1 : 1] != 1'b0)) ? 2'b11 : 2'b00);
  assign whole_bit_count_119 = 2'b10;
  assign left_bit_count_119 = 2'b01;
  assign _zz_367 = _zz_366[0 : 0];
  assign _zz_368 = _zz_367;
  assign all_zeros_238 = ((! (_zz_368 != 1'b0)) ? 1'b1 : 1'b0);
  assign all_left_zeros_238 = ((! (_zz_368[0 : 0] != 1'b0)) ? 1'b1 : 1'b0);
  assign left_all_zeros_count_118 = (all_left_zeros_237 & _zz_1405);
  assign _zz_369 = _zz_366[1 : 1];
  assign _zz_370 = _zz_369;
  assign all_zeros_239 = ((! (_zz_370 != 1'b0)) ? 1'b1 : 1'b0);
  assign all_left_zeros_239 = ((! (_zz_370[0 : 0] != 1'b0)) ? 1'b1 : 1'b0);
  assign left_non_all_zeros_count_113 = ((~ all_left_zeros_237) & _zz_1409);
  assign non_zeros_lzc_113 = (left_all_zeros_count_118 + left_non_all_zeros_count_113);
  assign left_non_all_zeros_count_114 = ((~ all_left_zeros_233) & _zz_1411);
  assign non_zeros_lzc_114 = (left_all_zeros_count_117 + left_non_all_zeros_count_114);
  assign left_non_all_zeros_count_115 = ((~ all_left_zeros_225) & _zz_1414);
  assign non_zeros_lzc_115 = (left_all_zeros_count_115 + left_non_all_zeros_count_115);
  assign left_all_zeros_count_119 = (all_left_zeros_224 & _zz_1416);
  assign _zz_371 = _zz_347[15 : 8];
  assign all_zeros_240 = ((! (_zz_371 != 8'h0)) ? 4'b1111 : 4'b0000);
  assign all_left_zeros_240 = ((! (_zz_371[7 : 4] != 4'b0000)) ? 4'b1111 : 4'b0000);
  assign whole_bit_count_120 = 4'b1000;
  assign left_bit_count_120 = 4'b0100;
  assign _zz_372 = _zz_371[3 : 0];
  assign all_zeros_241 = ((! (_zz_372 != 4'b0000)) ? 3'b111 : 3'b000);
  assign all_left_zeros_241 = ((! (_zz_372[3 : 2] != 2'b00)) ? 3'b111 : 3'b000);
  assign whole_bit_count_121 = 3'b100;
  assign left_bit_count_121 = 3'b010;
  assign _zz_373 = _zz_372[1 : 0];
  assign all_zeros_242 = ((! (_zz_373 != 2'b00)) ? 2'b11 : 2'b00);
  assign all_left_zeros_242 = ((! (_zz_373[1 : 1] != 1'b0)) ? 2'b11 : 2'b00);
  assign whole_bit_count_122 = 2'b10;
  assign left_bit_count_122 = 2'b01;
  assign _zz_374 = _zz_373[0 : 0];
  assign _zz_375 = _zz_374;
  assign all_zeros_243 = ((! (_zz_375 != 1'b0)) ? 1'b1 : 1'b0);
  assign all_left_zeros_243 = ((! (_zz_375[0 : 0] != 1'b0)) ? 1'b1 : 1'b0);
  assign left_all_zeros_count_120 = (all_left_zeros_242 & _zz_1420);
  assign _zz_376 = _zz_373[1 : 1];
  assign _zz_377 = _zz_376;
  assign all_zeros_244 = ((! (_zz_377 != 1'b0)) ? 1'b1 : 1'b0);
  assign all_left_zeros_244 = ((! (_zz_377[0 : 0] != 1'b0)) ? 1'b1 : 1'b0);
  assign left_non_all_zeros_count_116 = ((~ all_left_zeros_242) & _zz_1424);
  assign non_zeros_lzc_116 = (left_all_zeros_count_120 + left_non_all_zeros_count_116);
  assign left_all_zeros_count_121 = (all_left_zeros_241 & _zz_1425);
  assign _zz_378 = _zz_372[3 : 2];
  assign all_zeros_245 = ((! (_zz_378 != 2'b00)) ? 2'b11 : 2'b00);
  assign all_left_zeros_245 = ((! (_zz_378[1 : 1] != 1'b0)) ? 2'b11 : 2'b00);
  assign whole_bit_count_123 = 2'b10;
  assign left_bit_count_123 = 2'b01;
  assign _zz_379 = _zz_378[0 : 0];
  assign _zz_380 = _zz_379;
  assign all_zeros_246 = ((! (_zz_380 != 1'b0)) ? 1'b1 : 1'b0);
  assign all_left_zeros_246 = ((! (_zz_380[0 : 0] != 1'b0)) ? 1'b1 : 1'b0);
  assign left_all_zeros_count_122 = (all_left_zeros_245 & _zz_1429);
  assign _zz_381 = _zz_378[1 : 1];
  assign _zz_382 = _zz_381;
  assign all_zeros_247 = ((! (_zz_382 != 1'b0)) ? 1'b1 : 1'b0);
  assign all_left_zeros_247 = ((! (_zz_382[0 : 0] != 1'b0)) ? 1'b1 : 1'b0);
  assign left_non_all_zeros_count_117 = ((~ all_left_zeros_245) & _zz_1433);
  assign non_zeros_lzc_117 = (left_all_zeros_count_122 + left_non_all_zeros_count_117);
  assign left_non_all_zeros_count_118 = ((~ all_left_zeros_241) & _zz_1435);
  assign non_zeros_lzc_118 = (left_all_zeros_count_121 + left_non_all_zeros_count_118);
  assign left_all_zeros_count_123 = (all_left_zeros_240 & _zz_1437);
  assign _zz_383 = _zz_371[7 : 4];
  assign all_zeros_248 = ((! (_zz_383 != 4'b0000)) ? 3'b111 : 3'b000);
  assign all_left_zeros_248 = ((! (_zz_383[3 : 2] != 2'b00)) ? 3'b111 : 3'b000);
  assign whole_bit_count_124 = 3'b100;
  assign left_bit_count_124 = 3'b010;
  assign _zz_384 = _zz_383[1 : 0];
  assign all_zeros_249 = ((! (_zz_384 != 2'b00)) ? 2'b11 : 2'b00);
  assign all_left_zeros_249 = ((! (_zz_384[1 : 1] != 1'b0)) ? 2'b11 : 2'b00);
  assign whole_bit_count_125 = 2'b10;
  assign left_bit_count_125 = 2'b01;
  assign _zz_385 = _zz_384[0 : 0];
  assign _zz_386 = _zz_385;
  assign all_zeros_250 = ((! (_zz_386 != 1'b0)) ? 1'b1 : 1'b0);
  assign all_left_zeros_250 = ((! (_zz_386[0 : 0] != 1'b0)) ? 1'b1 : 1'b0);
  assign left_all_zeros_count_124 = (all_left_zeros_249 & _zz_1441);
  assign _zz_387 = _zz_384[1 : 1];
  assign _zz_388 = _zz_387;
  assign all_zeros_251 = ((! (_zz_388 != 1'b0)) ? 1'b1 : 1'b0);
  assign all_left_zeros_251 = ((! (_zz_388[0 : 0] != 1'b0)) ? 1'b1 : 1'b0);
  assign left_non_all_zeros_count_119 = ((~ all_left_zeros_249) & _zz_1445);
  assign non_zeros_lzc_119 = (left_all_zeros_count_124 + left_non_all_zeros_count_119);
  assign left_all_zeros_count_125 = (all_left_zeros_248 & _zz_1446);
  assign _zz_389 = _zz_383[3 : 2];
  assign all_zeros_252 = ((! (_zz_389 != 2'b00)) ? 2'b11 : 2'b00);
  assign all_left_zeros_252 = ((! (_zz_389[1 : 1] != 1'b0)) ? 2'b11 : 2'b00);
  assign whole_bit_count_126 = 2'b10;
  assign left_bit_count_126 = 2'b01;
  assign _zz_390 = _zz_389[0 : 0];
  assign _zz_391 = _zz_390;
  assign all_zeros_253 = ((! (_zz_391 != 1'b0)) ? 1'b1 : 1'b0);
  assign all_left_zeros_253 = ((! (_zz_391[0 : 0] != 1'b0)) ? 1'b1 : 1'b0);
  assign left_all_zeros_count_126 = (all_left_zeros_252 & _zz_1450);
  assign _zz_392 = _zz_389[1 : 1];
  assign _zz_393 = _zz_392;
  assign all_zeros_254 = ((! (_zz_393 != 1'b0)) ? 1'b1 : 1'b0);
  assign all_left_zeros_254 = ((! (_zz_393[0 : 0] != 1'b0)) ? 1'b1 : 1'b0);
  assign left_non_all_zeros_count_120 = ((~ all_left_zeros_252) & _zz_1454);
  assign non_zeros_lzc_120 = (left_all_zeros_count_126 + left_non_all_zeros_count_120);
  assign left_non_all_zeros_count_121 = ((~ all_left_zeros_248) & _zz_1456);
  assign non_zeros_lzc_121 = (left_all_zeros_count_125 + left_non_all_zeros_count_121);
  assign left_non_all_zeros_count_122 = ((~ all_left_zeros_240) & _zz_1459);
  assign non_zeros_lzc_122 = (left_all_zeros_count_123 + left_non_all_zeros_count_122);
  assign left_non_all_zeros_count_123 = ((~ all_left_zeros_224) & _zz_1462);
  assign non_zeros_lzc_123 = (left_all_zeros_count_119 + left_non_all_zeros_count_123);
  assign left_non_all_zeros_count_124 = ((~ all_left_zeros_192) & _zz_1465);
  assign non_zeros_lzc_124 = (left_all_zeros_count_111 + left_non_all_zeros_count_124);
  assign left_non_all_zeros_count_125 = ((~ all_left_zeros_128) & _zz_1468);
  assign non_zeros_lzc_125 = (left_all_zeros_count_95 + left_non_all_zeros_count_125);
  assign left_non_all_zeros_count_126 = ((~ all_left_zeros) & _zz_1471);
  assign non_zeros_lzc_126 = (left_all_zeros_count_63 + left_non_all_zeros_count_126);
  assign lzc = _zz_394[6:0];
  assign _zz_395 = (lzc - 7'h01);
  assign _zz_396 = _zz_1475[7 : 0];
  assign _zz_397 = _zz_448;
  assign _zz_398 = _zz_449;
  assign _zz_399 = ($signed(_zz_396) - $signed(_zz_1476));
  assign _zz_413 = ($signed(_zz_397) - $signed(_zz_451));
  assign _zz_414 = ($signed(_zz_398) - $signed(_zz_452));
  assign _zz_415 = _zz_1478;
  assign _zz_416 = _zz_399;
  assign _zz_400 = {{8{_zz_1480[7]}}, _zz_1480};
  assign _zz_417 = _zz_1481;
  assign _zz_418 = _zz_399;
  assign _zz_401 = {{8{_zz_1483[7]}}, _zz_1483};
  assign _zz_402 = ($signed(wd_prod) - $signed(_zz_396));
  assign _zz_403 = 8'h0;
  assign _zz_419 = ($signed(_zz_400) + $signed(_zz_401));
  assign _zz_420 = _zz_1484;
  assign _zz_421 = _zz_1486;
  assign _zz_422 = mulUnit_1_c[15 : 0];
  assign _zz_404 = _zz_1488[15 : 0];
  assign _zz_423 = ($signed(_zz_403) - $signed(_zz_402));
  assign _zz_424 = _zz_1489;
  assign _zz_425 = _zz_1491;
  assign _zz_426 = mulUnit_2_c[15 : 0];
  assign _zz_427 = ($signed(_zz_402) + $signed(_zz_403));
  assign _zz_428 = _zz_1493;
  assign _zz_429 = _zz_1495;
  assign _zz_430 = mulUnit_3_c[15 : 0];
  always @ (*) begin
    if(_zz_453)begin
      exp_wd_prod_real = _zz_405;
    end else begin
      if(_zz_454)begin
        exp_wd_prod_real = {{8{_zz_1511[23]}}, _zz_1511};
      end else begin
        exp_wd_prod_real = {{8{_zz_1513[23]}}, _zz_1513};
      end
    end
  end

  always @ (*) begin
    if(_zz_453)begin
      exp_wd_prod_imag = _zz_406;
    end else begin
      if(_zz_454)begin
        exp_wd_prod_imag = {{8{_zz_1512[23]}}, _zz_1512};
      end else begin
        exp_wd_prod_imag = {{8{_zz_1514[23]}}, _zz_1514};
      end
    end
  end

  assign _zz_407 = _zz_409;
  assign _zz_431 = _zz_1515;
  assign _zz_432 = _zz_407;
  assign _zz_433 = _zz_1517;
  assign _zz_434 = _zz_407;
  assign _zz_435 = ($signed(exp_wd_prod_divw_real) + $signed(exp_wd_prod_divw_imag));
  assign _zz_436 = _zz_1523;
  assign _zz_437 = _zz_1525;
  assign _zz_438 = mulUnit_4_c[31 : 0];
  assign _zz_410 = _zz_1527[31 : 0];
  assign _zz_439 = ($signed(timeshift_imag) - $signed(timeshift_real));
  assign _zz_440 = _zz_1528;
  assign _zz_441 = _zz_1530;
  assign _zz_442 = mulUnit_5_c[31 : 0];
  assign _zz_443 = ($signed(timeshift_real) + $signed(timeshift_imag));
  assign _zz_444 = _zz_1532;
  assign _zz_445 = _zz_1534;
  assign _zz_446 = mulUnit_6_c[31 : 0];
  assign io_coef_real = _zz_1544[15 : 0];
  assign io_coef_imag = _zz_1545[15 : 0];
  always @ (posedge clk) begin
    wave <= io_wave;
    distance <= io_distance;
    io_timeshift_regNext_real <= io_timeshift_real;
    io_timeshift_regNext_imag <= io_timeshift_imag;
    _zz_1 <= io_timeshift_regNext_real;
    _zz_2 <= io_timeshift_regNext_imag;
    _zz_3 <= _zz_1;
    _zz_4 <= _zz_2;
    _zz_5 <= _zz_3;
    _zz_6 <= _zz_4;
    _zz_7 <= _zz_5;
    _zz_8 <= _zz_6;
    _zz_9 <= ($signed(wave) * $signed(distance));
    _zz_394 <= ((all_zeros & _zz_1473) & non_zeros_lzc_126);
    wave_regNext <= wave;
    _zz_408 <= wave_regNext;
    _zz_409 <= _zz_408;
    exp_wd_prod_divw_real <= {{8{_zz_1519[23]}}, _zz_1519};
    exp_wd_prod_divw_imag <= {{8{_zz_1521[23]}}, _zz_1521};
    _zz_411 <= {{16{_zz_1536[47]}}, _zz_1536};
    _zz_412 <= {{16{_zz_1540[47]}}, _zz_1540};
  end

  always @ (posedge clk) begin
    _zz_405 <= ($signed(_zz_1498) + $signed(_zz_1503));
    _zz_406 <= ($signed(_zz_1505) + $signed(_zz_1510));
  end

  always @ (posedge clk) begin
    func_table_0_regNext_real <= func_table_0_real;
    func_table_0_regNext_imag <= func_table_0_imag;
  end

  always @ (posedge clk) begin
    func_table_127_regNext_real <= func_table_127_real;
    func_table_127_regNext_imag <= func_table_127_imag;
  end


endmodule

//SInt64fixTo39_24_ROUNDTOINF replaced by SInt64fixTo39_24_ROUNDTOINF

module SInt64fixTo39_24_ROUNDTOINF (
  input      [63:0]   din,
  output     [15:0]   dout
);
  wire       [64:0]   _zz_9;
  wire       [64:0]   _zz_10;
  wire       [23:0]   _zz_11;
  wire       [40:0]   _zz_12;
  wire       [40:0]   _zz_13;
  wire       [64:0]   _zz_14;
  wire       [64:0]   _zz_15;
  wire       [64:0]   _zz_16;
  wire       [25:0]   _zz_17;
  wire       [24:0]   _zz_18;
  reg        [40:0]   _zz_1;
  wire       [63:0]   _zz_2;
  wire       [63:0]   _zz_3;
  wire       [63:0]   _zz_4;
  wire       [64:0]   _zz_5;
  wire       [63:0]   _zz_6;
  reg        [40:0]   _zz_7;
  reg        [15:0]   _zz_8;

  assign _zz_9 = {_zz_4[63],_zz_4};
  assign _zz_10 = {_zz_3[63],_zz_3};
  assign _zz_11 = _zz_5[23 : 0];
  assign _zz_12 = _zz_5[64 : 24];
  assign _zz_13 = 41'h00000000001;
  assign _zz_14 = ($signed(_zz_15) + $signed(_zz_16));
  assign _zz_15 = {_zz_6[63],_zz_6};
  assign _zz_16 = {_zz_2[63],_zz_2};
  assign _zz_17 = _zz_1[40 : 15];
  assign _zz_18 = _zz_1[39 : 15];
  assign _zz_2 = {{40'h0,1'b1},23'h0};
  assign _zz_3 = {41'h1ffffffffff,23'h0};
  assign _zz_4 = din[63 : 0];
  assign _zz_5 = ($signed(_zz_9) + $signed(_zz_10));
  assign _zz_6 = din[63 : 0];
  always @ (*) begin
    if((_zz_11 != 24'h0))begin
      _zz_7 = ($signed(_zz_12) + $signed(_zz_13));
    end else begin
      _zz_7 = _zz_5[64 : 24];
    end
  end

  always @ (*) begin
    if(_zz_5[64])begin
      _zz_1 = _zz_7;
    end else begin
      _zz_1 = (_zz_14 >>> 24);
    end
  end

  always @ (*) begin
    if(_zz_1[40])begin
      if((! (_zz_17 == 26'h3ffffff)))begin
        _zz_8 = 16'h8000;
      end else begin
        _zz_8 = _zz_1[15 : 0];
      end
    end else begin
      if((_zz_18 != 25'h0))begin
        _zz_8 = 16'h7fff;
      end else begin
        _zz_8 = _zz_1[15 : 0];
      end
    end
  end

  assign dout = _zz_8;

endmodule

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt16fixTo31_0_ROUNDTOINF replaced by SInt16fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

//SInt16fixTo31_0_ROUNDTOINF replaced by SInt16fixTo31_0_ROUNDTOINF

//SInt32fixTo31_0_ROUNDTOINF replaced by SInt32fixTo31_0_ROUNDTOINF

module SInt16fixTo31_0_ROUNDTOINF (
  input      [15:0]   din,
  output     [31:0]   dout
);
  wire                _zz_1;
  wire       [0:0]    _zz_2;
  wire       [5:0]    _zz_3;

  assign _zz_1 = din[15];
  assign _zz_2 = din[15];
  assign _zz_3 = {din[15],{din[15],{din[15],{din[15],{din[15],din[15]}}}}};
  assign dout = {{din[15],{din[15],{din[15],{din[15],{din[15],{din[15],{din[15],{din[15],{_zz_1,{_zz_2,_zz_3}}}}}}}}}},din};

endmodule

module SInt32fixTo31_0_ROUNDTOINF (
  input      [31:0]   din,
  output     [31:0]   dout
);

  assign dout = din;

endmodule

//SInt32fixTo23_8_ROUNDTOINF replaced by SInt32fixTo23_8_ROUNDTOINF

module SInt32fixTo23_8_ROUNDTOINF (
  input      [31:0]   din,
  output     [15:0]   dout
);
  wire       [32:0]   _zz_9;
  wire       [32:0]   _zz_10;
  wire       [7:0]    _zz_11;
  wire       [24:0]   _zz_12;
  wire       [24:0]   _zz_13;
  wire       [32:0]   _zz_14;
  wire       [32:0]   _zz_15;
  wire       [32:0]   _zz_16;
  wire       [9:0]    _zz_17;
  wire       [8:0]    _zz_18;
  reg        [24:0]   _zz_1;
  wire       [31:0]   _zz_2;
  wire       [31:0]   _zz_3;
  wire       [31:0]   _zz_4;
  wire       [32:0]   _zz_5;
  wire       [31:0]   _zz_6;
  reg        [24:0]   _zz_7;
  reg        [15:0]   _zz_8;

  assign _zz_9 = {_zz_4[31],_zz_4};
  assign _zz_10 = {_zz_3[31],_zz_3};
  assign _zz_11 = _zz_5[7 : 0];
  assign _zz_12 = _zz_5[32 : 8];
  assign _zz_13 = 25'h0000001;
  assign _zz_14 = ($signed(_zz_15) + $signed(_zz_16));
  assign _zz_15 = {_zz_6[31],_zz_6};
  assign _zz_16 = {_zz_2[31],_zz_2};
  assign _zz_17 = _zz_1[24 : 15];
  assign _zz_18 = _zz_1[23 : 15];
  assign _zz_2 = {{24'h0,1'b1},7'h0};
  assign _zz_3 = {25'h1ffffff,7'h0};
  assign _zz_4 = din[31 : 0];
  assign _zz_5 = ($signed(_zz_9) + $signed(_zz_10));
  assign _zz_6 = din[31 : 0];
  always @ (*) begin
    if((_zz_11 != 8'h0))begin
      _zz_7 = ($signed(_zz_12) + $signed(_zz_13));
    end else begin
      _zz_7 = _zz_5[32 : 8];
    end
  end

  always @ (*) begin
    if(_zz_5[32])begin
      _zz_1 = _zz_7;
    end else begin
      _zz_1 = (_zz_14 >>> 8);
    end
  end

  always @ (*) begin
    if(_zz_1[24])begin
      if((! (_zz_17 == 10'h3ff)))begin
        _zz_8 = 16'h8000;
      end else begin
        _zz_8 = _zz_1[15 : 0];
      end
    end else begin
      if((_zz_18 != 9'h0))begin
        _zz_8 = 16'h7fff;
      end else begin
        _zz_8 = _zz_1[15 : 0];
      end
    end
  end

  assign dout = _zz_8;

endmodule

//SInt16fixTo15_0_ROUNDTOINF replaced by SInt16fixTo15_0_ROUNDTOINF

//SInt16fixTo15_0_ROUNDTOINF replaced by SInt16fixTo15_0_ROUNDTOINF

//SInt8fixTo15_0_ROUNDTOINF replaced by SInt8fixTo15_0_ROUNDTOINF

//SInt16fixTo15_0_ROUNDTOINF replaced by SInt16fixTo15_0_ROUNDTOINF

//SInt16fixTo15_0_ROUNDTOINF replaced by SInt16fixTo15_0_ROUNDTOINF

//SInt8fixTo15_0_ROUNDTOINF replaced by SInt8fixTo15_0_ROUNDTOINF

//SInt16fixTo15_0_ROUNDTOINF replaced by SInt16fixTo15_0_ROUNDTOINF

module SInt8fixTo15_0_ROUNDTOINF (
  input      [7:0]    din,
  output     [15:0]   dout
);

  assign dout = {{din[7],{din[7],{din[7],{din[7],{din[7],{din[7],{din[7],din[7]}}}}}}},din};

endmodule

module SInt16fixTo15_0_ROUNDTOINF (
  input      [15:0]   din,
  output     [15:0]   dout
);

  assign dout = din;

endmodule

//SInt16fixTo7_0_ROUNDTOINF replaced by SInt16fixTo7_0_ROUNDTOINF

module SInt16fixTo7_0_ROUNDTOINF (
  input      [15:0]   din,
  output     [7:0]    dout
);
  wire       [8:0]    _zz_2;
  wire       [7:0]    _zz_3;
  reg        [7:0]    _zz_1;

  assign _zz_2 = din[15 : 7];
  assign _zz_3 = din[14 : 7];
  always @ (*) begin
    if(din[15])begin
      if((! (_zz_2 == 9'h1ff)))begin
        _zz_1 = 8'h80;
      end else begin
        _zz_1 = din[7 : 0];
      end
    end else begin
      if((_zz_3 != 8'h0))begin
        _zz_1 = 8'h7f;
      end else begin
        _zz_1 = din[7 : 0];
      end
    end
  end

  assign dout = _zz_1;

endmodule

module SInt32fixTo15_8_ROUNDTOINF (
  input      [31:0]   din,
  output     [7:0]    dout
);
  wire       [32:0]   _zz_9;
  wire       [32:0]   _zz_10;
  wire       [7:0]    _zz_11;
  wire       [24:0]   _zz_12;
  wire       [24:0]   _zz_13;
  wire       [32:0]   _zz_14;
  wire       [32:0]   _zz_15;
  wire       [32:0]   _zz_16;
  wire       [17:0]   _zz_17;
  wire       [16:0]   _zz_18;
  reg        [24:0]   _zz_1;
  wire       [31:0]   _zz_2;
  wire       [31:0]   _zz_3;
  wire       [31:0]   _zz_4;
  wire       [32:0]   _zz_5;
  wire       [31:0]   _zz_6;
  reg        [24:0]   _zz_7;
  reg        [7:0]    _zz_8;

  assign _zz_9 = {_zz_4[31],_zz_4};
  assign _zz_10 = {_zz_3[31],_zz_3};
  assign _zz_11 = _zz_5[7 : 0];
  assign _zz_12 = _zz_5[32 : 8];
  assign _zz_13 = 25'h0000001;
  assign _zz_14 = ($signed(_zz_15) + $signed(_zz_16));
  assign _zz_15 = {_zz_6[31],_zz_6};
  assign _zz_16 = {_zz_2[31],_zz_2};
  assign _zz_17 = _zz_1[24 : 7];
  assign _zz_18 = _zz_1[23 : 7];
  assign _zz_2 = {{24'h0,1'b1},7'h0};
  assign _zz_3 = {25'h1ffffff,7'h0};
  assign _zz_4 = din[31 : 0];
  assign _zz_5 = ($signed(_zz_9) + $signed(_zz_10));
  assign _zz_6 = din[31 : 0];
  always @ (*) begin
    if((_zz_11 != 8'h0))begin
      _zz_7 = ($signed(_zz_12) + $signed(_zz_13));
    end else begin
      _zz_7 = _zz_5[32 : 8];
    end
  end

  always @ (*) begin
    if(_zz_5[32])begin
      _zz_1 = _zz_7;
    end else begin
      _zz_1 = (_zz_14 >>> 8);
    end
  end

  always @ (*) begin
    if(_zz_1[24])begin
      if((! (_zz_17 == 18'h3ffff)))begin
        _zz_8 = 8'h80;
      end else begin
        _zz_8 = _zz_1[7 : 0];
      end
    end else begin
      if((_zz_18 != 17'h0))begin
        _zz_8 = 8'h7f;
      end else begin
        _zz_8 = _zz_1[7 : 0];
      end
    end
  end

  assign dout = _zz_8;

endmodule
