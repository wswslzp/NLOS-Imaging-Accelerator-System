// Generator : SpinalHDL v1.4.1    git head : d1b4746673438bc5f242515335278fa39a666c38
// Component : Lzc
// Git hash  : 2a34fe18f42a28946060dbf37f9913e1060dc674



module Lzc (
  input      [15:0]   a,
  output     [15:0]   a_lzc
);
  wire       [1:0]    _zz_48;
  wire       [0:0]    _zz_49;
  wire       [1:0]    _zz_50;
  wire       [0:0]    _zz_51;
  wire       [1:0]    _zz_52;
  wire       [2:0]    _zz_53;
  wire       [1:0]    _zz_54;
  wire       [2:0]    _zz_55;
  wire       [1:0]    _zz_56;
  wire       [1:0]    _zz_57;
  wire       [0:0]    _zz_58;
  wire       [1:0]    _zz_59;
  wire       [0:0]    _zz_60;
  wire       [1:0]    _zz_61;
  wire       [1:0]    _zz_62;
  wire       [2:0]    _zz_63;
  wire       [1:0]    _zz_64;
  wire       [3:0]    _zz_65;
  wire       [2:0]    _zz_66;
  wire       [3:0]    _zz_67;
  wire       [2:0]    _zz_68;
  wire       [1:0]    _zz_69;
  wire       [0:0]    _zz_70;
  wire       [1:0]    _zz_71;
  wire       [0:0]    _zz_72;
  wire       [1:0]    _zz_73;
  wire       [2:0]    _zz_74;
  wire       [1:0]    _zz_75;
  wire       [2:0]    _zz_76;
  wire       [1:0]    _zz_77;
  wire       [1:0]    _zz_78;
  wire       [0:0]    _zz_79;
  wire       [1:0]    _zz_80;
  wire       [0:0]    _zz_81;
  wire       [1:0]    _zz_82;
  wire       [1:0]    _zz_83;
  wire       [2:0]    _zz_84;
  wire       [1:0]    _zz_85;
  wire       [2:0]    _zz_86;
  wire       [3:0]    _zz_87;
  wire       [2:0]    _zz_88;
  wire       [4:0]    _zz_89;
  wire       [3:0]    _zz_90;
  wire       [4:0]    _zz_91;
  wire       [3:0]    _zz_92;
  wire       [1:0]    _zz_93;
  wire       [0:0]    _zz_94;
  wire       [1:0]    _zz_95;
  wire       [0:0]    _zz_96;
  wire       [1:0]    _zz_97;
  wire       [2:0]    _zz_98;
  wire       [1:0]    _zz_99;
  wire       [2:0]    _zz_100;
  wire       [1:0]    _zz_101;
  wire       [1:0]    _zz_102;
  wire       [0:0]    _zz_103;
  wire       [1:0]    _zz_104;
  wire       [0:0]    _zz_105;
  wire       [1:0]    _zz_106;
  wire       [1:0]    _zz_107;
  wire       [2:0]    _zz_108;
  wire       [1:0]    _zz_109;
  wire       [3:0]    _zz_110;
  wire       [2:0]    _zz_111;
  wire       [3:0]    _zz_112;
  wire       [2:0]    _zz_113;
  wire       [1:0]    _zz_114;
  wire       [0:0]    _zz_115;
  wire       [1:0]    _zz_116;
  wire       [0:0]    _zz_117;
  wire       [1:0]    _zz_118;
  wire       [2:0]    _zz_119;
  wire       [1:0]    _zz_120;
  wire       [2:0]    _zz_121;
  wire       [1:0]    _zz_122;
  wire       [1:0]    _zz_123;
  wire       [0:0]    _zz_124;
  wire       [1:0]    _zz_125;
  wire       [0:0]    _zz_126;
  wire       [1:0]    _zz_127;
  wire       [1:0]    _zz_128;
  wire       [2:0]    _zz_129;
  wire       [1:0]    _zz_130;
  wire       [2:0]    _zz_131;
  wire       [3:0]    _zz_132;
  wire       [2:0]    _zz_133;
  wire       [3:0]    _zz_134;
  wire       [4:0]    _zz_135;
  wire       [3:0]    _zz_136;
  wire       [4:0]    _zz_137;
  wire       [4:0]    _zz_138;
  wire       [15:0]   _zz_1;
  wire       [4:0]    all_zeros;
  wire       [4:0]    all_left_zeros;
  wire       [4:0]    whole_bit_count;
  wire       [4:0]    left_bit_count;
  wire       [7:0]    _zz_2;
  wire       [3:0]    all_zeros_1;
  wire       [3:0]    all_left_zeros_1;
  wire       [3:0]    whole_bit_count_1;
  wire       [3:0]    left_bit_count_1;
  wire       [3:0]    _zz_3;
  wire       [2:0]    all_zeros_2;
  wire       [2:0]    all_left_zeros_2;
  wire       [2:0]    whole_bit_count_2;
  wire       [2:0]    left_bit_count_2;
  wire       [1:0]    _zz_4;
  wire       [1:0]    all_zeros_3;
  wire       [1:0]    all_left_zeros_3;
  wire       [1:0]    whole_bit_count_3;
  wire       [1:0]    left_bit_count_3;
  wire       [0:0]    _zz_5;
  wire       [0:0]    _zz_6;
  wire       [0:0]    all_zeros_4;
  wire       [0:0]    all_left_zeros_4;
  wire       [1:0]    left_all_zeros_count;
  wire       [0:0]    _zz_7;
  wire       [0:0]    _zz_8;
  wire       [0:0]    all_zeros_5;
  wire       [0:0]    all_left_zeros_5;
  wire       [1:0]    left_non_all_zeros_count;
  wire       [1:0]    non_zeros_lzc;
  wire       [2:0]    left_all_zeros_count_1;
  wire       [1:0]    _zz_9;
  wire       [1:0]    all_zeros_6;
  wire       [1:0]    all_left_zeros_6;
  wire       [1:0]    whole_bit_count_4;
  wire       [1:0]    left_bit_count_4;
  wire       [0:0]    _zz_10;
  wire       [0:0]    _zz_11;
  wire       [0:0]    all_zeros_7;
  wire       [0:0]    all_left_zeros_7;
  wire       [1:0]    left_all_zeros_count_2;
  wire       [0:0]    _zz_12;
  wire       [0:0]    _zz_13;
  wire       [0:0]    all_zeros_8;
  wire       [0:0]    all_left_zeros_8;
  wire       [1:0]    left_non_all_zeros_count_1;
  wire       [1:0]    non_zeros_lzc_1;
  wire       [2:0]    left_non_all_zeros_count_2;
  wire       [2:0]    non_zeros_lzc_2;
  wire       [3:0]    left_all_zeros_count_3;
  wire       [3:0]    _zz_14;
  wire       [2:0]    all_zeros_9;
  wire       [2:0]    all_left_zeros_9;
  wire       [2:0]    whole_bit_count_5;
  wire       [2:0]    left_bit_count_5;
  wire       [1:0]    _zz_15;
  wire       [1:0]    all_zeros_10;
  wire       [1:0]    all_left_zeros_10;
  wire       [1:0]    whole_bit_count_6;
  wire       [1:0]    left_bit_count_6;
  wire       [0:0]    _zz_16;
  wire       [0:0]    _zz_17;
  wire       [0:0]    all_zeros_11;
  wire       [0:0]    all_left_zeros_11;
  wire       [1:0]    left_all_zeros_count_4;
  wire       [0:0]    _zz_18;
  wire       [0:0]    _zz_19;
  wire       [0:0]    all_zeros_12;
  wire       [0:0]    all_left_zeros_12;
  wire       [1:0]    left_non_all_zeros_count_3;
  wire       [1:0]    non_zeros_lzc_3;
  wire       [2:0]    left_all_zeros_count_5;
  wire       [1:0]    _zz_20;
  wire       [1:0]    all_zeros_13;
  wire       [1:0]    all_left_zeros_13;
  wire       [1:0]    whole_bit_count_7;
  wire       [1:0]    left_bit_count_7;
  wire       [0:0]    _zz_21;
  wire       [0:0]    _zz_22;
  wire       [0:0]    all_zeros_14;
  wire       [0:0]    all_left_zeros_14;
  wire       [1:0]    left_all_zeros_count_6;
  wire       [0:0]    _zz_23;
  wire       [0:0]    _zz_24;
  wire       [0:0]    all_zeros_15;
  wire       [0:0]    all_left_zeros_15;
  wire       [1:0]    left_non_all_zeros_count_4;
  wire       [1:0]    non_zeros_lzc_4;
  wire       [2:0]    left_non_all_zeros_count_5;
  wire       [2:0]    non_zeros_lzc_5;
  wire       [3:0]    left_non_all_zeros_count_6;
  wire       [3:0]    non_zeros_lzc_6;
  wire       [4:0]    left_all_zeros_count_7;
  wire       [7:0]    _zz_25;
  wire       [3:0]    all_zeros_16;
  wire       [3:0]    all_left_zeros_16;
  wire       [3:0]    whole_bit_count_8;
  wire       [3:0]    left_bit_count_8;
  wire       [3:0]    _zz_26;
  wire       [2:0]    all_zeros_17;
  wire       [2:0]    all_left_zeros_17;
  wire       [2:0]    whole_bit_count_9;
  wire       [2:0]    left_bit_count_9;
  wire       [1:0]    _zz_27;
  wire       [1:0]    all_zeros_18;
  wire       [1:0]    all_left_zeros_18;
  wire       [1:0]    whole_bit_count_10;
  wire       [1:0]    left_bit_count_10;
  wire       [0:0]    _zz_28;
  wire       [0:0]    _zz_29;
  wire       [0:0]    all_zeros_19;
  wire       [0:0]    all_left_zeros_19;
  wire       [1:0]    left_all_zeros_count_8;
  wire       [0:0]    _zz_30;
  wire       [0:0]    _zz_31;
  wire       [0:0]    all_zeros_20;
  wire       [0:0]    all_left_zeros_20;
  wire       [1:0]    left_non_all_zeros_count_7;
  wire       [1:0]    non_zeros_lzc_7;
  wire       [2:0]    left_all_zeros_count_9;
  wire       [1:0]    _zz_32;
  wire       [1:0]    all_zeros_21;
  wire       [1:0]    all_left_zeros_21;
  wire       [1:0]    whole_bit_count_11;
  wire       [1:0]    left_bit_count_11;
  wire       [0:0]    _zz_33;
  wire       [0:0]    _zz_34;
  wire       [0:0]    all_zeros_22;
  wire       [0:0]    all_left_zeros_22;
  wire       [1:0]    left_all_zeros_count_10;
  wire       [0:0]    _zz_35;
  wire       [0:0]    _zz_36;
  wire       [0:0]    all_zeros_23;
  wire       [0:0]    all_left_zeros_23;
  wire       [1:0]    left_non_all_zeros_count_8;
  wire       [1:0]    non_zeros_lzc_8;
  wire       [2:0]    left_non_all_zeros_count_9;
  wire       [2:0]    non_zeros_lzc_9;
  wire       [3:0]    left_all_zeros_count_11;
  wire       [3:0]    _zz_37;
  wire       [2:0]    all_zeros_24;
  wire       [2:0]    all_left_zeros_24;
  wire       [2:0]    whole_bit_count_12;
  wire       [2:0]    left_bit_count_12;
  wire       [1:0]    _zz_38;
  wire       [1:0]    all_zeros_25;
  wire       [1:0]    all_left_zeros_25;
  wire       [1:0]    whole_bit_count_13;
  wire       [1:0]    left_bit_count_13;
  wire       [0:0]    _zz_39;
  wire       [0:0]    _zz_40;
  wire       [0:0]    all_zeros_26;
  wire       [0:0]    all_left_zeros_26;
  wire       [1:0]    left_all_zeros_count_12;
  wire       [0:0]    _zz_41;
  wire       [0:0]    _zz_42;
  wire       [0:0]    all_zeros_27;
  wire       [0:0]    all_left_zeros_27;
  wire       [1:0]    left_non_all_zeros_count_10;
  wire       [1:0]    non_zeros_lzc_10;
  wire       [2:0]    left_all_zeros_count_13;
  wire       [1:0]    _zz_43;
  wire       [1:0]    all_zeros_28;
  wire       [1:0]    all_left_zeros_28;
  wire       [1:0]    whole_bit_count_14;
  wire       [1:0]    left_bit_count_14;
  wire       [0:0]    _zz_44;
  wire       [0:0]    _zz_45;
  wire       [0:0]    all_zeros_29;
  wire       [0:0]    all_left_zeros_29;
  wire       [1:0]    left_all_zeros_count_14;
  wire       [0:0]    _zz_46;
  wire       [0:0]    _zz_47;
  wire       [0:0]    all_zeros_30;
  wire       [0:0]    all_left_zeros_30;
  wire       [1:0]    left_non_all_zeros_count_11;
  wire       [1:0]    non_zeros_lzc_11;
  wire       [2:0]    left_non_all_zeros_count_12;
  wire       [2:0]    non_zeros_lzc_12;
  wire       [3:0]    left_non_all_zeros_count_13;
  wire       [3:0]    non_zeros_lzc_13;
  wire       [4:0]    left_non_all_zeros_count_14;
  wire       [4:0]    non_zeros_lzc_14;

  assign _zz_48 = (left_bit_count_3 + _zz_50);
  assign _zz_49 = _zz_5[0];
  assign _zz_50 = {1'd0, _zz_49};
  assign _zz_51 = _zz_7[0];
  assign _zz_52 = {1'd0, _zz_51};
  assign _zz_53 = (left_bit_count_2 + _zz_55);
  assign _zz_54 = ((all_zeros_3 & _zz_56) & non_zeros_lzc);
  assign _zz_55 = {1'd0, _zz_54};
  assign _zz_56 = (whole_bit_count_3 + (~ all_zeros_3));
  assign _zz_57 = (left_bit_count_4 + _zz_59);
  assign _zz_58 = _zz_10[0];
  assign _zz_59 = {1'd0, _zz_58};
  assign _zz_60 = _zz_12[0];
  assign _zz_61 = {1'd0, _zz_60};
  assign _zz_62 = ((all_zeros_6 & _zz_64) & non_zeros_lzc_1);
  assign _zz_63 = {1'd0, _zz_62};
  assign _zz_64 = (whole_bit_count_4 + (~ all_zeros_6));
  assign _zz_65 = (left_bit_count_1 + _zz_67);
  assign _zz_66 = ((all_zeros_2 & _zz_68) & non_zeros_lzc_2);
  assign _zz_67 = {1'd0, _zz_66};
  assign _zz_68 = (whole_bit_count_2 + (~ all_zeros_2));
  assign _zz_69 = (left_bit_count_6 + _zz_71);
  assign _zz_70 = _zz_16[0];
  assign _zz_71 = {1'd0, _zz_70};
  assign _zz_72 = _zz_18[0];
  assign _zz_73 = {1'd0, _zz_72};
  assign _zz_74 = (left_bit_count_5 + _zz_76);
  assign _zz_75 = ((all_zeros_10 & _zz_77) & non_zeros_lzc_3);
  assign _zz_76 = {1'd0, _zz_75};
  assign _zz_77 = (whole_bit_count_6 + (~ all_zeros_10));
  assign _zz_78 = (left_bit_count_7 + _zz_80);
  assign _zz_79 = _zz_21[0];
  assign _zz_80 = {1'd0, _zz_79};
  assign _zz_81 = _zz_23[0];
  assign _zz_82 = {1'd0, _zz_81};
  assign _zz_83 = ((all_zeros_13 & _zz_85) & non_zeros_lzc_4);
  assign _zz_84 = {1'd0, _zz_83};
  assign _zz_85 = (whole_bit_count_7 + (~ all_zeros_13));
  assign _zz_86 = ((all_zeros_9 & _zz_88) & non_zeros_lzc_5);
  assign _zz_87 = {1'd0, _zz_86};
  assign _zz_88 = (whole_bit_count_5 + (~ all_zeros_9));
  assign _zz_89 = (left_bit_count + _zz_91);
  assign _zz_90 = ((all_zeros_1 & _zz_92) & non_zeros_lzc_6);
  assign _zz_91 = {1'd0, _zz_90};
  assign _zz_92 = (whole_bit_count_1 + (~ all_zeros_1));
  assign _zz_93 = (left_bit_count_10 + _zz_95);
  assign _zz_94 = _zz_28[0];
  assign _zz_95 = {1'd0, _zz_94};
  assign _zz_96 = _zz_30[0];
  assign _zz_97 = {1'd0, _zz_96};
  assign _zz_98 = (left_bit_count_9 + _zz_100);
  assign _zz_99 = ((all_zeros_18 & _zz_101) & non_zeros_lzc_7);
  assign _zz_100 = {1'd0, _zz_99};
  assign _zz_101 = (whole_bit_count_10 + (~ all_zeros_18));
  assign _zz_102 = (left_bit_count_11 + _zz_104);
  assign _zz_103 = _zz_33[0];
  assign _zz_104 = {1'd0, _zz_103};
  assign _zz_105 = _zz_35[0];
  assign _zz_106 = {1'd0, _zz_105};
  assign _zz_107 = ((all_zeros_21 & _zz_109) & non_zeros_lzc_8);
  assign _zz_108 = {1'd0, _zz_107};
  assign _zz_109 = (whole_bit_count_11 + (~ all_zeros_21));
  assign _zz_110 = (left_bit_count_8 + _zz_112);
  assign _zz_111 = ((all_zeros_17 & _zz_113) & non_zeros_lzc_9);
  assign _zz_112 = {1'd0, _zz_111};
  assign _zz_113 = (whole_bit_count_9 + (~ all_zeros_17));
  assign _zz_114 = (left_bit_count_13 + _zz_116);
  assign _zz_115 = _zz_39[0];
  assign _zz_116 = {1'd0, _zz_115};
  assign _zz_117 = _zz_41[0];
  assign _zz_118 = {1'd0, _zz_117};
  assign _zz_119 = (left_bit_count_12 + _zz_121);
  assign _zz_120 = ((all_zeros_25 & _zz_122) & non_zeros_lzc_10);
  assign _zz_121 = {1'd0, _zz_120};
  assign _zz_122 = (whole_bit_count_13 + (~ all_zeros_25));
  assign _zz_123 = (left_bit_count_14 + _zz_125);
  assign _zz_124 = _zz_44[0];
  assign _zz_125 = {1'd0, _zz_124};
  assign _zz_126 = _zz_46[0];
  assign _zz_127 = {1'd0, _zz_126};
  assign _zz_128 = ((all_zeros_28 & _zz_130) & non_zeros_lzc_11);
  assign _zz_129 = {1'd0, _zz_128};
  assign _zz_130 = (whole_bit_count_14 + (~ all_zeros_28));
  assign _zz_131 = ((all_zeros_24 & _zz_133) & non_zeros_lzc_12);
  assign _zz_132 = {1'd0, _zz_131};
  assign _zz_133 = (whole_bit_count_12 + (~ all_zeros_24));
  assign _zz_134 = ((all_zeros_16 & _zz_136) & non_zeros_lzc_13);
  assign _zz_135 = {1'd0, _zz_134};
  assign _zz_136 = (whole_bit_count_8 + (~ all_zeros_16));
  assign _zz_137 = ((all_zeros & _zz_138) & non_zeros_lzc_14);
  assign _zz_138 = (whole_bit_count + (~ all_zeros));
  assign _zz_1 = a;
  assign all_zeros = ((! (_zz_1 != 16'h0)) ? 5'h1f : 5'h0);
  assign all_left_zeros = ((! (_zz_1[15 : 8] != 8'h0)) ? 5'h1f : 5'h0);
  assign whole_bit_count = 5'h10;
  assign left_bit_count = 5'h08;
  assign _zz_2 = _zz_1[7 : 0];
  assign all_zeros_1 = ((! (_zz_2 != 8'h0)) ? 4'b1111 : 4'b0000);
  assign all_left_zeros_1 = ((! (_zz_2[7 : 4] != 4'b0000)) ? 4'b1111 : 4'b0000);
  assign whole_bit_count_1 = 4'b1000;
  assign left_bit_count_1 = 4'b0100;
  assign _zz_3 = _zz_2[3 : 0];
  assign all_zeros_2 = ((! (_zz_3 != 4'b0000)) ? 3'b111 : 3'b000);
  assign all_left_zeros_2 = ((! (_zz_3[3 : 2] != 2'b00)) ? 3'b111 : 3'b000);
  assign whole_bit_count_2 = 3'b100;
  assign left_bit_count_2 = 3'b010;
  assign _zz_4 = _zz_3[1 : 0];
  assign all_zeros_3 = ((! (_zz_4 != 2'b00)) ? 2'b11 : 2'b00);
  assign all_left_zeros_3 = ((! (_zz_4[1 : 1] != 1'b0)) ? 2'b11 : 2'b00);
  assign whole_bit_count_3 = 2'b10;
  assign left_bit_count_3 = 2'b01;
  assign _zz_5 = _zz_4[0 : 0];
  assign _zz_6 = _zz_5;
  assign all_zeros_4 = ((! (_zz_6 != 1'b0)) ? 1'b1 : 1'b0);
  assign all_left_zeros_4 = ((! (_zz_6[0 : 0] != 1'b0)) ? 1'b1 : 1'b0);
  assign left_all_zeros_count = (all_left_zeros_3 & _zz_48);
  assign _zz_7 = _zz_4[1 : 1];
  assign _zz_8 = _zz_7;
  assign all_zeros_5 = ((! (_zz_8 != 1'b0)) ? 1'b1 : 1'b0);
  assign all_left_zeros_5 = ((! (_zz_8[0 : 0] != 1'b0)) ? 1'b1 : 1'b0);
  assign left_non_all_zeros_count = ((~ all_left_zeros_3) & _zz_52);
  assign non_zeros_lzc = (left_all_zeros_count + left_non_all_zeros_count);
  assign left_all_zeros_count_1 = (all_left_zeros_2 & _zz_53);
  assign _zz_9 = _zz_3[3 : 2];
  assign all_zeros_6 = ((! (_zz_9 != 2'b00)) ? 2'b11 : 2'b00);
  assign all_left_zeros_6 = ((! (_zz_9[1 : 1] != 1'b0)) ? 2'b11 : 2'b00);
  assign whole_bit_count_4 = 2'b10;
  assign left_bit_count_4 = 2'b01;
  assign _zz_10 = _zz_9[0 : 0];
  assign _zz_11 = _zz_10;
  assign all_zeros_7 = ((! (_zz_11 != 1'b0)) ? 1'b1 : 1'b0);
  assign all_left_zeros_7 = ((! (_zz_11[0 : 0] != 1'b0)) ? 1'b1 : 1'b0);
  assign left_all_zeros_count_2 = (all_left_zeros_6 & _zz_57);
  assign _zz_12 = _zz_9[1 : 1];
  assign _zz_13 = _zz_12;
  assign all_zeros_8 = ((! (_zz_13 != 1'b0)) ? 1'b1 : 1'b0);
  assign all_left_zeros_8 = ((! (_zz_13[0 : 0] != 1'b0)) ? 1'b1 : 1'b0);
  assign left_non_all_zeros_count_1 = ((~ all_left_zeros_6) & _zz_61);
  assign non_zeros_lzc_1 = (left_all_zeros_count_2 + left_non_all_zeros_count_1);
  assign left_non_all_zeros_count_2 = ((~ all_left_zeros_2) & _zz_63);
  assign non_zeros_lzc_2 = (left_all_zeros_count_1 + left_non_all_zeros_count_2);
  assign left_all_zeros_count_3 = (all_left_zeros_1 & _zz_65);
  assign _zz_14 = _zz_2[7 : 4];
  assign all_zeros_9 = ((! (_zz_14 != 4'b0000)) ? 3'b111 : 3'b000);
  assign all_left_zeros_9 = ((! (_zz_14[3 : 2] != 2'b00)) ? 3'b111 : 3'b000);
  assign whole_bit_count_5 = 3'b100;
  assign left_bit_count_5 = 3'b010;
  assign _zz_15 = _zz_14[1 : 0];
  assign all_zeros_10 = ((! (_zz_15 != 2'b00)) ? 2'b11 : 2'b00);
  assign all_left_zeros_10 = ((! (_zz_15[1 : 1] != 1'b0)) ? 2'b11 : 2'b00);
  assign whole_bit_count_6 = 2'b10;
  assign left_bit_count_6 = 2'b01;
  assign _zz_16 = _zz_15[0 : 0];
  assign _zz_17 = _zz_16;
  assign all_zeros_11 = ((! (_zz_17 != 1'b0)) ? 1'b1 : 1'b0);
  assign all_left_zeros_11 = ((! (_zz_17[0 : 0] != 1'b0)) ? 1'b1 : 1'b0);
  assign left_all_zeros_count_4 = (all_left_zeros_10 & _zz_69);
  assign _zz_18 = _zz_15[1 : 1];
  assign _zz_19 = _zz_18;
  assign all_zeros_12 = ((! (_zz_19 != 1'b0)) ? 1'b1 : 1'b0);
  assign all_left_zeros_12 = ((! (_zz_19[0 : 0] != 1'b0)) ? 1'b1 : 1'b0);
  assign left_non_all_zeros_count_3 = ((~ all_left_zeros_10) & _zz_73);
  assign non_zeros_lzc_3 = (left_all_zeros_count_4 + left_non_all_zeros_count_3);
  assign left_all_zeros_count_5 = (all_left_zeros_9 & _zz_74);
  assign _zz_20 = _zz_14[3 : 2];
  assign all_zeros_13 = ((! (_zz_20 != 2'b00)) ? 2'b11 : 2'b00);
  assign all_left_zeros_13 = ((! (_zz_20[1 : 1] != 1'b0)) ? 2'b11 : 2'b00);
  assign whole_bit_count_7 = 2'b10;
  assign left_bit_count_7 = 2'b01;
  assign _zz_21 = _zz_20[0 : 0];
  assign _zz_22 = _zz_21;
  assign all_zeros_14 = ((! (_zz_22 != 1'b0)) ? 1'b1 : 1'b0);
  assign all_left_zeros_14 = ((! (_zz_22[0 : 0] != 1'b0)) ? 1'b1 : 1'b0);
  assign left_all_zeros_count_6 = (all_left_zeros_13 & _zz_78);
  assign _zz_23 = _zz_20[1 : 1];
  assign _zz_24 = _zz_23;
  assign all_zeros_15 = ((! (_zz_24 != 1'b0)) ? 1'b1 : 1'b0);
  assign all_left_zeros_15 = ((! (_zz_24[0 : 0] != 1'b0)) ? 1'b1 : 1'b0);
  assign left_non_all_zeros_count_4 = ((~ all_left_zeros_13) & _zz_82);
  assign non_zeros_lzc_4 = (left_all_zeros_count_6 + left_non_all_zeros_count_4);
  assign left_non_all_zeros_count_5 = ((~ all_left_zeros_9) & _zz_84);
  assign non_zeros_lzc_5 = (left_all_zeros_count_5 + left_non_all_zeros_count_5);
  assign left_non_all_zeros_count_6 = ((~ all_left_zeros_1) & _zz_87);
  assign non_zeros_lzc_6 = (left_all_zeros_count_3 + left_non_all_zeros_count_6);
  assign left_all_zeros_count_7 = (all_left_zeros & _zz_89);
  assign _zz_25 = _zz_1[15 : 8];
  assign all_zeros_16 = ((! (_zz_25 != 8'h0)) ? 4'b1111 : 4'b0000);
  assign all_left_zeros_16 = ((! (_zz_25[7 : 4] != 4'b0000)) ? 4'b1111 : 4'b0000);
  assign whole_bit_count_8 = 4'b1000;
  assign left_bit_count_8 = 4'b0100;
  assign _zz_26 = _zz_25[3 : 0];
  assign all_zeros_17 = ((! (_zz_26 != 4'b0000)) ? 3'b111 : 3'b000);
  assign all_left_zeros_17 = ((! (_zz_26[3 : 2] != 2'b00)) ? 3'b111 : 3'b000);
  assign whole_bit_count_9 = 3'b100;
  assign left_bit_count_9 = 3'b010;
  assign _zz_27 = _zz_26[1 : 0];
  assign all_zeros_18 = ((! (_zz_27 != 2'b00)) ? 2'b11 : 2'b00);
  assign all_left_zeros_18 = ((! (_zz_27[1 : 1] != 1'b0)) ? 2'b11 : 2'b00);
  assign whole_bit_count_10 = 2'b10;
  assign left_bit_count_10 = 2'b01;
  assign _zz_28 = _zz_27[0 : 0];
  assign _zz_29 = _zz_28;
  assign all_zeros_19 = ((! (_zz_29 != 1'b0)) ? 1'b1 : 1'b0);
  assign all_left_zeros_19 = ((! (_zz_29[0 : 0] != 1'b0)) ? 1'b1 : 1'b0);
  assign left_all_zeros_count_8 = (all_left_zeros_18 & _zz_93);
  assign _zz_30 = _zz_27[1 : 1];
  assign _zz_31 = _zz_30;
  assign all_zeros_20 = ((! (_zz_31 != 1'b0)) ? 1'b1 : 1'b0);
  assign all_left_zeros_20 = ((! (_zz_31[0 : 0] != 1'b0)) ? 1'b1 : 1'b0);
  assign left_non_all_zeros_count_7 = ((~ all_left_zeros_18) & _zz_97);
  assign non_zeros_lzc_7 = (left_all_zeros_count_8 + left_non_all_zeros_count_7);
  assign left_all_zeros_count_9 = (all_left_zeros_17 & _zz_98);
  assign _zz_32 = _zz_26[3 : 2];
  assign all_zeros_21 = ((! (_zz_32 != 2'b00)) ? 2'b11 : 2'b00);
  assign all_left_zeros_21 = ((! (_zz_32[1 : 1] != 1'b0)) ? 2'b11 : 2'b00);
  assign whole_bit_count_11 = 2'b10;
  assign left_bit_count_11 = 2'b01;
  assign _zz_33 = _zz_32[0 : 0];
  assign _zz_34 = _zz_33;
  assign all_zeros_22 = ((! (_zz_34 != 1'b0)) ? 1'b1 : 1'b0);
  assign all_left_zeros_22 = ((! (_zz_34[0 : 0] != 1'b0)) ? 1'b1 : 1'b0);
  assign left_all_zeros_count_10 = (all_left_zeros_21 & _zz_102);
  assign _zz_35 = _zz_32[1 : 1];
  assign _zz_36 = _zz_35;
  assign all_zeros_23 = ((! (_zz_36 != 1'b0)) ? 1'b1 : 1'b0);
  assign all_left_zeros_23 = ((! (_zz_36[0 : 0] != 1'b0)) ? 1'b1 : 1'b0);
  assign left_non_all_zeros_count_8 = ((~ all_left_zeros_21) & _zz_106);
  assign non_zeros_lzc_8 = (left_all_zeros_count_10 + left_non_all_zeros_count_8);
  assign left_non_all_zeros_count_9 = ((~ all_left_zeros_17) & _zz_108);
  assign non_zeros_lzc_9 = (left_all_zeros_count_9 + left_non_all_zeros_count_9);
  assign left_all_zeros_count_11 = (all_left_zeros_16 & _zz_110);
  assign _zz_37 = _zz_25[7 : 4];
  assign all_zeros_24 = ((! (_zz_37 != 4'b0000)) ? 3'b111 : 3'b000);
  assign all_left_zeros_24 = ((! (_zz_37[3 : 2] != 2'b00)) ? 3'b111 : 3'b000);
  assign whole_bit_count_12 = 3'b100;
  assign left_bit_count_12 = 3'b010;
  assign _zz_38 = _zz_37[1 : 0];
  assign all_zeros_25 = ((! (_zz_38 != 2'b00)) ? 2'b11 : 2'b00);
  assign all_left_zeros_25 = ((! (_zz_38[1 : 1] != 1'b0)) ? 2'b11 : 2'b00);
  assign whole_bit_count_13 = 2'b10;
  assign left_bit_count_13 = 2'b01;
  assign _zz_39 = _zz_38[0 : 0];
  assign _zz_40 = _zz_39;
  assign all_zeros_26 = ((! (_zz_40 != 1'b0)) ? 1'b1 : 1'b0);
  assign all_left_zeros_26 = ((! (_zz_40[0 : 0] != 1'b0)) ? 1'b1 : 1'b0);
  assign left_all_zeros_count_12 = (all_left_zeros_25 & _zz_114);
  assign _zz_41 = _zz_38[1 : 1];
  assign _zz_42 = _zz_41;
  assign all_zeros_27 = ((! (_zz_42 != 1'b0)) ? 1'b1 : 1'b0);
  assign all_left_zeros_27 = ((! (_zz_42[0 : 0] != 1'b0)) ? 1'b1 : 1'b0);
  assign left_non_all_zeros_count_10 = ((~ all_left_zeros_25) & _zz_118);
  assign non_zeros_lzc_10 = (left_all_zeros_count_12 + left_non_all_zeros_count_10);
  assign left_all_zeros_count_13 = (all_left_zeros_24 & _zz_119);
  assign _zz_43 = _zz_37[3 : 2];
  assign all_zeros_28 = ((! (_zz_43 != 2'b00)) ? 2'b11 : 2'b00);
  assign all_left_zeros_28 = ((! (_zz_43[1 : 1] != 1'b0)) ? 2'b11 : 2'b00);
  assign whole_bit_count_14 = 2'b10;
  assign left_bit_count_14 = 2'b01;
  assign _zz_44 = _zz_43[0 : 0];
  assign _zz_45 = _zz_44;
  assign all_zeros_29 = ((! (_zz_45 != 1'b0)) ? 1'b1 : 1'b0);
  assign all_left_zeros_29 = ((! (_zz_45[0 : 0] != 1'b0)) ? 1'b1 : 1'b0);
  assign left_all_zeros_count_14 = (all_left_zeros_28 & _zz_123);
  assign _zz_46 = _zz_43[1 : 1];
  assign _zz_47 = _zz_46;
  assign all_zeros_30 = ((! (_zz_47 != 1'b0)) ? 1'b1 : 1'b0);
  assign all_left_zeros_30 = ((! (_zz_47[0 : 0] != 1'b0)) ? 1'b1 : 1'b0);
  assign left_non_all_zeros_count_11 = ((~ all_left_zeros_28) & _zz_127);
  assign non_zeros_lzc_11 = (left_all_zeros_count_14 + left_non_all_zeros_count_11);
  assign left_non_all_zeros_count_12 = ((~ all_left_zeros_24) & _zz_129);
  assign non_zeros_lzc_12 = (left_all_zeros_count_13 + left_non_all_zeros_count_12);
  assign left_non_all_zeros_count_13 = ((~ all_left_zeros_16) & _zz_132);
  assign non_zeros_lzc_13 = (left_all_zeros_count_11 + left_non_all_zeros_count_13);
  assign left_non_all_zeros_count_14 = ((~ all_left_zeros) & _zz_135);
  assign non_zeros_lzc_14 = (left_all_zeros_count_7 + left_non_all_zeros_count_14);
  assign a_lzc = {11'd0, _zz_137};

endmodule
