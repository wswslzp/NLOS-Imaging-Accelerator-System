// Generator : SpinalHDL v1.4.0    git head : ecb5a80b713566f417ea3ea061f9969e73770a7f
// Date      : 20/05/2020, 21:49:53
// Component : CoefLoadUnit



module CoefLoadUnit (
  input               axi4_aw_valid,
  output              axi4_aw_ready,
  input      [31:0]   axi4_aw_payload_addr,
  input      [3:0]    axi4_aw_payload_id,
  input      [7:0]    axi4_aw_payload_len,
  input      [2:0]    axi4_aw_payload_size,
  input      [1:0]    axi4_aw_payload_burst,
  input               axi4_w_valid,
  output              axi4_w_ready,
  input      [31:0]   axi4_w_payload_data,
  input      [3:0]    axi4_w_payload_strb,
  input               axi4_w_payload_last,
  output              axi4_b_valid,
  input               axi4_b_ready,
  output     [3:0]    axi4_b_payload_id,
  output     [1:0]    axi4_b_payload_resp,
  output              io_coef_out_valid,
  output     [15:0]   io_coef_out_payload_0_0_0_real,
  output     [15:0]   io_coef_out_payload_0_0_0_imag,
  output     [15:0]   io_coef_out_payload_0_0_1_real,
  output     [15:0]   io_coef_out_payload_0_0_1_imag,
  output     [15:0]   io_coef_out_payload_0_0_2_real,
  output     [15:0]   io_coef_out_payload_0_0_2_imag,
  output     [15:0]   io_coef_out_payload_0_0_3_real,
  output     [15:0]   io_coef_out_payload_0_0_3_imag,
  output     [15:0]   io_coef_out_payload_0_0_4_real,
  output     [15:0]   io_coef_out_payload_0_0_4_imag,
  output     [15:0]   io_coef_out_payload_0_0_5_real,
  output     [15:0]   io_coef_out_payload_0_0_5_imag,
  output     [15:0]   io_coef_out_payload_0_0_6_real,
  output     [15:0]   io_coef_out_payload_0_0_6_imag,
  output     [15:0]   io_coef_out_payload_0_0_7_real,
  output     [15:0]   io_coef_out_payload_0_0_7_imag,
  output     [15:0]   io_coef_out_payload_0_0_8_real,
  output     [15:0]   io_coef_out_payload_0_0_8_imag,
  output     [15:0]   io_coef_out_payload_0_0_9_real,
  output     [15:0]   io_coef_out_payload_0_0_9_imag,
  output     [15:0]   io_coef_out_payload_0_0_10_real,
  output     [15:0]   io_coef_out_payload_0_0_10_imag,
  output     [15:0]   io_coef_out_payload_0_0_11_real,
  output     [15:0]   io_coef_out_payload_0_0_11_imag,
  output     [15:0]   io_coef_out_payload_0_0_12_real,
  output     [15:0]   io_coef_out_payload_0_0_12_imag,
  output     [15:0]   io_coef_out_payload_0_0_13_real,
  output     [15:0]   io_coef_out_payload_0_0_13_imag,
  output     [15:0]   io_coef_out_payload_0_0_14_real,
  output     [15:0]   io_coef_out_payload_0_0_14_imag,
  output     [15:0]   io_coef_out_payload_0_0_15_real,
  output     [15:0]   io_coef_out_payload_0_0_15_imag,
  output     [15:0]   io_coef_out_payload_0_0_16_real,
  output     [15:0]   io_coef_out_payload_0_0_16_imag,
  output     [15:0]   io_coef_out_payload_0_0_17_real,
  output     [15:0]   io_coef_out_payload_0_0_17_imag,
  output     [15:0]   io_coef_out_payload_0_0_18_real,
  output     [15:0]   io_coef_out_payload_0_0_18_imag,
  output     [15:0]   io_coef_out_payload_0_0_19_real,
  output     [15:0]   io_coef_out_payload_0_0_19_imag,
  output     [15:0]   io_coef_out_payload_0_0_20_real,
  output     [15:0]   io_coef_out_payload_0_0_20_imag,
  output     [15:0]   io_coef_out_payload_0_0_21_real,
  output     [15:0]   io_coef_out_payload_0_0_21_imag,
  output     [15:0]   io_coef_out_payload_0_0_22_real,
  output     [15:0]   io_coef_out_payload_0_0_22_imag,
  output     [15:0]   io_coef_out_payload_0_0_23_real,
  output     [15:0]   io_coef_out_payload_0_0_23_imag,
  output     [15:0]   io_coef_out_payload_0_0_24_real,
  output     [15:0]   io_coef_out_payload_0_0_24_imag,
  output     [15:0]   io_coef_out_payload_0_0_25_real,
  output     [15:0]   io_coef_out_payload_0_0_25_imag,
  output     [15:0]   io_coef_out_payload_0_0_26_real,
  output     [15:0]   io_coef_out_payload_0_0_26_imag,
  output     [15:0]   io_coef_out_payload_0_0_27_real,
  output     [15:0]   io_coef_out_payload_0_0_27_imag,
  output     [15:0]   io_coef_out_payload_0_0_28_real,
  output     [15:0]   io_coef_out_payload_0_0_28_imag,
  output     [15:0]   io_coef_out_payload_0_0_29_real,
  output     [15:0]   io_coef_out_payload_0_0_29_imag,
  output     [15:0]   io_coef_out_payload_0_0_30_real,
  output     [15:0]   io_coef_out_payload_0_0_30_imag,
  output     [15:0]   io_coef_out_payload_0_0_31_real,
  output     [15:0]   io_coef_out_payload_0_0_31_imag,
  output     [15:0]   io_coef_out_payload_0_0_32_real,
  output     [15:0]   io_coef_out_payload_0_0_32_imag,
  output     [15:0]   io_coef_out_payload_0_0_33_real,
  output     [15:0]   io_coef_out_payload_0_0_33_imag,
  output     [15:0]   io_coef_out_payload_0_0_34_real,
  output     [15:0]   io_coef_out_payload_0_0_34_imag,
  output     [15:0]   io_coef_out_payload_0_0_35_real,
  output     [15:0]   io_coef_out_payload_0_0_35_imag,
  output     [15:0]   io_coef_out_payload_0_0_36_real,
  output     [15:0]   io_coef_out_payload_0_0_36_imag,
  output     [15:0]   io_coef_out_payload_0_0_37_real,
  output     [15:0]   io_coef_out_payload_0_0_37_imag,
  output     [15:0]   io_coef_out_payload_0_0_38_real,
  output     [15:0]   io_coef_out_payload_0_0_38_imag,
  output     [15:0]   io_coef_out_payload_0_0_39_real,
  output     [15:0]   io_coef_out_payload_0_0_39_imag,
  output     [15:0]   io_coef_out_payload_0_0_40_real,
  output     [15:0]   io_coef_out_payload_0_0_40_imag,
  output     [15:0]   io_coef_out_payload_0_0_41_real,
  output     [15:0]   io_coef_out_payload_0_0_41_imag,
  output     [15:0]   io_coef_out_payload_0_0_42_real,
  output     [15:0]   io_coef_out_payload_0_0_42_imag,
  output     [15:0]   io_coef_out_payload_0_0_43_real,
  output     [15:0]   io_coef_out_payload_0_0_43_imag,
  output     [15:0]   io_coef_out_payload_0_0_44_real,
  output     [15:0]   io_coef_out_payload_0_0_44_imag,
  output     [15:0]   io_coef_out_payload_0_0_45_real,
  output     [15:0]   io_coef_out_payload_0_0_45_imag,
  output     [15:0]   io_coef_out_payload_0_0_46_real,
  output     [15:0]   io_coef_out_payload_0_0_46_imag,
  output     [15:0]   io_coef_out_payload_0_0_47_real,
  output     [15:0]   io_coef_out_payload_0_0_47_imag,
  output     [15:0]   io_coef_out_payload_0_0_48_real,
  output     [15:0]   io_coef_out_payload_0_0_48_imag,
  output     [15:0]   io_coef_out_payload_0_0_49_real,
  output     [15:0]   io_coef_out_payload_0_0_49_imag,
  output     [15:0]   io_coef_out_payload_0_1_0_real,
  output     [15:0]   io_coef_out_payload_0_1_0_imag,
  output     [15:0]   io_coef_out_payload_0_1_1_real,
  output     [15:0]   io_coef_out_payload_0_1_1_imag,
  output     [15:0]   io_coef_out_payload_0_1_2_real,
  output     [15:0]   io_coef_out_payload_0_1_2_imag,
  output     [15:0]   io_coef_out_payload_0_1_3_real,
  output     [15:0]   io_coef_out_payload_0_1_3_imag,
  output     [15:0]   io_coef_out_payload_0_1_4_real,
  output     [15:0]   io_coef_out_payload_0_1_4_imag,
  output     [15:0]   io_coef_out_payload_0_1_5_real,
  output     [15:0]   io_coef_out_payload_0_1_5_imag,
  output     [15:0]   io_coef_out_payload_0_1_6_real,
  output     [15:0]   io_coef_out_payload_0_1_6_imag,
  output     [15:0]   io_coef_out_payload_0_1_7_real,
  output     [15:0]   io_coef_out_payload_0_1_7_imag,
  output     [15:0]   io_coef_out_payload_0_1_8_real,
  output     [15:0]   io_coef_out_payload_0_1_8_imag,
  output     [15:0]   io_coef_out_payload_0_1_9_real,
  output     [15:0]   io_coef_out_payload_0_1_9_imag,
  output     [15:0]   io_coef_out_payload_0_1_10_real,
  output     [15:0]   io_coef_out_payload_0_1_10_imag,
  output     [15:0]   io_coef_out_payload_0_1_11_real,
  output     [15:0]   io_coef_out_payload_0_1_11_imag,
  output     [15:0]   io_coef_out_payload_0_1_12_real,
  output     [15:0]   io_coef_out_payload_0_1_12_imag,
  output     [15:0]   io_coef_out_payload_0_1_13_real,
  output     [15:0]   io_coef_out_payload_0_1_13_imag,
  output     [15:0]   io_coef_out_payload_0_1_14_real,
  output     [15:0]   io_coef_out_payload_0_1_14_imag,
  output     [15:0]   io_coef_out_payload_0_1_15_real,
  output     [15:0]   io_coef_out_payload_0_1_15_imag,
  output     [15:0]   io_coef_out_payload_0_1_16_real,
  output     [15:0]   io_coef_out_payload_0_1_16_imag,
  output     [15:0]   io_coef_out_payload_0_1_17_real,
  output     [15:0]   io_coef_out_payload_0_1_17_imag,
  output     [15:0]   io_coef_out_payload_0_1_18_real,
  output     [15:0]   io_coef_out_payload_0_1_18_imag,
  output     [15:0]   io_coef_out_payload_0_1_19_real,
  output     [15:0]   io_coef_out_payload_0_1_19_imag,
  output     [15:0]   io_coef_out_payload_0_1_20_real,
  output     [15:0]   io_coef_out_payload_0_1_20_imag,
  output     [15:0]   io_coef_out_payload_0_1_21_real,
  output     [15:0]   io_coef_out_payload_0_1_21_imag,
  output     [15:0]   io_coef_out_payload_0_1_22_real,
  output     [15:0]   io_coef_out_payload_0_1_22_imag,
  output     [15:0]   io_coef_out_payload_0_1_23_real,
  output     [15:0]   io_coef_out_payload_0_1_23_imag,
  output     [15:0]   io_coef_out_payload_0_1_24_real,
  output     [15:0]   io_coef_out_payload_0_1_24_imag,
  output     [15:0]   io_coef_out_payload_0_1_25_real,
  output     [15:0]   io_coef_out_payload_0_1_25_imag,
  output     [15:0]   io_coef_out_payload_0_1_26_real,
  output     [15:0]   io_coef_out_payload_0_1_26_imag,
  output     [15:0]   io_coef_out_payload_0_1_27_real,
  output     [15:0]   io_coef_out_payload_0_1_27_imag,
  output     [15:0]   io_coef_out_payload_0_1_28_real,
  output     [15:0]   io_coef_out_payload_0_1_28_imag,
  output     [15:0]   io_coef_out_payload_0_1_29_real,
  output     [15:0]   io_coef_out_payload_0_1_29_imag,
  output     [15:0]   io_coef_out_payload_0_1_30_real,
  output     [15:0]   io_coef_out_payload_0_1_30_imag,
  output     [15:0]   io_coef_out_payload_0_1_31_real,
  output     [15:0]   io_coef_out_payload_0_1_31_imag,
  output     [15:0]   io_coef_out_payload_0_1_32_real,
  output     [15:0]   io_coef_out_payload_0_1_32_imag,
  output     [15:0]   io_coef_out_payload_0_1_33_real,
  output     [15:0]   io_coef_out_payload_0_1_33_imag,
  output     [15:0]   io_coef_out_payload_0_1_34_real,
  output     [15:0]   io_coef_out_payload_0_1_34_imag,
  output     [15:0]   io_coef_out_payload_0_1_35_real,
  output     [15:0]   io_coef_out_payload_0_1_35_imag,
  output     [15:0]   io_coef_out_payload_0_1_36_real,
  output     [15:0]   io_coef_out_payload_0_1_36_imag,
  output     [15:0]   io_coef_out_payload_0_1_37_real,
  output     [15:0]   io_coef_out_payload_0_1_37_imag,
  output     [15:0]   io_coef_out_payload_0_1_38_real,
  output     [15:0]   io_coef_out_payload_0_1_38_imag,
  output     [15:0]   io_coef_out_payload_0_1_39_real,
  output     [15:0]   io_coef_out_payload_0_1_39_imag,
  output     [15:0]   io_coef_out_payload_0_1_40_real,
  output     [15:0]   io_coef_out_payload_0_1_40_imag,
  output     [15:0]   io_coef_out_payload_0_1_41_real,
  output     [15:0]   io_coef_out_payload_0_1_41_imag,
  output     [15:0]   io_coef_out_payload_0_1_42_real,
  output     [15:0]   io_coef_out_payload_0_1_42_imag,
  output     [15:0]   io_coef_out_payload_0_1_43_real,
  output     [15:0]   io_coef_out_payload_0_1_43_imag,
  output     [15:0]   io_coef_out_payload_0_1_44_real,
  output     [15:0]   io_coef_out_payload_0_1_44_imag,
  output     [15:0]   io_coef_out_payload_0_1_45_real,
  output     [15:0]   io_coef_out_payload_0_1_45_imag,
  output     [15:0]   io_coef_out_payload_0_1_46_real,
  output     [15:0]   io_coef_out_payload_0_1_46_imag,
  output     [15:0]   io_coef_out_payload_0_1_47_real,
  output     [15:0]   io_coef_out_payload_0_1_47_imag,
  output     [15:0]   io_coef_out_payload_0_1_48_real,
  output     [15:0]   io_coef_out_payload_0_1_48_imag,
  output     [15:0]   io_coef_out_payload_0_1_49_real,
  output     [15:0]   io_coef_out_payload_0_1_49_imag,
  output     [15:0]   io_coef_out_payload_0_2_0_real,
  output     [15:0]   io_coef_out_payload_0_2_0_imag,
  output     [15:0]   io_coef_out_payload_0_2_1_real,
  output     [15:0]   io_coef_out_payload_0_2_1_imag,
  output     [15:0]   io_coef_out_payload_0_2_2_real,
  output     [15:0]   io_coef_out_payload_0_2_2_imag,
  output     [15:0]   io_coef_out_payload_0_2_3_real,
  output     [15:0]   io_coef_out_payload_0_2_3_imag,
  output     [15:0]   io_coef_out_payload_0_2_4_real,
  output     [15:0]   io_coef_out_payload_0_2_4_imag,
  output     [15:0]   io_coef_out_payload_0_2_5_real,
  output     [15:0]   io_coef_out_payload_0_2_5_imag,
  output     [15:0]   io_coef_out_payload_0_2_6_real,
  output     [15:0]   io_coef_out_payload_0_2_6_imag,
  output     [15:0]   io_coef_out_payload_0_2_7_real,
  output     [15:0]   io_coef_out_payload_0_2_7_imag,
  output     [15:0]   io_coef_out_payload_0_2_8_real,
  output     [15:0]   io_coef_out_payload_0_2_8_imag,
  output     [15:0]   io_coef_out_payload_0_2_9_real,
  output     [15:0]   io_coef_out_payload_0_2_9_imag,
  output     [15:0]   io_coef_out_payload_0_2_10_real,
  output     [15:0]   io_coef_out_payload_0_2_10_imag,
  output     [15:0]   io_coef_out_payload_0_2_11_real,
  output     [15:0]   io_coef_out_payload_0_2_11_imag,
  output     [15:0]   io_coef_out_payload_0_2_12_real,
  output     [15:0]   io_coef_out_payload_0_2_12_imag,
  output     [15:0]   io_coef_out_payload_0_2_13_real,
  output     [15:0]   io_coef_out_payload_0_2_13_imag,
  output     [15:0]   io_coef_out_payload_0_2_14_real,
  output     [15:0]   io_coef_out_payload_0_2_14_imag,
  output     [15:0]   io_coef_out_payload_0_2_15_real,
  output     [15:0]   io_coef_out_payload_0_2_15_imag,
  output     [15:0]   io_coef_out_payload_0_2_16_real,
  output     [15:0]   io_coef_out_payload_0_2_16_imag,
  output     [15:0]   io_coef_out_payload_0_2_17_real,
  output     [15:0]   io_coef_out_payload_0_2_17_imag,
  output     [15:0]   io_coef_out_payload_0_2_18_real,
  output     [15:0]   io_coef_out_payload_0_2_18_imag,
  output     [15:0]   io_coef_out_payload_0_2_19_real,
  output     [15:0]   io_coef_out_payload_0_2_19_imag,
  output     [15:0]   io_coef_out_payload_0_2_20_real,
  output     [15:0]   io_coef_out_payload_0_2_20_imag,
  output     [15:0]   io_coef_out_payload_0_2_21_real,
  output     [15:0]   io_coef_out_payload_0_2_21_imag,
  output     [15:0]   io_coef_out_payload_0_2_22_real,
  output     [15:0]   io_coef_out_payload_0_2_22_imag,
  output     [15:0]   io_coef_out_payload_0_2_23_real,
  output     [15:0]   io_coef_out_payload_0_2_23_imag,
  output     [15:0]   io_coef_out_payload_0_2_24_real,
  output     [15:0]   io_coef_out_payload_0_2_24_imag,
  output     [15:0]   io_coef_out_payload_0_2_25_real,
  output     [15:0]   io_coef_out_payload_0_2_25_imag,
  output     [15:0]   io_coef_out_payload_0_2_26_real,
  output     [15:0]   io_coef_out_payload_0_2_26_imag,
  output     [15:0]   io_coef_out_payload_0_2_27_real,
  output     [15:0]   io_coef_out_payload_0_2_27_imag,
  output     [15:0]   io_coef_out_payload_0_2_28_real,
  output     [15:0]   io_coef_out_payload_0_2_28_imag,
  output     [15:0]   io_coef_out_payload_0_2_29_real,
  output     [15:0]   io_coef_out_payload_0_2_29_imag,
  output     [15:0]   io_coef_out_payload_0_2_30_real,
  output     [15:0]   io_coef_out_payload_0_2_30_imag,
  output     [15:0]   io_coef_out_payload_0_2_31_real,
  output     [15:0]   io_coef_out_payload_0_2_31_imag,
  output     [15:0]   io_coef_out_payload_0_2_32_real,
  output     [15:0]   io_coef_out_payload_0_2_32_imag,
  output     [15:0]   io_coef_out_payload_0_2_33_real,
  output     [15:0]   io_coef_out_payload_0_2_33_imag,
  output     [15:0]   io_coef_out_payload_0_2_34_real,
  output     [15:0]   io_coef_out_payload_0_2_34_imag,
  output     [15:0]   io_coef_out_payload_0_2_35_real,
  output     [15:0]   io_coef_out_payload_0_2_35_imag,
  output     [15:0]   io_coef_out_payload_0_2_36_real,
  output     [15:0]   io_coef_out_payload_0_2_36_imag,
  output     [15:0]   io_coef_out_payload_0_2_37_real,
  output     [15:0]   io_coef_out_payload_0_2_37_imag,
  output     [15:0]   io_coef_out_payload_0_2_38_real,
  output     [15:0]   io_coef_out_payload_0_2_38_imag,
  output     [15:0]   io_coef_out_payload_0_2_39_real,
  output     [15:0]   io_coef_out_payload_0_2_39_imag,
  output     [15:0]   io_coef_out_payload_0_2_40_real,
  output     [15:0]   io_coef_out_payload_0_2_40_imag,
  output     [15:0]   io_coef_out_payload_0_2_41_real,
  output     [15:0]   io_coef_out_payload_0_2_41_imag,
  output     [15:0]   io_coef_out_payload_0_2_42_real,
  output     [15:0]   io_coef_out_payload_0_2_42_imag,
  output     [15:0]   io_coef_out_payload_0_2_43_real,
  output     [15:0]   io_coef_out_payload_0_2_43_imag,
  output     [15:0]   io_coef_out_payload_0_2_44_real,
  output     [15:0]   io_coef_out_payload_0_2_44_imag,
  output     [15:0]   io_coef_out_payload_0_2_45_real,
  output     [15:0]   io_coef_out_payload_0_2_45_imag,
  output     [15:0]   io_coef_out_payload_0_2_46_real,
  output     [15:0]   io_coef_out_payload_0_2_46_imag,
  output     [15:0]   io_coef_out_payload_0_2_47_real,
  output     [15:0]   io_coef_out_payload_0_2_47_imag,
  output     [15:0]   io_coef_out_payload_0_2_48_real,
  output     [15:0]   io_coef_out_payload_0_2_48_imag,
  output     [15:0]   io_coef_out_payload_0_2_49_real,
  output     [15:0]   io_coef_out_payload_0_2_49_imag,
  output     [15:0]   io_coef_out_payload_0_3_0_real,
  output     [15:0]   io_coef_out_payload_0_3_0_imag,
  output     [15:0]   io_coef_out_payload_0_3_1_real,
  output     [15:0]   io_coef_out_payload_0_3_1_imag,
  output     [15:0]   io_coef_out_payload_0_3_2_real,
  output     [15:0]   io_coef_out_payload_0_3_2_imag,
  output     [15:0]   io_coef_out_payload_0_3_3_real,
  output     [15:0]   io_coef_out_payload_0_3_3_imag,
  output     [15:0]   io_coef_out_payload_0_3_4_real,
  output     [15:0]   io_coef_out_payload_0_3_4_imag,
  output     [15:0]   io_coef_out_payload_0_3_5_real,
  output     [15:0]   io_coef_out_payload_0_3_5_imag,
  output     [15:0]   io_coef_out_payload_0_3_6_real,
  output     [15:0]   io_coef_out_payload_0_3_6_imag,
  output     [15:0]   io_coef_out_payload_0_3_7_real,
  output     [15:0]   io_coef_out_payload_0_3_7_imag,
  output     [15:0]   io_coef_out_payload_0_3_8_real,
  output     [15:0]   io_coef_out_payload_0_3_8_imag,
  output     [15:0]   io_coef_out_payload_0_3_9_real,
  output     [15:0]   io_coef_out_payload_0_3_9_imag,
  output     [15:0]   io_coef_out_payload_0_3_10_real,
  output     [15:0]   io_coef_out_payload_0_3_10_imag,
  output     [15:0]   io_coef_out_payload_0_3_11_real,
  output     [15:0]   io_coef_out_payload_0_3_11_imag,
  output     [15:0]   io_coef_out_payload_0_3_12_real,
  output     [15:0]   io_coef_out_payload_0_3_12_imag,
  output     [15:0]   io_coef_out_payload_0_3_13_real,
  output     [15:0]   io_coef_out_payload_0_3_13_imag,
  output     [15:0]   io_coef_out_payload_0_3_14_real,
  output     [15:0]   io_coef_out_payload_0_3_14_imag,
  output     [15:0]   io_coef_out_payload_0_3_15_real,
  output     [15:0]   io_coef_out_payload_0_3_15_imag,
  output     [15:0]   io_coef_out_payload_0_3_16_real,
  output     [15:0]   io_coef_out_payload_0_3_16_imag,
  output     [15:0]   io_coef_out_payload_0_3_17_real,
  output     [15:0]   io_coef_out_payload_0_3_17_imag,
  output     [15:0]   io_coef_out_payload_0_3_18_real,
  output     [15:0]   io_coef_out_payload_0_3_18_imag,
  output     [15:0]   io_coef_out_payload_0_3_19_real,
  output     [15:0]   io_coef_out_payload_0_3_19_imag,
  output     [15:0]   io_coef_out_payload_0_3_20_real,
  output     [15:0]   io_coef_out_payload_0_3_20_imag,
  output     [15:0]   io_coef_out_payload_0_3_21_real,
  output     [15:0]   io_coef_out_payload_0_3_21_imag,
  output     [15:0]   io_coef_out_payload_0_3_22_real,
  output     [15:0]   io_coef_out_payload_0_3_22_imag,
  output     [15:0]   io_coef_out_payload_0_3_23_real,
  output     [15:0]   io_coef_out_payload_0_3_23_imag,
  output     [15:0]   io_coef_out_payload_0_3_24_real,
  output     [15:0]   io_coef_out_payload_0_3_24_imag,
  output     [15:0]   io_coef_out_payload_0_3_25_real,
  output     [15:0]   io_coef_out_payload_0_3_25_imag,
  output     [15:0]   io_coef_out_payload_0_3_26_real,
  output     [15:0]   io_coef_out_payload_0_3_26_imag,
  output     [15:0]   io_coef_out_payload_0_3_27_real,
  output     [15:0]   io_coef_out_payload_0_3_27_imag,
  output     [15:0]   io_coef_out_payload_0_3_28_real,
  output     [15:0]   io_coef_out_payload_0_3_28_imag,
  output     [15:0]   io_coef_out_payload_0_3_29_real,
  output     [15:0]   io_coef_out_payload_0_3_29_imag,
  output     [15:0]   io_coef_out_payload_0_3_30_real,
  output     [15:0]   io_coef_out_payload_0_3_30_imag,
  output     [15:0]   io_coef_out_payload_0_3_31_real,
  output     [15:0]   io_coef_out_payload_0_3_31_imag,
  output     [15:0]   io_coef_out_payload_0_3_32_real,
  output     [15:0]   io_coef_out_payload_0_3_32_imag,
  output     [15:0]   io_coef_out_payload_0_3_33_real,
  output     [15:0]   io_coef_out_payload_0_3_33_imag,
  output     [15:0]   io_coef_out_payload_0_3_34_real,
  output     [15:0]   io_coef_out_payload_0_3_34_imag,
  output     [15:0]   io_coef_out_payload_0_3_35_real,
  output     [15:0]   io_coef_out_payload_0_3_35_imag,
  output     [15:0]   io_coef_out_payload_0_3_36_real,
  output     [15:0]   io_coef_out_payload_0_3_36_imag,
  output     [15:0]   io_coef_out_payload_0_3_37_real,
  output     [15:0]   io_coef_out_payload_0_3_37_imag,
  output     [15:0]   io_coef_out_payload_0_3_38_real,
  output     [15:0]   io_coef_out_payload_0_3_38_imag,
  output     [15:0]   io_coef_out_payload_0_3_39_real,
  output     [15:0]   io_coef_out_payload_0_3_39_imag,
  output     [15:0]   io_coef_out_payload_0_3_40_real,
  output     [15:0]   io_coef_out_payload_0_3_40_imag,
  output     [15:0]   io_coef_out_payload_0_3_41_real,
  output     [15:0]   io_coef_out_payload_0_3_41_imag,
  output     [15:0]   io_coef_out_payload_0_3_42_real,
  output     [15:0]   io_coef_out_payload_0_3_42_imag,
  output     [15:0]   io_coef_out_payload_0_3_43_real,
  output     [15:0]   io_coef_out_payload_0_3_43_imag,
  output     [15:0]   io_coef_out_payload_0_3_44_real,
  output     [15:0]   io_coef_out_payload_0_3_44_imag,
  output     [15:0]   io_coef_out_payload_0_3_45_real,
  output     [15:0]   io_coef_out_payload_0_3_45_imag,
  output     [15:0]   io_coef_out_payload_0_3_46_real,
  output     [15:0]   io_coef_out_payload_0_3_46_imag,
  output     [15:0]   io_coef_out_payload_0_3_47_real,
  output     [15:0]   io_coef_out_payload_0_3_47_imag,
  output     [15:0]   io_coef_out_payload_0_3_48_real,
  output     [15:0]   io_coef_out_payload_0_3_48_imag,
  output     [15:0]   io_coef_out_payload_0_3_49_real,
  output     [15:0]   io_coef_out_payload_0_3_49_imag,
  output     [15:0]   io_coef_out_payload_0_4_0_real,
  output     [15:0]   io_coef_out_payload_0_4_0_imag,
  output     [15:0]   io_coef_out_payload_0_4_1_real,
  output     [15:0]   io_coef_out_payload_0_4_1_imag,
  output     [15:0]   io_coef_out_payload_0_4_2_real,
  output     [15:0]   io_coef_out_payload_0_4_2_imag,
  output     [15:0]   io_coef_out_payload_0_4_3_real,
  output     [15:0]   io_coef_out_payload_0_4_3_imag,
  output     [15:0]   io_coef_out_payload_0_4_4_real,
  output     [15:0]   io_coef_out_payload_0_4_4_imag,
  output     [15:0]   io_coef_out_payload_0_4_5_real,
  output     [15:0]   io_coef_out_payload_0_4_5_imag,
  output     [15:0]   io_coef_out_payload_0_4_6_real,
  output     [15:0]   io_coef_out_payload_0_4_6_imag,
  output     [15:0]   io_coef_out_payload_0_4_7_real,
  output     [15:0]   io_coef_out_payload_0_4_7_imag,
  output     [15:0]   io_coef_out_payload_0_4_8_real,
  output     [15:0]   io_coef_out_payload_0_4_8_imag,
  output     [15:0]   io_coef_out_payload_0_4_9_real,
  output     [15:0]   io_coef_out_payload_0_4_9_imag,
  output     [15:0]   io_coef_out_payload_0_4_10_real,
  output     [15:0]   io_coef_out_payload_0_4_10_imag,
  output     [15:0]   io_coef_out_payload_0_4_11_real,
  output     [15:0]   io_coef_out_payload_0_4_11_imag,
  output     [15:0]   io_coef_out_payload_0_4_12_real,
  output     [15:0]   io_coef_out_payload_0_4_12_imag,
  output     [15:0]   io_coef_out_payload_0_4_13_real,
  output     [15:0]   io_coef_out_payload_0_4_13_imag,
  output     [15:0]   io_coef_out_payload_0_4_14_real,
  output     [15:0]   io_coef_out_payload_0_4_14_imag,
  output     [15:0]   io_coef_out_payload_0_4_15_real,
  output     [15:0]   io_coef_out_payload_0_4_15_imag,
  output     [15:0]   io_coef_out_payload_0_4_16_real,
  output     [15:0]   io_coef_out_payload_0_4_16_imag,
  output     [15:0]   io_coef_out_payload_0_4_17_real,
  output     [15:0]   io_coef_out_payload_0_4_17_imag,
  output     [15:0]   io_coef_out_payload_0_4_18_real,
  output     [15:0]   io_coef_out_payload_0_4_18_imag,
  output     [15:0]   io_coef_out_payload_0_4_19_real,
  output     [15:0]   io_coef_out_payload_0_4_19_imag,
  output     [15:0]   io_coef_out_payload_0_4_20_real,
  output     [15:0]   io_coef_out_payload_0_4_20_imag,
  output     [15:0]   io_coef_out_payload_0_4_21_real,
  output     [15:0]   io_coef_out_payload_0_4_21_imag,
  output     [15:0]   io_coef_out_payload_0_4_22_real,
  output     [15:0]   io_coef_out_payload_0_4_22_imag,
  output     [15:0]   io_coef_out_payload_0_4_23_real,
  output     [15:0]   io_coef_out_payload_0_4_23_imag,
  output     [15:0]   io_coef_out_payload_0_4_24_real,
  output     [15:0]   io_coef_out_payload_0_4_24_imag,
  output     [15:0]   io_coef_out_payload_0_4_25_real,
  output     [15:0]   io_coef_out_payload_0_4_25_imag,
  output     [15:0]   io_coef_out_payload_0_4_26_real,
  output     [15:0]   io_coef_out_payload_0_4_26_imag,
  output     [15:0]   io_coef_out_payload_0_4_27_real,
  output     [15:0]   io_coef_out_payload_0_4_27_imag,
  output     [15:0]   io_coef_out_payload_0_4_28_real,
  output     [15:0]   io_coef_out_payload_0_4_28_imag,
  output     [15:0]   io_coef_out_payload_0_4_29_real,
  output     [15:0]   io_coef_out_payload_0_4_29_imag,
  output     [15:0]   io_coef_out_payload_0_4_30_real,
  output     [15:0]   io_coef_out_payload_0_4_30_imag,
  output     [15:0]   io_coef_out_payload_0_4_31_real,
  output     [15:0]   io_coef_out_payload_0_4_31_imag,
  output     [15:0]   io_coef_out_payload_0_4_32_real,
  output     [15:0]   io_coef_out_payload_0_4_32_imag,
  output     [15:0]   io_coef_out_payload_0_4_33_real,
  output     [15:0]   io_coef_out_payload_0_4_33_imag,
  output     [15:0]   io_coef_out_payload_0_4_34_real,
  output     [15:0]   io_coef_out_payload_0_4_34_imag,
  output     [15:0]   io_coef_out_payload_0_4_35_real,
  output     [15:0]   io_coef_out_payload_0_4_35_imag,
  output     [15:0]   io_coef_out_payload_0_4_36_real,
  output     [15:0]   io_coef_out_payload_0_4_36_imag,
  output     [15:0]   io_coef_out_payload_0_4_37_real,
  output     [15:0]   io_coef_out_payload_0_4_37_imag,
  output     [15:0]   io_coef_out_payload_0_4_38_real,
  output     [15:0]   io_coef_out_payload_0_4_38_imag,
  output     [15:0]   io_coef_out_payload_0_4_39_real,
  output     [15:0]   io_coef_out_payload_0_4_39_imag,
  output     [15:0]   io_coef_out_payload_0_4_40_real,
  output     [15:0]   io_coef_out_payload_0_4_40_imag,
  output     [15:0]   io_coef_out_payload_0_4_41_real,
  output     [15:0]   io_coef_out_payload_0_4_41_imag,
  output     [15:0]   io_coef_out_payload_0_4_42_real,
  output     [15:0]   io_coef_out_payload_0_4_42_imag,
  output     [15:0]   io_coef_out_payload_0_4_43_real,
  output     [15:0]   io_coef_out_payload_0_4_43_imag,
  output     [15:0]   io_coef_out_payload_0_4_44_real,
  output     [15:0]   io_coef_out_payload_0_4_44_imag,
  output     [15:0]   io_coef_out_payload_0_4_45_real,
  output     [15:0]   io_coef_out_payload_0_4_45_imag,
  output     [15:0]   io_coef_out_payload_0_4_46_real,
  output     [15:0]   io_coef_out_payload_0_4_46_imag,
  output     [15:0]   io_coef_out_payload_0_4_47_real,
  output     [15:0]   io_coef_out_payload_0_4_47_imag,
  output     [15:0]   io_coef_out_payload_0_4_48_real,
  output     [15:0]   io_coef_out_payload_0_4_48_imag,
  output     [15:0]   io_coef_out_payload_0_4_49_real,
  output     [15:0]   io_coef_out_payload_0_4_49_imag,
  output     [15:0]   io_coef_out_payload_0_5_0_real,
  output     [15:0]   io_coef_out_payload_0_5_0_imag,
  output     [15:0]   io_coef_out_payload_0_5_1_real,
  output     [15:0]   io_coef_out_payload_0_5_1_imag,
  output     [15:0]   io_coef_out_payload_0_5_2_real,
  output     [15:0]   io_coef_out_payload_0_5_2_imag,
  output     [15:0]   io_coef_out_payload_0_5_3_real,
  output     [15:0]   io_coef_out_payload_0_5_3_imag,
  output     [15:0]   io_coef_out_payload_0_5_4_real,
  output     [15:0]   io_coef_out_payload_0_5_4_imag,
  output     [15:0]   io_coef_out_payload_0_5_5_real,
  output     [15:0]   io_coef_out_payload_0_5_5_imag,
  output     [15:0]   io_coef_out_payload_0_5_6_real,
  output     [15:0]   io_coef_out_payload_0_5_6_imag,
  output     [15:0]   io_coef_out_payload_0_5_7_real,
  output     [15:0]   io_coef_out_payload_0_5_7_imag,
  output     [15:0]   io_coef_out_payload_0_5_8_real,
  output     [15:0]   io_coef_out_payload_0_5_8_imag,
  output     [15:0]   io_coef_out_payload_0_5_9_real,
  output     [15:0]   io_coef_out_payload_0_5_9_imag,
  output     [15:0]   io_coef_out_payload_0_5_10_real,
  output     [15:0]   io_coef_out_payload_0_5_10_imag,
  output     [15:0]   io_coef_out_payload_0_5_11_real,
  output     [15:0]   io_coef_out_payload_0_5_11_imag,
  output     [15:0]   io_coef_out_payload_0_5_12_real,
  output     [15:0]   io_coef_out_payload_0_5_12_imag,
  output     [15:0]   io_coef_out_payload_0_5_13_real,
  output     [15:0]   io_coef_out_payload_0_5_13_imag,
  output     [15:0]   io_coef_out_payload_0_5_14_real,
  output     [15:0]   io_coef_out_payload_0_5_14_imag,
  output     [15:0]   io_coef_out_payload_0_5_15_real,
  output     [15:0]   io_coef_out_payload_0_5_15_imag,
  output     [15:0]   io_coef_out_payload_0_5_16_real,
  output     [15:0]   io_coef_out_payload_0_5_16_imag,
  output     [15:0]   io_coef_out_payload_0_5_17_real,
  output     [15:0]   io_coef_out_payload_0_5_17_imag,
  output     [15:0]   io_coef_out_payload_0_5_18_real,
  output     [15:0]   io_coef_out_payload_0_5_18_imag,
  output     [15:0]   io_coef_out_payload_0_5_19_real,
  output     [15:0]   io_coef_out_payload_0_5_19_imag,
  output     [15:0]   io_coef_out_payload_0_5_20_real,
  output     [15:0]   io_coef_out_payload_0_5_20_imag,
  output     [15:0]   io_coef_out_payload_0_5_21_real,
  output     [15:0]   io_coef_out_payload_0_5_21_imag,
  output     [15:0]   io_coef_out_payload_0_5_22_real,
  output     [15:0]   io_coef_out_payload_0_5_22_imag,
  output     [15:0]   io_coef_out_payload_0_5_23_real,
  output     [15:0]   io_coef_out_payload_0_5_23_imag,
  output     [15:0]   io_coef_out_payload_0_5_24_real,
  output     [15:0]   io_coef_out_payload_0_5_24_imag,
  output     [15:0]   io_coef_out_payload_0_5_25_real,
  output     [15:0]   io_coef_out_payload_0_5_25_imag,
  output     [15:0]   io_coef_out_payload_0_5_26_real,
  output     [15:0]   io_coef_out_payload_0_5_26_imag,
  output     [15:0]   io_coef_out_payload_0_5_27_real,
  output     [15:0]   io_coef_out_payload_0_5_27_imag,
  output     [15:0]   io_coef_out_payload_0_5_28_real,
  output     [15:0]   io_coef_out_payload_0_5_28_imag,
  output     [15:0]   io_coef_out_payload_0_5_29_real,
  output     [15:0]   io_coef_out_payload_0_5_29_imag,
  output     [15:0]   io_coef_out_payload_0_5_30_real,
  output     [15:0]   io_coef_out_payload_0_5_30_imag,
  output     [15:0]   io_coef_out_payload_0_5_31_real,
  output     [15:0]   io_coef_out_payload_0_5_31_imag,
  output     [15:0]   io_coef_out_payload_0_5_32_real,
  output     [15:0]   io_coef_out_payload_0_5_32_imag,
  output     [15:0]   io_coef_out_payload_0_5_33_real,
  output     [15:0]   io_coef_out_payload_0_5_33_imag,
  output     [15:0]   io_coef_out_payload_0_5_34_real,
  output     [15:0]   io_coef_out_payload_0_5_34_imag,
  output     [15:0]   io_coef_out_payload_0_5_35_real,
  output     [15:0]   io_coef_out_payload_0_5_35_imag,
  output     [15:0]   io_coef_out_payload_0_5_36_real,
  output     [15:0]   io_coef_out_payload_0_5_36_imag,
  output     [15:0]   io_coef_out_payload_0_5_37_real,
  output     [15:0]   io_coef_out_payload_0_5_37_imag,
  output     [15:0]   io_coef_out_payload_0_5_38_real,
  output     [15:0]   io_coef_out_payload_0_5_38_imag,
  output     [15:0]   io_coef_out_payload_0_5_39_real,
  output     [15:0]   io_coef_out_payload_0_5_39_imag,
  output     [15:0]   io_coef_out_payload_0_5_40_real,
  output     [15:0]   io_coef_out_payload_0_5_40_imag,
  output     [15:0]   io_coef_out_payload_0_5_41_real,
  output     [15:0]   io_coef_out_payload_0_5_41_imag,
  output     [15:0]   io_coef_out_payload_0_5_42_real,
  output     [15:0]   io_coef_out_payload_0_5_42_imag,
  output     [15:0]   io_coef_out_payload_0_5_43_real,
  output     [15:0]   io_coef_out_payload_0_5_43_imag,
  output     [15:0]   io_coef_out_payload_0_5_44_real,
  output     [15:0]   io_coef_out_payload_0_5_44_imag,
  output     [15:0]   io_coef_out_payload_0_5_45_real,
  output     [15:0]   io_coef_out_payload_0_5_45_imag,
  output     [15:0]   io_coef_out_payload_0_5_46_real,
  output     [15:0]   io_coef_out_payload_0_5_46_imag,
  output     [15:0]   io_coef_out_payload_0_5_47_real,
  output     [15:0]   io_coef_out_payload_0_5_47_imag,
  output     [15:0]   io_coef_out_payload_0_5_48_real,
  output     [15:0]   io_coef_out_payload_0_5_48_imag,
  output     [15:0]   io_coef_out_payload_0_5_49_real,
  output     [15:0]   io_coef_out_payload_0_5_49_imag,
  output     [15:0]   io_coef_out_payload_0_6_0_real,
  output     [15:0]   io_coef_out_payload_0_6_0_imag,
  output     [15:0]   io_coef_out_payload_0_6_1_real,
  output     [15:0]   io_coef_out_payload_0_6_1_imag,
  output     [15:0]   io_coef_out_payload_0_6_2_real,
  output     [15:0]   io_coef_out_payload_0_6_2_imag,
  output     [15:0]   io_coef_out_payload_0_6_3_real,
  output     [15:0]   io_coef_out_payload_0_6_3_imag,
  output     [15:0]   io_coef_out_payload_0_6_4_real,
  output     [15:0]   io_coef_out_payload_0_6_4_imag,
  output     [15:0]   io_coef_out_payload_0_6_5_real,
  output     [15:0]   io_coef_out_payload_0_6_5_imag,
  output     [15:0]   io_coef_out_payload_0_6_6_real,
  output     [15:0]   io_coef_out_payload_0_6_6_imag,
  output     [15:0]   io_coef_out_payload_0_6_7_real,
  output     [15:0]   io_coef_out_payload_0_6_7_imag,
  output     [15:0]   io_coef_out_payload_0_6_8_real,
  output     [15:0]   io_coef_out_payload_0_6_8_imag,
  output     [15:0]   io_coef_out_payload_0_6_9_real,
  output     [15:0]   io_coef_out_payload_0_6_9_imag,
  output     [15:0]   io_coef_out_payload_0_6_10_real,
  output     [15:0]   io_coef_out_payload_0_6_10_imag,
  output     [15:0]   io_coef_out_payload_0_6_11_real,
  output     [15:0]   io_coef_out_payload_0_6_11_imag,
  output     [15:0]   io_coef_out_payload_0_6_12_real,
  output     [15:0]   io_coef_out_payload_0_6_12_imag,
  output     [15:0]   io_coef_out_payload_0_6_13_real,
  output     [15:0]   io_coef_out_payload_0_6_13_imag,
  output     [15:0]   io_coef_out_payload_0_6_14_real,
  output     [15:0]   io_coef_out_payload_0_6_14_imag,
  output     [15:0]   io_coef_out_payload_0_6_15_real,
  output     [15:0]   io_coef_out_payload_0_6_15_imag,
  output     [15:0]   io_coef_out_payload_0_6_16_real,
  output     [15:0]   io_coef_out_payload_0_6_16_imag,
  output     [15:0]   io_coef_out_payload_0_6_17_real,
  output     [15:0]   io_coef_out_payload_0_6_17_imag,
  output     [15:0]   io_coef_out_payload_0_6_18_real,
  output     [15:0]   io_coef_out_payload_0_6_18_imag,
  output     [15:0]   io_coef_out_payload_0_6_19_real,
  output     [15:0]   io_coef_out_payload_0_6_19_imag,
  output     [15:0]   io_coef_out_payload_0_6_20_real,
  output     [15:0]   io_coef_out_payload_0_6_20_imag,
  output     [15:0]   io_coef_out_payload_0_6_21_real,
  output     [15:0]   io_coef_out_payload_0_6_21_imag,
  output     [15:0]   io_coef_out_payload_0_6_22_real,
  output     [15:0]   io_coef_out_payload_0_6_22_imag,
  output     [15:0]   io_coef_out_payload_0_6_23_real,
  output     [15:0]   io_coef_out_payload_0_6_23_imag,
  output     [15:0]   io_coef_out_payload_0_6_24_real,
  output     [15:0]   io_coef_out_payload_0_6_24_imag,
  output     [15:0]   io_coef_out_payload_0_6_25_real,
  output     [15:0]   io_coef_out_payload_0_6_25_imag,
  output     [15:0]   io_coef_out_payload_0_6_26_real,
  output     [15:0]   io_coef_out_payload_0_6_26_imag,
  output     [15:0]   io_coef_out_payload_0_6_27_real,
  output     [15:0]   io_coef_out_payload_0_6_27_imag,
  output     [15:0]   io_coef_out_payload_0_6_28_real,
  output     [15:0]   io_coef_out_payload_0_6_28_imag,
  output     [15:0]   io_coef_out_payload_0_6_29_real,
  output     [15:0]   io_coef_out_payload_0_6_29_imag,
  output     [15:0]   io_coef_out_payload_0_6_30_real,
  output     [15:0]   io_coef_out_payload_0_6_30_imag,
  output     [15:0]   io_coef_out_payload_0_6_31_real,
  output     [15:0]   io_coef_out_payload_0_6_31_imag,
  output     [15:0]   io_coef_out_payload_0_6_32_real,
  output     [15:0]   io_coef_out_payload_0_6_32_imag,
  output     [15:0]   io_coef_out_payload_0_6_33_real,
  output     [15:0]   io_coef_out_payload_0_6_33_imag,
  output     [15:0]   io_coef_out_payload_0_6_34_real,
  output     [15:0]   io_coef_out_payload_0_6_34_imag,
  output     [15:0]   io_coef_out_payload_0_6_35_real,
  output     [15:0]   io_coef_out_payload_0_6_35_imag,
  output     [15:0]   io_coef_out_payload_0_6_36_real,
  output     [15:0]   io_coef_out_payload_0_6_36_imag,
  output     [15:0]   io_coef_out_payload_0_6_37_real,
  output     [15:0]   io_coef_out_payload_0_6_37_imag,
  output     [15:0]   io_coef_out_payload_0_6_38_real,
  output     [15:0]   io_coef_out_payload_0_6_38_imag,
  output     [15:0]   io_coef_out_payload_0_6_39_real,
  output     [15:0]   io_coef_out_payload_0_6_39_imag,
  output     [15:0]   io_coef_out_payload_0_6_40_real,
  output     [15:0]   io_coef_out_payload_0_6_40_imag,
  output     [15:0]   io_coef_out_payload_0_6_41_real,
  output     [15:0]   io_coef_out_payload_0_6_41_imag,
  output     [15:0]   io_coef_out_payload_0_6_42_real,
  output     [15:0]   io_coef_out_payload_0_6_42_imag,
  output     [15:0]   io_coef_out_payload_0_6_43_real,
  output     [15:0]   io_coef_out_payload_0_6_43_imag,
  output     [15:0]   io_coef_out_payload_0_6_44_real,
  output     [15:0]   io_coef_out_payload_0_6_44_imag,
  output     [15:0]   io_coef_out_payload_0_6_45_real,
  output     [15:0]   io_coef_out_payload_0_6_45_imag,
  output     [15:0]   io_coef_out_payload_0_6_46_real,
  output     [15:0]   io_coef_out_payload_0_6_46_imag,
  output     [15:0]   io_coef_out_payload_0_6_47_real,
  output     [15:0]   io_coef_out_payload_0_6_47_imag,
  output     [15:0]   io_coef_out_payload_0_6_48_real,
  output     [15:0]   io_coef_out_payload_0_6_48_imag,
  output     [15:0]   io_coef_out_payload_0_6_49_real,
  output     [15:0]   io_coef_out_payload_0_6_49_imag,
  output     [15:0]   io_coef_out_payload_0_7_0_real,
  output     [15:0]   io_coef_out_payload_0_7_0_imag,
  output     [15:0]   io_coef_out_payload_0_7_1_real,
  output     [15:0]   io_coef_out_payload_0_7_1_imag,
  output     [15:0]   io_coef_out_payload_0_7_2_real,
  output     [15:0]   io_coef_out_payload_0_7_2_imag,
  output     [15:0]   io_coef_out_payload_0_7_3_real,
  output     [15:0]   io_coef_out_payload_0_7_3_imag,
  output     [15:0]   io_coef_out_payload_0_7_4_real,
  output     [15:0]   io_coef_out_payload_0_7_4_imag,
  output     [15:0]   io_coef_out_payload_0_7_5_real,
  output     [15:0]   io_coef_out_payload_0_7_5_imag,
  output     [15:0]   io_coef_out_payload_0_7_6_real,
  output     [15:0]   io_coef_out_payload_0_7_6_imag,
  output     [15:0]   io_coef_out_payload_0_7_7_real,
  output     [15:0]   io_coef_out_payload_0_7_7_imag,
  output     [15:0]   io_coef_out_payload_0_7_8_real,
  output     [15:0]   io_coef_out_payload_0_7_8_imag,
  output     [15:0]   io_coef_out_payload_0_7_9_real,
  output     [15:0]   io_coef_out_payload_0_7_9_imag,
  output     [15:0]   io_coef_out_payload_0_7_10_real,
  output     [15:0]   io_coef_out_payload_0_7_10_imag,
  output     [15:0]   io_coef_out_payload_0_7_11_real,
  output     [15:0]   io_coef_out_payload_0_7_11_imag,
  output     [15:0]   io_coef_out_payload_0_7_12_real,
  output     [15:0]   io_coef_out_payload_0_7_12_imag,
  output     [15:0]   io_coef_out_payload_0_7_13_real,
  output     [15:0]   io_coef_out_payload_0_7_13_imag,
  output     [15:0]   io_coef_out_payload_0_7_14_real,
  output     [15:0]   io_coef_out_payload_0_7_14_imag,
  output     [15:0]   io_coef_out_payload_0_7_15_real,
  output     [15:0]   io_coef_out_payload_0_7_15_imag,
  output     [15:0]   io_coef_out_payload_0_7_16_real,
  output     [15:0]   io_coef_out_payload_0_7_16_imag,
  output     [15:0]   io_coef_out_payload_0_7_17_real,
  output     [15:0]   io_coef_out_payload_0_7_17_imag,
  output     [15:0]   io_coef_out_payload_0_7_18_real,
  output     [15:0]   io_coef_out_payload_0_7_18_imag,
  output     [15:0]   io_coef_out_payload_0_7_19_real,
  output     [15:0]   io_coef_out_payload_0_7_19_imag,
  output     [15:0]   io_coef_out_payload_0_7_20_real,
  output     [15:0]   io_coef_out_payload_0_7_20_imag,
  output     [15:0]   io_coef_out_payload_0_7_21_real,
  output     [15:0]   io_coef_out_payload_0_7_21_imag,
  output     [15:0]   io_coef_out_payload_0_7_22_real,
  output     [15:0]   io_coef_out_payload_0_7_22_imag,
  output     [15:0]   io_coef_out_payload_0_7_23_real,
  output     [15:0]   io_coef_out_payload_0_7_23_imag,
  output     [15:0]   io_coef_out_payload_0_7_24_real,
  output     [15:0]   io_coef_out_payload_0_7_24_imag,
  output     [15:0]   io_coef_out_payload_0_7_25_real,
  output     [15:0]   io_coef_out_payload_0_7_25_imag,
  output     [15:0]   io_coef_out_payload_0_7_26_real,
  output     [15:0]   io_coef_out_payload_0_7_26_imag,
  output     [15:0]   io_coef_out_payload_0_7_27_real,
  output     [15:0]   io_coef_out_payload_0_7_27_imag,
  output     [15:0]   io_coef_out_payload_0_7_28_real,
  output     [15:0]   io_coef_out_payload_0_7_28_imag,
  output     [15:0]   io_coef_out_payload_0_7_29_real,
  output     [15:0]   io_coef_out_payload_0_7_29_imag,
  output     [15:0]   io_coef_out_payload_0_7_30_real,
  output     [15:0]   io_coef_out_payload_0_7_30_imag,
  output     [15:0]   io_coef_out_payload_0_7_31_real,
  output     [15:0]   io_coef_out_payload_0_7_31_imag,
  output     [15:0]   io_coef_out_payload_0_7_32_real,
  output     [15:0]   io_coef_out_payload_0_7_32_imag,
  output     [15:0]   io_coef_out_payload_0_7_33_real,
  output     [15:0]   io_coef_out_payload_0_7_33_imag,
  output     [15:0]   io_coef_out_payload_0_7_34_real,
  output     [15:0]   io_coef_out_payload_0_7_34_imag,
  output     [15:0]   io_coef_out_payload_0_7_35_real,
  output     [15:0]   io_coef_out_payload_0_7_35_imag,
  output     [15:0]   io_coef_out_payload_0_7_36_real,
  output     [15:0]   io_coef_out_payload_0_7_36_imag,
  output     [15:0]   io_coef_out_payload_0_7_37_real,
  output     [15:0]   io_coef_out_payload_0_7_37_imag,
  output     [15:0]   io_coef_out_payload_0_7_38_real,
  output     [15:0]   io_coef_out_payload_0_7_38_imag,
  output     [15:0]   io_coef_out_payload_0_7_39_real,
  output     [15:0]   io_coef_out_payload_0_7_39_imag,
  output     [15:0]   io_coef_out_payload_0_7_40_real,
  output     [15:0]   io_coef_out_payload_0_7_40_imag,
  output     [15:0]   io_coef_out_payload_0_7_41_real,
  output     [15:0]   io_coef_out_payload_0_7_41_imag,
  output     [15:0]   io_coef_out_payload_0_7_42_real,
  output     [15:0]   io_coef_out_payload_0_7_42_imag,
  output     [15:0]   io_coef_out_payload_0_7_43_real,
  output     [15:0]   io_coef_out_payload_0_7_43_imag,
  output     [15:0]   io_coef_out_payload_0_7_44_real,
  output     [15:0]   io_coef_out_payload_0_7_44_imag,
  output     [15:0]   io_coef_out_payload_0_7_45_real,
  output     [15:0]   io_coef_out_payload_0_7_45_imag,
  output     [15:0]   io_coef_out_payload_0_7_46_real,
  output     [15:0]   io_coef_out_payload_0_7_46_imag,
  output     [15:0]   io_coef_out_payload_0_7_47_real,
  output     [15:0]   io_coef_out_payload_0_7_47_imag,
  output     [15:0]   io_coef_out_payload_0_7_48_real,
  output     [15:0]   io_coef_out_payload_0_7_48_imag,
  output     [15:0]   io_coef_out_payload_0_7_49_real,
  output     [15:0]   io_coef_out_payload_0_7_49_imag,
  output     [15:0]   io_coef_out_payload_0_8_0_real,
  output     [15:0]   io_coef_out_payload_0_8_0_imag,
  output     [15:0]   io_coef_out_payload_0_8_1_real,
  output     [15:0]   io_coef_out_payload_0_8_1_imag,
  output     [15:0]   io_coef_out_payload_0_8_2_real,
  output     [15:0]   io_coef_out_payload_0_8_2_imag,
  output     [15:0]   io_coef_out_payload_0_8_3_real,
  output     [15:0]   io_coef_out_payload_0_8_3_imag,
  output     [15:0]   io_coef_out_payload_0_8_4_real,
  output     [15:0]   io_coef_out_payload_0_8_4_imag,
  output     [15:0]   io_coef_out_payload_0_8_5_real,
  output     [15:0]   io_coef_out_payload_0_8_5_imag,
  output     [15:0]   io_coef_out_payload_0_8_6_real,
  output     [15:0]   io_coef_out_payload_0_8_6_imag,
  output     [15:0]   io_coef_out_payload_0_8_7_real,
  output     [15:0]   io_coef_out_payload_0_8_7_imag,
  output     [15:0]   io_coef_out_payload_0_8_8_real,
  output     [15:0]   io_coef_out_payload_0_8_8_imag,
  output     [15:0]   io_coef_out_payload_0_8_9_real,
  output     [15:0]   io_coef_out_payload_0_8_9_imag,
  output     [15:0]   io_coef_out_payload_0_8_10_real,
  output     [15:0]   io_coef_out_payload_0_8_10_imag,
  output     [15:0]   io_coef_out_payload_0_8_11_real,
  output     [15:0]   io_coef_out_payload_0_8_11_imag,
  output     [15:0]   io_coef_out_payload_0_8_12_real,
  output     [15:0]   io_coef_out_payload_0_8_12_imag,
  output     [15:0]   io_coef_out_payload_0_8_13_real,
  output     [15:0]   io_coef_out_payload_0_8_13_imag,
  output     [15:0]   io_coef_out_payload_0_8_14_real,
  output     [15:0]   io_coef_out_payload_0_8_14_imag,
  output     [15:0]   io_coef_out_payload_0_8_15_real,
  output     [15:0]   io_coef_out_payload_0_8_15_imag,
  output     [15:0]   io_coef_out_payload_0_8_16_real,
  output     [15:0]   io_coef_out_payload_0_8_16_imag,
  output     [15:0]   io_coef_out_payload_0_8_17_real,
  output     [15:0]   io_coef_out_payload_0_8_17_imag,
  output     [15:0]   io_coef_out_payload_0_8_18_real,
  output     [15:0]   io_coef_out_payload_0_8_18_imag,
  output     [15:0]   io_coef_out_payload_0_8_19_real,
  output     [15:0]   io_coef_out_payload_0_8_19_imag,
  output     [15:0]   io_coef_out_payload_0_8_20_real,
  output     [15:0]   io_coef_out_payload_0_8_20_imag,
  output     [15:0]   io_coef_out_payload_0_8_21_real,
  output     [15:0]   io_coef_out_payload_0_8_21_imag,
  output     [15:0]   io_coef_out_payload_0_8_22_real,
  output     [15:0]   io_coef_out_payload_0_8_22_imag,
  output     [15:0]   io_coef_out_payload_0_8_23_real,
  output     [15:0]   io_coef_out_payload_0_8_23_imag,
  output     [15:0]   io_coef_out_payload_0_8_24_real,
  output     [15:0]   io_coef_out_payload_0_8_24_imag,
  output     [15:0]   io_coef_out_payload_0_8_25_real,
  output     [15:0]   io_coef_out_payload_0_8_25_imag,
  output     [15:0]   io_coef_out_payload_0_8_26_real,
  output     [15:0]   io_coef_out_payload_0_8_26_imag,
  output     [15:0]   io_coef_out_payload_0_8_27_real,
  output     [15:0]   io_coef_out_payload_0_8_27_imag,
  output     [15:0]   io_coef_out_payload_0_8_28_real,
  output     [15:0]   io_coef_out_payload_0_8_28_imag,
  output     [15:0]   io_coef_out_payload_0_8_29_real,
  output     [15:0]   io_coef_out_payload_0_8_29_imag,
  output     [15:0]   io_coef_out_payload_0_8_30_real,
  output     [15:0]   io_coef_out_payload_0_8_30_imag,
  output     [15:0]   io_coef_out_payload_0_8_31_real,
  output     [15:0]   io_coef_out_payload_0_8_31_imag,
  output     [15:0]   io_coef_out_payload_0_8_32_real,
  output     [15:0]   io_coef_out_payload_0_8_32_imag,
  output     [15:0]   io_coef_out_payload_0_8_33_real,
  output     [15:0]   io_coef_out_payload_0_8_33_imag,
  output     [15:0]   io_coef_out_payload_0_8_34_real,
  output     [15:0]   io_coef_out_payload_0_8_34_imag,
  output     [15:0]   io_coef_out_payload_0_8_35_real,
  output     [15:0]   io_coef_out_payload_0_8_35_imag,
  output     [15:0]   io_coef_out_payload_0_8_36_real,
  output     [15:0]   io_coef_out_payload_0_8_36_imag,
  output     [15:0]   io_coef_out_payload_0_8_37_real,
  output     [15:0]   io_coef_out_payload_0_8_37_imag,
  output     [15:0]   io_coef_out_payload_0_8_38_real,
  output     [15:0]   io_coef_out_payload_0_8_38_imag,
  output     [15:0]   io_coef_out_payload_0_8_39_real,
  output     [15:0]   io_coef_out_payload_0_8_39_imag,
  output     [15:0]   io_coef_out_payload_0_8_40_real,
  output     [15:0]   io_coef_out_payload_0_8_40_imag,
  output     [15:0]   io_coef_out_payload_0_8_41_real,
  output     [15:0]   io_coef_out_payload_0_8_41_imag,
  output     [15:0]   io_coef_out_payload_0_8_42_real,
  output     [15:0]   io_coef_out_payload_0_8_42_imag,
  output     [15:0]   io_coef_out_payload_0_8_43_real,
  output     [15:0]   io_coef_out_payload_0_8_43_imag,
  output     [15:0]   io_coef_out_payload_0_8_44_real,
  output     [15:0]   io_coef_out_payload_0_8_44_imag,
  output     [15:0]   io_coef_out_payload_0_8_45_real,
  output     [15:0]   io_coef_out_payload_0_8_45_imag,
  output     [15:0]   io_coef_out_payload_0_8_46_real,
  output     [15:0]   io_coef_out_payload_0_8_46_imag,
  output     [15:0]   io_coef_out_payload_0_8_47_real,
  output     [15:0]   io_coef_out_payload_0_8_47_imag,
  output     [15:0]   io_coef_out_payload_0_8_48_real,
  output     [15:0]   io_coef_out_payload_0_8_48_imag,
  output     [15:0]   io_coef_out_payload_0_8_49_real,
  output     [15:0]   io_coef_out_payload_0_8_49_imag,
  output     [15:0]   io_coef_out_payload_0_9_0_real,
  output     [15:0]   io_coef_out_payload_0_9_0_imag,
  output     [15:0]   io_coef_out_payload_0_9_1_real,
  output     [15:0]   io_coef_out_payload_0_9_1_imag,
  output     [15:0]   io_coef_out_payload_0_9_2_real,
  output     [15:0]   io_coef_out_payload_0_9_2_imag,
  output     [15:0]   io_coef_out_payload_0_9_3_real,
  output     [15:0]   io_coef_out_payload_0_9_3_imag,
  output     [15:0]   io_coef_out_payload_0_9_4_real,
  output     [15:0]   io_coef_out_payload_0_9_4_imag,
  output     [15:0]   io_coef_out_payload_0_9_5_real,
  output     [15:0]   io_coef_out_payload_0_9_5_imag,
  output     [15:0]   io_coef_out_payload_0_9_6_real,
  output     [15:0]   io_coef_out_payload_0_9_6_imag,
  output     [15:0]   io_coef_out_payload_0_9_7_real,
  output     [15:0]   io_coef_out_payload_0_9_7_imag,
  output     [15:0]   io_coef_out_payload_0_9_8_real,
  output     [15:0]   io_coef_out_payload_0_9_8_imag,
  output     [15:0]   io_coef_out_payload_0_9_9_real,
  output     [15:0]   io_coef_out_payload_0_9_9_imag,
  output     [15:0]   io_coef_out_payload_0_9_10_real,
  output     [15:0]   io_coef_out_payload_0_9_10_imag,
  output     [15:0]   io_coef_out_payload_0_9_11_real,
  output     [15:0]   io_coef_out_payload_0_9_11_imag,
  output     [15:0]   io_coef_out_payload_0_9_12_real,
  output     [15:0]   io_coef_out_payload_0_9_12_imag,
  output     [15:0]   io_coef_out_payload_0_9_13_real,
  output     [15:0]   io_coef_out_payload_0_9_13_imag,
  output     [15:0]   io_coef_out_payload_0_9_14_real,
  output     [15:0]   io_coef_out_payload_0_9_14_imag,
  output     [15:0]   io_coef_out_payload_0_9_15_real,
  output     [15:0]   io_coef_out_payload_0_9_15_imag,
  output     [15:0]   io_coef_out_payload_0_9_16_real,
  output     [15:0]   io_coef_out_payload_0_9_16_imag,
  output     [15:0]   io_coef_out_payload_0_9_17_real,
  output     [15:0]   io_coef_out_payload_0_9_17_imag,
  output     [15:0]   io_coef_out_payload_0_9_18_real,
  output     [15:0]   io_coef_out_payload_0_9_18_imag,
  output     [15:0]   io_coef_out_payload_0_9_19_real,
  output     [15:0]   io_coef_out_payload_0_9_19_imag,
  output     [15:0]   io_coef_out_payload_0_9_20_real,
  output     [15:0]   io_coef_out_payload_0_9_20_imag,
  output     [15:0]   io_coef_out_payload_0_9_21_real,
  output     [15:0]   io_coef_out_payload_0_9_21_imag,
  output     [15:0]   io_coef_out_payload_0_9_22_real,
  output     [15:0]   io_coef_out_payload_0_9_22_imag,
  output     [15:0]   io_coef_out_payload_0_9_23_real,
  output     [15:0]   io_coef_out_payload_0_9_23_imag,
  output     [15:0]   io_coef_out_payload_0_9_24_real,
  output     [15:0]   io_coef_out_payload_0_9_24_imag,
  output     [15:0]   io_coef_out_payload_0_9_25_real,
  output     [15:0]   io_coef_out_payload_0_9_25_imag,
  output     [15:0]   io_coef_out_payload_0_9_26_real,
  output     [15:0]   io_coef_out_payload_0_9_26_imag,
  output     [15:0]   io_coef_out_payload_0_9_27_real,
  output     [15:0]   io_coef_out_payload_0_9_27_imag,
  output     [15:0]   io_coef_out_payload_0_9_28_real,
  output     [15:0]   io_coef_out_payload_0_9_28_imag,
  output     [15:0]   io_coef_out_payload_0_9_29_real,
  output     [15:0]   io_coef_out_payload_0_9_29_imag,
  output     [15:0]   io_coef_out_payload_0_9_30_real,
  output     [15:0]   io_coef_out_payload_0_9_30_imag,
  output     [15:0]   io_coef_out_payload_0_9_31_real,
  output     [15:0]   io_coef_out_payload_0_9_31_imag,
  output     [15:0]   io_coef_out_payload_0_9_32_real,
  output     [15:0]   io_coef_out_payload_0_9_32_imag,
  output     [15:0]   io_coef_out_payload_0_9_33_real,
  output     [15:0]   io_coef_out_payload_0_9_33_imag,
  output     [15:0]   io_coef_out_payload_0_9_34_real,
  output     [15:0]   io_coef_out_payload_0_9_34_imag,
  output     [15:0]   io_coef_out_payload_0_9_35_real,
  output     [15:0]   io_coef_out_payload_0_9_35_imag,
  output     [15:0]   io_coef_out_payload_0_9_36_real,
  output     [15:0]   io_coef_out_payload_0_9_36_imag,
  output     [15:0]   io_coef_out_payload_0_9_37_real,
  output     [15:0]   io_coef_out_payload_0_9_37_imag,
  output     [15:0]   io_coef_out_payload_0_9_38_real,
  output     [15:0]   io_coef_out_payload_0_9_38_imag,
  output     [15:0]   io_coef_out_payload_0_9_39_real,
  output     [15:0]   io_coef_out_payload_0_9_39_imag,
  output     [15:0]   io_coef_out_payload_0_9_40_real,
  output     [15:0]   io_coef_out_payload_0_9_40_imag,
  output     [15:0]   io_coef_out_payload_0_9_41_real,
  output     [15:0]   io_coef_out_payload_0_9_41_imag,
  output     [15:0]   io_coef_out_payload_0_9_42_real,
  output     [15:0]   io_coef_out_payload_0_9_42_imag,
  output     [15:0]   io_coef_out_payload_0_9_43_real,
  output     [15:0]   io_coef_out_payload_0_9_43_imag,
  output     [15:0]   io_coef_out_payload_0_9_44_real,
  output     [15:0]   io_coef_out_payload_0_9_44_imag,
  output     [15:0]   io_coef_out_payload_0_9_45_real,
  output     [15:0]   io_coef_out_payload_0_9_45_imag,
  output     [15:0]   io_coef_out_payload_0_9_46_real,
  output     [15:0]   io_coef_out_payload_0_9_46_imag,
  output     [15:0]   io_coef_out_payload_0_9_47_real,
  output     [15:0]   io_coef_out_payload_0_9_47_imag,
  output     [15:0]   io_coef_out_payload_0_9_48_real,
  output     [15:0]   io_coef_out_payload_0_9_48_imag,
  output     [15:0]   io_coef_out_payload_0_9_49_real,
  output     [15:0]   io_coef_out_payload_0_9_49_imag,
  output     [15:0]   io_coef_out_payload_0_10_0_real,
  output     [15:0]   io_coef_out_payload_0_10_0_imag,
  output     [15:0]   io_coef_out_payload_0_10_1_real,
  output     [15:0]   io_coef_out_payload_0_10_1_imag,
  output     [15:0]   io_coef_out_payload_0_10_2_real,
  output     [15:0]   io_coef_out_payload_0_10_2_imag,
  output     [15:0]   io_coef_out_payload_0_10_3_real,
  output     [15:0]   io_coef_out_payload_0_10_3_imag,
  output     [15:0]   io_coef_out_payload_0_10_4_real,
  output     [15:0]   io_coef_out_payload_0_10_4_imag,
  output     [15:0]   io_coef_out_payload_0_10_5_real,
  output     [15:0]   io_coef_out_payload_0_10_5_imag,
  output     [15:0]   io_coef_out_payload_0_10_6_real,
  output     [15:0]   io_coef_out_payload_0_10_6_imag,
  output     [15:0]   io_coef_out_payload_0_10_7_real,
  output     [15:0]   io_coef_out_payload_0_10_7_imag,
  output     [15:0]   io_coef_out_payload_0_10_8_real,
  output     [15:0]   io_coef_out_payload_0_10_8_imag,
  output     [15:0]   io_coef_out_payload_0_10_9_real,
  output     [15:0]   io_coef_out_payload_0_10_9_imag,
  output     [15:0]   io_coef_out_payload_0_10_10_real,
  output     [15:0]   io_coef_out_payload_0_10_10_imag,
  output     [15:0]   io_coef_out_payload_0_10_11_real,
  output     [15:0]   io_coef_out_payload_0_10_11_imag,
  output     [15:0]   io_coef_out_payload_0_10_12_real,
  output     [15:0]   io_coef_out_payload_0_10_12_imag,
  output     [15:0]   io_coef_out_payload_0_10_13_real,
  output     [15:0]   io_coef_out_payload_0_10_13_imag,
  output     [15:0]   io_coef_out_payload_0_10_14_real,
  output     [15:0]   io_coef_out_payload_0_10_14_imag,
  output     [15:0]   io_coef_out_payload_0_10_15_real,
  output     [15:0]   io_coef_out_payload_0_10_15_imag,
  output     [15:0]   io_coef_out_payload_0_10_16_real,
  output     [15:0]   io_coef_out_payload_0_10_16_imag,
  output     [15:0]   io_coef_out_payload_0_10_17_real,
  output     [15:0]   io_coef_out_payload_0_10_17_imag,
  output     [15:0]   io_coef_out_payload_0_10_18_real,
  output     [15:0]   io_coef_out_payload_0_10_18_imag,
  output     [15:0]   io_coef_out_payload_0_10_19_real,
  output     [15:0]   io_coef_out_payload_0_10_19_imag,
  output     [15:0]   io_coef_out_payload_0_10_20_real,
  output     [15:0]   io_coef_out_payload_0_10_20_imag,
  output     [15:0]   io_coef_out_payload_0_10_21_real,
  output     [15:0]   io_coef_out_payload_0_10_21_imag,
  output     [15:0]   io_coef_out_payload_0_10_22_real,
  output     [15:0]   io_coef_out_payload_0_10_22_imag,
  output     [15:0]   io_coef_out_payload_0_10_23_real,
  output     [15:0]   io_coef_out_payload_0_10_23_imag,
  output     [15:0]   io_coef_out_payload_0_10_24_real,
  output     [15:0]   io_coef_out_payload_0_10_24_imag,
  output     [15:0]   io_coef_out_payload_0_10_25_real,
  output     [15:0]   io_coef_out_payload_0_10_25_imag,
  output     [15:0]   io_coef_out_payload_0_10_26_real,
  output     [15:0]   io_coef_out_payload_0_10_26_imag,
  output     [15:0]   io_coef_out_payload_0_10_27_real,
  output     [15:0]   io_coef_out_payload_0_10_27_imag,
  output     [15:0]   io_coef_out_payload_0_10_28_real,
  output     [15:0]   io_coef_out_payload_0_10_28_imag,
  output     [15:0]   io_coef_out_payload_0_10_29_real,
  output     [15:0]   io_coef_out_payload_0_10_29_imag,
  output     [15:0]   io_coef_out_payload_0_10_30_real,
  output     [15:0]   io_coef_out_payload_0_10_30_imag,
  output     [15:0]   io_coef_out_payload_0_10_31_real,
  output     [15:0]   io_coef_out_payload_0_10_31_imag,
  output     [15:0]   io_coef_out_payload_0_10_32_real,
  output     [15:0]   io_coef_out_payload_0_10_32_imag,
  output     [15:0]   io_coef_out_payload_0_10_33_real,
  output     [15:0]   io_coef_out_payload_0_10_33_imag,
  output     [15:0]   io_coef_out_payload_0_10_34_real,
  output     [15:0]   io_coef_out_payload_0_10_34_imag,
  output     [15:0]   io_coef_out_payload_0_10_35_real,
  output     [15:0]   io_coef_out_payload_0_10_35_imag,
  output     [15:0]   io_coef_out_payload_0_10_36_real,
  output     [15:0]   io_coef_out_payload_0_10_36_imag,
  output     [15:0]   io_coef_out_payload_0_10_37_real,
  output     [15:0]   io_coef_out_payload_0_10_37_imag,
  output     [15:0]   io_coef_out_payload_0_10_38_real,
  output     [15:0]   io_coef_out_payload_0_10_38_imag,
  output     [15:0]   io_coef_out_payload_0_10_39_real,
  output     [15:0]   io_coef_out_payload_0_10_39_imag,
  output     [15:0]   io_coef_out_payload_0_10_40_real,
  output     [15:0]   io_coef_out_payload_0_10_40_imag,
  output     [15:0]   io_coef_out_payload_0_10_41_real,
  output     [15:0]   io_coef_out_payload_0_10_41_imag,
  output     [15:0]   io_coef_out_payload_0_10_42_real,
  output     [15:0]   io_coef_out_payload_0_10_42_imag,
  output     [15:0]   io_coef_out_payload_0_10_43_real,
  output     [15:0]   io_coef_out_payload_0_10_43_imag,
  output     [15:0]   io_coef_out_payload_0_10_44_real,
  output     [15:0]   io_coef_out_payload_0_10_44_imag,
  output     [15:0]   io_coef_out_payload_0_10_45_real,
  output     [15:0]   io_coef_out_payload_0_10_45_imag,
  output     [15:0]   io_coef_out_payload_0_10_46_real,
  output     [15:0]   io_coef_out_payload_0_10_46_imag,
  output     [15:0]   io_coef_out_payload_0_10_47_real,
  output     [15:0]   io_coef_out_payload_0_10_47_imag,
  output     [15:0]   io_coef_out_payload_0_10_48_real,
  output     [15:0]   io_coef_out_payload_0_10_48_imag,
  output     [15:0]   io_coef_out_payload_0_10_49_real,
  output     [15:0]   io_coef_out_payload_0_10_49_imag,
  output     [15:0]   io_coef_out_payload_0_11_0_real,
  output     [15:0]   io_coef_out_payload_0_11_0_imag,
  output     [15:0]   io_coef_out_payload_0_11_1_real,
  output     [15:0]   io_coef_out_payload_0_11_1_imag,
  output     [15:0]   io_coef_out_payload_0_11_2_real,
  output     [15:0]   io_coef_out_payload_0_11_2_imag,
  output     [15:0]   io_coef_out_payload_0_11_3_real,
  output     [15:0]   io_coef_out_payload_0_11_3_imag,
  output     [15:0]   io_coef_out_payload_0_11_4_real,
  output     [15:0]   io_coef_out_payload_0_11_4_imag,
  output     [15:0]   io_coef_out_payload_0_11_5_real,
  output     [15:0]   io_coef_out_payload_0_11_5_imag,
  output     [15:0]   io_coef_out_payload_0_11_6_real,
  output     [15:0]   io_coef_out_payload_0_11_6_imag,
  output     [15:0]   io_coef_out_payload_0_11_7_real,
  output     [15:0]   io_coef_out_payload_0_11_7_imag,
  output     [15:0]   io_coef_out_payload_0_11_8_real,
  output     [15:0]   io_coef_out_payload_0_11_8_imag,
  output     [15:0]   io_coef_out_payload_0_11_9_real,
  output     [15:0]   io_coef_out_payload_0_11_9_imag,
  output     [15:0]   io_coef_out_payload_0_11_10_real,
  output     [15:0]   io_coef_out_payload_0_11_10_imag,
  output     [15:0]   io_coef_out_payload_0_11_11_real,
  output     [15:0]   io_coef_out_payload_0_11_11_imag,
  output     [15:0]   io_coef_out_payload_0_11_12_real,
  output     [15:0]   io_coef_out_payload_0_11_12_imag,
  output     [15:0]   io_coef_out_payload_0_11_13_real,
  output     [15:0]   io_coef_out_payload_0_11_13_imag,
  output     [15:0]   io_coef_out_payload_0_11_14_real,
  output     [15:0]   io_coef_out_payload_0_11_14_imag,
  output     [15:0]   io_coef_out_payload_0_11_15_real,
  output     [15:0]   io_coef_out_payload_0_11_15_imag,
  output     [15:0]   io_coef_out_payload_0_11_16_real,
  output     [15:0]   io_coef_out_payload_0_11_16_imag,
  output     [15:0]   io_coef_out_payload_0_11_17_real,
  output     [15:0]   io_coef_out_payload_0_11_17_imag,
  output     [15:0]   io_coef_out_payload_0_11_18_real,
  output     [15:0]   io_coef_out_payload_0_11_18_imag,
  output     [15:0]   io_coef_out_payload_0_11_19_real,
  output     [15:0]   io_coef_out_payload_0_11_19_imag,
  output     [15:0]   io_coef_out_payload_0_11_20_real,
  output     [15:0]   io_coef_out_payload_0_11_20_imag,
  output     [15:0]   io_coef_out_payload_0_11_21_real,
  output     [15:0]   io_coef_out_payload_0_11_21_imag,
  output     [15:0]   io_coef_out_payload_0_11_22_real,
  output     [15:0]   io_coef_out_payload_0_11_22_imag,
  output     [15:0]   io_coef_out_payload_0_11_23_real,
  output     [15:0]   io_coef_out_payload_0_11_23_imag,
  output     [15:0]   io_coef_out_payload_0_11_24_real,
  output     [15:0]   io_coef_out_payload_0_11_24_imag,
  output     [15:0]   io_coef_out_payload_0_11_25_real,
  output     [15:0]   io_coef_out_payload_0_11_25_imag,
  output     [15:0]   io_coef_out_payload_0_11_26_real,
  output     [15:0]   io_coef_out_payload_0_11_26_imag,
  output     [15:0]   io_coef_out_payload_0_11_27_real,
  output     [15:0]   io_coef_out_payload_0_11_27_imag,
  output     [15:0]   io_coef_out_payload_0_11_28_real,
  output     [15:0]   io_coef_out_payload_0_11_28_imag,
  output     [15:0]   io_coef_out_payload_0_11_29_real,
  output     [15:0]   io_coef_out_payload_0_11_29_imag,
  output     [15:0]   io_coef_out_payload_0_11_30_real,
  output     [15:0]   io_coef_out_payload_0_11_30_imag,
  output     [15:0]   io_coef_out_payload_0_11_31_real,
  output     [15:0]   io_coef_out_payload_0_11_31_imag,
  output     [15:0]   io_coef_out_payload_0_11_32_real,
  output     [15:0]   io_coef_out_payload_0_11_32_imag,
  output     [15:0]   io_coef_out_payload_0_11_33_real,
  output     [15:0]   io_coef_out_payload_0_11_33_imag,
  output     [15:0]   io_coef_out_payload_0_11_34_real,
  output     [15:0]   io_coef_out_payload_0_11_34_imag,
  output     [15:0]   io_coef_out_payload_0_11_35_real,
  output     [15:0]   io_coef_out_payload_0_11_35_imag,
  output     [15:0]   io_coef_out_payload_0_11_36_real,
  output     [15:0]   io_coef_out_payload_0_11_36_imag,
  output     [15:0]   io_coef_out_payload_0_11_37_real,
  output     [15:0]   io_coef_out_payload_0_11_37_imag,
  output     [15:0]   io_coef_out_payload_0_11_38_real,
  output     [15:0]   io_coef_out_payload_0_11_38_imag,
  output     [15:0]   io_coef_out_payload_0_11_39_real,
  output     [15:0]   io_coef_out_payload_0_11_39_imag,
  output     [15:0]   io_coef_out_payload_0_11_40_real,
  output     [15:0]   io_coef_out_payload_0_11_40_imag,
  output     [15:0]   io_coef_out_payload_0_11_41_real,
  output     [15:0]   io_coef_out_payload_0_11_41_imag,
  output     [15:0]   io_coef_out_payload_0_11_42_real,
  output     [15:0]   io_coef_out_payload_0_11_42_imag,
  output     [15:0]   io_coef_out_payload_0_11_43_real,
  output     [15:0]   io_coef_out_payload_0_11_43_imag,
  output     [15:0]   io_coef_out_payload_0_11_44_real,
  output     [15:0]   io_coef_out_payload_0_11_44_imag,
  output     [15:0]   io_coef_out_payload_0_11_45_real,
  output     [15:0]   io_coef_out_payload_0_11_45_imag,
  output     [15:0]   io_coef_out_payload_0_11_46_real,
  output     [15:0]   io_coef_out_payload_0_11_46_imag,
  output     [15:0]   io_coef_out_payload_0_11_47_real,
  output     [15:0]   io_coef_out_payload_0_11_47_imag,
  output     [15:0]   io_coef_out_payload_0_11_48_real,
  output     [15:0]   io_coef_out_payload_0_11_48_imag,
  output     [15:0]   io_coef_out_payload_0_11_49_real,
  output     [15:0]   io_coef_out_payload_0_11_49_imag,
  output     [15:0]   io_coef_out_payload_0_12_0_real,
  output     [15:0]   io_coef_out_payload_0_12_0_imag,
  output     [15:0]   io_coef_out_payload_0_12_1_real,
  output     [15:0]   io_coef_out_payload_0_12_1_imag,
  output     [15:0]   io_coef_out_payload_0_12_2_real,
  output     [15:0]   io_coef_out_payload_0_12_2_imag,
  output     [15:0]   io_coef_out_payload_0_12_3_real,
  output     [15:0]   io_coef_out_payload_0_12_3_imag,
  output     [15:0]   io_coef_out_payload_0_12_4_real,
  output     [15:0]   io_coef_out_payload_0_12_4_imag,
  output     [15:0]   io_coef_out_payload_0_12_5_real,
  output     [15:0]   io_coef_out_payload_0_12_5_imag,
  output     [15:0]   io_coef_out_payload_0_12_6_real,
  output     [15:0]   io_coef_out_payload_0_12_6_imag,
  output     [15:0]   io_coef_out_payload_0_12_7_real,
  output     [15:0]   io_coef_out_payload_0_12_7_imag,
  output     [15:0]   io_coef_out_payload_0_12_8_real,
  output     [15:0]   io_coef_out_payload_0_12_8_imag,
  output     [15:0]   io_coef_out_payload_0_12_9_real,
  output     [15:0]   io_coef_out_payload_0_12_9_imag,
  output     [15:0]   io_coef_out_payload_0_12_10_real,
  output     [15:0]   io_coef_out_payload_0_12_10_imag,
  output     [15:0]   io_coef_out_payload_0_12_11_real,
  output     [15:0]   io_coef_out_payload_0_12_11_imag,
  output     [15:0]   io_coef_out_payload_0_12_12_real,
  output     [15:0]   io_coef_out_payload_0_12_12_imag,
  output     [15:0]   io_coef_out_payload_0_12_13_real,
  output     [15:0]   io_coef_out_payload_0_12_13_imag,
  output     [15:0]   io_coef_out_payload_0_12_14_real,
  output     [15:0]   io_coef_out_payload_0_12_14_imag,
  output     [15:0]   io_coef_out_payload_0_12_15_real,
  output     [15:0]   io_coef_out_payload_0_12_15_imag,
  output     [15:0]   io_coef_out_payload_0_12_16_real,
  output     [15:0]   io_coef_out_payload_0_12_16_imag,
  output     [15:0]   io_coef_out_payload_0_12_17_real,
  output     [15:0]   io_coef_out_payload_0_12_17_imag,
  output     [15:0]   io_coef_out_payload_0_12_18_real,
  output     [15:0]   io_coef_out_payload_0_12_18_imag,
  output     [15:0]   io_coef_out_payload_0_12_19_real,
  output     [15:0]   io_coef_out_payload_0_12_19_imag,
  output     [15:0]   io_coef_out_payload_0_12_20_real,
  output     [15:0]   io_coef_out_payload_0_12_20_imag,
  output     [15:0]   io_coef_out_payload_0_12_21_real,
  output     [15:0]   io_coef_out_payload_0_12_21_imag,
  output     [15:0]   io_coef_out_payload_0_12_22_real,
  output     [15:0]   io_coef_out_payload_0_12_22_imag,
  output     [15:0]   io_coef_out_payload_0_12_23_real,
  output     [15:0]   io_coef_out_payload_0_12_23_imag,
  output     [15:0]   io_coef_out_payload_0_12_24_real,
  output     [15:0]   io_coef_out_payload_0_12_24_imag,
  output     [15:0]   io_coef_out_payload_0_12_25_real,
  output     [15:0]   io_coef_out_payload_0_12_25_imag,
  output     [15:0]   io_coef_out_payload_0_12_26_real,
  output     [15:0]   io_coef_out_payload_0_12_26_imag,
  output     [15:0]   io_coef_out_payload_0_12_27_real,
  output     [15:0]   io_coef_out_payload_0_12_27_imag,
  output     [15:0]   io_coef_out_payload_0_12_28_real,
  output     [15:0]   io_coef_out_payload_0_12_28_imag,
  output     [15:0]   io_coef_out_payload_0_12_29_real,
  output     [15:0]   io_coef_out_payload_0_12_29_imag,
  output     [15:0]   io_coef_out_payload_0_12_30_real,
  output     [15:0]   io_coef_out_payload_0_12_30_imag,
  output     [15:0]   io_coef_out_payload_0_12_31_real,
  output     [15:0]   io_coef_out_payload_0_12_31_imag,
  output     [15:0]   io_coef_out_payload_0_12_32_real,
  output     [15:0]   io_coef_out_payload_0_12_32_imag,
  output     [15:0]   io_coef_out_payload_0_12_33_real,
  output     [15:0]   io_coef_out_payload_0_12_33_imag,
  output     [15:0]   io_coef_out_payload_0_12_34_real,
  output     [15:0]   io_coef_out_payload_0_12_34_imag,
  output     [15:0]   io_coef_out_payload_0_12_35_real,
  output     [15:0]   io_coef_out_payload_0_12_35_imag,
  output     [15:0]   io_coef_out_payload_0_12_36_real,
  output     [15:0]   io_coef_out_payload_0_12_36_imag,
  output     [15:0]   io_coef_out_payload_0_12_37_real,
  output     [15:0]   io_coef_out_payload_0_12_37_imag,
  output     [15:0]   io_coef_out_payload_0_12_38_real,
  output     [15:0]   io_coef_out_payload_0_12_38_imag,
  output     [15:0]   io_coef_out_payload_0_12_39_real,
  output     [15:0]   io_coef_out_payload_0_12_39_imag,
  output     [15:0]   io_coef_out_payload_0_12_40_real,
  output     [15:0]   io_coef_out_payload_0_12_40_imag,
  output     [15:0]   io_coef_out_payload_0_12_41_real,
  output     [15:0]   io_coef_out_payload_0_12_41_imag,
  output     [15:0]   io_coef_out_payload_0_12_42_real,
  output     [15:0]   io_coef_out_payload_0_12_42_imag,
  output     [15:0]   io_coef_out_payload_0_12_43_real,
  output     [15:0]   io_coef_out_payload_0_12_43_imag,
  output     [15:0]   io_coef_out_payload_0_12_44_real,
  output     [15:0]   io_coef_out_payload_0_12_44_imag,
  output     [15:0]   io_coef_out_payload_0_12_45_real,
  output     [15:0]   io_coef_out_payload_0_12_45_imag,
  output     [15:0]   io_coef_out_payload_0_12_46_real,
  output     [15:0]   io_coef_out_payload_0_12_46_imag,
  output     [15:0]   io_coef_out_payload_0_12_47_real,
  output     [15:0]   io_coef_out_payload_0_12_47_imag,
  output     [15:0]   io_coef_out_payload_0_12_48_real,
  output     [15:0]   io_coef_out_payload_0_12_48_imag,
  output     [15:0]   io_coef_out_payload_0_12_49_real,
  output     [15:0]   io_coef_out_payload_0_12_49_imag,
  output     [15:0]   io_coef_out_payload_0_13_0_real,
  output     [15:0]   io_coef_out_payload_0_13_0_imag,
  output     [15:0]   io_coef_out_payload_0_13_1_real,
  output     [15:0]   io_coef_out_payload_0_13_1_imag,
  output     [15:0]   io_coef_out_payload_0_13_2_real,
  output     [15:0]   io_coef_out_payload_0_13_2_imag,
  output     [15:0]   io_coef_out_payload_0_13_3_real,
  output     [15:0]   io_coef_out_payload_0_13_3_imag,
  output     [15:0]   io_coef_out_payload_0_13_4_real,
  output     [15:0]   io_coef_out_payload_0_13_4_imag,
  output     [15:0]   io_coef_out_payload_0_13_5_real,
  output     [15:0]   io_coef_out_payload_0_13_5_imag,
  output     [15:0]   io_coef_out_payload_0_13_6_real,
  output     [15:0]   io_coef_out_payload_0_13_6_imag,
  output     [15:0]   io_coef_out_payload_0_13_7_real,
  output     [15:0]   io_coef_out_payload_0_13_7_imag,
  output     [15:0]   io_coef_out_payload_0_13_8_real,
  output     [15:0]   io_coef_out_payload_0_13_8_imag,
  output     [15:0]   io_coef_out_payload_0_13_9_real,
  output     [15:0]   io_coef_out_payload_0_13_9_imag,
  output     [15:0]   io_coef_out_payload_0_13_10_real,
  output     [15:0]   io_coef_out_payload_0_13_10_imag,
  output     [15:0]   io_coef_out_payload_0_13_11_real,
  output     [15:0]   io_coef_out_payload_0_13_11_imag,
  output     [15:0]   io_coef_out_payload_0_13_12_real,
  output     [15:0]   io_coef_out_payload_0_13_12_imag,
  output     [15:0]   io_coef_out_payload_0_13_13_real,
  output     [15:0]   io_coef_out_payload_0_13_13_imag,
  output     [15:0]   io_coef_out_payload_0_13_14_real,
  output     [15:0]   io_coef_out_payload_0_13_14_imag,
  output     [15:0]   io_coef_out_payload_0_13_15_real,
  output     [15:0]   io_coef_out_payload_0_13_15_imag,
  output     [15:0]   io_coef_out_payload_0_13_16_real,
  output     [15:0]   io_coef_out_payload_0_13_16_imag,
  output     [15:0]   io_coef_out_payload_0_13_17_real,
  output     [15:0]   io_coef_out_payload_0_13_17_imag,
  output     [15:0]   io_coef_out_payload_0_13_18_real,
  output     [15:0]   io_coef_out_payload_0_13_18_imag,
  output     [15:0]   io_coef_out_payload_0_13_19_real,
  output     [15:0]   io_coef_out_payload_0_13_19_imag,
  output     [15:0]   io_coef_out_payload_0_13_20_real,
  output     [15:0]   io_coef_out_payload_0_13_20_imag,
  output     [15:0]   io_coef_out_payload_0_13_21_real,
  output     [15:0]   io_coef_out_payload_0_13_21_imag,
  output     [15:0]   io_coef_out_payload_0_13_22_real,
  output     [15:0]   io_coef_out_payload_0_13_22_imag,
  output     [15:0]   io_coef_out_payload_0_13_23_real,
  output     [15:0]   io_coef_out_payload_0_13_23_imag,
  output     [15:0]   io_coef_out_payload_0_13_24_real,
  output     [15:0]   io_coef_out_payload_0_13_24_imag,
  output     [15:0]   io_coef_out_payload_0_13_25_real,
  output     [15:0]   io_coef_out_payload_0_13_25_imag,
  output     [15:0]   io_coef_out_payload_0_13_26_real,
  output     [15:0]   io_coef_out_payload_0_13_26_imag,
  output     [15:0]   io_coef_out_payload_0_13_27_real,
  output     [15:0]   io_coef_out_payload_0_13_27_imag,
  output     [15:0]   io_coef_out_payload_0_13_28_real,
  output     [15:0]   io_coef_out_payload_0_13_28_imag,
  output     [15:0]   io_coef_out_payload_0_13_29_real,
  output     [15:0]   io_coef_out_payload_0_13_29_imag,
  output     [15:0]   io_coef_out_payload_0_13_30_real,
  output     [15:0]   io_coef_out_payload_0_13_30_imag,
  output     [15:0]   io_coef_out_payload_0_13_31_real,
  output     [15:0]   io_coef_out_payload_0_13_31_imag,
  output     [15:0]   io_coef_out_payload_0_13_32_real,
  output     [15:0]   io_coef_out_payload_0_13_32_imag,
  output     [15:0]   io_coef_out_payload_0_13_33_real,
  output     [15:0]   io_coef_out_payload_0_13_33_imag,
  output     [15:0]   io_coef_out_payload_0_13_34_real,
  output     [15:0]   io_coef_out_payload_0_13_34_imag,
  output     [15:0]   io_coef_out_payload_0_13_35_real,
  output     [15:0]   io_coef_out_payload_0_13_35_imag,
  output     [15:0]   io_coef_out_payload_0_13_36_real,
  output     [15:0]   io_coef_out_payload_0_13_36_imag,
  output     [15:0]   io_coef_out_payload_0_13_37_real,
  output     [15:0]   io_coef_out_payload_0_13_37_imag,
  output     [15:0]   io_coef_out_payload_0_13_38_real,
  output     [15:0]   io_coef_out_payload_0_13_38_imag,
  output     [15:0]   io_coef_out_payload_0_13_39_real,
  output     [15:0]   io_coef_out_payload_0_13_39_imag,
  output     [15:0]   io_coef_out_payload_0_13_40_real,
  output     [15:0]   io_coef_out_payload_0_13_40_imag,
  output     [15:0]   io_coef_out_payload_0_13_41_real,
  output     [15:0]   io_coef_out_payload_0_13_41_imag,
  output     [15:0]   io_coef_out_payload_0_13_42_real,
  output     [15:0]   io_coef_out_payload_0_13_42_imag,
  output     [15:0]   io_coef_out_payload_0_13_43_real,
  output     [15:0]   io_coef_out_payload_0_13_43_imag,
  output     [15:0]   io_coef_out_payload_0_13_44_real,
  output     [15:0]   io_coef_out_payload_0_13_44_imag,
  output     [15:0]   io_coef_out_payload_0_13_45_real,
  output     [15:0]   io_coef_out_payload_0_13_45_imag,
  output     [15:0]   io_coef_out_payload_0_13_46_real,
  output     [15:0]   io_coef_out_payload_0_13_46_imag,
  output     [15:0]   io_coef_out_payload_0_13_47_real,
  output     [15:0]   io_coef_out_payload_0_13_47_imag,
  output     [15:0]   io_coef_out_payload_0_13_48_real,
  output     [15:0]   io_coef_out_payload_0_13_48_imag,
  output     [15:0]   io_coef_out_payload_0_13_49_real,
  output     [15:0]   io_coef_out_payload_0_13_49_imag,
  output     [15:0]   io_coef_out_payload_0_14_0_real,
  output     [15:0]   io_coef_out_payload_0_14_0_imag,
  output     [15:0]   io_coef_out_payload_0_14_1_real,
  output     [15:0]   io_coef_out_payload_0_14_1_imag,
  output     [15:0]   io_coef_out_payload_0_14_2_real,
  output     [15:0]   io_coef_out_payload_0_14_2_imag,
  output     [15:0]   io_coef_out_payload_0_14_3_real,
  output     [15:0]   io_coef_out_payload_0_14_3_imag,
  output     [15:0]   io_coef_out_payload_0_14_4_real,
  output     [15:0]   io_coef_out_payload_0_14_4_imag,
  output     [15:0]   io_coef_out_payload_0_14_5_real,
  output     [15:0]   io_coef_out_payload_0_14_5_imag,
  output     [15:0]   io_coef_out_payload_0_14_6_real,
  output     [15:0]   io_coef_out_payload_0_14_6_imag,
  output     [15:0]   io_coef_out_payload_0_14_7_real,
  output     [15:0]   io_coef_out_payload_0_14_7_imag,
  output     [15:0]   io_coef_out_payload_0_14_8_real,
  output     [15:0]   io_coef_out_payload_0_14_8_imag,
  output     [15:0]   io_coef_out_payload_0_14_9_real,
  output     [15:0]   io_coef_out_payload_0_14_9_imag,
  output     [15:0]   io_coef_out_payload_0_14_10_real,
  output     [15:0]   io_coef_out_payload_0_14_10_imag,
  output     [15:0]   io_coef_out_payload_0_14_11_real,
  output     [15:0]   io_coef_out_payload_0_14_11_imag,
  output     [15:0]   io_coef_out_payload_0_14_12_real,
  output     [15:0]   io_coef_out_payload_0_14_12_imag,
  output     [15:0]   io_coef_out_payload_0_14_13_real,
  output     [15:0]   io_coef_out_payload_0_14_13_imag,
  output     [15:0]   io_coef_out_payload_0_14_14_real,
  output     [15:0]   io_coef_out_payload_0_14_14_imag,
  output     [15:0]   io_coef_out_payload_0_14_15_real,
  output     [15:0]   io_coef_out_payload_0_14_15_imag,
  output     [15:0]   io_coef_out_payload_0_14_16_real,
  output     [15:0]   io_coef_out_payload_0_14_16_imag,
  output     [15:0]   io_coef_out_payload_0_14_17_real,
  output     [15:0]   io_coef_out_payload_0_14_17_imag,
  output     [15:0]   io_coef_out_payload_0_14_18_real,
  output     [15:0]   io_coef_out_payload_0_14_18_imag,
  output     [15:0]   io_coef_out_payload_0_14_19_real,
  output     [15:0]   io_coef_out_payload_0_14_19_imag,
  output     [15:0]   io_coef_out_payload_0_14_20_real,
  output     [15:0]   io_coef_out_payload_0_14_20_imag,
  output     [15:0]   io_coef_out_payload_0_14_21_real,
  output     [15:0]   io_coef_out_payload_0_14_21_imag,
  output     [15:0]   io_coef_out_payload_0_14_22_real,
  output     [15:0]   io_coef_out_payload_0_14_22_imag,
  output     [15:0]   io_coef_out_payload_0_14_23_real,
  output     [15:0]   io_coef_out_payload_0_14_23_imag,
  output     [15:0]   io_coef_out_payload_0_14_24_real,
  output     [15:0]   io_coef_out_payload_0_14_24_imag,
  output     [15:0]   io_coef_out_payload_0_14_25_real,
  output     [15:0]   io_coef_out_payload_0_14_25_imag,
  output     [15:0]   io_coef_out_payload_0_14_26_real,
  output     [15:0]   io_coef_out_payload_0_14_26_imag,
  output     [15:0]   io_coef_out_payload_0_14_27_real,
  output     [15:0]   io_coef_out_payload_0_14_27_imag,
  output     [15:0]   io_coef_out_payload_0_14_28_real,
  output     [15:0]   io_coef_out_payload_0_14_28_imag,
  output     [15:0]   io_coef_out_payload_0_14_29_real,
  output     [15:0]   io_coef_out_payload_0_14_29_imag,
  output     [15:0]   io_coef_out_payload_0_14_30_real,
  output     [15:0]   io_coef_out_payload_0_14_30_imag,
  output     [15:0]   io_coef_out_payload_0_14_31_real,
  output     [15:0]   io_coef_out_payload_0_14_31_imag,
  output     [15:0]   io_coef_out_payload_0_14_32_real,
  output     [15:0]   io_coef_out_payload_0_14_32_imag,
  output     [15:0]   io_coef_out_payload_0_14_33_real,
  output     [15:0]   io_coef_out_payload_0_14_33_imag,
  output     [15:0]   io_coef_out_payload_0_14_34_real,
  output     [15:0]   io_coef_out_payload_0_14_34_imag,
  output     [15:0]   io_coef_out_payload_0_14_35_real,
  output     [15:0]   io_coef_out_payload_0_14_35_imag,
  output     [15:0]   io_coef_out_payload_0_14_36_real,
  output     [15:0]   io_coef_out_payload_0_14_36_imag,
  output     [15:0]   io_coef_out_payload_0_14_37_real,
  output     [15:0]   io_coef_out_payload_0_14_37_imag,
  output     [15:0]   io_coef_out_payload_0_14_38_real,
  output     [15:0]   io_coef_out_payload_0_14_38_imag,
  output     [15:0]   io_coef_out_payload_0_14_39_real,
  output     [15:0]   io_coef_out_payload_0_14_39_imag,
  output     [15:0]   io_coef_out_payload_0_14_40_real,
  output     [15:0]   io_coef_out_payload_0_14_40_imag,
  output     [15:0]   io_coef_out_payload_0_14_41_real,
  output     [15:0]   io_coef_out_payload_0_14_41_imag,
  output     [15:0]   io_coef_out_payload_0_14_42_real,
  output     [15:0]   io_coef_out_payload_0_14_42_imag,
  output     [15:0]   io_coef_out_payload_0_14_43_real,
  output     [15:0]   io_coef_out_payload_0_14_43_imag,
  output     [15:0]   io_coef_out_payload_0_14_44_real,
  output     [15:0]   io_coef_out_payload_0_14_44_imag,
  output     [15:0]   io_coef_out_payload_0_14_45_real,
  output     [15:0]   io_coef_out_payload_0_14_45_imag,
  output     [15:0]   io_coef_out_payload_0_14_46_real,
  output     [15:0]   io_coef_out_payload_0_14_46_imag,
  output     [15:0]   io_coef_out_payload_0_14_47_real,
  output     [15:0]   io_coef_out_payload_0_14_47_imag,
  output     [15:0]   io_coef_out_payload_0_14_48_real,
  output     [15:0]   io_coef_out_payload_0_14_48_imag,
  output     [15:0]   io_coef_out_payload_0_14_49_real,
  output     [15:0]   io_coef_out_payload_0_14_49_imag,
  output     [15:0]   io_coef_out_payload_0_15_0_real,
  output     [15:0]   io_coef_out_payload_0_15_0_imag,
  output     [15:0]   io_coef_out_payload_0_15_1_real,
  output     [15:0]   io_coef_out_payload_0_15_1_imag,
  output     [15:0]   io_coef_out_payload_0_15_2_real,
  output     [15:0]   io_coef_out_payload_0_15_2_imag,
  output     [15:0]   io_coef_out_payload_0_15_3_real,
  output     [15:0]   io_coef_out_payload_0_15_3_imag,
  output     [15:0]   io_coef_out_payload_0_15_4_real,
  output     [15:0]   io_coef_out_payload_0_15_4_imag,
  output     [15:0]   io_coef_out_payload_0_15_5_real,
  output     [15:0]   io_coef_out_payload_0_15_5_imag,
  output     [15:0]   io_coef_out_payload_0_15_6_real,
  output     [15:0]   io_coef_out_payload_0_15_6_imag,
  output     [15:0]   io_coef_out_payload_0_15_7_real,
  output     [15:0]   io_coef_out_payload_0_15_7_imag,
  output     [15:0]   io_coef_out_payload_0_15_8_real,
  output     [15:0]   io_coef_out_payload_0_15_8_imag,
  output     [15:0]   io_coef_out_payload_0_15_9_real,
  output     [15:0]   io_coef_out_payload_0_15_9_imag,
  output     [15:0]   io_coef_out_payload_0_15_10_real,
  output     [15:0]   io_coef_out_payload_0_15_10_imag,
  output     [15:0]   io_coef_out_payload_0_15_11_real,
  output     [15:0]   io_coef_out_payload_0_15_11_imag,
  output     [15:0]   io_coef_out_payload_0_15_12_real,
  output     [15:0]   io_coef_out_payload_0_15_12_imag,
  output     [15:0]   io_coef_out_payload_0_15_13_real,
  output     [15:0]   io_coef_out_payload_0_15_13_imag,
  output     [15:0]   io_coef_out_payload_0_15_14_real,
  output     [15:0]   io_coef_out_payload_0_15_14_imag,
  output     [15:0]   io_coef_out_payload_0_15_15_real,
  output     [15:0]   io_coef_out_payload_0_15_15_imag,
  output     [15:0]   io_coef_out_payload_0_15_16_real,
  output     [15:0]   io_coef_out_payload_0_15_16_imag,
  output     [15:0]   io_coef_out_payload_0_15_17_real,
  output     [15:0]   io_coef_out_payload_0_15_17_imag,
  output     [15:0]   io_coef_out_payload_0_15_18_real,
  output     [15:0]   io_coef_out_payload_0_15_18_imag,
  output     [15:0]   io_coef_out_payload_0_15_19_real,
  output     [15:0]   io_coef_out_payload_0_15_19_imag,
  output     [15:0]   io_coef_out_payload_0_15_20_real,
  output     [15:0]   io_coef_out_payload_0_15_20_imag,
  output     [15:0]   io_coef_out_payload_0_15_21_real,
  output     [15:0]   io_coef_out_payload_0_15_21_imag,
  output     [15:0]   io_coef_out_payload_0_15_22_real,
  output     [15:0]   io_coef_out_payload_0_15_22_imag,
  output     [15:0]   io_coef_out_payload_0_15_23_real,
  output     [15:0]   io_coef_out_payload_0_15_23_imag,
  output     [15:0]   io_coef_out_payload_0_15_24_real,
  output     [15:0]   io_coef_out_payload_0_15_24_imag,
  output     [15:0]   io_coef_out_payload_0_15_25_real,
  output     [15:0]   io_coef_out_payload_0_15_25_imag,
  output     [15:0]   io_coef_out_payload_0_15_26_real,
  output     [15:0]   io_coef_out_payload_0_15_26_imag,
  output     [15:0]   io_coef_out_payload_0_15_27_real,
  output     [15:0]   io_coef_out_payload_0_15_27_imag,
  output     [15:0]   io_coef_out_payload_0_15_28_real,
  output     [15:0]   io_coef_out_payload_0_15_28_imag,
  output     [15:0]   io_coef_out_payload_0_15_29_real,
  output     [15:0]   io_coef_out_payload_0_15_29_imag,
  output     [15:0]   io_coef_out_payload_0_15_30_real,
  output     [15:0]   io_coef_out_payload_0_15_30_imag,
  output     [15:0]   io_coef_out_payload_0_15_31_real,
  output     [15:0]   io_coef_out_payload_0_15_31_imag,
  output     [15:0]   io_coef_out_payload_0_15_32_real,
  output     [15:0]   io_coef_out_payload_0_15_32_imag,
  output     [15:0]   io_coef_out_payload_0_15_33_real,
  output     [15:0]   io_coef_out_payload_0_15_33_imag,
  output     [15:0]   io_coef_out_payload_0_15_34_real,
  output     [15:0]   io_coef_out_payload_0_15_34_imag,
  output     [15:0]   io_coef_out_payload_0_15_35_real,
  output     [15:0]   io_coef_out_payload_0_15_35_imag,
  output     [15:0]   io_coef_out_payload_0_15_36_real,
  output     [15:0]   io_coef_out_payload_0_15_36_imag,
  output     [15:0]   io_coef_out_payload_0_15_37_real,
  output     [15:0]   io_coef_out_payload_0_15_37_imag,
  output     [15:0]   io_coef_out_payload_0_15_38_real,
  output     [15:0]   io_coef_out_payload_0_15_38_imag,
  output     [15:0]   io_coef_out_payload_0_15_39_real,
  output     [15:0]   io_coef_out_payload_0_15_39_imag,
  output     [15:0]   io_coef_out_payload_0_15_40_real,
  output     [15:0]   io_coef_out_payload_0_15_40_imag,
  output     [15:0]   io_coef_out_payload_0_15_41_real,
  output     [15:0]   io_coef_out_payload_0_15_41_imag,
  output     [15:0]   io_coef_out_payload_0_15_42_real,
  output     [15:0]   io_coef_out_payload_0_15_42_imag,
  output     [15:0]   io_coef_out_payload_0_15_43_real,
  output     [15:0]   io_coef_out_payload_0_15_43_imag,
  output     [15:0]   io_coef_out_payload_0_15_44_real,
  output     [15:0]   io_coef_out_payload_0_15_44_imag,
  output     [15:0]   io_coef_out_payload_0_15_45_real,
  output     [15:0]   io_coef_out_payload_0_15_45_imag,
  output     [15:0]   io_coef_out_payload_0_15_46_real,
  output     [15:0]   io_coef_out_payload_0_15_46_imag,
  output     [15:0]   io_coef_out_payload_0_15_47_real,
  output     [15:0]   io_coef_out_payload_0_15_47_imag,
  output     [15:0]   io_coef_out_payload_0_15_48_real,
  output     [15:0]   io_coef_out_payload_0_15_48_imag,
  output     [15:0]   io_coef_out_payload_0_15_49_real,
  output     [15:0]   io_coef_out_payload_0_15_49_imag,
  output     [15:0]   io_coef_out_payload_0_16_0_real,
  output     [15:0]   io_coef_out_payload_0_16_0_imag,
  output     [15:0]   io_coef_out_payload_0_16_1_real,
  output     [15:0]   io_coef_out_payload_0_16_1_imag,
  output     [15:0]   io_coef_out_payload_0_16_2_real,
  output     [15:0]   io_coef_out_payload_0_16_2_imag,
  output     [15:0]   io_coef_out_payload_0_16_3_real,
  output     [15:0]   io_coef_out_payload_0_16_3_imag,
  output     [15:0]   io_coef_out_payload_0_16_4_real,
  output     [15:0]   io_coef_out_payload_0_16_4_imag,
  output     [15:0]   io_coef_out_payload_0_16_5_real,
  output     [15:0]   io_coef_out_payload_0_16_5_imag,
  output     [15:0]   io_coef_out_payload_0_16_6_real,
  output     [15:0]   io_coef_out_payload_0_16_6_imag,
  output     [15:0]   io_coef_out_payload_0_16_7_real,
  output     [15:0]   io_coef_out_payload_0_16_7_imag,
  output     [15:0]   io_coef_out_payload_0_16_8_real,
  output     [15:0]   io_coef_out_payload_0_16_8_imag,
  output     [15:0]   io_coef_out_payload_0_16_9_real,
  output     [15:0]   io_coef_out_payload_0_16_9_imag,
  output     [15:0]   io_coef_out_payload_0_16_10_real,
  output     [15:0]   io_coef_out_payload_0_16_10_imag,
  output     [15:0]   io_coef_out_payload_0_16_11_real,
  output     [15:0]   io_coef_out_payload_0_16_11_imag,
  output     [15:0]   io_coef_out_payload_0_16_12_real,
  output     [15:0]   io_coef_out_payload_0_16_12_imag,
  output     [15:0]   io_coef_out_payload_0_16_13_real,
  output     [15:0]   io_coef_out_payload_0_16_13_imag,
  output     [15:0]   io_coef_out_payload_0_16_14_real,
  output     [15:0]   io_coef_out_payload_0_16_14_imag,
  output     [15:0]   io_coef_out_payload_0_16_15_real,
  output     [15:0]   io_coef_out_payload_0_16_15_imag,
  output     [15:0]   io_coef_out_payload_0_16_16_real,
  output     [15:0]   io_coef_out_payload_0_16_16_imag,
  output     [15:0]   io_coef_out_payload_0_16_17_real,
  output     [15:0]   io_coef_out_payload_0_16_17_imag,
  output     [15:0]   io_coef_out_payload_0_16_18_real,
  output     [15:0]   io_coef_out_payload_0_16_18_imag,
  output     [15:0]   io_coef_out_payload_0_16_19_real,
  output     [15:0]   io_coef_out_payload_0_16_19_imag,
  output     [15:0]   io_coef_out_payload_0_16_20_real,
  output     [15:0]   io_coef_out_payload_0_16_20_imag,
  output     [15:0]   io_coef_out_payload_0_16_21_real,
  output     [15:0]   io_coef_out_payload_0_16_21_imag,
  output     [15:0]   io_coef_out_payload_0_16_22_real,
  output     [15:0]   io_coef_out_payload_0_16_22_imag,
  output     [15:0]   io_coef_out_payload_0_16_23_real,
  output     [15:0]   io_coef_out_payload_0_16_23_imag,
  output     [15:0]   io_coef_out_payload_0_16_24_real,
  output     [15:0]   io_coef_out_payload_0_16_24_imag,
  output     [15:0]   io_coef_out_payload_0_16_25_real,
  output     [15:0]   io_coef_out_payload_0_16_25_imag,
  output     [15:0]   io_coef_out_payload_0_16_26_real,
  output     [15:0]   io_coef_out_payload_0_16_26_imag,
  output     [15:0]   io_coef_out_payload_0_16_27_real,
  output     [15:0]   io_coef_out_payload_0_16_27_imag,
  output     [15:0]   io_coef_out_payload_0_16_28_real,
  output     [15:0]   io_coef_out_payload_0_16_28_imag,
  output     [15:0]   io_coef_out_payload_0_16_29_real,
  output     [15:0]   io_coef_out_payload_0_16_29_imag,
  output     [15:0]   io_coef_out_payload_0_16_30_real,
  output     [15:0]   io_coef_out_payload_0_16_30_imag,
  output     [15:0]   io_coef_out_payload_0_16_31_real,
  output     [15:0]   io_coef_out_payload_0_16_31_imag,
  output     [15:0]   io_coef_out_payload_0_16_32_real,
  output     [15:0]   io_coef_out_payload_0_16_32_imag,
  output     [15:0]   io_coef_out_payload_0_16_33_real,
  output     [15:0]   io_coef_out_payload_0_16_33_imag,
  output     [15:0]   io_coef_out_payload_0_16_34_real,
  output     [15:0]   io_coef_out_payload_0_16_34_imag,
  output     [15:0]   io_coef_out_payload_0_16_35_real,
  output     [15:0]   io_coef_out_payload_0_16_35_imag,
  output     [15:0]   io_coef_out_payload_0_16_36_real,
  output     [15:0]   io_coef_out_payload_0_16_36_imag,
  output     [15:0]   io_coef_out_payload_0_16_37_real,
  output     [15:0]   io_coef_out_payload_0_16_37_imag,
  output     [15:0]   io_coef_out_payload_0_16_38_real,
  output     [15:0]   io_coef_out_payload_0_16_38_imag,
  output     [15:0]   io_coef_out_payload_0_16_39_real,
  output     [15:0]   io_coef_out_payload_0_16_39_imag,
  output     [15:0]   io_coef_out_payload_0_16_40_real,
  output     [15:0]   io_coef_out_payload_0_16_40_imag,
  output     [15:0]   io_coef_out_payload_0_16_41_real,
  output     [15:0]   io_coef_out_payload_0_16_41_imag,
  output     [15:0]   io_coef_out_payload_0_16_42_real,
  output     [15:0]   io_coef_out_payload_0_16_42_imag,
  output     [15:0]   io_coef_out_payload_0_16_43_real,
  output     [15:0]   io_coef_out_payload_0_16_43_imag,
  output     [15:0]   io_coef_out_payload_0_16_44_real,
  output     [15:0]   io_coef_out_payload_0_16_44_imag,
  output     [15:0]   io_coef_out_payload_0_16_45_real,
  output     [15:0]   io_coef_out_payload_0_16_45_imag,
  output     [15:0]   io_coef_out_payload_0_16_46_real,
  output     [15:0]   io_coef_out_payload_0_16_46_imag,
  output     [15:0]   io_coef_out_payload_0_16_47_real,
  output     [15:0]   io_coef_out_payload_0_16_47_imag,
  output     [15:0]   io_coef_out_payload_0_16_48_real,
  output     [15:0]   io_coef_out_payload_0_16_48_imag,
  output     [15:0]   io_coef_out_payload_0_16_49_real,
  output     [15:0]   io_coef_out_payload_0_16_49_imag,
  output     [15:0]   io_coef_out_payload_0_17_0_real,
  output     [15:0]   io_coef_out_payload_0_17_0_imag,
  output     [15:0]   io_coef_out_payload_0_17_1_real,
  output     [15:0]   io_coef_out_payload_0_17_1_imag,
  output     [15:0]   io_coef_out_payload_0_17_2_real,
  output     [15:0]   io_coef_out_payload_0_17_2_imag,
  output     [15:0]   io_coef_out_payload_0_17_3_real,
  output     [15:0]   io_coef_out_payload_0_17_3_imag,
  output     [15:0]   io_coef_out_payload_0_17_4_real,
  output     [15:0]   io_coef_out_payload_0_17_4_imag,
  output     [15:0]   io_coef_out_payload_0_17_5_real,
  output     [15:0]   io_coef_out_payload_0_17_5_imag,
  output     [15:0]   io_coef_out_payload_0_17_6_real,
  output     [15:0]   io_coef_out_payload_0_17_6_imag,
  output     [15:0]   io_coef_out_payload_0_17_7_real,
  output     [15:0]   io_coef_out_payload_0_17_7_imag,
  output     [15:0]   io_coef_out_payload_0_17_8_real,
  output     [15:0]   io_coef_out_payload_0_17_8_imag,
  output     [15:0]   io_coef_out_payload_0_17_9_real,
  output     [15:0]   io_coef_out_payload_0_17_9_imag,
  output     [15:0]   io_coef_out_payload_0_17_10_real,
  output     [15:0]   io_coef_out_payload_0_17_10_imag,
  output     [15:0]   io_coef_out_payload_0_17_11_real,
  output     [15:0]   io_coef_out_payload_0_17_11_imag,
  output     [15:0]   io_coef_out_payload_0_17_12_real,
  output     [15:0]   io_coef_out_payload_0_17_12_imag,
  output     [15:0]   io_coef_out_payload_0_17_13_real,
  output     [15:0]   io_coef_out_payload_0_17_13_imag,
  output     [15:0]   io_coef_out_payload_0_17_14_real,
  output     [15:0]   io_coef_out_payload_0_17_14_imag,
  output     [15:0]   io_coef_out_payload_0_17_15_real,
  output     [15:0]   io_coef_out_payload_0_17_15_imag,
  output     [15:0]   io_coef_out_payload_0_17_16_real,
  output     [15:0]   io_coef_out_payload_0_17_16_imag,
  output     [15:0]   io_coef_out_payload_0_17_17_real,
  output     [15:0]   io_coef_out_payload_0_17_17_imag,
  output     [15:0]   io_coef_out_payload_0_17_18_real,
  output     [15:0]   io_coef_out_payload_0_17_18_imag,
  output     [15:0]   io_coef_out_payload_0_17_19_real,
  output     [15:0]   io_coef_out_payload_0_17_19_imag,
  output     [15:0]   io_coef_out_payload_0_17_20_real,
  output     [15:0]   io_coef_out_payload_0_17_20_imag,
  output     [15:0]   io_coef_out_payload_0_17_21_real,
  output     [15:0]   io_coef_out_payload_0_17_21_imag,
  output     [15:0]   io_coef_out_payload_0_17_22_real,
  output     [15:0]   io_coef_out_payload_0_17_22_imag,
  output     [15:0]   io_coef_out_payload_0_17_23_real,
  output     [15:0]   io_coef_out_payload_0_17_23_imag,
  output     [15:0]   io_coef_out_payload_0_17_24_real,
  output     [15:0]   io_coef_out_payload_0_17_24_imag,
  output     [15:0]   io_coef_out_payload_0_17_25_real,
  output     [15:0]   io_coef_out_payload_0_17_25_imag,
  output     [15:0]   io_coef_out_payload_0_17_26_real,
  output     [15:0]   io_coef_out_payload_0_17_26_imag,
  output     [15:0]   io_coef_out_payload_0_17_27_real,
  output     [15:0]   io_coef_out_payload_0_17_27_imag,
  output     [15:0]   io_coef_out_payload_0_17_28_real,
  output     [15:0]   io_coef_out_payload_0_17_28_imag,
  output     [15:0]   io_coef_out_payload_0_17_29_real,
  output     [15:0]   io_coef_out_payload_0_17_29_imag,
  output     [15:0]   io_coef_out_payload_0_17_30_real,
  output     [15:0]   io_coef_out_payload_0_17_30_imag,
  output     [15:0]   io_coef_out_payload_0_17_31_real,
  output     [15:0]   io_coef_out_payload_0_17_31_imag,
  output     [15:0]   io_coef_out_payload_0_17_32_real,
  output     [15:0]   io_coef_out_payload_0_17_32_imag,
  output     [15:0]   io_coef_out_payload_0_17_33_real,
  output     [15:0]   io_coef_out_payload_0_17_33_imag,
  output     [15:0]   io_coef_out_payload_0_17_34_real,
  output     [15:0]   io_coef_out_payload_0_17_34_imag,
  output     [15:0]   io_coef_out_payload_0_17_35_real,
  output     [15:0]   io_coef_out_payload_0_17_35_imag,
  output     [15:0]   io_coef_out_payload_0_17_36_real,
  output     [15:0]   io_coef_out_payload_0_17_36_imag,
  output     [15:0]   io_coef_out_payload_0_17_37_real,
  output     [15:0]   io_coef_out_payload_0_17_37_imag,
  output     [15:0]   io_coef_out_payload_0_17_38_real,
  output     [15:0]   io_coef_out_payload_0_17_38_imag,
  output     [15:0]   io_coef_out_payload_0_17_39_real,
  output     [15:0]   io_coef_out_payload_0_17_39_imag,
  output     [15:0]   io_coef_out_payload_0_17_40_real,
  output     [15:0]   io_coef_out_payload_0_17_40_imag,
  output     [15:0]   io_coef_out_payload_0_17_41_real,
  output     [15:0]   io_coef_out_payload_0_17_41_imag,
  output     [15:0]   io_coef_out_payload_0_17_42_real,
  output     [15:0]   io_coef_out_payload_0_17_42_imag,
  output     [15:0]   io_coef_out_payload_0_17_43_real,
  output     [15:0]   io_coef_out_payload_0_17_43_imag,
  output     [15:0]   io_coef_out_payload_0_17_44_real,
  output     [15:0]   io_coef_out_payload_0_17_44_imag,
  output     [15:0]   io_coef_out_payload_0_17_45_real,
  output     [15:0]   io_coef_out_payload_0_17_45_imag,
  output     [15:0]   io_coef_out_payload_0_17_46_real,
  output     [15:0]   io_coef_out_payload_0_17_46_imag,
  output     [15:0]   io_coef_out_payload_0_17_47_real,
  output     [15:0]   io_coef_out_payload_0_17_47_imag,
  output     [15:0]   io_coef_out_payload_0_17_48_real,
  output     [15:0]   io_coef_out_payload_0_17_48_imag,
  output     [15:0]   io_coef_out_payload_0_17_49_real,
  output     [15:0]   io_coef_out_payload_0_17_49_imag,
  output     [15:0]   io_coef_out_payload_0_18_0_real,
  output     [15:0]   io_coef_out_payload_0_18_0_imag,
  output     [15:0]   io_coef_out_payload_0_18_1_real,
  output     [15:0]   io_coef_out_payload_0_18_1_imag,
  output     [15:0]   io_coef_out_payload_0_18_2_real,
  output     [15:0]   io_coef_out_payload_0_18_2_imag,
  output     [15:0]   io_coef_out_payload_0_18_3_real,
  output     [15:0]   io_coef_out_payload_0_18_3_imag,
  output     [15:0]   io_coef_out_payload_0_18_4_real,
  output     [15:0]   io_coef_out_payload_0_18_4_imag,
  output     [15:0]   io_coef_out_payload_0_18_5_real,
  output     [15:0]   io_coef_out_payload_0_18_5_imag,
  output     [15:0]   io_coef_out_payload_0_18_6_real,
  output     [15:0]   io_coef_out_payload_0_18_6_imag,
  output     [15:0]   io_coef_out_payload_0_18_7_real,
  output     [15:0]   io_coef_out_payload_0_18_7_imag,
  output     [15:0]   io_coef_out_payload_0_18_8_real,
  output     [15:0]   io_coef_out_payload_0_18_8_imag,
  output     [15:0]   io_coef_out_payload_0_18_9_real,
  output     [15:0]   io_coef_out_payload_0_18_9_imag,
  output     [15:0]   io_coef_out_payload_0_18_10_real,
  output     [15:0]   io_coef_out_payload_0_18_10_imag,
  output     [15:0]   io_coef_out_payload_0_18_11_real,
  output     [15:0]   io_coef_out_payload_0_18_11_imag,
  output     [15:0]   io_coef_out_payload_0_18_12_real,
  output     [15:0]   io_coef_out_payload_0_18_12_imag,
  output     [15:0]   io_coef_out_payload_0_18_13_real,
  output     [15:0]   io_coef_out_payload_0_18_13_imag,
  output     [15:0]   io_coef_out_payload_0_18_14_real,
  output     [15:0]   io_coef_out_payload_0_18_14_imag,
  output     [15:0]   io_coef_out_payload_0_18_15_real,
  output     [15:0]   io_coef_out_payload_0_18_15_imag,
  output     [15:0]   io_coef_out_payload_0_18_16_real,
  output     [15:0]   io_coef_out_payload_0_18_16_imag,
  output     [15:0]   io_coef_out_payload_0_18_17_real,
  output     [15:0]   io_coef_out_payload_0_18_17_imag,
  output     [15:0]   io_coef_out_payload_0_18_18_real,
  output     [15:0]   io_coef_out_payload_0_18_18_imag,
  output     [15:0]   io_coef_out_payload_0_18_19_real,
  output     [15:0]   io_coef_out_payload_0_18_19_imag,
  output     [15:0]   io_coef_out_payload_0_18_20_real,
  output     [15:0]   io_coef_out_payload_0_18_20_imag,
  output     [15:0]   io_coef_out_payload_0_18_21_real,
  output     [15:0]   io_coef_out_payload_0_18_21_imag,
  output     [15:0]   io_coef_out_payload_0_18_22_real,
  output     [15:0]   io_coef_out_payload_0_18_22_imag,
  output     [15:0]   io_coef_out_payload_0_18_23_real,
  output     [15:0]   io_coef_out_payload_0_18_23_imag,
  output     [15:0]   io_coef_out_payload_0_18_24_real,
  output     [15:0]   io_coef_out_payload_0_18_24_imag,
  output     [15:0]   io_coef_out_payload_0_18_25_real,
  output     [15:0]   io_coef_out_payload_0_18_25_imag,
  output     [15:0]   io_coef_out_payload_0_18_26_real,
  output     [15:0]   io_coef_out_payload_0_18_26_imag,
  output     [15:0]   io_coef_out_payload_0_18_27_real,
  output     [15:0]   io_coef_out_payload_0_18_27_imag,
  output     [15:0]   io_coef_out_payload_0_18_28_real,
  output     [15:0]   io_coef_out_payload_0_18_28_imag,
  output     [15:0]   io_coef_out_payload_0_18_29_real,
  output     [15:0]   io_coef_out_payload_0_18_29_imag,
  output     [15:0]   io_coef_out_payload_0_18_30_real,
  output     [15:0]   io_coef_out_payload_0_18_30_imag,
  output     [15:0]   io_coef_out_payload_0_18_31_real,
  output     [15:0]   io_coef_out_payload_0_18_31_imag,
  output     [15:0]   io_coef_out_payload_0_18_32_real,
  output     [15:0]   io_coef_out_payload_0_18_32_imag,
  output     [15:0]   io_coef_out_payload_0_18_33_real,
  output     [15:0]   io_coef_out_payload_0_18_33_imag,
  output     [15:0]   io_coef_out_payload_0_18_34_real,
  output     [15:0]   io_coef_out_payload_0_18_34_imag,
  output     [15:0]   io_coef_out_payload_0_18_35_real,
  output     [15:0]   io_coef_out_payload_0_18_35_imag,
  output     [15:0]   io_coef_out_payload_0_18_36_real,
  output     [15:0]   io_coef_out_payload_0_18_36_imag,
  output     [15:0]   io_coef_out_payload_0_18_37_real,
  output     [15:0]   io_coef_out_payload_0_18_37_imag,
  output     [15:0]   io_coef_out_payload_0_18_38_real,
  output     [15:0]   io_coef_out_payload_0_18_38_imag,
  output     [15:0]   io_coef_out_payload_0_18_39_real,
  output     [15:0]   io_coef_out_payload_0_18_39_imag,
  output     [15:0]   io_coef_out_payload_0_18_40_real,
  output     [15:0]   io_coef_out_payload_0_18_40_imag,
  output     [15:0]   io_coef_out_payload_0_18_41_real,
  output     [15:0]   io_coef_out_payload_0_18_41_imag,
  output     [15:0]   io_coef_out_payload_0_18_42_real,
  output     [15:0]   io_coef_out_payload_0_18_42_imag,
  output     [15:0]   io_coef_out_payload_0_18_43_real,
  output     [15:0]   io_coef_out_payload_0_18_43_imag,
  output     [15:0]   io_coef_out_payload_0_18_44_real,
  output     [15:0]   io_coef_out_payload_0_18_44_imag,
  output     [15:0]   io_coef_out_payload_0_18_45_real,
  output     [15:0]   io_coef_out_payload_0_18_45_imag,
  output     [15:0]   io_coef_out_payload_0_18_46_real,
  output     [15:0]   io_coef_out_payload_0_18_46_imag,
  output     [15:0]   io_coef_out_payload_0_18_47_real,
  output     [15:0]   io_coef_out_payload_0_18_47_imag,
  output     [15:0]   io_coef_out_payload_0_18_48_real,
  output     [15:0]   io_coef_out_payload_0_18_48_imag,
  output     [15:0]   io_coef_out_payload_0_18_49_real,
  output     [15:0]   io_coef_out_payload_0_18_49_imag,
  output     [15:0]   io_coef_out_payload_0_19_0_real,
  output     [15:0]   io_coef_out_payload_0_19_0_imag,
  output     [15:0]   io_coef_out_payload_0_19_1_real,
  output     [15:0]   io_coef_out_payload_0_19_1_imag,
  output     [15:0]   io_coef_out_payload_0_19_2_real,
  output     [15:0]   io_coef_out_payload_0_19_2_imag,
  output     [15:0]   io_coef_out_payload_0_19_3_real,
  output     [15:0]   io_coef_out_payload_0_19_3_imag,
  output     [15:0]   io_coef_out_payload_0_19_4_real,
  output     [15:0]   io_coef_out_payload_0_19_4_imag,
  output     [15:0]   io_coef_out_payload_0_19_5_real,
  output     [15:0]   io_coef_out_payload_0_19_5_imag,
  output     [15:0]   io_coef_out_payload_0_19_6_real,
  output     [15:0]   io_coef_out_payload_0_19_6_imag,
  output     [15:0]   io_coef_out_payload_0_19_7_real,
  output     [15:0]   io_coef_out_payload_0_19_7_imag,
  output     [15:0]   io_coef_out_payload_0_19_8_real,
  output     [15:0]   io_coef_out_payload_0_19_8_imag,
  output     [15:0]   io_coef_out_payload_0_19_9_real,
  output     [15:0]   io_coef_out_payload_0_19_9_imag,
  output     [15:0]   io_coef_out_payload_0_19_10_real,
  output     [15:0]   io_coef_out_payload_0_19_10_imag,
  output     [15:0]   io_coef_out_payload_0_19_11_real,
  output     [15:0]   io_coef_out_payload_0_19_11_imag,
  output     [15:0]   io_coef_out_payload_0_19_12_real,
  output     [15:0]   io_coef_out_payload_0_19_12_imag,
  output     [15:0]   io_coef_out_payload_0_19_13_real,
  output     [15:0]   io_coef_out_payload_0_19_13_imag,
  output     [15:0]   io_coef_out_payload_0_19_14_real,
  output     [15:0]   io_coef_out_payload_0_19_14_imag,
  output     [15:0]   io_coef_out_payload_0_19_15_real,
  output     [15:0]   io_coef_out_payload_0_19_15_imag,
  output     [15:0]   io_coef_out_payload_0_19_16_real,
  output     [15:0]   io_coef_out_payload_0_19_16_imag,
  output     [15:0]   io_coef_out_payload_0_19_17_real,
  output     [15:0]   io_coef_out_payload_0_19_17_imag,
  output     [15:0]   io_coef_out_payload_0_19_18_real,
  output     [15:0]   io_coef_out_payload_0_19_18_imag,
  output     [15:0]   io_coef_out_payload_0_19_19_real,
  output     [15:0]   io_coef_out_payload_0_19_19_imag,
  output     [15:0]   io_coef_out_payload_0_19_20_real,
  output     [15:0]   io_coef_out_payload_0_19_20_imag,
  output     [15:0]   io_coef_out_payload_0_19_21_real,
  output     [15:0]   io_coef_out_payload_0_19_21_imag,
  output     [15:0]   io_coef_out_payload_0_19_22_real,
  output     [15:0]   io_coef_out_payload_0_19_22_imag,
  output     [15:0]   io_coef_out_payload_0_19_23_real,
  output     [15:0]   io_coef_out_payload_0_19_23_imag,
  output     [15:0]   io_coef_out_payload_0_19_24_real,
  output     [15:0]   io_coef_out_payload_0_19_24_imag,
  output     [15:0]   io_coef_out_payload_0_19_25_real,
  output     [15:0]   io_coef_out_payload_0_19_25_imag,
  output     [15:0]   io_coef_out_payload_0_19_26_real,
  output     [15:0]   io_coef_out_payload_0_19_26_imag,
  output     [15:0]   io_coef_out_payload_0_19_27_real,
  output     [15:0]   io_coef_out_payload_0_19_27_imag,
  output     [15:0]   io_coef_out_payload_0_19_28_real,
  output     [15:0]   io_coef_out_payload_0_19_28_imag,
  output     [15:0]   io_coef_out_payload_0_19_29_real,
  output     [15:0]   io_coef_out_payload_0_19_29_imag,
  output     [15:0]   io_coef_out_payload_0_19_30_real,
  output     [15:0]   io_coef_out_payload_0_19_30_imag,
  output     [15:0]   io_coef_out_payload_0_19_31_real,
  output     [15:0]   io_coef_out_payload_0_19_31_imag,
  output     [15:0]   io_coef_out_payload_0_19_32_real,
  output     [15:0]   io_coef_out_payload_0_19_32_imag,
  output     [15:0]   io_coef_out_payload_0_19_33_real,
  output     [15:0]   io_coef_out_payload_0_19_33_imag,
  output     [15:0]   io_coef_out_payload_0_19_34_real,
  output     [15:0]   io_coef_out_payload_0_19_34_imag,
  output     [15:0]   io_coef_out_payload_0_19_35_real,
  output     [15:0]   io_coef_out_payload_0_19_35_imag,
  output     [15:0]   io_coef_out_payload_0_19_36_real,
  output     [15:0]   io_coef_out_payload_0_19_36_imag,
  output     [15:0]   io_coef_out_payload_0_19_37_real,
  output     [15:0]   io_coef_out_payload_0_19_37_imag,
  output     [15:0]   io_coef_out_payload_0_19_38_real,
  output     [15:0]   io_coef_out_payload_0_19_38_imag,
  output     [15:0]   io_coef_out_payload_0_19_39_real,
  output     [15:0]   io_coef_out_payload_0_19_39_imag,
  output     [15:0]   io_coef_out_payload_0_19_40_real,
  output     [15:0]   io_coef_out_payload_0_19_40_imag,
  output     [15:0]   io_coef_out_payload_0_19_41_real,
  output     [15:0]   io_coef_out_payload_0_19_41_imag,
  output     [15:0]   io_coef_out_payload_0_19_42_real,
  output     [15:0]   io_coef_out_payload_0_19_42_imag,
  output     [15:0]   io_coef_out_payload_0_19_43_real,
  output     [15:0]   io_coef_out_payload_0_19_43_imag,
  output     [15:0]   io_coef_out_payload_0_19_44_real,
  output     [15:0]   io_coef_out_payload_0_19_44_imag,
  output     [15:0]   io_coef_out_payload_0_19_45_real,
  output     [15:0]   io_coef_out_payload_0_19_45_imag,
  output     [15:0]   io_coef_out_payload_0_19_46_real,
  output     [15:0]   io_coef_out_payload_0_19_46_imag,
  output     [15:0]   io_coef_out_payload_0_19_47_real,
  output     [15:0]   io_coef_out_payload_0_19_47_imag,
  output     [15:0]   io_coef_out_payload_0_19_48_real,
  output     [15:0]   io_coef_out_payload_0_19_48_imag,
  output     [15:0]   io_coef_out_payload_0_19_49_real,
  output     [15:0]   io_coef_out_payload_0_19_49_imag,
  output     [15:0]   io_coef_out_payload_0_20_0_real,
  output     [15:0]   io_coef_out_payload_0_20_0_imag,
  output     [15:0]   io_coef_out_payload_0_20_1_real,
  output     [15:0]   io_coef_out_payload_0_20_1_imag,
  output     [15:0]   io_coef_out_payload_0_20_2_real,
  output     [15:0]   io_coef_out_payload_0_20_2_imag,
  output     [15:0]   io_coef_out_payload_0_20_3_real,
  output     [15:0]   io_coef_out_payload_0_20_3_imag,
  output     [15:0]   io_coef_out_payload_0_20_4_real,
  output     [15:0]   io_coef_out_payload_0_20_4_imag,
  output     [15:0]   io_coef_out_payload_0_20_5_real,
  output     [15:0]   io_coef_out_payload_0_20_5_imag,
  output     [15:0]   io_coef_out_payload_0_20_6_real,
  output     [15:0]   io_coef_out_payload_0_20_6_imag,
  output     [15:0]   io_coef_out_payload_0_20_7_real,
  output     [15:0]   io_coef_out_payload_0_20_7_imag,
  output     [15:0]   io_coef_out_payload_0_20_8_real,
  output     [15:0]   io_coef_out_payload_0_20_8_imag,
  output     [15:0]   io_coef_out_payload_0_20_9_real,
  output     [15:0]   io_coef_out_payload_0_20_9_imag,
  output     [15:0]   io_coef_out_payload_0_20_10_real,
  output     [15:0]   io_coef_out_payload_0_20_10_imag,
  output     [15:0]   io_coef_out_payload_0_20_11_real,
  output     [15:0]   io_coef_out_payload_0_20_11_imag,
  output     [15:0]   io_coef_out_payload_0_20_12_real,
  output     [15:0]   io_coef_out_payload_0_20_12_imag,
  output     [15:0]   io_coef_out_payload_0_20_13_real,
  output     [15:0]   io_coef_out_payload_0_20_13_imag,
  output     [15:0]   io_coef_out_payload_0_20_14_real,
  output     [15:0]   io_coef_out_payload_0_20_14_imag,
  output     [15:0]   io_coef_out_payload_0_20_15_real,
  output     [15:0]   io_coef_out_payload_0_20_15_imag,
  output     [15:0]   io_coef_out_payload_0_20_16_real,
  output     [15:0]   io_coef_out_payload_0_20_16_imag,
  output     [15:0]   io_coef_out_payload_0_20_17_real,
  output     [15:0]   io_coef_out_payload_0_20_17_imag,
  output     [15:0]   io_coef_out_payload_0_20_18_real,
  output     [15:0]   io_coef_out_payload_0_20_18_imag,
  output     [15:0]   io_coef_out_payload_0_20_19_real,
  output     [15:0]   io_coef_out_payload_0_20_19_imag,
  output     [15:0]   io_coef_out_payload_0_20_20_real,
  output     [15:0]   io_coef_out_payload_0_20_20_imag,
  output     [15:0]   io_coef_out_payload_0_20_21_real,
  output     [15:0]   io_coef_out_payload_0_20_21_imag,
  output     [15:0]   io_coef_out_payload_0_20_22_real,
  output     [15:0]   io_coef_out_payload_0_20_22_imag,
  output     [15:0]   io_coef_out_payload_0_20_23_real,
  output     [15:0]   io_coef_out_payload_0_20_23_imag,
  output     [15:0]   io_coef_out_payload_0_20_24_real,
  output     [15:0]   io_coef_out_payload_0_20_24_imag,
  output     [15:0]   io_coef_out_payload_0_20_25_real,
  output     [15:0]   io_coef_out_payload_0_20_25_imag,
  output     [15:0]   io_coef_out_payload_0_20_26_real,
  output     [15:0]   io_coef_out_payload_0_20_26_imag,
  output     [15:0]   io_coef_out_payload_0_20_27_real,
  output     [15:0]   io_coef_out_payload_0_20_27_imag,
  output     [15:0]   io_coef_out_payload_0_20_28_real,
  output     [15:0]   io_coef_out_payload_0_20_28_imag,
  output     [15:0]   io_coef_out_payload_0_20_29_real,
  output     [15:0]   io_coef_out_payload_0_20_29_imag,
  output     [15:0]   io_coef_out_payload_0_20_30_real,
  output     [15:0]   io_coef_out_payload_0_20_30_imag,
  output     [15:0]   io_coef_out_payload_0_20_31_real,
  output     [15:0]   io_coef_out_payload_0_20_31_imag,
  output     [15:0]   io_coef_out_payload_0_20_32_real,
  output     [15:0]   io_coef_out_payload_0_20_32_imag,
  output     [15:0]   io_coef_out_payload_0_20_33_real,
  output     [15:0]   io_coef_out_payload_0_20_33_imag,
  output     [15:0]   io_coef_out_payload_0_20_34_real,
  output     [15:0]   io_coef_out_payload_0_20_34_imag,
  output     [15:0]   io_coef_out_payload_0_20_35_real,
  output     [15:0]   io_coef_out_payload_0_20_35_imag,
  output     [15:0]   io_coef_out_payload_0_20_36_real,
  output     [15:0]   io_coef_out_payload_0_20_36_imag,
  output     [15:0]   io_coef_out_payload_0_20_37_real,
  output     [15:0]   io_coef_out_payload_0_20_37_imag,
  output     [15:0]   io_coef_out_payload_0_20_38_real,
  output     [15:0]   io_coef_out_payload_0_20_38_imag,
  output     [15:0]   io_coef_out_payload_0_20_39_real,
  output     [15:0]   io_coef_out_payload_0_20_39_imag,
  output     [15:0]   io_coef_out_payload_0_20_40_real,
  output     [15:0]   io_coef_out_payload_0_20_40_imag,
  output     [15:0]   io_coef_out_payload_0_20_41_real,
  output     [15:0]   io_coef_out_payload_0_20_41_imag,
  output     [15:0]   io_coef_out_payload_0_20_42_real,
  output     [15:0]   io_coef_out_payload_0_20_42_imag,
  output     [15:0]   io_coef_out_payload_0_20_43_real,
  output     [15:0]   io_coef_out_payload_0_20_43_imag,
  output     [15:0]   io_coef_out_payload_0_20_44_real,
  output     [15:0]   io_coef_out_payload_0_20_44_imag,
  output     [15:0]   io_coef_out_payload_0_20_45_real,
  output     [15:0]   io_coef_out_payload_0_20_45_imag,
  output     [15:0]   io_coef_out_payload_0_20_46_real,
  output     [15:0]   io_coef_out_payload_0_20_46_imag,
  output     [15:0]   io_coef_out_payload_0_20_47_real,
  output     [15:0]   io_coef_out_payload_0_20_47_imag,
  output     [15:0]   io_coef_out_payload_0_20_48_real,
  output     [15:0]   io_coef_out_payload_0_20_48_imag,
  output     [15:0]   io_coef_out_payload_0_20_49_real,
  output     [15:0]   io_coef_out_payload_0_20_49_imag,
  output     [15:0]   io_coef_out_payload_0_21_0_real,
  output     [15:0]   io_coef_out_payload_0_21_0_imag,
  output     [15:0]   io_coef_out_payload_0_21_1_real,
  output     [15:0]   io_coef_out_payload_0_21_1_imag,
  output     [15:0]   io_coef_out_payload_0_21_2_real,
  output     [15:0]   io_coef_out_payload_0_21_2_imag,
  output     [15:0]   io_coef_out_payload_0_21_3_real,
  output     [15:0]   io_coef_out_payload_0_21_3_imag,
  output     [15:0]   io_coef_out_payload_0_21_4_real,
  output     [15:0]   io_coef_out_payload_0_21_4_imag,
  output     [15:0]   io_coef_out_payload_0_21_5_real,
  output     [15:0]   io_coef_out_payload_0_21_5_imag,
  output     [15:0]   io_coef_out_payload_0_21_6_real,
  output     [15:0]   io_coef_out_payload_0_21_6_imag,
  output     [15:0]   io_coef_out_payload_0_21_7_real,
  output     [15:0]   io_coef_out_payload_0_21_7_imag,
  output     [15:0]   io_coef_out_payload_0_21_8_real,
  output     [15:0]   io_coef_out_payload_0_21_8_imag,
  output     [15:0]   io_coef_out_payload_0_21_9_real,
  output     [15:0]   io_coef_out_payload_0_21_9_imag,
  output     [15:0]   io_coef_out_payload_0_21_10_real,
  output     [15:0]   io_coef_out_payload_0_21_10_imag,
  output     [15:0]   io_coef_out_payload_0_21_11_real,
  output     [15:0]   io_coef_out_payload_0_21_11_imag,
  output     [15:0]   io_coef_out_payload_0_21_12_real,
  output     [15:0]   io_coef_out_payload_0_21_12_imag,
  output     [15:0]   io_coef_out_payload_0_21_13_real,
  output     [15:0]   io_coef_out_payload_0_21_13_imag,
  output     [15:0]   io_coef_out_payload_0_21_14_real,
  output     [15:0]   io_coef_out_payload_0_21_14_imag,
  output     [15:0]   io_coef_out_payload_0_21_15_real,
  output     [15:0]   io_coef_out_payload_0_21_15_imag,
  output     [15:0]   io_coef_out_payload_0_21_16_real,
  output     [15:0]   io_coef_out_payload_0_21_16_imag,
  output     [15:0]   io_coef_out_payload_0_21_17_real,
  output     [15:0]   io_coef_out_payload_0_21_17_imag,
  output     [15:0]   io_coef_out_payload_0_21_18_real,
  output     [15:0]   io_coef_out_payload_0_21_18_imag,
  output     [15:0]   io_coef_out_payload_0_21_19_real,
  output     [15:0]   io_coef_out_payload_0_21_19_imag,
  output     [15:0]   io_coef_out_payload_0_21_20_real,
  output     [15:0]   io_coef_out_payload_0_21_20_imag,
  output     [15:0]   io_coef_out_payload_0_21_21_real,
  output     [15:0]   io_coef_out_payload_0_21_21_imag,
  output     [15:0]   io_coef_out_payload_0_21_22_real,
  output     [15:0]   io_coef_out_payload_0_21_22_imag,
  output     [15:0]   io_coef_out_payload_0_21_23_real,
  output     [15:0]   io_coef_out_payload_0_21_23_imag,
  output     [15:0]   io_coef_out_payload_0_21_24_real,
  output     [15:0]   io_coef_out_payload_0_21_24_imag,
  output     [15:0]   io_coef_out_payload_0_21_25_real,
  output     [15:0]   io_coef_out_payload_0_21_25_imag,
  output     [15:0]   io_coef_out_payload_0_21_26_real,
  output     [15:0]   io_coef_out_payload_0_21_26_imag,
  output     [15:0]   io_coef_out_payload_0_21_27_real,
  output     [15:0]   io_coef_out_payload_0_21_27_imag,
  output     [15:0]   io_coef_out_payload_0_21_28_real,
  output     [15:0]   io_coef_out_payload_0_21_28_imag,
  output     [15:0]   io_coef_out_payload_0_21_29_real,
  output     [15:0]   io_coef_out_payload_0_21_29_imag,
  output     [15:0]   io_coef_out_payload_0_21_30_real,
  output     [15:0]   io_coef_out_payload_0_21_30_imag,
  output     [15:0]   io_coef_out_payload_0_21_31_real,
  output     [15:0]   io_coef_out_payload_0_21_31_imag,
  output     [15:0]   io_coef_out_payload_0_21_32_real,
  output     [15:0]   io_coef_out_payload_0_21_32_imag,
  output     [15:0]   io_coef_out_payload_0_21_33_real,
  output     [15:0]   io_coef_out_payload_0_21_33_imag,
  output     [15:0]   io_coef_out_payload_0_21_34_real,
  output     [15:0]   io_coef_out_payload_0_21_34_imag,
  output     [15:0]   io_coef_out_payload_0_21_35_real,
  output     [15:0]   io_coef_out_payload_0_21_35_imag,
  output     [15:0]   io_coef_out_payload_0_21_36_real,
  output     [15:0]   io_coef_out_payload_0_21_36_imag,
  output     [15:0]   io_coef_out_payload_0_21_37_real,
  output     [15:0]   io_coef_out_payload_0_21_37_imag,
  output     [15:0]   io_coef_out_payload_0_21_38_real,
  output     [15:0]   io_coef_out_payload_0_21_38_imag,
  output     [15:0]   io_coef_out_payload_0_21_39_real,
  output     [15:0]   io_coef_out_payload_0_21_39_imag,
  output     [15:0]   io_coef_out_payload_0_21_40_real,
  output     [15:0]   io_coef_out_payload_0_21_40_imag,
  output     [15:0]   io_coef_out_payload_0_21_41_real,
  output     [15:0]   io_coef_out_payload_0_21_41_imag,
  output     [15:0]   io_coef_out_payload_0_21_42_real,
  output     [15:0]   io_coef_out_payload_0_21_42_imag,
  output     [15:0]   io_coef_out_payload_0_21_43_real,
  output     [15:0]   io_coef_out_payload_0_21_43_imag,
  output     [15:0]   io_coef_out_payload_0_21_44_real,
  output     [15:0]   io_coef_out_payload_0_21_44_imag,
  output     [15:0]   io_coef_out_payload_0_21_45_real,
  output     [15:0]   io_coef_out_payload_0_21_45_imag,
  output     [15:0]   io_coef_out_payload_0_21_46_real,
  output     [15:0]   io_coef_out_payload_0_21_46_imag,
  output     [15:0]   io_coef_out_payload_0_21_47_real,
  output     [15:0]   io_coef_out_payload_0_21_47_imag,
  output     [15:0]   io_coef_out_payload_0_21_48_real,
  output     [15:0]   io_coef_out_payload_0_21_48_imag,
  output     [15:0]   io_coef_out_payload_0_21_49_real,
  output     [15:0]   io_coef_out_payload_0_21_49_imag,
  output     [15:0]   io_coef_out_payload_0_22_0_real,
  output     [15:0]   io_coef_out_payload_0_22_0_imag,
  output     [15:0]   io_coef_out_payload_0_22_1_real,
  output     [15:0]   io_coef_out_payload_0_22_1_imag,
  output     [15:0]   io_coef_out_payload_0_22_2_real,
  output     [15:0]   io_coef_out_payload_0_22_2_imag,
  output     [15:0]   io_coef_out_payload_0_22_3_real,
  output     [15:0]   io_coef_out_payload_0_22_3_imag,
  output     [15:0]   io_coef_out_payload_0_22_4_real,
  output     [15:0]   io_coef_out_payload_0_22_4_imag,
  output     [15:0]   io_coef_out_payload_0_22_5_real,
  output     [15:0]   io_coef_out_payload_0_22_5_imag,
  output     [15:0]   io_coef_out_payload_0_22_6_real,
  output     [15:0]   io_coef_out_payload_0_22_6_imag,
  output     [15:0]   io_coef_out_payload_0_22_7_real,
  output     [15:0]   io_coef_out_payload_0_22_7_imag,
  output     [15:0]   io_coef_out_payload_0_22_8_real,
  output     [15:0]   io_coef_out_payload_0_22_8_imag,
  output     [15:0]   io_coef_out_payload_0_22_9_real,
  output     [15:0]   io_coef_out_payload_0_22_9_imag,
  output     [15:0]   io_coef_out_payload_0_22_10_real,
  output     [15:0]   io_coef_out_payload_0_22_10_imag,
  output     [15:0]   io_coef_out_payload_0_22_11_real,
  output     [15:0]   io_coef_out_payload_0_22_11_imag,
  output     [15:0]   io_coef_out_payload_0_22_12_real,
  output     [15:0]   io_coef_out_payload_0_22_12_imag,
  output     [15:0]   io_coef_out_payload_0_22_13_real,
  output     [15:0]   io_coef_out_payload_0_22_13_imag,
  output     [15:0]   io_coef_out_payload_0_22_14_real,
  output     [15:0]   io_coef_out_payload_0_22_14_imag,
  output     [15:0]   io_coef_out_payload_0_22_15_real,
  output     [15:0]   io_coef_out_payload_0_22_15_imag,
  output     [15:0]   io_coef_out_payload_0_22_16_real,
  output     [15:0]   io_coef_out_payload_0_22_16_imag,
  output     [15:0]   io_coef_out_payload_0_22_17_real,
  output     [15:0]   io_coef_out_payload_0_22_17_imag,
  output     [15:0]   io_coef_out_payload_0_22_18_real,
  output     [15:0]   io_coef_out_payload_0_22_18_imag,
  output     [15:0]   io_coef_out_payload_0_22_19_real,
  output     [15:0]   io_coef_out_payload_0_22_19_imag,
  output     [15:0]   io_coef_out_payload_0_22_20_real,
  output     [15:0]   io_coef_out_payload_0_22_20_imag,
  output     [15:0]   io_coef_out_payload_0_22_21_real,
  output     [15:0]   io_coef_out_payload_0_22_21_imag,
  output     [15:0]   io_coef_out_payload_0_22_22_real,
  output     [15:0]   io_coef_out_payload_0_22_22_imag,
  output     [15:0]   io_coef_out_payload_0_22_23_real,
  output     [15:0]   io_coef_out_payload_0_22_23_imag,
  output     [15:0]   io_coef_out_payload_0_22_24_real,
  output     [15:0]   io_coef_out_payload_0_22_24_imag,
  output     [15:0]   io_coef_out_payload_0_22_25_real,
  output     [15:0]   io_coef_out_payload_0_22_25_imag,
  output     [15:0]   io_coef_out_payload_0_22_26_real,
  output     [15:0]   io_coef_out_payload_0_22_26_imag,
  output     [15:0]   io_coef_out_payload_0_22_27_real,
  output     [15:0]   io_coef_out_payload_0_22_27_imag,
  output     [15:0]   io_coef_out_payload_0_22_28_real,
  output     [15:0]   io_coef_out_payload_0_22_28_imag,
  output     [15:0]   io_coef_out_payload_0_22_29_real,
  output     [15:0]   io_coef_out_payload_0_22_29_imag,
  output     [15:0]   io_coef_out_payload_0_22_30_real,
  output     [15:0]   io_coef_out_payload_0_22_30_imag,
  output     [15:0]   io_coef_out_payload_0_22_31_real,
  output     [15:0]   io_coef_out_payload_0_22_31_imag,
  output     [15:0]   io_coef_out_payload_0_22_32_real,
  output     [15:0]   io_coef_out_payload_0_22_32_imag,
  output     [15:0]   io_coef_out_payload_0_22_33_real,
  output     [15:0]   io_coef_out_payload_0_22_33_imag,
  output     [15:0]   io_coef_out_payload_0_22_34_real,
  output     [15:0]   io_coef_out_payload_0_22_34_imag,
  output     [15:0]   io_coef_out_payload_0_22_35_real,
  output     [15:0]   io_coef_out_payload_0_22_35_imag,
  output     [15:0]   io_coef_out_payload_0_22_36_real,
  output     [15:0]   io_coef_out_payload_0_22_36_imag,
  output     [15:0]   io_coef_out_payload_0_22_37_real,
  output     [15:0]   io_coef_out_payload_0_22_37_imag,
  output     [15:0]   io_coef_out_payload_0_22_38_real,
  output     [15:0]   io_coef_out_payload_0_22_38_imag,
  output     [15:0]   io_coef_out_payload_0_22_39_real,
  output     [15:0]   io_coef_out_payload_0_22_39_imag,
  output     [15:0]   io_coef_out_payload_0_22_40_real,
  output     [15:0]   io_coef_out_payload_0_22_40_imag,
  output     [15:0]   io_coef_out_payload_0_22_41_real,
  output     [15:0]   io_coef_out_payload_0_22_41_imag,
  output     [15:0]   io_coef_out_payload_0_22_42_real,
  output     [15:0]   io_coef_out_payload_0_22_42_imag,
  output     [15:0]   io_coef_out_payload_0_22_43_real,
  output     [15:0]   io_coef_out_payload_0_22_43_imag,
  output     [15:0]   io_coef_out_payload_0_22_44_real,
  output     [15:0]   io_coef_out_payload_0_22_44_imag,
  output     [15:0]   io_coef_out_payload_0_22_45_real,
  output     [15:0]   io_coef_out_payload_0_22_45_imag,
  output     [15:0]   io_coef_out_payload_0_22_46_real,
  output     [15:0]   io_coef_out_payload_0_22_46_imag,
  output     [15:0]   io_coef_out_payload_0_22_47_real,
  output     [15:0]   io_coef_out_payload_0_22_47_imag,
  output     [15:0]   io_coef_out_payload_0_22_48_real,
  output     [15:0]   io_coef_out_payload_0_22_48_imag,
  output     [15:0]   io_coef_out_payload_0_22_49_real,
  output     [15:0]   io_coef_out_payload_0_22_49_imag,
  output     [15:0]   io_coef_out_payload_0_23_0_real,
  output     [15:0]   io_coef_out_payload_0_23_0_imag,
  output     [15:0]   io_coef_out_payload_0_23_1_real,
  output     [15:0]   io_coef_out_payload_0_23_1_imag,
  output     [15:0]   io_coef_out_payload_0_23_2_real,
  output     [15:0]   io_coef_out_payload_0_23_2_imag,
  output     [15:0]   io_coef_out_payload_0_23_3_real,
  output     [15:0]   io_coef_out_payload_0_23_3_imag,
  output     [15:0]   io_coef_out_payload_0_23_4_real,
  output     [15:0]   io_coef_out_payload_0_23_4_imag,
  output     [15:0]   io_coef_out_payload_0_23_5_real,
  output     [15:0]   io_coef_out_payload_0_23_5_imag,
  output     [15:0]   io_coef_out_payload_0_23_6_real,
  output     [15:0]   io_coef_out_payload_0_23_6_imag,
  output     [15:0]   io_coef_out_payload_0_23_7_real,
  output     [15:0]   io_coef_out_payload_0_23_7_imag,
  output     [15:0]   io_coef_out_payload_0_23_8_real,
  output     [15:0]   io_coef_out_payload_0_23_8_imag,
  output     [15:0]   io_coef_out_payload_0_23_9_real,
  output     [15:0]   io_coef_out_payload_0_23_9_imag,
  output     [15:0]   io_coef_out_payload_0_23_10_real,
  output     [15:0]   io_coef_out_payload_0_23_10_imag,
  output     [15:0]   io_coef_out_payload_0_23_11_real,
  output     [15:0]   io_coef_out_payload_0_23_11_imag,
  output     [15:0]   io_coef_out_payload_0_23_12_real,
  output     [15:0]   io_coef_out_payload_0_23_12_imag,
  output     [15:0]   io_coef_out_payload_0_23_13_real,
  output     [15:0]   io_coef_out_payload_0_23_13_imag,
  output     [15:0]   io_coef_out_payload_0_23_14_real,
  output     [15:0]   io_coef_out_payload_0_23_14_imag,
  output     [15:0]   io_coef_out_payload_0_23_15_real,
  output     [15:0]   io_coef_out_payload_0_23_15_imag,
  output     [15:0]   io_coef_out_payload_0_23_16_real,
  output     [15:0]   io_coef_out_payload_0_23_16_imag,
  output     [15:0]   io_coef_out_payload_0_23_17_real,
  output     [15:0]   io_coef_out_payload_0_23_17_imag,
  output     [15:0]   io_coef_out_payload_0_23_18_real,
  output     [15:0]   io_coef_out_payload_0_23_18_imag,
  output     [15:0]   io_coef_out_payload_0_23_19_real,
  output     [15:0]   io_coef_out_payload_0_23_19_imag,
  output     [15:0]   io_coef_out_payload_0_23_20_real,
  output     [15:0]   io_coef_out_payload_0_23_20_imag,
  output     [15:0]   io_coef_out_payload_0_23_21_real,
  output     [15:0]   io_coef_out_payload_0_23_21_imag,
  output     [15:0]   io_coef_out_payload_0_23_22_real,
  output     [15:0]   io_coef_out_payload_0_23_22_imag,
  output     [15:0]   io_coef_out_payload_0_23_23_real,
  output     [15:0]   io_coef_out_payload_0_23_23_imag,
  output     [15:0]   io_coef_out_payload_0_23_24_real,
  output     [15:0]   io_coef_out_payload_0_23_24_imag,
  output     [15:0]   io_coef_out_payload_0_23_25_real,
  output     [15:0]   io_coef_out_payload_0_23_25_imag,
  output     [15:0]   io_coef_out_payload_0_23_26_real,
  output     [15:0]   io_coef_out_payload_0_23_26_imag,
  output     [15:0]   io_coef_out_payload_0_23_27_real,
  output     [15:0]   io_coef_out_payload_0_23_27_imag,
  output     [15:0]   io_coef_out_payload_0_23_28_real,
  output     [15:0]   io_coef_out_payload_0_23_28_imag,
  output     [15:0]   io_coef_out_payload_0_23_29_real,
  output     [15:0]   io_coef_out_payload_0_23_29_imag,
  output     [15:0]   io_coef_out_payload_0_23_30_real,
  output     [15:0]   io_coef_out_payload_0_23_30_imag,
  output     [15:0]   io_coef_out_payload_0_23_31_real,
  output     [15:0]   io_coef_out_payload_0_23_31_imag,
  output     [15:0]   io_coef_out_payload_0_23_32_real,
  output     [15:0]   io_coef_out_payload_0_23_32_imag,
  output     [15:0]   io_coef_out_payload_0_23_33_real,
  output     [15:0]   io_coef_out_payload_0_23_33_imag,
  output     [15:0]   io_coef_out_payload_0_23_34_real,
  output     [15:0]   io_coef_out_payload_0_23_34_imag,
  output     [15:0]   io_coef_out_payload_0_23_35_real,
  output     [15:0]   io_coef_out_payload_0_23_35_imag,
  output     [15:0]   io_coef_out_payload_0_23_36_real,
  output     [15:0]   io_coef_out_payload_0_23_36_imag,
  output     [15:0]   io_coef_out_payload_0_23_37_real,
  output     [15:0]   io_coef_out_payload_0_23_37_imag,
  output     [15:0]   io_coef_out_payload_0_23_38_real,
  output     [15:0]   io_coef_out_payload_0_23_38_imag,
  output     [15:0]   io_coef_out_payload_0_23_39_real,
  output     [15:0]   io_coef_out_payload_0_23_39_imag,
  output     [15:0]   io_coef_out_payload_0_23_40_real,
  output     [15:0]   io_coef_out_payload_0_23_40_imag,
  output     [15:0]   io_coef_out_payload_0_23_41_real,
  output     [15:0]   io_coef_out_payload_0_23_41_imag,
  output     [15:0]   io_coef_out_payload_0_23_42_real,
  output     [15:0]   io_coef_out_payload_0_23_42_imag,
  output     [15:0]   io_coef_out_payload_0_23_43_real,
  output     [15:0]   io_coef_out_payload_0_23_43_imag,
  output     [15:0]   io_coef_out_payload_0_23_44_real,
  output     [15:0]   io_coef_out_payload_0_23_44_imag,
  output     [15:0]   io_coef_out_payload_0_23_45_real,
  output     [15:0]   io_coef_out_payload_0_23_45_imag,
  output     [15:0]   io_coef_out_payload_0_23_46_real,
  output     [15:0]   io_coef_out_payload_0_23_46_imag,
  output     [15:0]   io_coef_out_payload_0_23_47_real,
  output     [15:0]   io_coef_out_payload_0_23_47_imag,
  output     [15:0]   io_coef_out_payload_0_23_48_real,
  output     [15:0]   io_coef_out_payload_0_23_48_imag,
  output     [15:0]   io_coef_out_payload_0_23_49_real,
  output     [15:0]   io_coef_out_payload_0_23_49_imag,
  output     [15:0]   io_coef_out_payload_0_24_0_real,
  output     [15:0]   io_coef_out_payload_0_24_0_imag,
  output     [15:0]   io_coef_out_payload_0_24_1_real,
  output     [15:0]   io_coef_out_payload_0_24_1_imag,
  output     [15:0]   io_coef_out_payload_0_24_2_real,
  output     [15:0]   io_coef_out_payload_0_24_2_imag,
  output     [15:0]   io_coef_out_payload_0_24_3_real,
  output     [15:0]   io_coef_out_payload_0_24_3_imag,
  output     [15:0]   io_coef_out_payload_0_24_4_real,
  output     [15:0]   io_coef_out_payload_0_24_4_imag,
  output     [15:0]   io_coef_out_payload_0_24_5_real,
  output     [15:0]   io_coef_out_payload_0_24_5_imag,
  output     [15:0]   io_coef_out_payload_0_24_6_real,
  output     [15:0]   io_coef_out_payload_0_24_6_imag,
  output     [15:0]   io_coef_out_payload_0_24_7_real,
  output     [15:0]   io_coef_out_payload_0_24_7_imag,
  output     [15:0]   io_coef_out_payload_0_24_8_real,
  output     [15:0]   io_coef_out_payload_0_24_8_imag,
  output     [15:0]   io_coef_out_payload_0_24_9_real,
  output     [15:0]   io_coef_out_payload_0_24_9_imag,
  output     [15:0]   io_coef_out_payload_0_24_10_real,
  output     [15:0]   io_coef_out_payload_0_24_10_imag,
  output     [15:0]   io_coef_out_payload_0_24_11_real,
  output     [15:0]   io_coef_out_payload_0_24_11_imag,
  output     [15:0]   io_coef_out_payload_0_24_12_real,
  output     [15:0]   io_coef_out_payload_0_24_12_imag,
  output     [15:0]   io_coef_out_payload_0_24_13_real,
  output     [15:0]   io_coef_out_payload_0_24_13_imag,
  output     [15:0]   io_coef_out_payload_0_24_14_real,
  output     [15:0]   io_coef_out_payload_0_24_14_imag,
  output     [15:0]   io_coef_out_payload_0_24_15_real,
  output     [15:0]   io_coef_out_payload_0_24_15_imag,
  output     [15:0]   io_coef_out_payload_0_24_16_real,
  output     [15:0]   io_coef_out_payload_0_24_16_imag,
  output     [15:0]   io_coef_out_payload_0_24_17_real,
  output     [15:0]   io_coef_out_payload_0_24_17_imag,
  output     [15:0]   io_coef_out_payload_0_24_18_real,
  output     [15:0]   io_coef_out_payload_0_24_18_imag,
  output     [15:0]   io_coef_out_payload_0_24_19_real,
  output     [15:0]   io_coef_out_payload_0_24_19_imag,
  output     [15:0]   io_coef_out_payload_0_24_20_real,
  output     [15:0]   io_coef_out_payload_0_24_20_imag,
  output     [15:0]   io_coef_out_payload_0_24_21_real,
  output     [15:0]   io_coef_out_payload_0_24_21_imag,
  output     [15:0]   io_coef_out_payload_0_24_22_real,
  output     [15:0]   io_coef_out_payload_0_24_22_imag,
  output     [15:0]   io_coef_out_payload_0_24_23_real,
  output     [15:0]   io_coef_out_payload_0_24_23_imag,
  output     [15:0]   io_coef_out_payload_0_24_24_real,
  output     [15:0]   io_coef_out_payload_0_24_24_imag,
  output     [15:0]   io_coef_out_payload_0_24_25_real,
  output     [15:0]   io_coef_out_payload_0_24_25_imag,
  output     [15:0]   io_coef_out_payload_0_24_26_real,
  output     [15:0]   io_coef_out_payload_0_24_26_imag,
  output     [15:0]   io_coef_out_payload_0_24_27_real,
  output     [15:0]   io_coef_out_payload_0_24_27_imag,
  output     [15:0]   io_coef_out_payload_0_24_28_real,
  output     [15:0]   io_coef_out_payload_0_24_28_imag,
  output     [15:0]   io_coef_out_payload_0_24_29_real,
  output     [15:0]   io_coef_out_payload_0_24_29_imag,
  output     [15:0]   io_coef_out_payload_0_24_30_real,
  output     [15:0]   io_coef_out_payload_0_24_30_imag,
  output     [15:0]   io_coef_out_payload_0_24_31_real,
  output     [15:0]   io_coef_out_payload_0_24_31_imag,
  output     [15:0]   io_coef_out_payload_0_24_32_real,
  output     [15:0]   io_coef_out_payload_0_24_32_imag,
  output     [15:0]   io_coef_out_payload_0_24_33_real,
  output     [15:0]   io_coef_out_payload_0_24_33_imag,
  output     [15:0]   io_coef_out_payload_0_24_34_real,
  output     [15:0]   io_coef_out_payload_0_24_34_imag,
  output     [15:0]   io_coef_out_payload_0_24_35_real,
  output     [15:0]   io_coef_out_payload_0_24_35_imag,
  output     [15:0]   io_coef_out_payload_0_24_36_real,
  output     [15:0]   io_coef_out_payload_0_24_36_imag,
  output     [15:0]   io_coef_out_payload_0_24_37_real,
  output     [15:0]   io_coef_out_payload_0_24_37_imag,
  output     [15:0]   io_coef_out_payload_0_24_38_real,
  output     [15:0]   io_coef_out_payload_0_24_38_imag,
  output     [15:0]   io_coef_out_payload_0_24_39_real,
  output     [15:0]   io_coef_out_payload_0_24_39_imag,
  output     [15:0]   io_coef_out_payload_0_24_40_real,
  output     [15:0]   io_coef_out_payload_0_24_40_imag,
  output     [15:0]   io_coef_out_payload_0_24_41_real,
  output     [15:0]   io_coef_out_payload_0_24_41_imag,
  output     [15:0]   io_coef_out_payload_0_24_42_real,
  output     [15:0]   io_coef_out_payload_0_24_42_imag,
  output     [15:0]   io_coef_out_payload_0_24_43_real,
  output     [15:0]   io_coef_out_payload_0_24_43_imag,
  output     [15:0]   io_coef_out_payload_0_24_44_real,
  output     [15:0]   io_coef_out_payload_0_24_44_imag,
  output     [15:0]   io_coef_out_payload_0_24_45_real,
  output     [15:0]   io_coef_out_payload_0_24_45_imag,
  output     [15:0]   io_coef_out_payload_0_24_46_real,
  output     [15:0]   io_coef_out_payload_0_24_46_imag,
  output     [15:0]   io_coef_out_payload_0_24_47_real,
  output     [15:0]   io_coef_out_payload_0_24_47_imag,
  output     [15:0]   io_coef_out_payload_0_24_48_real,
  output     [15:0]   io_coef_out_payload_0_24_48_imag,
  output     [15:0]   io_coef_out_payload_0_24_49_real,
  output     [15:0]   io_coef_out_payload_0_24_49_imag,
  output     [15:0]   io_coef_out_payload_0_25_0_real,
  output     [15:0]   io_coef_out_payload_0_25_0_imag,
  output     [15:0]   io_coef_out_payload_0_25_1_real,
  output     [15:0]   io_coef_out_payload_0_25_1_imag,
  output     [15:0]   io_coef_out_payload_0_25_2_real,
  output     [15:0]   io_coef_out_payload_0_25_2_imag,
  output     [15:0]   io_coef_out_payload_0_25_3_real,
  output     [15:0]   io_coef_out_payload_0_25_3_imag,
  output     [15:0]   io_coef_out_payload_0_25_4_real,
  output     [15:0]   io_coef_out_payload_0_25_4_imag,
  output     [15:0]   io_coef_out_payload_0_25_5_real,
  output     [15:0]   io_coef_out_payload_0_25_5_imag,
  output     [15:0]   io_coef_out_payload_0_25_6_real,
  output     [15:0]   io_coef_out_payload_0_25_6_imag,
  output     [15:0]   io_coef_out_payload_0_25_7_real,
  output     [15:0]   io_coef_out_payload_0_25_7_imag,
  output     [15:0]   io_coef_out_payload_0_25_8_real,
  output     [15:0]   io_coef_out_payload_0_25_8_imag,
  output     [15:0]   io_coef_out_payload_0_25_9_real,
  output     [15:0]   io_coef_out_payload_0_25_9_imag,
  output     [15:0]   io_coef_out_payload_0_25_10_real,
  output     [15:0]   io_coef_out_payload_0_25_10_imag,
  output     [15:0]   io_coef_out_payload_0_25_11_real,
  output     [15:0]   io_coef_out_payload_0_25_11_imag,
  output     [15:0]   io_coef_out_payload_0_25_12_real,
  output     [15:0]   io_coef_out_payload_0_25_12_imag,
  output     [15:0]   io_coef_out_payload_0_25_13_real,
  output     [15:0]   io_coef_out_payload_0_25_13_imag,
  output     [15:0]   io_coef_out_payload_0_25_14_real,
  output     [15:0]   io_coef_out_payload_0_25_14_imag,
  output     [15:0]   io_coef_out_payload_0_25_15_real,
  output     [15:0]   io_coef_out_payload_0_25_15_imag,
  output     [15:0]   io_coef_out_payload_0_25_16_real,
  output     [15:0]   io_coef_out_payload_0_25_16_imag,
  output     [15:0]   io_coef_out_payload_0_25_17_real,
  output     [15:0]   io_coef_out_payload_0_25_17_imag,
  output     [15:0]   io_coef_out_payload_0_25_18_real,
  output     [15:0]   io_coef_out_payload_0_25_18_imag,
  output     [15:0]   io_coef_out_payload_0_25_19_real,
  output     [15:0]   io_coef_out_payload_0_25_19_imag,
  output     [15:0]   io_coef_out_payload_0_25_20_real,
  output     [15:0]   io_coef_out_payload_0_25_20_imag,
  output     [15:0]   io_coef_out_payload_0_25_21_real,
  output     [15:0]   io_coef_out_payload_0_25_21_imag,
  output     [15:0]   io_coef_out_payload_0_25_22_real,
  output     [15:0]   io_coef_out_payload_0_25_22_imag,
  output     [15:0]   io_coef_out_payload_0_25_23_real,
  output     [15:0]   io_coef_out_payload_0_25_23_imag,
  output     [15:0]   io_coef_out_payload_0_25_24_real,
  output     [15:0]   io_coef_out_payload_0_25_24_imag,
  output     [15:0]   io_coef_out_payload_0_25_25_real,
  output     [15:0]   io_coef_out_payload_0_25_25_imag,
  output     [15:0]   io_coef_out_payload_0_25_26_real,
  output     [15:0]   io_coef_out_payload_0_25_26_imag,
  output     [15:0]   io_coef_out_payload_0_25_27_real,
  output     [15:0]   io_coef_out_payload_0_25_27_imag,
  output     [15:0]   io_coef_out_payload_0_25_28_real,
  output     [15:0]   io_coef_out_payload_0_25_28_imag,
  output     [15:0]   io_coef_out_payload_0_25_29_real,
  output     [15:0]   io_coef_out_payload_0_25_29_imag,
  output     [15:0]   io_coef_out_payload_0_25_30_real,
  output     [15:0]   io_coef_out_payload_0_25_30_imag,
  output     [15:0]   io_coef_out_payload_0_25_31_real,
  output     [15:0]   io_coef_out_payload_0_25_31_imag,
  output     [15:0]   io_coef_out_payload_0_25_32_real,
  output     [15:0]   io_coef_out_payload_0_25_32_imag,
  output     [15:0]   io_coef_out_payload_0_25_33_real,
  output     [15:0]   io_coef_out_payload_0_25_33_imag,
  output     [15:0]   io_coef_out_payload_0_25_34_real,
  output     [15:0]   io_coef_out_payload_0_25_34_imag,
  output     [15:0]   io_coef_out_payload_0_25_35_real,
  output     [15:0]   io_coef_out_payload_0_25_35_imag,
  output     [15:0]   io_coef_out_payload_0_25_36_real,
  output     [15:0]   io_coef_out_payload_0_25_36_imag,
  output     [15:0]   io_coef_out_payload_0_25_37_real,
  output     [15:0]   io_coef_out_payload_0_25_37_imag,
  output     [15:0]   io_coef_out_payload_0_25_38_real,
  output     [15:0]   io_coef_out_payload_0_25_38_imag,
  output     [15:0]   io_coef_out_payload_0_25_39_real,
  output     [15:0]   io_coef_out_payload_0_25_39_imag,
  output     [15:0]   io_coef_out_payload_0_25_40_real,
  output     [15:0]   io_coef_out_payload_0_25_40_imag,
  output     [15:0]   io_coef_out_payload_0_25_41_real,
  output     [15:0]   io_coef_out_payload_0_25_41_imag,
  output     [15:0]   io_coef_out_payload_0_25_42_real,
  output     [15:0]   io_coef_out_payload_0_25_42_imag,
  output     [15:0]   io_coef_out_payload_0_25_43_real,
  output     [15:0]   io_coef_out_payload_0_25_43_imag,
  output     [15:0]   io_coef_out_payload_0_25_44_real,
  output     [15:0]   io_coef_out_payload_0_25_44_imag,
  output     [15:0]   io_coef_out_payload_0_25_45_real,
  output     [15:0]   io_coef_out_payload_0_25_45_imag,
  output     [15:0]   io_coef_out_payload_0_25_46_real,
  output     [15:0]   io_coef_out_payload_0_25_46_imag,
  output     [15:0]   io_coef_out_payload_0_25_47_real,
  output     [15:0]   io_coef_out_payload_0_25_47_imag,
  output     [15:0]   io_coef_out_payload_0_25_48_real,
  output     [15:0]   io_coef_out_payload_0_25_48_imag,
  output     [15:0]   io_coef_out_payload_0_25_49_real,
  output     [15:0]   io_coef_out_payload_0_25_49_imag,
  output     [15:0]   io_coef_out_payload_0_26_0_real,
  output     [15:0]   io_coef_out_payload_0_26_0_imag,
  output     [15:0]   io_coef_out_payload_0_26_1_real,
  output     [15:0]   io_coef_out_payload_0_26_1_imag,
  output     [15:0]   io_coef_out_payload_0_26_2_real,
  output     [15:0]   io_coef_out_payload_0_26_2_imag,
  output     [15:0]   io_coef_out_payload_0_26_3_real,
  output     [15:0]   io_coef_out_payload_0_26_3_imag,
  output     [15:0]   io_coef_out_payload_0_26_4_real,
  output     [15:0]   io_coef_out_payload_0_26_4_imag,
  output     [15:0]   io_coef_out_payload_0_26_5_real,
  output     [15:0]   io_coef_out_payload_0_26_5_imag,
  output     [15:0]   io_coef_out_payload_0_26_6_real,
  output     [15:0]   io_coef_out_payload_0_26_6_imag,
  output     [15:0]   io_coef_out_payload_0_26_7_real,
  output     [15:0]   io_coef_out_payload_0_26_7_imag,
  output     [15:0]   io_coef_out_payload_0_26_8_real,
  output     [15:0]   io_coef_out_payload_0_26_8_imag,
  output     [15:0]   io_coef_out_payload_0_26_9_real,
  output     [15:0]   io_coef_out_payload_0_26_9_imag,
  output     [15:0]   io_coef_out_payload_0_26_10_real,
  output     [15:0]   io_coef_out_payload_0_26_10_imag,
  output     [15:0]   io_coef_out_payload_0_26_11_real,
  output     [15:0]   io_coef_out_payload_0_26_11_imag,
  output     [15:0]   io_coef_out_payload_0_26_12_real,
  output     [15:0]   io_coef_out_payload_0_26_12_imag,
  output     [15:0]   io_coef_out_payload_0_26_13_real,
  output     [15:0]   io_coef_out_payload_0_26_13_imag,
  output     [15:0]   io_coef_out_payload_0_26_14_real,
  output     [15:0]   io_coef_out_payload_0_26_14_imag,
  output     [15:0]   io_coef_out_payload_0_26_15_real,
  output     [15:0]   io_coef_out_payload_0_26_15_imag,
  output     [15:0]   io_coef_out_payload_0_26_16_real,
  output     [15:0]   io_coef_out_payload_0_26_16_imag,
  output     [15:0]   io_coef_out_payload_0_26_17_real,
  output     [15:0]   io_coef_out_payload_0_26_17_imag,
  output     [15:0]   io_coef_out_payload_0_26_18_real,
  output     [15:0]   io_coef_out_payload_0_26_18_imag,
  output     [15:0]   io_coef_out_payload_0_26_19_real,
  output     [15:0]   io_coef_out_payload_0_26_19_imag,
  output     [15:0]   io_coef_out_payload_0_26_20_real,
  output     [15:0]   io_coef_out_payload_0_26_20_imag,
  output     [15:0]   io_coef_out_payload_0_26_21_real,
  output     [15:0]   io_coef_out_payload_0_26_21_imag,
  output     [15:0]   io_coef_out_payload_0_26_22_real,
  output     [15:0]   io_coef_out_payload_0_26_22_imag,
  output     [15:0]   io_coef_out_payload_0_26_23_real,
  output     [15:0]   io_coef_out_payload_0_26_23_imag,
  output     [15:0]   io_coef_out_payload_0_26_24_real,
  output     [15:0]   io_coef_out_payload_0_26_24_imag,
  output     [15:0]   io_coef_out_payload_0_26_25_real,
  output     [15:0]   io_coef_out_payload_0_26_25_imag,
  output     [15:0]   io_coef_out_payload_0_26_26_real,
  output     [15:0]   io_coef_out_payload_0_26_26_imag,
  output     [15:0]   io_coef_out_payload_0_26_27_real,
  output     [15:0]   io_coef_out_payload_0_26_27_imag,
  output     [15:0]   io_coef_out_payload_0_26_28_real,
  output     [15:0]   io_coef_out_payload_0_26_28_imag,
  output     [15:0]   io_coef_out_payload_0_26_29_real,
  output     [15:0]   io_coef_out_payload_0_26_29_imag,
  output     [15:0]   io_coef_out_payload_0_26_30_real,
  output     [15:0]   io_coef_out_payload_0_26_30_imag,
  output     [15:0]   io_coef_out_payload_0_26_31_real,
  output     [15:0]   io_coef_out_payload_0_26_31_imag,
  output     [15:0]   io_coef_out_payload_0_26_32_real,
  output     [15:0]   io_coef_out_payload_0_26_32_imag,
  output     [15:0]   io_coef_out_payload_0_26_33_real,
  output     [15:0]   io_coef_out_payload_0_26_33_imag,
  output     [15:0]   io_coef_out_payload_0_26_34_real,
  output     [15:0]   io_coef_out_payload_0_26_34_imag,
  output     [15:0]   io_coef_out_payload_0_26_35_real,
  output     [15:0]   io_coef_out_payload_0_26_35_imag,
  output     [15:0]   io_coef_out_payload_0_26_36_real,
  output     [15:0]   io_coef_out_payload_0_26_36_imag,
  output     [15:0]   io_coef_out_payload_0_26_37_real,
  output     [15:0]   io_coef_out_payload_0_26_37_imag,
  output     [15:0]   io_coef_out_payload_0_26_38_real,
  output     [15:0]   io_coef_out_payload_0_26_38_imag,
  output     [15:0]   io_coef_out_payload_0_26_39_real,
  output     [15:0]   io_coef_out_payload_0_26_39_imag,
  output     [15:0]   io_coef_out_payload_0_26_40_real,
  output     [15:0]   io_coef_out_payload_0_26_40_imag,
  output     [15:0]   io_coef_out_payload_0_26_41_real,
  output     [15:0]   io_coef_out_payload_0_26_41_imag,
  output     [15:0]   io_coef_out_payload_0_26_42_real,
  output     [15:0]   io_coef_out_payload_0_26_42_imag,
  output     [15:0]   io_coef_out_payload_0_26_43_real,
  output     [15:0]   io_coef_out_payload_0_26_43_imag,
  output     [15:0]   io_coef_out_payload_0_26_44_real,
  output     [15:0]   io_coef_out_payload_0_26_44_imag,
  output     [15:0]   io_coef_out_payload_0_26_45_real,
  output     [15:0]   io_coef_out_payload_0_26_45_imag,
  output     [15:0]   io_coef_out_payload_0_26_46_real,
  output     [15:0]   io_coef_out_payload_0_26_46_imag,
  output     [15:0]   io_coef_out_payload_0_26_47_real,
  output     [15:0]   io_coef_out_payload_0_26_47_imag,
  output     [15:0]   io_coef_out_payload_0_26_48_real,
  output     [15:0]   io_coef_out_payload_0_26_48_imag,
  output     [15:0]   io_coef_out_payload_0_26_49_real,
  output     [15:0]   io_coef_out_payload_0_26_49_imag,
  output     [15:0]   io_coef_out_payload_0_27_0_real,
  output     [15:0]   io_coef_out_payload_0_27_0_imag,
  output     [15:0]   io_coef_out_payload_0_27_1_real,
  output     [15:0]   io_coef_out_payload_0_27_1_imag,
  output     [15:0]   io_coef_out_payload_0_27_2_real,
  output     [15:0]   io_coef_out_payload_0_27_2_imag,
  output     [15:0]   io_coef_out_payload_0_27_3_real,
  output     [15:0]   io_coef_out_payload_0_27_3_imag,
  output     [15:0]   io_coef_out_payload_0_27_4_real,
  output     [15:0]   io_coef_out_payload_0_27_4_imag,
  output     [15:0]   io_coef_out_payload_0_27_5_real,
  output     [15:0]   io_coef_out_payload_0_27_5_imag,
  output     [15:0]   io_coef_out_payload_0_27_6_real,
  output     [15:0]   io_coef_out_payload_0_27_6_imag,
  output     [15:0]   io_coef_out_payload_0_27_7_real,
  output     [15:0]   io_coef_out_payload_0_27_7_imag,
  output     [15:0]   io_coef_out_payload_0_27_8_real,
  output     [15:0]   io_coef_out_payload_0_27_8_imag,
  output     [15:0]   io_coef_out_payload_0_27_9_real,
  output     [15:0]   io_coef_out_payload_0_27_9_imag,
  output     [15:0]   io_coef_out_payload_0_27_10_real,
  output     [15:0]   io_coef_out_payload_0_27_10_imag,
  output     [15:0]   io_coef_out_payload_0_27_11_real,
  output     [15:0]   io_coef_out_payload_0_27_11_imag,
  output     [15:0]   io_coef_out_payload_0_27_12_real,
  output     [15:0]   io_coef_out_payload_0_27_12_imag,
  output     [15:0]   io_coef_out_payload_0_27_13_real,
  output     [15:0]   io_coef_out_payload_0_27_13_imag,
  output     [15:0]   io_coef_out_payload_0_27_14_real,
  output     [15:0]   io_coef_out_payload_0_27_14_imag,
  output     [15:0]   io_coef_out_payload_0_27_15_real,
  output     [15:0]   io_coef_out_payload_0_27_15_imag,
  output     [15:0]   io_coef_out_payload_0_27_16_real,
  output     [15:0]   io_coef_out_payload_0_27_16_imag,
  output     [15:0]   io_coef_out_payload_0_27_17_real,
  output     [15:0]   io_coef_out_payload_0_27_17_imag,
  output     [15:0]   io_coef_out_payload_0_27_18_real,
  output     [15:0]   io_coef_out_payload_0_27_18_imag,
  output     [15:0]   io_coef_out_payload_0_27_19_real,
  output     [15:0]   io_coef_out_payload_0_27_19_imag,
  output     [15:0]   io_coef_out_payload_0_27_20_real,
  output     [15:0]   io_coef_out_payload_0_27_20_imag,
  output     [15:0]   io_coef_out_payload_0_27_21_real,
  output     [15:0]   io_coef_out_payload_0_27_21_imag,
  output     [15:0]   io_coef_out_payload_0_27_22_real,
  output     [15:0]   io_coef_out_payload_0_27_22_imag,
  output     [15:0]   io_coef_out_payload_0_27_23_real,
  output     [15:0]   io_coef_out_payload_0_27_23_imag,
  output     [15:0]   io_coef_out_payload_0_27_24_real,
  output     [15:0]   io_coef_out_payload_0_27_24_imag,
  output     [15:0]   io_coef_out_payload_0_27_25_real,
  output     [15:0]   io_coef_out_payload_0_27_25_imag,
  output     [15:0]   io_coef_out_payload_0_27_26_real,
  output     [15:0]   io_coef_out_payload_0_27_26_imag,
  output     [15:0]   io_coef_out_payload_0_27_27_real,
  output     [15:0]   io_coef_out_payload_0_27_27_imag,
  output     [15:0]   io_coef_out_payload_0_27_28_real,
  output     [15:0]   io_coef_out_payload_0_27_28_imag,
  output     [15:0]   io_coef_out_payload_0_27_29_real,
  output     [15:0]   io_coef_out_payload_0_27_29_imag,
  output     [15:0]   io_coef_out_payload_0_27_30_real,
  output     [15:0]   io_coef_out_payload_0_27_30_imag,
  output     [15:0]   io_coef_out_payload_0_27_31_real,
  output     [15:0]   io_coef_out_payload_0_27_31_imag,
  output     [15:0]   io_coef_out_payload_0_27_32_real,
  output     [15:0]   io_coef_out_payload_0_27_32_imag,
  output     [15:0]   io_coef_out_payload_0_27_33_real,
  output     [15:0]   io_coef_out_payload_0_27_33_imag,
  output     [15:0]   io_coef_out_payload_0_27_34_real,
  output     [15:0]   io_coef_out_payload_0_27_34_imag,
  output     [15:0]   io_coef_out_payload_0_27_35_real,
  output     [15:0]   io_coef_out_payload_0_27_35_imag,
  output     [15:0]   io_coef_out_payload_0_27_36_real,
  output     [15:0]   io_coef_out_payload_0_27_36_imag,
  output     [15:0]   io_coef_out_payload_0_27_37_real,
  output     [15:0]   io_coef_out_payload_0_27_37_imag,
  output     [15:0]   io_coef_out_payload_0_27_38_real,
  output     [15:0]   io_coef_out_payload_0_27_38_imag,
  output     [15:0]   io_coef_out_payload_0_27_39_real,
  output     [15:0]   io_coef_out_payload_0_27_39_imag,
  output     [15:0]   io_coef_out_payload_0_27_40_real,
  output     [15:0]   io_coef_out_payload_0_27_40_imag,
  output     [15:0]   io_coef_out_payload_0_27_41_real,
  output     [15:0]   io_coef_out_payload_0_27_41_imag,
  output     [15:0]   io_coef_out_payload_0_27_42_real,
  output     [15:0]   io_coef_out_payload_0_27_42_imag,
  output     [15:0]   io_coef_out_payload_0_27_43_real,
  output     [15:0]   io_coef_out_payload_0_27_43_imag,
  output     [15:0]   io_coef_out_payload_0_27_44_real,
  output     [15:0]   io_coef_out_payload_0_27_44_imag,
  output     [15:0]   io_coef_out_payload_0_27_45_real,
  output     [15:0]   io_coef_out_payload_0_27_45_imag,
  output     [15:0]   io_coef_out_payload_0_27_46_real,
  output     [15:0]   io_coef_out_payload_0_27_46_imag,
  output     [15:0]   io_coef_out_payload_0_27_47_real,
  output     [15:0]   io_coef_out_payload_0_27_47_imag,
  output     [15:0]   io_coef_out_payload_0_27_48_real,
  output     [15:0]   io_coef_out_payload_0_27_48_imag,
  output     [15:0]   io_coef_out_payload_0_27_49_real,
  output     [15:0]   io_coef_out_payload_0_27_49_imag,
  output     [15:0]   io_coef_out_payload_0_28_0_real,
  output     [15:0]   io_coef_out_payload_0_28_0_imag,
  output     [15:0]   io_coef_out_payload_0_28_1_real,
  output     [15:0]   io_coef_out_payload_0_28_1_imag,
  output     [15:0]   io_coef_out_payload_0_28_2_real,
  output     [15:0]   io_coef_out_payload_0_28_2_imag,
  output     [15:0]   io_coef_out_payload_0_28_3_real,
  output     [15:0]   io_coef_out_payload_0_28_3_imag,
  output     [15:0]   io_coef_out_payload_0_28_4_real,
  output     [15:0]   io_coef_out_payload_0_28_4_imag,
  output     [15:0]   io_coef_out_payload_0_28_5_real,
  output     [15:0]   io_coef_out_payload_0_28_5_imag,
  output     [15:0]   io_coef_out_payload_0_28_6_real,
  output     [15:0]   io_coef_out_payload_0_28_6_imag,
  output     [15:0]   io_coef_out_payload_0_28_7_real,
  output     [15:0]   io_coef_out_payload_0_28_7_imag,
  output     [15:0]   io_coef_out_payload_0_28_8_real,
  output     [15:0]   io_coef_out_payload_0_28_8_imag,
  output     [15:0]   io_coef_out_payload_0_28_9_real,
  output     [15:0]   io_coef_out_payload_0_28_9_imag,
  output     [15:0]   io_coef_out_payload_0_28_10_real,
  output     [15:0]   io_coef_out_payload_0_28_10_imag,
  output     [15:0]   io_coef_out_payload_0_28_11_real,
  output     [15:0]   io_coef_out_payload_0_28_11_imag,
  output     [15:0]   io_coef_out_payload_0_28_12_real,
  output     [15:0]   io_coef_out_payload_0_28_12_imag,
  output     [15:0]   io_coef_out_payload_0_28_13_real,
  output     [15:0]   io_coef_out_payload_0_28_13_imag,
  output     [15:0]   io_coef_out_payload_0_28_14_real,
  output     [15:0]   io_coef_out_payload_0_28_14_imag,
  output     [15:0]   io_coef_out_payload_0_28_15_real,
  output     [15:0]   io_coef_out_payload_0_28_15_imag,
  output     [15:0]   io_coef_out_payload_0_28_16_real,
  output     [15:0]   io_coef_out_payload_0_28_16_imag,
  output     [15:0]   io_coef_out_payload_0_28_17_real,
  output     [15:0]   io_coef_out_payload_0_28_17_imag,
  output     [15:0]   io_coef_out_payload_0_28_18_real,
  output     [15:0]   io_coef_out_payload_0_28_18_imag,
  output     [15:0]   io_coef_out_payload_0_28_19_real,
  output     [15:0]   io_coef_out_payload_0_28_19_imag,
  output     [15:0]   io_coef_out_payload_0_28_20_real,
  output     [15:0]   io_coef_out_payload_0_28_20_imag,
  output     [15:0]   io_coef_out_payload_0_28_21_real,
  output     [15:0]   io_coef_out_payload_0_28_21_imag,
  output     [15:0]   io_coef_out_payload_0_28_22_real,
  output     [15:0]   io_coef_out_payload_0_28_22_imag,
  output     [15:0]   io_coef_out_payload_0_28_23_real,
  output     [15:0]   io_coef_out_payload_0_28_23_imag,
  output     [15:0]   io_coef_out_payload_0_28_24_real,
  output     [15:0]   io_coef_out_payload_0_28_24_imag,
  output     [15:0]   io_coef_out_payload_0_28_25_real,
  output     [15:0]   io_coef_out_payload_0_28_25_imag,
  output     [15:0]   io_coef_out_payload_0_28_26_real,
  output     [15:0]   io_coef_out_payload_0_28_26_imag,
  output     [15:0]   io_coef_out_payload_0_28_27_real,
  output     [15:0]   io_coef_out_payload_0_28_27_imag,
  output     [15:0]   io_coef_out_payload_0_28_28_real,
  output     [15:0]   io_coef_out_payload_0_28_28_imag,
  output     [15:0]   io_coef_out_payload_0_28_29_real,
  output     [15:0]   io_coef_out_payload_0_28_29_imag,
  output     [15:0]   io_coef_out_payload_0_28_30_real,
  output     [15:0]   io_coef_out_payload_0_28_30_imag,
  output     [15:0]   io_coef_out_payload_0_28_31_real,
  output     [15:0]   io_coef_out_payload_0_28_31_imag,
  output     [15:0]   io_coef_out_payload_0_28_32_real,
  output     [15:0]   io_coef_out_payload_0_28_32_imag,
  output     [15:0]   io_coef_out_payload_0_28_33_real,
  output     [15:0]   io_coef_out_payload_0_28_33_imag,
  output     [15:0]   io_coef_out_payload_0_28_34_real,
  output     [15:0]   io_coef_out_payload_0_28_34_imag,
  output     [15:0]   io_coef_out_payload_0_28_35_real,
  output     [15:0]   io_coef_out_payload_0_28_35_imag,
  output     [15:0]   io_coef_out_payload_0_28_36_real,
  output     [15:0]   io_coef_out_payload_0_28_36_imag,
  output     [15:0]   io_coef_out_payload_0_28_37_real,
  output     [15:0]   io_coef_out_payload_0_28_37_imag,
  output     [15:0]   io_coef_out_payload_0_28_38_real,
  output     [15:0]   io_coef_out_payload_0_28_38_imag,
  output     [15:0]   io_coef_out_payload_0_28_39_real,
  output     [15:0]   io_coef_out_payload_0_28_39_imag,
  output     [15:0]   io_coef_out_payload_0_28_40_real,
  output     [15:0]   io_coef_out_payload_0_28_40_imag,
  output     [15:0]   io_coef_out_payload_0_28_41_real,
  output     [15:0]   io_coef_out_payload_0_28_41_imag,
  output     [15:0]   io_coef_out_payload_0_28_42_real,
  output     [15:0]   io_coef_out_payload_0_28_42_imag,
  output     [15:0]   io_coef_out_payload_0_28_43_real,
  output     [15:0]   io_coef_out_payload_0_28_43_imag,
  output     [15:0]   io_coef_out_payload_0_28_44_real,
  output     [15:0]   io_coef_out_payload_0_28_44_imag,
  output     [15:0]   io_coef_out_payload_0_28_45_real,
  output     [15:0]   io_coef_out_payload_0_28_45_imag,
  output     [15:0]   io_coef_out_payload_0_28_46_real,
  output     [15:0]   io_coef_out_payload_0_28_46_imag,
  output     [15:0]   io_coef_out_payload_0_28_47_real,
  output     [15:0]   io_coef_out_payload_0_28_47_imag,
  output     [15:0]   io_coef_out_payload_0_28_48_real,
  output     [15:0]   io_coef_out_payload_0_28_48_imag,
  output     [15:0]   io_coef_out_payload_0_28_49_real,
  output     [15:0]   io_coef_out_payload_0_28_49_imag,
  output     [15:0]   io_coef_out_payload_0_29_0_real,
  output     [15:0]   io_coef_out_payload_0_29_0_imag,
  output     [15:0]   io_coef_out_payload_0_29_1_real,
  output     [15:0]   io_coef_out_payload_0_29_1_imag,
  output     [15:0]   io_coef_out_payload_0_29_2_real,
  output     [15:0]   io_coef_out_payload_0_29_2_imag,
  output     [15:0]   io_coef_out_payload_0_29_3_real,
  output     [15:0]   io_coef_out_payload_0_29_3_imag,
  output     [15:0]   io_coef_out_payload_0_29_4_real,
  output     [15:0]   io_coef_out_payload_0_29_4_imag,
  output     [15:0]   io_coef_out_payload_0_29_5_real,
  output     [15:0]   io_coef_out_payload_0_29_5_imag,
  output     [15:0]   io_coef_out_payload_0_29_6_real,
  output     [15:0]   io_coef_out_payload_0_29_6_imag,
  output     [15:0]   io_coef_out_payload_0_29_7_real,
  output     [15:0]   io_coef_out_payload_0_29_7_imag,
  output     [15:0]   io_coef_out_payload_0_29_8_real,
  output     [15:0]   io_coef_out_payload_0_29_8_imag,
  output     [15:0]   io_coef_out_payload_0_29_9_real,
  output     [15:0]   io_coef_out_payload_0_29_9_imag,
  output     [15:0]   io_coef_out_payload_0_29_10_real,
  output     [15:0]   io_coef_out_payload_0_29_10_imag,
  output     [15:0]   io_coef_out_payload_0_29_11_real,
  output     [15:0]   io_coef_out_payload_0_29_11_imag,
  output     [15:0]   io_coef_out_payload_0_29_12_real,
  output     [15:0]   io_coef_out_payload_0_29_12_imag,
  output     [15:0]   io_coef_out_payload_0_29_13_real,
  output     [15:0]   io_coef_out_payload_0_29_13_imag,
  output     [15:0]   io_coef_out_payload_0_29_14_real,
  output     [15:0]   io_coef_out_payload_0_29_14_imag,
  output     [15:0]   io_coef_out_payload_0_29_15_real,
  output     [15:0]   io_coef_out_payload_0_29_15_imag,
  output     [15:0]   io_coef_out_payload_0_29_16_real,
  output     [15:0]   io_coef_out_payload_0_29_16_imag,
  output     [15:0]   io_coef_out_payload_0_29_17_real,
  output     [15:0]   io_coef_out_payload_0_29_17_imag,
  output     [15:0]   io_coef_out_payload_0_29_18_real,
  output     [15:0]   io_coef_out_payload_0_29_18_imag,
  output     [15:0]   io_coef_out_payload_0_29_19_real,
  output     [15:0]   io_coef_out_payload_0_29_19_imag,
  output     [15:0]   io_coef_out_payload_0_29_20_real,
  output     [15:0]   io_coef_out_payload_0_29_20_imag,
  output     [15:0]   io_coef_out_payload_0_29_21_real,
  output     [15:0]   io_coef_out_payload_0_29_21_imag,
  output     [15:0]   io_coef_out_payload_0_29_22_real,
  output     [15:0]   io_coef_out_payload_0_29_22_imag,
  output     [15:0]   io_coef_out_payload_0_29_23_real,
  output     [15:0]   io_coef_out_payload_0_29_23_imag,
  output     [15:0]   io_coef_out_payload_0_29_24_real,
  output     [15:0]   io_coef_out_payload_0_29_24_imag,
  output     [15:0]   io_coef_out_payload_0_29_25_real,
  output     [15:0]   io_coef_out_payload_0_29_25_imag,
  output     [15:0]   io_coef_out_payload_0_29_26_real,
  output     [15:0]   io_coef_out_payload_0_29_26_imag,
  output     [15:0]   io_coef_out_payload_0_29_27_real,
  output     [15:0]   io_coef_out_payload_0_29_27_imag,
  output     [15:0]   io_coef_out_payload_0_29_28_real,
  output     [15:0]   io_coef_out_payload_0_29_28_imag,
  output     [15:0]   io_coef_out_payload_0_29_29_real,
  output     [15:0]   io_coef_out_payload_0_29_29_imag,
  output     [15:0]   io_coef_out_payload_0_29_30_real,
  output     [15:0]   io_coef_out_payload_0_29_30_imag,
  output     [15:0]   io_coef_out_payload_0_29_31_real,
  output     [15:0]   io_coef_out_payload_0_29_31_imag,
  output     [15:0]   io_coef_out_payload_0_29_32_real,
  output     [15:0]   io_coef_out_payload_0_29_32_imag,
  output     [15:0]   io_coef_out_payload_0_29_33_real,
  output     [15:0]   io_coef_out_payload_0_29_33_imag,
  output     [15:0]   io_coef_out_payload_0_29_34_real,
  output     [15:0]   io_coef_out_payload_0_29_34_imag,
  output     [15:0]   io_coef_out_payload_0_29_35_real,
  output     [15:0]   io_coef_out_payload_0_29_35_imag,
  output     [15:0]   io_coef_out_payload_0_29_36_real,
  output     [15:0]   io_coef_out_payload_0_29_36_imag,
  output     [15:0]   io_coef_out_payload_0_29_37_real,
  output     [15:0]   io_coef_out_payload_0_29_37_imag,
  output     [15:0]   io_coef_out_payload_0_29_38_real,
  output     [15:0]   io_coef_out_payload_0_29_38_imag,
  output     [15:0]   io_coef_out_payload_0_29_39_real,
  output     [15:0]   io_coef_out_payload_0_29_39_imag,
  output     [15:0]   io_coef_out_payload_0_29_40_real,
  output     [15:0]   io_coef_out_payload_0_29_40_imag,
  output     [15:0]   io_coef_out_payload_0_29_41_real,
  output     [15:0]   io_coef_out_payload_0_29_41_imag,
  output     [15:0]   io_coef_out_payload_0_29_42_real,
  output     [15:0]   io_coef_out_payload_0_29_42_imag,
  output     [15:0]   io_coef_out_payload_0_29_43_real,
  output     [15:0]   io_coef_out_payload_0_29_43_imag,
  output     [15:0]   io_coef_out_payload_0_29_44_real,
  output     [15:0]   io_coef_out_payload_0_29_44_imag,
  output     [15:0]   io_coef_out_payload_0_29_45_real,
  output     [15:0]   io_coef_out_payload_0_29_45_imag,
  output     [15:0]   io_coef_out_payload_0_29_46_real,
  output     [15:0]   io_coef_out_payload_0_29_46_imag,
  output     [15:0]   io_coef_out_payload_0_29_47_real,
  output     [15:0]   io_coef_out_payload_0_29_47_imag,
  output     [15:0]   io_coef_out_payload_0_29_48_real,
  output     [15:0]   io_coef_out_payload_0_29_48_imag,
  output     [15:0]   io_coef_out_payload_0_29_49_real,
  output     [15:0]   io_coef_out_payload_0_29_49_imag,
  output     [15:0]   io_coef_out_payload_0_30_0_real,
  output     [15:0]   io_coef_out_payload_0_30_0_imag,
  output     [15:0]   io_coef_out_payload_0_30_1_real,
  output     [15:0]   io_coef_out_payload_0_30_1_imag,
  output     [15:0]   io_coef_out_payload_0_30_2_real,
  output     [15:0]   io_coef_out_payload_0_30_2_imag,
  output     [15:0]   io_coef_out_payload_0_30_3_real,
  output     [15:0]   io_coef_out_payload_0_30_3_imag,
  output     [15:0]   io_coef_out_payload_0_30_4_real,
  output     [15:0]   io_coef_out_payload_0_30_4_imag,
  output     [15:0]   io_coef_out_payload_0_30_5_real,
  output     [15:0]   io_coef_out_payload_0_30_5_imag,
  output     [15:0]   io_coef_out_payload_0_30_6_real,
  output     [15:0]   io_coef_out_payload_0_30_6_imag,
  output     [15:0]   io_coef_out_payload_0_30_7_real,
  output     [15:0]   io_coef_out_payload_0_30_7_imag,
  output     [15:0]   io_coef_out_payload_0_30_8_real,
  output     [15:0]   io_coef_out_payload_0_30_8_imag,
  output     [15:0]   io_coef_out_payload_0_30_9_real,
  output     [15:0]   io_coef_out_payload_0_30_9_imag,
  output     [15:0]   io_coef_out_payload_0_30_10_real,
  output     [15:0]   io_coef_out_payload_0_30_10_imag,
  output     [15:0]   io_coef_out_payload_0_30_11_real,
  output     [15:0]   io_coef_out_payload_0_30_11_imag,
  output     [15:0]   io_coef_out_payload_0_30_12_real,
  output     [15:0]   io_coef_out_payload_0_30_12_imag,
  output     [15:0]   io_coef_out_payload_0_30_13_real,
  output     [15:0]   io_coef_out_payload_0_30_13_imag,
  output     [15:0]   io_coef_out_payload_0_30_14_real,
  output     [15:0]   io_coef_out_payload_0_30_14_imag,
  output     [15:0]   io_coef_out_payload_0_30_15_real,
  output     [15:0]   io_coef_out_payload_0_30_15_imag,
  output     [15:0]   io_coef_out_payload_0_30_16_real,
  output     [15:0]   io_coef_out_payload_0_30_16_imag,
  output     [15:0]   io_coef_out_payload_0_30_17_real,
  output     [15:0]   io_coef_out_payload_0_30_17_imag,
  output     [15:0]   io_coef_out_payload_0_30_18_real,
  output     [15:0]   io_coef_out_payload_0_30_18_imag,
  output     [15:0]   io_coef_out_payload_0_30_19_real,
  output     [15:0]   io_coef_out_payload_0_30_19_imag,
  output     [15:0]   io_coef_out_payload_0_30_20_real,
  output     [15:0]   io_coef_out_payload_0_30_20_imag,
  output     [15:0]   io_coef_out_payload_0_30_21_real,
  output     [15:0]   io_coef_out_payload_0_30_21_imag,
  output     [15:0]   io_coef_out_payload_0_30_22_real,
  output     [15:0]   io_coef_out_payload_0_30_22_imag,
  output     [15:0]   io_coef_out_payload_0_30_23_real,
  output     [15:0]   io_coef_out_payload_0_30_23_imag,
  output     [15:0]   io_coef_out_payload_0_30_24_real,
  output     [15:0]   io_coef_out_payload_0_30_24_imag,
  output     [15:0]   io_coef_out_payload_0_30_25_real,
  output     [15:0]   io_coef_out_payload_0_30_25_imag,
  output     [15:0]   io_coef_out_payload_0_30_26_real,
  output     [15:0]   io_coef_out_payload_0_30_26_imag,
  output     [15:0]   io_coef_out_payload_0_30_27_real,
  output     [15:0]   io_coef_out_payload_0_30_27_imag,
  output     [15:0]   io_coef_out_payload_0_30_28_real,
  output     [15:0]   io_coef_out_payload_0_30_28_imag,
  output     [15:0]   io_coef_out_payload_0_30_29_real,
  output     [15:0]   io_coef_out_payload_0_30_29_imag,
  output     [15:0]   io_coef_out_payload_0_30_30_real,
  output     [15:0]   io_coef_out_payload_0_30_30_imag,
  output     [15:0]   io_coef_out_payload_0_30_31_real,
  output     [15:0]   io_coef_out_payload_0_30_31_imag,
  output     [15:0]   io_coef_out_payload_0_30_32_real,
  output     [15:0]   io_coef_out_payload_0_30_32_imag,
  output     [15:0]   io_coef_out_payload_0_30_33_real,
  output     [15:0]   io_coef_out_payload_0_30_33_imag,
  output     [15:0]   io_coef_out_payload_0_30_34_real,
  output     [15:0]   io_coef_out_payload_0_30_34_imag,
  output     [15:0]   io_coef_out_payload_0_30_35_real,
  output     [15:0]   io_coef_out_payload_0_30_35_imag,
  output     [15:0]   io_coef_out_payload_0_30_36_real,
  output     [15:0]   io_coef_out_payload_0_30_36_imag,
  output     [15:0]   io_coef_out_payload_0_30_37_real,
  output     [15:0]   io_coef_out_payload_0_30_37_imag,
  output     [15:0]   io_coef_out_payload_0_30_38_real,
  output     [15:0]   io_coef_out_payload_0_30_38_imag,
  output     [15:0]   io_coef_out_payload_0_30_39_real,
  output     [15:0]   io_coef_out_payload_0_30_39_imag,
  output     [15:0]   io_coef_out_payload_0_30_40_real,
  output     [15:0]   io_coef_out_payload_0_30_40_imag,
  output     [15:0]   io_coef_out_payload_0_30_41_real,
  output     [15:0]   io_coef_out_payload_0_30_41_imag,
  output     [15:0]   io_coef_out_payload_0_30_42_real,
  output     [15:0]   io_coef_out_payload_0_30_42_imag,
  output     [15:0]   io_coef_out_payload_0_30_43_real,
  output     [15:0]   io_coef_out_payload_0_30_43_imag,
  output     [15:0]   io_coef_out_payload_0_30_44_real,
  output     [15:0]   io_coef_out_payload_0_30_44_imag,
  output     [15:0]   io_coef_out_payload_0_30_45_real,
  output     [15:0]   io_coef_out_payload_0_30_45_imag,
  output     [15:0]   io_coef_out_payload_0_30_46_real,
  output     [15:0]   io_coef_out_payload_0_30_46_imag,
  output     [15:0]   io_coef_out_payload_0_30_47_real,
  output     [15:0]   io_coef_out_payload_0_30_47_imag,
  output     [15:0]   io_coef_out_payload_0_30_48_real,
  output     [15:0]   io_coef_out_payload_0_30_48_imag,
  output     [15:0]   io_coef_out_payload_0_30_49_real,
  output     [15:0]   io_coef_out_payload_0_30_49_imag,
  output     [15:0]   io_coef_out_payload_0_31_0_real,
  output     [15:0]   io_coef_out_payload_0_31_0_imag,
  output     [15:0]   io_coef_out_payload_0_31_1_real,
  output     [15:0]   io_coef_out_payload_0_31_1_imag,
  output     [15:0]   io_coef_out_payload_0_31_2_real,
  output     [15:0]   io_coef_out_payload_0_31_2_imag,
  output     [15:0]   io_coef_out_payload_0_31_3_real,
  output     [15:0]   io_coef_out_payload_0_31_3_imag,
  output     [15:0]   io_coef_out_payload_0_31_4_real,
  output     [15:0]   io_coef_out_payload_0_31_4_imag,
  output     [15:0]   io_coef_out_payload_0_31_5_real,
  output     [15:0]   io_coef_out_payload_0_31_5_imag,
  output     [15:0]   io_coef_out_payload_0_31_6_real,
  output     [15:0]   io_coef_out_payload_0_31_6_imag,
  output     [15:0]   io_coef_out_payload_0_31_7_real,
  output     [15:0]   io_coef_out_payload_0_31_7_imag,
  output     [15:0]   io_coef_out_payload_0_31_8_real,
  output     [15:0]   io_coef_out_payload_0_31_8_imag,
  output     [15:0]   io_coef_out_payload_0_31_9_real,
  output     [15:0]   io_coef_out_payload_0_31_9_imag,
  output     [15:0]   io_coef_out_payload_0_31_10_real,
  output     [15:0]   io_coef_out_payload_0_31_10_imag,
  output     [15:0]   io_coef_out_payload_0_31_11_real,
  output     [15:0]   io_coef_out_payload_0_31_11_imag,
  output     [15:0]   io_coef_out_payload_0_31_12_real,
  output     [15:0]   io_coef_out_payload_0_31_12_imag,
  output     [15:0]   io_coef_out_payload_0_31_13_real,
  output     [15:0]   io_coef_out_payload_0_31_13_imag,
  output     [15:0]   io_coef_out_payload_0_31_14_real,
  output     [15:0]   io_coef_out_payload_0_31_14_imag,
  output     [15:0]   io_coef_out_payload_0_31_15_real,
  output     [15:0]   io_coef_out_payload_0_31_15_imag,
  output     [15:0]   io_coef_out_payload_0_31_16_real,
  output     [15:0]   io_coef_out_payload_0_31_16_imag,
  output     [15:0]   io_coef_out_payload_0_31_17_real,
  output     [15:0]   io_coef_out_payload_0_31_17_imag,
  output     [15:0]   io_coef_out_payload_0_31_18_real,
  output     [15:0]   io_coef_out_payload_0_31_18_imag,
  output     [15:0]   io_coef_out_payload_0_31_19_real,
  output     [15:0]   io_coef_out_payload_0_31_19_imag,
  output     [15:0]   io_coef_out_payload_0_31_20_real,
  output     [15:0]   io_coef_out_payload_0_31_20_imag,
  output     [15:0]   io_coef_out_payload_0_31_21_real,
  output     [15:0]   io_coef_out_payload_0_31_21_imag,
  output     [15:0]   io_coef_out_payload_0_31_22_real,
  output     [15:0]   io_coef_out_payload_0_31_22_imag,
  output     [15:0]   io_coef_out_payload_0_31_23_real,
  output     [15:0]   io_coef_out_payload_0_31_23_imag,
  output     [15:0]   io_coef_out_payload_0_31_24_real,
  output     [15:0]   io_coef_out_payload_0_31_24_imag,
  output     [15:0]   io_coef_out_payload_0_31_25_real,
  output     [15:0]   io_coef_out_payload_0_31_25_imag,
  output     [15:0]   io_coef_out_payload_0_31_26_real,
  output     [15:0]   io_coef_out_payload_0_31_26_imag,
  output     [15:0]   io_coef_out_payload_0_31_27_real,
  output     [15:0]   io_coef_out_payload_0_31_27_imag,
  output     [15:0]   io_coef_out_payload_0_31_28_real,
  output     [15:0]   io_coef_out_payload_0_31_28_imag,
  output     [15:0]   io_coef_out_payload_0_31_29_real,
  output     [15:0]   io_coef_out_payload_0_31_29_imag,
  output     [15:0]   io_coef_out_payload_0_31_30_real,
  output     [15:0]   io_coef_out_payload_0_31_30_imag,
  output     [15:0]   io_coef_out_payload_0_31_31_real,
  output     [15:0]   io_coef_out_payload_0_31_31_imag,
  output     [15:0]   io_coef_out_payload_0_31_32_real,
  output     [15:0]   io_coef_out_payload_0_31_32_imag,
  output     [15:0]   io_coef_out_payload_0_31_33_real,
  output     [15:0]   io_coef_out_payload_0_31_33_imag,
  output     [15:0]   io_coef_out_payload_0_31_34_real,
  output     [15:0]   io_coef_out_payload_0_31_34_imag,
  output     [15:0]   io_coef_out_payload_0_31_35_real,
  output     [15:0]   io_coef_out_payload_0_31_35_imag,
  output     [15:0]   io_coef_out_payload_0_31_36_real,
  output     [15:0]   io_coef_out_payload_0_31_36_imag,
  output     [15:0]   io_coef_out_payload_0_31_37_real,
  output     [15:0]   io_coef_out_payload_0_31_37_imag,
  output     [15:0]   io_coef_out_payload_0_31_38_real,
  output     [15:0]   io_coef_out_payload_0_31_38_imag,
  output     [15:0]   io_coef_out_payload_0_31_39_real,
  output     [15:0]   io_coef_out_payload_0_31_39_imag,
  output     [15:0]   io_coef_out_payload_0_31_40_real,
  output     [15:0]   io_coef_out_payload_0_31_40_imag,
  output     [15:0]   io_coef_out_payload_0_31_41_real,
  output     [15:0]   io_coef_out_payload_0_31_41_imag,
  output     [15:0]   io_coef_out_payload_0_31_42_real,
  output     [15:0]   io_coef_out_payload_0_31_42_imag,
  output     [15:0]   io_coef_out_payload_0_31_43_real,
  output     [15:0]   io_coef_out_payload_0_31_43_imag,
  output     [15:0]   io_coef_out_payload_0_31_44_real,
  output     [15:0]   io_coef_out_payload_0_31_44_imag,
  output     [15:0]   io_coef_out_payload_0_31_45_real,
  output     [15:0]   io_coef_out_payload_0_31_45_imag,
  output     [15:0]   io_coef_out_payload_0_31_46_real,
  output     [15:0]   io_coef_out_payload_0_31_46_imag,
  output     [15:0]   io_coef_out_payload_0_31_47_real,
  output     [15:0]   io_coef_out_payload_0_31_47_imag,
  output     [15:0]   io_coef_out_payload_0_31_48_real,
  output     [15:0]   io_coef_out_payload_0_31_48_imag,
  output     [15:0]   io_coef_out_payload_0_31_49_real,
  output     [15:0]   io_coef_out_payload_0_31_49_imag,
  output     [15:0]   io_coef_out_payload_0_32_0_real,
  output     [15:0]   io_coef_out_payload_0_32_0_imag,
  output     [15:0]   io_coef_out_payload_0_32_1_real,
  output     [15:0]   io_coef_out_payload_0_32_1_imag,
  output     [15:0]   io_coef_out_payload_0_32_2_real,
  output     [15:0]   io_coef_out_payload_0_32_2_imag,
  output     [15:0]   io_coef_out_payload_0_32_3_real,
  output     [15:0]   io_coef_out_payload_0_32_3_imag,
  output     [15:0]   io_coef_out_payload_0_32_4_real,
  output     [15:0]   io_coef_out_payload_0_32_4_imag,
  output     [15:0]   io_coef_out_payload_0_32_5_real,
  output     [15:0]   io_coef_out_payload_0_32_5_imag,
  output     [15:0]   io_coef_out_payload_0_32_6_real,
  output     [15:0]   io_coef_out_payload_0_32_6_imag,
  output     [15:0]   io_coef_out_payload_0_32_7_real,
  output     [15:0]   io_coef_out_payload_0_32_7_imag,
  output     [15:0]   io_coef_out_payload_0_32_8_real,
  output     [15:0]   io_coef_out_payload_0_32_8_imag,
  output     [15:0]   io_coef_out_payload_0_32_9_real,
  output     [15:0]   io_coef_out_payload_0_32_9_imag,
  output     [15:0]   io_coef_out_payload_0_32_10_real,
  output     [15:0]   io_coef_out_payload_0_32_10_imag,
  output     [15:0]   io_coef_out_payload_0_32_11_real,
  output     [15:0]   io_coef_out_payload_0_32_11_imag,
  output     [15:0]   io_coef_out_payload_0_32_12_real,
  output     [15:0]   io_coef_out_payload_0_32_12_imag,
  output     [15:0]   io_coef_out_payload_0_32_13_real,
  output     [15:0]   io_coef_out_payload_0_32_13_imag,
  output     [15:0]   io_coef_out_payload_0_32_14_real,
  output     [15:0]   io_coef_out_payload_0_32_14_imag,
  output     [15:0]   io_coef_out_payload_0_32_15_real,
  output     [15:0]   io_coef_out_payload_0_32_15_imag,
  output     [15:0]   io_coef_out_payload_0_32_16_real,
  output     [15:0]   io_coef_out_payload_0_32_16_imag,
  output     [15:0]   io_coef_out_payload_0_32_17_real,
  output     [15:0]   io_coef_out_payload_0_32_17_imag,
  output     [15:0]   io_coef_out_payload_0_32_18_real,
  output     [15:0]   io_coef_out_payload_0_32_18_imag,
  output     [15:0]   io_coef_out_payload_0_32_19_real,
  output     [15:0]   io_coef_out_payload_0_32_19_imag,
  output     [15:0]   io_coef_out_payload_0_32_20_real,
  output     [15:0]   io_coef_out_payload_0_32_20_imag,
  output     [15:0]   io_coef_out_payload_0_32_21_real,
  output     [15:0]   io_coef_out_payload_0_32_21_imag,
  output     [15:0]   io_coef_out_payload_0_32_22_real,
  output     [15:0]   io_coef_out_payload_0_32_22_imag,
  output     [15:0]   io_coef_out_payload_0_32_23_real,
  output     [15:0]   io_coef_out_payload_0_32_23_imag,
  output     [15:0]   io_coef_out_payload_0_32_24_real,
  output     [15:0]   io_coef_out_payload_0_32_24_imag,
  output     [15:0]   io_coef_out_payload_0_32_25_real,
  output     [15:0]   io_coef_out_payload_0_32_25_imag,
  output     [15:0]   io_coef_out_payload_0_32_26_real,
  output     [15:0]   io_coef_out_payload_0_32_26_imag,
  output     [15:0]   io_coef_out_payload_0_32_27_real,
  output     [15:0]   io_coef_out_payload_0_32_27_imag,
  output     [15:0]   io_coef_out_payload_0_32_28_real,
  output     [15:0]   io_coef_out_payload_0_32_28_imag,
  output     [15:0]   io_coef_out_payload_0_32_29_real,
  output     [15:0]   io_coef_out_payload_0_32_29_imag,
  output     [15:0]   io_coef_out_payload_0_32_30_real,
  output     [15:0]   io_coef_out_payload_0_32_30_imag,
  output     [15:0]   io_coef_out_payload_0_32_31_real,
  output     [15:0]   io_coef_out_payload_0_32_31_imag,
  output     [15:0]   io_coef_out_payload_0_32_32_real,
  output     [15:0]   io_coef_out_payload_0_32_32_imag,
  output     [15:0]   io_coef_out_payload_0_32_33_real,
  output     [15:0]   io_coef_out_payload_0_32_33_imag,
  output     [15:0]   io_coef_out_payload_0_32_34_real,
  output     [15:0]   io_coef_out_payload_0_32_34_imag,
  output     [15:0]   io_coef_out_payload_0_32_35_real,
  output     [15:0]   io_coef_out_payload_0_32_35_imag,
  output     [15:0]   io_coef_out_payload_0_32_36_real,
  output     [15:0]   io_coef_out_payload_0_32_36_imag,
  output     [15:0]   io_coef_out_payload_0_32_37_real,
  output     [15:0]   io_coef_out_payload_0_32_37_imag,
  output     [15:0]   io_coef_out_payload_0_32_38_real,
  output     [15:0]   io_coef_out_payload_0_32_38_imag,
  output     [15:0]   io_coef_out_payload_0_32_39_real,
  output     [15:0]   io_coef_out_payload_0_32_39_imag,
  output     [15:0]   io_coef_out_payload_0_32_40_real,
  output     [15:0]   io_coef_out_payload_0_32_40_imag,
  output     [15:0]   io_coef_out_payload_0_32_41_real,
  output     [15:0]   io_coef_out_payload_0_32_41_imag,
  output     [15:0]   io_coef_out_payload_0_32_42_real,
  output     [15:0]   io_coef_out_payload_0_32_42_imag,
  output     [15:0]   io_coef_out_payload_0_32_43_real,
  output     [15:0]   io_coef_out_payload_0_32_43_imag,
  output     [15:0]   io_coef_out_payload_0_32_44_real,
  output     [15:0]   io_coef_out_payload_0_32_44_imag,
  output     [15:0]   io_coef_out_payload_0_32_45_real,
  output     [15:0]   io_coef_out_payload_0_32_45_imag,
  output     [15:0]   io_coef_out_payload_0_32_46_real,
  output     [15:0]   io_coef_out_payload_0_32_46_imag,
  output     [15:0]   io_coef_out_payload_0_32_47_real,
  output     [15:0]   io_coef_out_payload_0_32_47_imag,
  output     [15:0]   io_coef_out_payload_0_32_48_real,
  output     [15:0]   io_coef_out_payload_0_32_48_imag,
  output     [15:0]   io_coef_out_payload_0_32_49_real,
  output     [15:0]   io_coef_out_payload_0_32_49_imag,
  output     [15:0]   io_coef_out_payload_0_33_0_real,
  output     [15:0]   io_coef_out_payload_0_33_0_imag,
  output     [15:0]   io_coef_out_payload_0_33_1_real,
  output     [15:0]   io_coef_out_payload_0_33_1_imag,
  output     [15:0]   io_coef_out_payload_0_33_2_real,
  output     [15:0]   io_coef_out_payload_0_33_2_imag,
  output     [15:0]   io_coef_out_payload_0_33_3_real,
  output     [15:0]   io_coef_out_payload_0_33_3_imag,
  output     [15:0]   io_coef_out_payload_0_33_4_real,
  output     [15:0]   io_coef_out_payload_0_33_4_imag,
  output     [15:0]   io_coef_out_payload_0_33_5_real,
  output     [15:0]   io_coef_out_payload_0_33_5_imag,
  output     [15:0]   io_coef_out_payload_0_33_6_real,
  output     [15:0]   io_coef_out_payload_0_33_6_imag,
  output     [15:0]   io_coef_out_payload_0_33_7_real,
  output     [15:0]   io_coef_out_payload_0_33_7_imag,
  output     [15:0]   io_coef_out_payload_0_33_8_real,
  output     [15:0]   io_coef_out_payload_0_33_8_imag,
  output     [15:0]   io_coef_out_payload_0_33_9_real,
  output     [15:0]   io_coef_out_payload_0_33_9_imag,
  output     [15:0]   io_coef_out_payload_0_33_10_real,
  output     [15:0]   io_coef_out_payload_0_33_10_imag,
  output     [15:0]   io_coef_out_payload_0_33_11_real,
  output     [15:0]   io_coef_out_payload_0_33_11_imag,
  output     [15:0]   io_coef_out_payload_0_33_12_real,
  output     [15:0]   io_coef_out_payload_0_33_12_imag,
  output     [15:0]   io_coef_out_payload_0_33_13_real,
  output     [15:0]   io_coef_out_payload_0_33_13_imag,
  output     [15:0]   io_coef_out_payload_0_33_14_real,
  output     [15:0]   io_coef_out_payload_0_33_14_imag,
  output     [15:0]   io_coef_out_payload_0_33_15_real,
  output     [15:0]   io_coef_out_payload_0_33_15_imag,
  output     [15:0]   io_coef_out_payload_0_33_16_real,
  output     [15:0]   io_coef_out_payload_0_33_16_imag,
  output     [15:0]   io_coef_out_payload_0_33_17_real,
  output     [15:0]   io_coef_out_payload_0_33_17_imag,
  output     [15:0]   io_coef_out_payload_0_33_18_real,
  output     [15:0]   io_coef_out_payload_0_33_18_imag,
  output     [15:0]   io_coef_out_payload_0_33_19_real,
  output     [15:0]   io_coef_out_payload_0_33_19_imag,
  output     [15:0]   io_coef_out_payload_0_33_20_real,
  output     [15:0]   io_coef_out_payload_0_33_20_imag,
  output     [15:0]   io_coef_out_payload_0_33_21_real,
  output     [15:0]   io_coef_out_payload_0_33_21_imag,
  output     [15:0]   io_coef_out_payload_0_33_22_real,
  output     [15:0]   io_coef_out_payload_0_33_22_imag,
  output     [15:0]   io_coef_out_payload_0_33_23_real,
  output     [15:0]   io_coef_out_payload_0_33_23_imag,
  output     [15:0]   io_coef_out_payload_0_33_24_real,
  output     [15:0]   io_coef_out_payload_0_33_24_imag,
  output     [15:0]   io_coef_out_payload_0_33_25_real,
  output     [15:0]   io_coef_out_payload_0_33_25_imag,
  output     [15:0]   io_coef_out_payload_0_33_26_real,
  output     [15:0]   io_coef_out_payload_0_33_26_imag,
  output     [15:0]   io_coef_out_payload_0_33_27_real,
  output     [15:0]   io_coef_out_payload_0_33_27_imag,
  output     [15:0]   io_coef_out_payload_0_33_28_real,
  output     [15:0]   io_coef_out_payload_0_33_28_imag,
  output     [15:0]   io_coef_out_payload_0_33_29_real,
  output     [15:0]   io_coef_out_payload_0_33_29_imag,
  output     [15:0]   io_coef_out_payload_0_33_30_real,
  output     [15:0]   io_coef_out_payload_0_33_30_imag,
  output     [15:0]   io_coef_out_payload_0_33_31_real,
  output     [15:0]   io_coef_out_payload_0_33_31_imag,
  output     [15:0]   io_coef_out_payload_0_33_32_real,
  output     [15:0]   io_coef_out_payload_0_33_32_imag,
  output     [15:0]   io_coef_out_payload_0_33_33_real,
  output     [15:0]   io_coef_out_payload_0_33_33_imag,
  output     [15:0]   io_coef_out_payload_0_33_34_real,
  output     [15:0]   io_coef_out_payload_0_33_34_imag,
  output     [15:0]   io_coef_out_payload_0_33_35_real,
  output     [15:0]   io_coef_out_payload_0_33_35_imag,
  output     [15:0]   io_coef_out_payload_0_33_36_real,
  output     [15:0]   io_coef_out_payload_0_33_36_imag,
  output     [15:0]   io_coef_out_payload_0_33_37_real,
  output     [15:0]   io_coef_out_payload_0_33_37_imag,
  output     [15:0]   io_coef_out_payload_0_33_38_real,
  output     [15:0]   io_coef_out_payload_0_33_38_imag,
  output     [15:0]   io_coef_out_payload_0_33_39_real,
  output     [15:0]   io_coef_out_payload_0_33_39_imag,
  output     [15:0]   io_coef_out_payload_0_33_40_real,
  output     [15:0]   io_coef_out_payload_0_33_40_imag,
  output     [15:0]   io_coef_out_payload_0_33_41_real,
  output     [15:0]   io_coef_out_payload_0_33_41_imag,
  output     [15:0]   io_coef_out_payload_0_33_42_real,
  output     [15:0]   io_coef_out_payload_0_33_42_imag,
  output     [15:0]   io_coef_out_payload_0_33_43_real,
  output     [15:0]   io_coef_out_payload_0_33_43_imag,
  output     [15:0]   io_coef_out_payload_0_33_44_real,
  output     [15:0]   io_coef_out_payload_0_33_44_imag,
  output     [15:0]   io_coef_out_payload_0_33_45_real,
  output     [15:0]   io_coef_out_payload_0_33_45_imag,
  output     [15:0]   io_coef_out_payload_0_33_46_real,
  output     [15:0]   io_coef_out_payload_0_33_46_imag,
  output     [15:0]   io_coef_out_payload_0_33_47_real,
  output     [15:0]   io_coef_out_payload_0_33_47_imag,
  output     [15:0]   io_coef_out_payload_0_33_48_real,
  output     [15:0]   io_coef_out_payload_0_33_48_imag,
  output     [15:0]   io_coef_out_payload_0_33_49_real,
  output     [15:0]   io_coef_out_payload_0_33_49_imag,
  output     [15:0]   io_coef_out_payload_0_34_0_real,
  output     [15:0]   io_coef_out_payload_0_34_0_imag,
  output     [15:0]   io_coef_out_payload_0_34_1_real,
  output     [15:0]   io_coef_out_payload_0_34_1_imag,
  output     [15:0]   io_coef_out_payload_0_34_2_real,
  output     [15:0]   io_coef_out_payload_0_34_2_imag,
  output     [15:0]   io_coef_out_payload_0_34_3_real,
  output     [15:0]   io_coef_out_payload_0_34_3_imag,
  output     [15:0]   io_coef_out_payload_0_34_4_real,
  output     [15:0]   io_coef_out_payload_0_34_4_imag,
  output     [15:0]   io_coef_out_payload_0_34_5_real,
  output     [15:0]   io_coef_out_payload_0_34_5_imag,
  output     [15:0]   io_coef_out_payload_0_34_6_real,
  output     [15:0]   io_coef_out_payload_0_34_6_imag,
  output     [15:0]   io_coef_out_payload_0_34_7_real,
  output     [15:0]   io_coef_out_payload_0_34_7_imag,
  output     [15:0]   io_coef_out_payload_0_34_8_real,
  output     [15:0]   io_coef_out_payload_0_34_8_imag,
  output     [15:0]   io_coef_out_payload_0_34_9_real,
  output     [15:0]   io_coef_out_payload_0_34_9_imag,
  output     [15:0]   io_coef_out_payload_0_34_10_real,
  output     [15:0]   io_coef_out_payload_0_34_10_imag,
  output     [15:0]   io_coef_out_payload_0_34_11_real,
  output     [15:0]   io_coef_out_payload_0_34_11_imag,
  output     [15:0]   io_coef_out_payload_0_34_12_real,
  output     [15:0]   io_coef_out_payload_0_34_12_imag,
  output     [15:0]   io_coef_out_payload_0_34_13_real,
  output     [15:0]   io_coef_out_payload_0_34_13_imag,
  output     [15:0]   io_coef_out_payload_0_34_14_real,
  output     [15:0]   io_coef_out_payload_0_34_14_imag,
  output     [15:0]   io_coef_out_payload_0_34_15_real,
  output     [15:0]   io_coef_out_payload_0_34_15_imag,
  output     [15:0]   io_coef_out_payload_0_34_16_real,
  output     [15:0]   io_coef_out_payload_0_34_16_imag,
  output     [15:0]   io_coef_out_payload_0_34_17_real,
  output     [15:0]   io_coef_out_payload_0_34_17_imag,
  output     [15:0]   io_coef_out_payload_0_34_18_real,
  output     [15:0]   io_coef_out_payload_0_34_18_imag,
  output     [15:0]   io_coef_out_payload_0_34_19_real,
  output     [15:0]   io_coef_out_payload_0_34_19_imag,
  output     [15:0]   io_coef_out_payload_0_34_20_real,
  output     [15:0]   io_coef_out_payload_0_34_20_imag,
  output     [15:0]   io_coef_out_payload_0_34_21_real,
  output     [15:0]   io_coef_out_payload_0_34_21_imag,
  output     [15:0]   io_coef_out_payload_0_34_22_real,
  output     [15:0]   io_coef_out_payload_0_34_22_imag,
  output     [15:0]   io_coef_out_payload_0_34_23_real,
  output     [15:0]   io_coef_out_payload_0_34_23_imag,
  output     [15:0]   io_coef_out_payload_0_34_24_real,
  output     [15:0]   io_coef_out_payload_0_34_24_imag,
  output     [15:0]   io_coef_out_payload_0_34_25_real,
  output     [15:0]   io_coef_out_payload_0_34_25_imag,
  output     [15:0]   io_coef_out_payload_0_34_26_real,
  output     [15:0]   io_coef_out_payload_0_34_26_imag,
  output     [15:0]   io_coef_out_payload_0_34_27_real,
  output     [15:0]   io_coef_out_payload_0_34_27_imag,
  output     [15:0]   io_coef_out_payload_0_34_28_real,
  output     [15:0]   io_coef_out_payload_0_34_28_imag,
  output     [15:0]   io_coef_out_payload_0_34_29_real,
  output     [15:0]   io_coef_out_payload_0_34_29_imag,
  output     [15:0]   io_coef_out_payload_0_34_30_real,
  output     [15:0]   io_coef_out_payload_0_34_30_imag,
  output     [15:0]   io_coef_out_payload_0_34_31_real,
  output     [15:0]   io_coef_out_payload_0_34_31_imag,
  output     [15:0]   io_coef_out_payload_0_34_32_real,
  output     [15:0]   io_coef_out_payload_0_34_32_imag,
  output     [15:0]   io_coef_out_payload_0_34_33_real,
  output     [15:0]   io_coef_out_payload_0_34_33_imag,
  output     [15:0]   io_coef_out_payload_0_34_34_real,
  output     [15:0]   io_coef_out_payload_0_34_34_imag,
  output     [15:0]   io_coef_out_payload_0_34_35_real,
  output     [15:0]   io_coef_out_payload_0_34_35_imag,
  output     [15:0]   io_coef_out_payload_0_34_36_real,
  output     [15:0]   io_coef_out_payload_0_34_36_imag,
  output     [15:0]   io_coef_out_payload_0_34_37_real,
  output     [15:0]   io_coef_out_payload_0_34_37_imag,
  output     [15:0]   io_coef_out_payload_0_34_38_real,
  output     [15:0]   io_coef_out_payload_0_34_38_imag,
  output     [15:0]   io_coef_out_payload_0_34_39_real,
  output     [15:0]   io_coef_out_payload_0_34_39_imag,
  output     [15:0]   io_coef_out_payload_0_34_40_real,
  output     [15:0]   io_coef_out_payload_0_34_40_imag,
  output     [15:0]   io_coef_out_payload_0_34_41_real,
  output     [15:0]   io_coef_out_payload_0_34_41_imag,
  output     [15:0]   io_coef_out_payload_0_34_42_real,
  output     [15:0]   io_coef_out_payload_0_34_42_imag,
  output     [15:0]   io_coef_out_payload_0_34_43_real,
  output     [15:0]   io_coef_out_payload_0_34_43_imag,
  output     [15:0]   io_coef_out_payload_0_34_44_real,
  output     [15:0]   io_coef_out_payload_0_34_44_imag,
  output     [15:0]   io_coef_out_payload_0_34_45_real,
  output     [15:0]   io_coef_out_payload_0_34_45_imag,
  output     [15:0]   io_coef_out_payload_0_34_46_real,
  output     [15:0]   io_coef_out_payload_0_34_46_imag,
  output     [15:0]   io_coef_out_payload_0_34_47_real,
  output     [15:0]   io_coef_out_payload_0_34_47_imag,
  output     [15:0]   io_coef_out_payload_0_34_48_real,
  output     [15:0]   io_coef_out_payload_0_34_48_imag,
  output     [15:0]   io_coef_out_payload_0_34_49_real,
  output     [15:0]   io_coef_out_payload_0_34_49_imag,
  output     [15:0]   io_coef_out_payload_0_35_0_real,
  output     [15:0]   io_coef_out_payload_0_35_0_imag,
  output     [15:0]   io_coef_out_payload_0_35_1_real,
  output     [15:0]   io_coef_out_payload_0_35_1_imag,
  output     [15:0]   io_coef_out_payload_0_35_2_real,
  output     [15:0]   io_coef_out_payload_0_35_2_imag,
  output     [15:0]   io_coef_out_payload_0_35_3_real,
  output     [15:0]   io_coef_out_payload_0_35_3_imag,
  output     [15:0]   io_coef_out_payload_0_35_4_real,
  output     [15:0]   io_coef_out_payload_0_35_4_imag,
  output     [15:0]   io_coef_out_payload_0_35_5_real,
  output     [15:0]   io_coef_out_payload_0_35_5_imag,
  output     [15:0]   io_coef_out_payload_0_35_6_real,
  output     [15:0]   io_coef_out_payload_0_35_6_imag,
  output     [15:0]   io_coef_out_payload_0_35_7_real,
  output     [15:0]   io_coef_out_payload_0_35_7_imag,
  output     [15:0]   io_coef_out_payload_0_35_8_real,
  output     [15:0]   io_coef_out_payload_0_35_8_imag,
  output     [15:0]   io_coef_out_payload_0_35_9_real,
  output     [15:0]   io_coef_out_payload_0_35_9_imag,
  output     [15:0]   io_coef_out_payload_0_35_10_real,
  output     [15:0]   io_coef_out_payload_0_35_10_imag,
  output     [15:0]   io_coef_out_payload_0_35_11_real,
  output     [15:0]   io_coef_out_payload_0_35_11_imag,
  output     [15:0]   io_coef_out_payload_0_35_12_real,
  output     [15:0]   io_coef_out_payload_0_35_12_imag,
  output     [15:0]   io_coef_out_payload_0_35_13_real,
  output     [15:0]   io_coef_out_payload_0_35_13_imag,
  output     [15:0]   io_coef_out_payload_0_35_14_real,
  output     [15:0]   io_coef_out_payload_0_35_14_imag,
  output     [15:0]   io_coef_out_payload_0_35_15_real,
  output     [15:0]   io_coef_out_payload_0_35_15_imag,
  output     [15:0]   io_coef_out_payload_0_35_16_real,
  output     [15:0]   io_coef_out_payload_0_35_16_imag,
  output     [15:0]   io_coef_out_payload_0_35_17_real,
  output     [15:0]   io_coef_out_payload_0_35_17_imag,
  output     [15:0]   io_coef_out_payload_0_35_18_real,
  output     [15:0]   io_coef_out_payload_0_35_18_imag,
  output     [15:0]   io_coef_out_payload_0_35_19_real,
  output     [15:0]   io_coef_out_payload_0_35_19_imag,
  output     [15:0]   io_coef_out_payload_0_35_20_real,
  output     [15:0]   io_coef_out_payload_0_35_20_imag,
  output     [15:0]   io_coef_out_payload_0_35_21_real,
  output     [15:0]   io_coef_out_payload_0_35_21_imag,
  output     [15:0]   io_coef_out_payload_0_35_22_real,
  output     [15:0]   io_coef_out_payload_0_35_22_imag,
  output     [15:0]   io_coef_out_payload_0_35_23_real,
  output     [15:0]   io_coef_out_payload_0_35_23_imag,
  output     [15:0]   io_coef_out_payload_0_35_24_real,
  output     [15:0]   io_coef_out_payload_0_35_24_imag,
  output     [15:0]   io_coef_out_payload_0_35_25_real,
  output     [15:0]   io_coef_out_payload_0_35_25_imag,
  output     [15:0]   io_coef_out_payload_0_35_26_real,
  output     [15:0]   io_coef_out_payload_0_35_26_imag,
  output     [15:0]   io_coef_out_payload_0_35_27_real,
  output     [15:0]   io_coef_out_payload_0_35_27_imag,
  output     [15:0]   io_coef_out_payload_0_35_28_real,
  output     [15:0]   io_coef_out_payload_0_35_28_imag,
  output     [15:0]   io_coef_out_payload_0_35_29_real,
  output     [15:0]   io_coef_out_payload_0_35_29_imag,
  output     [15:0]   io_coef_out_payload_0_35_30_real,
  output     [15:0]   io_coef_out_payload_0_35_30_imag,
  output     [15:0]   io_coef_out_payload_0_35_31_real,
  output     [15:0]   io_coef_out_payload_0_35_31_imag,
  output     [15:0]   io_coef_out_payload_0_35_32_real,
  output     [15:0]   io_coef_out_payload_0_35_32_imag,
  output     [15:0]   io_coef_out_payload_0_35_33_real,
  output     [15:0]   io_coef_out_payload_0_35_33_imag,
  output     [15:0]   io_coef_out_payload_0_35_34_real,
  output     [15:0]   io_coef_out_payload_0_35_34_imag,
  output     [15:0]   io_coef_out_payload_0_35_35_real,
  output     [15:0]   io_coef_out_payload_0_35_35_imag,
  output     [15:0]   io_coef_out_payload_0_35_36_real,
  output     [15:0]   io_coef_out_payload_0_35_36_imag,
  output     [15:0]   io_coef_out_payload_0_35_37_real,
  output     [15:0]   io_coef_out_payload_0_35_37_imag,
  output     [15:0]   io_coef_out_payload_0_35_38_real,
  output     [15:0]   io_coef_out_payload_0_35_38_imag,
  output     [15:0]   io_coef_out_payload_0_35_39_real,
  output     [15:0]   io_coef_out_payload_0_35_39_imag,
  output     [15:0]   io_coef_out_payload_0_35_40_real,
  output     [15:0]   io_coef_out_payload_0_35_40_imag,
  output     [15:0]   io_coef_out_payload_0_35_41_real,
  output     [15:0]   io_coef_out_payload_0_35_41_imag,
  output     [15:0]   io_coef_out_payload_0_35_42_real,
  output     [15:0]   io_coef_out_payload_0_35_42_imag,
  output     [15:0]   io_coef_out_payload_0_35_43_real,
  output     [15:0]   io_coef_out_payload_0_35_43_imag,
  output     [15:0]   io_coef_out_payload_0_35_44_real,
  output     [15:0]   io_coef_out_payload_0_35_44_imag,
  output     [15:0]   io_coef_out_payload_0_35_45_real,
  output     [15:0]   io_coef_out_payload_0_35_45_imag,
  output     [15:0]   io_coef_out_payload_0_35_46_real,
  output     [15:0]   io_coef_out_payload_0_35_46_imag,
  output     [15:0]   io_coef_out_payload_0_35_47_real,
  output     [15:0]   io_coef_out_payload_0_35_47_imag,
  output     [15:0]   io_coef_out_payload_0_35_48_real,
  output     [15:0]   io_coef_out_payload_0_35_48_imag,
  output     [15:0]   io_coef_out_payload_0_35_49_real,
  output     [15:0]   io_coef_out_payload_0_35_49_imag,
  output     [15:0]   io_coef_out_payload_0_36_0_real,
  output     [15:0]   io_coef_out_payload_0_36_0_imag,
  output     [15:0]   io_coef_out_payload_0_36_1_real,
  output     [15:0]   io_coef_out_payload_0_36_1_imag,
  output     [15:0]   io_coef_out_payload_0_36_2_real,
  output     [15:0]   io_coef_out_payload_0_36_2_imag,
  output     [15:0]   io_coef_out_payload_0_36_3_real,
  output     [15:0]   io_coef_out_payload_0_36_3_imag,
  output     [15:0]   io_coef_out_payload_0_36_4_real,
  output     [15:0]   io_coef_out_payload_0_36_4_imag,
  output     [15:0]   io_coef_out_payload_0_36_5_real,
  output     [15:0]   io_coef_out_payload_0_36_5_imag,
  output     [15:0]   io_coef_out_payload_0_36_6_real,
  output     [15:0]   io_coef_out_payload_0_36_6_imag,
  output     [15:0]   io_coef_out_payload_0_36_7_real,
  output     [15:0]   io_coef_out_payload_0_36_7_imag,
  output     [15:0]   io_coef_out_payload_0_36_8_real,
  output     [15:0]   io_coef_out_payload_0_36_8_imag,
  output     [15:0]   io_coef_out_payload_0_36_9_real,
  output     [15:0]   io_coef_out_payload_0_36_9_imag,
  output     [15:0]   io_coef_out_payload_0_36_10_real,
  output     [15:0]   io_coef_out_payload_0_36_10_imag,
  output     [15:0]   io_coef_out_payload_0_36_11_real,
  output     [15:0]   io_coef_out_payload_0_36_11_imag,
  output     [15:0]   io_coef_out_payload_0_36_12_real,
  output     [15:0]   io_coef_out_payload_0_36_12_imag,
  output     [15:0]   io_coef_out_payload_0_36_13_real,
  output     [15:0]   io_coef_out_payload_0_36_13_imag,
  output     [15:0]   io_coef_out_payload_0_36_14_real,
  output     [15:0]   io_coef_out_payload_0_36_14_imag,
  output     [15:0]   io_coef_out_payload_0_36_15_real,
  output     [15:0]   io_coef_out_payload_0_36_15_imag,
  output     [15:0]   io_coef_out_payload_0_36_16_real,
  output     [15:0]   io_coef_out_payload_0_36_16_imag,
  output     [15:0]   io_coef_out_payload_0_36_17_real,
  output     [15:0]   io_coef_out_payload_0_36_17_imag,
  output     [15:0]   io_coef_out_payload_0_36_18_real,
  output     [15:0]   io_coef_out_payload_0_36_18_imag,
  output     [15:0]   io_coef_out_payload_0_36_19_real,
  output     [15:0]   io_coef_out_payload_0_36_19_imag,
  output     [15:0]   io_coef_out_payload_0_36_20_real,
  output     [15:0]   io_coef_out_payload_0_36_20_imag,
  output     [15:0]   io_coef_out_payload_0_36_21_real,
  output     [15:0]   io_coef_out_payload_0_36_21_imag,
  output     [15:0]   io_coef_out_payload_0_36_22_real,
  output     [15:0]   io_coef_out_payload_0_36_22_imag,
  output     [15:0]   io_coef_out_payload_0_36_23_real,
  output     [15:0]   io_coef_out_payload_0_36_23_imag,
  output     [15:0]   io_coef_out_payload_0_36_24_real,
  output     [15:0]   io_coef_out_payload_0_36_24_imag,
  output     [15:0]   io_coef_out_payload_0_36_25_real,
  output     [15:0]   io_coef_out_payload_0_36_25_imag,
  output     [15:0]   io_coef_out_payload_0_36_26_real,
  output     [15:0]   io_coef_out_payload_0_36_26_imag,
  output     [15:0]   io_coef_out_payload_0_36_27_real,
  output     [15:0]   io_coef_out_payload_0_36_27_imag,
  output     [15:0]   io_coef_out_payload_0_36_28_real,
  output     [15:0]   io_coef_out_payload_0_36_28_imag,
  output     [15:0]   io_coef_out_payload_0_36_29_real,
  output     [15:0]   io_coef_out_payload_0_36_29_imag,
  output     [15:0]   io_coef_out_payload_0_36_30_real,
  output     [15:0]   io_coef_out_payload_0_36_30_imag,
  output     [15:0]   io_coef_out_payload_0_36_31_real,
  output     [15:0]   io_coef_out_payload_0_36_31_imag,
  output     [15:0]   io_coef_out_payload_0_36_32_real,
  output     [15:0]   io_coef_out_payload_0_36_32_imag,
  output     [15:0]   io_coef_out_payload_0_36_33_real,
  output     [15:0]   io_coef_out_payload_0_36_33_imag,
  output     [15:0]   io_coef_out_payload_0_36_34_real,
  output     [15:0]   io_coef_out_payload_0_36_34_imag,
  output     [15:0]   io_coef_out_payload_0_36_35_real,
  output     [15:0]   io_coef_out_payload_0_36_35_imag,
  output     [15:0]   io_coef_out_payload_0_36_36_real,
  output     [15:0]   io_coef_out_payload_0_36_36_imag,
  output     [15:0]   io_coef_out_payload_0_36_37_real,
  output     [15:0]   io_coef_out_payload_0_36_37_imag,
  output     [15:0]   io_coef_out_payload_0_36_38_real,
  output     [15:0]   io_coef_out_payload_0_36_38_imag,
  output     [15:0]   io_coef_out_payload_0_36_39_real,
  output     [15:0]   io_coef_out_payload_0_36_39_imag,
  output     [15:0]   io_coef_out_payload_0_36_40_real,
  output     [15:0]   io_coef_out_payload_0_36_40_imag,
  output     [15:0]   io_coef_out_payload_0_36_41_real,
  output     [15:0]   io_coef_out_payload_0_36_41_imag,
  output     [15:0]   io_coef_out_payload_0_36_42_real,
  output     [15:0]   io_coef_out_payload_0_36_42_imag,
  output     [15:0]   io_coef_out_payload_0_36_43_real,
  output     [15:0]   io_coef_out_payload_0_36_43_imag,
  output     [15:0]   io_coef_out_payload_0_36_44_real,
  output     [15:0]   io_coef_out_payload_0_36_44_imag,
  output     [15:0]   io_coef_out_payload_0_36_45_real,
  output     [15:0]   io_coef_out_payload_0_36_45_imag,
  output     [15:0]   io_coef_out_payload_0_36_46_real,
  output     [15:0]   io_coef_out_payload_0_36_46_imag,
  output     [15:0]   io_coef_out_payload_0_36_47_real,
  output     [15:0]   io_coef_out_payload_0_36_47_imag,
  output     [15:0]   io_coef_out_payload_0_36_48_real,
  output     [15:0]   io_coef_out_payload_0_36_48_imag,
  output     [15:0]   io_coef_out_payload_0_36_49_real,
  output     [15:0]   io_coef_out_payload_0_36_49_imag,
  output     [15:0]   io_coef_out_payload_0_37_0_real,
  output     [15:0]   io_coef_out_payload_0_37_0_imag,
  output     [15:0]   io_coef_out_payload_0_37_1_real,
  output     [15:0]   io_coef_out_payload_0_37_1_imag,
  output     [15:0]   io_coef_out_payload_0_37_2_real,
  output     [15:0]   io_coef_out_payload_0_37_2_imag,
  output     [15:0]   io_coef_out_payload_0_37_3_real,
  output     [15:0]   io_coef_out_payload_0_37_3_imag,
  output     [15:0]   io_coef_out_payload_0_37_4_real,
  output     [15:0]   io_coef_out_payload_0_37_4_imag,
  output     [15:0]   io_coef_out_payload_0_37_5_real,
  output     [15:0]   io_coef_out_payload_0_37_5_imag,
  output     [15:0]   io_coef_out_payload_0_37_6_real,
  output     [15:0]   io_coef_out_payload_0_37_6_imag,
  output     [15:0]   io_coef_out_payload_0_37_7_real,
  output     [15:0]   io_coef_out_payload_0_37_7_imag,
  output     [15:0]   io_coef_out_payload_0_37_8_real,
  output     [15:0]   io_coef_out_payload_0_37_8_imag,
  output     [15:0]   io_coef_out_payload_0_37_9_real,
  output     [15:0]   io_coef_out_payload_0_37_9_imag,
  output     [15:0]   io_coef_out_payload_0_37_10_real,
  output     [15:0]   io_coef_out_payload_0_37_10_imag,
  output     [15:0]   io_coef_out_payload_0_37_11_real,
  output     [15:0]   io_coef_out_payload_0_37_11_imag,
  output     [15:0]   io_coef_out_payload_0_37_12_real,
  output     [15:0]   io_coef_out_payload_0_37_12_imag,
  output     [15:0]   io_coef_out_payload_0_37_13_real,
  output     [15:0]   io_coef_out_payload_0_37_13_imag,
  output     [15:0]   io_coef_out_payload_0_37_14_real,
  output     [15:0]   io_coef_out_payload_0_37_14_imag,
  output     [15:0]   io_coef_out_payload_0_37_15_real,
  output     [15:0]   io_coef_out_payload_0_37_15_imag,
  output     [15:0]   io_coef_out_payload_0_37_16_real,
  output     [15:0]   io_coef_out_payload_0_37_16_imag,
  output     [15:0]   io_coef_out_payload_0_37_17_real,
  output     [15:0]   io_coef_out_payload_0_37_17_imag,
  output     [15:0]   io_coef_out_payload_0_37_18_real,
  output     [15:0]   io_coef_out_payload_0_37_18_imag,
  output     [15:0]   io_coef_out_payload_0_37_19_real,
  output     [15:0]   io_coef_out_payload_0_37_19_imag,
  output     [15:0]   io_coef_out_payload_0_37_20_real,
  output     [15:0]   io_coef_out_payload_0_37_20_imag,
  output     [15:0]   io_coef_out_payload_0_37_21_real,
  output     [15:0]   io_coef_out_payload_0_37_21_imag,
  output     [15:0]   io_coef_out_payload_0_37_22_real,
  output     [15:0]   io_coef_out_payload_0_37_22_imag,
  output     [15:0]   io_coef_out_payload_0_37_23_real,
  output     [15:0]   io_coef_out_payload_0_37_23_imag,
  output     [15:0]   io_coef_out_payload_0_37_24_real,
  output     [15:0]   io_coef_out_payload_0_37_24_imag,
  output     [15:0]   io_coef_out_payload_0_37_25_real,
  output     [15:0]   io_coef_out_payload_0_37_25_imag,
  output     [15:0]   io_coef_out_payload_0_37_26_real,
  output     [15:0]   io_coef_out_payload_0_37_26_imag,
  output     [15:0]   io_coef_out_payload_0_37_27_real,
  output     [15:0]   io_coef_out_payload_0_37_27_imag,
  output     [15:0]   io_coef_out_payload_0_37_28_real,
  output     [15:0]   io_coef_out_payload_0_37_28_imag,
  output     [15:0]   io_coef_out_payload_0_37_29_real,
  output     [15:0]   io_coef_out_payload_0_37_29_imag,
  output     [15:0]   io_coef_out_payload_0_37_30_real,
  output     [15:0]   io_coef_out_payload_0_37_30_imag,
  output     [15:0]   io_coef_out_payload_0_37_31_real,
  output     [15:0]   io_coef_out_payload_0_37_31_imag,
  output     [15:0]   io_coef_out_payload_0_37_32_real,
  output     [15:0]   io_coef_out_payload_0_37_32_imag,
  output     [15:0]   io_coef_out_payload_0_37_33_real,
  output     [15:0]   io_coef_out_payload_0_37_33_imag,
  output     [15:0]   io_coef_out_payload_0_37_34_real,
  output     [15:0]   io_coef_out_payload_0_37_34_imag,
  output     [15:0]   io_coef_out_payload_0_37_35_real,
  output     [15:0]   io_coef_out_payload_0_37_35_imag,
  output     [15:0]   io_coef_out_payload_0_37_36_real,
  output     [15:0]   io_coef_out_payload_0_37_36_imag,
  output     [15:0]   io_coef_out_payload_0_37_37_real,
  output     [15:0]   io_coef_out_payload_0_37_37_imag,
  output     [15:0]   io_coef_out_payload_0_37_38_real,
  output     [15:0]   io_coef_out_payload_0_37_38_imag,
  output     [15:0]   io_coef_out_payload_0_37_39_real,
  output     [15:0]   io_coef_out_payload_0_37_39_imag,
  output     [15:0]   io_coef_out_payload_0_37_40_real,
  output     [15:0]   io_coef_out_payload_0_37_40_imag,
  output     [15:0]   io_coef_out_payload_0_37_41_real,
  output     [15:0]   io_coef_out_payload_0_37_41_imag,
  output     [15:0]   io_coef_out_payload_0_37_42_real,
  output     [15:0]   io_coef_out_payload_0_37_42_imag,
  output     [15:0]   io_coef_out_payload_0_37_43_real,
  output     [15:0]   io_coef_out_payload_0_37_43_imag,
  output     [15:0]   io_coef_out_payload_0_37_44_real,
  output     [15:0]   io_coef_out_payload_0_37_44_imag,
  output     [15:0]   io_coef_out_payload_0_37_45_real,
  output     [15:0]   io_coef_out_payload_0_37_45_imag,
  output     [15:0]   io_coef_out_payload_0_37_46_real,
  output     [15:0]   io_coef_out_payload_0_37_46_imag,
  output     [15:0]   io_coef_out_payload_0_37_47_real,
  output     [15:0]   io_coef_out_payload_0_37_47_imag,
  output     [15:0]   io_coef_out_payload_0_37_48_real,
  output     [15:0]   io_coef_out_payload_0_37_48_imag,
  output     [15:0]   io_coef_out_payload_0_37_49_real,
  output     [15:0]   io_coef_out_payload_0_37_49_imag,
  output     [15:0]   io_coef_out_payload_0_38_0_real,
  output     [15:0]   io_coef_out_payload_0_38_0_imag,
  output     [15:0]   io_coef_out_payload_0_38_1_real,
  output     [15:0]   io_coef_out_payload_0_38_1_imag,
  output     [15:0]   io_coef_out_payload_0_38_2_real,
  output     [15:0]   io_coef_out_payload_0_38_2_imag,
  output     [15:0]   io_coef_out_payload_0_38_3_real,
  output     [15:0]   io_coef_out_payload_0_38_3_imag,
  output     [15:0]   io_coef_out_payload_0_38_4_real,
  output     [15:0]   io_coef_out_payload_0_38_4_imag,
  output     [15:0]   io_coef_out_payload_0_38_5_real,
  output     [15:0]   io_coef_out_payload_0_38_5_imag,
  output     [15:0]   io_coef_out_payload_0_38_6_real,
  output     [15:0]   io_coef_out_payload_0_38_6_imag,
  output     [15:0]   io_coef_out_payload_0_38_7_real,
  output     [15:0]   io_coef_out_payload_0_38_7_imag,
  output     [15:0]   io_coef_out_payload_0_38_8_real,
  output     [15:0]   io_coef_out_payload_0_38_8_imag,
  output     [15:0]   io_coef_out_payload_0_38_9_real,
  output     [15:0]   io_coef_out_payload_0_38_9_imag,
  output     [15:0]   io_coef_out_payload_0_38_10_real,
  output     [15:0]   io_coef_out_payload_0_38_10_imag,
  output     [15:0]   io_coef_out_payload_0_38_11_real,
  output     [15:0]   io_coef_out_payload_0_38_11_imag,
  output     [15:0]   io_coef_out_payload_0_38_12_real,
  output     [15:0]   io_coef_out_payload_0_38_12_imag,
  output     [15:0]   io_coef_out_payload_0_38_13_real,
  output     [15:0]   io_coef_out_payload_0_38_13_imag,
  output     [15:0]   io_coef_out_payload_0_38_14_real,
  output     [15:0]   io_coef_out_payload_0_38_14_imag,
  output     [15:0]   io_coef_out_payload_0_38_15_real,
  output     [15:0]   io_coef_out_payload_0_38_15_imag,
  output     [15:0]   io_coef_out_payload_0_38_16_real,
  output     [15:0]   io_coef_out_payload_0_38_16_imag,
  output     [15:0]   io_coef_out_payload_0_38_17_real,
  output     [15:0]   io_coef_out_payload_0_38_17_imag,
  output     [15:0]   io_coef_out_payload_0_38_18_real,
  output     [15:0]   io_coef_out_payload_0_38_18_imag,
  output     [15:0]   io_coef_out_payload_0_38_19_real,
  output     [15:0]   io_coef_out_payload_0_38_19_imag,
  output     [15:0]   io_coef_out_payload_0_38_20_real,
  output     [15:0]   io_coef_out_payload_0_38_20_imag,
  output     [15:0]   io_coef_out_payload_0_38_21_real,
  output     [15:0]   io_coef_out_payload_0_38_21_imag,
  output     [15:0]   io_coef_out_payload_0_38_22_real,
  output     [15:0]   io_coef_out_payload_0_38_22_imag,
  output     [15:0]   io_coef_out_payload_0_38_23_real,
  output     [15:0]   io_coef_out_payload_0_38_23_imag,
  output     [15:0]   io_coef_out_payload_0_38_24_real,
  output     [15:0]   io_coef_out_payload_0_38_24_imag,
  output     [15:0]   io_coef_out_payload_0_38_25_real,
  output     [15:0]   io_coef_out_payload_0_38_25_imag,
  output     [15:0]   io_coef_out_payload_0_38_26_real,
  output     [15:0]   io_coef_out_payload_0_38_26_imag,
  output     [15:0]   io_coef_out_payload_0_38_27_real,
  output     [15:0]   io_coef_out_payload_0_38_27_imag,
  output     [15:0]   io_coef_out_payload_0_38_28_real,
  output     [15:0]   io_coef_out_payload_0_38_28_imag,
  output     [15:0]   io_coef_out_payload_0_38_29_real,
  output     [15:0]   io_coef_out_payload_0_38_29_imag,
  output     [15:0]   io_coef_out_payload_0_38_30_real,
  output     [15:0]   io_coef_out_payload_0_38_30_imag,
  output     [15:0]   io_coef_out_payload_0_38_31_real,
  output     [15:0]   io_coef_out_payload_0_38_31_imag,
  output     [15:0]   io_coef_out_payload_0_38_32_real,
  output     [15:0]   io_coef_out_payload_0_38_32_imag,
  output     [15:0]   io_coef_out_payload_0_38_33_real,
  output     [15:0]   io_coef_out_payload_0_38_33_imag,
  output     [15:0]   io_coef_out_payload_0_38_34_real,
  output     [15:0]   io_coef_out_payload_0_38_34_imag,
  output     [15:0]   io_coef_out_payload_0_38_35_real,
  output     [15:0]   io_coef_out_payload_0_38_35_imag,
  output     [15:0]   io_coef_out_payload_0_38_36_real,
  output     [15:0]   io_coef_out_payload_0_38_36_imag,
  output     [15:0]   io_coef_out_payload_0_38_37_real,
  output     [15:0]   io_coef_out_payload_0_38_37_imag,
  output     [15:0]   io_coef_out_payload_0_38_38_real,
  output     [15:0]   io_coef_out_payload_0_38_38_imag,
  output     [15:0]   io_coef_out_payload_0_38_39_real,
  output     [15:0]   io_coef_out_payload_0_38_39_imag,
  output     [15:0]   io_coef_out_payload_0_38_40_real,
  output     [15:0]   io_coef_out_payload_0_38_40_imag,
  output     [15:0]   io_coef_out_payload_0_38_41_real,
  output     [15:0]   io_coef_out_payload_0_38_41_imag,
  output     [15:0]   io_coef_out_payload_0_38_42_real,
  output     [15:0]   io_coef_out_payload_0_38_42_imag,
  output     [15:0]   io_coef_out_payload_0_38_43_real,
  output     [15:0]   io_coef_out_payload_0_38_43_imag,
  output     [15:0]   io_coef_out_payload_0_38_44_real,
  output     [15:0]   io_coef_out_payload_0_38_44_imag,
  output     [15:0]   io_coef_out_payload_0_38_45_real,
  output     [15:0]   io_coef_out_payload_0_38_45_imag,
  output     [15:0]   io_coef_out_payload_0_38_46_real,
  output     [15:0]   io_coef_out_payload_0_38_46_imag,
  output     [15:0]   io_coef_out_payload_0_38_47_real,
  output     [15:0]   io_coef_out_payload_0_38_47_imag,
  output     [15:0]   io_coef_out_payload_0_38_48_real,
  output     [15:0]   io_coef_out_payload_0_38_48_imag,
  output     [15:0]   io_coef_out_payload_0_38_49_real,
  output     [15:0]   io_coef_out_payload_0_38_49_imag,
  output     [15:0]   io_coef_out_payload_0_39_0_real,
  output     [15:0]   io_coef_out_payload_0_39_0_imag,
  output     [15:0]   io_coef_out_payload_0_39_1_real,
  output     [15:0]   io_coef_out_payload_0_39_1_imag,
  output     [15:0]   io_coef_out_payload_0_39_2_real,
  output     [15:0]   io_coef_out_payload_0_39_2_imag,
  output     [15:0]   io_coef_out_payload_0_39_3_real,
  output     [15:0]   io_coef_out_payload_0_39_3_imag,
  output     [15:0]   io_coef_out_payload_0_39_4_real,
  output     [15:0]   io_coef_out_payload_0_39_4_imag,
  output     [15:0]   io_coef_out_payload_0_39_5_real,
  output     [15:0]   io_coef_out_payload_0_39_5_imag,
  output     [15:0]   io_coef_out_payload_0_39_6_real,
  output     [15:0]   io_coef_out_payload_0_39_6_imag,
  output     [15:0]   io_coef_out_payload_0_39_7_real,
  output     [15:0]   io_coef_out_payload_0_39_7_imag,
  output     [15:0]   io_coef_out_payload_0_39_8_real,
  output     [15:0]   io_coef_out_payload_0_39_8_imag,
  output     [15:0]   io_coef_out_payload_0_39_9_real,
  output     [15:0]   io_coef_out_payload_0_39_9_imag,
  output     [15:0]   io_coef_out_payload_0_39_10_real,
  output     [15:0]   io_coef_out_payload_0_39_10_imag,
  output     [15:0]   io_coef_out_payload_0_39_11_real,
  output     [15:0]   io_coef_out_payload_0_39_11_imag,
  output     [15:0]   io_coef_out_payload_0_39_12_real,
  output     [15:0]   io_coef_out_payload_0_39_12_imag,
  output     [15:0]   io_coef_out_payload_0_39_13_real,
  output     [15:0]   io_coef_out_payload_0_39_13_imag,
  output     [15:0]   io_coef_out_payload_0_39_14_real,
  output     [15:0]   io_coef_out_payload_0_39_14_imag,
  output     [15:0]   io_coef_out_payload_0_39_15_real,
  output     [15:0]   io_coef_out_payload_0_39_15_imag,
  output     [15:0]   io_coef_out_payload_0_39_16_real,
  output     [15:0]   io_coef_out_payload_0_39_16_imag,
  output     [15:0]   io_coef_out_payload_0_39_17_real,
  output     [15:0]   io_coef_out_payload_0_39_17_imag,
  output     [15:0]   io_coef_out_payload_0_39_18_real,
  output     [15:0]   io_coef_out_payload_0_39_18_imag,
  output     [15:0]   io_coef_out_payload_0_39_19_real,
  output     [15:0]   io_coef_out_payload_0_39_19_imag,
  output     [15:0]   io_coef_out_payload_0_39_20_real,
  output     [15:0]   io_coef_out_payload_0_39_20_imag,
  output     [15:0]   io_coef_out_payload_0_39_21_real,
  output     [15:0]   io_coef_out_payload_0_39_21_imag,
  output     [15:0]   io_coef_out_payload_0_39_22_real,
  output     [15:0]   io_coef_out_payload_0_39_22_imag,
  output     [15:0]   io_coef_out_payload_0_39_23_real,
  output     [15:0]   io_coef_out_payload_0_39_23_imag,
  output     [15:0]   io_coef_out_payload_0_39_24_real,
  output     [15:0]   io_coef_out_payload_0_39_24_imag,
  output     [15:0]   io_coef_out_payload_0_39_25_real,
  output     [15:0]   io_coef_out_payload_0_39_25_imag,
  output     [15:0]   io_coef_out_payload_0_39_26_real,
  output     [15:0]   io_coef_out_payload_0_39_26_imag,
  output     [15:0]   io_coef_out_payload_0_39_27_real,
  output     [15:0]   io_coef_out_payload_0_39_27_imag,
  output     [15:0]   io_coef_out_payload_0_39_28_real,
  output     [15:0]   io_coef_out_payload_0_39_28_imag,
  output     [15:0]   io_coef_out_payload_0_39_29_real,
  output     [15:0]   io_coef_out_payload_0_39_29_imag,
  output     [15:0]   io_coef_out_payload_0_39_30_real,
  output     [15:0]   io_coef_out_payload_0_39_30_imag,
  output     [15:0]   io_coef_out_payload_0_39_31_real,
  output     [15:0]   io_coef_out_payload_0_39_31_imag,
  output     [15:0]   io_coef_out_payload_0_39_32_real,
  output     [15:0]   io_coef_out_payload_0_39_32_imag,
  output     [15:0]   io_coef_out_payload_0_39_33_real,
  output     [15:0]   io_coef_out_payload_0_39_33_imag,
  output     [15:0]   io_coef_out_payload_0_39_34_real,
  output     [15:0]   io_coef_out_payload_0_39_34_imag,
  output     [15:0]   io_coef_out_payload_0_39_35_real,
  output     [15:0]   io_coef_out_payload_0_39_35_imag,
  output     [15:0]   io_coef_out_payload_0_39_36_real,
  output     [15:0]   io_coef_out_payload_0_39_36_imag,
  output     [15:0]   io_coef_out_payload_0_39_37_real,
  output     [15:0]   io_coef_out_payload_0_39_37_imag,
  output     [15:0]   io_coef_out_payload_0_39_38_real,
  output     [15:0]   io_coef_out_payload_0_39_38_imag,
  output     [15:0]   io_coef_out_payload_0_39_39_real,
  output     [15:0]   io_coef_out_payload_0_39_39_imag,
  output     [15:0]   io_coef_out_payload_0_39_40_real,
  output     [15:0]   io_coef_out_payload_0_39_40_imag,
  output     [15:0]   io_coef_out_payload_0_39_41_real,
  output     [15:0]   io_coef_out_payload_0_39_41_imag,
  output     [15:0]   io_coef_out_payload_0_39_42_real,
  output     [15:0]   io_coef_out_payload_0_39_42_imag,
  output     [15:0]   io_coef_out_payload_0_39_43_real,
  output     [15:0]   io_coef_out_payload_0_39_43_imag,
  output     [15:0]   io_coef_out_payload_0_39_44_real,
  output     [15:0]   io_coef_out_payload_0_39_44_imag,
  output     [15:0]   io_coef_out_payload_0_39_45_real,
  output     [15:0]   io_coef_out_payload_0_39_45_imag,
  output     [15:0]   io_coef_out_payload_0_39_46_real,
  output     [15:0]   io_coef_out_payload_0_39_46_imag,
  output     [15:0]   io_coef_out_payload_0_39_47_real,
  output     [15:0]   io_coef_out_payload_0_39_47_imag,
  output     [15:0]   io_coef_out_payload_0_39_48_real,
  output     [15:0]   io_coef_out_payload_0_39_48_imag,
  output     [15:0]   io_coef_out_payload_0_39_49_real,
  output     [15:0]   io_coef_out_payload_0_39_49_imag,
  output     [15:0]   io_coef_out_payload_0_40_0_real,
  output     [15:0]   io_coef_out_payload_0_40_0_imag,
  output     [15:0]   io_coef_out_payload_0_40_1_real,
  output     [15:0]   io_coef_out_payload_0_40_1_imag,
  output     [15:0]   io_coef_out_payload_0_40_2_real,
  output     [15:0]   io_coef_out_payload_0_40_2_imag,
  output     [15:0]   io_coef_out_payload_0_40_3_real,
  output     [15:0]   io_coef_out_payload_0_40_3_imag,
  output     [15:0]   io_coef_out_payload_0_40_4_real,
  output     [15:0]   io_coef_out_payload_0_40_4_imag,
  output     [15:0]   io_coef_out_payload_0_40_5_real,
  output     [15:0]   io_coef_out_payload_0_40_5_imag,
  output     [15:0]   io_coef_out_payload_0_40_6_real,
  output     [15:0]   io_coef_out_payload_0_40_6_imag,
  output     [15:0]   io_coef_out_payload_0_40_7_real,
  output     [15:0]   io_coef_out_payload_0_40_7_imag,
  output     [15:0]   io_coef_out_payload_0_40_8_real,
  output     [15:0]   io_coef_out_payload_0_40_8_imag,
  output     [15:0]   io_coef_out_payload_0_40_9_real,
  output     [15:0]   io_coef_out_payload_0_40_9_imag,
  output     [15:0]   io_coef_out_payload_0_40_10_real,
  output     [15:0]   io_coef_out_payload_0_40_10_imag,
  output     [15:0]   io_coef_out_payload_0_40_11_real,
  output     [15:0]   io_coef_out_payload_0_40_11_imag,
  output     [15:0]   io_coef_out_payload_0_40_12_real,
  output     [15:0]   io_coef_out_payload_0_40_12_imag,
  output     [15:0]   io_coef_out_payload_0_40_13_real,
  output     [15:0]   io_coef_out_payload_0_40_13_imag,
  output     [15:0]   io_coef_out_payload_0_40_14_real,
  output     [15:0]   io_coef_out_payload_0_40_14_imag,
  output     [15:0]   io_coef_out_payload_0_40_15_real,
  output     [15:0]   io_coef_out_payload_0_40_15_imag,
  output     [15:0]   io_coef_out_payload_0_40_16_real,
  output     [15:0]   io_coef_out_payload_0_40_16_imag,
  output     [15:0]   io_coef_out_payload_0_40_17_real,
  output     [15:0]   io_coef_out_payload_0_40_17_imag,
  output     [15:0]   io_coef_out_payload_0_40_18_real,
  output     [15:0]   io_coef_out_payload_0_40_18_imag,
  output     [15:0]   io_coef_out_payload_0_40_19_real,
  output     [15:0]   io_coef_out_payload_0_40_19_imag,
  output     [15:0]   io_coef_out_payload_0_40_20_real,
  output     [15:0]   io_coef_out_payload_0_40_20_imag,
  output     [15:0]   io_coef_out_payload_0_40_21_real,
  output     [15:0]   io_coef_out_payload_0_40_21_imag,
  output     [15:0]   io_coef_out_payload_0_40_22_real,
  output     [15:0]   io_coef_out_payload_0_40_22_imag,
  output     [15:0]   io_coef_out_payload_0_40_23_real,
  output     [15:0]   io_coef_out_payload_0_40_23_imag,
  output     [15:0]   io_coef_out_payload_0_40_24_real,
  output     [15:0]   io_coef_out_payload_0_40_24_imag,
  output     [15:0]   io_coef_out_payload_0_40_25_real,
  output     [15:0]   io_coef_out_payload_0_40_25_imag,
  output     [15:0]   io_coef_out_payload_0_40_26_real,
  output     [15:0]   io_coef_out_payload_0_40_26_imag,
  output     [15:0]   io_coef_out_payload_0_40_27_real,
  output     [15:0]   io_coef_out_payload_0_40_27_imag,
  output     [15:0]   io_coef_out_payload_0_40_28_real,
  output     [15:0]   io_coef_out_payload_0_40_28_imag,
  output     [15:0]   io_coef_out_payload_0_40_29_real,
  output     [15:0]   io_coef_out_payload_0_40_29_imag,
  output     [15:0]   io_coef_out_payload_0_40_30_real,
  output     [15:0]   io_coef_out_payload_0_40_30_imag,
  output     [15:0]   io_coef_out_payload_0_40_31_real,
  output     [15:0]   io_coef_out_payload_0_40_31_imag,
  output     [15:0]   io_coef_out_payload_0_40_32_real,
  output     [15:0]   io_coef_out_payload_0_40_32_imag,
  output     [15:0]   io_coef_out_payload_0_40_33_real,
  output     [15:0]   io_coef_out_payload_0_40_33_imag,
  output     [15:0]   io_coef_out_payload_0_40_34_real,
  output     [15:0]   io_coef_out_payload_0_40_34_imag,
  output     [15:0]   io_coef_out_payload_0_40_35_real,
  output     [15:0]   io_coef_out_payload_0_40_35_imag,
  output     [15:0]   io_coef_out_payload_0_40_36_real,
  output     [15:0]   io_coef_out_payload_0_40_36_imag,
  output     [15:0]   io_coef_out_payload_0_40_37_real,
  output     [15:0]   io_coef_out_payload_0_40_37_imag,
  output     [15:0]   io_coef_out_payload_0_40_38_real,
  output     [15:0]   io_coef_out_payload_0_40_38_imag,
  output     [15:0]   io_coef_out_payload_0_40_39_real,
  output     [15:0]   io_coef_out_payload_0_40_39_imag,
  output     [15:0]   io_coef_out_payload_0_40_40_real,
  output     [15:0]   io_coef_out_payload_0_40_40_imag,
  output     [15:0]   io_coef_out_payload_0_40_41_real,
  output     [15:0]   io_coef_out_payload_0_40_41_imag,
  output     [15:0]   io_coef_out_payload_0_40_42_real,
  output     [15:0]   io_coef_out_payload_0_40_42_imag,
  output     [15:0]   io_coef_out_payload_0_40_43_real,
  output     [15:0]   io_coef_out_payload_0_40_43_imag,
  output     [15:0]   io_coef_out_payload_0_40_44_real,
  output     [15:0]   io_coef_out_payload_0_40_44_imag,
  output     [15:0]   io_coef_out_payload_0_40_45_real,
  output     [15:0]   io_coef_out_payload_0_40_45_imag,
  output     [15:0]   io_coef_out_payload_0_40_46_real,
  output     [15:0]   io_coef_out_payload_0_40_46_imag,
  output     [15:0]   io_coef_out_payload_0_40_47_real,
  output     [15:0]   io_coef_out_payload_0_40_47_imag,
  output     [15:0]   io_coef_out_payload_0_40_48_real,
  output     [15:0]   io_coef_out_payload_0_40_48_imag,
  output     [15:0]   io_coef_out_payload_0_40_49_real,
  output     [15:0]   io_coef_out_payload_0_40_49_imag,
  output     [15:0]   io_coef_out_payload_0_41_0_real,
  output     [15:0]   io_coef_out_payload_0_41_0_imag,
  output     [15:0]   io_coef_out_payload_0_41_1_real,
  output     [15:0]   io_coef_out_payload_0_41_1_imag,
  output     [15:0]   io_coef_out_payload_0_41_2_real,
  output     [15:0]   io_coef_out_payload_0_41_2_imag,
  output     [15:0]   io_coef_out_payload_0_41_3_real,
  output     [15:0]   io_coef_out_payload_0_41_3_imag,
  output     [15:0]   io_coef_out_payload_0_41_4_real,
  output     [15:0]   io_coef_out_payload_0_41_4_imag,
  output     [15:0]   io_coef_out_payload_0_41_5_real,
  output     [15:0]   io_coef_out_payload_0_41_5_imag,
  output     [15:0]   io_coef_out_payload_0_41_6_real,
  output     [15:0]   io_coef_out_payload_0_41_6_imag,
  output     [15:0]   io_coef_out_payload_0_41_7_real,
  output     [15:0]   io_coef_out_payload_0_41_7_imag,
  output     [15:0]   io_coef_out_payload_0_41_8_real,
  output     [15:0]   io_coef_out_payload_0_41_8_imag,
  output     [15:0]   io_coef_out_payload_0_41_9_real,
  output     [15:0]   io_coef_out_payload_0_41_9_imag,
  output     [15:0]   io_coef_out_payload_0_41_10_real,
  output     [15:0]   io_coef_out_payload_0_41_10_imag,
  output     [15:0]   io_coef_out_payload_0_41_11_real,
  output     [15:0]   io_coef_out_payload_0_41_11_imag,
  output     [15:0]   io_coef_out_payload_0_41_12_real,
  output     [15:0]   io_coef_out_payload_0_41_12_imag,
  output     [15:0]   io_coef_out_payload_0_41_13_real,
  output     [15:0]   io_coef_out_payload_0_41_13_imag,
  output     [15:0]   io_coef_out_payload_0_41_14_real,
  output     [15:0]   io_coef_out_payload_0_41_14_imag,
  output     [15:0]   io_coef_out_payload_0_41_15_real,
  output     [15:0]   io_coef_out_payload_0_41_15_imag,
  output     [15:0]   io_coef_out_payload_0_41_16_real,
  output     [15:0]   io_coef_out_payload_0_41_16_imag,
  output     [15:0]   io_coef_out_payload_0_41_17_real,
  output     [15:0]   io_coef_out_payload_0_41_17_imag,
  output     [15:0]   io_coef_out_payload_0_41_18_real,
  output     [15:0]   io_coef_out_payload_0_41_18_imag,
  output     [15:0]   io_coef_out_payload_0_41_19_real,
  output     [15:0]   io_coef_out_payload_0_41_19_imag,
  output     [15:0]   io_coef_out_payload_0_41_20_real,
  output     [15:0]   io_coef_out_payload_0_41_20_imag,
  output     [15:0]   io_coef_out_payload_0_41_21_real,
  output     [15:0]   io_coef_out_payload_0_41_21_imag,
  output     [15:0]   io_coef_out_payload_0_41_22_real,
  output     [15:0]   io_coef_out_payload_0_41_22_imag,
  output     [15:0]   io_coef_out_payload_0_41_23_real,
  output     [15:0]   io_coef_out_payload_0_41_23_imag,
  output     [15:0]   io_coef_out_payload_0_41_24_real,
  output     [15:0]   io_coef_out_payload_0_41_24_imag,
  output     [15:0]   io_coef_out_payload_0_41_25_real,
  output     [15:0]   io_coef_out_payload_0_41_25_imag,
  output     [15:0]   io_coef_out_payload_0_41_26_real,
  output     [15:0]   io_coef_out_payload_0_41_26_imag,
  output     [15:0]   io_coef_out_payload_0_41_27_real,
  output     [15:0]   io_coef_out_payload_0_41_27_imag,
  output     [15:0]   io_coef_out_payload_0_41_28_real,
  output     [15:0]   io_coef_out_payload_0_41_28_imag,
  output     [15:0]   io_coef_out_payload_0_41_29_real,
  output     [15:0]   io_coef_out_payload_0_41_29_imag,
  output     [15:0]   io_coef_out_payload_0_41_30_real,
  output     [15:0]   io_coef_out_payload_0_41_30_imag,
  output     [15:0]   io_coef_out_payload_0_41_31_real,
  output     [15:0]   io_coef_out_payload_0_41_31_imag,
  output     [15:0]   io_coef_out_payload_0_41_32_real,
  output     [15:0]   io_coef_out_payload_0_41_32_imag,
  output     [15:0]   io_coef_out_payload_0_41_33_real,
  output     [15:0]   io_coef_out_payload_0_41_33_imag,
  output     [15:0]   io_coef_out_payload_0_41_34_real,
  output     [15:0]   io_coef_out_payload_0_41_34_imag,
  output     [15:0]   io_coef_out_payload_0_41_35_real,
  output     [15:0]   io_coef_out_payload_0_41_35_imag,
  output     [15:0]   io_coef_out_payload_0_41_36_real,
  output     [15:0]   io_coef_out_payload_0_41_36_imag,
  output     [15:0]   io_coef_out_payload_0_41_37_real,
  output     [15:0]   io_coef_out_payload_0_41_37_imag,
  output     [15:0]   io_coef_out_payload_0_41_38_real,
  output     [15:0]   io_coef_out_payload_0_41_38_imag,
  output     [15:0]   io_coef_out_payload_0_41_39_real,
  output     [15:0]   io_coef_out_payload_0_41_39_imag,
  output     [15:0]   io_coef_out_payload_0_41_40_real,
  output     [15:0]   io_coef_out_payload_0_41_40_imag,
  output     [15:0]   io_coef_out_payload_0_41_41_real,
  output     [15:0]   io_coef_out_payload_0_41_41_imag,
  output     [15:0]   io_coef_out_payload_0_41_42_real,
  output     [15:0]   io_coef_out_payload_0_41_42_imag,
  output     [15:0]   io_coef_out_payload_0_41_43_real,
  output     [15:0]   io_coef_out_payload_0_41_43_imag,
  output     [15:0]   io_coef_out_payload_0_41_44_real,
  output     [15:0]   io_coef_out_payload_0_41_44_imag,
  output     [15:0]   io_coef_out_payload_0_41_45_real,
  output     [15:0]   io_coef_out_payload_0_41_45_imag,
  output     [15:0]   io_coef_out_payload_0_41_46_real,
  output     [15:0]   io_coef_out_payload_0_41_46_imag,
  output     [15:0]   io_coef_out_payload_0_41_47_real,
  output     [15:0]   io_coef_out_payload_0_41_47_imag,
  output     [15:0]   io_coef_out_payload_0_41_48_real,
  output     [15:0]   io_coef_out_payload_0_41_48_imag,
  output     [15:0]   io_coef_out_payload_0_41_49_real,
  output     [15:0]   io_coef_out_payload_0_41_49_imag,
  output     [15:0]   io_coef_out_payload_0_42_0_real,
  output     [15:0]   io_coef_out_payload_0_42_0_imag,
  output     [15:0]   io_coef_out_payload_0_42_1_real,
  output     [15:0]   io_coef_out_payload_0_42_1_imag,
  output     [15:0]   io_coef_out_payload_0_42_2_real,
  output     [15:0]   io_coef_out_payload_0_42_2_imag,
  output     [15:0]   io_coef_out_payload_0_42_3_real,
  output     [15:0]   io_coef_out_payload_0_42_3_imag,
  output     [15:0]   io_coef_out_payload_0_42_4_real,
  output     [15:0]   io_coef_out_payload_0_42_4_imag,
  output     [15:0]   io_coef_out_payload_0_42_5_real,
  output     [15:0]   io_coef_out_payload_0_42_5_imag,
  output     [15:0]   io_coef_out_payload_0_42_6_real,
  output     [15:0]   io_coef_out_payload_0_42_6_imag,
  output     [15:0]   io_coef_out_payload_0_42_7_real,
  output     [15:0]   io_coef_out_payload_0_42_7_imag,
  output     [15:0]   io_coef_out_payload_0_42_8_real,
  output     [15:0]   io_coef_out_payload_0_42_8_imag,
  output     [15:0]   io_coef_out_payload_0_42_9_real,
  output     [15:0]   io_coef_out_payload_0_42_9_imag,
  output     [15:0]   io_coef_out_payload_0_42_10_real,
  output     [15:0]   io_coef_out_payload_0_42_10_imag,
  output     [15:0]   io_coef_out_payload_0_42_11_real,
  output     [15:0]   io_coef_out_payload_0_42_11_imag,
  output     [15:0]   io_coef_out_payload_0_42_12_real,
  output     [15:0]   io_coef_out_payload_0_42_12_imag,
  output     [15:0]   io_coef_out_payload_0_42_13_real,
  output     [15:0]   io_coef_out_payload_0_42_13_imag,
  output     [15:0]   io_coef_out_payload_0_42_14_real,
  output     [15:0]   io_coef_out_payload_0_42_14_imag,
  output     [15:0]   io_coef_out_payload_0_42_15_real,
  output     [15:0]   io_coef_out_payload_0_42_15_imag,
  output     [15:0]   io_coef_out_payload_0_42_16_real,
  output     [15:0]   io_coef_out_payload_0_42_16_imag,
  output     [15:0]   io_coef_out_payload_0_42_17_real,
  output     [15:0]   io_coef_out_payload_0_42_17_imag,
  output     [15:0]   io_coef_out_payload_0_42_18_real,
  output     [15:0]   io_coef_out_payload_0_42_18_imag,
  output     [15:0]   io_coef_out_payload_0_42_19_real,
  output     [15:0]   io_coef_out_payload_0_42_19_imag,
  output     [15:0]   io_coef_out_payload_0_42_20_real,
  output     [15:0]   io_coef_out_payload_0_42_20_imag,
  output     [15:0]   io_coef_out_payload_0_42_21_real,
  output     [15:0]   io_coef_out_payload_0_42_21_imag,
  output     [15:0]   io_coef_out_payload_0_42_22_real,
  output     [15:0]   io_coef_out_payload_0_42_22_imag,
  output     [15:0]   io_coef_out_payload_0_42_23_real,
  output     [15:0]   io_coef_out_payload_0_42_23_imag,
  output     [15:0]   io_coef_out_payload_0_42_24_real,
  output     [15:0]   io_coef_out_payload_0_42_24_imag,
  output     [15:0]   io_coef_out_payload_0_42_25_real,
  output     [15:0]   io_coef_out_payload_0_42_25_imag,
  output     [15:0]   io_coef_out_payload_0_42_26_real,
  output     [15:0]   io_coef_out_payload_0_42_26_imag,
  output     [15:0]   io_coef_out_payload_0_42_27_real,
  output     [15:0]   io_coef_out_payload_0_42_27_imag,
  output     [15:0]   io_coef_out_payload_0_42_28_real,
  output     [15:0]   io_coef_out_payload_0_42_28_imag,
  output     [15:0]   io_coef_out_payload_0_42_29_real,
  output     [15:0]   io_coef_out_payload_0_42_29_imag,
  output     [15:0]   io_coef_out_payload_0_42_30_real,
  output     [15:0]   io_coef_out_payload_0_42_30_imag,
  output     [15:0]   io_coef_out_payload_0_42_31_real,
  output     [15:0]   io_coef_out_payload_0_42_31_imag,
  output     [15:0]   io_coef_out_payload_0_42_32_real,
  output     [15:0]   io_coef_out_payload_0_42_32_imag,
  output     [15:0]   io_coef_out_payload_0_42_33_real,
  output     [15:0]   io_coef_out_payload_0_42_33_imag,
  output     [15:0]   io_coef_out_payload_0_42_34_real,
  output     [15:0]   io_coef_out_payload_0_42_34_imag,
  output     [15:0]   io_coef_out_payload_0_42_35_real,
  output     [15:0]   io_coef_out_payload_0_42_35_imag,
  output     [15:0]   io_coef_out_payload_0_42_36_real,
  output     [15:0]   io_coef_out_payload_0_42_36_imag,
  output     [15:0]   io_coef_out_payload_0_42_37_real,
  output     [15:0]   io_coef_out_payload_0_42_37_imag,
  output     [15:0]   io_coef_out_payload_0_42_38_real,
  output     [15:0]   io_coef_out_payload_0_42_38_imag,
  output     [15:0]   io_coef_out_payload_0_42_39_real,
  output     [15:0]   io_coef_out_payload_0_42_39_imag,
  output     [15:0]   io_coef_out_payload_0_42_40_real,
  output     [15:0]   io_coef_out_payload_0_42_40_imag,
  output     [15:0]   io_coef_out_payload_0_42_41_real,
  output     [15:0]   io_coef_out_payload_0_42_41_imag,
  output     [15:0]   io_coef_out_payload_0_42_42_real,
  output     [15:0]   io_coef_out_payload_0_42_42_imag,
  output     [15:0]   io_coef_out_payload_0_42_43_real,
  output     [15:0]   io_coef_out_payload_0_42_43_imag,
  output     [15:0]   io_coef_out_payload_0_42_44_real,
  output     [15:0]   io_coef_out_payload_0_42_44_imag,
  output     [15:0]   io_coef_out_payload_0_42_45_real,
  output     [15:0]   io_coef_out_payload_0_42_45_imag,
  output     [15:0]   io_coef_out_payload_0_42_46_real,
  output     [15:0]   io_coef_out_payload_0_42_46_imag,
  output     [15:0]   io_coef_out_payload_0_42_47_real,
  output     [15:0]   io_coef_out_payload_0_42_47_imag,
  output     [15:0]   io_coef_out_payload_0_42_48_real,
  output     [15:0]   io_coef_out_payload_0_42_48_imag,
  output     [15:0]   io_coef_out_payload_0_42_49_real,
  output     [15:0]   io_coef_out_payload_0_42_49_imag,
  output     [15:0]   io_coef_out_payload_0_43_0_real,
  output     [15:0]   io_coef_out_payload_0_43_0_imag,
  output     [15:0]   io_coef_out_payload_0_43_1_real,
  output     [15:0]   io_coef_out_payload_0_43_1_imag,
  output     [15:0]   io_coef_out_payload_0_43_2_real,
  output     [15:0]   io_coef_out_payload_0_43_2_imag,
  output     [15:0]   io_coef_out_payload_0_43_3_real,
  output     [15:0]   io_coef_out_payload_0_43_3_imag,
  output     [15:0]   io_coef_out_payload_0_43_4_real,
  output     [15:0]   io_coef_out_payload_0_43_4_imag,
  output     [15:0]   io_coef_out_payload_0_43_5_real,
  output     [15:0]   io_coef_out_payload_0_43_5_imag,
  output     [15:0]   io_coef_out_payload_0_43_6_real,
  output     [15:0]   io_coef_out_payload_0_43_6_imag,
  output     [15:0]   io_coef_out_payload_0_43_7_real,
  output     [15:0]   io_coef_out_payload_0_43_7_imag,
  output     [15:0]   io_coef_out_payload_0_43_8_real,
  output     [15:0]   io_coef_out_payload_0_43_8_imag,
  output     [15:0]   io_coef_out_payload_0_43_9_real,
  output     [15:0]   io_coef_out_payload_0_43_9_imag,
  output     [15:0]   io_coef_out_payload_0_43_10_real,
  output     [15:0]   io_coef_out_payload_0_43_10_imag,
  output     [15:0]   io_coef_out_payload_0_43_11_real,
  output     [15:0]   io_coef_out_payload_0_43_11_imag,
  output     [15:0]   io_coef_out_payload_0_43_12_real,
  output     [15:0]   io_coef_out_payload_0_43_12_imag,
  output     [15:0]   io_coef_out_payload_0_43_13_real,
  output     [15:0]   io_coef_out_payload_0_43_13_imag,
  output     [15:0]   io_coef_out_payload_0_43_14_real,
  output     [15:0]   io_coef_out_payload_0_43_14_imag,
  output     [15:0]   io_coef_out_payload_0_43_15_real,
  output     [15:0]   io_coef_out_payload_0_43_15_imag,
  output     [15:0]   io_coef_out_payload_0_43_16_real,
  output     [15:0]   io_coef_out_payload_0_43_16_imag,
  output     [15:0]   io_coef_out_payload_0_43_17_real,
  output     [15:0]   io_coef_out_payload_0_43_17_imag,
  output     [15:0]   io_coef_out_payload_0_43_18_real,
  output     [15:0]   io_coef_out_payload_0_43_18_imag,
  output     [15:0]   io_coef_out_payload_0_43_19_real,
  output     [15:0]   io_coef_out_payload_0_43_19_imag,
  output     [15:0]   io_coef_out_payload_0_43_20_real,
  output     [15:0]   io_coef_out_payload_0_43_20_imag,
  output     [15:0]   io_coef_out_payload_0_43_21_real,
  output     [15:0]   io_coef_out_payload_0_43_21_imag,
  output     [15:0]   io_coef_out_payload_0_43_22_real,
  output     [15:0]   io_coef_out_payload_0_43_22_imag,
  output     [15:0]   io_coef_out_payload_0_43_23_real,
  output     [15:0]   io_coef_out_payload_0_43_23_imag,
  output     [15:0]   io_coef_out_payload_0_43_24_real,
  output     [15:0]   io_coef_out_payload_0_43_24_imag,
  output     [15:0]   io_coef_out_payload_0_43_25_real,
  output     [15:0]   io_coef_out_payload_0_43_25_imag,
  output     [15:0]   io_coef_out_payload_0_43_26_real,
  output     [15:0]   io_coef_out_payload_0_43_26_imag,
  output     [15:0]   io_coef_out_payload_0_43_27_real,
  output     [15:0]   io_coef_out_payload_0_43_27_imag,
  output     [15:0]   io_coef_out_payload_0_43_28_real,
  output     [15:0]   io_coef_out_payload_0_43_28_imag,
  output     [15:0]   io_coef_out_payload_0_43_29_real,
  output     [15:0]   io_coef_out_payload_0_43_29_imag,
  output     [15:0]   io_coef_out_payload_0_43_30_real,
  output     [15:0]   io_coef_out_payload_0_43_30_imag,
  output     [15:0]   io_coef_out_payload_0_43_31_real,
  output     [15:0]   io_coef_out_payload_0_43_31_imag,
  output     [15:0]   io_coef_out_payload_0_43_32_real,
  output     [15:0]   io_coef_out_payload_0_43_32_imag,
  output     [15:0]   io_coef_out_payload_0_43_33_real,
  output     [15:0]   io_coef_out_payload_0_43_33_imag,
  output     [15:0]   io_coef_out_payload_0_43_34_real,
  output     [15:0]   io_coef_out_payload_0_43_34_imag,
  output     [15:0]   io_coef_out_payload_0_43_35_real,
  output     [15:0]   io_coef_out_payload_0_43_35_imag,
  output     [15:0]   io_coef_out_payload_0_43_36_real,
  output     [15:0]   io_coef_out_payload_0_43_36_imag,
  output     [15:0]   io_coef_out_payload_0_43_37_real,
  output     [15:0]   io_coef_out_payload_0_43_37_imag,
  output     [15:0]   io_coef_out_payload_0_43_38_real,
  output     [15:0]   io_coef_out_payload_0_43_38_imag,
  output     [15:0]   io_coef_out_payload_0_43_39_real,
  output     [15:0]   io_coef_out_payload_0_43_39_imag,
  output     [15:0]   io_coef_out_payload_0_43_40_real,
  output     [15:0]   io_coef_out_payload_0_43_40_imag,
  output     [15:0]   io_coef_out_payload_0_43_41_real,
  output     [15:0]   io_coef_out_payload_0_43_41_imag,
  output     [15:0]   io_coef_out_payload_0_43_42_real,
  output     [15:0]   io_coef_out_payload_0_43_42_imag,
  output     [15:0]   io_coef_out_payload_0_43_43_real,
  output     [15:0]   io_coef_out_payload_0_43_43_imag,
  output     [15:0]   io_coef_out_payload_0_43_44_real,
  output     [15:0]   io_coef_out_payload_0_43_44_imag,
  output     [15:0]   io_coef_out_payload_0_43_45_real,
  output     [15:0]   io_coef_out_payload_0_43_45_imag,
  output     [15:0]   io_coef_out_payload_0_43_46_real,
  output     [15:0]   io_coef_out_payload_0_43_46_imag,
  output     [15:0]   io_coef_out_payload_0_43_47_real,
  output     [15:0]   io_coef_out_payload_0_43_47_imag,
  output     [15:0]   io_coef_out_payload_0_43_48_real,
  output     [15:0]   io_coef_out_payload_0_43_48_imag,
  output     [15:0]   io_coef_out_payload_0_43_49_real,
  output     [15:0]   io_coef_out_payload_0_43_49_imag,
  output     [15:0]   io_coef_out_payload_0_44_0_real,
  output     [15:0]   io_coef_out_payload_0_44_0_imag,
  output     [15:0]   io_coef_out_payload_0_44_1_real,
  output     [15:0]   io_coef_out_payload_0_44_1_imag,
  output     [15:0]   io_coef_out_payload_0_44_2_real,
  output     [15:0]   io_coef_out_payload_0_44_2_imag,
  output     [15:0]   io_coef_out_payload_0_44_3_real,
  output     [15:0]   io_coef_out_payload_0_44_3_imag,
  output     [15:0]   io_coef_out_payload_0_44_4_real,
  output     [15:0]   io_coef_out_payload_0_44_4_imag,
  output     [15:0]   io_coef_out_payload_0_44_5_real,
  output     [15:0]   io_coef_out_payload_0_44_5_imag,
  output     [15:0]   io_coef_out_payload_0_44_6_real,
  output     [15:0]   io_coef_out_payload_0_44_6_imag,
  output     [15:0]   io_coef_out_payload_0_44_7_real,
  output     [15:0]   io_coef_out_payload_0_44_7_imag,
  output     [15:0]   io_coef_out_payload_0_44_8_real,
  output     [15:0]   io_coef_out_payload_0_44_8_imag,
  output     [15:0]   io_coef_out_payload_0_44_9_real,
  output     [15:0]   io_coef_out_payload_0_44_9_imag,
  output     [15:0]   io_coef_out_payload_0_44_10_real,
  output     [15:0]   io_coef_out_payload_0_44_10_imag,
  output     [15:0]   io_coef_out_payload_0_44_11_real,
  output     [15:0]   io_coef_out_payload_0_44_11_imag,
  output     [15:0]   io_coef_out_payload_0_44_12_real,
  output     [15:0]   io_coef_out_payload_0_44_12_imag,
  output     [15:0]   io_coef_out_payload_0_44_13_real,
  output     [15:0]   io_coef_out_payload_0_44_13_imag,
  output     [15:0]   io_coef_out_payload_0_44_14_real,
  output     [15:0]   io_coef_out_payload_0_44_14_imag,
  output     [15:0]   io_coef_out_payload_0_44_15_real,
  output     [15:0]   io_coef_out_payload_0_44_15_imag,
  output     [15:0]   io_coef_out_payload_0_44_16_real,
  output     [15:0]   io_coef_out_payload_0_44_16_imag,
  output     [15:0]   io_coef_out_payload_0_44_17_real,
  output     [15:0]   io_coef_out_payload_0_44_17_imag,
  output     [15:0]   io_coef_out_payload_0_44_18_real,
  output     [15:0]   io_coef_out_payload_0_44_18_imag,
  output     [15:0]   io_coef_out_payload_0_44_19_real,
  output     [15:0]   io_coef_out_payload_0_44_19_imag,
  output     [15:0]   io_coef_out_payload_0_44_20_real,
  output     [15:0]   io_coef_out_payload_0_44_20_imag,
  output     [15:0]   io_coef_out_payload_0_44_21_real,
  output     [15:0]   io_coef_out_payload_0_44_21_imag,
  output     [15:0]   io_coef_out_payload_0_44_22_real,
  output     [15:0]   io_coef_out_payload_0_44_22_imag,
  output     [15:0]   io_coef_out_payload_0_44_23_real,
  output     [15:0]   io_coef_out_payload_0_44_23_imag,
  output     [15:0]   io_coef_out_payload_0_44_24_real,
  output     [15:0]   io_coef_out_payload_0_44_24_imag,
  output     [15:0]   io_coef_out_payload_0_44_25_real,
  output     [15:0]   io_coef_out_payload_0_44_25_imag,
  output     [15:0]   io_coef_out_payload_0_44_26_real,
  output     [15:0]   io_coef_out_payload_0_44_26_imag,
  output     [15:0]   io_coef_out_payload_0_44_27_real,
  output     [15:0]   io_coef_out_payload_0_44_27_imag,
  output     [15:0]   io_coef_out_payload_0_44_28_real,
  output     [15:0]   io_coef_out_payload_0_44_28_imag,
  output     [15:0]   io_coef_out_payload_0_44_29_real,
  output     [15:0]   io_coef_out_payload_0_44_29_imag,
  output     [15:0]   io_coef_out_payload_0_44_30_real,
  output     [15:0]   io_coef_out_payload_0_44_30_imag,
  output     [15:0]   io_coef_out_payload_0_44_31_real,
  output     [15:0]   io_coef_out_payload_0_44_31_imag,
  output     [15:0]   io_coef_out_payload_0_44_32_real,
  output     [15:0]   io_coef_out_payload_0_44_32_imag,
  output     [15:0]   io_coef_out_payload_0_44_33_real,
  output     [15:0]   io_coef_out_payload_0_44_33_imag,
  output     [15:0]   io_coef_out_payload_0_44_34_real,
  output     [15:0]   io_coef_out_payload_0_44_34_imag,
  output     [15:0]   io_coef_out_payload_0_44_35_real,
  output     [15:0]   io_coef_out_payload_0_44_35_imag,
  output     [15:0]   io_coef_out_payload_0_44_36_real,
  output     [15:0]   io_coef_out_payload_0_44_36_imag,
  output     [15:0]   io_coef_out_payload_0_44_37_real,
  output     [15:0]   io_coef_out_payload_0_44_37_imag,
  output     [15:0]   io_coef_out_payload_0_44_38_real,
  output     [15:0]   io_coef_out_payload_0_44_38_imag,
  output     [15:0]   io_coef_out_payload_0_44_39_real,
  output     [15:0]   io_coef_out_payload_0_44_39_imag,
  output     [15:0]   io_coef_out_payload_0_44_40_real,
  output     [15:0]   io_coef_out_payload_0_44_40_imag,
  output     [15:0]   io_coef_out_payload_0_44_41_real,
  output     [15:0]   io_coef_out_payload_0_44_41_imag,
  output     [15:0]   io_coef_out_payload_0_44_42_real,
  output     [15:0]   io_coef_out_payload_0_44_42_imag,
  output     [15:0]   io_coef_out_payload_0_44_43_real,
  output     [15:0]   io_coef_out_payload_0_44_43_imag,
  output     [15:0]   io_coef_out_payload_0_44_44_real,
  output     [15:0]   io_coef_out_payload_0_44_44_imag,
  output     [15:0]   io_coef_out_payload_0_44_45_real,
  output     [15:0]   io_coef_out_payload_0_44_45_imag,
  output     [15:0]   io_coef_out_payload_0_44_46_real,
  output     [15:0]   io_coef_out_payload_0_44_46_imag,
  output     [15:0]   io_coef_out_payload_0_44_47_real,
  output     [15:0]   io_coef_out_payload_0_44_47_imag,
  output     [15:0]   io_coef_out_payload_0_44_48_real,
  output     [15:0]   io_coef_out_payload_0_44_48_imag,
  output     [15:0]   io_coef_out_payload_0_44_49_real,
  output     [15:0]   io_coef_out_payload_0_44_49_imag,
  output     [15:0]   io_coef_out_payload_0_45_0_real,
  output     [15:0]   io_coef_out_payload_0_45_0_imag,
  output     [15:0]   io_coef_out_payload_0_45_1_real,
  output     [15:0]   io_coef_out_payload_0_45_1_imag,
  output     [15:0]   io_coef_out_payload_0_45_2_real,
  output     [15:0]   io_coef_out_payload_0_45_2_imag,
  output     [15:0]   io_coef_out_payload_0_45_3_real,
  output     [15:0]   io_coef_out_payload_0_45_3_imag,
  output     [15:0]   io_coef_out_payload_0_45_4_real,
  output     [15:0]   io_coef_out_payload_0_45_4_imag,
  output     [15:0]   io_coef_out_payload_0_45_5_real,
  output     [15:0]   io_coef_out_payload_0_45_5_imag,
  output     [15:0]   io_coef_out_payload_0_45_6_real,
  output     [15:0]   io_coef_out_payload_0_45_6_imag,
  output     [15:0]   io_coef_out_payload_0_45_7_real,
  output     [15:0]   io_coef_out_payload_0_45_7_imag,
  output     [15:0]   io_coef_out_payload_0_45_8_real,
  output     [15:0]   io_coef_out_payload_0_45_8_imag,
  output     [15:0]   io_coef_out_payload_0_45_9_real,
  output     [15:0]   io_coef_out_payload_0_45_9_imag,
  output     [15:0]   io_coef_out_payload_0_45_10_real,
  output     [15:0]   io_coef_out_payload_0_45_10_imag,
  output     [15:0]   io_coef_out_payload_0_45_11_real,
  output     [15:0]   io_coef_out_payload_0_45_11_imag,
  output     [15:0]   io_coef_out_payload_0_45_12_real,
  output     [15:0]   io_coef_out_payload_0_45_12_imag,
  output     [15:0]   io_coef_out_payload_0_45_13_real,
  output     [15:0]   io_coef_out_payload_0_45_13_imag,
  output     [15:0]   io_coef_out_payload_0_45_14_real,
  output     [15:0]   io_coef_out_payload_0_45_14_imag,
  output     [15:0]   io_coef_out_payload_0_45_15_real,
  output     [15:0]   io_coef_out_payload_0_45_15_imag,
  output     [15:0]   io_coef_out_payload_0_45_16_real,
  output     [15:0]   io_coef_out_payload_0_45_16_imag,
  output     [15:0]   io_coef_out_payload_0_45_17_real,
  output     [15:0]   io_coef_out_payload_0_45_17_imag,
  output     [15:0]   io_coef_out_payload_0_45_18_real,
  output     [15:0]   io_coef_out_payload_0_45_18_imag,
  output     [15:0]   io_coef_out_payload_0_45_19_real,
  output     [15:0]   io_coef_out_payload_0_45_19_imag,
  output     [15:0]   io_coef_out_payload_0_45_20_real,
  output     [15:0]   io_coef_out_payload_0_45_20_imag,
  output     [15:0]   io_coef_out_payload_0_45_21_real,
  output     [15:0]   io_coef_out_payload_0_45_21_imag,
  output     [15:0]   io_coef_out_payload_0_45_22_real,
  output     [15:0]   io_coef_out_payload_0_45_22_imag,
  output     [15:0]   io_coef_out_payload_0_45_23_real,
  output     [15:0]   io_coef_out_payload_0_45_23_imag,
  output     [15:0]   io_coef_out_payload_0_45_24_real,
  output     [15:0]   io_coef_out_payload_0_45_24_imag,
  output     [15:0]   io_coef_out_payload_0_45_25_real,
  output     [15:0]   io_coef_out_payload_0_45_25_imag,
  output     [15:0]   io_coef_out_payload_0_45_26_real,
  output     [15:0]   io_coef_out_payload_0_45_26_imag,
  output     [15:0]   io_coef_out_payload_0_45_27_real,
  output     [15:0]   io_coef_out_payload_0_45_27_imag,
  output     [15:0]   io_coef_out_payload_0_45_28_real,
  output     [15:0]   io_coef_out_payload_0_45_28_imag,
  output     [15:0]   io_coef_out_payload_0_45_29_real,
  output     [15:0]   io_coef_out_payload_0_45_29_imag,
  output     [15:0]   io_coef_out_payload_0_45_30_real,
  output     [15:0]   io_coef_out_payload_0_45_30_imag,
  output     [15:0]   io_coef_out_payload_0_45_31_real,
  output     [15:0]   io_coef_out_payload_0_45_31_imag,
  output     [15:0]   io_coef_out_payload_0_45_32_real,
  output     [15:0]   io_coef_out_payload_0_45_32_imag,
  output     [15:0]   io_coef_out_payload_0_45_33_real,
  output     [15:0]   io_coef_out_payload_0_45_33_imag,
  output     [15:0]   io_coef_out_payload_0_45_34_real,
  output     [15:0]   io_coef_out_payload_0_45_34_imag,
  output     [15:0]   io_coef_out_payload_0_45_35_real,
  output     [15:0]   io_coef_out_payload_0_45_35_imag,
  output     [15:0]   io_coef_out_payload_0_45_36_real,
  output     [15:0]   io_coef_out_payload_0_45_36_imag,
  output     [15:0]   io_coef_out_payload_0_45_37_real,
  output     [15:0]   io_coef_out_payload_0_45_37_imag,
  output     [15:0]   io_coef_out_payload_0_45_38_real,
  output     [15:0]   io_coef_out_payload_0_45_38_imag,
  output     [15:0]   io_coef_out_payload_0_45_39_real,
  output     [15:0]   io_coef_out_payload_0_45_39_imag,
  output     [15:0]   io_coef_out_payload_0_45_40_real,
  output     [15:0]   io_coef_out_payload_0_45_40_imag,
  output     [15:0]   io_coef_out_payload_0_45_41_real,
  output     [15:0]   io_coef_out_payload_0_45_41_imag,
  output     [15:0]   io_coef_out_payload_0_45_42_real,
  output     [15:0]   io_coef_out_payload_0_45_42_imag,
  output     [15:0]   io_coef_out_payload_0_45_43_real,
  output     [15:0]   io_coef_out_payload_0_45_43_imag,
  output     [15:0]   io_coef_out_payload_0_45_44_real,
  output     [15:0]   io_coef_out_payload_0_45_44_imag,
  output     [15:0]   io_coef_out_payload_0_45_45_real,
  output     [15:0]   io_coef_out_payload_0_45_45_imag,
  output     [15:0]   io_coef_out_payload_0_45_46_real,
  output     [15:0]   io_coef_out_payload_0_45_46_imag,
  output     [15:0]   io_coef_out_payload_0_45_47_real,
  output     [15:0]   io_coef_out_payload_0_45_47_imag,
  output     [15:0]   io_coef_out_payload_0_45_48_real,
  output     [15:0]   io_coef_out_payload_0_45_48_imag,
  output     [15:0]   io_coef_out_payload_0_45_49_real,
  output     [15:0]   io_coef_out_payload_0_45_49_imag,
  output     [15:0]   io_coef_out_payload_0_46_0_real,
  output     [15:0]   io_coef_out_payload_0_46_0_imag,
  output     [15:0]   io_coef_out_payload_0_46_1_real,
  output     [15:0]   io_coef_out_payload_0_46_1_imag,
  output     [15:0]   io_coef_out_payload_0_46_2_real,
  output     [15:0]   io_coef_out_payload_0_46_2_imag,
  output     [15:0]   io_coef_out_payload_0_46_3_real,
  output     [15:0]   io_coef_out_payload_0_46_3_imag,
  output     [15:0]   io_coef_out_payload_0_46_4_real,
  output     [15:0]   io_coef_out_payload_0_46_4_imag,
  output     [15:0]   io_coef_out_payload_0_46_5_real,
  output     [15:0]   io_coef_out_payload_0_46_5_imag,
  output     [15:0]   io_coef_out_payload_0_46_6_real,
  output     [15:0]   io_coef_out_payload_0_46_6_imag,
  output     [15:0]   io_coef_out_payload_0_46_7_real,
  output     [15:0]   io_coef_out_payload_0_46_7_imag,
  output     [15:0]   io_coef_out_payload_0_46_8_real,
  output     [15:0]   io_coef_out_payload_0_46_8_imag,
  output     [15:0]   io_coef_out_payload_0_46_9_real,
  output     [15:0]   io_coef_out_payload_0_46_9_imag,
  output     [15:0]   io_coef_out_payload_0_46_10_real,
  output     [15:0]   io_coef_out_payload_0_46_10_imag,
  output     [15:0]   io_coef_out_payload_0_46_11_real,
  output     [15:0]   io_coef_out_payload_0_46_11_imag,
  output     [15:0]   io_coef_out_payload_0_46_12_real,
  output     [15:0]   io_coef_out_payload_0_46_12_imag,
  output     [15:0]   io_coef_out_payload_0_46_13_real,
  output     [15:0]   io_coef_out_payload_0_46_13_imag,
  output     [15:0]   io_coef_out_payload_0_46_14_real,
  output     [15:0]   io_coef_out_payload_0_46_14_imag,
  output     [15:0]   io_coef_out_payload_0_46_15_real,
  output     [15:0]   io_coef_out_payload_0_46_15_imag,
  output     [15:0]   io_coef_out_payload_0_46_16_real,
  output     [15:0]   io_coef_out_payload_0_46_16_imag,
  output     [15:0]   io_coef_out_payload_0_46_17_real,
  output     [15:0]   io_coef_out_payload_0_46_17_imag,
  output     [15:0]   io_coef_out_payload_0_46_18_real,
  output     [15:0]   io_coef_out_payload_0_46_18_imag,
  output     [15:0]   io_coef_out_payload_0_46_19_real,
  output     [15:0]   io_coef_out_payload_0_46_19_imag,
  output     [15:0]   io_coef_out_payload_0_46_20_real,
  output     [15:0]   io_coef_out_payload_0_46_20_imag,
  output     [15:0]   io_coef_out_payload_0_46_21_real,
  output     [15:0]   io_coef_out_payload_0_46_21_imag,
  output     [15:0]   io_coef_out_payload_0_46_22_real,
  output     [15:0]   io_coef_out_payload_0_46_22_imag,
  output     [15:0]   io_coef_out_payload_0_46_23_real,
  output     [15:0]   io_coef_out_payload_0_46_23_imag,
  output     [15:0]   io_coef_out_payload_0_46_24_real,
  output     [15:0]   io_coef_out_payload_0_46_24_imag,
  output     [15:0]   io_coef_out_payload_0_46_25_real,
  output     [15:0]   io_coef_out_payload_0_46_25_imag,
  output     [15:0]   io_coef_out_payload_0_46_26_real,
  output     [15:0]   io_coef_out_payload_0_46_26_imag,
  output     [15:0]   io_coef_out_payload_0_46_27_real,
  output     [15:0]   io_coef_out_payload_0_46_27_imag,
  output     [15:0]   io_coef_out_payload_0_46_28_real,
  output     [15:0]   io_coef_out_payload_0_46_28_imag,
  output     [15:0]   io_coef_out_payload_0_46_29_real,
  output     [15:0]   io_coef_out_payload_0_46_29_imag,
  output     [15:0]   io_coef_out_payload_0_46_30_real,
  output     [15:0]   io_coef_out_payload_0_46_30_imag,
  output     [15:0]   io_coef_out_payload_0_46_31_real,
  output     [15:0]   io_coef_out_payload_0_46_31_imag,
  output     [15:0]   io_coef_out_payload_0_46_32_real,
  output     [15:0]   io_coef_out_payload_0_46_32_imag,
  output     [15:0]   io_coef_out_payload_0_46_33_real,
  output     [15:0]   io_coef_out_payload_0_46_33_imag,
  output     [15:0]   io_coef_out_payload_0_46_34_real,
  output     [15:0]   io_coef_out_payload_0_46_34_imag,
  output     [15:0]   io_coef_out_payload_0_46_35_real,
  output     [15:0]   io_coef_out_payload_0_46_35_imag,
  output     [15:0]   io_coef_out_payload_0_46_36_real,
  output     [15:0]   io_coef_out_payload_0_46_36_imag,
  output     [15:0]   io_coef_out_payload_0_46_37_real,
  output     [15:0]   io_coef_out_payload_0_46_37_imag,
  output     [15:0]   io_coef_out_payload_0_46_38_real,
  output     [15:0]   io_coef_out_payload_0_46_38_imag,
  output     [15:0]   io_coef_out_payload_0_46_39_real,
  output     [15:0]   io_coef_out_payload_0_46_39_imag,
  output     [15:0]   io_coef_out_payload_0_46_40_real,
  output     [15:0]   io_coef_out_payload_0_46_40_imag,
  output     [15:0]   io_coef_out_payload_0_46_41_real,
  output     [15:0]   io_coef_out_payload_0_46_41_imag,
  output     [15:0]   io_coef_out_payload_0_46_42_real,
  output     [15:0]   io_coef_out_payload_0_46_42_imag,
  output     [15:0]   io_coef_out_payload_0_46_43_real,
  output     [15:0]   io_coef_out_payload_0_46_43_imag,
  output     [15:0]   io_coef_out_payload_0_46_44_real,
  output     [15:0]   io_coef_out_payload_0_46_44_imag,
  output     [15:0]   io_coef_out_payload_0_46_45_real,
  output     [15:0]   io_coef_out_payload_0_46_45_imag,
  output     [15:0]   io_coef_out_payload_0_46_46_real,
  output     [15:0]   io_coef_out_payload_0_46_46_imag,
  output     [15:0]   io_coef_out_payload_0_46_47_real,
  output     [15:0]   io_coef_out_payload_0_46_47_imag,
  output     [15:0]   io_coef_out_payload_0_46_48_real,
  output     [15:0]   io_coef_out_payload_0_46_48_imag,
  output     [15:0]   io_coef_out_payload_0_46_49_real,
  output     [15:0]   io_coef_out_payload_0_46_49_imag,
  output     [15:0]   io_coef_out_payload_0_47_0_real,
  output     [15:0]   io_coef_out_payload_0_47_0_imag,
  output     [15:0]   io_coef_out_payload_0_47_1_real,
  output     [15:0]   io_coef_out_payload_0_47_1_imag,
  output     [15:0]   io_coef_out_payload_0_47_2_real,
  output     [15:0]   io_coef_out_payload_0_47_2_imag,
  output     [15:0]   io_coef_out_payload_0_47_3_real,
  output     [15:0]   io_coef_out_payload_0_47_3_imag,
  output     [15:0]   io_coef_out_payload_0_47_4_real,
  output     [15:0]   io_coef_out_payload_0_47_4_imag,
  output     [15:0]   io_coef_out_payload_0_47_5_real,
  output     [15:0]   io_coef_out_payload_0_47_5_imag,
  output     [15:0]   io_coef_out_payload_0_47_6_real,
  output     [15:0]   io_coef_out_payload_0_47_6_imag,
  output     [15:0]   io_coef_out_payload_0_47_7_real,
  output     [15:0]   io_coef_out_payload_0_47_7_imag,
  output     [15:0]   io_coef_out_payload_0_47_8_real,
  output     [15:0]   io_coef_out_payload_0_47_8_imag,
  output     [15:0]   io_coef_out_payload_0_47_9_real,
  output     [15:0]   io_coef_out_payload_0_47_9_imag,
  output     [15:0]   io_coef_out_payload_0_47_10_real,
  output     [15:0]   io_coef_out_payload_0_47_10_imag,
  output     [15:0]   io_coef_out_payload_0_47_11_real,
  output     [15:0]   io_coef_out_payload_0_47_11_imag,
  output     [15:0]   io_coef_out_payload_0_47_12_real,
  output     [15:0]   io_coef_out_payload_0_47_12_imag,
  output     [15:0]   io_coef_out_payload_0_47_13_real,
  output     [15:0]   io_coef_out_payload_0_47_13_imag,
  output     [15:0]   io_coef_out_payload_0_47_14_real,
  output     [15:0]   io_coef_out_payload_0_47_14_imag,
  output     [15:0]   io_coef_out_payload_0_47_15_real,
  output     [15:0]   io_coef_out_payload_0_47_15_imag,
  output     [15:0]   io_coef_out_payload_0_47_16_real,
  output     [15:0]   io_coef_out_payload_0_47_16_imag,
  output     [15:0]   io_coef_out_payload_0_47_17_real,
  output     [15:0]   io_coef_out_payload_0_47_17_imag,
  output     [15:0]   io_coef_out_payload_0_47_18_real,
  output     [15:0]   io_coef_out_payload_0_47_18_imag,
  output     [15:0]   io_coef_out_payload_0_47_19_real,
  output     [15:0]   io_coef_out_payload_0_47_19_imag,
  output     [15:0]   io_coef_out_payload_0_47_20_real,
  output     [15:0]   io_coef_out_payload_0_47_20_imag,
  output     [15:0]   io_coef_out_payload_0_47_21_real,
  output     [15:0]   io_coef_out_payload_0_47_21_imag,
  output     [15:0]   io_coef_out_payload_0_47_22_real,
  output     [15:0]   io_coef_out_payload_0_47_22_imag,
  output     [15:0]   io_coef_out_payload_0_47_23_real,
  output     [15:0]   io_coef_out_payload_0_47_23_imag,
  output     [15:0]   io_coef_out_payload_0_47_24_real,
  output     [15:0]   io_coef_out_payload_0_47_24_imag,
  output     [15:0]   io_coef_out_payload_0_47_25_real,
  output     [15:0]   io_coef_out_payload_0_47_25_imag,
  output     [15:0]   io_coef_out_payload_0_47_26_real,
  output     [15:0]   io_coef_out_payload_0_47_26_imag,
  output     [15:0]   io_coef_out_payload_0_47_27_real,
  output     [15:0]   io_coef_out_payload_0_47_27_imag,
  output     [15:0]   io_coef_out_payload_0_47_28_real,
  output     [15:0]   io_coef_out_payload_0_47_28_imag,
  output     [15:0]   io_coef_out_payload_0_47_29_real,
  output     [15:0]   io_coef_out_payload_0_47_29_imag,
  output     [15:0]   io_coef_out_payload_0_47_30_real,
  output     [15:0]   io_coef_out_payload_0_47_30_imag,
  output     [15:0]   io_coef_out_payload_0_47_31_real,
  output     [15:0]   io_coef_out_payload_0_47_31_imag,
  output     [15:0]   io_coef_out_payload_0_47_32_real,
  output     [15:0]   io_coef_out_payload_0_47_32_imag,
  output     [15:0]   io_coef_out_payload_0_47_33_real,
  output     [15:0]   io_coef_out_payload_0_47_33_imag,
  output     [15:0]   io_coef_out_payload_0_47_34_real,
  output     [15:0]   io_coef_out_payload_0_47_34_imag,
  output     [15:0]   io_coef_out_payload_0_47_35_real,
  output     [15:0]   io_coef_out_payload_0_47_35_imag,
  output     [15:0]   io_coef_out_payload_0_47_36_real,
  output     [15:0]   io_coef_out_payload_0_47_36_imag,
  output     [15:0]   io_coef_out_payload_0_47_37_real,
  output     [15:0]   io_coef_out_payload_0_47_37_imag,
  output     [15:0]   io_coef_out_payload_0_47_38_real,
  output     [15:0]   io_coef_out_payload_0_47_38_imag,
  output     [15:0]   io_coef_out_payload_0_47_39_real,
  output     [15:0]   io_coef_out_payload_0_47_39_imag,
  output     [15:0]   io_coef_out_payload_0_47_40_real,
  output     [15:0]   io_coef_out_payload_0_47_40_imag,
  output     [15:0]   io_coef_out_payload_0_47_41_real,
  output     [15:0]   io_coef_out_payload_0_47_41_imag,
  output     [15:0]   io_coef_out_payload_0_47_42_real,
  output     [15:0]   io_coef_out_payload_0_47_42_imag,
  output     [15:0]   io_coef_out_payload_0_47_43_real,
  output     [15:0]   io_coef_out_payload_0_47_43_imag,
  output     [15:0]   io_coef_out_payload_0_47_44_real,
  output     [15:0]   io_coef_out_payload_0_47_44_imag,
  output     [15:0]   io_coef_out_payload_0_47_45_real,
  output     [15:0]   io_coef_out_payload_0_47_45_imag,
  output     [15:0]   io_coef_out_payload_0_47_46_real,
  output     [15:0]   io_coef_out_payload_0_47_46_imag,
  output     [15:0]   io_coef_out_payload_0_47_47_real,
  output     [15:0]   io_coef_out_payload_0_47_47_imag,
  output     [15:0]   io_coef_out_payload_0_47_48_real,
  output     [15:0]   io_coef_out_payload_0_47_48_imag,
  output     [15:0]   io_coef_out_payload_0_47_49_real,
  output     [15:0]   io_coef_out_payload_0_47_49_imag,
  output     [15:0]   io_coef_out_payload_0_48_0_real,
  output     [15:0]   io_coef_out_payload_0_48_0_imag,
  output     [15:0]   io_coef_out_payload_0_48_1_real,
  output     [15:0]   io_coef_out_payload_0_48_1_imag,
  output     [15:0]   io_coef_out_payload_0_48_2_real,
  output     [15:0]   io_coef_out_payload_0_48_2_imag,
  output     [15:0]   io_coef_out_payload_0_48_3_real,
  output     [15:0]   io_coef_out_payload_0_48_3_imag,
  output     [15:0]   io_coef_out_payload_0_48_4_real,
  output     [15:0]   io_coef_out_payload_0_48_4_imag,
  output     [15:0]   io_coef_out_payload_0_48_5_real,
  output     [15:0]   io_coef_out_payload_0_48_5_imag,
  output     [15:0]   io_coef_out_payload_0_48_6_real,
  output     [15:0]   io_coef_out_payload_0_48_6_imag,
  output     [15:0]   io_coef_out_payload_0_48_7_real,
  output     [15:0]   io_coef_out_payload_0_48_7_imag,
  output     [15:0]   io_coef_out_payload_0_48_8_real,
  output     [15:0]   io_coef_out_payload_0_48_8_imag,
  output     [15:0]   io_coef_out_payload_0_48_9_real,
  output     [15:0]   io_coef_out_payload_0_48_9_imag,
  output     [15:0]   io_coef_out_payload_0_48_10_real,
  output     [15:0]   io_coef_out_payload_0_48_10_imag,
  output     [15:0]   io_coef_out_payload_0_48_11_real,
  output     [15:0]   io_coef_out_payload_0_48_11_imag,
  output     [15:0]   io_coef_out_payload_0_48_12_real,
  output     [15:0]   io_coef_out_payload_0_48_12_imag,
  output     [15:0]   io_coef_out_payload_0_48_13_real,
  output     [15:0]   io_coef_out_payload_0_48_13_imag,
  output     [15:0]   io_coef_out_payload_0_48_14_real,
  output     [15:0]   io_coef_out_payload_0_48_14_imag,
  output     [15:0]   io_coef_out_payload_0_48_15_real,
  output     [15:0]   io_coef_out_payload_0_48_15_imag,
  output     [15:0]   io_coef_out_payload_0_48_16_real,
  output     [15:0]   io_coef_out_payload_0_48_16_imag,
  output     [15:0]   io_coef_out_payload_0_48_17_real,
  output     [15:0]   io_coef_out_payload_0_48_17_imag,
  output     [15:0]   io_coef_out_payload_0_48_18_real,
  output     [15:0]   io_coef_out_payload_0_48_18_imag,
  output     [15:0]   io_coef_out_payload_0_48_19_real,
  output     [15:0]   io_coef_out_payload_0_48_19_imag,
  output     [15:0]   io_coef_out_payload_0_48_20_real,
  output     [15:0]   io_coef_out_payload_0_48_20_imag,
  output     [15:0]   io_coef_out_payload_0_48_21_real,
  output     [15:0]   io_coef_out_payload_0_48_21_imag,
  output     [15:0]   io_coef_out_payload_0_48_22_real,
  output     [15:0]   io_coef_out_payload_0_48_22_imag,
  output     [15:0]   io_coef_out_payload_0_48_23_real,
  output     [15:0]   io_coef_out_payload_0_48_23_imag,
  output     [15:0]   io_coef_out_payload_0_48_24_real,
  output     [15:0]   io_coef_out_payload_0_48_24_imag,
  output     [15:0]   io_coef_out_payload_0_48_25_real,
  output     [15:0]   io_coef_out_payload_0_48_25_imag,
  output     [15:0]   io_coef_out_payload_0_48_26_real,
  output     [15:0]   io_coef_out_payload_0_48_26_imag,
  output     [15:0]   io_coef_out_payload_0_48_27_real,
  output     [15:0]   io_coef_out_payload_0_48_27_imag,
  output     [15:0]   io_coef_out_payload_0_48_28_real,
  output     [15:0]   io_coef_out_payload_0_48_28_imag,
  output     [15:0]   io_coef_out_payload_0_48_29_real,
  output     [15:0]   io_coef_out_payload_0_48_29_imag,
  output     [15:0]   io_coef_out_payload_0_48_30_real,
  output     [15:0]   io_coef_out_payload_0_48_30_imag,
  output     [15:0]   io_coef_out_payload_0_48_31_real,
  output     [15:0]   io_coef_out_payload_0_48_31_imag,
  output     [15:0]   io_coef_out_payload_0_48_32_real,
  output     [15:0]   io_coef_out_payload_0_48_32_imag,
  output     [15:0]   io_coef_out_payload_0_48_33_real,
  output     [15:0]   io_coef_out_payload_0_48_33_imag,
  output     [15:0]   io_coef_out_payload_0_48_34_real,
  output     [15:0]   io_coef_out_payload_0_48_34_imag,
  output     [15:0]   io_coef_out_payload_0_48_35_real,
  output     [15:0]   io_coef_out_payload_0_48_35_imag,
  output     [15:0]   io_coef_out_payload_0_48_36_real,
  output     [15:0]   io_coef_out_payload_0_48_36_imag,
  output     [15:0]   io_coef_out_payload_0_48_37_real,
  output     [15:0]   io_coef_out_payload_0_48_37_imag,
  output     [15:0]   io_coef_out_payload_0_48_38_real,
  output     [15:0]   io_coef_out_payload_0_48_38_imag,
  output     [15:0]   io_coef_out_payload_0_48_39_real,
  output     [15:0]   io_coef_out_payload_0_48_39_imag,
  output     [15:0]   io_coef_out_payload_0_48_40_real,
  output     [15:0]   io_coef_out_payload_0_48_40_imag,
  output     [15:0]   io_coef_out_payload_0_48_41_real,
  output     [15:0]   io_coef_out_payload_0_48_41_imag,
  output     [15:0]   io_coef_out_payload_0_48_42_real,
  output     [15:0]   io_coef_out_payload_0_48_42_imag,
  output     [15:0]   io_coef_out_payload_0_48_43_real,
  output     [15:0]   io_coef_out_payload_0_48_43_imag,
  output     [15:0]   io_coef_out_payload_0_48_44_real,
  output     [15:0]   io_coef_out_payload_0_48_44_imag,
  output     [15:0]   io_coef_out_payload_0_48_45_real,
  output     [15:0]   io_coef_out_payload_0_48_45_imag,
  output     [15:0]   io_coef_out_payload_0_48_46_real,
  output     [15:0]   io_coef_out_payload_0_48_46_imag,
  output     [15:0]   io_coef_out_payload_0_48_47_real,
  output     [15:0]   io_coef_out_payload_0_48_47_imag,
  output     [15:0]   io_coef_out_payload_0_48_48_real,
  output     [15:0]   io_coef_out_payload_0_48_48_imag,
  output     [15:0]   io_coef_out_payload_0_48_49_real,
  output     [15:0]   io_coef_out_payload_0_48_49_imag,
  output     [15:0]   io_coef_out_payload_0_49_0_real,
  output     [15:0]   io_coef_out_payload_0_49_0_imag,
  output     [15:0]   io_coef_out_payload_0_49_1_real,
  output     [15:0]   io_coef_out_payload_0_49_1_imag,
  output     [15:0]   io_coef_out_payload_0_49_2_real,
  output     [15:0]   io_coef_out_payload_0_49_2_imag,
  output     [15:0]   io_coef_out_payload_0_49_3_real,
  output     [15:0]   io_coef_out_payload_0_49_3_imag,
  output     [15:0]   io_coef_out_payload_0_49_4_real,
  output     [15:0]   io_coef_out_payload_0_49_4_imag,
  output     [15:0]   io_coef_out_payload_0_49_5_real,
  output     [15:0]   io_coef_out_payload_0_49_5_imag,
  output     [15:0]   io_coef_out_payload_0_49_6_real,
  output     [15:0]   io_coef_out_payload_0_49_6_imag,
  output     [15:0]   io_coef_out_payload_0_49_7_real,
  output     [15:0]   io_coef_out_payload_0_49_7_imag,
  output     [15:0]   io_coef_out_payload_0_49_8_real,
  output     [15:0]   io_coef_out_payload_0_49_8_imag,
  output     [15:0]   io_coef_out_payload_0_49_9_real,
  output     [15:0]   io_coef_out_payload_0_49_9_imag,
  output     [15:0]   io_coef_out_payload_0_49_10_real,
  output     [15:0]   io_coef_out_payload_0_49_10_imag,
  output     [15:0]   io_coef_out_payload_0_49_11_real,
  output     [15:0]   io_coef_out_payload_0_49_11_imag,
  output     [15:0]   io_coef_out_payload_0_49_12_real,
  output     [15:0]   io_coef_out_payload_0_49_12_imag,
  output     [15:0]   io_coef_out_payload_0_49_13_real,
  output     [15:0]   io_coef_out_payload_0_49_13_imag,
  output     [15:0]   io_coef_out_payload_0_49_14_real,
  output     [15:0]   io_coef_out_payload_0_49_14_imag,
  output     [15:0]   io_coef_out_payload_0_49_15_real,
  output     [15:0]   io_coef_out_payload_0_49_15_imag,
  output     [15:0]   io_coef_out_payload_0_49_16_real,
  output     [15:0]   io_coef_out_payload_0_49_16_imag,
  output     [15:0]   io_coef_out_payload_0_49_17_real,
  output     [15:0]   io_coef_out_payload_0_49_17_imag,
  output     [15:0]   io_coef_out_payload_0_49_18_real,
  output     [15:0]   io_coef_out_payload_0_49_18_imag,
  output     [15:0]   io_coef_out_payload_0_49_19_real,
  output     [15:0]   io_coef_out_payload_0_49_19_imag,
  output     [15:0]   io_coef_out_payload_0_49_20_real,
  output     [15:0]   io_coef_out_payload_0_49_20_imag,
  output     [15:0]   io_coef_out_payload_0_49_21_real,
  output     [15:0]   io_coef_out_payload_0_49_21_imag,
  output     [15:0]   io_coef_out_payload_0_49_22_real,
  output     [15:0]   io_coef_out_payload_0_49_22_imag,
  output     [15:0]   io_coef_out_payload_0_49_23_real,
  output     [15:0]   io_coef_out_payload_0_49_23_imag,
  output     [15:0]   io_coef_out_payload_0_49_24_real,
  output     [15:0]   io_coef_out_payload_0_49_24_imag,
  output     [15:0]   io_coef_out_payload_0_49_25_real,
  output     [15:0]   io_coef_out_payload_0_49_25_imag,
  output     [15:0]   io_coef_out_payload_0_49_26_real,
  output     [15:0]   io_coef_out_payload_0_49_26_imag,
  output     [15:0]   io_coef_out_payload_0_49_27_real,
  output     [15:0]   io_coef_out_payload_0_49_27_imag,
  output     [15:0]   io_coef_out_payload_0_49_28_real,
  output     [15:0]   io_coef_out_payload_0_49_28_imag,
  output     [15:0]   io_coef_out_payload_0_49_29_real,
  output     [15:0]   io_coef_out_payload_0_49_29_imag,
  output     [15:0]   io_coef_out_payload_0_49_30_real,
  output     [15:0]   io_coef_out_payload_0_49_30_imag,
  output     [15:0]   io_coef_out_payload_0_49_31_real,
  output     [15:0]   io_coef_out_payload_0_49_31_imag,
  output     [15:0]   io_coef_out_payload_0_49_32_real,
  output     [15:0]   io_coef_out_payload_0_49_32_imag,
  output     [15:0]   io_coef_out_payload_0_49_33_real,
  output     [15:0]   io_coef_out_payload_0_49_33_imag,
  output     [15:0]   io_coef_out_payload_0_49_34_real,
  output     [15:0]   io_coef_out_payload_0_49_34_imag,
  output     [15:0]   io_coef_out_payload_0_49_35_real,
  output     [15:0]   io_coef_out_payload_0_49_35_imag,
  output     [15:0]   io_coef_out_payload_0_49_36_real,
  output     [15:0]   io_coef_out_payload_0_49_36_imag,
  output     [15:0]   io_coef_out_payload_0_49_37_real,
  output     [15:0]   io_coef_out_payload_0_49_37_imag,
  output     [15:0]   io_coef_out_payload_0_49_38_real,
  output     [15:0]   io_coef_out_payload_0_49_38_imag,
  output     [15:0]   io_coef_out_payload_0_49_39_real,
  output     [15:0]   io_coef_out_payload_0_49_39_imag,
  output     [15:0]   io_coef_out_payload_0_49_40_real,
  output     [15:0]   io_coef_out_payload_0_49_40_imag,
  output     [15:0]   io_coef_out_payload_0_49_41_real,
  output     [15:0]   io_coef_out_payload_0_49_41_imag,
  output     [15:0]   io_coef_out_payload_0_49_42_real,
  output     [15:0]   io_coef_out_payload_0_49_42_imag,
  output     [15:0]   io_coef_out_payload_0_49_43_real,
  output     [15:0]   io_coef_out_payload_0_49_43_imag,
  output     [15:0]   io_coef_out_payload_0_49_44_real,
  output     [15:0]   io_coef_out_payload_0_49_44_imag,
  output     [15:0]   io_coef_out_payload_0_49_45_real,
  output     [15:0]   io_coef_out_payload_0_49_45_imag,
  output     [15:0]   io_coef_out_payload_0_49_46_real,
  output     [15:0]   io_coef_out_payload_0_49_46_imag,
  output     [15:0]   io_coef_out_payload_0_49_47_real,
  output     [15:0]   io_coef_out_payload_0_49_47_imag,
  output     [15:0]   io_coef_out_payload_0_49_48_real,
  output     [15:0]   io_coef_out_payload_0_49_48_imag,
  output     [15:0]   io_coef_out_payload_0_49_49_real,
  output     [15:0]   io_coef_out_payload_0_49_49_imag,
  input               clk,
  input               reset 
);
  reg        [11:0]   _zz_2752_;
  reg        [15:0]   _zz_2753_;
  reg        [15:0]   _zz_2754_;
  reg        [15:0]   _zz_2755_;
  reg        [15:0]   _zz_2756_;
  reg        [15:0]   _zz_2757_;
  reg        [15:0]   _zz_2758_;
  reg        [15:0]   _zz_2759_;
  reg        [15:0]   _zz_2760_;
  reg        [15:0]   _zz_2761_;
  reg        [15:0]   _zz_2762_;
  reg        [15:0]   _zz_2763_;
  reg        [15:0]   _zz_2764_;
  reg        [15:0]   _zz_2765_;
  reg        [15:0]   _zz_2766_;
  reg        [15:0]   _zz_2767_;
  reg        [15:0]   _zz_2768_;
  reg        [15:0]   _zz_2769_;
  reg        [15:0]   _zz_2770_;
  reg        [15:0]   _zz_2771_;
  reg        [15:0]   _zz_2772_;
  reg        [15:0]   _zz_2773_;
  reg        [15:0]   _zz_2774_;
  reg        [15:0]   _zz_2775_;
  reg        [15:0]   _zz_2776_;
  reg        [15:0]   _zz_2777_;
  reg        [15:0]   _zz_2778_;
  reg        [15:0]   _zz_2779_;
  reg        [15:0]   _zz_2780_;
  reg        [15:0]   _zz_2781_;
  reg        [15:0]   _zz_2782_;
  reg        [15:0]   _zz_2783_;
  reg        [15:0]   _zz_2784_;
  reg        [15:0]   _zz_2785_;
  reg        [15:0]   _zz_2786_;
  reg        [15:0]   _zz_2787_;
  reg        [15:0]   _zz_2788_;
  reg        [15:0]   _zz_2789_;
  reg        [15:0]   _zz_2790_;
  reg        [15:0]   _zz_2791_;
  reg        [15:0]   _zz_2792_;
  reg        [15:0]   _zz_2793_;
  reg        [15:0]   _zz_2794_;
  reg        [15:0]   _zz_2795_;
  reg        [15:0]   _zz_2796_;
  reg        [15:0]   _zz_2797_;
  reg        [15:0]   _zz_2798_;
  reg        [15:0]   _zz_2799_;
  reg        [15:0]   _zz_2800_;
  reg        [15:0]   _zz_2801_;
  reg        [15:0]   _zz_2802_;
  reg        [15:0]   _zz_2803_;
  reg        [15:0]   _zz_2804_;
  reg        [15:0]   _zz_2805_;
  reg        [15:0]   _zz_2806_;
  reg        [15:0]   _zz_2807_;
  reg        [15:0]   _zz_2808_;
  reg        [15:0]   _zz_2809_;
  reg        [15:0]   _zz_2810_;
  reg        [15:0]   _zz_2811_;
  reg        [15:0]   _zz_2812_;
  reg        [15:0]   _zz_2813_;
  reg        [15:0]   _zz_2814_;
  reg        [15:0]   _zz_2815_;
  reg        [15:0]   _zz_2816_;
  reg        [15:0]   _zz_2817_;
  reg        [15:0]   _zz_2818_;
  reg        [15:0]   _zz_2819_;
  reg        [15:0]   _zz_2820_;
  reg        [15:0]   _zz_2821_;
  reg        [15:0]   _zz_2822_;
  reg        [15:0]   _zz_2823_;
  reg        [15:0]   _zz_2824_;
  reg        [15:0]   _zz_2825_;
  reg        [15:0]   _zz_2826_;
  reg        [15:0]   _zz_2827_;
  reg        [15:0]   _zz_2828_;
  reg        [15:0]   _zz_2829_;
  reg        [15:0]   _zz_2830_;
  reg        [15:0]   _zz_2831_;
  reg        [15:0]   _zz_2832_;
  reg        [15:0]   _zz_2833_;
  reg        [15:0]   _zz_2834_;
  reg        [15:0]   _zz_2835_;
  reg        [15:0]   _zz_2836_;
  reg        [15:0]   _zz_2837_;
  reg        [15:0]   _zz_2838_;
  reg        [15:0]   _zz_2839_;
  reg        [15:0]   _zz_2840_;
  reg        [15:0]   _zz_2841_;
  reg        [15:0]   _zz_2842_;
  reg        [15:0]   _zz_2843_;
  reg        [15:0]   _zz_2844_;
  reg        [15:0]   _zz_2845_;
  reg        [15:0]   _zz_2846_;
  reg        [15:0]   _zz_2847_;
  reg        [15:0]   _zz_2848_;
  reg        [15:0]   _zz_2849_;
  reg        [15:0]   _zz_2850_;
  reg        [15:0]   _zz_2851_;
  reg        [15:0]   _zz_2852_;
  wire       [11:0]   _zz_2853_;
  wire       [11:0]   _zz_2854_;
  wire       [11:0]   _zz_2855_;
  wire       [0:0]    _zz_2856_;
  wire       [31:0]   _zz_2857_;
  wire       [31:0]   _zz_2858_;
  wire       [31:0]   _zz_2859_;
  wire       [31:0]   _zz_2860_;
  wire       [31:0]   _zz_2861_;
  wire       [31:0]   _zz_2862_;
  wire       [31:0]   _zz_2863_;
  wire       [31:0]   _zz_2864_;
  wire       [31:0]   _zz_2865_;
  wire       [31:0]   _zz_2866_;
  wire       [31:0]   _zz_2867_;
  wire       [31:0]   _zz_2868_;
  wire       [31:0]   _zz_2869_;
  wire       [31:0]   _zz_2870_;
  wire       [31:0]   _zz_2871_;
  wire       [31:0]   _zz_2872_;
  wire       [31:0]   _zz_2873_;
  wire       [31:0]   _zz_2874_;
  wire       [31:0]   _zz_2875_;
  wire       [31:0]   _zz_2876_;
  wire       [31:0]   _zz_2877_;
  wire       [31:0]   _zz_2878_;
  wire       [31:0]   _zz_2879_;
  wire       [31:0]   _zz_2880_;
  wire       [31:0]   _zz_2881_;
  wire       [31:0]   _zz_2882_;
  wire       [31:0]   _zz_2883_;
  wire       [31:0]   _zz_2884_;
  wire       [31:0]   _zz_2885_;
  wire       [31:0]   _zz_2886_;
  wire       [31:0]   _zz_2887_;
  wire       [31:0]   _zz_2888_;
  wire       [31:0]   _zz_2889_;
  wire       [31:0]   _zz_2890_;
  wire       [31:0]   _zz_2891_;
  wire       [31:0]   _zz_2892_;
  wire       [31:0]   _zz_2893_;
  wire       [31:0]   _zz_2894_;
  wire       [31:0]   _zz_2895_;
  wire       [31:0]   _zz_2896_;
  wire       [31:0]   _zz_2897_;
  wire       [31:0]   _zz_2898_;
  wire       [31:0]   _zz_2899_;
  wire       [31:0]   _zz_2900_;
  wire       [31:0]   _zz_2901_;
  wire       [31:0]   _zz_2902_;
  wire       [31:0]   _zz_2903_;
  wire       [31:0]   _zz_2904_;
  wire       [31:0]   _zz_2905_;
  wire       [31:0]   _zz_2906_;
  reg        [31:0]   aw_area_awaddr_r;
  reg        [7:0]    aw_area_awlen_r;
  reg        [2:0]    aw_area_awsize_r;
  reg        [3:0]    aw_area_awid_r;
  reg                 transfer_done;
  reg        [15:0]   int_reg_array_40_0_real;
  reg        [15:0]   int_reg_array_40_0_imag;
  reg        [15:0]   int_reg_array_40_1_real;
  reg        [15:0]   int_reg_array_40_1_imag;
  reg        [15:0]   int_reg_array_40_2_real;
  reg        [15:0]   int_reg_array_40_2_imag;
  reg        [15:0]   int_reg_array_40_3_real;
  reg        [15:0]   int_reg_array_40_3_imag;
  reg        [15:0]   int_reg_array_40_4_real;
  reg        [15:0]   int_reg_array_40_4_imag;
  reg        [15:0]   int_reg_array_40_5_real;
  reg        [15:0]   int_reg_array_40_5_imag;
  reg        [15:0]   int_reg_array_40_6_real;
  reg        [15:0]   int_reg_array_40_6_imag;
  reg        [15:0]   int_reg_array_40_7_real;
  reg        [15:0]   int_reg_array_40_7_imag;
  reg        [15:0]   int_reg_array_40_8_real;
  reg        [15:0]   int_reg_array_40_8_imag;
  reg        [15:0]   int_reg_array_40_9_real;
  reg        [15:0]   int_reg_array_40_9_imag;
  reg        [15:0]   int_reg_array_40_10_real;
  reg        [15:0]   int_reg_array_40_10_imag;
  reg        [15:0]   int_reg_array_40_11_real;
  reg        [15:0]   int_reg_array_40_11_imag;
  reg        [15:0]   int_reg_array_40_12_real;
  reg        [15:0]   int_reg_array_40_12_imag;
  reg        [15:0]   int_reg_array_40_13_real;
  reg        [15:0]   int_reg_array_40_13_imag;
  reg        [15:0]   int_reg_array_40_14_real;
  reg        [15:0]   int_reg_array_40_14_imag;
  reg        [15:0]   int_reg_array_40_15_real;
  reg        [15:0]   int_reg_array_40_15_imag;
  reg        [15:0]   int_reg_array_40_16_real;
  reg        [15:0]   int_reg_array_40_16_imag;
  reg        [15:0]   int_reg_array_40_17_real;
  reg        [15:0]   int_reg_array_40_17_imag;
  reg        [15:0]   int_reg_array_40_18_real;
  reg        [15:0]   int_reg_array_40_18_imag;
  reg        [15:0]   int_reg_array_40_19_real;
  reg        [15:0]   int_reg_array_40_19_imag;
  reg        [15:0]   int_reg_array_40_20_real;
  reg        [15:0]   int_reg_array_40_20_imag;
  reg        [15:0]   int_reg_array_40_21_real;
  reg        [15:0]   int_reg_array_40_21_imag;
  reg        [15:0]   int_reg_array_40_22_real;
  reg        [15:0]   int_reg_array_40_22_imag;
  reg        [15:0]   int_reg_array_40_23_real;
  reg        [15:0]   int_reg_array_40_23_imag;
  reg        [15:0]   int_reg_array_40_24_real;
  reg        [15:0]   int_reg_array_40_24_imag;
  reg        [15:0]   int_reg_array_40_25_real;
  reg        [15:0]   int_reg_array_40_25_imag;
  reg        [15:0]   int_reg_array_40_26_real;
  reg        [15:0]   int_reg_array_40_26_imag;
  reg        [15:0]   int_reg_array_40_27_real;
  reg        [15:0]   int_reg_array_40_27_imag;
  reg        [15:0]   int_reg_array_40_28_real;
  reg        [15:0]   int_reg_array_40_28_imag;
  reg        [15:0]   int_reg_array_40_29_real;
  reg        [15:0]   int_reg_array_40_29_imag;
  reg        [15:0]   int_reg_array_40_30_real;
  reg        [15:0]   int_reg_array_40_30_imag;
  reg        [15:0]   int_reg_array_40_31_real;
  reg        [15:0]   int_reg_array_40_31_imag;
  reg        [15:0]   int_reg_array_40_32_real;
  reg        [15:0]   int_reg_array_40_32_imag;
  reg        [15:0]   int_reg_array_40_33_real;
  reg        [15:0]   int_reg_array_40_33_imag;
  reg        [15:0]   int_reg_array_40_34_real;
  reg        [15:0]   int_reg_array_40_34_imag;
  reg        [15:0]   int_reg_array_40_35_real;
  reg        [15:0]   int_reg_array_40_35_imag;
  reg        [15:0]   int_reg_array_40_36_real;
  reg        [15:0]   int_reg_array_40_36_imag;
  reg        [15:0]   int_reg_array_40_37_real;
  reg        [15:0]   int_reg_array_40_37_imag;
  reg        [15:0]   int_reg_array_40_38_real;
  reg        [15:0]   int_reg_array_40_38_imag;
  reg        [15:0]   int_reg_array_40_39_real;
  reg        [15:0]   int_reg_array_40_39_imag;
  reg        [15:0]   int_reg_array_40_40_real;
  reg        [15:0]   int_reg_array_40_40_imag;
  reg        [15:0]   int_reg_array_40_41_real;
  reg        [15:0]   int_reg_array_40_41_imag;
  reg        [15:0]   int_reg_array_40_42_real;
  reg        [15:0]   int_reg_array_40_42_imag;
  reg        [15:0]   int_reg_array_40_43_real;
  reg        [15:0]   int_reg_array_40_43_imag;
  reg        [15:0]   int_reg_array_40_44_real;
  reg        [15:0]   int_reg_array_40_44_imag;
  reg        [15:0]   int_reg_array_40_45_real;
  reg        [15:0]   int_reg_array_40_45_imag;
  reg        [15:0]   int_reg_array_40_46_real;
  reg        [15:0]   int_reg_array_40_46_imag;
  reg        [15:0]   int_reg_array_40_47_real;
  reg        [15:0]   int_reg_array_40_47_imag;
  reg        [15:0]   int_reg_array_40_48_real;
  reg        [15:0]   int_reg_array_40_48_imag;
  reg        [15:0]   int_reg_array_40_49_real;
  reg        [15:0]   int_reg_array_40_49_imag;
  reg        [15:0]   int_reg_array_37_0_real;
  reg        [15:0]   int_reg_array_37_0_imag;
  reg        [15:0]   int_reg_array_37_1_real;
  reg        [15:0]   int_reg_array_37_1_imag;
  reg        [15:0]   int_reg_array_37_2_real;
  reg        [15:0]   int_reg_array_37_2_imag;
  reg        [15:0]   int_reg_array_37_3_real;
  reg        [15:0]   int_reg_array_37_3_imag;
  reg        [15:0]   int_reg_array_37_4_real;
  reg        [15:0]   int_reg_array_37_4_imag;
  reg        [15:0]   int_reg_array_37_5_real;
  reg        [15:0]   int_reg_array_37_5_imag;
  reg        [15:0]   int_reg_array_37_6_real;
  reg        [15:0]   int_reg_array_37_6_imag;
  reg        [15:0]   int_reg_array_37_7_real;
  reg        [15:0]   int_reg_array_37_7_imag;
  reg        [15:0]   int_reg_array_37_8_real;
  reg        [15:0]   int_reg_array_37_8_imag;
  reg        [15:0]   int_reg_array_37_9_real;
  reg        [15:0]   int_reg_array_37_9_imag;
  reg        [15:0]   int_reg_array_37_10_real;
  reg        [15:0]   int_reg_array_37_10_imag;
  reg        [15:0]   int_reg_array_37_11_real;
  reg        [15:0]   int_reg_array_37_11_imag;
  reg        [15:0]   int_reg_array_37_12_real;
  reg        [15:0]   int_reg_array_37_12_imag;
  reg        [15:0]   int_reg_array_37_13_real;
  reg        [15:0]   int_reg_array_37_13_imag;
  reg        [15:0]   int_reg_array_37_14_real;
  reg        [15:0]   int_reg_array_37_14_imag;
  reg        [15:0]   int_reg_array_37_15_real;
  reg        [15:0]   int_reg_array_37_15_imag;
  reg        [15:0]   int_reg_array_37_16_real;
  reg        [15:0]   int_reg_array_37_16_imag;
  reg        [15:0]   int_reg_array_37_17_real;
  reg        [15:0]   int_reg_array_37_17_imag;
  reg        [15:0]   int_reg_array_37_18_real;
  reg        [15:0]   int_reg_array_37_18_imag;
  reg        [15:0]   int_reg_array_37_19_real;
  reg        [15:0]   int_reg_array_37_19_imag;
  reg        [15:0]   int_reg_array_37_20_real;
  reg        [15:0]   int_reg_array_37_20_imag;
  reg        [15:0]   int_reg_array_37_21_real;
  reg        [15:0]   int_reg_array_37_21_imag;
  reg        [15:0]   int_reg_array_37_22_real;
  reg        [15:0]   int_reg_array_37_22_imag;
  reg        [15:0]   int_reg_array_37_23_real;
  reg        [15:0]   int_reg_array_37_23_imag;
  reg        [15:0]   int_reg_array_37_24_real;
  reg        [15:0]   int_reg_array_37_24_imag;
  reg        [15:0]   int_reg_array_37_25_real;
  reg        [15:0]   int_reg_array_37_25_imag;
  reg        [15:0]   int_reg_array_37_26_real;
  reg        [15:0]   int_reg_array_37_26_imag;
  reg        [15:0]   int_reg_array_37_27_real;
  reg        [15:0]   int_reg_array_37_27_imag;
  reg        [15:0]   int_reg_array_37_28_real;
  reg        [15:0]   int_reg_array_37_28_imag;
  reg        [15:0]   int_reg_array_37_29_real;
  reg        [15:0]   int_reg_array_37_29_imag;
  reg        [15:0]   int_reg_array_37_30_real;
  reg        [15:0]   int_reg_array_37_30_imag;
  reg        [15:0]   int_reg_array_37_31_real;
  reg        [15:0]   int_reg_array_37_31_imag;
  reg        [15:0]   int_reg_array_37_32_real;
  reg        [15:0]   int_reg_array_37_32_imag;
  reg        [15:0]   int_reg_array_37_33_real;
  reg        [15:0]   int_reg_array_37_33_imag;
  reg        [15:0]   int_reg_array_37_34_real;
  reg        [15:0]   int_reg_array_37_34_imag;
  reg        [15:0]   int_reg_array_37_35_real;
  reg        [15:0]   int_reg_array_37_35_imag;
  reg        [15:0]   int_reg_array_37_36_real;
  reg        [15:0]   int_reg_array_37_36_imag;
  reg        [15:0]   int_reg_array_37_37_real;
  reg        [15:0]   int_reg_array_37_37_imag;
  reg        [15:0]   int_reg_array_37_38_real;
  reg        [15:0]   int_reg_array_37_38_imag;
  reg        [15:0]   int_reg_array_37_39_real;
  reg        [15:0]   int_reg_array_37_39_imag;
  reg        [15:0]   int_reg_array_37_40_real;
  reg        [15:0]   int_reg_array_37_40_imag;
  reg        [15:0]   int_reg_array_37_41_real;
  reg        [15:0]   int_reg_array_37_41_imag;
  reg        [15:0]   int_reg_array_37_42_real;
  reg        [15:0]   int_reg_array_37_42_imag;
  reg        [15:0]   int_reg_array_37_43_real;
  reg        [15:0]   int_reg_array_37_43_imag;
  reg        [15:0]   int_reg_array_37_44_real;
  reg        [15:0]   int_reg_array_37_44_imag;
  reg        [15:0]   int_reg_array_37_45_real;
  reg        [15:0]   int_reg_array_37_45_imag;
  reg        [15:0]   int_reg_array_37_46_real;
  reg        [15:0]   int_reg_array_37_46_imag;
  reg        [15:0]   int_reg_array_37_47_real;
  reg        [15:0]   int_reg_array_37_47_imag;
  reg        [15:0]   int_reg_array_37_48_real;
  reg        [15:0]   int_reg_array_37_48_imag;
  reg        [15:0]   int_reg_array_37_49_real;
  reg        [15:0]   int_reg_array_37_49_imag;
  reg        [15:0]   int_reg_array_0_0_real;
  reg        [15:0]   int_reg_array_0_0_imag;
  reg        [15:0]   int_reg_array_0_1_real;
  reg        [15:0]   int_reg_array_0_1_imag;
  reg        [15:0]   int_reg_array_0_2_real;
  reg        [15:0]   int_reg_array_0_2_imag;
  reg        [15:0]   int_reg_array_0_3_real;
  reg        [15:0]   int_reg_array_0_3_imag;
  reg        [15:0]   int_reg_array_0_4_real;
  reg        [15:0]   int_reg_array_0_4_imag;
  reg        [15:0]   int_reg_array_0_5_real;
  reg        [15:0]   int_reg_array_0_5_imag;
  reg        [15:0]   int_reg_array_0_6_real;
  reg        [15:0]   int_reg_array_0_6_imag;
  reg        [15:0]   int_reg_array_0_7_real;
  reg        [15:0]   int_reg_array_0_7_imag;
  reg        [15:0]   int_reg_array_0_8_real;
  reg        [15:0]   int_reg_array_0_8_imag;
  reg        [15:0]   int_reg_array_0_9_real;
  reg        [15:0]   int_reg_array_0_9_imag;
  reg        [15:0]   int_reg_array_0_10_real;
  reg        [15:0]   int_reg_array_0_10_imag;
  reg        [15:0]   int_reg_array_0_11_real;
  reg        [15:0]   int_reg_array_0_11_imag;
  reg        [15:0]   int_reg_array_0_12_real;
  reg        [15:0]   int_reg_array_0_12_imag;
  reg        [15:0]   int_reg_array_0_13_real;
  reg        [15:0]   int_reg_array_0_13_imag;
  reg        [15:0]   int_reg_array_0_14_real;
  reg        [15:0]   int_reg_array_0_14_imag;
  reg        [15:0]   int_reg_array_0_15_real;
  reg        [15:0]   int_reg_array_0_15_imag;
  reg        [15:0]   int_reg_array_0_16_real;
  reg        [15:0]   int_reg_array_0_16_imag;
  reg        [15:0]   int_reg_array_0_17_real;
  reg        [15:0]   int_reg_array_0_17_imag;
  reg        [15:0]   int_reg_array_0_18_real;
  reg        [15:0]   int_reg_array_0_18_imag;
  reg        [15:0]   int_reg_array_0_19_real;
  reg        [15:0]   int_reg_array_0_19_imag;
  reg        [15:0]   int_reg_array_0_20_real;
  reg        [15:0]   int_reg_array_0_20_imag;
  reg        [15:0]   int_reg_array_0_21_real;
  reg        [15:0]   int_reg_array_0_21_imag;
  reg        [15:0]   int_reg_array_0_22_real;
  reg        [15:0]   int_reg_array_0_22_imag;
  reg        [15:0]   int_reg_array_0_23_real;
  reg        [15:0]   int_reg_array_0_23_imag;
  reg        [15:0]   int_reg_array_0_24_real;
  reg        [15:0]   int_reg_array_0_24_imag;
  reg        [15:0]   int_reg_array_0_25_real;
  reg        [15:0]   int_reg_array_0_25_imag;
  reg        [15:0]   int_reg_array_0_26_real;
  reg        [15:0]   int_reg_array_0_26_imag;
  reg        [15:0]   int_reg_array_0_27_real;
  reg        [15:0]   int_reg_array_0_27_imag;
  reg        [15:0]   int_reg_array_0_28_real;
  reg        [15:0]   int_reg_array_0_28_imag;
  reg        [15:0]   int_reg_array_0_29_real;
  reg        [15:0]   int_reg_array_0_29_imag;
  reg        [15:0]   int_reg_array_0_30_real;
  reg        [15:0]   int_reg_array_0_30_imag;
  reg        [15:0]   int_reg_array_0_31_real;
  reg        [15:0]   int_reg_array_0_31_imag;
  reg        [15:0]   int_reg_array_0_32_real;
  reg        [15:0]   int_reg_array_0_32_imag;
  reg        [15:0]   int_reg_array_0_33_real;
  reg        [15:0]   int_reg_array_0_33_imag;
  reg        [15:0]   int_reg_array_0_34_real;
  reg        [15:0]   int_reg_array_0_34_imag;
  reg        [15:0]   int_reg_array_0_35_real;
  reg        [15:0]   int_reg_array_0_35_imag;
  reg        [15:0]   int_reg_array_0_36_real;
  reg        [15:0]   int_reg_array_0_36_imag;
  reg        [15:0]   int_reg_array_0_37_real;
  reg        [15:0]   int_reg_array_0_37_imag;
  reg        [15:0]   int_reg_array_0_38_real;
  reg        [15:0]   int_reg_array_0_38_imag;
  reg        [15:0]   int_reg_array_0_39_real;
  reg        [15:0]   int_reg_array_0_39_imag;
  reg        [15:0]   int_reg_array_0_40_real;
  reg        [15:0]   int_reg_array_0_40_imag;
  reg        [15:0]   int_reg_array_0_41_real;
  reg        [15:0]   int_reg_array_0_41_imag;
  reg        [15:0]   int_reg_array_0_42_real;
  reg        [15:0]   int_reg_array_0_42_imag;
  reg        [15:0]   int_reg_array_0_43_real;
  reg        [15:0]   int_reg_array_0_43_imag;
  reg        [15:0]   int_reg_array_0_44_real;
  reg        [15:0]   int_reg_array_0_44_imag;
  reg        [15:0]   int_reg_array_0_45_real;
  reg        [15:0]   int_reg_array_0_45_imag;
  reg        [15:0]   int_reg_array_0_46_real;
  reg        [15:0]   int_reg_array_0_46_imag;
  reg        [15:0]   int_reg_array_0_47_real;
  reg        [15:0]   int_reg_array_0_47_imag;
  reg        [15:0]   int_reg_array_0_48_real;
  reg        [15:0]   int_reg_array_0_48_imag;
  reg        [15:0]   int_reg_array_0_49_real;
  reg        [15:0]   int_reg_array_0_49_imag;
  reg        [15:0]   int_reg_array_26_0_real;
  reg        [15:0]   int_reg_array_26_0_imag;
  reg        [15:0]   int_reg_array_26_1_real;
  reg        [15:0]   int_reg_array_26_1_imag;
  reg        [15:0]   int_reg_array_26_2_real;
  reg        [15:0]   int_reg_array_26_2_imag;
  reg        [15:0]   int_reg_array_26_3_real;
  reg        [15:0]   int_reg_array_26_3_imag;
  reg        [15:0]   int_reg_array_26_4_real;
  reg        [15:0]   int_reg_array_26_4_imag;
  reg        [15:0]   int_reg_array_26_5_real;
  reg        [15:0]   int_reg_array_26_5_imag;
  reg        [15:0]   int_reg_array_26_6_real;
  reg        [15:0]   int_reg_array_26_6_imag;
  reg        [15:0]   int_reg_array_26_7_real;
  reg        [15:0]   int_reg_array_26_7_imag;
  reg        [15:0]   int_reg_array_26_8_real;
  reg        [15:0]   int_reg_array_26_8_imag;
  reg        [15:0]   int_reg_array_26_9_real;
  reg        [15:0]   int_reg_array_26_9_imag;
  reg        [15:0]   int_reg_array_26_10_real;
  reg        [15:0]   int_reg_array_26_10_imag;
  reg        [15:0]   int_reg_array_26_11_real;
  reg        [15:0]   int_reg_array_26_11_imag;
  reg        [15:0]   int_reg_array_26_12_real;
  reg        [15:0]   int_reg_array_26_12_imag;
  reg        [15:0]   int_reg_array_26_13_real;
  reg        [15:0]   int_reg_array_26_13_imag;
  reg        [15:0]   int_reg_array_26_14_real;
  reg        [15:0]   int_reg_array_26_14_imag;
  reg        [15:0]   int_reg_array_26_15_real;
  reg        [15:0]   int_reg_array_26_15_imag;
  reg        [15:0]   int_reg_array_26_16_real;
  reg        [15:0]   int_reg_array_26_16_imag;
  reg        [15:0]   int_reg_array_26_17_real;
  reg        [15:0]   int_reg_array_26_17_imag;
  reg        [15:0]   int_reg_array_26_18_real;
  reg        [15:0]   int_reg_array_26_18_imag;
  reg        [15:0]   int_reg_array_26_19_real;
  reg        [15:0]   int_reg_array_26_19_imag;
  reg        [15:0]   int_reg_array_26_20_real;
  reg        [15:0]   int_reg_array_26_20_imag;
  reg        [15:0]   int_reg_array_26_21_real;
  reg        [15:0]   int_reg_array_26_21_imag;
  reg        [15:0]   int_reg_array_26_22_real;
  reg        [15:0]   int_reg_array_26_22_imag;
  reg        [15:0]   int_reg_array_26_23_real;
  reg        [15:0]   int_reg_array_26_23_imag;
  reg        [15:0]   int_reg_array_26_24_real;
  reg        [15:0]   int_reg_array_26_24_imag;
  reg        [15:0]   int_reg_array_26_25_real;
  reg        [15:0]   int_reg_array_26_25_imag;
  reg        [15:0]   int_reg_array_26_26_real;
  reg        [15:0]   int_reg_array_26_26_imag;
  reg        [15:0]   int_reg_array_26_27_real;
  reg        [15:0]   int_reg_array_26_27_imag;
  reg        [15:0]   int_reg_array_26_28_real;
  reg        [15:0]   int_reg_array_26_28_imag;
  reg        [15:0]   int_reg_array_26_29_real;
  reg        [15:0]   int_reg_array_26_29_imag;
  reg        [15:0]   int_reg_array_26_30_real;
  reg        [15:0]   int_reg_array_26_30_imag;
  reg        [15:0]   int_reg_array_26_31_real;
  reg        [15:0]   int_reg_array_26_31_imag;
  reg        [15:0]   int_reg_array_26_32_real;
  reg        [15:0]   int_reg_array_26_32_imag;
  reg        [15:0]   int_reg_array_26_33_real;
  reg        [15:0]   int_reg_array_26_33_imag;
  reg        [15:0]   int_reg_array_26_34_real;
  reg        [15:0]   int_reg_array_26_34_imag;
  reg        [15:0]   int_reg_array_26_35_real;
  reg        [15:0]   int_reg_array_26_35_imag;
  reg        [15:0]   int_reg_array_26_36_real;
  reg        [15:0]   int_reg_array_26_36_imag;
  reg        [15:0]   int_reg_array_26_37_real;
  reg        [15:0]   int_reg_array_26_37_imag;
  reg        [15:0]   int_reg_array_26_38_real;
  reg        [15:0]   int_reg_array_26_38_imag;
  reg        [15:0]   int_reg_array_26_39_real;
  reg        [15:0]   int_reg_array_26_39_imag;
  reg        [15:0]   int_reg_array_26_40_real;
  reg        [15:0]   int_reg_array_26_40_imag;
  reg        [15:0]   int_reg_array_26_41_real;
  reg        [15:0]   int_reg_array_26_41_imag;
  reg        [15:0]   int_reg_array_26_42_real;
  reg        [15:0]   int_reg_array_26_42_imag;
  reg        [15:0]   int_reg_array_26_43_real;
  reg        [15:0]   int_reg_array_26_43_imag;
  reg        [15:0]   int_reg_array_26_44_real;
  reg        [15:0]   int_reg_array_26_44_imag;
  reg        [15:0]   int_reg_array_26_45_real;
  reg        [15:0]   int_reg_array_26_45_imag;
  reg        [15:0]   int_reg_array_26_46_real;
  reg        [15:0]   int_reg_array_26_46_imag;
  reg        [15:0]   int_reg_array_26_47_real;
  reg        [15:0]   int_reg_array_26_47_imag;
  reg        [15:0]   int_reg_array_26_48_real;
  reg        [15:0]   int_reg_array_26_48_imag;
  reg        [15:0]   int_reg_array_26_49_real;
  reg        [15:0]   int_reg_array_26_49_imag;
  reg        [15:0]   int_reg_array_36_0_real;
  reg        [15:0]   int_reg_array_36_0_imag;
  reg        [15:0]   int_reg_array_36_1_real;
  reg        [15:0]   int_reg_array_36_1_imag;
  reg        [15:0]   int_reg_array_36_2_real;
  reg        [15:0]   int_reg_array_36_2_imag;
  reg        [15:0]   int_reg_array_36_3_real;
  reg        [15:0]   int_reg_array_36_3_imag;
  reg        [15:0]   int_reg_array_36_4_real;
  reg        [15:0]   int_reg_array_36_4_imag;
  reg        [15:0]   int_reg_array_36_5_real;
  reg        [15:0]   int_reg_array_36_5_imag;
  reg        [15:0]   int_reg_array_36_6_real;
  reg        [15:0]   int_reg_array_36_6_imag;
  reg        [15:0]   int_reg_array_36_7_real;
  reg        [15:0]   int_reg_array_36_7_imag;
  reg        [15:0]   int_reg_array_36_8_real;
  reg        [15:0]   int_reg_array_36_8_imag;
  reg        [15:0]   int_reg_array_36_9_real;
  reg        [15:0]   int_reg_array_36_9_imag;
  reg        [15:0]   int_reg_array_36_10_real;
  reg        [15:0]   int_reg_array_36_10_imag;
  reg        [15:0]   int_reg_array_36_11_real;
  reg        [15:0]   int_reg_array_36_11_imag;
  reg        [15:0]   int_reg_array_36_12_real;
  reg        [15:0]   int_reg_array_36_12_imag;
  reg        [15:0]   int_reg_array_36_13_real;
  reg        [15:0]   int_reg_array_36_13_imag;
  reg        [15:0]   int_reg_array_36_14_real;
  reg        [15:0]   int_reg_array_36_14_imag;
  reg        [15:0]   int_reg_array_36_15_real;
  reg        [15:0]   int_reg_array_36_15_imag;
  reg        [15:0]   int_reg_array_36_16_real;
  reg        [15:0]   int_reg_array_36_16_imag;
  reg        [15:0]   int_reg_array_36_17_real;
  reg        [15:0]   int_reg_array_36_17_imag;
  reg        [15:0]   int_reg_array_36_18_real;
  reg        [15:0]   int_reg_array_36_18_imag;
  reg        [15:0]   int_reg_array_36_19_real;
  reg        [15:0]   int_reg_array_36_19_imag;
  reg        [15:0]   int_reg_array_36_20_real;
  reg        [15:0]   int_reg_array_36_20_imag;
  reg        [15:0]   int_reg_array_36_21_real;
  reg        [15:0]   int_reg_array_36_21_imag;
  reg        [15:0]   int_reg_array_36_22_real;
  reg        [15:0]   int_reg_array_36_22_imag;
  reg        [15:0]   int_reg_array_36_23_real;
  reg        [15:0]   int_reg_array_36_23_imag;
  reg        [15:0]   int_reg_array_36_24_real;
  reg        [15:0]   int_reg_array_36_24_imag;
  reg        [15:0]   int_reg_array_36_25_real;
  reg        [15:0]   int_reg_array_36_25_imag;
  reg        [15:0]   int_reg_array_36_26_real;
  reg        [15:0]   int_reg_array_36_26_imag;
  reg        [15:0]   int_reg_array_36_27_real;
  reg        [15:0]   int_reg_array_36_27_imag;
  reg        [15:0]   int_reg_array_36_28_real;
  reg        [15:0]   int_reg_array_36_28_imag;
  reg        [15:0]   int_reg_array_36_29_real;
  reg        [15:0]   int_reg_array_36_29_imag;
  reg        [15:0]   int_reg_array_36_30_real;
  reg        [15:0]   int_reg_array_36_30_imag;
  reg        [15:0]   int_reg_array_36_31_real;
  reg        [15:0]   int_reg_array_36_31_imag;
  reg        [15:0]   int_reg_array_36_32_real;
  reg        [15:0]   int_reg_array_36_32_imag;
  reg        [15:0]   int_reg_array_36_33_real;
  reg        [15:0]   int_reg_array_36_33_imag;
  reg        [15:0]   int_reg_array_36_34_real;
  reg        [15:0]   int_reg_array_36_34_imag;
  reg        [15:0]   int_reg_array_36_35_real;
  reg        [15:0]   int_reg_array_36_35_imag;
  reg        [15:0]   int_reg_array_36_36_real;
  reg        [15:0]   int_reg_array_36_36_imag;
  reg        [15:0]   int_reg_array_36_37_real;
  reg        [15:0]   int_reg_array_36_37_imag;
  reg        [15:0]   int_reg_array_36_38_real;
  reg        [15:0]   int_reg_array_36_38_imag;
  reg        [15:0]   int_reg_array_36_39_real;
  reg        [15:0]   int_reg_array_36_39_imag;
  reg        [15:0]   int_reg_array_36_40_real;
  reg        [15:0]   int_reg_array_36_40_imag;
  reg        [15:0]   int_reg_array_36_41_real;
  reg        [15:0]   int_reg_array_36_41_imag;
  reg        [15:0]   int_reg_array_36_42_real;
  reg        [15:0]   int_reg_array_36_42_imag;
  reg        [15:0]   int_reg_array_36_43_real;
  reg        [15:0]   int_reg_array_36_43_imag;
  reg        [15:0]   int_reg_array_36_44_real;
  reg        [15:0]   int_reg_array_36_44_imag;
  reg        [15:0]   int_reg_array_36_45_real;
  reg        [15:0]   int_reg_array_36_45_imag;
  reg        [15:0]   int_reg_array_36_46_real;
  reg        [15:0]   int_reg_array_36_46_imag;
  reg        [15:0]   int_reg_array_36_47_real;
  reg        [15:0]   int_reg_array_36_47_imag;
  reg        [15:0]   int_reg_array_36_48_real;
  reg        [15:0]   int_reg_array_36_48_imag;
  reg        [15:0]   int_reg_array_36_49_real;
  reg        [15:0]   int_reg_array_36_49_imag;
  reg        [15:0]   int_reg_array_46_0_real;
  reg        [15:0]   int_reg_array_46_0_imag;
  reg        [15:0]   int_reg_array_46_1_real;
  reg        [15:0]   int_reg_array_46_1_imag;
  reg        [15:0]   int_reg_array_46_2_real;
  reg        [15:0]   int_reg_array_46_2_imag;
  reg        [15:0]   int_reg_array_46_3_real;
  reg        [15:0]   int_reg_array_46_3_imag;
  reg        [15:0]   int_reg_array_46_4_real;
  reg        [15:0]   int_reg_array_46_4_imag;
  reg        [15:0]   int_reg_array_46_5_real;
  reg        [15:0]   int_reg_array_46_5_imag;
  reg        [15:0]   int_reg_array_46_6_real;
  reg        [15:0]   int_reg_array_46_6_imag;
  reg        [15:0]   int_reg_array_46_7_real;
  reg        [15:0]   int_reg_array_46_7_imag;
  reg        [15:0]   int_reg_array_46_8_real;
  reg        [15:0]   int_reg_array_46_8_imag;
  reg        [15:0]   int_reg_array_46_9_real;
  reg        [15:0]   int_reg_array_46_9_imag;
  reg        [15:0]   int_reg_array_46_10_real;
  reg        [15:0]   int_reg_array_46_10_imag;
  reg        [15:0]   int_reg_array_46_11_real;
  reg        [15:0]   int_reg_array_46_11_imag;
  reg        [15:0]   int_reg_array_46_12_real;
  reg        [15:0]   int_reg_array_46_12_imag;
  reg        [15:0]   int_reg_array_46_13_real;
  reg        [15:0]   int_reg_array_46_13_imag;
  reg        [15:0]   int_reg_array_46_14_real;
  reg        [15:0]   int_reg_array_46_14_imag;
  reg        [15:0]   int_reg_array_46_15_real;
  reg        [15:0]   int_reg_array_46_15_imag;
  reg        [15:0]   int_reg_array_46_16_real;
  reg        [15:0]   int_reg_array_46_16_imag;
  reg        [15:0]   int_reg_array_46_17_real;
  reg        [15:0]   int_reg_array_46_17_imag;
  reg        [15:0]   int_reg_array_46_18_real;
  reg        [15:0]   int_reg_array_46_18_imag;
  reg        [15:0]   int_reg_array_46_19_real;
  reg        [15:0]   int_reg_array_46_19_imag;
  reg        [15:0]   int_reg_array_46_20_real;
  reg        [15:0]   int_reg_array_46_20_imag;
  reg        [15:0]   int_reg_array_46_21_real;
  reg        [15:0]   int_reg_array_46_21_imag;
  reg        [15:0]   int_reg_array_46_22_real;
  reg        [15:0]   int_reg_array_46_22_imag;
  reg        [15:0]   int_reg_array_46_23_real;
  reg        [15:0]   int_reg_array_46_23_imag;
  reg        [15:0]   int_reg_array_46_24_real;
  reg        [15:0]   int_reg_array_46_24_imag;
  reg        [15:0]   int_reg_array_46_25_real;
  reg        [15:0]   int_reg_array_46_25_imag;
  reg        [15:0]   int_reg_array_46_26_real;
  reg        [15:0]   int_reg_array_46_26_imag;
  reg        [15:0]   int_reg_array_46_27_real;
  reg        [15:0]   int_reg_array_46_27_imag;
  reg        [15:0]   int_reg_array_46_28_real;
  reg        [15:0]   int_reg_array_46_28_imag;
  reg        [15:0]   int_reg_array_46_29_real;
  reg        [15:0]   int_reg_array_46_29_imag;
  reg        [15:0]   int_reg_array_46_30_real;
  reg        [15:0]   int_reg_array_46_30_imag;
  reg        [15:0]   int_reg_array_46_31_real;
  reg        [15:0]   int_reg_array_46_31_imag;
  reg        [15:0]   int_reg_array_46_32_real;
  reg        [15:0]   int_reg_array_46_32_imag;
  reg        [15:0]   int_reg_array_46_33_real;
  reg        [15:0]   int_reg_array_46_33_imag;
  reg        [15:0]   int_reg_array_46_34_real;
  reg        [15:0]   int_reg_array_46_34_imag;
  reg        [15:0]   int_reg_array_46_35_real;
  reg        [15:0]   int_reg_array_46_35_imag;
  reg        [15:0]   int_reg_array_46_36_real;
  reg        [15:0]   int_reg_array_46_36_imag;
  reg        [15:0]   int_reg_array_46_37_real;
  reg        [15:0]   int_reg_array_46_37_imag;
  reg        [15:0]   int_reg_array_46_38_real;
  reg        [15:0]   int_reg_array_46_38_imag;
  reg        [15:0]   int_reg_array_46_39_real;
  reg        [15:0]   int_reg_array_46_39_imag;
  reg        [15:0]   int_reg_array_46_40_real;
  reg        [15:0]   int_reg_array_46_40_imag;
  reg        [15:0]   int_reg_array_46_41_real;
  reg        [15:0]   int_reg_array_46_41_imag;
  reg        [15:0]   int_reg_array_46_42_real;
  reg        [15:0]   int_reg_array_46_42_imag;
  reg        [15:0]   int_reg_array_46_43_real;
  reg        [15:0]   int_reg_array_46_43_imag;
  reg        [15:0]   int_reg_array_46_44_real;
  reg        [15:0]   int_reg_array_46_44_imag;
  reg        [15:0]   int_reg_array_46_45_real;
  reg        [15:0]   int_reg_array_46_45_imag;
  reg        [15:0]   int_reg_array_46_46_real;
  reg        [15:0]   int_reg_array_46_46_imag;
  reg        [15:0]   int_reg_array_46_47_real;
  reg        [15:0]   int_reg_array_46_47_imag;
  reg        [15:0]   int_reg_array_46_48_real;
  reg        [15:0]   int_reg_array_46_48_imag;
  reg        [15:0]   int_reg_array_46_49_real;
  reg        [15:0]   int_reg_array_46_49_imag;
  reg        [15:0]   int_reg_array_49_0_real;
  reg        [15:0]   int_reg_array_49_0_imag;
  reg        [15:0]   int_reg_array_49_1_real;
  reg        [15:0]   int_reg_array_49_1_imag;
  reg        [15:0]   int_reg_array_49_2_real;
  reg        [15:0]   int_reg_array_49_2_imag;
  reg        [15:0]   int_reg_array_49_3_real;
  reg        [15:0]   int_reg_array_49_3_imag;
  reg        [15:0]   int_reg_array_49_4_real;
  reg        [15:0]   int_reg_array_49_4_imag;
  reg        [15:0]   int_reg_array_49_5_real;
  reg        [15:0]   int_reg_array_49_5_imag;
  reg        [15:0]   int_reg_array_49_6_real;
  reg        [15:0]   int_reg_array_49_6_imag;
  reg        [15:0]   int_reg_array_49_7_real;
  reg        [15:0]   int_reg_array_49_7_imag;
  reg        [15:0]   int_reg_array_49_8_real;
  reg        [15:0]   int_reg_array_49_8_imag;
  reg        [15:0]   int_reg_array_49_9_real;
  reg        [15:0]   int_reg_array_49_9_imag;
  reg        [15:0]   int_reg_array_49_10_real;
  reg        [15:0]   int_reg_array_49_10_imag;
  reg        [15:0]   int_reg_array_49_11_real;
  reg        [15:0]   int_reg_array_49_11_imag;
  reg        [15:0]   int_reg_array_49_12_real;
  reg        [15:0]   int_reg_array_49_12_imag;
  reg        [15:0]   int_reg_array_49_13_real;
  reg        [15:0]   int_reg_array_49_13_imag;
  reg        [15:0]   int_reg_array_49_14_real;
  reg        [15:0]   int_reg_array_49_14_imag;
  reg        [15:0]   int_reg_array_49_15_real;
  reg        [15:0]   int_reg_array_49_15_imag;
  reg        [15:0]   int_reg_array_49_16_real;
  reg        [15:0]   int_reg_array_49_16_imag;
  reg        [15:0]   int_reg_array_49_17_real;
  reg        [15:0]   int_reg_array_49_17_imag;
  reg        [15:0]   int_reg_array_49_18_real;
  reg        [15:0]   int_reg_array_49_18_imag;
  reg        [15:0]   int_reg_array_49_19_real;
  reg        [15:0]   int_reg_array_49_19_imag;
  reg        [15:0]   int_reg_array_49_20_real;
  reg        [15:0]   int_reg_array_49_20_imag;
  reg        [15:0]   int_reg_array_49_21_real;
  reg        [15:0]   int_reg_array_49_21_imag;
  reg        [15:0]   int_reg_array_49_22_real;
  reg        [15:0]   int_reg_array_49_22_imag;
  reg        [15:0]   int_reg_array_49_23_real;
  reg        [15:0]   int_reg_array_49_23_imag;
  reg        [15:0]   int_reg_array_49_24_real;
  reg        [15:0]   int_reg_array_49_24_imag;
  reg        [15:0]   int_reg_array_49_25_real;
  reg        [15:0]   int_reg_array_49_25_imag;
  reg        [15:0]   int_reg_array_49_26_real;
  reg        [15:0]   int_reg_array_49_26_imag;
  reg        [15:0]   int_reg_array_49_27_real;
  reg        [15:0]   int_reg_array_49_27_imag;
  reg        [15:0]   int_reg_array_49_28_real;
  reg        [15:0]   int_reg_array_49_28_imag;
  reg        [15:0]   int_reg_array_49_29_real;
  reg        [15:0]   int_reg_array_49_29_imag;
  reg        [15:0]   int_reg_array_49_30_real;
  reg        [15:0]   int_reg_array_49_30_imag;
  reg        [15:0]   int_reg_array_49_31_real;
  reg        [15:0]   int_reg_array_49_31_imag;
  reg        [15:0]   int_reg_array_49_32_real;
  reg        [15:0]   int_reg_array_49_32_imag;
  reg        [15:0]   int_reg_array_49_33_real;
  reg        [15:0]   int_reg_array_49_33_imag;
  reg        [15:0]   int_reg_array_49_34_real;
  reg        [15:0]   int_reg_array_49_34_imag;
  reg        [15:0]   int_reg_array_49_35_real;
  reg        [15:0]   int_reg_array_49_35_imag;
  reg        [15:0]   int_reg_array_49_36_real;
  reg        [15:0]   int_reg_array_49_36_imag;
  reg        [15:0]   int_reg_array_49_37_real;
  reg        [15:0]   int_reg_array_49_37_imag;
  reg        [15:0]   int_reg_array_49_38_real;
  reg        [15:0]   int_reg_array_49_38_imag;
  reg        [15:0]   int_reg_array_49_39_real;
  reg        [15:0]   int_reg_array_49_39_imag;
  reg        [15:0]   int_reg_array_49_40_real;
  reg        [15:0]   int_reg_array_49_40_imag;
  reg        [15:0]   int_reg_array_49_41_real;
  reg        [15:0]   int_reg_array_49_41_imag;
  reg        [15:0]   int_reg_array_49_42_real;
  reg        [15:0]   int_reg_array_49_42_imag;
  reg        [15:0]   int_reg_array_49_43_real;
  reg        [15:0]   int_reg_array_49_43_imag;
  reg        [15:0]   int_reg_array_49_44_real;
  reg        [15:0]   int_reg_array_49_44_imag;
  reg        [15:0]   int_reg_array_49_45_real;
  reg        [15:0]   int_reg_array_49_45_imag;
  reg        [15:0]   int_reg_array_49_46_real;
  reg        [15:0]   int_reg_array_49_46_imag;
  reg        [15:0]   int_reg_array_49_47_real;
  reg        [15:0]   int_reg_array_49_47_imag;
  reg        [15:0]   int_reg_array_49_48_real;
  reg        [15:0]   int_reg_array_49_48_imag;
  reg        [15:0]   int_reg_array_49_49_real;
  reg        [15:0]   int_reg_array_49_49_imag;
  reg        [15:0]   int_reg_array_28_0_real;
  reg        [15:0]   int_reg_array_28_0_imag;
  reg        [15:0]   int_reg_array_28_1_real;
  reg        [15:0]   int_reg_array_28_1_imag;
  reg        [15:0]   int_reg_array_28_2_real;
  reg        [15:0]   int_reg_array_28_2_imag;
  reg        [15:0]   int_reg_array_28_3_real;
  reg        [15:0]   int_reg_array_28_3_imag;
  reg        [15:0]   int_reg_array_28_4_real;
  reg        [15:0]   int_reg_array_28_4_imag;
  reg        [15:0]   int_reg_array_28_5_real;
  reg        [15:0]   int_reg_array_28_5_imag;
  reg        [15:0]   int_reg_array_28_6_real;
  reg        [15:0]   int_reg_array_28_6_imag;
  reg        [15:0]   int_reg_array_28_7_real;
  reg        [15:0]   int_reg_array_28_7_imag;
  reg        [15:0]   int_reg_array_28_8_real;
  reg        [15:0]   int_reg_array_28_8_imag;
  reg        [15:0]   int_reg_array_28_9_real;
  reg        [15:0]   int_reg_array_28_9_imag;
  reg        [15:0]   int_reg_array_28_10_real;
  reg        [15:0]   int_reg_array_28_10_imag;
  reg        [15:0]   int_reg_array_28_11_real;
  reg        [15:0]   int_reg_array_28_11_imag;
  reg        [15:0]   int_reg_array_28_12_real;
  reg        [15:0]   int_reg_array_28_12_imag;
  reg        [15:0]   int_reg_array_28_13_real;
  reg        [15:0]   int_reg_array_28_13_imag;
  reg        [15:0]   int_reg_array_28_14_real;
  reg        [15:0]   int_reg_array_28_14_imag;
  reg        [15:0]   int_reg_array_28_15_real;
  reg        [15:0]   int_reg_array_28_15_imag;
  reg        [15:0]   int_reg_array_28_16_real;
  reg        [15:0]   int_reg_array_28_16_imag;
  reg        [15:0]   int_reg_array_28_17_real;
  reg        [15:0]   int_reg_array_28_17_imag;
  reg        [15:0]   int_reg_array_28_18_real;
  reg        [15:0]   int_reg_array_28_18_imag;
  reg        [15:0]   int_reg_array_28_19_real;
  reg        [15:0]   int_reg_array_28_19_imag;
  reg        [15:0]   int_reg_array_28_20_real;
  reg        [15:0]   int_reg_array_28_20_imag;
  reg        [15:0]   int_reg_array_28_21_real;
  reg        [15:0]   int_reg_array_28_21_imag;
  reg        [15:0]   int_reg_array_28_22_real;
  reg        [15:0]   int_reg_array_28_22_imag;
  reg        [15:0]   int_reg_array_28_23_real;
  reg        [15:0]   int_reg_array_28_23_imag;
  reg        [15:0]   int_reg_array_28_24_real;
  reg        [15:0]   int_reg_array_28_24_imag;
  reg        [15:0]   int_reg_array_28_25_real;
  reg        [15:0]   int_reg_array_28_25_imag;
  reg        [15:0]   int_reg_array_28_26_real;
  reg        [15:0]   int_reg_array_28_26_imag;
  reg        [15:0]   int_reg_array_28_27_real;
  reg        [15:0]   int_reg_array_28_27_imag;
  reg        [15:0]   int_reg_array_28_28_real;
  reg        [15:0]   int_reg_array_28_28_imag;
  reg        [15:0]   int_reg_array_28_29_real;
  reg        [15:0]   int_reg_array_28_29_imag;
  reg        [15:0]   int_reg_array_28_30_real;
  reg        [15:0]   int_reg_array_28_30_imag;
  reg        [15:0]   int_reg_array_28_31_real;
  reg        [15:0]   int_reg_array_28_31_imag;
  reg        [15:0]   int_reg_array_28_32_real;
  reg        [15:0]   int_reg_array_28_32_imag;
  reg        [15:0]   int_reg_array_28_33_real;
  reg        [15:0]   int_reg_array_28_33_imag;
  reg        [15:0]   int_reg_array_28_34_real;
  reg        [15:0]   int_reg_array_28_34_imag;
  reg        [15:0]   int_reg_array_28_35_real;
  reg        [15:0]   int_reg_array_28_35_imag;
  reg        [15:0]   int_reg_array_28_36_real;
  reg        [15:0]   int_reg_array_28_36_imag;
  reg        [15:0]   int_reg_array_28_37_real;
  reg        [15:0]   int_reg_array_28_37_imag;
  reg        [15:0]   int_reg_array_28_38_real;
  reg        [15:0]   int_reg_array_28_38_imag;
  reg        [15:0]   int_reg_array_28_39_real;
  reg        [15:0]   int_reg_array_28_39_imag;
  reg        [15:0]   int_reg_array_28_40_real;
  reg        [15:0]   int_reg_array_28_40_imag;
  reg        [15:0]   int_reg_array_28_41_real;
  reg        [15:0]   int_reg_array_28_41_imag;
  reg        [15:0]   int_reg_array_28_42_real;
  reg        [15:0]   int_reg_array_28_42_imag;
  reg        [15:0]   int_reg_array_28_43_real;
  reg        [15:0]   int_reg_array_28_43_imag;
  reg        [15:0]   int_reg_array_28_44_real;
  reg        [15:0]   int_reg_array_28_44_imag;
  reg        [15:0]   int_reg_array_28_45_real;
  reg        [15:0]   int_reg_array_28_45_imag;
  reg        [15:0]   int_reg_array_28_46_real;
  reg        [15:0]   int_reg_array_28_46_imag;
  reg        [15:0]   int_reg_array_28_47_real;
  reg        [15:0]   int_reg_array_28_47_imag;
  reg        [15:0]   int_reg_array_28_48_real;
  reg        [15:0]   int_reg_array_28_48_imag;
  reg        [15:0]   int_reg_array_28_49_real;
  reg        [15:0]   int_reg_array_28_49_imag;
  reg        [15:0]   int_reg_array_30_0_real;
  reg        [15:0]   int_reg_array_30_0_imag;
  reg        [15:0]   int_reg_array_30_1_real;
  reg        [15:0]   int_reg_array_30_1_imag;
  reg        [15:0]   int_reg_array_30_2_real;
  reg        [15:0]   int_reg_array_30_2_imag;
  reg        [15:0]   int_reg_array_30_3_real;
  reg        [15:0]   int_reg_array_30_3_imag;
  reg        [15:0]   int_reg_array_30_4_real;
  reg        [15:0]   int_reg_array_30_4_imag;
  reg        [15:0]   int_reg_array_30_5_real;
  reg        [15:0]   int_reg_array_30_5_imag;
  reg        [15:0]   int_reg_array_30_6_real;
  reg        [15:0]   int_reg_array_30_6_imag;
  reg        [15:0]   int_reg_array_30_7_real;
  reg        [15:0]   int_reg_array_30_7_imag;
  reg        [15:0]   int_reg_array_30_8_real;
  reg        [15:0]   int_reg_array_30_8_imag;
  reg        [15:0]   int_reg_array_30_9_real;
  reg        [15:0]   int_reg_array_30_9_imag;
  reg        [15:0]   int_reg_array_30_10_real;
  reg        [15:0]   int_reg_array_30_10_imag;
  reg        [15:0]   int_reg_array_30_11_real;
  reg        [15:0]   int_reg_array_30_11_imag;
  reg        [15:0]   int_reg_array_30_12_real;
  reg        [15:0]   int_reg_array_30_12_imag;
  reg        [15:0]   int_reg_array_30_13_real;
  reg        [15:0]   int_reg_array_30_13_imag;
  reg        [15:0]   int_reg_array_30_14_real;
  reg        [15:0]   int_reg_array_30_14_imag;
  reg        [15:0]   int_reg_array_30_15_real;
  reg        [15:0]   int_reg_array_30_15_imag;
  reg        [15:0]   int_reg_array_30_16_real;
  reg        [15:0]   int_reg_array_30_16_imag;
  reg        [15:0]   int_reg_array_30_17_real;
  reg        [15:0]   int_reg_array_30_17_imag;
  reg        [15:0]   int_reg_array_30_18_real;
  reg        [15:0]   int_reg_array_30_18_imag;
  reg        [15:0]   int_reg_array_30_19_real;
  reg        [15:0]   int_reg_array_30_19_imag;
  reg        [15:0]   int_reg_array_30_20_real;
  reg        [15:0]   int_reg_array_30_20_imag;
  reg        [15:0]   int_reg_array_30_21_real;
  reg        [15:0]   int_reg_array_30_21_imag;
  reg        [15:0]   int_reg_array_30_22_real;
  reg        [15:0]   int_reg_array_30_22_imag;
  reg        [15:0]   int_reg_array_30_23_real;
  reg        [15:0]   int_reg_array_30_23_imag;
  reg        [15:0]   int_reg_array_30_24_real;
  reg        [15:0]   int_reg_array_30_24_imag;
  reg        [15:0]   int_reg_array_30_25_real;
  reg        [15:0]   int_reg_array_30_25_imag;
  reg        [15:0]   int_reg_array_30_26_real;
  reg        [15:0]   int_reg_array_30_26_imag;
  reg        [15:0]   int_reg_array_30_27_real;
  reg        [15:0]   int_reg_array_30_27_imag;
  reg        [15:0]   int_reg_array_30_28_real;
  reg        [15:0]   int_reg_array_30_28_imag;
  reg        [15:0]   int_reg_array_30_29_real;
  reg        [15:0]   int_reg_array_30_29_imag;
  reg        [15:0]   int_reg_array_30_30_real;
  reg        [15:0]   int_reg_array_30_30_imag;
  reg        [15:0]   int_reg_array_30_31_real;
  reg        [15:0]   int_reg_array_30_31_imag;
  reg        [15:0]   int_reg_array_30_32_real;
  reg        [15:0]   int_reg_array_30_32_imag;
  reg        [15:0]   int_reg_array_30_33_real;
  reg        [15:0]   int_reg_array_30_33_imag;
  reg        [15:0]   int_reg_array_30_34_real;
  reg        [15:0]   int_reg_array_30_34_imag;
  reg        [15:0]   int_reg_array_30_35_real;
  reg        [15:0]   int_reg_array_30_35_imag;
  reg        [15:0]   int_reg_array_30_36_real;
  reg        [15:0]   int_reg_array_30_36_imag;
  reg        [15:0]   int_reg_array_30_37_real;
  reg        [15:0]   int_reg_array_30_37_imag;
  reg        [15:0]   int_reg_array_30_38_real;
  reg        [15:0]   int_reg_array_30_38_imag;
  reg        [15:0]   int_reg_array_30_39_real;
  reg        [15:0]   int_reg_array_30_39_imag;
  reg        [15:0]   int_reg_array_30_40_real;
  reg        [15:0]   int_reg_array_30_40_imag;
  reg        [15:0]   int_reg_array_30_41_real;
  reg        [15:0]   int_reg_array_30_41_imag;
  reg        [15:0]   int_reg_array_30_42_real;
  reg        [15:0]   int_reg_array_30_42_imag;
  reg        [15:0]   int_reg_array_30_43_real;
  reg        [15:0]   int_reg_array_30_43_imag;
  reg        [15:0]   int_reg_array_30_44_real;
  reg        [15:0]   int_reg_array_30_44_imag;
  reg        [15:0]   int_reg_array_30_45_real;
  reg        [15:0]   int_reg_array_30_45_imag;
  reg        [15:0]   int_reg_array_30_46_real;
  reg        [15:0]   int_reg_array_30_46_imag;
  reg        [15:0]   int_reg_array_30_47_real;
  reg        [15:0]   int_reg_array_30_47_imag;
  reg        [15:0]   int_reg_array_30_48_real;
  reg        [15:0]   int_reg_array_30_48_imag;
  reg        [15:0]   int_reg_array_30_49_real;
  reg        [15:0]   int_reg_array_30_49_imag;
  reg        [15:0]   int_reg_array_29_0_real;
  reg        [15:0]   int_reg_array_29_0_imag;
  reg        [15:0]   int_reg_array_29_1_real;
  reg        [15:0]   int_reg_array_29_1_imag;
  reg        [15:0]   int_reg_array_29_2_real;
  reg        [15:0]   int_reg_array_29_2_imag;
  reg        [15:0]   int_reg_array_29_3_real;
  reg        [15:0]   int_reg_array_29_3_imag;
  reg        [15:0]   int_reg_array_29_4_real;
  reg        [15:0]   int_reg_array_29_4_imag;
  reg        [15:0]   int_reg_array_29_5_real;
  reg        [15:0]   int_reg_array_29_5_imag;
  reg        [15:0]   int_reg_array_29_6_real;
  reg        [15:0]   int_reg_array_29_6_imag;
  reg        [15:0]   int_reg_array_29_7_real;
  reg        [15:0]   int_reg_array_29_7_imag;
  reg        [15:0]   int_reg_array_29_8_real;
  reg        [15:0]   int_reg_array_29_8_imag;
  reg        [15:0]   int_reg_array_29_9_real;
  reg        [15:0]   int_reg_array_29_9_imag;
  reg        [15:0]   int_reg_array_29_10_real;
  reg        [15:0]   int_reg_array_29_10_imag;
  reg        [15:0]   int_reg_array_29_11_real;
  reg        [15:0]   int_reg_array_29_11_imag;
  reg        [15:0]   int_reg_array_29_12_real;
  reg        [15:0]   int_reg_array_29_12_imag;
  reg        [15:0]   int_reg_array_29_13_real;
  reg        [15:0]   int_reg_array_29_13_imag;
  reg        [15:0]   int_reg_array_29_14_real;
  reg        [15:0]   int_reg_array_29_14_imag;
  reg        [15:0]   int_reg_array_29_15_real;
  reg        [15:0]   int_reg_array_29_15_imag;
  reg        [15:0]   int_reg_array_29_16_real;
  reg        [15:0]   int_reg_array_29_16_imag;
  reg        [15:0]   int_reg_array_29_17_real;
  reg        [15:0]   int_reg_array_29_17_imag;
  reg        [15:0]   int_reg_array_29_18_real;
  reg        [15:0]   int_reg_array_29_18_imag;
  reg        [15:0]   int_reg_array_29_19_real;
  reg        [15:0]   int_reg_array_29_19_imag;
  reg        [15:0]   int_reg_array_29_20_real;
  reg        [15:0]   int_reg_array_29_20_imag;
  reg        [15:0]   int_reg_array_29_21_real;
  reg        [15:0]   int_reg_array_29_21_imag;
  reg        [15:0]   int_reg_array_29_22_real;
  reg        [15:0]   int_reg_array_29_22_imag;
  reg        [15:0]   int_reg_array_29_23_real;
  reg        [15:0]   int_reg_array_29_23_imag;
  reg        [15:0]   int_reg_array_29_24_real;
  reg        [15:0]   int_reg_array_29_24_imag;
  reg        [15:0]   int_reg_array_29_25_real;
  reg        [15:0]   int_reg_array_29_25_imag;
  reg        [15:0]   int_reg_array_29_26_real;
  reg        [15:0]   int_reg_array_29_26_imag;
  reg        [15:0]   int_reg_array_29_27_real;
  reg        [15:0]   int_reg_array_29_27_imag;
  reg        [15:0]   int_reg_array_29_28_real;
  reg        [15:0]   int_reg_array_29_28_imag;
  reg        [15:0]   int_reg_array_29_29_real;
  reg        [15:0]   int_reg_array_29_29_imag;
  reg        [15:0]   int_reg_array_29_30_real;
  reg        [15:0]   int_reg_array_29_30_imag;
  reg        [15:0]   int_reg_array_29_31_real;
  reg        [15:0]   int_reg_array_29_31_imag;
  reg        [15:0]   int_reg_array_29_32_real;
  reg        [15:0]   int_reg_array_29_32_imag;
  reg        [15:0]   int_reg_array_29_33_real;
  reg        [15:0]   int_reg_array_29_33_imag;
  reg        [15:0]   int_reg_array_29_34_real;
  reg        [15:0]   int_reg_array_29_34_imag;
  reg        [15:0]   int_reg_array_29_35_real;
  reg        [15:0]   int_reg_array_29_35_imag;
  reg        [15:0]   int_reg_array_29_36_real;
  reg        [15:0]   int_reg_array_29_36_imag;
  reg        [15:0]   int_reg_array_29_37_real;
  reg        [15:0]   int_reg_array_29_37_imag;
  reg        [15:0]   int_reg_array_29_38_real;
  reg        [15:0]   int_reg_array_29_38_imag;
  reg        [15:0]   int_reg_array_29_39_real;
  reg        [15:0]   int_reg_array_29_39_imag;
  reg        [15:0]   int_reg_array_29_40_real;
  reg        [15:0]   int_reg_array_29_40_imag;
  reg        [15:0]   int_reg_array_29_41_real;
  reg        [15:0]   int_reg_array_29_41_imag;
  reg        [15:0]   int_reg_array_29_42_real;
  reg        [15:0]   int_reg_array_29_42_imag;
  reg        [15:0]   int_reg_array_29_43_real;
  reg        [15:0]   int_reg_array_29_43_imag;
  reg        [15:0]   int_reg_array_29_44_real;
  reg        [15:0]   int_reg_array_29_44_imag;
  reg        [15:0]   int_reg_array_29_45_real;
  reg        [15:0]   int_reg_array_29_45_imag;
  reg        [15:0]   int_reg_array_29_46_real;
  reg        [15:0]   int_reg_array_29_46_imag;
  reg        [15:0]   int_reg_array_29_47_real;
  reg        [15:0]   int_reg_array_29_47_imag;
  reg        [15:0]   int_reg_array_29_48_real;
  reg        [15:0]   int_reg_array_29_48_imag;
  reg        [15:0]   int_reg_array_29_49_real;
  reg        [15:0]   int_reg_array_29_49_imag;
  reg        [15:0]   int_reg_array_8_0_real;
  reg        [15:0]   int_reg_array_8_0_imag;
  reg        [15:0]   int_reg_array_8_1_real;
  reg        [15:0]   int_reg_array_8_1_imag;
  reg        [15:0]   int_reg_array_8_2_real;
  reg        [15:0]   int_reg_array_8_2_imag;
  reg        [15:0]   int_reg_array_8_3_real;
  reg        [15:0]   int_reg_array_8_3_imag;
  reg        [15:0]   int_reg_array_8_4_real;
  reg        [15:0]   int_reg_array_8_4_imag;
  reg        [15:0]   int_reg_array_8_5_real;
  reg        [15:0]   int_reg_array_8_5_imag;
  reg        [15:0]   int_reg_array_8_6_real;
  reg        [15:0]   int_reg_array_8_6_imag;
  reg        [15:0]   int_reg_array_8_7_real;
  reg        [15:0]   int_reg_array_8_7_imag;
  reg        [15:0]   int_reg_array_8_8_real;
  reg        [15:0]   int_reg_array_8_8_imag;
  reg        [15:0]   int_reg_array_8_9_real;
  reg        [15:0]   int_reg_array_8_9_imag;
  reg        [15:0]   int_reg_array_8_10_real;
  reg        [15:0]   int_reg_array_8_10_imag;
  reg        [15:0]   int_reg_array_8_11_real;
  reg        [15:0]   int_reg_array_8_11_imag;
  reg        [15:0]   int_reg_array_8_12_real;
  reg        [15:0]   int_reg_array_8_12_imag;
  reg        [15:0]   int_reg_array_8_13_real;
  reg        [15:0]   int_reg_array_8_13_imag;
  reg        [15:0]   int_reg_array_8_14_real;
  reg        [15:0]   int_reg_array_8_14_imag;
  reg        [15:0]   int_reg_array_8_15_real;
  reg        [15:0]   int_reg_array_8_15_imag;
  reg        [15:0]   int_reg_array_8_16_real;
  reg        [15:0]   int_reg_array_8_16_imag;
  reg        [15:0]   int_reg_array_8_17_real;
  reg        [15:0]   int_reg_array_8_17_imag;
  reg        [15:0]   int_reg_array_8_18_real;
  reg        [15:0]   int_reg_array_8_18_imag;
  reg        [15:0]   int_reg_array_8_19_real;
  reg        [15:0]   int_reg_array_8_19_imag;
  reg        [15:0]   int_reg_array_8_20_real;
  reg        [15:0]   int_reg_array_8_20_imag;
  reg        [15:0]   int_reg_array_8_21_real;
  reg        [15:0]   int_reg_array_8_21_imag;
  reg        [15:0]   int_reg_array_8_22_real;
  reg        [15:0]   int_reg_array_8_22_imag;
  reg        [15:0]   int_reg_array_8_23_real;
  reg        [15:0]   int_reg_array_8_23_imag;
  reg        [15:0]   int_reg_array_8_24_real;
  reg        [15:0]   int_reg_array_8_24_imag;
  reg        [15:0]   int_reg_array_8_25_real;
  reg        [15:0]   int_reg_array_8_25_imag;
  reg        [15:0]   int_reg_array_8_26_real;
  reg        [15:0]   int_reg_array_8_26_imag;
  reg        [15:0]   int_reg_array_8_27_real;
  reg        [15:0]   int_reg_array_8_27_imag;
  reg        [15:0]   int_reg_array_8_28_real;
  reg        [15:0]   int_reg_array_8_28_imag;
  reg        [15:0]   int_reg_array_8_29_real;
  reg        [15:0]   int_reg_array_8_29_imag;
  reg        [15:0]   int_reg_array_8_30_real;
  reg        [15:0]   int_reg_array_8_30_imag;
  reg        [15:0]   int_reg_array_8_31_real;
  reg        [15:0]   int_reg_array_8_31_imag;
  reg        [15:0]   int_reg_array_8_32_real;
  reg        [15:0]   int_reg_array_8_32_imag;
  reg        [15:0]   int_reg_array_8_33_real;
  reg        [15:0]   int_reg_array_8_33_imag;
  reg        [15:0]   int_reg_array_8_34_real;
  reg        [15:0]   int_reg_array_8_34_imag;
  reg        [15:0]   int_reg_array_8_35_real;
  reg        [15:0]   int_reg_array_8_35_imag;
  reg        [15:0]   int_reg_array_8_36_real;
  reg        [15:0]   int_reg_array_8_36_imag;
  reg        [15:0]   int_reg_array_8_37_real;
  reg        [15:0]   int_reg_array_8_37_imag;
  reg        [15:0]   int_reg_array_8_38_real;
  reg        [15:0]   int_reg_array_8_38_imag;
  reg        [15:0]   int_reg_array_8_39_real;
  reg        [15:0]   int_reg_array_8_39_imag;
  reg        [15:0]   int_reg_array_8_40_real;
  reg        [15:0]   int_reg_array_8_40_imag;
  reg        [15:0]   int_reg_array_8_41_real;
  reg        [15:0]   int_reg_array_8_41_imag;
  reg        [15:0]   int_reg_array_8_42_real;
  reg        [15:0]   int_reg_array_8_42_imag;
  reg        [15:0]   int_reg_array_8_43_real;
  reg        [15:0]   int_reg_array_8_43_imag;
  reg        [15:0]   int_reg_array_8_44_real;
  reg        [15:0]   int_reg_array_8_44_imag;
  reg        [15:0]   int_reg_array_8_45_real;
  reg        [15:0]   int_reg_array_8_45_imag;
  reg        [15:0]   int_reg_array_8_46_real;
  reg        [15:0]   int_reg_array_8_46_imag;
  reg        [15:0]   int_reg_array_8_47_real;
  reg        [15:0]   int_reg_array_8_47_imag;
  reg        [15:0]   int_reg_array_8_48_real;
  reg        [15:0]   int_reg_array_8_48_imag;
  reg        [15:0]   int_reg_array_8_49_real;
  reg        [15:0]   int_reg_array_8_49_imag;
  reg        [15:0]   int_reg_array_7_0_real;
  reg        [15:0]   int_reg_array_7_0_imag;
  reg        [15:0]   int_reg_array_7_1_real;
  reg        [15:0]   int_reg_array_7_1_imag;
  reg        [15:0]   int_reg_array_7_2_real;
  reg        [15:0]   int_reg_array_7_2_imag;
  reg        [15:0]   int_reg_array_7_3_real;
  reg        [15:0]   int_reg_array_7_3_imag;
  reg        [15:0]   int_reg_array_7_4_real;
  reg        [15:0]   int_reg_array_7_4_imag;
  reg        [15:0]   int_reg_array_7_5_real;
  reg        [15:0]   int_reg_array_7_5_imag;
  reg        [15:0]   int_reg_array_7_6_real;
  reg        [15:0]   int_reg_array_7_6_imag;
  reg        [15:0]   int_reg_array_7_7_real;
  reg        [15:0]   int_reg_array_7_7_imag;
  reg        [15:0]   int_reg_array_7_8_real;
  reg        [15:0]   int_reg_array_7_8_imag;
  reg        [15:0]   int_reg_array_7_9_real;
  reg        [15:0]   int_reg_array_7_9_imag;
  reg        [15:0]   int_reg_array_7_10_real;
  reg        [15:0]   int_reg_array_7_10_imag;
  reg        [15:0]   int_reg_array_7_11_real;
  reg        [15:0]   int_reg_array_7_11_imag;
  reg        [15:0]   int_reg_array_7_12_real;
  reg        [15:0]   int_reg_array_7_12_imag;
  reg        [15:0]   int_reg_array_7_13_real;
  reg        [15:0]   int_reg_array_7_13_imag;
  reg        [15:0]   int_reg_array_7_14_real;
  reg        [15:0]   int_reg_array_7_14_imag;
  reg        [15:0]   int_reg_array_7_15_real;
  reg        [15:0]   int_reg_array_7_15_imag;
  reg        [15:0]   int_reg_array_7_16_real;
  reg        [15:0]   int_reg_array_7_16_imag;
  reg        [15:0]   int_reg_array_7_17_real;
  reg        [15:0]   int_reg_array_7_17_imag;
  reg        [15:0]   int_reg_array_7_18_real;
  reg        [15:0]   int_reg_array_7_18_imag;
  reg        [15:0]   int_reg_array_7_19_real;
  reg        [15:0]   int_reg_array_7_19_imag;
  reg        [15:0]   int_reg_array_7_20_real;
  reg        [15:0]   int_reg_array_7_20_imag;
  reg        [15:0]   int_reg_array_7_21_real;
  reg        [15:0]   int_reg_array_7_21_imag;
  reg        [15:0]   int_reg_array_7_22_real;
  reg        [15:0]   int_reg_array_7_22_imag;
  reg        [15:0]   int_reg_array_7_23_real;
  reg        [15:0]   int_reg_array_7_23_imag;
  reg        [15:0]   int_reg_array_7_24_real;
  reg        [15:0]   int_reg_array_7_24_imag;
  reg        [15:0]   int_reg_array_7_25_real;
  reg        [15:0]   int_reg_array_7_25_imag;
  reg        [15:0]   int_reg_array_7_26_real;
  reg        [15:0]   int_reg_array_7_26_imag;
  reg        [15:0]   int_reg_array_7_27_real;
  reg        [15:0]   int_reg_array_7_27_imag;
  reg        [15:0]   int_reg_array_7_28_real;
  reg        [15:0]   int_reg_array_7_28_imag;
  reg        [15:0]   int_reg_array_7_29_real;
  reg        [15:0]   int_reg_array_7_29_imag;
  reg        [15:0]   int_reg_array_7_30_real;
  reg        [15:0]   int_reg_array_7_30_imag;
  reg        [15:0]   int_reg_array_7_31_real;
  reg        [15:0]   int_reg_array_7_31_imag;
  reg        [15:0]   int_reg_array_7_32_real;
  reg        [15:0]   int_reg_array_7_32_imag;
  reg        [15:0]   int_reg_array_7_33_real;
  reg        [15:0]   int_reg_array_7_33_imag;
  reg        [15:0]   int_reg_array_7_34_real;
  reg        [15:0]   int_reg_array_7_34_imag;
  reg        [15:0]   int_reg_array_7_35_real;
  reg        [15:0]   int_reg_array_7_35_imag;
  reg        [15:0]   int_reg_array_7_36_real;
  reg        [15:0]   int_reg_array_7_36_imag;
  reg        [15:0]   int_reg_array_7_37_real;
  reg        [15:0]   int_reg_array_7_37_imag;
  reg        [15:0]   int_reg_array_7_38_real;
  reg        [15:0]   int_reg_array_7_38_imag;
  reg        [15:0]   int_reg_array_7_39_real;
  reg        [15:0]   int_reg_array_7_39_imag;
  reg        [15:0]   int_reg_array_7_40_real;
  reg        [15:0]   int_reg_array_7_40_imag;
  reg        [15:0]   int_reg_array_7_41_real;
  reg        [15:0]   int_reg_array_7_41_imag;
  reg        [15:0]   int_reg_array_7_42_real;
  reg        [15:0]   int_reg_array_7_42_imag;
  reg        [15:0]   int_reg_array_7_43_real;
  reg        [15:0]   int_reg_array_7_43_imag;
  reg        [15:0]   int_reg_array_7_44_real;
  reg        [15:0]   int_reg_array_7_44_imag;
  reg        [15:0]   int_reg_array_7_45_real;
  reg        [15:0]   int_reg_array_7_45_imag;
  reg        [15:0]   int_reg_array_7_46_real;
  reg        [15:0]   int_reg_array_7_46_imag;
  reg        [15:0]   int_reg_array_7_47_real;
  reg        [15:0]   int_reg_array_7_47_imag;
  reg        [15:0]   int_reg_array_7_48_real;
  reg        [15:0]   int_reg_array_7_48_imag;
  reg        [15:0]   int_reg_array_7_49_real;
  reg        [15:0]   int_reg_array_7_49_imag;
  reg        [15:0]   int_reg_array_20_0_real;
  reg        [15:0]   int_reg_array_20_0_imag;
  reg        [15:0]   int_reg_array_20_1_real;
  reg        [15:0]   int_reg_array_20_1_imag;
  reg        [15:0]   int_reg_array_20_2_real;
  reg        [15:0]   int_reg_array_20_2_imag;
  reg        [15:0]   int_reg_array_20_3_real;
  reg        [15:0]   int_reg_array_20_3_imag;
  reg        [15:0]   int_reg_array_20_4_real;
  reg        [15:0]   int_reg_array_20_4_imag;
  reg        [15:0]   int_reg_array_20_5_real;
  reg        [15:0]   int_reg_array_20_5_imag;
  reg        [15:0]   int_reg_array_20_6_real;
  reg        [15:0]   int_reg_array_20_6_imag;
  reg        [15:0]   int_reg_array_20_7_real;
  reg        [15:0]   int_reg_array_20_7_imag;
  reg        [15:0]   int_reg_array_20_8_real;
  reg        [15:0]   int_reg_array_20_8_imag;
  reg        [15:0]   int_reg_array_20_9_real;
  reg        [15:0]   int_reg_array_20_9_imag;
  reg        [15:0]   int_reg_array_20_10_real;
  reg        [15:0]   int_reg_array_20_10_imag;
  reg        [15:0]   int_reg_array_20_11_real;
  reg        [15:0]   int_reg_array_20_11_imag;
  reg        [15:0]   int_reg_array_20_12_real;
  reg        [15:0]   int_reg_array_20_12_imag;
  reg        [15:0]   int_reg_array_20_13_real;
  reg        [15:0]   int_reg_array_20_13_imag;
  reg        [15:0]   int_reg_array_20_14_real;
  reg        [15:0]   int_reg_array_20_14_imag;
  reg        [15:0]   int_reg_array_20_15_real;
  reg        [15:0]   int_reg_array_20_15_imag;
  reg        [15:0]   int_reg_array_20_16_real;
  reg        [15:0]   int_reg_array_20_16_imag;
  reg        [15:0]   int_reg_array_20_17_real;
  reg        [15:0]   int_reg_array_20_17_imag;
  reg        [15:0]   int_reg_array_20_18_real;
  reg        [15:0]   int_reg_array_20_18_imag;
  reg        [15:0]   int_reg_array_20_19_real;
  reg        [15:0]   int_reg_array_20_19_imag;
  reg        [15:0]   int_reg_array_20_20_real;
  reg        [15:0]   int_reg_array_20_20_imag;
  reg        [15:0]   int_reg_array_20_21_real;
  reg        [15:0]   int_reg_array_20_21_imag;
  reg        [15:0]   int_reg_array_20_22_real;
  reg        [15:0]   int_reg_array_20_22_imag;
  reg        [15:0]   int_reg_array_20_23_real;
  reg        [15:0]   int_reg_array_20_23_imag;
  reg        [15:0]   int_reg_array_20_24_real;
  reg        [15:0]   int_reg_array_20_24_imag;
  reg        [15:0]   int_reg_array_20_25_real;
  reg        [15:0]   int_reg_array_20_25_imag;
  reg        [15:0]   int_reg_array_20_26_real;
  reg        [15:0]   int_reg_array_20_26_imag;
  reg        [15:0]   int_reg_array_20_27_real;
  reg        [15:0]   int_reg_array_20_27_imag;
  reg        [15:0]   int_reg_array_20_28_real;
  reg        [15:0]   int_reg_array_20_28_imag;
  reg        [15:0]   int_reg_array_20_29_real;
  reg        [15:0]   int_reg_array_20_29_imag;
  reg        [15:0]   int_reg_array_20_30_real;
  reg        [15:0]   int_reg_array_20_30_imag;
  reg        [15:0]   int_reg_array_20_31_real;
  reg        [15:0]   int_reg_array_20_31_imag;
  reg        [15:0]   int_reg_array_20_32_real;
  reg        [15:0]   int_reg_array_20_32_imag;
  reg        [15:0]   int_reg_array_20_33_real;
  reg        [15:0]   int_reg_array_20_33_imag;
  reg        [15:0]   int_reg_array_20_34_real;
  reg        [15:0]   int_reg_array_20_34_imag;
  reg        [15:0]   int_reg_array_20_35_real;
  reg        [15:0]   int_reg_array_20_35_imag;
  reg        [15:0]   int_reg_array_20_36_real;
  reg        [15:0]   int_reg_array_20_36_imag;
  reg        [15:0]   int_reg_array_20_37_real;
  reg        [15:0]   int_reg_array_20_37_imag;
  reg        [15:0]   int_reg_array_20_38_real;
  reg        [15:0]   int_reg_array_20_38_imag;
  reg        [15:0]   int_reg_array_20_39_real;
  reg        [15:0]   int_reg_array_20_39_imag;
  reg        [15:0]   int_reg_array_20_40_real;
  reg        [15:0]   int_reg_array_20_40_imag;
  reg        [15:0]   int_reg_array_20_41_real;
  reg        [15:0]   int_reg_array_20_41_imag;
  reg        [15:0]   int_reg_array_20_42_real;
  reg        [15:0]   int_reg_array_20_42_imag;
  reg        [15:0]   int_reg_array_20_43_real;
  reg        [15:0]   int_reg_array_20_43_imag;
  reg        [15:0]   int_reg_array_20_44_real;
  reg        [15:0]   int_reg_array_20_44_imag;
  reg        [15:0]   int_reg_array_20_45_real;
  reg        [15:0]   int_reg_array_20_45_imag;
  reg        [15:0]   int_reg_array_20_46_real;
  reg        [15:0]   int_reg_array_20_46_imag;
  reg        [15:0]   int_reg_array_20_47_real;
  reg        [15:0]   int_reg_array_20_47_imag;
  reg        [15:0]   int_reg_array_20_48_real;
  reg        [15:0]   int_reg_array_20_48_imag;
  reg        [15:0]   int_reg_array_20_49_real;
  reg        [15:0]   int_reg_array_20_49_imag;
  reg        [15:0]   int_reg_array_1_0_real;
  reg        [15:0]   int_reg_array_1_0_imag;
  reg        [15:0]   int_reg_array_1_1_real;
  reg        [15:0]   int_reg_array_1_1_imag;
  reg        [15:0]   int_reg_array_1_2_real;
  reg        [15:0]   int_reg_array_1_2_imag;
  reg        [15:0]   int_reg_array_1_3_real;
  reg        [15:0]   int_reg_array_1_3_imag;
  reg        [15:0]   int_reg_array_1_4_real;
  reg        [15:0]   int_reg_array_1_4_imag;
  reg        [15:0]   int_reg_array_1_5_real;
  reg        [15:0]   int_reg_array_1_5_imag;
  reg        [15:0]   int_reg_array_1_6_real;
  reg        [15:0]   int_reg_array_1_6_imag;
  reg        [15:0]   int_reg_array_1_7_real;
  reg        [15:0]   int_reg_array_1_7_imag;
  reg        [15:0]   int_reg_array_1_8_real;
  reg        [15:0]   int_reg_array_1_8_imag;
  reg        [15:0]   int_reg_array_1_9_real;
  reg        [15:0]   int_reg_array_1_9_imag;
  reg        [15:0]   int_reg_array_1_10_real;
  reg        [15:0]   int_reg_array_1_10_imag;
  reg        [15:0]   int_reg_array_1_11_real;
  reg        [15:0]   int_reg_array_1_11_imag;
  reg        [15:0]   int_reg_array_1_12_real;
  reg        [15:0]   int_reg_array_1_12_imag;
  reg        [15:0]   int_reg_array_1_13_real;
  reg        [15:0]   int_reg_array_1_13_imag;
  reg        [15:0]   int_reg_array_1_14_real;
  reg        [15:0]   int_reg_array_1_14_imag;
  reg        [15:0]   int_reg_array_1_15_real;
  reg        [15:0]   int_reg_array_1_15_imag;
  reg        [15:0]   int_reg_array_1_16_real;
  reg        [15:0]   int_reg_array_1_16_imag;
  reg        [15:0]   int_reg_array_1_17_real;
  reg        [15:0]   int_reg_array_1_17_imag;
  reg        [15:0]   int_reg_array_1_18_real;
  reg        [15:0]   int_reg_array_1_18_imag;
  reg        [15:0]   int_reg_array_1_19_real;
  reg        [15:0]   int_reg_array_1_19_imag;
  reg        [15:0]   int_reg_array_1_20_real;
  reg        [15:0]   int_reg_array_1_20_imag;
  reg        [15:0]   int_reg_array_1_21_real;
  reg        [15:0]   int_reg_array_1_21_imag;
  reg        [15:0]   int_reg_array_1_22_real;
  reg        [15:0]   int_reg_array_1_22_imag;
  reg        [15:0]   int_reg_array_1_23_real;
  reg        [15:0]   int_reg_array_1_23_imag;
  reg        [15:0]   int_reg_array_1_24_real;
  reg        [15:0]   int_reg_array_1_24_imag;
  reg        [15:0]   int_reg_array_1_25_real;
  reg        [15:0]   int_reg_array_1_25_imag;
  reg        [15:0]   int_reg_array_1_26_real;
  reg        [15:0]   int_reg_array_1_26_imag;
  reg        [15:0]   int_reg_array_1_27_real;
  reg        [15:0]   int_reg_array_1_27_imag;
  reg        [15:0]   int_reg_array_1_28_real;
  reg        [15:0]   int_reg_array_1_28_imag;
  reg        [15:0]   int_reg_array_1_29_real;
  reg        [15:0]   int_reg_array_1_29_imag;
  reg        [15:0]   int_reg_array_1_30_real;
  reg        [15:0]   int_reg_array_1_30_imag;
  reg        [15:0]   int_reg_array_1_31_real;
  reg        [15:0]   int_reg_array_1_31_imag;
  reg        [15:0]   int_reg_array_1_32_real;
  reg        [15:0]   int_reg_array_1_32_imag;
  reg        [15:0]   int_reg_array_1_33_real;
  reg        [15:0]   int_reg_array_1_33_imag;
  reg        [15:0]   int_reg_array_1_34_real;
  reg        [15:0]   int_reg_array_1_34_imag;
  reg        [15:0]   int_reg_array_1_35_real;
  reg        [15:0]   int_reg_array_1_35_imag;
  reg        [15:0]   int_reg_array_1_36_real;
  reg        [15:0]   int_reg_array_1_36_imag;
  reg        [15:0]   int_reg_array_1_37_real;
  reg        [15:0]   int_reg_array_1_37_imag;
  reg        [15:0]   int_reg_array_1_38_real;
  reg        [15:0]   int_reg_array_1_38_imag;
  reg        [15:0]   int_reg_array_1_39_real;
  reg        [15:0]   int_reg_array_1_39_imag;
  reg        [15:0]   int_reg_array_1_40_real;
  reg        [15:0]   int_reg_array_1_40_imag;
  reg        [15:0]   int_reg_array_1_41_real;
  reg        [15:0]   int_reg_array_1_41_imag;
  reg        [15:0]   int_reg_array_1_42_real;
  reg        [15:0]   int_reg_array_1_42_imag;
  reg        [15:0]   int_reg_array_1_43_real;
  reg        [15:0]   int_reg_array_1_43_imag;
  reg        [15:0]   int_reg_array_1_44_real;
  reg        [15:0]   int_reg_array_1_44_imag;
  reg        [15:0]   int_reg_array_1_45_real;
  reg        [15:0]   int_reg_array_1_45_imag;
  reg        [15:0]   int_reg_array_1_46_real;
  reg        [15:0]   int_reg_array_1_46_imag;
  reg        [15:0]   int_reg_array_1_47_real;
  reg        [15:0]   int_reg_array_1_47_imag;
  reg        [15:0]   int_reg_array_1_48_real;
  reg        [15:0]   int_reg_array_1_48_imag;
  reg        [15:0]   int_reg_array_1_49_real;
  reg        [15:0]   int_reg_array_1_49_imag;
  reg        [15:0]   int_reg_array_2_0_real;
  reg        [15:0]   int_reg_array_2_0_imag;
  reg        [15:0]   int_reg_array_2_1_real;
  reg        [15:0]   int_reg_array_2_1_imag;
  reg        [15:0]   int_reg_array_2_2_real;
  reg        [15:0]   int_reg_array_2_2_imag;
  reg        [15:0]   int_reg_array_2_3_real;
  reg        [15:0]   int_reg_array_2_3_imag;
  reg        [15:0]   int_reg_array_2_4_real;
  reg        [15:0]   int_reg_array_2_4_imag;
  reg        [15:0]   int_reg_array_2_5_real;
  reg        [15:0]   int_reg_array_2_5_imag;
  reg        [15:0]   int_reg_array_2_6_real;
  reg        [15:0]   int_reg_array_2_6_imag;
  reg        [15:0]   int_reg_array_2_7_real;
  reg        [15:0]   int_reg_array_2_7_imag;
  reg        [15:0]   int_reg_array_2_8_real;
  reg        [15:0]   int_reg_array_2_8_imag;
  reg        [15:0]   int_reg_array_2_9_real;
  reg        [15:0]   int_reg_array_2_9_imag;
  reg        [15:0]   int_reg_array_2_10_real;
  reg        [15:0]   int_reg_array_2_10_imag;
  reg        [15:0]   int_reg_array_2_11_real;
  reg        [15:0]   int_reg_array_2_11_imag;
  reg        [15:0]   int_reg_array_2_12_real;
  reg        [15:0]   int_reg_array_2_12_imag;
  reg        [15:0]   int_reg_array_2_13_real;
  reg        [15:0]   int_reg_array_2_13_imag;
  reg        [15:0]   int_reg_array_2_14_real;
  reg        [15:0]   int_reg_array_2_14_imag;
  reg        [15:0]   int_reg_array_2_15_real;
  reg        [15:0]   int_reg_array_2_15_imag;
  reg        [15:0]   int_reg_array_2_16_real;
  reg        [15:0]   int_reg_array_2_16_imag;
  reg        [15:0]   int_reg_array_2_17_real;
  reg        [15:0]   int_reg_array_2_17_imag;
  reg        [15:0]   int_reg_array_2_18_real;
  reg        [15:0]   int_reg_array_2_18_imag;
  reg        [15:0]   int_reg_array_2_19_real;
  reg        [15:0]   int_reg_array_2_19_imag;
  reg        [15:0]   int_reg_array_2_20_real;
  reg        [15:0]   int_reg_array_2_20_imag;
  reg        [15:0]   int_reg_array_2_21_real;
  reg        [15:0]   int_reg_array_2_21_imag;
  reg        [15:0]   int_reg_array_2_22_real;
  reg        [15:0]   int_reg_array_2_22_imag;
  reg        [15:0]   int_reg_array_2_23_real;
  reg        [15:0]   int_reg_array_2_23_imag;
  reg        [15:0]   int_reg_array_2_24_real;
  reg        [15:0]   int_reg_array_2_24_imag;
  reg        [15:0]   int_reg_array_2_25_real;
  reg        [15:0]   int_reg_array_2_25_imag;
  reg        [15:0]   int_reg_array_2_26_real;
  reg        [15:0]   int_reg_array_2_26_imag;
  reg        [15:0]   int_reg_array_2_27_real;
  reg        [15:0]   int_reg_array_2_27_imag;
  reg        [15:0]   int_reg_array_2_28_real;
  reg        [15:0]   int_reg_array_2_28_imag;
  reg        [15:0]   int_reg_array_2_29_real;
  reg        [15:0]   int_reg_array_2_29_imag;
  reg        [15:0]   int_reg_array_2_30_real;
  reg        [15:0]   int_reg_array_2_30_imag;
  reg        [15:0]   int_reg_array_2_31_real;
  reg        [15:0]   int_reg_array_2_31_imag;
  reg        [15:0]   int_reg_array_2_32_real;
  reg        [15:0]   int_reg_array_2_32_imag;
  reg        [15:0]   int_reg_array_2_33_real;
  reg        [15:0]   int_reg_array_2_33_imag;
  reg        [15:0]   int_reg_array_2_34_real;
  reg        [15:0]   int_reg_array_2_34_imag;
  reg        [15:0]   int_reg_array_2_35_real;
  reg        [15:0]   int_reg_array_2_35_imag;
  reg        [15:0]   int_reg_array_2_36_real;
  reg        [15:0]   int_reg_array_2_36_imag;
  reg        [15:0]   int_reg_array_2_37_real;
  reg        [15:0]   int_reg_array_2_37_imag;
  reg        [15:0]   int_reg_array_2_38_real;
  reg        [15:0]   int_reg_array_2_38_imag;
  reg        [15:0]   int_reg_array_2_39_real;
  reg        [15:0]   int_reg_array_2_39_imag;
  reg        [15:0]   int_reg_array_2_40_real;
  reg        [15:0]   int_reg_array_2_40_imag;
  reg        [15:0]   int_reg_array_2_41_real;
  reg        [15:0]   int_reg_array_2_41_imag;
  reg        [15:0]   int_reg_array_2_42_real;
  reg        [15:0]   int_reg_array_2_42_imag;
  reg        [15:0]   int_reg_array_2_43_real;
  reg        [15:0]   int_reg_array_2_43_imag;
  reg        [15:0]   int_reg_array_2_44_real;
  reg        [15:0]   int_reg_array_2_44_imag;
  reg        [15:0]   int_reg_array_2_45_real;
  reg        [15:0]   int_reg_array_2_45_imag;
  reg        [15:0]   int_reg_array_2_46_real;
  reg        [15:0]   int_reg_array_2_46_imag;
  reg        [15:0]   int_reg_array_2_47_real;
  reg        [15:0]   int_reg_array_2_47_imag;
  reg        [15:0]   int_reg_array_2_48_real;
  reg        [15:0]   int_reg_array_2_48_imag;
  reg        [15:0]   int_reg_array_2_49_real;
  reg        [15:0]   int_reg_array_2_49_imag;
  reg        [15:0]   int_reg_array_38_0_real;
  reg        [15:0]   int_reg_array_38_0_imag;
  reg        [15:0]   int_reg_array_38_1_real;
  reg        [15:0]   int_reg_array_38_1_imag;
  reg        [15:0]   int_reg_array_38_2_real;
  reg        [15:0]   int_reg_array_38_2_imag;
  reg        [15:0]   int_reg_array_38_3_real;
  reg        [15:0]   int_reg_array_38_3_imag;
  reg        [15:0]   int_reg_array_38_4_real;
  reg        [15:0]   int_reg_array_38_4_imag;
  reg        [15:0]   int_reg_array_38_5_real;
  reg        [15:0]   int_reg_array_38_5_imag;
  reg        [15:0]   int_reg_array_38_6_real;
  reg        [15:0]   int_reg_array_38_6_imag;
  reg        [15:0]   int_reg_array_38_7_real;
  reg        [15:0]   int_reg_array_38_7_imag;
  reg        [15:0]   int_reg_array_38_8_real;
  reg        [15:0]   int_reg_array_38_8_imag;
  reg        [15:0]   int_reg_array_38_9_real;
  reg        [15:0]   int_reg_array_38_9_imag;
  reg        [15:0]   int_reg_array_38_10_real;
  reg        [15:0]   int_reg_array_38_10_imag;
  reg        [15:0]   int_reg_array_38_11_real;
  reg        [15:0]   int_reg_array_38_11_imag;
  reg        [15:0]   int_reg_array_38_12_real;
  reg        [15:0]   int_reg_array_38_12_imag;
  reg        [15:0]   int_reg_array_38_13_real;
  reg        [15:0]   int_reg_array_38_13_imag;
  reg        [15:0]   int_reg_array_38_14_real;
  reg        [15:0]   int_reg_array_38_14_imag;
  reg        [15:0]   int_reg_array_38_15_real;
  reg        [15:0]   int_reg_array_38_15_imag;
  reg        [15:0]   int_reg_array_38_16_real;
  reg        [15:0]   int_reg_array_38_16_imag;
  reg        [15:0]   int_reg_array_38_17_real;
  reg        [15:0]   int_reg_array_38_17_imag;
  reg        [15:0]   int_reg_array_38_18_real;
  reg        [15:0]   int_reg_array_38_18_imag;
  reg        [15:0]   int_reg_array_38_19_real;
  reg        [15:0]   int_reg_array_38_19_imag;
  reg        [15:0]   int_reg_array_38_20_real;
  reg        [15:0]   int_reg_array_38_20_imag;
  reg        [15:0]   int_reg_array_38_21_real;
  reg        [15:0]   int_reg_array_38_21_imag;
  reg        [15:0]   int_reg_array_38_22_real;
  reg        [15:0]   int_reg_array_38_22_imag;
  reg        [15:0]   int_reg_array_38_23_real;
  reg        [15:0]   int_reg_array_38_23_imag;
  reg        [15:0]   int_reg_array_38_24_real;
  reg        [15:0]   int_reg_array_38_24_imag;
  reg        [15:0]   int_reg_array_38_25_real;
  reg        [15:0]   int_reg_array_38_25_imag;
  reg        [15:0]   int_reg_array_38_26_real;
  reg        [15:0]   int_reg_array_38_26_imag;
  reg        [15:0]   int_reg_array_38_27_real;
  reg        [15:0]   int_reg_array_38_27_imag;
  reg        [15:0]   int_reg_array_38_28_real;
  reg        [15:0]   int_reg_array_38_28_imag;
  reg        [15:0]   int_reg_array_38_29_real;
  reg        [15:0]   int_reg_array_38_29_imag;
  reg        [15:0]   int_reg_array_38_30_real;
  reg        [15:0]   int_reg_array_38_30_imag;
  reg        [15:0]   int_reg_array_38_31_real;
  reg        [15:0]   int_reg_array_38_31_imag;
  reg        [15:0]   int_reg_array_38_32_real;
  reg        [15:0]   int_reg_array_38_32_imag;
  reg        [15:0]   int_reg_array_38_33_real;
  reg        [15:0]   int_reg_array_38_33_imag;
  reg        [15:0]   int_reg_array_38_34_real;
  reg        [15:0]   int_reg_array_38_34_imag;
  reg        [15:0]   int_reg_array_38_35_real;
  reg        [15:0]   int_reg_array_38_35_imag;
  reg        [15:0]   int_reg_array_38_36_real;
  reg        [15:0]   int_reg_array_38_36_imag;
  reg        [15:0]   int_reg_array_38_37_real;
  reg        [15:0]   int_reg_array_38_37_imag;
  reg        [15:0]   int_reg_array_38_38_real;
  reg        [15:0]   int_reg_array_38_38_imag;
  reg        [15:0]   int_reg_array_38_39_real;
  reg        [15:0]   int_reg_array_38_39_imag;
  reg        [15:0]   int_reg_array_38_40_real;
  reg        [15:0]   int_reg_array_38_40_imag;
  reg        [15:0]   int_reg_array_38_41_real;
  reg        [15:0]   int_reg_array_38_41_imag;
  reg        [15:0]   int_reg_array_38_42_real;
  reg        [15:0]   int_reg_array_38_42_imag;
  reg        [15:0]   int_reg_array_38_43_real;
  reg        [15:0]   int_reg_array_38_43_imag;
  reg        [15:0]   int_reg_array_38_44_real;
  reg        [15:0]   int_reg_array_38_44_imag;
  reg        [15:0]   int_reg_array_38_45_real;
  reg        [15:0]   int_reg_array_38_45_imag;
  reg        [15:0]   int_reg_array_38_46_real;
  reg        [15:0]   int_reg_array_38_46_imag;
  reg        [15:0]   int_reg_array_38_47_real;
  reg        [15:0]   int_reg_array_38_47_imag;
  reg        [15:0]   int_reg_array_38_48_real;
  reg        [15:0]   int_reg_array_38_48_imag;
  reg        [15:0]   int_reg_array_38_49_real;
  reg        [15:0]   int_reg_array_38_49_imag;
  reg        [15:0]   int_reg_array_6_0_real;
  reg        [15:0]   int_reg_array_6_0_imag;
  reg        [15:0]   int_reg_array_6_1_real;
  reg        [15:0]   int_reg_array_6_1_imag;
  reg        [15:0]   int_reg_array_6_2_real;
  reg        [15:0]   int_reg_array_6_2_imag;
  reg        [15:0]   int_reg_array_6_3_real;
  reg        [15:0]   int_reg_array_6_3_imag;
  reg        [15:0]   int_reg_array_6_4_real;
  reg        [15:0]   int_reg_array_6_4_imag;
  reg        [15:0]   int_reg_array_6_5_real;
  reg        [15:0]   int_reg_array_6_5_imag;
  reg        [15:0]   int_reg_array_6_6_real;
  reg        [15:0]   int_reg_array_6_6_imag;
  reg        [15:0]   int_reg_array_6_7_real;
  reg        [15:0]   int_reg_array_6_7_imag;
  reg        [15:0]   int_reg_array_6_8_real;
  reg        [15:0]   int_reg_array_6_8_imag;
  reg        [15:0]   int_reg_array_6_9_real;
  reg        [15:0]   int_reg_array_6_9_imag;
  reg        [15:0]   int_reg_array_6_10_real;
  reg        [15:0]   int_reg_array_6_10_imag;
  reg        [15:0]   int_reg_array_6_11_real;
  reg        [15:0]   int_reg_array_6_11_imag;
  reg        [15:0]   int_reg_array_6_12_real;
  reg        [15:0]   int_reg_array_6_12_imag;
  reg        [15:0]   int_reg_array_6_13_real;
  reg        [15:0]   int_reg_array_6_13_imag;
  reg        [15:0]   int_reg_array_6_14_real;
  reg        [15:0]   int_reg_array_6_14_imag;
  reg        [15:0]   int_reg_array_6_15_real;
  reg        [15:0]   int_reg_array_6_15_imag;
  reg        [15:0]   int_reg_array_6_16_real;
  reg        [15:0]   int_reg_array_6_16_imag;
  reg        [15:0]   int_reg_array_6_17_real;
  reg        [15:0]   int_reg_array_6_17_imag;
  reg        [15:0]   int_reg_array_6_18_real;
  reg        [15:0]   int_reg_array_6_18_imag;
  reg        [15:0]   int_reg_array_6_19_real;
  reg        [15:0]   int_reg_array_6_19_imag;
  reg        [15:0]   int_reg_array_6_20_real;
  reg        [15:0]   int_reg_array_6_20_imag;
  reg        [15:0]   int_reg_array_6_21_real;
  reg        [15:0]   int_reg_array_6_21_imag;
  reg        [15:0]   int_reg_array_6_22_real;
  reg        [15:0]   int_reg_array_6_22_imag;
  reg        [15:0]   int_reg_array_6_23_real;
  reg        [15:0]   int_reg_array_6_23_imag;
  reg        [15:0]   int_reg_array_6_24_real;
  reg        [15:0]   int_reg_array_6_24_imag;
  reg        [15:0]   int_reg_array_6_25_real;
  reg        [15:0]   int_reg_array_6_25_imag;
  reg        [15:0]   int_reg_array_6_26_real;
  reg        [15:0]   int_reg_array_6_26_imag;
  reg        [15:0]   int_reg_array_6_27_real;
  reg        [15:0]   int_reg_array_6_27_imag;
  reg        [15:0]   int_reg_array_6_28_real;
  reg        [15:0]   int_reg_array_6_28_imag;
  reg        [15:0]   int_reg_array_6_29_real;
  reg        [15:0]   int_reg_array_6_29_imag;
  reg        [15:0]   int_reg_array_6_30_real;
  reg        [15:0]   int_reg_array_6_30_imag;
  reg        [15:0]   int_reg_array_6_31_real;
  reg        [15:0]   int_reg_array_6_31_imag;
  reg        [15:0]   int_reg_array_6_32_real;
  reg        [15:0]   int_reg_array_6_32_imag;
  reg        [15:0]   int_reg_array_6_33_real;
  reg        [15:0]   int_reg_array_6_33_imag;
  reg        [15:0]   int_reg_array_6_34_real;
  reg        [15:0]   int_reg_array_6_34_imag;
  reg        [15:0]   int_reg_array_6_35_real;
  reg        [15:0]   int_reg_array_6_35_imag;
  reg        [15:0]   int_reg_array_6_36_real;
  reg        [15:0]   int_reg_array_6_36_imag;
  reg        [15:0]   int_reg_array_6_37_real;
  reg        [15:0]   int_reg_array_6_37_imag;
  reg        [15:0]   int_reg_array_6_38_real;
  reg        [15:0]   int_reg_array_6_38_imag;
  reg        [15:0]   int_reg_array_6_39_real;
  reg        [15:0]   int_reg_array_6_39_imag;
  reg        [15:0]   int_reg_array_6_40_real;
  reg        [15:0]   int_reg_array_6_40_imag;
  reg        [15:0]   int_reg_array_6_41_real;
  reg        [15:0]   int_reg_array_6_41_imag;
  reg        [15:0]   int_reg_array_6_42_real;
  reg        [15:0]   int_reg_array_6_42_imag;
  reg        [15:0]   int_reg_array_6_43_real;
  reg        [15:0]   int_reg_array_6_43_imag;
  reg        [15:0]   int_reg_array_6_44_real;
  reg        [15:0]   int_reg_array_6_44_imag;
  reg        [15:0]   int_reg_array_6_45_real;
  reg        [15:0]   int_reg_array_6_45_imag;
  reg        [15:0]   int_reg_array_6_46_real;
  reg        [15:0]   int_reg_array_6_46_imag;
  reg        [15:0]   int_reg_array_6_47_real;
  reg        [15:0]   int_reg_array_6_47_imag;
  reg        [15:0]   int_reg_array_6_48_real;
  reg        [15:0]   int_reg_array_6_48_imag;
  reg        [15:0]   int_reg_array_6_49_real;
  reg        [15:0]   int_reg_array_6_49_imag;
  reg        [15:0]   int_reg_array_5_0_real;
  reg        [15:0]   int_reg_array_5_0_imag;
  reg        [15:0]   int_reg_array_5_1_real;
  reg        [15:0]   int_reg_array_5_1_imag;
  reg        [15:0]   int_reg_array_5_2_real;
  reg        [15:0]   int_reg_array_5_2_imag;
  reg        [15:0]   int_reg_array_5_3_real;
  reg        [15:0]   int_reg_array_5_3_imag;
  reg        [15:0]   int_reg_array_5_4_real;
  reg        [15:0]   int_reg_array_5_4_imag;
  reg        [15:0]   int_reg_array_5_5_real;
  reg        [15:0]   int_reg_array_5_5_imag;
  reg        [15:0]   int_reg_array_5_6_real;
  reg        [15:0]   int_reg_array_5_6_imag;
  reg        [15:0]   int_reg_array_5_7_real;
  reg        [15:0]   int_reg_array_5_7_imag;
  reg        [15:0]   int_reg_array_5_8_real;
  reg        [15:0]   int_reg_array_5_8_imag;
  reg        [15:0]   int_reg_array_5_9_real;
  reg        [15:0]   int_reg_array_5_9_imag;
  reg        [15:0]   int_reg_array_5_10_real;
  reg        [15:0]   int_reg_array_5_10_imag;
  reg        [15:0]   int_reg_array_5_11_real;
  reg        [15:0]   int_reg_array_5_11_imag;
  reg        [15:0]   int_reg_array_5_12_real;
  reg        [15:0]   int_reg_array_5_12_imag;
  reg        [15:0]   int_reg_array_5_13_real;
  reg        [15:0]   int_reg_array_5_13_imag;
  reg        [15:0]   int_reg_array_5_14_real;
  reg        [15:0]   int_reg_array_5_14_imag;
  reg        [15:0]   int_reg_array_5_15_real;
  reg        [15:0]   int_reg_array_5_15_imag;
  reg        [15:0]   int_reg_array_5_16_real;
  reg        [15:0]   int_reg_array_5_16_imag;
  reg        [15:0]   int_reg_array_5_17_real;
  reg        [15:0]   int_reg_array_5_17_imag;
  reg        [15:0]   int_reg_array_5_18_real;
  reg        [15:0]   int_reg_array_5_18_imag;
  reg        [15:0]   int_reg_array_5_19_real;
  reg        [15:0]   int_reg_array_5_19_imag;
  reg        [15:0]   int_reg_array_5_20_real;
  reg        [15:0]   int_reg_array_5_20_imag;
  reg        [15:0]   int_reg_array_5_21_real;
  reg        [15:0]   int_reg_array_5_21_imag;
  reg        [15:0]   int_reg_array_5_22_real;
  reg        [15:0]   int_reg_array_5_22_imag;
  reg        [15:0]   int_reg_array_5_23_real;
  reg        [15:0]   int_reg_array_5_23_imag;
  reg        [15:0]   int_reg_array_5_24_real;
  reg        [15:0]   int_reg_array_5_24_imag;
  reg        [15:0]   int_reg_array_5_25_real;
  reg        [15:0]   int_reg_array_5_25_imag;
  reg        [15:0]   int_reg_array_5_26_real;
  reg        [15:0]   int_reg_array_5_26_imag;
  reg        [15:0]   int_reg_array_5_27_real;
  reg        [15:0]   int_reg_array_5_27_imag;
  reg        [15:0]   int_reg_array_5_28_real;
  reg        [15:0]   int_reg_array_5_28_imag;
  reg        [15:0]   int_reg_array_5_29_real;
  reg        [15:0]   int_reg_array_5_29_imag;
  reg        [15:0]   int_reg_array_5_30_real;
  reg        [15:0]   int_reg_array_5_30_imag;
  reg        [15:0]   int_reg_array_5_31_real;
  reg        [15:0]   int_reg_array_5_31_imag;
  reg        [15:0]   int_reg_array_5_32_real;
  reg        [15:0]   int_reg_array_5_32_imag;
  reg        [15:0]   int_reg_array_5_33_real;
  reg        [15:0]   int_reg_array_5_33_imag;
  reg        [15:0]   int_reg_array_5_34_real;
  reg        [15:0]   int_reg_array_5_34_imag;
  reg        [15:0]   int_reg_array_5_35_real;
  reg        [15:0]   int_reg_array_5_35_imag;
  reg        [15:0]   int_reg_array_5_36_real;
  reg        [15:0]   int_reg_array_5_36_imag;
  reg        [15:0]   int_reg_array_5_37_real;
  reg        [15:0]   int_reg_array_5_37_imag;
  reg        [15:0]   int_reg_array_5_38_real;
  reg        [15:0]   int_reg_array_5_38_imag;
  reg        [15:0]   int_reg_array_5_39_real;
  reg        [15:0]   int_reg_array_5_39_imag;
  reg        [15:0]   int_reg_array_5_40_real;
  reg        [15:0]   int_reg_array_5_40_imag;
  reg        [15:0]   int_reg_array_5_41_real;
  reg        [15:0]   int_reg_array_5_41_imag;
  reg        [15:0]   int_reg_array_5_42_real;
  reg        [15:0]   int_reg_array_5_42_imag;
  reg        [15:0]   int_reg_array_5_43_real;
  reg        [15:0]   int_reg_array_5_43_imag;
  reg        [15:0]   int_reg_array_5_44_real;
  reg        [15:0]   int_reg_array_5_44_imag;
  reg        [15:0]   int_reg_array_5_45_real;
  reg        [15:0]   int_reg_array_5_45_imag;
  reg        [15:0]   int_reg_array_5_46_real;
  reg        [15:0]   int_reg_array_5_46_imag;
  reg        [15:0]   int_reg_array_5_47_real;
  reg        [15:0]   int_reg_array_5_47_imag;
  reg        [15:0]   int_reg_array_5_48_real;
  reg        [15:0]   int_reg_array_5_48_imag;
  reg        [15:0]   int_reg_array_5_49_real;
  reg        [15:0]   int_reg_array_5_49_imag;
  reg        [15:0]   int_reg_array_31_0_real;
  reg        [15:0]   int_reg_array_31_0_imag;
  reg        [15:0]   int_reg_array_31_1_real;
  reg        [15:0]   int_reg_array_31_1_imag;
  reg        [15:0]   int_reg_array_31_2_real;
  reg        [15:0]   int_reg_array_31_2_imag;
  reg        [15:0]   int_reg_array_31_3_real;
  reg        [15:0]   int_reg_array_31_3_imag;
  reg        [15:0]   int_reg_array_31_4_real;
  reg        [15:0]   int_reg_array_31_4_imag;
  reg        [15:0]   int_reg_array_31_5_real;
  reg        [15:0]   int_reg_array_31_5_imag;
  reg        [15:0]   int_reg_array_31_6_real;
  reg        [15:0]   int_reg_array_31_6_imag;
  reg        [15:0]   int_reg_array_31_7_real;
  reg        [15:0]   int_reg_array_31_7_imag;
  reg        [15:0]   int_reg_array_31_8_real;
  reg        [15:0]   int_reg_array_31_8_imag;
  reg        [15:0]   int_reg_array_31_9_real;
  reg        [15:0]   int_reg_array_31_9_imag;
  reg        [15:0]   int_reg_array_31_10_real;
  reg        [15:0]   int_reg_array_31_10_imag;
  reg        [15:0]   int_reg_array_31_11_real;
  reg        [15:0]   int_reg_array_31_11_imag;
  reg        [15:0]   int_reg_array_31_12_real;
  reg        [15:0]   int_reg_array_31_12_imag;
  reg        [15:0]   int_reg_array_31_13_real;
  reg        [15:0]   int_reg_array_31_13_imag;
  reg        [15:0]   int_reg_array_31_14_real;
  reg        [15:0]   int_reg_array_31_14_imag;
  reg        [15:0]   int_reg_array_31_15_real;
  reg        [15:0]   int_reg_array_31_15_imag;
  reg        [15:0]   int_reg_array_31_16_real;
  reg        [15:0]   int_reg_array_31_16_imag;
  reg        [15:0]   int_reg_array_31_17_real;
  reg        [15:0]   int_reg_array_31_17_imag;
  reg        [15:0]   int_reg_array_31_18_real;
  reg        [15:0]   int_reg_array_31_18_imag;
  reg        [15:0]   int_reg_array_31_19_real;
  reg        [15:0]   int_reg_array_31_19_imag;
  reg        [15:0]   int_reg_array_31_20_real;
  reg        [15:0]   int_reg_array_31_20_imag;
  reg        [15:0]   int_reg_array_31_21_real;
  reg        [15:0]   int_reg_array_31_21_imag;
  reg        [15:0]   int_reg_array_31_22_real;
  reg        [15:0]   int_reg_array_31_22_imag;
  reg        [15:0]   int_reg_array_31_23_real;
  reg        [15:0]   int_reg_array_31_23_imag;
  reg        [15:0]   int_reg_array_31_24_real;
  reg        [15:0]   int_reg_array_31_24_imag;
  reg        [15:0]   int_reg_array_31_25_real;
  reg        [15:0]   int_reg_array_31_25_imag;
  reg        [15:0]   int_reg_array_31_26_real;
  reg        [15:0]   int_reg_array_31_26_imag;
  reg        [15:0]   int_reg_array_31_27_real;
  reg        [15:0]   int_reg_array_31_27_imag;
  reg        [15:0]   int_reg_array_31_28_real;
  reg        [15:0]   int_reg_array_31_28_imag;
  reg        [15:0]   int_reg_array_31_29_real;
  reg        [15:0]   int_reg_array_31_29_imag;
  reg        [15:0]   int_reg_array_31_30_real;
  reg        [15:0]   int_reg_array_31_30_imag;
  reg        [15:0]   int_reg_array_31_31_real;
  reg        [15:0]   int_reg_array_31_31_imag;
  reg        [15:0]   int_reg_array_31_32_real;
  reg        [15:0]   int_reg_array_31_32_imag;
  reg        [15:0]   int_reg_array_31_33_real;
  reg        [15:0]   int_reg_array_31_33_imag;
  reg        [15:0]   int_reg_array_31_34_real;
  reg        [15:0]   int_reg_array_31_34_imag;
  reg        [15:0]   int_reg_array_31_35_real;
  reg        [15:0]   int_reg_array_31_35_imag;
  reg        [15:0]   int_reg_array_31_36_real;
  reg        [15:0]   int_reg_array_31_36_imag;
  reg        [15:0]   int_reg_array_31_37_real;
  reg        [15:0]   int_reg_array_31_37_imag;
  reg        [15:0]   int_reg_array_31_38_real;
  reg        [15:0]   int_reg_array_31_38_imag;
  reg        [15:0]   int_reg_array_31_39_real;
  reg        [15:0]   int_reg_array_31_39_imag;
  reg        [15:0]   int_reg_array_31_40_real;
  reg        [15:0]   int_reg_array_31_40_imag;
  reg        [15:0]   int_reg_array_31_41_real;
  reg        [15:0]   int_reg_array_31_41_imag;
  reg        [15:0]   int_reg_array_31_42_real;
  reg        [15:0]   int_reg_array_31_42_imag;
  reg        [15:0]   int_reg_array_31_43_real;
  reg        [15:0]   int_reg_array_31_43_imag;
  reg        [15:0]   int_reg_array_31_44_real;
  reg        [15:0]   int_reg_array_31_44_imag;
  reg        [15:0]   int_reg_array_31_45_real;
  reg        [15:0]   int_reg_array_31_45_imag;
  reg        [15:0]   int_reg_array_31_46_real;
  reg        [15:0]   int_reg_array_31_46_imag;
  reg        [15:0]   int_reg_array_31_47_real;
  reg        [15:0]   int_reg_array_31_47_imag;
  reg        [15:0]   int_reg_array_31_48_real;
  reg        [15:0]   int_reg_array_31_48_imag;
  reg        [15:0]   int_reg_array_31_49_real;
  reg        [15:0]   int_reg_array_31_49_imag;
  reg        [15:0]   int_reg_array_3_0_real;
  reg        [15:0]   int_reg_array_3_0_imag;
  reg        [15:0]   int_reg_array_3_1_real;
  reg        [15:0]   int_reg_array_3_1_imag;
  reg        [15:0]   int_reg_array_3_2_real;
  reg        [15:0]   int_reg_array_3_2_imag;
  reg        [15:0]   int_reg_array_3_3_real;
  reg        [15:0]   int_reg_array_3_3_imag;
  reg        [15:0]   int_reg_array_3_4_real;
  reg        [15:0]   int_reg_array_3_4_imag;
  reg        [15:0]   int_reg_array_3_5_real;
  reg        [15:0]   int_reg_array_3_5_imag;
  reg        [15:0]   int_reg_array_3_6_real;
  reg        [15:0]   int_reg_array_3_6_imag;
  reg        [15:0]   int_reg_array_3_7_real;
  reg        [15:0]   int_reg_array_3_7_imag;
  reg        [15:0]   int_reg_array_3_8_real;
  reg        [15:0]   int_reg_array_3_8_imag;
  reg        [15:0]   int_reg_array_3_9_real;
  reg        [15:0]   int_reg_array_3_9_imag;
  reg        [15:0]   int_reg_array_3_10_real;
  reg        [15:0]   int_reg_array_3_10_imag;
  reg        [15:0]   int_reg_array_3_11_real;
  reg        [15:0]   int_reg_array_3_11_imag;
  reg        [15:0]   int_reg_array_3_12_real;
  reg        [15:0]   int_reg_array_3_12_imag;
  reg        [15:0]   int_reg_array_3_13_real;
  reg        [15:0]   int_reg_array_3_13_imag;
  reg        [15:0]   int_reg_array_3_14_real;
  reg        [15:0]   int_reg_array_3_14_imag;
  reg        [15:0]   int_reg_array_3_15_real;
  reg        [15:0]   int_reg_array_3_15_imag;
  reg        [15:0]   int_reg_array_3_16_real;
  reg        [15:0]   int_reg_array_3_16_imag;
  reg        [15:0]   int_reg_array_3_17_real;
  reg        [15:0]   int_reg_array_3_17_imag;
  reg        [15:0]   int_reg_array_3_18_real;
  reg        [15:0]   int_reg_array_3_18_imag;
  reg        [15:0]   int_reg_array_3_19_real;
  reg        [15:0]   int_reg_array_3_19_imag;
  reg        [15:0]   int_reg_array_3_20_real;
  reg        [15:0]   int_reg_array_3_20_imag;
  reg        [15:0]   int_reg_array_3_21_real;
  reg        [15:0]   int_reg_array_3_21_imag;
  reg        [15:0]   int_reg_array_3_22_real;
  reg        [15:0]   int_reg_array_3_22_imag;
  reg        [15:0]   int_reg_array_3_23_real;
  reg        [15:0]   int_reg_array_3_23_imag;
  reg        [15:0]   int_reg_array_3_24_real;
  reg        [15:0]   int_reg_array_3_24_imag;
  reg        [15:0]   int_reg_array_3_25_real;
  reg        [15:0]   int_reg_array_3_25_imag;
  reg        [15:0]   int_reg_array_3_26_real;
  reg        [15:0]   int_reg_array_3_26_imag;
  reg        [15:0]   int_reg_array_3_27_real;
  reg        [15:0]   int_reg_array_3_27_imag;
  reg        [15:0]   int_reg_array_3_28_real;
  reg        [15:0]   int_reg_array_3_28_imag;
  reg        [15:0]   int_reg_array_3_29_real;
  reg        [15:0]   int_reg_array_3_29_imag;
  reg        [15:0]   int_reg_array_3_30_real;
  reg        [15:0]   int_reg_array_3_30_imag;
  reg        [15:0]   int_reg_array_3_31_real;
  reg        [15:0]   int_reg_array_3_31_imag;
  reg        [15:0]   int_reg_array_3_32_real;
  reg        [15:0]   int_reg_array_3_32_imag;
  reg        [15:0]   int_reg_array_3_33_real;
  reg        [15:0]   int_reg_array_3_33_imag;
  reg        [15:0]   int_reg_array_3_34_real;
  reg        [15:0]   int_reg_array_3_34_imag;
  reg        [15:0]   int_reg_array_3_35_real;
  reg        [15:0]   int_reg_array_3_35_imag;
  reg        [15:0]   int_reg_array_3_36_real;
  reg        [15:0]   int_reg_array_3_36_imag;
  reg        [15:0]   int_reg_array_3_37_real;
  reg        [15:0]   int_reg_array_3_37_imag;
  reg        [15:0]   int_reg_array_3_38_real;
  reg        [15:0]   int_reg_array_3_38_imag;
  reg        [15:0]   int_reg_array_3_39_real;
  reg        [15:0]   int_reg_array_3_39_imag;
  reg        [15:0]   int_reg_array_3_40_real;
  reg        [15:0]   int_reg_array_3_40_imag;
  reg        [15:0]   int_reg_array_3_41_real;
  reg        [15:0]   int_reg_array_3_41_imag;
  reg        [15:0]   int_reg_array_3_42_real;
  reg        [15:0]   int_reg_array_3_42_imag;
  reg        [15:0]   int_reg_array_3_43_real;
  reg        [15:0]   int_reg_array_3_43_imag;
  reg        [15:0]   int_reg_array_3_44_real;
  reg        [15:0]   int_reg_array_3_44_imag;
  reg        [15:0]   int_reg_array_3_45_real;
  reg        [15:0]   int_reg_array_3_45_imag;
  reg        [15:0]   int_reg_array_3_46_real;
  reg        [15:0]   int_reg_array_3_46_imag;
  reg        [15:0]   int_reg_array_3_47_real;
  reg        [15:0]   int_reg_array_3_47_imag;
  reg        [15:0]   int_reg_array_3_48_real;
  reg        [15:0]   int_reg_array_3_48_imag;
  reg        [15:0]   int_reg_array_3_49_real;
  reg        [15:0]   int_reg_array_3_49_imag;
  reg        [15:0]   int_reg_array_22_0_real;
  reg        [15:0]   int_reg_array_22_0_imag;
  reg        [15:0]   int_reg_array_22_1_real;
  reg        [15:0]   int_reg_array_22_1_imag;
  reg        [15:0]   int_reg_array_22_2_real;
  reg        [15:0]   int_reg_array_22_2_imag;
  reg        [15:0]   int_reg_array_22_3_real;
  reg        [15:0]   int_reg_array_22_3_imag;
  reg        [15:0]   int_reg_array_22_4_real;
  reg        [15:0]   int_reg_array_22_4_imag;
  reg        [15:0]   int_reg_array_22_5_real;
  reg        [15:0]   int_reg_array_22_5_imag;
  reg        [15:0]   int_reg_array_22_6_real;
  reg        [15:0]   int_reg_array_22_6_imag;
  reg        [15:0]   int_reg_array_22_7_real;
  reg        [15:0]   int_reg_array_22_7_imag;
  reg        [15:0]   int_reg_array_22_8_real;
  reg        [15:0]   int_reg_array_22_8_imag;
  reg        [15:0]   int_reg_array_22_9_real;
  reg        [15:0]   int_reg_array_22_9_imag;
  reg        [15:0]   int_reg_array_22_10_real;
  reg        [15:0]   int_reg_array_22_10_imag;
  reg        [15:0]   int_reg_array_22_11_real;
  reg        [15:0]   int_reg_array_22_11_imag;
  reg        [15:0]   int_reg_array_22_12_real;
  reg        [15:0]   int_reg_array_22_12_imag;
  reg        [15:0]   int_reg_array_22_13_real;
  reg        [15:0]   int_reg_array_22_13_imag;
  reg        [15:0]   int_reg_array_22_14_real;
  reg        [15:0]   int_reg_array_22_14_imag;
  reg        [15:0]   int_reg_array_22_15_real;
  reg        [15:0]   int_reg_array_22_15_imag;
  reg        [15:0]   int_reg_array_22_16_real;
  reg        [15:0]   int_reg_array_22_16_imag;
  reg        [15:0]   int_reg_array_22_17_real;
  reg        [15:0]   int_reg_array_22_17_imag;
  reg        [15:0]   int_reg_array_22_18_real;
  reg        [15:0]   int_reg_array_22_18_imag;
  reg        [15:0]   int_reg_array_22_19_real;
  reg        [15:0]   int_reg_array_22_19_imag;
  reg        [15:0]   int_reg_array_22_20_real;
  reg        [15:0]   int_reg_array_22_20_imag;
  reg        [15:0]   int_reg_array_22_21_real;
  reg        [15:0]   int_reg_array_22_21_imag;
  reg        [15:0]   int_reg_array_22_22_real;
  reg        [15:0]   int_reg_array_22_22_imag;
  reg        [15:0]   int_reg_array_22_23_real;
  reg        [15:0]   int_reg_array_22_23_imag;
  reg        [15:0]   int_reg_array_22_24_real;
  reg        [15:0]   int_reg_array_22_24_imag;
  reg        [15:0]   int_reg_array_22_25_real;
  reg        [15:0]   int_reg_array_22_25_imag;
  reg        [15:0]   int_reg_array_22_26_real;
  reg        [15:0]   int_reg_array_22_26_imag;
  reg        [15:0]   int_reg_array_22_27_real;
  reg        [15:0]   int_reg_array_22_27_imag;
  reg        [15:0]   int_reg_array_22_28_real;
  reg        [15:0]   int_reg_array_22_28_imag;
  reg        [15:0]   int_reg_array_22_29_real;
  reg        [15:0]   int_reg_array_22_29_imag;
  reg        [15:0]   int_reg_array_22_30_real;
  reg        [15:0]   int_reg_array_22_30_imag;
  reg        [15:0]   int_reg_array_22_31_real;
  reg        [15:0]   int_reg_array_22_31_imag;
  reg        [15:0]   int_reg_array_22_32_real;
  reg        [15:0]   int_reg_array_22_32_imag;
  reg        [15:0]   int_reg_array_22_33_real;
  reg        [15:0]   int_reg_array_22_33_imag;
  reg        [15:0]   int_reg_array_22_34_real;
  reg        [15:0]   int_reg_array_22_34_imag;
  reg        [15:0]   int_reg_array_22_35_real;
  reg        [15:0]   int_reg_array_22_35_imag;
  reg        [15:0]   int_reg_array_22_36_real;
  reg        [15:0]   int_reg_array_22_36_imag;
  reg        [15:0]   int_reg_array_22_37_real;
  reg        [15:0]   int_reg_array_22_37_imag;
  reg        [15:0]   int_reg_array_22_38_real;
  reg        [15:0]   int_reg_array_22_38_imag;
  reg        [15:0]   int_reg_array_22_39_real;
  reg        [15:0]   int_reg_array_22_39_imag;
  reg        [15:0]   int_reg_array_22_40_real;
  reg        [15:0]   int_reg_array_22_40_imag;
  reg        [15:0]   int_reg_array_22_41_real;
  reg        [15:0]   int_reg_array_22_41_imag;
  reg        [15:0]   int_reg_array_22_42_real;
  reg        [15:0]   int_reg_array_22_42_imag;
  reg        [15:0]   int_reg_array_22_43_real;
  reg        [15:0]   int_reg_array_22_43_imag;
  reg        [15:0]   int_reg_array_22_44_real;
  reg        [15:0]   int_reg_array_22_44_imag;
  reg        [15:0]   int_reg_array_22_45_real;
  reg        [15:0]   int_reg_array_22_45_imag;
  reg        [15:0]   int_reg_array_22_46_real;
  reg        [15:0]   int_reg_array_22_46_imag;
  reg        [15:0]   int_reg_array_22_47_real;
  reg        [15:0]   int_reg_array_22_47_imag;
  reg        [15:0]   int_reg_array_22_48_real;
  reg        [15:0]   int_reg_array_22_48_imag;
  reg        [15:0]   int_reg_array_22_49_real;
  reg        [15:0]   int_reg_array_22_49_imag;
  reg        [15:0]   int_reg_array_11_0_real;
  reg        [15:0]   int_reg_array_11_0_imag;
  reg        [15:0]   int_reg_array_11_1_real;
  reg        [15:0]   int_reg_array_11_1_imag;
  reg        [15:0]   int_reg_array_11_2_real;
  reg        [15:0]   int_reg_array_11_2_imag;
  reg        [15:0]   int_reg_array_11_3_real;
  reg        [15:0]   int_reg_array_11_3_imag;
  reg        [15:0]   int_reg_array_11_4_real;
  reg        [15:0]   int_reg_array_11_4_imag;
  reg        [15:0]   int_reg_array_11_5_real;
  reg        [15:0]   int_reg_array_11_5_imag;
  reg        [15:0]   int_reg_array_11_6_real;
  reg        [15:0]   int_reg_array_11_6_imag;
  reg        [15:0]   int_reg_array_11_7_real;
  reg        [15:0]   int_reg_array_11_7_imag;
  reg        [15:0]   int_reg_array_11_8_real;
  reg        [15:0]   int_reg_array_11_8_imag;
  reg        [15:0]   int_reg_array_11_9_real;
  reg        [15:0]   int_reg_array_11_9_imag;
  reg        [15:0]   int_reg_array_11_10_real;
  reg        [15:0]   int_reg_array_11_10_imag;
  reg        [15:0]   int_reg_array_11_11_real;
  reg        [15:0]   int_reg_array_11_11_imag;
  reg        [15:0]   int_reg_array_11_12_real;
  reg        [15:0]   int_reg_array_11_12_imag;
  reg        [15:0]   int_reg_array_11_13_real;
  reg        [15:0]   int_reg_array_11_13_imag;
  reg        [15:0]   int_reg_array_11_14_real;
  reg        [15:0]   int_reg_array_11_14_imag;
  reg        [15:0]   int_reg_array_11_15_real;
  reg        [15:0]   int_reg_array_11_15_imag;
  reg        [15:0]   int_reg_array_11_16_real;
  reg        [15:0]   int_reg_array_11_16_imag;
  reg        [15:0]   int_reg_array_11_17_real;
  reg        [15:0]   int_reg_array_11_17_imag;
  reg        [15:0]   int_reg_array_11_18_real;
  reg        [15:0]   int_reg_array_11_18_imag;
  reg        [15:0]   int_reg_array_11_19_real;
  reg        [15:0]   int_reg_array_11_19_imag;
  reg        [15:0]   int_reg_array_11_20_real;
  reg        [15:0]   int_reg_array_11_20_imag;
  reg        [15:0]   int_reg_array_11_21_real;
  reg        [15:0]   int_reg_array_11_21_imag;
  reg        [15:0]   int_reg_array_11_22_real;
  reg        [15:0]   int_reg_array_11_22_imag;
  reg        [15:0]   int_reg_array_11_23_real;
  reg        [15:0]   int_reg_array_11_23_imag;
  reg        [15:0]   int_reg_array_11_24_real;
  reg        [15:0]   int_reg_array_11_24_imag;
  reg        [15:0]   int_reg_array_11_25_real;
  reg        [15:0]   int_reg_array_11_25_imag;
  reg        [15:0]   int_reg_array_11_26_real;
  reg        [15:0]   int_reg_array_11_26_imag;
  reg        [15:0]   int_reg_array_11_27_real;
  reg        [15:0]   int_reg_array_11_27_imag;
  reg        [15:0]   int_reg_array_11_28_real;
  reg        [15:0]   int_reg_array_11_28_imag;
  reg        [15:0]   int_reg_array_11_29_real;
  reg        [15:0]   int_reg_array_11_29_imag;
  reg        [15:0]   int_reg_array_11_30_real;
  reg        [15:0]   int_reg_array_11_30_imag;
  reg        [15:0]   int_reg_array_11_31_real;
  reg        [15:0]   int_reg_array_11_31_imag;
  reg        [15:0]   int_reg_array_11_32_real;
  reg        [15:0]   int_reg_array_11_32_imag;
  reg        [15:0]   int_reg_array_11_33_real;
  reg        [15:0]   int_reg_array_11_33_imag;
  reg        [15:0]   int_reg_array_11_34_real;
  reg        [15:0]   int_reg_array_11_34_imag;
  reg        [15:0]   int_reg_array_11_35_real;
  reg        [15:0]   int_reg_array_11_35_imag;
  reg        [15:0]   int_reg_array_11_36_real;
  reg        [15:0]   int_reg_array_11_36_imag;
  reg        [15:0]   int_reg_array_11_37_real;
  reg        [15:0]   int_reg_array_11_37_imag;
  reg        [15:0]   int_reg_array_11_38_real;
  reg        [15:0]   int_reg_array_11_38_imag;
  reg        [15:0]   int_reg_array_11_39_real;
  reg        [15:0]   int_reg_array_11_39_imag;
  reg        [15:0]   int_reg_array_11_40_real;
  reg        [15:0]   int_reg_array_11_40_imag;
  reg        [15:0]   int_reg_array_11_41_real;
  reg        [15:0]   int_reg_array_11_41_imag;
  reg        [15:0]   int_reg_array_11_42_real;
  reg        [15:0]   int_reg_array_11_42_imag;
  reg        [15:0]   int_reg_array_11_43_real;
  reg        [15:0]   int_reg_array_11_43_imag;
  reg        [15:0]   int_reg_array_11_44_real;
  reg        [15:0]   int_reg_array_11_44_imag;
  reg        [15:0]   int_reg_array_11_45_real;
  reg        [15:0]   int_reg_array_11_45_imag;
  reg        [15:0]   int_reg_array_11_46_real;
  reg        [15:0]   int_reg_array_11_46_imag;
  reg        [15:0]   int_reg_array_11_47_real;
  reg        [15:0]   int_reg_array_11_47_imag;
  reg        [15:0]   int_reg_array_11_48_real;
  reg        [15:0]   int_reg_array_11_48_imag;
  reg        [15:0]   int_reg_array_11_49_real;
  reg        [15:0]   int_reg_array_11_49_imag;
  reg        [15:0]   int_reg_array_41_0_real;
  reg        [15:0]   int_reg_array_41_0_imag;
  reg        [15:0]   int_reg_array_41_1_real;
  reg        [15:0]   int_reg_array_41_1_imag;
  reg        [15:0]   int_reg_array_41_2_real;
  reg        [15:0]   int_reg_array_41_2_imag;
  reg        [15:0]   int_reg_array_41_3_real;
  reg        [15:0]   int_reg_array_41_3_imag;
  reg        [15:0]   int_reg_array_41_4_real;
  reg        [15:0]   int_reg_array_41_4_imag;
  reg        [15:0]   int_reg_array_41_5_real;
  reg        [15:0]   int_reg_array_41_5_imag;
  reg        [15:0]   int_reg_array_41_6_real;
  reg        [15:0]   int_reg_array_41_6_imag;
  reg        [15:0]   int_reg_array_41_7_real;
  reg        [15:0]   int_reg_array_41_7_imag;
  reg        [15:0]   int_reg_array_41_8_real;
  reg        [15:0]   int_reg_array_41_8_imag;
  reg        [15:0]   int_reg_array_41_9_real;
  reg        [15:0]   int_reg_array_41_9_imag;
  reg        [15:0]   int_reg_array_41_10_real;
  reg        [15:0]   int_reg_array_41_10_imag;
  reg        [15:0]   int_reg_array_41_11_real;
  reg        [15:0]   int_reg_array_41_11_imag;
  reg        [15:0]   int_reg_array_41_12_real;
  reg        [15:0]   int_reg_array_41_12_imag;
  reg        [15:0]   int_reg_array_41_13_real;
  reg        [15:0]   int_reg_array_41_13_imag;
  reg        [15:0]   int_reg_array_41_14_real;
  reg        [15:0]   int_reg_array_41_14_imag;
  reg        [15:0]   int_reg_array_41_15_real;
  reg        [15:0]   int_reg_array_41_15_imag;
  reg        [15:0]   int_reg_array_41_16_real;
  reg        [15:0]   int_reg_array_41_16_imag;
  reg        [15:0]   int_reg_array_41_17_real;
  reg        [15:0]   int_reg_array_41_17_imag;
  reg        [15:0]   int_reg_array_41_18_real;
  reg        [15:0]   int_reg_array_41_18_imag;
  reg        [15:0]   int_reg_array_41_19_real;
  reg        [15:0]   int_reg_array_41_19_imag;
  reg        [15:0]   int_reg_array_41_20_real;
  reg        [15:0]   int_reg_array_41_20_imag;
  reg        [15:0]   int_reg_array_41_21_real;
  reg        [15:0]   int_reg_array_41_21_imag;
  reg        [15:0]   int_reg_array_41_22_real;
  reg        [15:0]   int_reg_array_41_22_imag;
  reg        [15:0]   int_reg_array_41_23_real;
  reg        [15:0]   int_reg_array_41_23_imag;
  reg        [15:0]   int_reg_array_41_24_real;
  reg        [15:0]   int_reg_array_41_24_imag;
  reg        [15:0]   int_reg_array_41_25_real;
  reg        [15:0]   int_reg_array_41_25_imag;
  reg        [15:0]   int_reg_array_41_26_real;
  reg        [15:0]   int_reg_array_41_26_imag;
  reg        [15:0]   int_reg_array_41_27_real;
  reg        [15:0]   int_reg_array_41_27_imag;
  reg        [15:0]   int_reg_array_41_28_real;
  reg        [15:0]   int_reg_array_41_28_imag;
  reg        [15:0]   int_reg_array_41_29_real;
  reg        [15:0]   int_reg_array_41_29_imag;
  reg        [15:0]   int_reg_array_41_30_real;
  reg        [15:0]   int_reg_array_41_30_imag;
  reg        [15:0]   int_reg_array_41_31_real;
  reg        [15:0]   int_reg_array_41_31_imag;
  reg        [15:0]   int_reg_array_41_32_real;
  reg        [15:0]   int_reg_array_41_32_imag;
  reg        [15:0]   int_reg_array_41_33_real;
  reg        [15:0]   int_reg_array_41_33_imag;
  reg        [15:0]   int_reg_array_41_34_real;
  reg        [15:0]   int_reg_array_41_34_imag;
  reg        [15:0]   int_reg_array_41_35_real;
  reg        [15:0]   int_reg_array_41_35_imag;
  reg        [15:0]   int_reg_array_41_36_real;
  reg        [15:0]   int_reg_array_41_36_imag;
  reg        [15:0]   int_reg_array_41_37_real;
  reg        [15:0]   int_reg_array_41_37_imag;
  reg        [15:0]   int_reg_array_41_38_real;
  reg        [15:0]   int_reg_array_41_38_imag;
  reg        [15:0]   int_reg_array_41_39_real;
  reg        [15:0]   int_reg_array_41_39_imag;
  reg        [15:0]   int_reg_array_41_40_real;
  reg        [15:0]   int_reg_array_41_40_imag;
  reg        [15:0]   int_reg_array_41_41_real;
  reg        [15:0]   int_reg_array_41_41_imag;
  reg        [15:0]   int_reg_array_41_42_real;
  reg        [15:0]   int_reg_array_41_42_imag;
  reg        [15:0]   int_reg_array_41_43_real;
  reg        [15:0]   int_reg_array_41_43_imag;
  reg        [15:0]   int_reg_array_41_44_real;
  reg        [15:0]   int_reg_array_41_44_imag;
  reg        [15:0]   int_reg_array_41_45_real;
  reg        [15:0]   int_reg_array_41_45_imag;
  reg        [15:0]   int_reg_array_41_46_real;
  reg        [15:0]   int_reg_array_41_46_imag;
  reg        [15:0]   int_reg_array_41_47_real;
  reg        [15:0]   int_reg_array_41_47_imag;
  reg        [15:0]   int_reg_array_41_48_real;
  reg        [15:0]   int_reg_array_41_48_imag;
  reg        [15:0]   int_reg_array_41_49_real;
  reg        [15:0]   int_reg_array_41_49_imag;
  reg        [15:0]   int_reg_array_10_0_real;
  reg        [15:0]   int_reg_array_10_0_imag;
  reg        [15:0]   int_reg_array_10_1_real;
  reg        [15:0]   int_reg_array_10_1_imag;
  reg        [15:0]   int_reg_array_10_2_real;
  reg        [15:0]   int_reg_array_10_2_imag;
  reg        [15:0]   int_reg_array_10_3_real;
  reg        [15:0]   int_reg_array_10_3_imag;
  reg        [15:0]   int_reg_array_10_4_real;
  reg        [15:0]   int_reg_array_10_4_imag;
  reg        [15:0]   int_reg_array_10_5_real;
  reg        [15:0]   int_reg_array_10_5_imag;
  reg        [15:0]   int_reg_array_10_6_real;
  reg        [15:0]   int_reg_array_10_6_imag;
  reg        [15:0]   int_reg_array_10_7_real;
  reg        [15:0]   int_reg_array_10_7_imag;
  reg        [15:0]   int_reg_array_10_8_real;
  reg        [15:0]   int_reg_array_10_8_imag;
  reg        [15:0]   int_reg_array_10_9_real;
  reg        [15:0]   int_reg_array_10_9_imag;
  reg        [15:0]   int_reg_array_10_10_real;
  reg        [15:0]   int_reg_array_10_10_imag;
  reg        [15:0]   int_reg_array_10_11_real;
  reg        [15:0]   int_reg_array_10_11_imag;
  reg        [15:0]   int_reg_array_10_12_real;
  reg        [15:0]   int_reg_array_10_12_imag;
  reg        [15:0]   int_reg_array_10_13_real;
  reg        [15:0]   int_reg_array_10_13_imag;
  reg        [15:0]   int_reg_array_10_14_real;
  reg        [15:0]   int_reg_array_10_14_imag;
  reg        [15:0]   int_reg_array_10_15_real;
  reg        [15:0]   int_reg_array_10_15_imag;
  reg        [15:0]   int_reg_array_10_16_real;
  reg        [15:0]   int_reg_array_10_16_imag;
  reg        [15:0]   int_reg_array_10_17_real;
  reg        [15:0]   int_reg_array_10_17_imag;
  reg        [15:0]   int_reg_array_10_18_real;
  reg        [15:0]   int_reg_array_10_18_imag;
  reg        [15:0]   int_reg_array_10_19_real;
  reg        [15:0]   int_reg_array_10_19_imag;
  reg        [15:0]   int_reg_array_10_20_real;
  reg        [15:0]   int_reg_array_10_20_imag;
  reg        [15:0]   int_reg_array_10_21_real;
  reg        [15:0]   int_reg_array_10_21_imag;
  reg        [15:0]   int_reg_array_10_22_real;
  reg        [15:0]   int_reg_array_10_22_imag;
  reg        [15:0]   int_reg_array_10_23_real;
  reg        [15:0]   int_reg_array_10_23_imag;
  reg        [15:0]   int_reg_array_10_24_real;
  reg        [15:0]   int_reg_array_10_24_imag;
  reg        [15:0]   int_reg_array_10_25_real;
  reg        [15:0]   int_reg_array_10_25_imag;
  reg        [15:0]   int_reg_array_10_26_real;
  reg        [15:0]   int_reg_array_10_26_imag;
  reg        [15:0]   int_reg_array_10_27_real;
  reg        [15:0]   int_reg_array_10_27_imag;
  reg        [15:0]   int_reg_array_10_28_real;
  reg        [15:0]   int_reg_array_10_28_imag;
  reg        [15:0]   int_reg_array_10_29_real;
  reg        [15:0]   int_reg_array_10_29_imag;
  reg        [15:0]   int_reg_array_10_30_real;
  reg        [15:0]   int_reg_array_10_30_imag;
  reg        [15:0]   int_reg_array_10_31_real;
  reg        [15:0]   int_reg_array_10_31_imag;
  reg        [15:0]   int_reg_array_10_32_real;
  reg        [15:0]   int_reg_array_10_32_imag;
  reg        [15:0]   int_reg_array_10_33_real;
  reg        [15:0]   int_reg_array_10_33_imag;
  reg        [15:0]   int_reg_array_10_34_real;
  reg        [15:0]   int_reg_array_10_34_imag;
  reg        [15:0]   int_reg_array_10_35_real;
  reg        [15:0]   int_reg_array_10_35_imag;
  reg        [15:0]   int_reg_array_10_36_real;
  reg        [15:0]   int_reg_array_10_36_imag;
  reg        [15:0]   int_reg_array_10_37_real;
  reg        [15:0]   int_reg_array_10_37_imag;
  reg        [15:0]   int_reg_array_10_38_real;
  reg        [15:0]   int_reg_array_10_38_imag;
  reg        [15:0]   int_reg_array_10_39_real;
  reg        [15:0]   int_reg_array_10_39_imag;
  reg        [15:0]   int_reg_array_10_40_real;
  reg        [15:0]   int_reg_array_10_40_imag;
  reg        [15:0]   int_reg_array_10_41_real;
  reg        [15:0]   int_reg_array_10_41_imag;
  reg        [15:0]   int_reg_array_10_42_real;
  reg        [15:0]   int_reg_array_10_42_imag;
  reg        [15:0]   int_reg_array_10_43_real;
  reg        [15:0]   int_reg_array_10_43_imag;
  reg        [15:0]   int_reg_array_10_44_real;
  reg        [15:0]   int_reg_array_10_44_imag;
  reg        [15:0]   int_reg_array_10_45_real;
  reg        [15:0]   int_reg_array_10_45_imag;
  reg        [15:0]   int_reg_array_10_46_real;
  reg        [15:0]   int_reg_array_10_46_imag;
  reg        [15:0]   int_reg_array_10_47_real;
  reg        [15:0]   int_reg_array_10_47_imag;
  reg        [15:0]   int_reg_array_10_48_real;
  reg        [15:0]   int_reg_array_10_48_imag;
  reg        [15:0]   int_reg_array_10_49_real;
  reg        [15:0]   int_reg_array_10_49_imag;
  reg        [15:0]   int_reg_array_14_0_real;
  reg        [15:0]   int_reg_array_14_0_imag;
  reg        [15:0]   int_reg_array_14_1_real;
  reg        [15:0]   int_reg_array_14_1_imag;
  reg        [15:0]   int_reg_array_14_2_real;
  reg        [15:0]   int_reg_array_14_2_imag;
  reg        [15:0]   int_reg_array_14_3_real;
  reg        [15:0]   int_reg_array_14_3_imag;
  reg        [15:0]   int_reg_array_14_4_real;
  reg        [15:0]   int_reg_array_14_4_imag;
  reg        [15:0]   int_reg_array_14_5_real;
  reg        [15:0]   int_reg_array_14_5_imag;
  reg        [15:0]   int_reg_array_14_6_real;
  reg        [15:0]   int_reg_array_14_6_imag;
  reg        [15:0]   int_reg_array_14_7_real;
  reg        [15:0]   int_reg_array_14_7_imag;
  reg        [15:0]   int_reg_array_14_8_real;
  reg        [15:0]   int_reg_array_14_8_imag;
  reg        [15:0]   int_reg_array_14_9_real;
  reg        [15:0]   int_reg_array_14_9_imag;
  reg        [15:0]   int_reg_array_14_10_real;
  reg        [15:0]   int_reg_array_14_10_imag;
  reg        [15:0]   int_reg_array_14_11_real;
  reg        [15:0]   int_reg_array_14_11_imag;
  reg        [15:0]   int_reg_array_14_12_real;
  reg        [15:0]   int_reg_array_14_12_imag;
  reg        [15:0]   int_reg_array_14_13_real;
  reg        [15:0]   int_reg_array_14_13_imag;
  reg        [15:0]   int_reg_array_14_14_real;
  reg        [15:0]   int_reg_array_14_14_imag;
  reg        [15:0]   int_reg_array_14_15_real;
  reg        [15:0]   int_reg_array_14_15_imag;
  reg        [15:0]   int_reg_array_14_16_real;
  reg        [15:0]   int_reg_array_14_16_imag;
  reg        [15:0]   int_reg_array_14_17_real;
  reg        [15:0]   int_reg_array_14_17_imag;
  reg        [15:0]   int_reg_array_14_18_real;
  reg        [15:0]   int_reg_array_14_18_imag;
  reg        [15:0]   int_reg_array_14_19_real;
  reg        [15:0]   int_reg_array_14_19_imag;
  reg        [15:0]   int_reg_array_14_20_real;
  reg        [15:0]   int_reg_array_14_20_imag;
  reg        [15:0]   int_reg_array_14_21_real;
  reg        [15:0]   int_reg_array_14_21_imag;
  reg        [15:0]   int_reg_array_14_22_real;
  reg        [15:0]   int_reg_array_14_22_imag;
  reg        [15:0]   int_reg_array_14_23_real;
  reg        [15:0]   int_reg_array_14_23_imag;
  reg        [15:0]   int_reg_array_14_24_real;
  reg        [15:0]   int_reg_array_14_24_imag;
  reg        [15:0]   int_reg_array_14_25_real;
  reg        [15:0]   int_reg_array_14_25_imag;
  reg        [15:0]   int_reg_array_14_26_real;
  reg        [15:0]   int_reg_array_14_26_imag;
  reg        [15:0]   int_reg_array_14_27_real;
  reg        [15:0]   int_reg_array_14_27_imag;
  reg        [15:0]   int_reg_array_14_28_real;
  reg        [15:0]   int_reg_array_14_28_imag;
  reg        [15:0]   int_reg_array_14_29_real;
  reg        [15:0]   int_reg_array_14_29_imag;
  reg        [15:0]   int_reg_array_14_30_real;
  reg        [15:0]   int_reg_array_14_30_imag;
  reg        [15:0]   int_reg_array_14_31_real;
  reg        [15:0]   int_reg_array_14_31_imag;
  reg        [15:0]   int_reg_array_14_32_real;
  reg        [15:0]   int_reg_array_14_32_imag;
  reg        [15:0]   int_reg_array_14_33_real;
  reg        [15:0]   int_reg_array_14_33_imag;
  reg        [15:0]   int_reg_array_14_34_real;
  reg        [15:0]   int_reg_array_14_34_imag;
  reg        [15:0]   int_reg_array_14_35_real;
  reg        [15:0]   int_reg_array_14_35_imag;
  reg        [15:0]   int_reg_array_14_36_real;
  reg        [15:0]   int_reg_array_14_36_imag;
  reg        [15:0]   int_reg_array_14_37_real;
  reg        [15:0]   int_reg_array_14_37_imag;
  reg        [15:0]   int_reg_array_14_38_real;
  reg        [15:0]   int_reg_array_14_38_imag;
  reg        [15:0]   int_reg_array_14_39_real;
  reg        [15:0]   int_reg_array_14_39_imag;
  reg        [15:0]   int_reg_array_14_40_real;
  reg        [15:0]   int_reg_array_14_40_imag;
  reg        [15:0]   int_reg_array_14_41_real;
  reg        [15:0]   int_reg_array_14_41_imag;
  reg        [15:0]   int_reg_array_14_42_real;
  reg        [15:0]   int_reg_array_14_42_imag;
  reg        [15:0]   int_reg_array_14_43_real;
  reg        [15:0]   int_reg_array_14_43_imag;
  reg        [15:0]   int_reg_array_14_44_real;
  reg        [15:0]   int_reg_array_14_44_imag;
  reg        [15:0]   int_reg_array_14_45_real;
  reg        [15:0]   int_reg_array_14_45_imag;
  reg        [15:0]   int_reg_array_14_46_real;
  reg        [15:0]   int_reg_array_14_46_imag;
  reg        [15:0]   int_reg_array_14_47_real;
  reg        [15:0]   int_reg_array_14_47_imag;
  reg        [15:0]   int_reg_array_14_48_real;
  reg        [15:0]   int_reg_array_14_48_imag;
  reg        [15:0]   int_reg_array_14_49_real;
  reg        [15:0]   int_reg_array_14_49_imag;
  reg        [15:0]   int_reg_array_19_0_real;
  reg        [15:0]   int_reg_array_19_0_imag;
  reg        [15:0]   int_reg_array_19_1_real;
  reg        [15:0]   int_reg_array_19_1_imag;
  reg        [15:0]   int_reg_array_19_2_real;
  reg        [15:0]   int_reg_array_19_2_imag;
  reg        [15:0]   int_reg_array_19_3_real;
  reg        [15:0]   int_reg_array_19_3_imag;
  reg        [15:0]   int_reg_array_19_4_real;
  reg        [15:0]   int_reg_array_19_4_imag;
  reg        [15:0]   int_reg_array_19_5_real;
  reg        [15:0]   int_reg_array_19_5_imag;
  reg        [15:0]   int_reg_array_19_6_real;
  reg        [15:0]   int_reg_array_19_6_imag;
  reg        [15:0]   int_reg_array_19_7_real;
  reg        [15:0]   int_reg_array_19_7_imag;
  reg        [15:0]   int_reg_array_19_8_real;
  reg        [15:0]   int_reg_array_19_8_imag;
  reg        [15:0]   int_reg_array_19_9_real;
  reg        [15:0]   int_reg_array_19_9_imag;
  reg        [15:0]   int_reg_array_19_10_real;
  reg        [15:0]   int_reg_array_19_10_imag;
  reg        [15:0]   int_reg_array_19_11_real;
  reg        [15:0]   int_reg_array_19_11_imag;
  reg        [15:0]   int_reg_array_19_12_real;
  reg        [15:0]   int_reg_array_19_12_imag;
  reg        [15:0]   int_reg_array_19_13_real;
  reg        [15:0]   int_reg_array_19_13_imag;
  reg        [15:0]   int_reg_array_19_14_real;
  reg        [15:0]   int_reg_array_19_14_imag;
  reg        [15:0]   int_reg_array_19_15_real;
  reg        [15:0]   int_reg_array_19_15_imag;
  reg        [15:0]   int_reg_array_19_16_real;
  reg        [15:0]   int_reg_array_19_16_imag;
  reg        [15:0]   int_reg_array_19_17_real;
  reg        [15:0]   int_reg_array_19_17_imag;
  reg        [15:0]   int_reg_array_19_18_real;
  reg        [15:0]   int_reg_array_19_18_imag;
  reg        [15:0]   int_reg_array_19_19_real;
  reg        [15:0]   int_reg_array_19_19_imag;
  reg        [15:0]   int_reg_array_19_20_real;
  reg        [15:0]   int_reg_array_19_20_imag;
  reg        [15:0]   int_reg_array_19_21_real;
  reg        [15:0]   int_reg_array_19_21_imag;
  reg        [15:0]   int_reg_array_19_22_real;
  reg        [15:0]   int_reg_array_19_22_imag;
  reg        [15:0]   int_reg_array_19_23_real;
  reg        [15:0]   int_reg_array_19_23_imag;
  reg        [15:0]   int_reg_array_19_24_real;
  reg        [15:0]   int_reg_array_19_24_imag;
  reg        [15:0]   int_reg_array_19_25_real;
  reg        [15:0]   int_reg_array_19_25_imag;
  reg        [15:0]   int_reg_array_19_26_real;
  reg        [15:0]   int_reg_array_19_26_imag;
  reg        [15:0]   int_reg_array_19_27_real;
  reg        [15:0]   int_reg_array_19_27_imag;
  reg        [15:0]   int_reg_array_19_28_real;
  reg        [15:0]   int_reg_array_19_28_imag;
  reg        [15:0]   int_reg_array_19_29_real;
  reg        [15:0]   int_reg_array_19_29_imag;
  reg        [15:0]   int_reg_array_19_30_real;
  reg        [15:0]   int_reg_array_19_30_imag;
  reg        [15:0]   int_reg_array_19_31_real;
  reg        [15:0]   int_reg_array_19_31_imag;
  reg        [15:0]   int_reg_array_19_32_real;
  reg        [15:0]   int_reg_array_19_32_imag;
  reg        [15:0]   int_reg_array_19_33_real;
  reg        [15:0]   int_reg_array_19_33_imag;
  reg        [15:0]   int_reg_array_19_34_real;
  reg        [15:0]   int_reg_array_19_34_imag;
  reg        [15:0]   int_reg_array_19_35_real;
  reg        [15:0]   int_reg_array_19_35_imag;
  reg        [15:0]   int_reg_array_19_36_real;
  reg        [15:0]   int_reg_array_19_36_imag;
  reg        [15:0]   int_reg_array_19_37_real;
  reg        [15:0]   int_reg_array_19_37_imag;
  reg        [15:0]   int_reg_array_19_38_real;
  reg        [15:0]   int_reg_array_19_38_imag;
  reg        [15:0]   int_reg_array_19_39_real;
  reg        [15:0]   int_reg_array_19_39_imag;
  reg        [15:0]   int_reg_array_19_40_real;
  reg        [15:0]   int_reg_array_19_40_imag;
  reg        [15:0]   int_reg_array_19_41_real;
  reg        [15:0]   int_reg_array_19_41_imag;
  reg        [15:0]   int_reg_array_19_42_real;
  reg        [15:0]   int_reg_array_19_42_imag;
  reg        [15:0]   int_reg_array_19_43_real;
  reg        [15:0]   int_reg_array_19_43_imag;
  reg        [15:0]   int_reg_array_19_44_real;
  reg        [15:0]   int_reg_array_19_44_imag;
  reg        [15:0]   int_reg_array_19_45_real;
  reg        [15:0]   int_reg_array_19_45_imag;
  reg        [15:0]   int_reg_array_19_46_real;
  reg        [15:0]   int_reg_array_19_46_imag;
  reg        [15:0]   int_reg_array_19_47_real;
  reg        [15:0]   int_reg_array_19_47_imag;
  reg        [15:0]   int_reg_array_19_48_real;
  reg        [15:0]   int_reg_array_19_48_imag;
  reg        [15:0]   int_reg_array_19_49_real;
  reg        [15:0]   int_reg_array_19_49_imag;
  reg        [15:0]   int_reg_array_42_0_real;
  reg        [15:0]   int_reg_array_42_0_imag;
  reg        [15:0]   int_reg_array_42_1_real;
  reg        [15:0]   int_reg_array_42_1_imag;
  reg        [15:0]   int_reg_array_42_2_real;
  reg        [15:0]   int_reg_array_42_2_imag;
  reg        [15:0]   int_reg_array_42_3_real;
  reg        [15:0]   int_reg_array_42_3_imag;
  reg        [15:0]   int_reg_array_42_4_real;
  reg        [15:0]   int_reg_array_42_4_imag;
  reg        [15:0]   int_reg_array_42_5_real;
  reg        [15:0]   int_reg_array_42_5_imag;
  reg        [15:0]   int_reg_array_42_6_real;
  reg        [15:0]   int_reg_array_42_6_imag;
  reg        [15:0]   int_reg_array_42_7_real;
  reg        [15:0]   int_reg_array_42_7_imag;
  reg        [15:0]   int_reg_array_42_8_real;
  reg        [15:0]   int_reg_array_42_8_imag;
  reg        [15:0]   int_reg_array_42_9_real;
  reg        [15:0]   int_reg_array_42_9_imag;
  reg        [15:0]   int_reg_array_42_10_real;
  reg        [15:0]   int_reg_array_42_10_imag;
  reg        [15:0]   int_reg_array_42_11_real;
  reg        [15:0]   int_reg_array_42_11_imag;
  reg        [15:0]   int_reg_array_42_12_real;
  reg        [15:0]   int_reg_array_42_12_imag;
  reg        [15:0]   int_reg_array_42_13_real;
  reg        [15:0]   int_reg_array_42_13_imag;
  reg        [15:0]   int_reg_array_42_14_real;
  reg        [15:0]   int_reg_array_42_14_imag;
  reg        [15:0]   int_reg_array_42_15_real;
  reg        [15:0]   int_reg_array_42_15_imag;
  reg        [15:0]   int_reg_array_42_16_real;
  reg        [15:0]   int_reg_array_42_16_imag;
  reg        [15:0]   int_reg_array_42_17_real;
  reg        [15:0]   int_reg_array_42_17_imag;
  reg        [15:0]   int_reg_array_42_18_real;
  reg        [15:0]   int_reg_array_42_18_imag;
  reg        [15:0]   int_reg_array_42_19_real;
  reg        [15:0]   int_reg_array_42_19_imag;
  reg        [15:0]   int_reg_array_42_20_real;
  reg        [15:0]   int_reg_array_42_20_imag;
  reg        [15:0]   int_reg_array_42_21_real;
  reg        [15:0]   int_reg_array_42_21_imag;
  reg        [15:0]   int_reg_array_42_22_real;
  reg        [15:0]   int_reg_array_42_22_imag;
  reg        [15:0]   int_reg_array_42_23_real;
  reg        [15:0]   int_reg_array_42_23_imag;
  reg        [15:0]   int_reg_array_42_24_real;
  reg        [15:0]   int_reg_array_42_24_imag;
  reg        [15:0]   int_reg_array_42_25_real;
  reg        [15:0]   int_reg_array_42_25_imag;
  reg        [15:0]   int_reg_array_42_26_real;
  reg        [15:0]   int_reg_array_42_26_imag;
  reg        [15:0]   int_reg_array_42_27_real;
  reg        [15:0]   int_reg_array_42_27_imag;
  reg        [15:0]   int_reg_array_42_28_real;
  reg        [15:0]   int_reg_array_42_28_imag;
  reg        [15:0]   int_reg_array_42_29_real;
  reg        [15:0]   int_reg_array_42_29_imag;
  reg        [15:0]   int_reg_array_42_30_real;
  reg        [15:0]   int_reg_array_42_30_imag;
  reg        [15:0]   int_reg_array_42_31_real;
  reg        [15:0]   int_reg_array_42_31_imag;
  reg        [15:0]   int_reg_array_42_32_real;
  reg        [15:0]   int_reg_array_42_32_imag;
  reg        [15:0]   int_reg_array_42_33_real;
  reg        [15:0]   int_reg_array_42_33_imag;
  reg        [15:0]   int_reg_array_42_34_real;
  reg        [15:0]   int_reg_array_42_34_imag;
  reg        [15:0]   int_reg_array_42_35_real;
  reg        [15:0]   int_reg_array_42_35_imag;
  reg        [15:0]   int_reg_array_42_36_real;
  reg        [15:0]   int_reg_array_42_36_imag;
  reg        [15:0]   int_reg_array_42_37_real;
  reg        [15:0]   int_reg_array_42_37_imag;
  reg        [15:0]   int_reg_array_42_38_real;
  reg        [15:0]   int_reg_array_42_38_imag;
  reg        [15:0]   int_reg_array_42_39_real;
  reg        [15:0]   int_reg_array_42_39_imag;
  reg        [15:0]   int_reg_array_42_40_real;
  reg        [15:0]   int_reg_array_42_40_imag;
  reg        [15:0]   int_reg_array_42_41_real;
  reg        [15:0]   int_reg_array_42_41_imag;
  reg        [15:0]   int_reg_array_42_42_real;
  reg        [15:0]   int_reg_array_42_42_imag;
  reg        [15:0]   int_reg_array_42_43_real;
  reg        [15:0]   int_reg_array_42_43_imag;
  reg        [15:0]   int_reg_array_42_44_real;
  reg        [15:0]   int_reg_array_42_44_imag;
  reg        [15:0]   int_reg_array_42_45_real;
  reg        [15:0]   int_reg_array_42_45_imag;
  reg        [15:0]   int_reg_array_42_46_real;
  reg        [15:0]   int_reg_array_42_46_imag;
  reg        [15:0]   int_reg_array_42_47_real;
  reg        [15:0]   int_reg_array_42_47_imag;
  reg        [15:0]   int_reg_array_42_48_real;
  reg        [15:0]   int_reg_array_42_48_imag;
  reg        [15:0]   int_reg_array_42_49_real;
  reg        [15:0]   int_reg_array_42_49_imag;
  reg        [15:0]   int_reg_array_18_0_real;
  reg        [15:0]   int_reg_array_18_0_imag;
  reg        [15:0]   int_reg_array_18_1_real;
  reg        [15:0]   int_reg_array_18_1_imag;
  reg        [15:0]   int_reg_array_18_2_real;
  reg        [15:0]   int_reg_array_18_2_imag;
  reg        [15:0]   int_reg_array_18_3_real;
  reg        [15:0]   int_reg_array_18_3_imag;
  reg        [15:0]   int_reg_array_18_4_real;
  reg        [15:0]   int_reg_array_18_4_imag;
  reg        [15:0]   int_reg_array_18_5_real;
  reg        [15:0]   int_reg_array_18_5_imag;
  reg        [15:0]   int_reg_array_18_6_real;
  reg        [15:0]   int_reg_array_18_6_imag;
  reg        [15:0]   int_reg_array_18_7_real;
  reg        [15:0]   int_reg_array_18_7_imag;
  reg        [15:0]   int_reg_array_18_8_real;
  reg        [15:0]   int_reg_array_18_8_imag;
  reg        [15:0]   int_reg_array_18_9_real;
  reg        [15:0]   int_reg_array_18_9_imag;
  reg        [15:0]   int_reg_array_18_10_real;
  reg        [15:0]   int_reg_array_18_10_imag;
  reg        [15:0]   int_reg_array_18_11_real;
  reg        [15:0]   int_reg_array_18_11_imag;
  reg        [15:0]   int_reg_array_18_12_real;
  reg        [15:0]   int_reg_array_18_12_imag;
  reg        [15:0]   int_reg_array_18_13_real;
  reg        [15:0]   int_reg_array_18_13_imag;
  reg        [15:0]   int_reg_array_18_14_real;
  reg        [15:0]   int_reg_array_18_14_imag;
  reg        [15:0]   int_reg_array_18_15_real;
  reg        [15:0]   int_reg_array_18_15_imag;
  reg        [15:0]   int_reg_array_18_16_real;
  reg        [15:0]   int_reg_array_18_16_imag;
  reg        [15:0]   int_reg_array_18_17_real;
  reg        [15:0]   int_reg_array_18_17_imag;
  reg        [15:0]   int_reg_array_18_18_real;
  reg        [15:0]   int_reg_array_18_18_imag;
  reg        [15:0]   int_reg_array_18_19_real;
  reg        [15:0]   int_reg_array_18_19_imag;
  reg        [15:0]   int_reg_array_18_20_real;
  reg        [15:0]   int_reg_array_18_20_imag;
  reg        [15:0]   int_reg_array_18_21_real;
  reg        [15:0]   int_reg_array_18_21_imag;
  reg        [15:0]   int_reg_array_18_22_real;
  reg        [15:0]   int_reg_array_18_22_imag;
  reg        [15:0]   int_reg_array_18_23_real;
  reg        [15:0]   int_reg_array_18_23_imag;
  reg        [15:0]   int_reg_array_18_24_real;
  reg        [15:0]   int_reg_array_18_24_imag;
  reg        [15:0]   int_reg_array_18_25_real;
  reg        [15:0]   int_reg_array_18_25_imag;
  reg        [15:0]   int_reg_array_18_26_real;
  reg        [15:0]   int_reg_array_18_26_imag;
  reg        [15:0]   int_reg_array_18_27_real;
  reg        [15:0]   int_reg_array_18_27_imag;
  reg        [15:0]   int_reg_array_18_28_real;
  reg        [15:0]   int_reg_array_18_28_imag;
  reg        [15:0]   int_reg_array_18_29_real;
  reg        [15:0]   int_reg_array_18_29_imag;
  reg        [15:0]   int_reg_array_18_30_real;
  reg        [15:0]   int_reg_array_18_30_imag;
  reg        [15:0]   int_reg_array_18_31_real;
  reg        [15:0]   int_reg_array_18_31_imag;
  reg        [15:0]   int_reg_array_18_32_real;
  reg        [15:0]   int_reg_array_18_32_imag;
  reg        [15:0]   int_reg_array_18_33_real;
  reg        [15:0]   int_reg_array_18_33_imag;
  reg        [15:0]   int_reg_array_18_34_real;
  reg        [15:0]   int_reg_array_18_34_imag;
  reg        [15:0]   int_reg_array_18_35_real;
  reg        [15:0]   int_reg_array_18_35_imag;
  reg        [15:0]   int_reg_array_18_36_real;
  reg        [15:0]   int_reg_array_18_36_imag;
  reg        [15:0]   int_reg_array_18_37_real;
  reg        [15:0]   int_reg_array_18_37_imag;
  reg        [15:0]   int_reg_array_18_38_real;
  reg        [15:0]   int_reg_array_18_38_imag;
  reg        [15:0]   int_reg_array_18_39_real;
  reg        [15:0]   int_reg_array_18_39_imag;
  reg        [15:0]   int_reg_array_18_40_real;
  reg        [15:0]   int_reg_array_18_40_imag;
  reg        [15:0]   int_reg_array_18_41_real;
  reg        [15:0]   int_reg_array_18_41_imag;
  reg        [15:0]   int_reg_array_18_42_real;
  reg        [15:0]   int_reg_array_18_42_imag;
  reg        [15:0]   int_reg_array_18_43_real;
  reg        [15:0]   int_reg_array_18_43_imag;
  reg        [15:0]   int_reg_array_18_44_real;
  reg        [15:0]   int_reg_array_18_44_imag;
  reg        [15:0]   int_reg_array_18_45_real;
  reg        [15:0]   int_reg_array_18_45_imag;
  reg        [15:0]   int_reg_array_18_46_real;
  reg        [15:0]   int_reg_array_18_46_imag;
  reg        [15:0]   int_reg_array_18_47_real;
  reg        [15:0]   int_reg_array_18_47_imag;
  reg        [15:0]   int_reg_array_18_48_real;
  reg        [15:0]   int_reg_array_18_48_imag;
  reg        [15:0]   int_reg_array_18_49_real;
  reg        [15:0]   int_reg_array_18_49_imag;
  reg        [15:0]   int_reg_array_34_0_real;
  reg        [15:0]   int_reg_array_34_0_imag;
  reg        [15:0]   int_reg_array_34_1_real;
  reg        [15:0]   int_reg_array_34_1_imag;
  reg        [15:0]   int_reg_array_34_2_real;
  reg        [15:0]   int_reg_array_34_2_imag;
  reg        [15:0]   int_reg_array_34_3_real;
  reg        [15:0]   int_reg_array_34_3_imag;
  reg        [15:0]   int_reg_array_34_4_real;
  reg        [15:0]   int_reg_array_34_4_imag;
  reg        [15:0]   int_reg_array_34_5_real;
  reg        [15:0]   int_reg_array_34_5_imag;
  reg        [15:0]   int_reg_array_34_6_real;
  reg        [15:0]   int_reg_array_34_6_imag;
  reg        [15:0]   int_reg_array_34_7_real;
  reg        [15:0]   int_reg_array_34_7_imag;
  reg        [15:0]   int_reg_array_34_8_real;
  reg        [15:0]   int_reg_array_34_8_imag;
  reg        [15:0]   int_reg_array_34_9_real;
  reg        [15:0]   int_reg_array_34_9_imag;
  reg        [15:0]   int_reg_array_34_10_real;
  reg        [15:0]   int_reg_array_34_10_imag;
  reg        [15:0]   int_reg_array_34_11_real;
  reg        [15:0]   int_reg_array_34_11_imag;
  reg        [15:0]   int_reg_array_34_12_real;
  reg        [15:0]   int_reg_array_34_12_imag;
  reg        [15:0]   int_reg_array_34_13_real;
  reg        [15:0]   int_reg_array_34_13_imag;
  reg        [15:0]   int_reg_array_34_14_real;
  reg        [15:0]   int_reg_array_34_14_imag;
  reg        [15:0]   int_reg_array_34_15_real;
  reg        [15:0]   int_reg_array_34_15_imag;
  reg        [15:0]   int_reg_array_34_16_real;
  reg        [15:0]   int_reg_array_34_16_imag;
  reg        [15:0]   int_reg_array_34_17_real;
  reg        [15:0]   int_reg_array_34_17_imag;
  reg        [15:0]   int_reg_array_34_18_real;
  reg        [15:0]   int_reg_array_34_18_imag;
  reg        [15:0]   int_reg_array_34_19_real;
  reg        [15:0]   int_reg_array_34_19_imag;
  reg        [15:0]   int_reg_array_34_20_real;
  reg        [15:0]   int_reg_array_34_20_imag;
  reg        [15:0]   int_reg_array_34_21_real;
  reg        [15:0]   int_reg_array_34_21_imag;
  reg        [15:0]   int_reg_array_34_22_real;
  reg        [15:0]   int_reg_array_34_22_imag;
  reg        [15:0]   int_reg_array_34_23_real;
  reg        [15:0]   int_reg_array_34_23_imag;
  reg        [15:0]   int_reg_array_34_24_real;
  reg        [15:0]   int_reg_array_34_24_imag;
  reg        [15:0]   int_reg_array_34_25_real;
  reg        [15:0]   int_reg_array_34_25_imag;
  reg        [15:0]   int_reg_array_34_26_real;
  reg        [15:0]   int_reg_array_34_26_imag;
  reg        [15:0]   int_reg_array_34_27_real;
  reg        [15:0]   int_reg_array_34_27_imag;
  reg        [15:0]   int_reg_array_34_28_real;
  reg        [15:0]   int_reg_array_34_28_imag;
  reg        [15:0]   int_reg_array_34_29_real;
  reg        [15:0]   int_reg_array_34_29_imag;
  reg        [15:0]   int_reg_array_34_30_real;
  reg        [15:0]   int_reg_array_34_30_imag;
  reg        [15:0]   int_reg_array_34_31_real;
  reg        [15:0]   int_reg_array_34_31_imag;
  reg        [15:0]   int_reg_array_34_32_real;
  reg        [15:0]   int_reg_array_34_32_imag;
  reg        [15:0]   int_reg_array_34_33_real;
  reg        [15:0]   int_reg_array_34_33_imag;
  reg        [15:0]   int_reg_array_34_34_real;
  reg        [15:0]   int_reg_array_34_34_imag;
  reg        [15:0]   int_reg_array_34_35_real;
  reg        [15:0]   int_reg_array_34_35_imag;
  reg        [15:0]   int_reg_array_34_36_real;
  reg        [15:0]   int_reg_array_34_36_imag;
  reg        [15:0]   int_reg_array_34_37_real;
  reg        [15:0]   int_reg_array_34_37_imag;
  reg        [15:0]   int_reg_array_34_38_real;
  reg        [15:0]   int_reg_array_34_38_imag;
  reg        [15:0]   int_reg_array_34_39_real;
  reg        [15:0]   int_reg_array_34_39_imag;
  reg        [15:0]   int_reg_array_34_40_real;
  reg        [15:0]   int_reg_array_34_40_imag;
  reg        [15:0]   int_reg_array_34_41_real;
  reg        [15:0]   int_reg_array_34_41_imag;
  reg        [15:0]   int_reg_array_34_42_real;
  reg        [15:0]   int_reg_array_34_42_imag;
  reg        [15:0]   int_reg_array_34_43_real;
  reg        [15:0]   int_reg_array_34_43_imag;
  reg        [15:0]   int_reg_array_34_44_real;
  reg        [15:0]   int_reg_array_34_44_imag;
  reg        [15:0]   int_reg_array_34_45_real;
  reg        [15:0]   int_reg_array_34_45_imag;
  reg        [15:0]   int_reg_array_34_46_real;
  reg        [15:0]   int_reg_array_34_46_imag;
  reg        [15:0]   int_reg_array_34_47_real;
  reg        [15:0]   int_reg_array_34_47_imag;
  reg        [15:0]   int_reg_array_34_48_real;
  reg        [15:0]   int_reg_array_34_48_imag;
  reg        [15:0]   int_reg_array_34_49_real;
  reg        [15:0]   int_reg_array_34_49_imag;
  reg        [15:0]   int_reg_array_23_0_real;
  reg        [15:0]   int_reg_array_23_0_imag;
  reg        [15:0]   int_reg_array_23_1_real;
  reg        [15:0]   int_reg_array_23_1_imag;
  reg        [15:0]   int_reg_array_23_2_real;
  reg        [15:0]   int_reg_array_23_2_imag;
  reg        [15:0]   int_reg_array_23_3_real;
  reg        [15:0]   int_reg_array_23_3_imag;
  reg        [15:0]   int_reg_array_23_4_real;
  reg        [15:0]   int_reg_array_23_4_imag;
  reg        [15:0]   int_reg_array_23_5_real;
  reg        [15:0]   int_reg_array_23_5_imag;
  reg        [15:0]   int_reg_array_23_6_real;
  reg        [15:0]   int_reg_array_23_6_imag;
  reg        [15:0]   int_reg_array_23_7_real;
  reg        [15:0]   int_reg_array_23_7_imag;
  reg        [15:0]   int_reg_array_23_8_real;
  reg        [15:0]   int_reg_array_23_8_imag;
  reg        [15:0]   int_reg_array_23_9_real;
  reg        [15:0]   int_reg_array_23_9_imag;
  reg        [15:0]   int_reg_array_23_10_real;
  reg        [15:0]   int_reg_array_23_10_imag;
  reg        [15:0]   int_reg_array_23_11_real;
  reg        [15:0]   int_reg_array_23_11_imag;
  reg        [15:0]   int_reg_array_23_12_real;
  reg        [15:0]   int_reg_array_23_12_imag;
  reg        [15:0]   int_reg_array_23_13_real;
  reg        [15:0]   int_reg_array_23_13_imag;
  reg        [15:0]   int_reg_array_23_14_real;
  reg        [15:0]   int_reg_array_23_14_imag;
  reg        [15:0]   int_reg_array_23_15_real;
  reg        [15:0]   int_reg_array_23_15_imag;
  reg        [15:0]   int_reg_array_23_16_real;
  reg        [15:0]   int_reg_array_23_16_imag;
  reg        [15:0]   int_reg_array_23_17_real;
  reg        [15:0]   int_reg_array_23_17_imag;
  reg        [15:0]   int_reg_array_23_18_real;
  reg        [15:0]   int_reg_array_23_18_imag;
  reg        [15:0]   int_reg_array_23_19_real;
  reg        [15:0]   int_reg_array_23_19_imag;
  reg        [15:0]   int_reg_array_23_20_real;
  reg        [15:0]   int_reg_array_23_20_imag;
  reg        [15:0]   int_reg_array_23_21_real;
  reg        [15:0]   int_reg_array_23_21_imag;
  reg        [15:0]   int_reg_array_23_22_real;
  reg        [15:0]   int_reg_array_23_22_imag;
  reg        [15:0]   int_reg_array_23_23_real;
  reg        [15:0]   int_reg_array_23_23_imag;
  reg        [15:0]   int_reg_array_23_24_real;
  reg        [15:0]   int_reg_array_23_24_imag;
  reg        [15:0]   int_reg_array_23_25_real;
  reg        [15:0]   int_reg_array_23_25_imag;
  reg        [15:0]   int_reg_array_23_26_real;
  reg        [15:0]   int_reg_array_23_26_imag;
  reg        [15:0]   int_reg_array_23_27_real;
  reg        [15:0]   int_reg_array_23_27_imag;
  reg        [15:0]   int_reg_array_23_28_real;
  reg        [15:0]   int_reg_array_23_28_imag;
  reg        [15:0]   int_reg_array_23_29_real;
  reg        [15:0]   int_reg_array_23_29_imag;
  reg        [15:0]   int_reg_array_23_30_real;
  reg        [15:0]   int_reg_array_23_30_imag;
  reg        [15:0]   int_reg_array_23_31_real;
  reg        [15:0]   int_reg_array_23_31_imag;
  reg        [15:0]   int_reg_array_23_32_real;
  reg        [15:0]   int_reg_array_23_32_imag;
  reg        [15:0]   int_reg_array_23_33_real;
  reg        [15:0]   int_reg_array_23_33_imag;
  reg        [15:0]   int_reg_array_23_34_real;
  reg        [15:0]   int_reg_array_23_34_imag;
  reg        [15:0]   int_reg_array_23_35_real;
  reg        [15:0]   int_reg_array_23_35_imag;
  reg        [15:0]   int_reg_array_23_36_real;
  reg        [15:0]   int_reg_array_23_36_imag;
  reg        [15:0]   int_reg_array_23_37_real;
  reg        [15:0]   int_reg_array_23_37_imag;
  reg        [15:0]   int_reg_array_23_38_real;
  reg        [15:0]   int_reg_array_23_38_imag;
  reg        [15:0]   int_reg_array_23_39_real;
  reg        [15:0]   int_reg_array_23_39_imag;
  reg        [15:0]   int_reg_array_23_40_real;
  reg        [15:0]   int_reg_array_23_40_imag;
  reg        [15:0]   int_reg_array_23_41_real;
  reg        [15:0]   int_reg_array_23_41_imag;
  reg        [15:0]   int_reg_array_23_42_real;
  reg        [15:0]   int_reg_array_23_42_imag;
  reg        [15:0]   int_reg_array_23_43_real;
  reg        [15:0]   int_reg_array_23_43_imag;
  reg        [15:0]   int_reg_array_23_44_real;
  reg        [15:0]   int_reg_array_23_44_imag;
  reg        [15:0]   int_reg_array_23_45_real;
  reg        [15:0]   int_reg_array_23_45_imag;
  reg        [15:0]   int_reg_array_23_46_real;
  reg        [15:0]   int_reg_array_23_46_imag;
  reg        [15:0]   int_reg_array_23_47_real;
  reg        [15:0]   int_reg_array_23_47_imag;
  reg        [15:0]   int_reg_array_23_48_real;
  reg        [15:0]   int_reg_array_23_48_imag;
  reg        [15:0]   int_reg_array_23_49_real;
  reg        [15:0]   int_reg_array_23_49_imag;
  reg        [15:0]   int_reg_array_16_0_real;
  reg        [15:0]   int_reg_array_16_0_imag;
  reg        [15:0]   int_reg_array_16_1_real;
  reg        [15:0]   int_reg_array_16_1_imag;
  reg        [15:0]   int_reg_array_16_2_real;
  reg        [15:0]   int_reg_array_16_2_imag;
  reg        [15:0]   int_reg_array_16_3_real;
  reg        [15:0]   int_reg_array_16_3_imag;
  reg        [15:0]   int_reg_array_16_4_real;
  reg        [15:0]   int_reg_array_16_4_imag;
  reg        [15:0]   int_reg_array_16_5_real;
  reg        [15:0]   int_reg_array_16_5_imag;
  reg        [15:0]   int_reg_array_16_6_real;
  reg        [15:0]   int_reg_array_16_6_imag;
  reg        [15:0]   int_reg_array_16_7_real;
  reg        [15:0]   int_reg_array_16_7_imag;
  reg        [15:0]   int_reg_array_16_8_real;
  reg        [15:0]   int_reg_array_16_8_imag;
  reg        [15:0]   int_reg_array_16_9_real;
  reg        [15:0]   int_reg_array_16_9_imag;
  reg        [15:0]   int_reg_array_16_10_real;
  reg        [15:0]   int_reg_array_16_10_imag;
  reg        [15:0]   int_reg_array_16_11_real;
  reg        [15:0]   int_reg_array_16_11_imag;
  reg        [15:0]   int_reg_array_16_12_real;
  reg        [15:0]   int_reg_array_16_12_imag;
  reg        [15:0]   int_reg_array_16_13_real;
  reg        [15:0]   int_reg_array_16_13_imag;
  reg        [15:0]   int_reg_array_16_14_real;
  reg        [15:0]   int_reg_array_16_14_imag;
  reg        [15:0]   int_reg_array_16_15_real;
  reg        [15:0]   int_reg_array_16_15_imag;
  reg        [15:0]   int_reg_array_16_16_real;
  reg        [15:0]   int_reg_array_16_16_imag;
  reg        [15:0]   int_reg_array_16_17_real;
  reg        [15:0]   int_reg_array_16_17_imag;
  reg        [15:0]   int_reg_array_16_18_real;
  reg        [15:0]   int_reg_array_16_18_imag;
  reg        [15:0]   int_reg_array_16_19_real;
  reg        [15:0]   int_reg_array_16_19_imag;
  reg        [15:0]   int_reg_array_16_20_real;
  reg        [15:0]   int_reg_array_16_20_imag;
  reg        [15:0]   int_reg_array_16_21_real;
  reg        [15:0]   int_reg_array_16_21_imag;
  reg        [15:0]   int_reg_array_16_22_real;
  reg        [15:0]   int_reg_array_16_22_imag;
  reg        [15:0]   int_reg_array_16_23_real;
  reg        [15:0]   int_reg_array_16_23_imag;
  reg        [15:0]   int_reg_array_16_24_real;
  reg        [15:0]   int_reg_array_16_24_imag;
  reg        [15:0]   int_reg_array_16_25_real;
  reg        [15:0]   int_reg_array_16_25_imag;
  reg        [15:0]   int_reg_array_16_26_real;
  reg        [15:0]   int_reg_array_16_26_imag;
  reg        [15:0]   int_reg_array_16_27_real;
  reg        [15:0]   int_reg_array_16_27_imag;
  reg        [15:0]   int_reg_array_16_28_real;
  reg        [15:0]   int_reg_array_16_28_imag;
  reg        [15:0]   int_reg_array_16_29_real;
  reg        [15:0]   int_reg_array_16_29_imag;
  reg        [15:0]   int_reg_array_16_30_real;
  reg        [15:0]   int_reg_array_16_30_imag;
  reg        [15:0]   int_reg_array_16_31_real;
  reg        [15:0]   int_reg_array_16_31_imag;
  reg        [15:0]   int_reg_array_16_32_real;
  reg        [15:0]   int_reg_array_16_32_imag;
  reg        [15:0]   int_reg_array_16_33_real;
  reg        [15:0]   int_reg_array_16_33_imag;
  reg        [15:0]   int_reg_array_16_34_real;
  reg        [15:0]   int_reg_array_16_34_imag;
  reg        [15:0]   int_reg_array_16_35_real;
  reg        [15:0]   int_reg_array_16_35_imag;
  reg        [15:0]   int_reg_array_16_36_real;
  reg        [15:0]   int_reg_array_16_36_imag;
  reg        [15:0]   int_reg_array_16_37_real;
  reg        [15:0]   int_reg_array_16_37_imag;
  reg        [15:0]   int_reg_array_16_38_real;
  reg        [15:0]   int_reg_array_16_38_imag;
  reg        [15:0]   int_reg_array_16_39_real;
  reg        [15:0]   int_reg_array_16_39_imag;
  reg        [15:0]   int_reg_array_16_40_real;
  reg        [15:0]   int_reg_array_16_40_imag;
  reg        [15:0]   int_reg_array_16_41_real;
  reg        [15:0]   int_reg_array_16_41_imag;
  reg        [15:0]   int_reg_array_16_42_real;
  reg        [15:0]   int_reg_array_16_42_imag;
  reg        [15:0]   int_reg_array_16_43_real;
  reg        [15:0]   int_reg_array_16_43_imag;
  reg        [15:0]   int_reg_array_16_44_real;
  reg        [15:0]   int_reg_array_16_44_imag;
  reg        [15:0]   int_reg_array_16_45_real;
  reg        [15:0]   int_reg_array_16_45_imag;
  reg        [15:0]   int_reg_array_16_46_real;
  reg        [15:0]   int_reg_array_16_46_imag;
  reg        [15:0]   int_reg_array_16_47_real;
  reg        [15:0]   int_reg_array_16_47_imag;
  reg        [15:0]   int_reg_array_16_48_real;
  reg        [15:0]   int_reg_array_16_48_imag;
  reg        [15:0]   int_reg_array_16_49_real;
  reg        [15:0]   int_reg_array_16_49_imag;
  reg        [15:0]   int_reg_array_45_0_real;
  reg        [15:0]   int_reg_array_45_0_imag;
  reg        [15:0]   int_reg_array_45_1_real;
  reg        [15:0]   int_reg_array_45_1_imag;
  reg        [15:0]   int_reg_array_45_2_real;
  reg        [15:0]   int_reg_array_45_2_imag;
  reg        [15:0]   int_reg_array_45_3_real;
  reg        [15:0]   int_reg_array_45_3_imag;
  reg        [15:0]   int_reg_array_45_4_real;
  reg        [15:0]   int_reg_array_45_4_imag;
  reg        [15:0]   int_reg_array_45_5_real;
  reg        [15:0]   int_reg_array_45_5_imag;
  reg        [15:0]   int_reg_array_45_6_real;
  reg        [15:0]   int_reg_array_45_6_imag;
  reg        [15:0]   int_reg_array_45_7_real;
  reg        [15:0]   int_reg_array_45_7_imag;
  reg        [15:0]   int_reg_array_45_8_real;
  reg        [15:0]   int_reg_array_45_8_imag;
  reg        [15:0]   int_reg_array_45_9_real;
  reg        [15:0]   int_reg_array_45_9_imag;
  reg        [15:0]   int_reg_array_45_10_real;
  reg        [15:0]   int_reg_array_45_10_imag;
  reg        [15:0]   int_reg_array_45_11_real;
  reg        [15:0]   int_reg_array_45_11_imag;
  reg        [15:0]   int_reg_array_45_12_real;
  reg        [15:0]   int_reg_array_45_12_imag;
  reg        [15:0]   int_reg_array_45_13_real;
  reg        [15:0]   int_reg_array_45_13_imag;
  reg        [15:0]   int_reg_array_45_14_real;
  reg        [15:0]   int_reg_array_45_14_imag;
  reg        [15:0]   int_reg_array_45_15_real;
  reg        [15:0]   int_reg_array_45_15_imag;
  reg        [15:0]   int_reg_array_45_16_real;
  reg        [15:0]   int_reg_array_45_16_imag;
  reg        [15:0]   int_reg_array_45_17_real;
  reg        [15:0]   int_reg_array_45_17_imag;
  reg        [15:0]   int_reg_array_45_18_real;
  reg        [15:0]   int_reg_array_45_18_imag;
  reg        [15:0]   int_reg_array_45_19_real;
  reg        [15:0]   int_reg_array_45_19_imag;
  reg        [15:0]   int_reg_array_45_20_real;
  reg        [15:0]   int_reg_array_45_20_imag;
  reg        [15:0]   int_reg_array_45_21_real;
  reg        [15:0]   int_reg_array_45_21_imag;
  reg        [15:0]   int_reg_array_45_22_real;
  reg        [15:0]   int_reg_array_45_22_imag;
  reg        [15:0]   int_reg_array_45_23_real;
  reg        [15:0]   int_reg_array_45_23_imag;
  reg        [15:0]   int_reg_array_45_24_real;
  reg        [15:0]   int_reg_array_45_24_imag;
  reg        [15:0]   int_reg_array_45_25_real;
  reg        [15:0]   int_reg_array_45_25_imag;
  reg        [15:0]   int_reg_array_45_26_real;
  reg        [15:0]   int_reg_array_45_26_imag;
  reg        [15:0]   int_reg_array_45_27_real;
  reg        [15:0]   int_reg_array_45_27_imag;
  reg        [15:0]   int_reg_array_45_28_real;
  reg        [15:0]   int_reg_array_45_28_imag;
  reg        [15:0]   int_reg_array_45_29_real;
  reg        [15:0]   int_reg_array_45_29_imag;
  reg        [15:0]   int_reg_array_45_30_real;
  reg        [15:0]   int_reg_array_45_30_imag;
  reg        [15:0]   int_reg_array_45_31_real;
  reg        [15:0]   int_reg_array_45_31_imag;
  reg        [15:0]   int_reg_array_45_32_real;
  reg        [15:0]   int_reg_array_45_32_imag;
  reg        [15:0]   int_reg_array_45_33_real;
  reg        [15:0]   int_reg_array_45_33_imag;
  reg        [15:0]   int_reg_array_45_34_real;
  reg        [15:0]   int_reg_array_45_34_imag;
  reg        [15:0]   int_reg_array_45_35_real;
  reg        [15:0]   int_reg_array_45_35_imag;
  reg        [15:0]   int_reg_array_45_36_real;
  reg        [15:0]   int_reg_array_45_36_imag;
  reg        [15:0]   int_reg_array_45_37_real;
  reg        [15:0]   int_reg_array_45_37_imag;
  reg        [15:0]   int_reg_array_45_38_real;
  reg        [15:0]   int_reg_array_45_38_imag;
  reg        [15:0]   int_reg_array_45_39_real;
  reg        [15:0]   int_reg_array_45_39_imag;
  reg        [15:0]   int_reg_array_45_40_real;
  reg        [15:0]   int_reg_array_45_40_imag;
  reg        [15:0]   int_reg_array_45_41_real;
  reg        [15:0]   int_reg_array_45_41_imag;
  reg        [15:0]   int_reg_array_45_42_real;
  reg        [15:0]   int_reg_array_45_42_imag;
  reg        [15:0]   int_reg_array_45_43_real;
  reg        [15:0]   int_reg_array_45_43_imag;
  reg        [15:0]   int_reg_array_45_44_real;
  reg        [15:0]   int_reg_array_45_44_imag;
  reg        [15:0]   int_reg_array_45_45_real;
  reg        [15:0]   int_reg_array_45_45_imag;
  reg        [15:0]   int_reg_array_45_46_real;
  reg        [15:0]   int_reg_array_45_46_imag;
  reg        [15:0]   int_reg_array_45_47_real;
  reg        [15:0]   int_reg_array_45_47_imag;
  reg        [15:0]   int_reg_array_45_48_real;
  reg        [15:0]   int_reg_array_45_48_imag;
  reg        [15:0]   int_reg_array_45_49_real;
  reg        [15:0]   int_reg_array_45_49_imag;
  reg        [15:0]   int_reg_array_17_0_real;
  reg        [15:0]   int_reg_array_17_0_imag;
  reg        [15:0]   int_reg_array_17_1_real;
  reg        [15:0]   int_reg_array_17_1_imag;
  reg        [15:0]   int_reg_array_17_2_real;
  reg        [15:0]   int_reg_array_17_2_imag;
  reg        [15:0]   int_reg_array_17_3_real;
  reg        [15:0]   int_reg_array_17_3_imag;
  reg        [15:0]   int_reg_array_17_4_real;
  reg        [15:0]   int_reg_array_17_4_imag;
  reg        [15:0]   int_reg_array_17_5_real;
  reg        [15:0]   int_reg_array_17_5_imag;
  reg        [15:0]   int_reg_array_17_6_real;
  reg        [15:0]   int_reg_array_17_6_imag;
  reg        [15:0]   int_reg_array_17_7_real;
  reg        [15:0]   int_reg_array_17_7_imag;
  reg        [15:0]   int_reg_array_17_8_real;
  reg        [15:0]   int_reg_array_17_8_imag;
  reg        [15:0]   int_reg_array_17_9_real;
  reg        [15:0]   int_reg_array_17_9_imag;
  reg        [15:0]   int_reg_array_17_10_real;
  reg        [15:0]   int_reg_array_17_10_imag;
  reg        [15:0]   int_reg_array_17_11_real;
  reg        [15:0]   int_reg_array_17_11_imag;
  reg        [15:0]   int_reg_array_17_12_real;
  reg        [15:0]   int_reg_array_17_12_imag;
  reg        [15:0]   int_reg_array_17_13_real;
  reg        [15:0]   int_reg_array_17_13_imag;
  reg        [15:0]   int_reg_array_17_14_real;
  reg        [15:0]   int_reg_array_17_14_imag;
  reg        [15:0]   int_reg_array_17_15_real;
  reg        [15:0]   int_reg_array_17_15_imag;
  reg        [15:0]   int_reg_array_17_16_real;
  reg        [15:0]   int_reg_array_17_16_imag;
  reg        [15:0]   int_reg_array_17_17_real;
  reg        [15:0]   int_reg_array_17_17_imag;
  reg        [15:0]   int_reg_array_17_18_real;
  reg        [15:0]   int_reg_array_17_18_imag;
  reg        [15:0]   int_reg_array_17_19_real;
  reg        [15:0]   int_reg_array_17_19_imag;
  reg        [15:0]   int_reg_array_17_20_real;
  reg        [15:0]   int_reg_array_17_20_imag;
  reg        [15:0]   int_reg_array_17_21_real;
  reg        [15:0]   int_reg_array_17_21_imag;
  reg        [15:0]   int_reg_array_17_22_real;
  reg        [15:0]   int_reg_array_17_22_imag;
  reg        [15:0]   int_reg_array_17_23_real;
  reg        [15:0]   int_reg_array_17_23_imag;
  reg        [15:0]   int_reg_array_17_24_real;
  reg        [15:0]   int_reg_array_17_24_imag;
  reg        [15:0]   int_reg_array_17_25_real;
  reg        [15:0]   int_reg_array_17_25_imag;
  reg        [15:0]   int_reg_array_17_26_real;
  reg        [15:0]   int_reg_array_17_26_imag;
  reg        [15:0]   int_reg_array_17_27_real;
  reg        [15:0]   int_reg_array_17_27_imag;
  reg        [15:0]   int_reg_array_17_28_real;
  reg        [15:0]   int_reg_array_17_28_imag;
  reg        [15:0]   int_reg_array_17_29_real;
  reg        [15:0]   int_reg_array_17_29_imag;
  reg        [15:0]   int_reg_array_17_30_real;
  reg        [15:0]   int_reg_array_17_30_imag;
  reg        [15:0]   int_reg_array_17_31_real;
  reg        [15:0]   int_reg_array_17_31_imag;
  reg        [15:0]   int_reg_array_17_32_real;
  reg        [15:0]   int_reg_array_17_32_imag;
  reg        [15:0]   int_reg_array_17_33_real;
  reg        [15:0]   int_reg_array_17_33_imag;
  reg        [15:0]   int_reg_array_17_34_real;
  reg        [15:0]   int_reg_array_17_34_imag;
  reg        [15:0]   int_reg_array_17_35_real;
  reg        [15:0]   int_reg_array_17_35_imag;
  reg        [15:0]   int_reg_array_17_36_real;
  reg        [15:0]   int_reg_array_17_36_imag;
  reg        [15:0]   int_reg_array_17_37_real;
  reg        [15:0]   int_reg_array_17_37_imag;
  reg        [15:0]   int_reg_array_17_38_real;
  reg        [15:0]   int_reg_array_17_38_imag;
  reg        [15:0]   int_reg_array_17_39_real;
  reg        [15:0]   int_reg_array_17_39_imag;
  reg        [15:0]   int_reg_array_17_40_real;
  reg        [15:0]   int_reg_array_17_40_imag;
  reg        [15:0]   int_reg_array_17_41_real;
  reg        [15:0]   int_reg_array_17_41_imag;
  reg        [15:0]   int_reg_array_17_42_real;
  reg        [15:0]   int_reg_array_17_42_imag;
  reg        [15:0]   int_reg_array_17_43_real;
  reg        [15:0]   int_reg_array_17_43_imag;
  reg        [15:0]   int_reg_array_17_44_real;
  reg        [15:0]   int_reg_array_17_44_imag;
  reg        [15:0]   int_reg_array_17_45_real;
  reg        [15:0]   int_reg_array_17_45_imag;
  reg        [15:0]   int_reg_array_17_46_real;
  reg        [15:0]   int_reg_array_17_46_imag;
  reg        [15:0]   int_reg_array_17_47_real;
  reg        [15:0]   int_reg_array_17_47_imag;
  reg        [15:0]   int_reg_array_17_48_real;
  reg        [15:0]   int_reg_array_17_48_imag;
  reg        [15:0]   int_reg_array_17_49_real;
  reg        [15:0]   int_reg_array_17_49_imag;
  reg        [15:0]   int_reg_array_4_0_real;
  reg        [15:0]   int_reg_array_4_0_imag;
  reg        [15:0]   int_reg_array_4_1_real;
  reg        [15:0]   int_reg_array_4_1_imag;
  reg        [15:0]   int_reg_array_4_2_real;
  reg        [15:0]   int_reg_array_4_2_imag;
  reg        [15:0]   int_reg_array_4_3_real;
  reg        [15:0]   int_reg_array_4_3_imag;
  reg        [15:0]   int_reg_array_4_4_real;
  reg        [15:0]   int_reg_array_4_4_imag;
  reg        [15:0]   int_reg_array_4_5_real;
  reg        [15:0]   int_reg_array_4_5_imag;
  reg        [15:0]   int_reg_array_4_6_real;
  reg        [15:0]   int_reg_array_4_6_imag;
  reg        [15:0]   int_reg_array_4_7_real;
  reg        [15:0]   int_reg_array_4_7_imag;
  reg        [15:0]   int_reg_array_4_8_real;
  reg        [15:0]   int_reg_array_4_8_imag;
  reg        [15:0]   int_reg_array_4_9_real;
  reg        [15:0]   int_reg_array_4_9_imag;
  reg        [15:0]   int_reg_array_4_10_real;
  reg        [15:0]   int_reg_array_4_10_imag;
  reg        [15:0]   int_reg_array_4_11_real;
  reg        [15:0]   int_reg_array_4_11_imag;
  reg        [15:0]   int_reg_array_4_12_real;
  reg        [15:0]   int_reg_array_4_12_imag;
  reg        [15:0]   int_reg_array_4_13_real;
  reg        [15:0]   int_reg_array_4_13_imag;
  reg        [15:0]   int_reg_array_4_14_real;
  reg        [15:0]   int_reg_array_4_14_imag;
  reg        [15:0]   int_reg_array_4_15_real;
  reg        [15:0]   int_reg_array_4_15_imag;
  reg        [15:0]   int_reg_array_4_16_real;
  reg        [15:0]   int_reg_array_4_16_imag;
  reg        [15:0]   int_reg_array_4_17_real;
  reg        [15:0]   int_reg_array_4_17_imag;
  reg        [15:0]   int_reg_array_4_18_real;
  reg        [15:0]   int_reg_array_4_18_imag;
  reg        [15:0]   int_reg_array_4_19_real;
  reg        [15:0]   int_reg_array_4_19_imag;
  reg        [15:0]   int_reg_array_4_20_real;
  reg        [15:0]   int_reg_array_4_20_imag;
  reg        [15:0]   int_reg_array_4_21_real;
  reg        [15:0]   int_reg_array_4_21_imag;
  reg        [15:0]   int_reg_array_4_22_real;
  reg        [15:0]   int_reg_array_4_22_imag;
  reg        [15:0]   int_reg_array_4_23_real;
  reg        [15:0]   int_reg_array_4_23_imag;
  reg        [15:0]   int_reg_array_4_24_real;
  reg        [15:0]   int_reg_array_4_24_imag;
  reg        [15:0]   int_reg_array_4_25_real;
  reg        [15:0]   int_reg_array_4_25_imag;
  reg        [15:0]   int_reg_array_4_26_real;
  reg        [15:0]   int_reg_array_4_26_imag;
  reg        [15:0]   int_reg_array_4_27_real;
  reg        [15:0]   int_reg_array_4_27_imag;
  reg        [15:0]   int_reg_array_4_28_real;
  reg        [15:0]   int_reg_array_4_28_imag;
  reg        [15:0]   int_reg_array_4_29_real;
  reg        [15:0]   int_reg_array_4_29_imag;
  reg        [15:0]   int_reg_array_4_30_real;
  reg        [15:0]   int_reg_array_4_30_imag;
  reg        [15:0]   int_reg_array_4_31_real;
  reg        [15:0]   int_reg_array_4_31_imag;
  reg        [15:0]   int_reg_array_4_32_real;
  reg        [15:0]   int_reg_array_4_32_imag;
  reg        [15:0]   int_reg_array_4_33_real;
  reg        [15:0]   int_reg_array_4_33_imag;
  reg        [15:0]   int_reg_array_4_34_real;
  reg        [15:0]   int_reg_array_4_34_imag;
  reg        [15:0]   int_reg_array_4_35_real;
  reg        [15:0]   int_reg_array_4_35_imag;
  reg        [15:0]   int_reg_array_4_36_real;
  reg        [15:0]   int_reg_array_4_36_imag;
  reg        [15:0]   int_reg_array_4_37_real;
  reg        [15:0]   int_reg_array_4_37_imag;
  reg        [15:0]   int_reg_array_4_38_real;
  reg        [15:0]   int_reg_array_4_38_imag;
  reg        [15:0]   int_reg_array_4_39_real;
  reg        [15:0]   int_reg_array_4_39_imag;
  reg        [15:0]   int_reg_array_4_40_real;
  reg        [15:0]   int_reg_array_4_40_imag;
  reg        [15:0]   int_reg_array_4_41_real;
  reg        [15:0]   int_reg_array_4_41_imag;
  reg        [15:0]   int_reg_array_4_42_real;
  reg        [15:0]   int_reg_array_4_42_imag;
  reg        [15:0]   int_reg_array_4_43_real;
  reg        [15:0]   int_reg_array_4_43_imag;
  reg        [15:0]   int_reg_array_4_44_real;
  reg        [15:0]   int_reg_array_4_44_imag;
  reg        [15:0]   int_reg_array_4_45_real;
  reg        [15:0]   int_reg_array_4_45_imag;
  reg        [15:0]   int_reg_array_4_46_real;
  reg        [15:0]   int_reg_array_4_46_imag;
  reg        [15:0]   int_reg_array_4_47_real;
  reg        [15:0]   int_reg_array_4_47_imag;
  reg        [15:0]   int_reg_array_4_48_real;
  reg        [15:0]   int_reg_array_4_48_imag;
  reg        [15:0]   int_reg_array_4_49_real;
  reg        [15:0]   int_reg_array_4_49_imag;
  reg        [15:0]   int_reg_array_27_0_real;
  reg        [15:0]   int_reg_array_27_0_imag;
  reg        [15:0]   int_reg_array_27_1_real;
  reg        [15:0]   int_reg_array_27_1_imag;
  reg        [15:0]   int_reg_array_27_2_real;
  reg        [15:0]   int_reg_array_27_2_imag;
  reg        [15:0]   int_reg_array_27_3_real;
  reg        [15:0]   int_reg_array_27_3_imag;
  reg        [15:0]   int_reg_array_27_4_real;
  reg        [15:0]   int_reg_array_27_4_imag;
  reg        [15:0]   int_reg_array_27_5_real;
  reg        [15:0]   int_reg_array_27_5_imag;
  reg        [15:0]   int_reg_array_27_6_real;
  reg        [15:0]   int_reg_array_27_6_imag;
  reg        [15:0]   int_reg_array_27_7_real;
  reg        [15:0]   int_reg_array_27_7_imag;
  reg        [15:0]   int_reg_array_27_8_real;
  reg        [15:0]   int_reg_array_27_8_imag;
  reg        [15:0]   int_reg_array_27_9_real;
  reg        [15:0]   int_reg_array_27_9_imag;
  reg        [15:0]   int_reg_array_27_10_real;
  reg        [15:0]   int_reg_array_27_10_imag;
  reg        [15:0]   int_reg_array_27_11_real;
  reg        [15:0]   int_reg_array_27_11_imag;
  reg        [15:0]   int_reg_array_27_12_real;
  reg        [15:0]   int_reg_array_27_12_imag;
  reg        [15:0]   int_reg_array_27_13_real;
  reg        [15:0]   int_reg_array_27_13_imag;
  reg        [15:0]   int_reg_array_27_14_real;
  reg        [15:0]   int_reg_array_27_14_imag;
  reg        [15:0]   int_reg_array_27_15_real;
  reg        [15:0]   int_reg_array_27_15_imag;
  reg        [15:0]   int_reg_array_27_16_real;
  reg        [15:0]   int_reg_array_27_16_imag;
  reg        [15:0]   int_reg_array_27_17_real;
  reg        [15:0]   int_reg_array_27_17_imag;
  reg        [15:0]   int_reg_array_27_18_real;
  reg        [15:0]   int_reg_array_27_18_imag;
  reg        [15:0]   int_reg_array_27_19_real;
  reg        [15:0]   int_reg_array_27_19_imag;
  reg        [15:0]   int_reg_array_27_20_real;
  reg        [15:0]   int_reg_array_27_20_imag;
  reg        [15:0]   int_reg_array_27_21_real;
  reg        [15:0]   int_reg_array_27_21_imag;
  reg        [15:0]   int_reg_array_27_22_real;
  reg        [15:0]   int_reg_array_27_22_imag;
  reg        [15:0]   int_reg_array_27_23_real;
  reg        [15:0]   int_reg_array_27_23_imag;
  reg        [15:0]   int_reg_array_27_24_real;
  reg        [15:0]   int_reg_array_27_24_imag;
  reg        [15:0]   int_reg_array_27_25_real;
  reg        [15:0]   int_reg_array_27_25_imag;
  reg        [15:0]   int_reg_array_27_26_real;
  reg        [15:0]   int_reg_array_27_26_imag;
  reg        [15:0]   int_reg_array_27_27_real;
  reg        [15:0]   int_reg_array_27_27_imag;
  reg        [15:0]   int_reg_array_27_28_real;
  reg        [15:0]   int_reg_array_27_28_imag;
  reg        [15:0]   int_reg_array_27_29_real;
  reg        [15:0]   int_reg_array_27_29_imag;
  reg        [15:0]   int_reg_array_27_30_real;
  reg        [15:0]   int_reg_array_27_30_imag;
  reg        [15:0]   int_reg_array_27_31_real;
  reg        [15:0]   int_reg_array_27_31_imag;
  reg        [15:0]   int_reg_array_27_32_real;
  reg        [15:0]   int_reg_array_27_32_imag;
  reg        [15:0]   int_reg_array_27_33_real;
  reg        [15:0]   int_reg_array_27_33_imag;
  reg        [15:0]   int_reg_array_27_34_real;
  reg        [15:0]   int_reg_array_27_34_imag;
  reg        [15:0]   int_reg_array_27_35_real;
  reg        [15:0]   int_reg_array_27_35_imag;
  reg        [15:0]   int_reg_array_27_36_real;
  reg        [15:0]   int_reg_array_27_36_imag;
  reg        [15:0]   int_reg_array_27_37_real;
  reg        [15:0]   int_reg_array_27_37_imag;
  reg        [15:0]   int_reg_array_27_38_real;
  reg        [15:0]   int_reg_array_27_38_imag;
  reg        [15:0]   int_reg_array_27_39_real;
  reg        [15:0]   int_reg_array_27_39_imag;
  reg        [15:0]   int_reg_array_27_40_real;
  reg        [15:0]   int_reg_array_27_40_imag;
  reg        [15:0]   int_reg_array_27_41_real;
  reg        [15:0]   int_reg_array_27_41_imag;
  reg        [15:0]   int_reg_array_27_42_real;
  reg        [15:0]   int_reg_array_27_42_imag;
  reg        [15:0]   int_reg_array_27_43_real;
  reg        [15:0]   int_reg_array_27_43_imag;
  reg        [15:0]   int_reg_array_27_44_real;
  reg        [15:0]   int_reg_array_27_44_imag;
  reg        [15:0]   int_reg_array_27_45_real;
  reg        [15:0]   int_reg_array_27_45_imag;
  reg        [15:0]   int_reg_array_27_46_real;
  reg        [15:0]   int_reg_array_27_46_imag;
  reg        [15:0]   int_reg_array_27_47_real;
  reg        [15:0]   int_reg_array_27_47_imag;
  reg        [15:0]   int_reg_array_27_48_real;
  reg        [15:0]   int_reg_array_27_48_imag;
  reg        [15:0]   int_reg_array_27_49_real;
  reg        [15:0]   int_reg_array_27_49_imag;
  reg        [15:0]   int_reg_array_35_0_real;
  reg        [15:0]   int_reg_array_35_0_imag;
  reg        [15:0]   int_reg_array_35_1_real;
  reg        [15:0]   int_reg_array_35_1_imag;
  reg        [15:0]   int_reg_array_35_2_real;
  reg        [15:0]   int_reg_array_35_2_imag;
  reg        [15:0]   int_reg_array_35_3_real;
  reg        [15:0]   int_reg_array_35_3_imag;
  reg        [15:0]   int_reg_array_35_4_real;
  reg        [15:0]   int_reg_array_35_4_imag;
  reg        [15:0]   int_reg_array_35_5_real;
  reg        [15:0]   int_reg_array_35_5_imag;
  reg        [15:0]   int_reg_array_35_6_real;
  reg        [15:0]   int_reg_array_35_6_imag;
  reg        [15:0]   int_reg_array_35_7_real;
  reg        [15:0]   int_reg_array_35_7_imag;
  reg        [15:0]   int_reg_array_35_8_real;
  reg        [15:0]   int_reg_array_35_8_imag;
  reg        [15:0]   int_reg_array_35_9_real;
  reg        [15:0]   int_reg_array_35_9_imag;
  reg        [15:0]   int_reg_array_35_10_real;
  reg        [15:0]   int_reg_array_35_10_imag;
  reg        [15:0]   int_reg_array_35_11_real;
  reg        [15:0]   int_reg_array_35_11_imag;
  reg        [15:0]   int_reg_array_35_12_real;
  reg        [15:0]   int_reg_array_35_12_imag;
  reg        [15:0]   int_reg_array_35_13_real;
  reg        [15:0]   int_reg_array_35_13_imag;
  reg        [15:0]   int_reg_array_35_14_real;
  reg        [15:0]   int_reg_array_35_14_imag;
  reg        [15:0]   int_reg_array_35_15_real;
  reg        [15:0]   int_reg_array_35_15_imag;
  reg        [15:0]   int_reg_array_35_16_real;
  reg        [15:0]   int_reg_array_35_16_imag;
  reg        [15:0]   int_reg_array_35_17_real;
  reg        [15:0]   int_reg_array_35_17_imag;
  reg        [15:0]   int_reg_array_35_18_real;
  reg        [15:0]   int_reg_array_35_18_imag;
  reg        [15:0]   int_reg_array_35_19_real;
  reg        [15:0]   int_reg_array_35_19_imag;
  reg        [15:0]   int_reg_array_35_20_real;
  reg        [15:0]   int_reg_array_35_20_imag;
  reg        [15:0]   int_reg_array_35_21_real;
  reg        [15:0]   int_reg_array_35_21_imag;
  reg        [15:0]   int_reg_array_35_22_real;
  reg        [15:0]   int_reg_array_35_22_imag;
  reg        [15:0]   int_reg_array_35_23_real;
  reg        [15:0]   int_reg_array_35_23_imag;
  reg        [15:0]   int_reg_array_35_24_real;
  reg        [15:0]   int_reg_array_35_24_imag;
  reg        [15:0]   int_reg_array_35_25_real;
  reg        [15:0]   int_reg_array_35_25_imag;
  reg        [15:0]   int_reg_array_35_26_real;
  reg        [15:0]   int_reg_array_35_26_imag;
  reg        [15:0]   int_reg_array_35_27_real;
  reg        [15:0]   int_reg_array_35_27_imag;
  reg        [15:0]   int_reg_array_35_28_real;
  reg        [15:0]   int_reg_array_35_28_imag;
  reg        [15:0]   int_reg_array_35_29_real;
  reg        [15:0]   int_reg_array_35_29_imag;
  reg        [15:0]   int_reg_array_35_30_real;
  reg        [15:0]   int_reg_array_35_30_imag;
  reg        [15:0]   int_reg_array_35_31_real;
  reg        [15:0]   int_reg_array_35_31_imag;
  reg        [15:0]   int_reg_array_35_32_real;
  reg        [15:0]   int_reg_array_35_32_imag;
  reg        [15:0]   int_reg_array_35_33_real;
  reg        [15:0]   int_reg_array_35_33_imag;
  reg        [15:0]   int_reg_array_35_34_real;
  reg        [15:0]   int_reg_array_35_34_imag;
  reg        [15:0]   int_reg_array_35_35_real;
  reg        [15:0]   int_reg_array_35_35_imag;
  reg        [15:0]   int_reg_array_35_36_real;
  reg        [15:0]   int_reg_array_35_36_imag;
  reg        [15:0]   int_reg_array_35_37_real;
  reg        [15:0]   int_reg_array_35_37_imag;
  reg        [15:0]   int_reg_array_35_38_real;
  reg        [15:0]   int_reg_array_35_38_imag;
  reg        [15:0]   int_reg_array_35_39_real;
  reg        [15:0]   int_reg_array_35_39_imag;
  reg        [15:0]   int_reg_array_35_40_real;
  reg        [15:0]   int_reg_array_35_40_imag;
  reg        [15:0]   int_reg_array_35_41_real;
  reg        [15:0]   int_reg_array_35_41_imag;
  reg        [15:0]   int_reg_array_35_42_real;
  reg        [15:0]   int_reg_array_35_42_imag;
  reg        [15:0]   int_reg_array_35_43_real;
  reg        [15:0]   int_reg_array_35_43_imag;
  reg        [15:0]   int_reg_array_35_44_real;
  reg        [15:0]   int_reg_array_35_44_imag;
  reg        [15:0]   int_reg_array_35_45_real;
  reg        [15:0]   int_reg_array_35_45_imag;
  reg        [15:0]   int_reg_array_35_46_real;
  reg        [15:0]   int_reg_array_35_46_imag;
  reg        [15:0]   int_reg_array_35_47_real;
  reg        [15:0]   int_reg_array_35_47_imag;
  reg        [15:0]   int_reg_array_35_48_real;
  reg        [15:0]   int_reg_array_35_48_imag;
  reg        [15:0]   int_reg_array_35_49_real;
  reg        [15:0]   int_reg_array_35_49_imag;
  reg        [15:0]   int_reg_array_44_0_real;
  reg        [15:0]   int_reg_array_44_0_imag;
  reg        [15:0]   int_reg_array_44_1_real;
  reg        [15:0]   int_reg_array_44_1_imag;
  reg        [15:0]   int_reg_array_44_2_real;
  reg        [15:0]   int_reg_array_44_2_imag;
  reg        [15:0]   int_reg_array_44_3_real;
  reg        [15:0]   int_reg_array_44_3_imag;
  reg        [15:0]   int_reg_array_44_4_real;
  reg        [15:0]   int_reg_array_44_4_imag;
  reg        [15:0]   int_reg_array_44_5_real;
  reg        [15:0]   int_reg_array_44_5_imag;
  reg        [15:0]   int_reg_array_44_6_real;
  reg        [15:0]   int_reg_array_44_6_imag;
  reg        [15:0]   int_reg_array_44_7_real;
  reg        [15:0]   int_reg_array_44_7_imag;
  reg        [15:0]   int_reg_array_44_8_real;
  reg        [15:0]   int_reg_array_44_8_imag;
  reg        [15:0]   int_reg_array_44_9_real;
  reg        [15:0]   int_reg_array_44_9_imag;
  reg        [15:0]   int_reg_array_44_10_real;
  reg        [15:0]   int_reg_array_44_10_imag;
  reg        [15:0]   int_reg_array_44_11_real;
  reg        [15:0]   int_reg_array_44_11_imag;
  reg        [15:0]   int_reg_array_44_12_real;
  reg        [15:0]   int_reg_array_44_12_imag;
  reg        [15:0]   int_reg_array_44_13_real;
  reg        [15:0]   int_reg_array_44_13_imag;
  reg        [15:0]   int_reg_array_44_14_real;
  reg        [15:0]   int_reg_array_44_14_imag;
  reg        [15:0]   int_reg_array_44_15_real;
  reg        [15:0]   int_reg_array_44_15_imag;
  reg        [15:0]   int_reg_array_44_16_real;
  reg        [15:0]   int_reg_array_44_16_imag;
  reg        [15:0]   int_reg_array_44_17_real;
  reg        [15:0]   int_reg_array_44_17_imag;
  reg        [15:0]   int_reg_array_44_18_real;
  reg        [15:0]   int_reg_array_44_18_imag;
  reg        [15:0]   int_reg_array_44_19_real;
  reg        [15:0]   int_reg_array_44_19_imag;
  reg        [15:0]   int_reg_array_44_20_real;
  reg        [15:0]   int_reg_array_44_20_imag;
  reg        [15:0]   int_reg_array_44_21_real;
  reg        [15:0]   int_reg_array_44_21_imag;
  reg        [15:0]   int_reg_array_44_22_real;
  reg        [15:0]   int_reg_array_44_22_imag;
  reg        [15:0]   int_reg_array_44_23_real;
  reg        [15:0]   int_reg_array_44_23_imag;
  reg        [15:0]   int_reg_array_44_24_real;
  reg        [15:0]   int_reg_array_44_24_imag;
  reg        [15:0]   int_reg_array_44_25_real;
  reg        [15:0]   int_reg_array_44_25_imag;
  reg        [15:0]   int_reg_array_44_26_real;
  reg        [15:0]   int_reg_array_44_26_imag;
  reg        [15:0]   int_reg_array_44_27_real;
  reg        [15:0]   int_reg_array_44_27_imag;
  reg        [15:0]   int_reg_array_44_28_real;
  reg        [15:0]   int_reg_array_44_28_imag;
  reg        [15:0]   int_reg_array_44_29_real;
  reg        [15:0]   int_reg_array_44_29_imag;
  reg        [15:0]   int_reg_array_44_30_real;
  reg        [15:0]   int_reg_array_44_30_imag;
  reg        [15:0]   int_reg_array_44_31_real;
  reg        [15:0]   int_reg_array_44_31_imag;
  reg        [15:0]   int_reg_array_44_32_real;
  reg        [15:0]   int_reg_array_44_32_imag;
  reg        [15:0]   int_reg_array_44_33_real;
  reg        [15:0]   int_reg_array_44_33_imag;
  reg        [15:0]   int_reg_array_44_34_real;
  reg        [15:0]   int_reg_array_44_34_imag;
  reg        [15:0]   int_reg_array_44_35_real;
  reg        [15:0]   int_reg_array_44_35_imag;
  reg        [15:0]   int_reg_array_44_36_real;
  reg        [15:0]   int_reg_array_44_36_imag;
  reg        [15:0]   int_reg_array_44_37_real;
  reg        [15:0]   int_reg_array_44_37_imag;
  reg        [15:0]   int_reg_array_44_38_real;
  reg        [15:0]   int_reg_array_44_38_imag;
  reg        [15:0]   int_reg_array_44_39_real;
  reg        [15:0]   int_reg_array_44_39_imag;
  reg        [15:0]   int_reg_array_44_40_real;
  reg        [15:0]   int_reg_array_44_40_imag;
  reg        [15:0]   int_reg_array_44_41_real;
  reg        [15:0]   int_reg_array_44_41_imag;
  reg        [15:0]   int_reg_array_44_42_real;
  reg        [15:0]   int_reg_array_44_42_imag;
  reg        [15:0]   int_reg_array_44_43_real;
  reg        [15:0]   int_reg_array_44_43_imag;
  reg        [15:0]   int_reg_array_44_44_real;
  reg        [15:0]   int_reg_array_44_44_imag;
  reg        [15:0]   int_reg_array_44_45_real;
  reg        [15:0]   int_reg_array_44_45_imag;
  reg        [15:0]   int_reg_array_44_46_real;
  reg        [15:0]   int_reg_array_44_46_imag;
  reg        [15:0]   int_reg_array_44_47_real;
  reg        [15:0]   int_reg_array_44_47_imag;
  reg        [15:0]   int_reg_array_44_48_real;
  reg        [15:0]   int_reg_array_44_48_imag;
  reg        [15:0]   int_reg_array_44_49_real;
  reg        [15:0]   int_reg_array_44_49_imag;
  reg        [15:0]   int_reg_array_9_0_real;
  reg        [15:0]   int_reg_array_9_0_imag;
  reg        [15:0]   int_reg_array_9_1_real;
  reg        [15:0]   int_reg_array_9_1_imag;
  reg        [15:0]   int_reg_array_9_2_real;
  reg        [15:0]   int_reg_array_9_2_imag;
  reg        [15:0]   int_reg_array_9_3_real;
  reg        [15:0]   int_reg_array_9_3_imag;
  reg        [15:0]   int_reg_array_9_4_real;
  reg        [15:0]   int_reg_array_9_4_imag;
  reg        [15:0]   int_reg_array_9_5_real;
  reg        [15:0]   int_reg_array_9_5_imag;
  reg        [15:0]   int_reg_array_9_6_real;
  reg        [15:0]   int_reg_array_9_6_imag;
  reg        [15:0]   int_reg_array_9_7_real;
  reg        [15:0]   int_reg_array_9_7_imag;
  reg        [15:0]   int_reg_array_9_8_real;
  reg        [15:0]   int_reg_array_9_8_imag;
  reg        [15:0]   int_reg_array_9_9_real;
  reg        [15:0]   int_reg_array_9_9_imag;
  reg        [15:0]   int_reg_array_9_10_real;
  reg        [15:0]   int_reg_array_9_10_imag;
  reg        [15:0]   int_reg_array_9_11_real;
  reg        [15:0]   int_reg_array_9_11_imag;
  reg        [15:0]   int_reg_array_9_12_real;
  reg        [15:0]   int_reg_array_9_12_imag;
  reg        [15:0]   int_reg_array_9_13_real;
  reg        [15:0]   int_reg_array_9_13_imag;
  reg        [15:0]   int_reg_array_9_14_real;
  reg        [15:0]   int_reg_array_9_14_imag;
  reg        [15:0]   int_reg_array_9_15_real;
  reg        [15:0]   int_reg_array_9_15_imag;
  reg        [15:0]   int_reg_array_9_16_real;
  reg        [15:0]   int_reg_array_9_16_imag;
  reg        [15:0]   int_reg_array_9_17_real;
  reg        [15:0]   int_reg_array_9_17_imag;
  reg        [15:0]   int_reg_array_9_18_real;
  reg        [15:0]   int_reg_array_9_18_imag;
  reg        [15:0]   int_reg_array_9_19_real;
  reg        [15:0]   int_reg_array_9_19_imag;
  reg        [15:0]   int_reg_array_9_20_real;
  reg        [15:0]   int_reg_array_9_20_imag;
  reg        [15:0]   int_reg_array_9_21_real;
  reg        [15:0]   int_reg_array_9_21_imag;
  reg        [15:0]   int_reg_array_9_22_real;
  reg        [15:0]   int_reg_array_9_22_imag;
  reg        [15:0]   int_reg_array_9_23_real;
  reg        [15:0]   int_reg_array_9_23_imag;
  reg        [15:0]   int_reg_array_9_24_real;
  reg        [15:0]   int_reg_array_9_24_imag;
  reg        [15:0]   int_reg_array_9_25_real;
  reg        [15:0]   int_reg_array_9_25_imag;
  reg        [15:0]   int_reg_array_9_26_real;
  reg        [15:0]   int_reg_array_9_26_imag;
  reg        [15:0]   int_reg_array_9_27_real;
  reg        [15:0]   int_reg_array_9_27_imag;
  reg        [15:0]   int_reg_array_9_28_real;
  reg        [15:0]   int_reg_array_9_28_imag;
  reg        [15:0]   int_reg_array_9_29_real;
  reg        [15:0]   int_reg_array_9_29_imag;
  reg        [15:0]   int_reg_array_9_30_real;
  reg        [15:0]   int_reg_array_9_30_imag;
  reg        [15:0]   int_reg_array_9_31_real;
  reg        [15:0]   int_reg_array_9_31_imag;
  reg        [15:0]   int_reg_array_9_32_real;
  reg        [15:0]   int_reg_array_9_32_imag;
  reg        [15:0]   int_reg_array_9_33_real;
  reg        [15:0]   int_reg_array_9_33_imag;
  reg        [15:0]   int_reg_array_9_34_real;
  reg        [15:0]   int_reg_array_9_34_imag;
  reg        [15:0]   int_reg_array_9_35_real;
  reg        [15:0]   int_reg_array_9_35_imag;
  reg        [15:0]   int_reg_array_9_36_real;
  reg        [15:0]   int_reg_array_9_36_imag;
  reg        [15:0]   int_reg_array_9_37_real;
  reg        [15:0]   int_reg_array_9_37_imag;
  reg        [15:0]   int_reg_array_9_38_real;
  reg        [15:0]   int_reg_array_9_38_imag;
  reg        [15:0]   int_reg_array_9_39_real;
  reg        [15:0]   int_reg_array_9_39_imag;
  reg        [15:0]   int_reg_array_9_40_real;
  reg        [15:0]   int_reg_array_9_40_imag;
  reg        [15:0]   int_reg_array_9_41_real;
  reg        [15:0]   int_reg_array_9_41_imag;
  reg        [15:0]   int_reg_array_9_42_real;
  reg        [15:0]   int_reg_array_9_42_imag;
  reg        [15:0]   int_reg_array_9_43_real;
  reg        [15:0]   int_reg_array_9_43_imag;
  reg        [15:0]   int_reg_array_9_44_real;
  reg        [15:0]   int_reg_array_9_44_imag;
  reg        [15:0]   int_reg_array_9_45_real;
  reg        [15:0]   int_reg_array_9_45_imag;
  reg        [15:0]   int_reg_array_9_46_real;
  reg        [15:0]   int_reg_array_9_46_imag;
  reg        [15:0]   int_reg_array_9_47_real;
  reg        [15:0]   int_reg_array_9_47_imag;
  reg        [15:0]   int_reg_array_9_48_real;
  reg        [15:0]   int_reg_array_9_48_imag;
  reg        [15:0]   int_reg_array_9_49_real;
  reg        [15:0]   int_reg_array_9_49_imag;
  reg        [15:0]   int_reg_array_25_0_real;
  reg        [15:0]   int_reg_array_25_0_imag;
  reg        [15:0]   int_reg_array_25_1_real;
  reg        [15:0]   int_reg_array_25_1_imag;
  reg        [15:0]   int_reg_array_25_2_real;
  reg        [15:0]   int_reg_array_25_2_imag;
  reg        [15:0]   int_reg_array_25_3_real;
  reg        [15:0]   int_reg_array_25_3_imag;
  reg        [15:0]   int_reg_array_25_4_real;
  reg        [15:0]   int_reg_array_25_4_imag;
  reg        [15:0]   int_reg_array_25_5_real;
  reg        [15:0]   int_reg_array_25_5_imag;
  reg        [15:0]   int_reg_array_25_6_real;
  reg        [15:0]   int_reg_array_25_6_imag;
  reg        [15:0]   int_reg_array_25_7_real;
  reg        [15:0]   int_reg_array_25_7_imag;
  reg        [15:0]   int_reg_array_25_8_real;
  reg        [15:0]   int_reg_array_25_8_imag;
  reg        [15:0]   int_reg_array_25_9_real;
  reg        [15:0]   int_reg_array_25_9_imag;
  reg        [15:0]   int_reg_array_25_10_real;
  reg        [15:0]   int_reg_array_25_10_imag;
  reg        [15:0]   int_reg_array_25_11_real;
  reg        [15:0]   int_reg_array_25_11_imag;
  reg        [15:0]   int_reg_array_25_12_real;
  reg        [15:0]   int_reg_array_25_12_imag;
  reg        [15:0]   int_reg_array_25_13_real;
  reg        [15:0]   int_reg_array_25_13_imag;
  reg        [15:0]   int_reg_array_25_14_real;
  reg        [15:0]   int_reg_array_25_14_imag;
  reg        [15:0]   int_reg_array_25_15_real;
  reg        [15:0]   int_reg_array_25_15_imag;
  reg        [15:0]   int_reg_array_25_16_real;
  reg        [15:0]   int_reg_array_25_16_imag;
  reg        [15:0]   int_reg_array_25_17_real;
  reg        [15:0]   int_reg_array_25_17_imag;
  reg        [15:0]   int_reg_array_25_18_real;
  reg        [15:0]   int_reg_array_25_18_imag;
  reg        [15:0]   int_reg_array_25_19_real;
  reg        [15:0]   int_reg_array_25_19_imag;
  reg        [15:0]   int_reg_array_25_20_real;
  reg        [15:0]   int_reg_array_25_20_imag;
  reg        [15:0]   int_reg_array_25_21_real;
  reg        [15:0]   int_reg_array_25_21_imag;
  reg        [15:0]   int_reg_array_25_22_real;
  reg        [15:0]   int_reg_array_25_22_imag;
  reg        [15:0]   int_reg_array_25_23_real;
  reg        [15:0]   int_reg_array_25_23_imag;
  reg        [15:0]   int_reg_array_25_24_real;
  reg        [15:0]   int_reg_array_25_24_imag;
  reg        [15:0]   int_reg_array_25_25_real;
  reg        [15:0]   int_reg_array_25_25_imag;
  reg        [15:0]   int_reg_array_25_26_real;
  reg        [15:0]   int_reg_array_25_26_imag;
  reg        [15:0]   int_reg_array_25_27_real;
  reg        [15:0]   int_reg_array_25_27_imag;
  reg        [15:0]   int_reg_array_25_28_real;
  reg        [15:0]   int_reg_array_25_28_imag;
  reg        [15:0]   int_reg_array_25_29_real;
  reg        [15:0]   int_reg_array_25_29_imag;
  reg        [15:0]   int_reg_array_25_30_real;
  reg        [15:0]   int_reg_array_25_30_imag;
  reg        [15:0]   int_reg_array_25_31_real;
  reg        [15:0]   int_reg_array_25_31_imag;
  reg        [15:0]   int_reg_array_25_32_real;
  reg        [15:0]   int_reg_array_25_32_imag;
  reg        [15:0]   int_reg_array_25_33_real;
  reg        [15:0]   int_reg_array_25_33_imag;
  reg        [15:0]   int_reg_array_25_34_real;
  reg        [15:0]   int_reg_array_25_34_imag;
  reg        [15:0]   int_reg_array_25_35_real;
  reg        [15:0]   int_reg_array_25_35_imag;
  reg        [15:0]   int_reg_array_25_36_real;
  reg        [15:0]   int_reg_array_25_36_imag;
  reg        [15:0]   int_reg_array_25_37_real;
  reg        [15:0]   int_reg_array_25_37_imag;
  reg        [15:0]   int_reg_array_25_38_real;
  reg        [15:0]   int_reg_array_25_38_imag;
  reg        [15:0]   int_reg_array_25_39_real;
  reg        [15:0]   int_reg_array_25_39_imag;
  reg        [15:0]   int_reg_array_25_40_real;
  reg        [15:0]   int_reg_array_25_40_imag;
  reg        [15:0]   int_reg_array_25_41_real;
  reg        [15:0]   int_reg_array_25_41_imag;
  reg        [15:0]   int_reg_array_25_42_real;
  reg        [15:0]   int_reg_array_25_42_imag;
  reg        [15:0]   int_reg_array_25_43_real;
  reg        [15:0]   int_reg_array_25_43_imag;
  reg        [15:0]   int_reg_array_25_44_real;
  reg        [15:0]   int_reg_array_25_44_imag;
  reg        [15:0]   int_reg_array_25_45_real;
  reg        [15:0]   int_reg_array_25_45_imag;
  reg        [15:0]   int_reg_array_25_46_real;
  reg        [15:0]   int_reg_array_25_46_imag;
  reg        [15:0]   int_reg_array_25_47_real;
  reg        [15:0]   int_reg_array_25_47_imag;
  reg        [15:0]   int_reg_array_25_48_real;
  reg        [15:0]   int_reg_array_25_48_imag;
  reg        [15:0]   int_reg_array_25_49_real;
  reg        [15:0]   int_reg_array_25_49_imag;
  reg        [15:0]   int_reg_array_48_0_real;
  reg        [15:0]   int_reg_array_48_0_imag;
  reg        [15:0]   int_reg_array_48_1_real;
  reg        [15:0]   int_reg_array_48_1_imag;
  reg        [15:0]   int_reg_array_48_2_real;
  reg        [15:0]   int_reg_array_48_2_imag;
  reg        [15:0]   int_reg_array_48_3_real;
  reg        [15:0]   int_reg_array_48_3_imag;
  reg        [15:0]   int_reg_array_48_4_real;
  reg        [15:0]   int_reg_array_48_4_imag;
  reg        [15:0]   int_reg_array_48_5_real;
  reg        [15:0]   int_reg_array_48_5_imag;
  reg        [15:0]   int_reg_array_48_6_real;
  reg        [15:0]   int_reg_array_48_6_imag;
  reg        [15:0]   int_reg_array_48_7_real;
  reg        [15:0]   int_reg_array_48_7_imag;
  reg        [15:0]   int_reg_array_48_8_real;
  reg        [15:0]   int_reg_array_48_8_imag;
  reg        [15:0]   int_reg_array_48_9_real;
  reg        [15:0]   int_reg_array_48_9_imag;
  reg        [15:0]   int_reg_array_48_10_real;
  reg        [15:0]   int_reg_array_48_10_imag;
  reg        [15:0]   int_reg_array_48_11_real;
  reg        [15:0]   int_reg_array_48_11_imag;
  reg        [15:0]   int_reg_array_48_12_real;
  reg        [15:0]   int_reg_array_48_12_imag;
  reg        [15:0]   int_reg_array_48_13_real;
  reg        [15:0]   int_reg_array_48_13_imag;
  reg        [15:0]   int_reg_array_48_14_real;
  reg        [15:0]   int_reg_array_48_14_imag;
  reg        [15:0]   int_reg_array_48_15_real;
  reg        [15:0]   int_reg_array_48_15_imag;
  reg        [15:0]   int_reg_array_48_16_real;
  reg        [15:0]   int_reg_array_48_16_imag;
  reg        [15:0]   int_reg_array_48_17_real;
  reg        [15:0]   int_reg_array_48_17_imag;
  reg        [15:0]   int_reg_array_48_18_real;
  reg        [15:0]   int_reg_array_48_18_imag;
  reg        [15:0]   int_reg_array_48_19_real;
  reg        [15:0]   int_reg_array_48_19_imag;
  reg        [15:0]   int_reg_array_48_20_real;
  reg        [15:0]   int_reg_array_48_20_imag;
  reg        [15:0]   int_reg_array_48_21_real;
  reg        [15:0]   int_reg_array_48_21_imag;
  reg        [15:0]   int_reg_array_48_22_real;
  reg        [15:0]   int_reg_array_48_22_imag;
  reg        [15:0]   int_reg_array_48_23_real;
  reg        [15:0]   int_reg_array_48_23_imag;
  reg        [15:0]   int_reg_array_48_24_real;
  reg        [15:0]   int_reg_array_48_24_imag;
  reg        [15:0]   int_reg_array_48_25_real;
  reg        [15:0]   int_reg_array_48_25_imag;
  reg        [15:0]   int_reg_array_48_26_real;
  reg        [15:0]   int_reg_array_48_26_imag;
  reg        [15:0]   int_reg_array_48_27_real;
  reg        [15:0]   int_reg_array_48_27_imag;
  reg        [15:0]   int_reg_array_48_28_real;
  reg        [15:0]   int_reg_array_48_28_imag;
  reg        [15:0]   int_reg_array_48_29_real;
  reg        [15:0]   int_reg_array_48_29_imag;
  reg        [15:0]   int_reg_array_48_30_real;
  reg        [15:0]   int_reg_array_48_30_imag;
  reg        [15:0]   int_reg_array_48_31_real;
  reg        [15:0]   int_reg_array_48_31_imag;
  reg        [15:0]   int_reg_array_48_32_real;
  reg        [15:0]   int_reg_array_48_32_imag;
  reg        [15:0]   int_reg_array_48_33_real;
  reg        [15:0]   int_reg_array_48_33_imag;
  reg        [15:0]   int_reg_array_48_34_real;
  reg        [15:0]   int_reg_array_48_34_imag;
  reg        [15:0]   int_reg_array_48_35_real;
  reg        [15:0]   int_reg_array_48_35_imag;
  reg        [15:0]   int_reg_array_48_36_real;
  reg        [15:0]   int_reg_array_48_36_imag;
  reg        [15:0]   int_reg_array_48_37_real;
  reg        [15:0]   int_reg_array_48_37_imag;
  reg        [15:0]   int_reg_array_48_38_real;
  reg        [15:0]   int_reg_array_48_38_imag;
  reg        [15:0]   int_reg_array_48_39_real;
  reg        [15:0]   int_reg_array_48_39_imag;
  reg        [15:0]   int_reg_array_48_40_real;
  reg        [15:0]   int_reg_array_48_40_imag;
  reg        [15:0]   int_reg_array_48_41_real;
  reg        [15:0]   int_reg_array_48_41_imag;
  reg        [15:0]   int_reg_array_48_42_real;
  reg        [15:0]   int_reg_array_48_42_imag;
  reg        [15:0]   int_reg_array_48_43_real;
  reg        [15:0]   int_reg_array_48_43_imag;
  reg        [15:0]   int_reg_array_48_44_real;
  reg        [15:0]   int_reg_array_48_44_imag;
  reg        [15:0]   int_reg_array_48_45_real;
  reg        [15:0]   int_reg_array_48_45_imag;
  reg        [15:0]   int_reg_array_48_46_real;
  reg        [15:0]   int_reg_array_48_46_imag;
  reg        [15:0]   int_reg_array_48_47_real;
  reg        [15:0]   int_reg_array_48_47_imag;
  reg        [15:0]   int_reg_array_48_48_real;
  reg        [15:0]   int_reg_array_48_48_imag;
  reg        [15:0]   int_reg_array_48_49_real;
  reg        [15:0]   int_reg_array_48_49_imag;
  reg        [15:0]   int_reg_array_47_0_real;
  reg        [15:0]   int_reg_array_47_0_imag;
  reg        [15:0]   int_reg_array_47_1_real;
  reg        [15:0]   int_reg_array_47_1_imag;
  reg        [15:0]   int_reg_array_47_2_real;
  reg        [15:0]   int_reg_array_47_2_imag;
  reg        [15:0]   int_reg_array_47_3_real;
  reg        [15:0]   int_reg_array_47_3_imag;
  reg        [15:0]   int_reg_array_47_4_real;
  reg        [15:0]   int_reg_array_47_4_imag;
  reg        [15:0]   int_reg_array_47_5_real;
  reg        [15:0]   int_reg_array_47_5_imag;
  reg        [15:0]   int_reg_array_47_6_real;
  reg        [15:0]   int_reg_array_47_6_imag;
  reg        [15:0]   int_reg_array_47_7_real;
  reg        [15:0]   int_reg_array_47_7_imag;
  reg        [15:0]   int_reg_array_47_8_real;
  reg        [15:0]   int_reg_array_47_8_imag;
  reg        [15:0]   int_reg_array_47_9_real;
  reg        [15:0]   int_reg_array_47_9_imag;
  reg        [15:0]   int_reg_array_47_10_real;
  reg        [15:0]   int_reg_array_47_10_imag;
  reg        [15:0]   int_reg_array_47_11_real;
  reg        [15:0]   int_reg_array_47_11_imag;
  reg        [15:0]   int_reg_array_47_12_real;
  reg        [15:0]   int_reg_array_47_12_imag;
  reg        [15:0]   int_reg_array_47_13_real;
  reg        [15:0]   int_reg_array_47_13_imag;
  reg        [15:0]   int_reg_array_47_14_real;
  reg        [15:0]   int_reg_array_47_14_imag;
  reg        [15:0]   int_reg_array_47_15_real;
  reg        [15:0]   int_reg_array_47_15_imag;
  reg        [15:0]   int_reg_array_47_16_real;
  reg        [15:0]   int_reg_array_47_16_imag;
  reg        [15:0]   int_reg_array_47_17_real;
  reg        [15:0]   int_reg_array_47_17_imag;
  reg        [15:0]   int_reg_array_47_18_real;
  reg        [15:0]   int_reg_array_47_18_imag;
  reg        [15:0]   int_reg_array_47_19_real;
  reg        [15:0]   int_reg_array_47_19_imag;
  reg        [15:0]   int_reg_array_47_20_real;
  reg        [15:0]   int_reg_array_47_20_imag;
  reg        [15:0]   int_reg_array_47_21_real;
  reg        [15:0]   int_reg_array_47_21_imag;
  reg        [15:0]   int_reg_array_47_22_real;
  reg        [15:0]   int_reg_array_47_22_imag;
  reg        [15:0]   int_reg_array_47_23_real;
  reg        [15:0]   int_reg_array_47_23_imag;
  reg        [15:0]   int_reg_array_47_24_real;
  reg        [15:0]   int_reg_array_47_24_imag;
  reg        [15:0]   int_reg_array_47_25_real;
  reg        [15:0]   int_reg_array_47_25_imag;
  reg        [15:0]   int_reg_array_47_26_real;
  reg        [15:0]   int_reg_array_47_26_imag;
  reg        [15:0]   int_reg_array_47_27_real;
  reg        [15:0]   int_reg_array_47_27_imag;
  reg        [15:0]   int_reg_array_47_28_real;
  reg        [15:0]   int_reg_array_47_28_imag;
  reg        [15:0]   int_reg_array_47_29_real;
  reg        [15:0]   int_reg_array_47_29_imag;
  reg        [15:0]   int_reg_array_47_30_real;
  reg        [15:0]   int_reg_array_47_30_imag;
  reg        [15:0]   int_reg_array_47_31_real;
  reg        [15:0]   int_reg_array_47_31_imag;
  reg        [15:0]   int_reg_array_47_32_real;
  reg        [15:0]   int_reg_array_47_32_imag;
  reg        [15:0]   int_reg_array_47_33_real;
  reg        [15:0]   int_reg_array_47_33_imag;
  reg        [15:0]   int_reg_array_47_34_real;
  reg        [15:0]   int_reg_array_47_34_imag;
  reg        [15:0]   int_reg_array_47_35_real;
  reg        [15:0]   int_reg_array_47_35_imag;
  reg        [15:0]   int_reg_array_47_36_real;
  reg        [15:0]   int_reg_array_47_36_imag;
  reg        [15:0]   int_reg_array_47_37_real;
  reg        [15:0]   int_reg_array_47_37_imag;
  reg        [15:0]   int_reg_array_47_38_real;
  reg        [15:0]   int_reg_array_47_38_imag;
  reg        [15:0]   int_reg_array_47_39_real;
  reg        [15:0]   int_reg_array_47_39_imag;
  reg        [15:0]   int_reg_array_47_40_real;
  reg        [15:0]   int_reg_array_47_40_imag;
  reg        [15:0]   int_reg_array_47_41_real;
  reg        [15:0]   int_reg_array_47_41_imag;
  reg        [15:0]   int_reg_array_47_42_real;
  reg        [15:0]   int_reg_array_47_42_imag;
  reg        [15:0]   int_reg_array_47_43_real;
  reg        [15:0]   int_reg_array_47_43_imag;
  reg        [15:0]   int_reg_array_47_44_real;
  reg        [15:0]   int_reg_array_47_44_imag;
  reg        [15:0]   int_reg_array_47_45_real;
  reg        [15:0]   int_reg_array_47_45_imag;
  reg        [15:0]   int_reg_array_47_46_real;
  reg        [15:0]   int_reg_array_47_46_imag;
  reg        [15:0]   int_reg_array_47_47_real;
  reg        [15:0]   int_reg_array_47_47_imag;
  reg        [15:0]   int_reg_array_47_48_real;
  reg        [15:0]   int_reg_array_47_48_imag;
  reg        [15:0]   int_reg_array_47_49_real;
  reg        [15:0]   int_reg_array_47_49_imag;
  reg        [15:0]   int_reg_array_24_0_real;
  reg        [15:0]   int_reg_array_24_0_imag;
  reg        [15:0]   int_reg_array_24_1_real;
  reg        [15:0]   int_reg_array_24_1_imag;
  reg        [15:0]   int_reg_array_24_2_real;
  reg        [15:0]   int_reg_array_24_2_imag;
  reg        [15:0]   int_reg_array_24_3_real;
  reg        [15:0]   int_reg_array_24_3_imag;
  reg        [15:0]   int_reg_array_24_4_real;
  reg        [15:0]   int_reg_array_24_4_imag;
  reg        [15:0]   int_reg_array_24_5_real;
  reg        [15:0]   int_reg_array_24_5_imag;
  reg        [15:0]   int_reg_array_24_6_real;
  reg        [15:0]   int_reg_array_24_6_imag;
  reg        [15:0]   int_reg_array_24_7_real;
  reg        [15:0]   int_reg_array_24_7_imag;
  reg        [15:0]   int_reg_array_24_8_real;
  reg        [15:0]   int_reg_array_24_8_imag;
  reg        [15:0]   int_reg_array_24_9_real;
  reg        [15:0]   int_reg_array_24_9_imag;
  reg        [15:0]   int_reg_array_24_10_real;
  reg        [15:0]   int_reg_array_24_10_imag;
  reg        [15:0]   int_reg_array_24_11_real;
  reg        [15:0]   int_reg_array_24_11_imag;
  reg        [15:0]   int_reg_array_24_12_real;
  reg        [15:0]   int_reg_array_24_12_imag;
  reg        [15:0]   int_reg_array_24_13_real;
  reg        [15:0]   int_reg_array_24_13_imag;
  reg        [15:0]   int_reg_array_24_14_real;
  reg        [15:0]   int_reg_array_24_14_imag;
  reg        [15:0]   int_reg_array_24_15_real;
  reg        [15:0]   int_reg_array_24_15_imag;
  reg        [15:0]   int_reg_array_24_16_real;
  reg        [15:0]   int_reg_array_24_16_imag;
  reg        [15:0]   int_reg_array_24_17_real;
  reg        [15:0]   int_reg_array_24_17_imag;
  reg        [15:0]   int_reg_array_24_18_real;
  reg        [15:0]   int_reg_array_24_18_imag;
  reg        [15:0]   int_reg_array_24_19_real;
  reg        [15:0]   int_reg_array_24_19_imag;
  reg        [15:0]   int_reg_array_24_20_real;
  reg        [15:0]   int_reg_array_24_20_imag;
  reg        [15:0]   int_reg_array_24_21_real;
  reg        [15:0]   int_reg_array_24_21_imag;
  reg        [15:0]   int_reg_array_24_22_real;
  reg        [15:0]   int_reg_array_24_22_imag;
  reg        [15:0]   int_reg_array_24_23_real;
  reg        [15:0]   int_reg_array_24_23_imag;
  reg        [15:0]   int_reg_array_24_24_real;
  reg        [15:0]   int_reg_array_24_24_imag;
  reg        [15:0]   int_reg_array_24_25_real;
  reg        [15:0]   int_reg_array_24_25_imag;
  reg        [15:0]   int_reg_array_24_26_real;
  reg        [15:0]   int_reg_array_24_26_imag;
  reg        [15:0]   int_reg_array_24_27_real;
  reg        [15:0]   int_reg_array_24_27_imag;
  reg        [15:0]   int_reg_array_24_28_real;
  reg        [15:0]   int_reg_array_24_28_imag;
  reg        [15:0]   int_reg_array_24_29_real;
  reg        [15:0]   int_reg_array_24_29_imag;
  reg        [15:0]   int_reg_array_24_30_real;
  reg        [15:0]   int_reg_array_24_30_imag;
  reg        [15:0]   int_reg_array_24_31_real;
  reg        [15:0]   int_reg_array_24_31_imag;
  reg        [15:0]   int_reg_array_24_32_real;
  reg        [15:0]   int_reg_array_24_32_imag;
  reg        [15:0]   int_reg_array_24_33_real;
  reg        [15:0]   int_reg_array_24_33_imag;
  reg        [15:0]   int_reg_array_24_34_real;
  reg        [15:0]   int_reg_array_24_34_imag;
  reg        [15:0]   int_reg_array_24_35_real;
  reg        [15:0]   int_reg_array_24_35_imag;
  reg        [15:0]   int_reg_array_24_36_real;
  reg        [15:0]   int_reg_array_24_36_imag;
  reg        [15:0]   int_reg_array_24_37_real;
  reg        [15:0]   int_reg_array_24_37_imag;
  reg        [15:0]   int_reg_array_24_38_real;
  reg        [15:0]   int_reg_array_24_38_imag;
  reg        [15:0]   int_reg_array_24_39_real;
  reg        [15:0]   int_reg_array_24_39_imag;
  reg        [15:0]   int_reg_array_24_40_real;
  reg        [15:0]   int_reg_array_24_40_imag;
  reg        [15:0]   int_reg_array_24_41_real;
  reg        [15:0]   int_reg_array_24_41_imag;
  reg        [15:0]   int_reg_array_24_42_real;
  reg        [15:0]   int_reg_array_24_42_imag;
  reg        [15:0]   int_reg_array_24_43_real;
  reg        [15:0]   int_reg_array_24_43_imag;
  reg        [15:0]   int_reg_array_24_44_real;
  reg        [15:0]   int_reg_array_24_44_imag;
  reg        [15:0]   int_reg_array_24_45_real;
  reg        [15:0]   int_reg_array_24_45_imag;
  reg        [15:0]   int_reg_array_24_46_real;
  reg        [15:0]   int_reg_array_24_46_imag;
  reg        [15:0]   int_reg_array_24_47_real;
  reg        [15:0]   int_reg_array_24_47_imag;
  reg        [15:0]   int_reg_array_24_48_real;
  reg        [15:0]   int_reg_array_24_48_imag;
  reg        [15:0]   int_reg_array_24_49_real;
  reg        [15:0]   int_reg_array_24_49_imag;
  reg        [15:0]   int_reg_array_15_0_real;
  reg        [15:0]   int_reg_array_15_0_imag;
  reg        [15:0]   int_reg_array_15_1_real;
  reg        [15:0]   int_reg_array_15_1_imag;
  reg        [15:0]   int_reg_array_15_2_real;
  reg        [15:0]   int_reg_array_15_2_imag;
  reg        [15:0]   int_reg_array_15_3_real;
  reg        [15:0]   int_reg_array_15_3_imag;
  reg        [15:0]   int_reg_array_15_4_real;
  reg        [15:0]   int_reg_array_15_4_imag;
  reg        [15:0]   int_reg_array_15_5_real;
  reg        [15:0]   int_reg_array_15_5_imag;
  reg        [15:0]   int_reg_array_15_6_real;
  reg        [15:0]   int_reg_array_15_6_imag;
  reg        [15:0]   int_reg_array_15_7_real;
  reg        [15:0]   int_reg_array_15_7_imag;
  reg        [15:0]   int_reg_array_15_8_real;
  reg        [15:0]   int_reg_array_15_8_imag;
  reg        [15:0]   int_reg_array_15_9_real;
  reg        [15:0]   int_reg_array_15_9_imag;
  reg        [15:0]   int_reg_array_15_10_real;
  reg        [15:0]   int_reg_array_15_10_imag;
  reg        [15:0]   int_reg_array_15_11_real;
  reg        [15:0]   int_reg_array_15_11_imag;
  reg        [15:0]   int_reg_array_15_12_real;
  reg        [15:0]   int_reg_array_15_12_imag;
  reg        [15:0]   int_reg_array_15_13_real;
  reg        [15:0]   int_reg_array_15_13_imag;
  reg        [15:0]   int_reg_array_15_14_real;
  reg        [15:0]   int_reg_array_15_14_imag;
  reg        [15:0]   int_reg_array_15_15_real;
  reg        [15:0]   int_reg_array_15_15_imag;
  reg        [15:0]   int_reg_array_15_16_real;
  reg        [15:0]   int_reg_array_15_16_imag;
  reg        [15:0]   int_reg_array_15_17_real;
  reg        [15:0]   int_reg_array_15_17_imag;
  reg        [15:0]   int_reg_array_15_18_real;
  reg        [15:0]   int_reg_array_15_18_imag;
  reg        [15:0]   int_reg_array_15_19_real;
  reg        [15:0]   int_reg_array_15_19_imag;
  reg        [15:0]   int_reg_array_15_20_real;
  reg        [15:0]   int_reg_array_15_20_imag;
  reg        [15:0]   int_reg_array_15_21_real;
  reg        [15:0]   int_reg_array_15_21_imag;
  reg        [15:0]   int_reg_array_15_22_real;
  reg        [15:0]   int_reg_array_15_22_imag;
  reg        [15:0]   int_reg_array_15_23_real;
  reg        [15:0]   int_reg_array_15_23_imag;
  reg        [15:0]   int_reg_array_15_24_real;
  reg        [15:0]   int_reg_array_15_24_imag;
  reg        [15:0]   int_reg_array_15_25_real;
  reg        [15:0]   int_reg_array_15_25_imag;
  reg        [15:0]   int_reg_array_15_26_real;
  reg        [15:0]   int_reg_array_15_26_imag;
  reg        [15:0]   int_reg_array_15_27_real;
  reg        [15:0]   int_reg_array_15_27_imag;
  reg        [15:0]   int_reg_array_15_28_real;
  reg        [15:0]   int_reg_array_15_28_imag;
  reg        [15:0]   int_reg_array_15_29_real;
  reg        [15:0]   int_reg_array_15_29_imag;
  reg        [15:0]   int_reg_array_15_30_real;
  reg        [15:0]   int_reg_array_15_30_imag;
  reg        [15:0]   int_reg_array_15_31_real;
  reg        [15:0]   int_reg_array_15_31_imag;
  reg        [15:0]   int_reg_array_15_32_real;
  reg        [15:0]   int_reg_array_15_32_imag;
  reg        [15:0]   int_reg_array_15_33_real;
  reg        [15:0]   int_reg_array_15_33_imag;
  reg        [15:0]   int_reg_array_15_34_real;
  reg        [15:0]   int_reg_array_15_34_imag;
  reg        [15:0]   int_reg_array_15_35_real;
  reg        [15:0]   int_reg_array_15_35_imag;
  reg        [15:0]   int_reg_array_15_36_real;
  reg        [15:0]   int_reg_array_15_36_imag;
  reg        [15:0]   int_reg_array_15_37_real;
  reg        [15:0]   int_reg_array_15_37_imag;
  reg        [15:0]   int_reg_array_15_38_real;
  reg        [15:0]   int_reg_array_15_38_imag;
  reg        [15:0]   int_reg_array_15_39_real;
  reg        [15:0]   int_reg_array_15_39_imag;
  reg        [15:0]   int_reg_array_15_40_real;
  reg        [15:0]   int_reg_array_15_40_imag;
  reg        [15:0]   int_reg_array_15_41_real;
  reg        [15:0]   int_reg_array_15_41_imag;
  reg        [15:0]   int_reg_array_15_42_real;
  reg        [15:0]   int_reg_array_15_42_imag;
  reg        [15:0]   int_reg_array_15_43_real;
  reg        [15:0]   int_reg_array_15_43_imag;
  reg        [15:0]   int_reg_array_15_44_real;
  reg        [15:0]   int_reg_array_15_44_imag;
  reg        [15:0]   int_reg_array_15_45_real;
  reg        [15:0]   int_reg_array_15_45_imag;
  reg        [15:0]   int_reg_array_15_46_real;
  reg        [15:0]   int_reg_array_15_46_imag;
  reg        [15:0]   int_reg_array_15_47_real;
  reg        [15:0]   int_reg_array_15_47_imag;
  reg        [15:0]   int_reg_array_15_48_real;
  reg        [15:0]   int_reg_array_15_48_imag;
  reg        [15:0]   int_reg_array_15_49_real;
  reg        [15:0]   int_reg_array_15_49_imag;
  reg        [15:0]   int_reg_array_32_0_real;
  reg        [15:0]   int_reg_array_32_0_imag;
  reg        [15:0]   int_reg_array_32_1_real;
  reg        [15:0]   int_reg_array_32_1_imag;
  reg        [15:0]   int_reg_array_32_2_real;
  reg        [15:0]   int_reg_array_32_2_imag;
  reg        [15:0]   int_reg_array_32_3_real;
  reg        [15:0]   int_reg_array_32_3_imag;
  reg        [15:0]   int_reg_array_32_4_real;
  reg        [15:0]   int_reg_array_32_4_imag;
  reg        [15:0]   int_reg_array_32_5_real;
  reg        [15:0]   int_reg_array_32_5_imag;
  reg        [15:0]   int_reg_array_32_6_real;
  reg        [15:0]   int_reg_array_32_6_imag;
  reg        [15:0]   int_reg_array_32_7_real;
  reg        [15:0]   int_reg_array_32_7_imag;
  reg        [15:0]   int_reg_array_32_8_real;
  reg        [15:0]   int_reg_array_32_8_imag;
  reg        [15:0]   int_reg_array_32_9_real;
  reg        [15:0]   int_reg_array_32_9_imag;
  reg        [15:0]   int_reg_array_32_10_real;
  reg        [15:0]   int_reg_array_32_10_imag;
  reg        [15:0]   int_reg_array_32_11_real;
  reg        [15:0]   int_reg_array_32_11_imag;
  reg        [15:0]   int_reg_array_32_12_real;
  reg        [15:0]   int_reg_array_32_12_imag;
  reg        [15:0]   int_reg_array_32_13_real;
  reg        [15:0]   int_reg_array_32_13_imag;
  reg        [15:0]   int_reg_array_32_14_real;
  reg        [15:0]   int_reg_array_32_14_imag;
  reg        [15:0]   int_reg_array_32_15_real;
  reg        [15:0]   int_reg_array_32_15_imag;
  reg        [15:0]   int_reg_array_32_16_real;
  reg        [15:0]   int_reg_array_32_16_imag;
  reg        [15:0]   int_reg_array_32_17_real;
  reg        [15:0]   int_reg_array_32_17_imag;
  reg        [15:0]   int_reg_array_32_18_real;
  reg        [15:0]   int_reg_array_32_18_imag;
  reg        [15:0]   int_reg_array_32_19_real;
  reg        [15:0]   int_reg_array_32_19_imag;
  reg        [15:0]   int_reg_array_32_20_real;
  reg        [15:0]   int_reg_array_32_20_imag;
  reg        [15:0]   int_reg_array_32_21_real;
  reg        [15:0]   int_reg_array_32_21_imag;
  reg        [15:0]   int_reg_array_32_22_real;
  reg        [15:0]   int_reg_array_32_22_imag;
  reg        [15:0]   int_reg_array_32_23_real;
  reg        [15:0]   int_reg_array_32_23_imag;
  reg        [15:0]   int_reg_array_32_24_real;
  reg        [15:0]   int_reg_array_32_24_imag;
  reg        [15:0]   int_reg_array_32_25_real;
  reg        [15:0]   int_reg_array_32_25_imag;
  reg        [15:0]   int_reg_array_32_26_real;
  reg        [15:0]   int_reg_array_32_26_imag;
  reg        [15:0]   int_reg_array_32_27_real;
  reg        [15:0]   int_reg_array_32_27_imag;
  reg        [15:0]   int_reg_array_32_28_real;
  reg        [15:0]   int_reg_array_32_28_imag;
  reg        [15:0]   int_reg_array_32_29_real;
  reg        [15:0]   int_reg_array_32_29_imag;
  reg        [15:0]   int_reg_array_32_30_real;
  reg        [15:0]   int_reg_array_32_30_imag;
  reg        [15:0]   int_reg_array_32_31_real;
  reg        [15:0]   int_reg_array_32_31_imag;
  reg        [15:0]   int_reg_array_32_32_real;
  reg        [15:0]   int_reg_array_32_32_imag;
  reg        [15:0]   int_reg_array_32_33_real;
  reg        [15:0]   int_reg_array_32_33_imag;
  reg        [15:0]   int_reg_array_32_34_real;
  reg        [15:0]   int_reg_array_32_34_imag;
  reg        [15:0]   int_reg_array_32_35_real;
  reg        [15:0]   int_reg_array_32_35_imag;
  reg        [15:0]   int_reg_array_32_36_real;
  reg        [15:0]   int_reg_array_32_36_imag;
  reg        [15:0]   int_reg_array_32_37_real;
  reg        [15:0]   int_reg_array_32_37_imag;
  reg        [15:0]   int_reg_array_32_38_real;
  reg        [15:0]   int_reg_array_32_38_imag;
  reg        [15:0]   int_reg_array_32_39_real;
  reg        [15:0]   int_reg_array_32_39_imag;
  reg        [15:0]   int_reg_array_32_40_real;
  reg        [15:0]   int_reg_array_32_40_imag;
  reg        [15:0]   int_reg_array_32_41_real;
  reg        [15:0]   int_reg_array_32_41_imag;
  reg        [15:0]   int_reg_array_32_42_real;
  reg        [15:0]   int_reg_array_32_42_imag;
  reg        [15:0]   int_reg_array_32_43_real;
  reg        [15:0]   int_reg_array_32_43_imag;
  reg        [15:0]   int_reg_array_32_44_real;
  reg        [15:0]   int_reg_array_32_44_imag;
  reg        [15:0]   int_reg_array_32_45_real;
  reg        [15:0]   int_reg_array_32_45_imag;
  reg        [15:0]   int_reg_array_32_46_real;
  reg        [15:0]   int_reg_array_32_46_imag;
  reg        [15:0]   int_reg_array_32_47_real;
  reg        [15:0]   int_reg_array_32_47_imag;
  reg        [15:0]   int_reg_array_32_48_real;
  reg        [15:0]   int_reg_array_32_48_imag;
  reg        [15:0]   int_reg_array_32_49_real;
  reg        [15:0]   int_reg_array_32_49_imag;
  reg        [15:0]   int_reg_array_13_0_real;
  reg        [15:0]   int_reg_array_13_0_imag;
  reg        [15:0]   int_reg_array_13_1_real;
  reg        [15:0]   int_reg_array_13_1_imag;
  reg        [15:0]   int_reg_array_13_2_real;
  reg        [15:0]   int_reg_array_13_2_imag;
  reg        [15:0]   int_reg_array_13_3_real;
  reg        [15:0]   int_reg_array_13_3_imag;
  reg        [15:0]   int_reg_array_13_4_real;
  reg        [15:0]   int_reg_array_13_4_imag;
  reg        [15:0]   int_reg_array_13_5_real;
  reg        [15:0]   int_reg_array_13_5_imag;
  reg        [15:0]   int_reg_array_13_6_real;
  reg        [15:0]   int_reg_array_13_6_imag;
  reg        [15:0]   int_reg_array_13_7_real;
  reg        [15:0]   int_reg_array_13_7_imag;
  reg        [15:0]   int_reg_array_13_8_real;
  reg        [15:0]   int_reg_array_13_8_imag;
  reg        [15:0]   int_reg_array_13_9_real;
  reg        [15:0]   int_reg_array_13_9_imag;
  reg        [15:0]   int_reg_array_13_10_real;
  reg        [15:0]   int_reg_array_13_10_imag;
  reg        [15:0]   int_reg_array_13_11_real;
  reg        [15:0]   int_reg_array_13_11_imag;
  reg        [15:0]   int_reg_array_13_12_real;
  reg        [15:0]   int_reg_array_13_12_imag;
  reg        [15:0]   int_reg_array_13_13_real;
  reg        [15:0]   int_reg_array_13_13_imag;
  reg        [15:0]   int_reg_array_13_14_real;
  reg        [15:0]   int_reg_array_13_14_imag;
  reg        [15:0]   int_reg_array_13_15_real;
  reg        [15:0]   int_reg_array_13_15_imag;
  reg        [15:0]   int_reg_array_13_16_real;
  reg        [15:0]   int_reg_array_13_16_imag;
  reg        [15:0]   int_reg_array_13_17_real;
  reg        [15:0]   int_reg_array_13_17_imag;
  reg        [15:0]   int_reg_array_13_18_real;
  reg        [15:0]   int_reg_array_13_18_imag;
  reg        [15:0]   int_reg_array_13_19_real;
  reg        [15:0]   int_reg_array_13_19_imag;
  reg        [15:0]   int_reg_array_13_20_real;
  reg        [15:0]   int_reg_array_13_20_imag;
  reg        [15:0]   int_reg_array_13_21_real;
  reg        [15:0]   int_reg_array_13_21_imag;
  reg        [15:0]   int_reg_array_13_22_real;
  reg        [15:0]   int_reg_array_13_22_imag;
  reg        [15:0]   int_reg_array_13_23_real;
  reg        [15:0]   int_reg_array_13_23_imag;
  reg        [15:0]   int_reg_array_13_24_real;
  reg        [15:0]   int_reg_array_13_24_imag;
  reg        [15:0]   int_reg_array_13_25_real;
  reg        [15:0]   int_reg_array_13_25_imag;
  reg        [15:0]   int_reg_array_13_26_real;
  reg        [15:0]   int_reg_array_13_26_imag;
  reg        [15:0]   int_reg_array_13_27_real;
  reg        [15:0]   int_reg_array_13_27_imag;
  reg        [15:0]   int_reg_array_13_28_real;
  reg        [15:0]   int_reg_array_13_28_imag;
  reg        [15:0]   int_reg_array_13_29_real;
  reg        [15:0]   int_reg_array_13_29_imag;
  reg        [15:0]   int_reg_array_13_30_real;
  reg        [15:0]   int_reg_array_13_30_imag;
  reg        [15:0]   int_reg_array_13_31_real;
  reg        [15:0]   int_reg_array_13_31_imag;
  reg        [15:0]   int_reg_array_13_32_real;
  reg        [15:0]   int_reg_array_13_32_imag;
  reg        [15:0]   int_reg_array_13_33_real;
  reg        [15:0]   int_reg_array_13_33_imag;
  reg        [15:0]   int_reg_array_13_34_real;
  reg        [15:0]   int_reg_array_13_34_imag;
  reg        [15:0]   int_reg_array_13_35_real;
  reg        [15:0]   int_reg_array_13_35_imag;
  reg        [15:0]   int_reg_array_13_36_real;
  reg        [15:0]   int_reg_array_13_36_imag;
  reg        [15:0]   int_reg_array_13_37_real;
  reg        [15:0]   int_reg_array_13_37_imag;
  reg        [15:0]   int_reg_array_13_38_real;
  reg        [15:0]   int_reg_array_13_38_imag;
  reg        [15:0]   int_reg_array_13_39_real;
  reg        [15:0]   int_reg_array_13_39_imag;
  reg        [15:0]   int_reg_array_13_40_real;
  reg        [15:0]   int_reg_array_13_40_imag;
  reg        [15:0]   int_reg_array_13_41_real;
  reg        [15:0]   int_reg_array_13_41_imag;
  reg        [15:0]   int_reg_array_13_42_real;
  reg        [15:0]   int_reg_array_13_42_imag;
  reg        [15:0]   int_reg_array_13_43_real;
  reg        [15:0]   int_reg_array_13_43_imag;
  reg        [15:0]   int_reg_array_13_44_real;
  reg        [15:0]   int_reg_array_13_44_imag;
  reg        [15:0]   int_reg_array_13_45_real;
  reg        [15:0]   int_reg_array_13_45_imag;
  reg        [15:0]   int_reg_array_13_46_real;
  reg        [15:0]   int_reg_array_13_46_imag;
  reg        [15:0]   int_reg_array_13_47_real;
  reg        [15:0]   int_reg_array_13_47_imag;
  reg        [15:0]   int_reg_array_13_48_real;
  reg        [15:0]   int_reg_array_13_48_imag;
  reg        [15:0]   int_reg_array_13_49_real;
  reg        [15:0]   int_reg_array_13_49_imag;
  reg        [15:0]   int_reg_array_12_0_real;
  reg        [15:0]   int_reg_array_12_0_imag;
  reg        [15:0]   int_reg_array_12_1_real;
  reg        [15:0]   int_reg_array_12_1_imag;
  reg        [15:0]   int_reg_array_12_2_real;
  reg        [15:0]   int_reg_array_12_2_imag;
  reg        [15:0]   int_reg_array_12_3_real;
  reg        [15:0]   int_reg_array_12_3_imag;
  reg        [15:0]   int_reg_array_12_4_real;
  reg        [15:0]   int_reg_array_12_4_imag;
  reg        [15:0]   int_reg_array_12_5_real;
  reg        [15:0]   int_reg_array_12_5_imag;
  reg        [15:0]   int_reg_array_12_6_real;
  reg        [15:0]   int_reg_array_12_6_imag;
  reg        [15:0]   int_reg_array_12_7_real;
  reg        [15:0]   int_reg_array_12_7_imag;
  reg        [15:0]   int_reg_array_12_8_real;
  reg        [15:0]   int_reg_array_12_8_imag;
  reg        [15:0]   int_reg_array_12_9_real;
  reg        [15:0]   int_reg_array_12_9_imag;
  reg        [15:0]   int_reg_array_12_10_real;
  reg        [15:0]   int_reg_array_12_10_imag;
  reg        [15:0]   int_reg_array_12_11_real;
  reg        [15:0]   int_reg_array_12_11_imag;
  reg        [15:0]   int_reg_array_12_12_real;
  reg        [15:0]   int_reg_array_12_12_imag;
  reg        [15:0]   int_reg_array_12_13_real;
  reg        [15:0]   int_reg_array_12_13_imag;
  reg        [15:0]   int_reg_array_12_14_real;
  reg        [15:0]   int_reg_array_12_14_imag;
  reg        [15:0]   int_reg_array_12_15_real;
  reg        [15:0]   int_reg_array_12_15_imag;
  reg        [15:0]   int_reg_array_12_16_real;
  reg        [15:0]   int_reg_array_12_16_imag;
  reg        [15:0]   int_reg_array_12_17_real;
  reg        [15:0]   int_reg_array_12_17_imag;
  reg        [15:0]   int_reg_array_12_18_real;
  reg        [15:0]   int_reg_array_12_18_imag;
  reg        [15:0]   int_reg_array_12_19_real;
  reg        [15:0]   int_reg_array_12_19_imag;
  reg        [15:0]   int_reg_array_12_20_real;
  reg        [15:0]   int_reg_array_12_20_imag;
  reg        [15:0]   int_reg_array_12_21_real;
  reg        [15:0]   int_reg_array_12_21_imag;
  reg        [15:0]   int_reg_array_12_22_real;
  reg        [15:0]   int_reg_array_12_22_imag;
  reg        [15:0]   int_reg_array_12_23_real;
  reg        [15:0]   int_reg_array_12_23_imag;
  reg        [15:0]   int_reg_array_12_24_real;
  reg        [15:0]   int_reg_array_12_24_imag;
  reg        [15:0]   int_reg_array_12_25_real;
  reg        [15:0]   int_reg_array_12_25_imag;
  reg        [15:0]   int_reg_array_12_26_real;
  reg        [15:0]   int_reg_array_12_26_imag;
  reg        [15:0]   int_reg_array_12_27_real;
  reg        [15:0]   int_reg_array_12_27_imag;
  reg        [15:0]   int_reg_array_12_28_real;
  reg        [15:0]   int_reg_array_12_28_imag;
  reg        [15:0]   int_reg_array_12_29_real;
  reg        [15:0]   int_reg_array_12_29_imag;
  reg        [15:0]   int_reg_array_12_30_real;
  reg        [15:0]   int_reg_array_12_30_imag;
  reg        [15:0]   int_reg_array_12_31_real;
  reg        [15:0]   int_reg_array_12_31_imag;
  reg        [15:0]   int_reg_array_12_32_real;
  reg        [15:0]   int_reg_array_12_32_imag;
  reg        [15:0]   int_reg_array_12_33_real;
  reg        [15:0]   int_reg_array_12_33_imag;
  reg        [15:0]   int_reg_array_12_34_real;
  reg        [15:0]   int_reg_array_12_34_imag;
  reg        [15:0]   int_reg_array_12_35_real;
  reg        [15:0]   int_reg_array_12_35_imag;
  reg        [15:0]   int_reg_array_12_36_real;
  reg        [15:0]   int_reg_array_12_36_imag;
  reg        [15:0]   int_reg_array_12_37_real;
  reg        [15:0]   int_reg_array_12_37_imag;
  reg        [15:0]   int_reg_array_12_38_real;
  reg        [15:0]   int_reg_array_12_38_imag;
  reg        [15:0]   int_reg_array_12_39_real;
  reg        [15:0]   int_reg_array_12_39_imag;
  reg        [15:0]   int_reg_array_12_40_real;
  reg        [15:0]   int_reg_array_12_40_imag;
  reg        [15:0]   int_reg_array_12_41_real;
  reg        [15:0]   int_reg_array_12_41_imag;
  reg        [15:0]   int_reg_array_12_42_real;
  reg        [15:0]   int_reg_array_12_42_imag;
  reg        [15:0]   int_reg_array_12_43_real;
  reg        [15:0]   int_reg_array_12_43_imag;
  reg        [15:0]   int_reg_array_12_44_real;
  reg        [15:0]   int_reg_array_12_44_imag;
  reg        [15:0]   int_reg_array_12_45_real;
  reg        [15:0]   int_reg_array_12_45_imag;
  reg        [15:0]   int_reg_array_12_46_real;
  reg        [15:0]   int_reg_array_12_46_imag;
  reg        [15:0]   int_reg_array_12_47_real;
  reg        [15:0]   int_reg_array_12_47_imag;
  reg        [15:0]   int_reg_array_12_48_real;
  reg        [15:0]   int_reg_array_12_48_imag;
  reg        [15:0]   int_reg_array_12_49_real;
  reg        [15:0]   int_reg_array_12_49_imag;
  reg        [15:0]   int_reg_array_39_0_real;
  reg        [15:0]   int_reg_array_39_0_imag;
  reg        [15:0]   int_reg_array_39_1_real;
  reg        [15:0]   int_reg_array_39_1_imag;
  reg        [15:0]   int_reg_array_39_2_real;
  reg        [15:0]   int_reg_array_39_2_imag;
  reg        [15:0]   int_reg_array_39_3_real;
  reg        [15:0]   int_reg_array_39_3_imag;
  reg        [15:0]   int_reg_array_39_4_real;
  reg        [15:0]   int_reg_array_39_4_imag;
  reg        [15:0]   int_reg_array_39_5_real;
  reg        [15:0]   int_reg_array_39_5_imag;
  reg        [15:0]   int_reg_array_39_6_real;
  reg        [15:0]   int_reg_array_39_6_imag;
  reg        [15:0]   int_reg_array_39_7_real;
  reg        [15:0]   int_reg_array_39_7_imag;
  reg        [15:0]   int_reg_array_39_8_real;
  reg        [15:0]   int_reg_array_39_8_imag;
  reg        [15:0]   int_reg_array_39_9_real;
  reg        [15:0]   int_reg_array_39_9_imag;
  reg        [15:0]   int_reg_array_39_10_real;
  reg        [15:0]   int_reg_array_39_10_imag;
  reg        [15:0]   int_reg_array_39_11_real;
  reg        [15:0]   int_reg_array_39_11_imag;
  reg        [15:0]   int_reg_array_39_12_real;
  reg        [15:0]   int_reg_array_39_12_imag;
  reg        [15:0]   int_reg_array_39_13_real;
  reg        [15:0]   int_reg_array_39_13_imag;
  reg        [15:0]   int_reg_array_39_14_real;
  reg        [15:0]   int_reg_array_39_14_imag;
  reg        [15:0]   int_reg_array_39_15_real;
  reg        [15:0]   int_reg_array_39_15_imag;
  reg        [15:0]   int_reg_array_39_16_real;
  reg        [15:0]   int_reg_array_39_16_imag;
  reg        [15:0]   int_reg_array_39_17_real;
  reg        [15:0]   int_reg_array_39_17_imag;
  reg        [15:0]   int_reg_array_39_18_real;
  reg        [15:0]   int_reg_array_39_18_imag;
  reg        [15:0]   int_reg_array_39_19_real;
  reg        [15:0]   int_reg_array_39_19_imag;
  reg        [15:0]   int_reg_array_39_20_real;
  reg        [15:0]   int_reg_array_39_20_imag;
  reg        [15:0]   int_reg_array_39_21_real;
  reg        [15:0]   int_reg_array_39_21_imag;
  reg        [15:0]   int_reg_array_39_22_real;
  reg        [15:0]   int_reg_array_39_22_imag;
  reg        [15:0]   int_reg_array_39_23_real;
  reg        [15:0]   int_reg_array_39_23_imag;
  reg        [15:0]   int_reg_array_39_24_real;
  reg        [15:0]   int_reg_array_39_24_imag;
  reg        [15:0]   int_reg_array_39_25_real;
  reg        [15:0]   int_reg_array_39_25_imag;
  reg        [15:0]   int_reg_array_39_26_real;
  reg        [15:0]   int_reg_array_39_26_imag;
  reg        [15:0]   int_reg_array_39_27_real;
  reg        [15:0]   int_reg_array_39_27_imag;
  reg        [15:0]   int_reg_array_39_28_real;
  reg        [15:0]   int_reg_array_39_28_imag;
  reg        [15:0]   int_reg_array_39_29_real;
  reg        [15:0]   int_reg_array_39_29_imag;
  reg        [15:0]   int_reg_array_39_30_real;
  reg        [15:0]   int_reg_array_39_30_imag;
  reg        [15:0]   int_reg_array_39_31_real;
  reg        [15:0]   int_reg_array_39_31_imag;
  reg        [15:0]   int_reg_array_39_32_real;
  reg        [15:0]   int_reg_array_39_32_imag;
  reg        [15:0]   int_reg_array_39_33_real;
  reg        [15:0]   int_reg_array_39_33_imag;
  reg        [15:0]   int_reg_array_39_34_real;
  reg        [15:0]   int_reg_array_39_34_imag;
  reg        [15:0]   int_reg_array_39_35_real;
  reg        [15:0]   int_reg_array_39_35_imag;
  reg        [15:0]   int_reg_array_39_36_real;
  reg        [15:0]   int_reg_array_39_36_imag;
  reg        [15:0]   int_reg_array_39_37_real;
  reg        [15:0]   int_reg_array_39_37_imag;
  reg        [15:0]   int_reg_array_39_38_real;
  reg        [15:0]   int_reg_array_39_38_imag;
  reg        [15:0]   int_reg_array_39_39_real;
  reg        [15:0]   int_reg_array_39_39_imag;
  reg        [15:0]   int_reg_array_39_40_real;
  reg        [15:0]   int_reg_array_39_40_imag;
  reg        [15:0]   int_reg_array_39_41_real;
  reg        [15:0]   int_reg_array_39_41_imag;
  reg        [15:0]   int_reg_array_39_42_real;
  reg        [15:0]   int_reg_array_39_42_imag;
  reg        [15:0]   int_reg_array_39_43_real;
  reg        [15:0]   int_reg_array_39_43_imag;
  reg        [15:0]   int_reg_array_39_44_real;
  reg        [15:0]   int_reg_array_39_44_imag;
  reg        [15:0]   int_reg_array_39_45_real;
  reg        [15:0]   int_reg_array_39_45_imag;
  reg        [15:0]   int_reg_array_39_46_real;
  reg        [15:0]   int_reg_array_39_46_imag;
  reg        [15:0]   int_reg_array_39_47_real;
  reg        [15:0]   int_reg_array_39_47_imag;
  reg        [15:0]   int_reg_array_39_48_real;
  reg        [15:0]   int_reg_array_39_48_imag;
  reg        [15:0]   int_reg_array_39_49_real;
  reg        [15:0]   int_reg_array_39_49_imag;
  reg        [15:0]   int_reg_array_43_0_real;
  reg        [15:0]   int_reg_array_43_0_imag;
  reg        [15:0]   int_reg_array_43_1_real;
  reg        [15:0]   int_reg_array_43_1_imag;
  reg        [15:0]   int_reg_array_43_2_real;
  reg        [15:0]   int_reg_array_43_2_imag;
  reg        [15:0]   int_reg_array_43_3_real;
  reg        [15:0]   int_reg_array_43_3_imag;
  reg        [15:0]   int_reg_array_43_4_real;
  reg        [15:0]   int_reg_array_43_4_imag;
  reg        [15:0]   int_reg_array_43_5_real;
  reg        [15:0]   int_reg_array_43_5_imag;
  reg        [15:0]   int_reg_array_43_6_real;
  reg        [15:0]   int_reg_array_43_6_imag;
  reg        [15:0]   int_reg_array_43_7_real;
  reg        [15:0]   int_reg_array_43_7_imag;
  reg        [15:0]   int_reg_array_43_8_real;
  reg        [15:0]   int_reg_array_43_8_imag;
  reg        [15:0]   int_reg_array_43_9_real;
  reg        [15:0]   int_reg_array_43_9_imag;
  reg        [15:0]   int_reg_array_43_10_real;
  reg        [15:0]   int_reg_array_43_10_imag;
  reg        [15:0]   int_reg_array_43_11_real;
  reg        [15:0]   int_reg_array_43_11_imag;
  reg        [15:0]   int_reg_array_43_12_real;
  reg        [15:0]   int_reg_array_43_12_imag;
  reg        [15:0]   int_reg_array_43_13_real;
  reg        [15:0]   int_reg_array_43_13_imag;
  reg        [15:0]   int_reg_array_43_14_real;
  reg        [15:0]   int_reg_array_43_14_imag;
  reg        [15:0]   int_reg_array_43_15_real;
  reg        [15:0]   int_reg_array_43_15_imag;
  reg        [15:0]   int_reg_array_43_16_real;
  reg        [15:0]   int_reg_array_43_16_imag;
  reg        [15:0]   int_reg_array_43_17_real;
  reg        [15:0]   int_reg_array_43_17_imag;
  reg        [15:0]   int_reg_array_43_18_real;
  reg        [15:0]   int_reg_array_43_18_imag;
  reg        [15:0]   int_reg_array_43_19_real;
  reg        [15:0]   int_reg_array_43_19_imag;
  reg        [15:0]   int_reg_array_43_20_real;
  reg        [15:0]   int_reg_array_43_20_imag;
  reg        [15:0]   int_reg_array_43_21_real;
  reg        [15:0]   int_reg_array_43_21_imag;
  reg        [15:0]   int_reg_array_43_22_real;
  reg        [15:0]   int_reg_array_43_22_imag;
  reg        [15:0]   int_reg_array_43_23_real;
  reg        [15:0]   int_reg_array_43_23_imag;
  reg        [15:0]   int_reg_array_43_24_real;
  reg        [15:0]   int_reg_array_43_24_imag;
  reg        [15:0]   int_reg_array_43_25_real;
  reg        [15:0]   int_reg_array_43_25_imag;
  reg        [15:0]   int_reg_array_43_26_real;
  reg        [15:0]   int_reg_array_43_26_imag;
  reg        [15:0]   int_reg_array_43_27_real;
  reg        [15:0]   int_reg_array_43_27_imag;
  reg        [15:0]   int_reg_array_43_28_real;
  reg        [15:0]   int_reg_array_43_28_imag;
  reg        [15:0]   int_reg_array_43_29_real;
  reg        [15:0]   int_reg_array_43_29_imag;
  reg        [15:0]   int_reg_array_43_30_real;
  reg        [15:0]   int_reg_array_43_30_imag;
  reg        [15:0]   int_reg_array_43_31_real;
  reg        [15:0]   int_reg_array_43_31_imag;
  reg        [15:0]   int_reg_array_43_32_real;
  reg        [15:0]   int_reg_array_43_32_imag;
  reg        [15:0]   int_reg_array_43_33_real;
  reg        [15:0]   int_reg_array_43_33_imag;
  reg        [15:0]   int_reg_array_43_34_real;
  reg        [15:0]   int_reg_array_43_34_imag;
  reg        [15:0]   int_reg_array_43_35_real;
  reg        [15:0]   int_reg_array_43_35_imag;
  reg        [15:0]   int_reg_array_43_36_real;
  reg        [15:0]   int_reg_array_43_36_imag;
  reg        [15:0]   int_reg_array_43_37_real;
  reg        [15:0]   int_reg_array_43_37_imag;
  reg        [15:0]   int_reg_array_43_38_real;
  reg        [15:0]   int_reg_array_43_38_imag;
  reg        [15:0]   int_reg_array_43_39_real;
  reg        [15:0]   int_reg_array_43_39_imag;
  reg        [15:0]   int_reg_array_43_40_real;
  reg        [15:0]   int_reg_array_43_40_imag;
  reg        [15:0]   int_reg_array_43_41_real;
  reg        [15:0]   int_reg_array_43_41_imag;
  reg        [15:0]   int_reg_array_43_42_real;
  reg        [15:0]   int_reg_array_43_42_imag;
  reg        [15:0]   int_reg_array_43_43_real;
  reg        [15:0]   int_reg_array_43_43_imag;
  reg        [15:0]   int_reg_array_43_44_real;
  reg        [15:0]   int_reg_array_43_44_imag;
  reg        [15:0]   int_reg_array_43_45_real;
  reg        [15:0]   int_reg_array_43_45_imag;
  reg        [15:0]   int_reg_array_43_46_real;
  reg        [15:0]   int_reg_array_43_46_imag;
  reg        [15:0]   int_reg_array_43_47_real;
  reg        [15:0]   int_reg_array_43_47_imag;
  reg        [15:0]   int_reg_array_43_48_real;
  reg        [15:0]   int_reg_array_43_48_imag;
  reg        [15:0]   int_reg_array_43_49_real;
  reg        [15:0]   int_reg_array_43_49_imag;
  reg        [15:0]   int_reg_array_33_0_real;
  reg        [15:0]   int_reg_array_33_0_imag;
  reg        [15:0]   int_reg_array_33_1_real;
  reg        [15:0]   int_reg_array_33_1_imag;
  reg        [15:0]   int_reg_array_33_2_real;
  reg        [15:0]   int_reg_array_33_2_imag;
  reg        [15:0]   int_reg_array_33_3_real;
  reg        [15:0]   int_reg_array_33_3_imag;
  reg        [15:0]   int_reg_array_33_4_real;
  reg        [15:0]   int_reg_array_33_4_imag;
  reg        [15:0]   int_reg_array_33_5_real;
  reg        [15:0]   int_reg_array_33_5_imag;
  reg        [15:0]   int_reg_array_33_6_real;
  reg        [15:0]   int_reg_array_33_6_imag;
  reg        [15:0]   int_reg_array_33_7_real;
  reg        [15:0]   int_reg_array_33_7_imag;
  reg        [15:0]   int_reg_array_33_8_real;
  reg        [15:0]   int_reg_array_33_8_imag;
  reg        [15:0]   int_reg_array_33_9_real;
  reg        [15:0]   int_reg_array_33_9_imag;
  reg        [15:0]   int_reg_array_33_10_real;
  reg        [15:0]   int_reg_array_33_10_imag;
  reg        [15:0]   int_reg_array_33_11_real;
  reg        [15:0]   int_reg_array_33_11_imag;
  reg        [15:0]   int_reg_array_33_12_real;
  reg        [15:0]   int_reg_array_33_12_imag;
  reg        [15:0]   int_reg_array_33_13_real;
  reg        [15:0]   int_reg_array_33_13_imag;
  reg        [15:0]   int_reg_array_33_14_real;
  reg        [15:0]   int_reg_array_33_14_imag;
  reg        [15:0]   int_reg_array_33_15_real;
  reg        [15:0]   int_reg_array_33_15_imag;
  reg        [15:0]   int_reg_array_33_16_real;
  reg        [15:0]   int_reg_array_33_16_imag;
  reg        [15:0]   int_reg_array_33_17_real;
  reg        [15:0]   int_reg_array_33_17_imag;
  reg        [15:0]   int_reg_array_33_18_real;
  reg        [15:0]   int_reg_array_33_18_imag;
  reg        [15:0]   int_reg_array_33_19_real;
  reg        [15:0]   int_reg_array_33_19_imag;
  reg        [15:0]   int_reg_array_33_20_real;
  reg        [15:0]   int_reg_array_33_20_imag;
  reg        [15:0]   int_reg_array_33_21_real;
  reg        [15:0]   int_reg_array_33_21_imag;
  reg        [15:0]   int_reg_array_33_22_real;
  reg        [15:0]   int_reg_array_33_22_imag;
  reg        [15:0]   int_reg_array_33_23_real;
  reg        [15:0]   int_reg_array_33_23_imag;
  reg        [15:0]   int_reg_array_33_24_real;
  reg        [15:0]   int_reg_array_33_24_imag;
  reg        [15:0]   int_reg_array_33_25_real;
  reg        [15:0]   int_reg_array_33_25_imag;
  reg        [15:0]   int_reg_array_33_26_real;
  reg        [15:0]   int_reg_array_33_26_imag;
  reg        [15:0]   int_reg_array_33_27_real;
  reg        [15:0]   int_reg_array_33_27_imag;
  reg        [15:0]   int_reg_array_33_28_real;
  reg        [15:0]   int_reg_array_33_28_imag;
  reg        [15:0]   int_reg_array_33_29_real;
  reg        [15:0]   int_reg_array_33_29_imag;
  reg        [15:0]   int_reg_array_33_30_real;
  reg        [15:0]   int_reg_array_33_30_imag;
  reg        [15:0]   int_reg_array_33_31_real;
  reg        [15:0]   int_reg_array_33_31_imag;
  reg        [15:0]   int_reg_array_33_32_real;
  reg        [15:0]   int_reg_array_33_32_imag;
  reg        [15:0]   int_reg_array_33_33_real;
  reg        [15:0]   int_reg_array_33_33_imag;
  reg        [15:0]   int_reg_array_33_34_real;
  reg        [15:0]   int_reg_array_33_34_imag;
  reg        [15:0]   int_reg_array_33_35_real;
  reg        [15:0]   int_reg_array_33_35_imag;
  reg        [15:0]   int_reg_array_33_36_real;
  reg        [15:0]   int_reg_array_33_36_imag;
  reg        [15:0]   int_reg_array_33_37_real;
  reg        [15:0]   int_reg_array_33_37_imag;
  reg        [15:0]   int_reg_array_33_38_real;
  reg        [15:0]   int_reg_array_33_38_imag;
  reg        [15:0]   int_reg_array_33_39_real;
  reg        [15:0]   int_reg_array_33_39_imag;
  reg        [15:0]   int_reg_array_33_40_real;
  reg        [15:0]   int_reg_array_33_40_imag;
  reg        [15:0]   int_reg_array_33_41_real;
  reg        [15:0]   int_reg_array_33_41_imag;
  reg        [15:0]   int_reg_array_33_42_real;
  reg        [15:0]   int_reg_array_33_42_imag;
  reg        [15:0]   int_reg_array_33_43_real;
  reg        [15:0]   int_reg_array_33_43_imag;
  reg        [15:0]   int_reg_array_33_44_real;
  reg        [15:0]   int_reg_array_33_44_imag;
  reg        [15:0]   int_reg_array_33_45_real;
  reg        [15:0]   int_reg_array_33_45_imag;
  reg        [15:0]   int_reg_array_33_46_real;
  reg        [15:0]   int_reg_array_33_46_imag;
  reg        [15:0]   int_reg_array_33_47_real;
  reg        [15:0]   int_reg_array_33_47_imag;
  reg        [15:0]   int_reg_array_33_48_real;
  reg        [15:0]   int_reg_array_33_48_imag;
  reg        [15:0]   int_reg_array_33_49_real;
  reg        [15:0]   int_reg_array_33_49_imag;
  reg        [15:0]   int_reg_array_21_0_real;
  reg        [15:0]   int_reg_array_21_0_imag;
  reg        [15:0]   int_reg_array_21_1_real;
  reg        [15:0]   int_reg_array_21_1_imag;
  reg        [15:0]   int_reg_array_21_2_real;
  reg        [15:0]   int_reg_array_21_2_imag;
  reg        [15:0]   int_reg_array_21_3_real;
  reg        [15:0]   int_reg_array_21_3_imag;
  reg        [15:0]   int_reg_array_21_4_real;
  reg        [15:0]   int_reg_array_21_4_imag;
  reg        [15:0]   int_reg_array_21_5_real;
  reg        [15:0]   int_reg_array_21_5_imag;
  reg        [15:0]   int_reg_array_21_6_real;
  reg        [15:0]   int_reg_array_21_6_imag;
  reg        [15:0]   int_reg_array_21_7_real;
  reg        [15:0]   int_reg_array_21_7_imag;
  reg        [15:0]   int_reg_array_21_8_real;
  reg        [15:0]   int_reg_array_21_8_imag;
  reg        [15:0]   int_reg_array_21_9_real;
  reg        [15:0]   int_reg_array_21_9_imag;
  reg        [15:0]   int_reg_array_21_10_real;
  reg        [15:0]   int_reg_array_21_10_imag;
  reg        [15:0]   int_reg_array_21_11_real;
  reg        [15:0]   int_reg_array_21_11_imag;
  reg        [15:0]   int_reg_array_21_12_real;
  reg        [15:0]   int_reg_array_21_12_imag;
  reg        [15:0]   int_reg_array_21_13_real;
  reg        [15:0]   int_reg_array_21_13_imag;
  reg        [15:0]   int_reg_array_21_14_real;
  reg        [15:0]   int_reg_array_21_14_imag;
  reg        [15:0]   int_reg_array_21_15_real;
  reg        [15:0]   int_reg_array_21_15_imag;
  reg        [15:0]   int_reg_array_21_16_real;
  reg        [15:0]   int_reg_array_21_16_imag;
  reg        [15:0]   int_reg_array_21_17_real;
  reg        [15:0]   int_reg_array_21_17_imag;
  reg        [15:0]   int_reg_array_21_18_real;
  reg        [15:0]   int_reg_array_21_18_imag;
  reg        [15:0]   int_reg_array_21_19_real;
  reg        [15:0]   int_reg_array_21_19_imag;
  reg        [15:0]   int_reg_array_21_20_real;
  reg        [15:0]   int_reg_array_21_20_imag;
  reg        [15:0]   int_reg_array_21_21_real;
  reg        [15:0]   int_reg_array_21_21_imag;
  reg        [15:0]   int_reg_array_21_22_real;
  reg        [15:0]   int_reg_array_21_22_imag;
  reg        [15:0]   int_reg_array_21_23_real;
  reg        [15:0]   int_reg_array_21_23_imag;
  reg        [15:0]   int_reg_array_21_24_real;
  reg        [15:0]   int_reg_array_21_24_imag;
  reg        [15:0]   int_reg_array_21_25_real;
  reg        [15:0]   int_reg_array_21_25_imag;
  reg        [15:0]   int_reg_array_21_26_real;
  reg        [15:0]   int_reg_array_21_26_imag;
  reg        [15:0]   int_reg_array_21_27_real;
  reg        [15:0]   int_reg_array_21_27_imag;
  reg        [15:0]   int_reg_array_21_28_real;
  reg        [15:0]   int_reg_array_21_28_imag;
  reg        [15:0]   int_reg_array_21_29_real;
  reg        [15:0]   int_reg_array_21_29_imag;
  reg        [15:0]   int_reg_array_21_30_real;
  reg        [15:0]   int_reg_array_21_30_imag;
  reg        [15:0]   int_reg_array_21_31_real;
  reg        [15:0]   int_reg_array_21_31_imag;
  reg        [15:0]   int_reg_array_21_32_real;
  reg        [15:0]   int_reg_array_21_32_imag;
  reg        [15:0]   int_reg_array_21_33_real;
  reg        [15:0]   int_reg_array_21_33_imag;
  reg        [15:0]   int_reg_array_21_34_real;
  reg        [15:0]   int_reg_array_21_34_imag;
  reg        [15:0]   int_reg_array_21_35_real;
  reg        [15:0]   int_reg_array_21_35_imag;
  reg        [15:0]   int_reg_array_21_36_real;
  reg        [15:0]   int_reg_array_21_36_imag;
  reg        [15:0]   int_reg_array_21_37_real;
  reg        [15:0]   int_reg_array_21_37_imag;
  reg        [15:0]   int_reg_array_21_38_real;
  reg        [15:0]   int_reg_array_21_38_imag;
  reg        [15:0]   int_reg_array_21_39_real;
  reg        [15:0]   int_reg_array_21_39_imag;
  reg        [15:0]   int_reg_array_21_40_real;
  reg        [15:0]   int_reg_array_21_40_imag;
  reg        [15:0]   int_reg_array_21_41_real;
  reg        [15:0]   int_reg_array_21_41_imag;
  reg        [15:0]   int_reg_array_21_42_real;
  reg        [15:0]   int_reg_array_21_42_imag;
  reg        [15:0]   int_reg_array_21_43_real;
  reg        [15:0]   int_reg_array_21_43_imag;
  reg        [15:0]   int_reg_array_21_44_real;
  reg        [15:0]   int_reg_array_21_44_imag;
  reg        [15:0]   int_reg_array_21_45_real;
  reg        [15:0]   int_reg_array_21_45_imag;
  reg        [15:0]   int_reg_array_21_46_real;
  reg        [15:0]   int_reg_array_21_46_imag;
  reg        [15:0]   int_reg_array_21_47_real;
  reg        [15:0]   int_reg_array_21_47_imag;
  reg        [15:0]   int_reg_array_21_48_real;
  reg        [15:0]   int_reg_array_21_48_imag;
  reg        [15:0]   int_reg_array_21_49_real;
  reg        [15:0]   int_reg_array_21_49_imag;
  reg        [31:0]   load_data_area_current_addr;
  reg        [31:0]   Axi4Incr_result;
  wire       [19:0]   Axi4Incr_highCat;
  wire       [0:0]    Axi4Incr_sizeValue;
  wire       [11:0]   Axi4Incr_alignMask;
  wire       [11:0]   Axi4Incr_base;
  wire       [11:0]   Axi4Incr_baseIncr;
  reg        [1:0]    _zz_1_;
  wire       [1:0]    Axi4Incr_wrapCase;
  reg        [31:0]   axi4_w_payload_data_regNext;
  wire       [5:0]    _zz_2_;
  wire       [63:0]   _zz_3_;
  wire                _zz_4_;
  wire                _zz_5_;
  wire                _zz_6_;
  wire                _zz_7_;
  wire                _zz_8_;
  wire                _zz_9_;
  wire                _zz_10_;
  wire                _zz_11_;
  wire                _zz_12_;
  wire                _zz_13_;
  wire                _zz_14_;
  wire                _zz_15_;
  wire                _zz_16_;
  wire                _zz_17_;
  wire                _zz_18_;
  wire                _zz_19_;
  wire                _zz_20_;
  wire                _zz_21_;
  wire                _zz_22_;
  wire                _zz_23_;
  wire                _zz_24_;
  wire                _zz_25_;
  wire                _zz_26_;
  wire                _zz_27_;
  wire                _zz_28_;
  wire                _zz_29_;
  wire                _zz_30_;
  wire                _zz_31_;
  wire                _zz_32_;
  wire                _zz_33_;
  wire                _zz_34_;
  wire                _zz_35_;
  wire                _zz_36_;
  wire                _zz_37_;
  wire                _zz_38_;
  wire                _zz_39_;
  wire                _zz_40_;
  wire                _zz_41_;
  wire                _zz_42_;
  wire                _zz_43_;
  wire                _zz_44_;
  wire                _zz_45_;
  wire                _zz_46_;
  wire                _zz_47_;
  wire                _zz_48_;
  wire                _zz_49_;
  wire                _zz_50_;
  wire                _zz_51_;
  wire                _zz_52_;
  wire                _zz_53_;
  wire       [31:0]   _zz_54_;
  wire       [15:0]   _zz_55_;
  wire       [15:0]   _zz_56_;
  wire       [5:0]    _zz_57_;
  wire       [63:0]   _zz_58_;
  wire                _zz_59_;
  wire                _zz_60_;
  wire                _zz_61_;
  wire                _zz_62_;
  wire                _zz_63_;
  wire                _zz_64_;
  wire                _zz_65_;
  wire                _zz_66_;
  wire                _zz_67_;
  wire                _zz_68_;
  wire                _zz_69_;
  wire                _zz_70_;
  wire                _zz_71_;
  wire                _zz_72_;
  wire                _zz_73_;
  wire                _zz_74_;
  wire                _zz_75_;
  wire                _zz_76_;
  wire                _zz_77_;
  wire                _zz_78_;
  wire                _zz_79_;
  wire                _zz_80_;
  wire                _zz_81_;
  wire                _zz_82_;
  wire                _zz_83_;
  wire                _zz_84_;
  wire                _zz_85_;
  wire                _zz_86_;
  wire                _zz_87_;
  wire                _zz_88_;
  wire                _zz_89_;
  wire                _zz_90_;
  wire                _zz_91_;
  wire                _zz_92_;
  wire                _zz_93_;
  wire                _zz_94_;
  wire                _zz_95_;
  wire                _zz_96_;
  wire                _zz_97_;
  wire                _zz_98_;
  wire                _zz_99_;
  wire                _zz_100_;
  wire                _zz_101_;
  wire                _zz_102_;
  wire                _zz_103_;
  wire                _zz_104_;
  wire                _zz_105_;
  wire                _zz_106_;
  wire                _zz_107_;
  wire                _zz_108_;
  wire       [31:0]   _zz_109_;
  wire       [15:0]   _zz_110_;
  wire       [15:0]   _zz_111_;
  wire       [5:0]    _zz_112_;
  wire       [63:0]   _zz_113_;
  wire                _zz_114_;
  wire                _zz_115_;
  wire                _zz_116_;
  wire                _zz_117_;
  wire                _zz_118_;
  wire                _zz_119_;
  wire                _zz_120_;
  wire                _zz_121_;
  wire                _zz_122_;
  wire                _zz_123_;
  wire                _zz_124_;
  wire                _zz_125_;
  wire                _zz_126_;
  wire                _zz_127_;
  wire                _zz_128_;
  wire                _zz_129_;
  wire                _zz_130_;
  wire                _zz_131_;
  wire                _zz_132_;
  wire                _zz_133_;
  wire                _zz_134_;
  wire                _zz_135_;
  wire                _zz_136_;
  wire                _zz_137_;
  wire                _zz_138_;
  wire                _zz_139_;
  wire                _zz_140_;
  wire                _zz_141_;
  wire                _zz_142_;
  wire                _zz_143_;
  wire                _zz_144_;
  wire                _zz_145_;
  wire                _zz_146_;
  wire                _zz_147_;
  wire                _zz_148_;
  wire                _zz_149_;
  wire                _zz_150_;
  wire                _zz_151_;
  wire                _zz_152_;
  wire                _zz_153_;
  wire                _zz_154_;
  wire                _zz_155_;
  wire                _zz_156_;
  wire                _zz_157_;
  wire                _zz_158_;
  wire                _zz_159_;
  wire                _zz_160_;
  wire                _zz_161_;
  wire                _zz_162_;
  wire                _zz_163_;
  wire       [31:0]   _zz_164_;
  wire       [15:0]   _zz_165_;
  wire       [15:0]   _zz_166_;
  wire       [5:0]    _zz_167_;
  wire       [63:0]   _zz_168_;
  wire                _zz_169_;
  wire                _zz_170_;
  wire                _zz_171_;
  wire                _zz_172_;
  wire                _zz_173_;
  wire                _zz_174_;
  wire                _zz_175_;
  wire                _zz_176_;
  wire                _zz_177_;
  wire                _zz_178_;
  wire                _zz_179_;
  wire                _zz_180_;
  wire                _zz_181_;
  wire                _zz_182_;
  wire                _zz_183_;
  wire                _zz_184_;
  wire                _zz_185_;
  wire                _zz_186_;
  wire                _zz_187_;
  wire                _zz_188_;
  wire                _zz_189_;
  wire                _zz_190_;
  wire                _zz_191_;
  wire                _zz_192_;
  wire                _zz_193_;
  wire                _zz_194_;
  wire                _zz_195_;
  wire                _zz_196_;
  wire                _zz_197_;
  wire                _zz_198_;
  wire                _zz_199_;
  wire                _zz_200_;
  wire                _zz_201_;
  wire                _zz_202_;
  wire                _zz_203_;
  wire                _zz_204_;
  wire                _zz_205_;
  wire                _zz_206_;
  wire                _zz_207_;
  wire                _zz_208_;
  wire                _zz_209_;
  wire                _zz_210_;
  wire                _zz_211_;
  wire                _zz_212_;
  wire                _zz_213_;
  wire                _zz_214_;
  wire                _zz_215_;
  wire                _zz_216_;
  wire                _zz_217_;
  wire                _zz_218_;
  wire       [31:0]   _zz_219_;
  wire       [15:0]   _zz_220_;
  wire       [15:0]   _zz_221_;
  wire       [5:0]    _zz_222_;
  wire       [63:0]   _zz_223_;
  wire                _zz_224_;
  wire                _zz_225_;
  wire                _zz_226_;
  wire                _zz_227_;
  wire                _zz_228_;
  wire                _zz_229_;
  wire                _zz_230_;
  wire                _zz_231_;
  wire                _zz_232_;
  wire                _zz_233_;
  wire                _zz_234_;
  wire                _zz_235_;
  wire                _zz_236_;
  wire                _zz_237_;
  wire                _zz_238_;
  wire                _zz_239_;
  wire                _zz_240_;
  wire                _zz_241_;
  wire                _zz_242_;
  wire                _zz_243_;
  wire                _zz_244_;
  wire                _zz_245_;
  wire                _zz_246_;
  wire                _zz_247_;
  wire                _zz_248_;
  wire                _zz_249_;
  wire                _zz_250_;
  wire                _zz_251_;
  wire                _zz_252_;
  wire                _zz_253_;
  wire                _zz_254_;
  wire                _zz_255_;
  wire                _zz_256_;
  wire                _zz_257_;
  wire                _zz_258_;
  wire                _zz_259_;
  wire                _zz_260_;
  wire                _zz_261_;
  wire                _zz_262_;
  wire                _zz_263_;
  wire                _zz_264_;
  wire                _zz_265_;
  wire                _zz_266_;
  wire                _zz_267_;
  wire                _zz_268_;
  wire                _zz_269_;
  wire                _zz_270_;
  wire                _zz_271_;
  wire                _zz_272_;
  wire                _zz_273_;
  wire       [31:0]   _zz_274_;
  wire       [15:0]   _zz_275_;
  wire       [15:0]   _zz_276_;
  wire       [5:0]    _zz_277_;
  wire       [63:0]   _zz_278_;
  wire                _zz_279_;
  wire                _zz_280_;
  wire                _zz_281_;
  wire                _zz_282_;
  wire                _zz_283_;
  wire                _zz_284_;
  wire                _zz_285_;
  wire                _zz_286_;
  wire                _zz_287_;
  wire                _zz_288_;
  wire                _zz_289_;
  wire                _zz_290_;
  wire                _zz_291_;
  wire                _zz_292_;
  wire                _zz_293_;
  wire                _zz_294_;
  wire                _zz_295_;
  wire                _zz_296_;
  wire                _zz_297_;
  wire                _zz_298_;
  wire                _zz_299_;
  wire                _zz_300_;
  wire                _zz_301_;
  wire                _zz_302_;
  wire                _zz_303_;
  wire                _zz_304_;
  wire                _zz_305_;
  wire                _zz_306_;
  wire                _zz_307_;
  wire                _zz_308_;
  wire                _zz_309_;
  wire                _zz_310_;
  wire                _zz_311_;
  wire                _zz_312_;
  wire                _zz_313_;
  wire                _zz_314_;
  wire                _zz_315_;
  wire                _zz_316_;
  wire                _zz_317_;
  wire                _zz_318_;
  wire                _zz_319_;
  wire                _zz_320_;
  wire                _zz_321_;
  wire                _zz_322_;
  wire                _zz_323_;
  wire                _zz_324_;
  wire                _zz_325_;
  wire                _zz_326_;
  wire                _zz_327_;
  wire                _zz_328_;
  wire       [31:0]   _zz_329_;
  wire       [15:0]   _zz_330_;
  wire       [15:0]   _zz_331_;
  wire       [5:0]    _zz_332_;
  wire       [63:0]   _zz_333_;
  wire                _zz_334_;
  wire                _zz_335_;
  wire                _zz_336_;
  wire                _zz_337_;
  wire                _zz_338_;
  wire                _zz_339_;
  wire                _zz_340_;
  wire                _zz_341_;
  wire                _zz_342_;
  wire                _zz_343_;
  wire                _zz_344_;
  wire                _zz_345_;
  wire                _zz_346_;
  wire                _zz_347_;
  wire                _zz_348_;
  wire                _zz_349_;
  wire                _zz_350_;
  wire                _zz_351_;
  wire                _zz_352_;
  wire                _zz_353_;
  wire                _zz_354_;
  wire                _zz_355_;
  wire                _zz_356_;
  wire                _zz_357_;
  wire                _zz_358_;
  wire                _zz_359_;
  wire                _zz_360_;
  wire                _zz_361_;
  wire                _zz_362_;
  wire                _zz_363_;
  wire                _zz_364_;
  wire                _zz_365_;
  wire                _zz_366_;
  wire                _zz_367_;
  wire                _zz_368_;
  wire                _zz_369_;
  wire                _zz_370_;
  wire                _zz_371_;
  wire                _zz_372_;
  wire                _zz_373_;
  wire                _zz_374_;
  wire                _zz_375_;
  wire                _zz_376_;
  wire                _zz_377_;
  wire                _zz_378_;
  wire                _zz_379_;
  wire                _zz_380_;
  wire                _zz_381_;
  wire                _zz_382_;
  wire                _zz_383_;
  wire       [31:0]   _zz_384_;
  wire       [15:0]   _zz_385_;
  wire       [15:0]   _zz_386_;
  wire       [5:0]    _zz_387_;
  wire       [63:0]   _zz_388_;
  wire                _zz_389_;
  wire                _zz_390_;
  wire                _zz_391_;
  wire                _zz_392_;
  wire                _zz_393_;
  wire                _zz_394_;
  wire                _zz_395_;
  wire                _zz_396_;
  wire                _zz_397_;
  wire                _zz_398_;
  wire                _zz_399_;
  wire                _zz_400_;
  wire                _zz_401_;
  wire                _zz_402_;
  wire                _zz_403_;
  wire                _zz_404_;
  wire                _zz_405_;
  wire                _zz_406_;
  wire                _zz_407_;
  wire                _zz_408_;
  wire                _zz_409_;
  wire                _zz_410_;
  wire                _zz_411_;
  wire                _zz_412_;
  wire                _zz_413_;
  wire                _zz_414_;
  wire                _zz_415_;
  wire                _zz_416_;
  wire                _zz_417_;
  wire                _zz_418_;
  wire                _zz_419_;
  wire                _zz_420_;
  wire                _zz_421_;
  wire                _zz_422_;
  wire                _zz_423_;
  wire                _zz_424_;
  wire                _zz_425_;
  wire                _zz_426_;
  wire                _zz_427_;
  wire                _zz_428_;
  wire                _zz_429_;
  wire                _zz_430_;
  wire                _zz_431_;
  wire                _zz_432_;
  wire                _zz_433_;
  wire                _zz_434_;
  wire                _zz_435_;
  wire                _zz_436_;
  wire                _zz_437_;
  wire                _zz_438_;
  wire       [31:0]   _zz_439_;
  wire       [15:0]   _zz_440_;
  wire       [15:0]   _zz_441_;
  wire       [5:0]    _zz_442_;
  wire       [63:0]   _zz_443_;
  wire                _zz_444_;
  wire                _zz_445_;
  wire                _zz_446_;
  wire                _zz_447_;
  wire                _zz_448_;
  wire                _zz_449_;
  wire                _zz_450_;
  wire                _zz_451_;
  wire                _zz_452_;
  wire                _zz_453_;
  wire                _zz_454_;
  wire                _zz_455_;
  wire                _zz_456_;
  wire                _zz_457_;
  wire                _zz_458_;
  wire                _zz_459_;
  wire                _zz_460_;
  wire                _zz_461_;
  wire                _zz_462_;
  wire                _zz_463_;
  wire                _zz_464_;
  wire                _zz_465_;
  wire                _zz_466_;
  wire                _zz_467_;
  wire                _zz_468_;
  wire                _zz_469_;
  wire                _zz_470_;
  wire                _zz_471_;
  wire                _zz_472_;
  wire                _zz_473_;
  wire                _zz_474_;
  wire                _zz_475_;
  wire                _zz_476_;
  wire                _zz_477_;
  wire                _zz_478_;
  wire                _zz_479_;
  wire                _zz_480_;
  wire                _zz_481_;
  wire                _zz_482_;
  wire                _zz_483_;
  wire                _zz_484_;
  wire                _zz_485_;
  wire                _zz_486_;
  wire                _zz_487_;
  wire                _zz_488_;
  wire                _zz_489_;
  wire                _zz_490_;
  wire                _zz_491_;
  wire                _zz_492_;
  wire                _zz_493_;
  wire       [31:0]   _zz_494_;
  wire       [15:0]   _zz_495_;
  wire       [15:0]   _zz_496_;
  wire       [5:0]    _zz_497_;
  wire       [63:0]   _zz_498_;
  wire                _zz_499_;
  wire                _zz_500_;
  wire                _zz_501_;
  wire                _zz_502_;
  wire                _zz_503_;
  wire                _zz_504_;
  wire                _zz_505_;
  wire                _zz_506_;
  wire                _zz_507_;
  wire                _zz_508_;
  wire                _zz_509_;
  wire                _zz_510_;
  wire                _zz_511_;
  wire                _zz_512_;
  wire                _zz_513_;
  wire                _zz_514_;
  wire                _zz_515_;
  wire                _zz_516_;
  wire                _zz_517_;
  wire                _zz_518_;
  wire                _zz_519_;
  wire                _zz_520_;
  wire                _zz_521_;
  wire                _zz_522_;
  wire                _zz_523_;
  wire                _zz_524_;
  wire                _zz_525_;
  wire                _zz_526_;
  wire                _zz_527_;
  wire                _zz_528_;
  wire                _zz_529_;
  wire                _zz_530_;
  wire                _zz_531_;
  wire                _zz_532_;
  wire                _zz_533_;
  wire                _zz_534_;
  wire                _zz_535_;
  wire                _zz_536_;
  wire                _zz_537_;
  wire                _zz_538_;
  wire                _zz_539_;
  wire                _zz_540_;
  wire                _zz_541_;
  wire                _zz_542_;
  wire                _zz_543_;
  wire                _zz_544_;
  wire                _zz_545_;
  wire                _zz_546_;
  wire                _zz_547_;
  wire                _zz_548_;
  wire       [31:0]   _zz_549_;
  wire       [15:0]   _zz_550_;
  wire       [15:0]   _zz_551_;
  wire       [5:0]    _zz_552_;
  wire       [63:0]   _zz_553_;
  wire                _zz_554_;
  wire                _zz_555_;
  wire                _zz_556_;
  wire                _zz_557_;
  wire                _zz_558_;
  wire                _zz_559_;
  wire                _zz_560_;
  wire                _zz_561_;
  wire                _zz_562_;
  wire                _zz_563_;
  wire                _zz_564_;
  wire                _zz_565_;
  wire                _zz_566_;
  wire                _zz_567_;
  wire                _zz_568_;
  wire                _zz_569_;
  wire                _zz_570_;
  wire                _zz_571_;
  wire                _zz_572_;
  wire                _zz_573_;
  wire                _zz_574_;
  wire                _zz_575_;
  wire                _zz_576_;
  wire                _zz_577_;
  wire                _zz_578_;
  wire                _zz_579_;
  wire                _zz_580_;
  wire                _zz_581_;
  wire                _zz_582_;
  wire                _zz_583_;
  wire                _zz_584_;
  wire                _zz_585_;
  wire                _zz_586_;
  wire                _zz_587_;
  wire                _zz_588_;
  wire                _zz_589_;
  wire                _zz_590_;
  wire                _zz_591_;
  wire                _zz_592_;
  wire                _zz_593_;
  wire                _zz_594_;
  wire                _zz_595_;
  wire                _zz_596_;
  wire                _zz_597_;
  wire                _zz_598_;
  wire                _zz_599_;
  wire                _zz_600_;
  wire                _zz_601_;
  wire                _zz_602_;
  wire                _zz_603_;
  wire       [31:0]   _zz_604_;
  wire       [15:0]   _zz_605_;
  wire       [15:0]   _zz_606_;
  wire       [5:0]    _zz_607_;
  wire       [63:0]   _zz_608_;
  wire                _zz_609_;
  wire                _zz_610_;
  wire                _zz_611_;
  wire                _zz_612_;
  wire                _zz_613_;
  wire                _zz_614_;
  wire                _zz_615_;
  wire                _zz_616_;
  wire                _zz_617_;
  wire                _zz_618_;
  wire                _zz_619_;
  wire                _zz_620_;
  wire                _zz_621_;
  wire                _zz_622_;
  wire                _zz_623_;
  wire                _zz_624_;
  wire                _zz_625_;
  wire                _zz_626_;
  wire                _zz_627_;
  wire                _zz_628_;
  wire                _zz_629_;
  wire                _zz_630_;
  wire                _zz_631_;
  wire                _zz_632_;
  wire                _zz_633_;
  wire                _zz_634_;
  wire                _zz_635_;
  wire                _zz_636_;
  wire                _zz_637_;
  wire                _zz_638_;
  wire                _zz_639_;
  wire                _zz_640_;
  wire                _zz_641_;
  wire                _zz_642_;
  wire                _zz_643_;
  wire                _zz_644_;
  wire                _zz_645_;
  wire                _zz_646_;
  wire                _zz_647_;
  wire                _zz_648_;
  wire                _zz_649_;
  wire                _zz_650_;
  wire                _zz_651_;
  wire                _zz_652_;
  wire                _zz_653_;
  wire                _zz_654_;
  wire                _zz_655_;
  wire                _zz_656_;
  wire                _zz_657_;
  wire                _zz_658_;
  wire       [31:0]   _zz_659_;
  wire       [15:0]   _zz_660_;
  wire       [15:0]   _zz_661_;
  wire       [5:0]    _zz_662_;
  wire       [63:0]   _zz_663_;
  wire                _zz_664_;
  wire                _zz_665_;
  wire                _zz_666_;
  wire                _zz_667_;
  wire                _zz_668_;
  wire                _zz_669_;
  wire                _zz_670_;
  wire                _zz_671_;
  wire                _zz_672_;
  wire                _zz_673_;
  wire                _zz_674_;
  wire                _zz_675_;
  wire                _zz_676_;
  wire                _zz_677_;
  wire                _zz_678_;
  wire                _zz_679_;
  wire                _zz_680_;
  wire                _zz_681_;
  wire                _zz_682_;
  wire                _zz_683_;
  wire                _zz_684_;
  wire                _zz_685_;
  wire                _zz_686_;
  wire                _zz_687_;
  wire                _zz_688_;
  wire                _zz_689_;
  wire                _zz_690_;
  wire                _zz_691_;
  wire                _zz_692_;
  wire                _zz_693_;
  wire                _zz_694_;
  wire                _zz_695_;
  wire                _zz_696_;
  wire                _zz_697_;
  wire                _zz_698_;
  wire                _zz_699_;
  wire                _zz_700_;
  wire                _zz_701_;
  wire                _zz_702_;
  wire                _zz_703_;
  wire                _zz_704_;
  wire                _zz_705_;
  wire                _zz_706_;
  wire                _zz_707_;
  wire                _zz_708_;
  wire                _zz_709_;
  wire                _zz_710_;
  wire                _zz_711_;
  wire                _zz_712_;
  wire                _zz_713_;
  wire       [31:0]   _zz_714_;
  wire       [15:0]   _zz_715_;
  wire       [15:0]   _zz_716_;
  wire       [5:0]    _zz_717_;
  wire       [63:0]   _zz_718_;
  wire                _zz_719_;
  wire                _zz_720_;
  wire                _zz_721_;
  wire                _zz_722_;
  wire                _zz_723_;
  wire                _zz_724_;
  wire                _zz_725_;
  wire                _zz_726_;
  wire                _zz_727_;
  wire                _zz_728_;
  wire                _zz_729_;
  wire                _zz_730_;
  wire                _zz_731_;
  wire                _zz_732_;
  wire                _zz_733_;
  wire                _zz_734_;
  wire                _zz_735_;
  wire                _zz_736_;
  wire                _zz_737_;
  wire                _zz_738_;
  wire                _zz_739_;
  wire                _zz_740_;
  wire                _zz_741_;
  wire                _zz_742_;
  wire                _zz_743_;
  wire                _zz_744_;
  wire                _zz_745_;
  wire                _zz_746_;
  wire                _zz_747_;
  wire                _zz_748_;
  wire                _zz_749_;
  wire                _zz_750_;
  wire                _zz_751_;
  wire                _zz_752_;
  wire                _zz_753_;
  wire                _zz_754_;
  wire                _zz_755_;
  wire                _zz_756_;
  wire                _zz_757_;
  wire                _zz_758_;
  wire                _zz_759_;
  wire                _zz_760_;
  wire                _zz_761_;
  wire                _zz_762_;
  wire                _zz_763_;
  wire                _zz_764_;
  wire                _zz_765_;
  wire                _zz_766_;
  wire                _zz_767_;
  wire                _zz_768_;
  wire       [31:0]   _zz_769_;
  wire       [15:0]   _zz_770_;
  wire       [15:0]   _zz_771_;
  wire       [5:0]    _zz_772_;
  wire       [63:0]   _zz_773_;
  wire                _zz_774_;
  wire                _zz_775_;
  wire                _zz_776_;
  wire                _zz_777_;
  wire                _zz_778_;
  wire                _zz_779_;
  wire                _zz_780_;
  wire                _zz_781_;
  wire                _zz_782_;
  wire                _zz_783_;
  wire                _zz_784_;
  wire                _zz_785_;
  wire                _zz_786_;
  wire                _zz_787_;
  wire                _zz_788_;
  wire                _zz_789_;
  wire                _zz_790_;
  wire                _zz_791_;
  wire                _zz_792_;
  wire                _zz_793_;
  wire                _zz_794_;
  wire                _zz_795_;
  wire                _zz_796_;
  wire                _zz_797_;
  wire                _zz_798_;
  wire                _zz_799_;
  wire                _zz_800_;
  wire                _zz_801_;
  wire                _zz_802_;
  wire                _zz_803_;
  wire                _zz_804_;
  wire                _zz_805_;
  wire                _zz_806_;
  wire                _zz_807_;
  wire                _zz_808_;
  wire                _zz_809_;
  wire                _zz_810_;
  wire                _zz_811_;
  wire                _zz_812_;
  wire                _zz_813_;
  wire                _zz_814_;
  wire                _zz_815_;
  wire                _zz_816_;
  wire                _zz_817_;
  wire                _zz_818_;
  wire                _zz_819_;
  wire                _zz_820_;
  wire                _zz_821_;
  wire                _zz_822_;
  wire                _zz_823_;
  wire       [31:0]   _zz_824_;
  wire       [15:0]   _zz_825_;
  wire       [15:0]   _zz_826_;
  wire       [5:0]    _zz_827_;
  wire       [63:0]   _zz_828_;
  wire                _zz_829_;
  wire                _zz_830_;
  wire                _zz_831_;
  wire                _zz_832_;
  wire                _zz_833_;
  wire                _zz_834_;
  wire                _zz_835_;
  wire                _zz_836_;
  wire                _zz_837_;
  wire                _zz_838_;
  wire                _zz_839_;
  wire                _zz_840_;
  wire                _zz_841_;
  wire                _zz_842_;
  wire                _zz_843_;
  wire                _zz_844_;
  wire                _zz_845_;
  wire                _zz_846_;
  wire                _zz_847_;
  wire                _zz_848_;
  wire                _zz_849_;
  wire                _zz_850_;
  wire                _zz_851_;
  wire                _zz_852_;
  wire                _zz_853_;
  wire                _zz_854_;
  wire                _zz_855_;
  wire                _zz_856_;
  wire                _zz_857_;
  wire                _zz_858_;
  wire                _zz_859_;
  wire                _zz_860_;
  wire                _zz_861_;
  wire                _zz_862_;
  wire                _zz_863_;
  wire                _zz_864_;
  wire                _zz_865_;
  wire                _zz_866_;
  wire                _zz_867_;
  wire                _zz_868_;
  wire                _zz_869_;
  wire                _zz_870_;
  wire                _zz_871_;
  wire                _zz_872_;
  wire                _zz_873_;
  wire                _zz_874_;
  wire                _zz_875_;
  wire                _zz_876_;
  wire                _zz_877_;
  wire                _zz_878_;
  wire       [31:0]   _zz_879_;
  wire       [15:0]   _zz_880_;
  wire       [15:0]   _zz_881_;
  wire       [5:0]    _zz_882_;
  wire       [63:0]   _zz_883_;
  wire                _zz_884_;
  wire                _zz_885_;
  wire                _zz_886_;
  wire                _zz_887_;
  wire                _zz_888_;
  wire                _zz_889_;
  wire                _zz_890_;
  wire                _zz_891_;
  wire                _zz_892_;
  wire                _zz_893_;
  wire                _zz_894_;
  wire                _zz_895_;
  wire                _zz_896_;
  wire                _zz_897_;
  wire                _zz_898_;
  wire                _zz_899_;
  wire                _zz_900_;
  wire                _zz_901_;
  wire                _zz_902_;
  wire                _zz_903_;
  wire                _zz_904_;
  wire                _zz_905_;
  wire                _zz_906_;
  wire                _zz_907_;
  wire                _zz_908_;
  wire                _zz_909_;
  wire                _zz_910_;
  wire                _zz_911_;
  wire                _zz_912_;
  wire                _zz_913_;
  wire                _zz_914_;
  wire                _zz_915_;
  wire                _zz_916_;
  wire                _zz_917_;
  wire                _zz_918_;
  wire                _zz_919_;
  wire                _zz_920_;
  wire                _zz_921_;
  wire                _zz_922_;
  wire                _zz_923_;
  wire                _zz_924_;
  wire                _zz_925_;
  wire                _zz_926_;
  wire                _zz_927_;
  wire                _zz_928_;
  wire                _zz_929_;
  wire                _zz_930_;
  wire                _zz_931_;
  wire                _zz_932_;
  wire                _zz_933_;
  wire       [31:0]   _zz_934_;
  wire       [15:0]   _zz_935_;
  wire       [15:0]   _zz_936_;
  wire       [5:0]    _zz_937_;
  wire       [63:0]   _zz_938_;
  wire                _zz_939_;
  wire                _zz_940_;
  wire                _zz_941_;
  wire                _zz_942_;
  wire                _zz_943_;
  wire                _zz_944_;
  wire                _zz_945_;
  wire                _zz_946_;
  wire                _zz_947_;
  wire                _zz_948_;
  wire                _zz_949_;
  wire                _zz_950_;
  wire                _zz_951_;
  wire                _zz_952_;
  wire                _zz_953_;
  wire                _zz_954_;
  wire                _zz_955_;
  wire                _zz_956_;
  wire                _zz_957_;
  wire                _zz_958_;
  wire                _zz_959_;
  wire                _zz_960_;
  wire                _zz_961_;
  wire                _zz_962_;
  wire                _zz_963_;
  wire                _zz_964_;
  wire                _zz_965_;
  wire                _zz_966_;
  wire                _zz_967_;
  wire                _zz_968_;
  wire                _zz_969_;
  wire                _zz_970_;
  wire                _zz_971_;
  wire                _zz_972_;
  wire                _zz_973_;
  wire                _zz_974_;
  wire                _zz_975_;
  wire                _zz_976_;
  wire                _zz_977_;
  wire                _zz_978_;
  wire                _zz_979_;
  wire                _zz_980_;
  wire                _zz_981_;
  wire                _zz_982_;
  wire                _zz_983_;
  wire                _zz_984_;
  wire                _zz_985_;
  wire                _zz_986_;
  wire                _zz_987_;
  wire                _zz_988_;
  wire       [31:0]   _zz_989_;
  wire       [15:0]   _zz_990_;
  wire       [15:0]   _zz_991_;
  wire       [5:0]    _zz_992_;
  wire       [63:0]   _zz_993_;
  wire                _zz_994_;
  wire                _zz_995_;
  wire                _zz_996_;
  wire                _zz_997_;
  wire                _zz_998_;
  wire                _zz_999_;
  wire                _zz_1000_;
  wire                _zz_1001_;
  wire                _zz_1002_;
  wire                _zz_1003_;
  wire                _zz_1004_;
  wire                _zz_1005_;
  wire                _zz_1006_;
  wire                _zz_1007_;
  wire                _zz_1008_;
  wire                _zz_1009_;
  wire                _zz_1010_;
  wire                _zz_1011_;
  wire                _zz_1012_;
  wire                _zz_1013_;
  wire                _zz_1014_;
  wire                _zz_1015_;
  wire                _zz_1016_;
  wire                _zz_1017_;
  wire                _zz_1018_;
  wire                _zz_1019_;
  wire                _zz_1020_;
  wire                _zz_1021_;
  wire                _zz_1022_;
  wire                _zz_1023_;
  wire                _zz_1024_;
  wire                _zz_1025_;
  wire                _zz_1026_;
  wire                _zz_1027_;
  wire                _zz_1028_;
  wire                _zz_1029_;
  wire                _zz_1030_;
  wire                _zz_1031_;
  wire                _zz_1032_;
  wire                _zz_1033_;
  wire                _zz_1034_;
  wire                _zz_1035_;
  wire                _zz_1036_;
  wire                _zz_1037_;
  wire                _zz_1038_;
  wire                _zz_1039_;
  wire                _zz_1040_;
  wire                _zz_1041_;
  wire                _zz_1042_;
  wire                _zz_1043_;
  wire       [31:0]   _zz_1044_;
  wire       [15:0]   _zz_1045_;
  wire       [15:0]   _zz_1046_;
  wire       [5:0]    _zz_1047_;
  wire       [63:0]   _zz_1048_;
  wire                _zz_1049_;
  wire                _zz_1050_;
  wire                _zz_1051_;
  wire                _zz_1052_;
  wire                _zz_1053_;
  wire                _zz_1054_;
  wire                _zz_1055_;
  wire                _zz_1056_;
  wire                _zz_1057_;
  wire                _zz_1058_;
  wire                _zz_1059_;
  wire                _zz_1060_;
  wire                _zz_1061_;
  wire                _zz_1062_;
  wire                _zz_1063_;
  wire                _zz_1064_;
  wire                _zz_1065_;
  wire                _zz_1066_;
  wire                _zz_1067_;
  wire                _zz_1068_;
  wire                _zz_1069_;
  wire                _zz_1070_;
  wire                _zz_1071_;
  wire                _zz_1072_;
  wire                _zz_1073_;
  wire                _zz_1074_;
  wire                _zz_1075_;
  wire                _zz_1076_;
  wire                _zz_1077_;
  wire                _zz_1078_;
  wire                _zz_1079_;
  wire                _zz_1080_;
  wire                _zz_1081_;
  wire                _zz_1082_;
  wire                _zz_1083_;
  wire                _zz_1084_;
  wire                _zz_1085_;
  wire                _zz_1086_;
  wire                _zz_1087_;
  wire                _zz_1088_;
  wire                _zz_1089_;
  wire                _zz_1090_;
  wire                _zz_1091_;
  wire                _zz_1092_;
  wire                _zz_1093_;
  wire                _zz_1094_;
  wire                _zz_1095_;
  wire                _zz_1096_;
  wire                _zz_1097_;
  wire                _zz_1098_;
  wire       [31:0]   _zz_1099_;
  wire       [15:0]   _zz_1100_;
  wire       [15:0]   _zz_1101_;
  wire       [5:0]    _zz_1102_;
  wire       [63:0]   _zz_1103_;
  wire                _zz_1104_;
  wire                _zz_1105_;
  wire                _zz_1106_;
  wire                _zz_1107_;
  wire                _zz_1108_;
  wire                _zz_1109_;
  wire                _zz_1110_;
  wire                _zz_1111_;
  wire                _zz_1112_;
  wire                _zz_1113_;
  wire                _zz_1114_;
  wire                _zz_1115_;
  wire                _zz_1116_;
  wire                _zz_1117_;
  wire                _zz_1118_;
  wire                _zz_1119_;
  wire                _zz_1120_;
  wire                _zz_1121_;
  wire                _zz_1122_;
  wire                _zz_1123_;
  wire                _zz_1124_;
  wire                _zz_1125_;
  wire                _zz_1126_;
  wire                _zz_1127_;
  wire                _zz_1128_;
  wire                _zz_1129_;
  wire                _zz_1130_;
  wire                _zz_1131_;
  wire                _zz_1132_;
  wire                _zz_1133_;
  wire                _zz_1134_;
  wire                _zz_1135_;
  wire                _zz_1136_;
  wire                _zz_1137_;
  wire                _zz_1138_;
  wire                _zz_1139_;
  wire                _zz_1140_;
  wire                _zz_1141_;
  wire                _zz_1142_;
  wire                _zz_1143_;
  wire                _zz_1144_;
  wire                _zz_1145_;
  wire                _zz_1146_;
  wire                _zz_1147_;
  wire                _zz_1148_;
  wire                _zz_1149_;
  wire                _zz_1150_;
  wire                _zz_1151_;
  wire                _zz_1152_;
  wire                _zz_1153_;
  wire       [31:0]   _zz_1154_;
  wire       [15:0]   _zz_1155_;
  wire       [15:0]   _zz_1156_;
  wire       [5:0]    _zz_1157_;
  wire       [63:0]   _zz_1158_;
  wire                _zz_1159_;
  wire                _zz_1160_;
  wire                _zz_1161_;
  wire                _zz_1162_;
  wire                _zz_1163_;
  wire                _zz_1164_;
  wire                _zz_1165_;
  wire                _zz_1166_;
  wire                _zz_1167_;
  wire                _zz_1168_;
  wire                _zz_1169_;
  wire                _zz_1170_;
  wire                _zz_1171_;
  wire                _zz_1172_;
  wire                _zz_1173_;
  wire                _zz_1174_;
  wire                _zz_1175_;
  wire                _zz_1176_;
  wire                _zz_1177_;
  wire                _zz_1178_;
  wire                _zz_1179_;
  wire                _zz_1180_;
  wire                _zz_1181_;
  wire                _zz_1182_;
  wire                _zz_1183_;
  wire                _zz_1184_;
  wire                _zz_1185_;
  wire                _zz_1186_;
  wire                _zz_1187_;
  wire                _zz_1188_;
  wire                _zz_1189_;
  wire                _zz_1190_;
  wire                _zz_1191_;
  wire                _zz_1192_;
  wire                _zz_1193_;
  wire                _zz_1194_;
  wire                _zz_1195_;
  wire                _zz_1196_;
  wire                _zz_1197_;
  wire                _zz_1198_;
  wire                _zz_1199_;
  wire                _zz_1200_;
  wire                _zz_1201_;
  wire                _zz_1202_;
  wire                _zz_1203_;
  wire                _zz_1204_;
  wire                _zz_1205_;
  wire                _zz_1206_;
  wire                _zz_1207_;
  wire                _zz_1208_;
  wire       [31:0]   _zz_1209_;
  wire       [15:0]   _zz_1210_;
  wire       [15:0]   _zz_1211_;
  wire       [5:0]    _zz_1212_;
  wire       [63:0]   _zz_1213_;
  wire                _zz_1214_;
  wire                _zz_1215_;
  wire                _zz_1216_;
  wire                _zz_1217_;
  wire                _zz_1218_;
  wire                _zz_1219_;
  wire                _zz_1220_;
  wire                _zz_1221_;
  wire                _zz_1222_;
  wire                _zz_1223_;
  wire                _zz_1224_;
  wire                _zz_1225_;
  wire                _zz_1226_;
  wire                _zz_1227_;
  wire                _zz_1228_;
  wire                _zz_1229_;
  wire                _zz_1230_;
  wire                _zz_1231_;
  wire                _zz_1232_;
  wire                _zz_1233_;
  wire                _zz_1234_;
  wire                _zz_1235_;
  wire                _zz_1236_;
  wire                _zz_1237_;
  wire                _zz_1238_;
  wire                _zz_1239_;
  wire                _zz_1240_;
  wire                _zz_1241_;
  wire                _zz_1242_;
  wire                _zz_1243_;
  wire                _zz_1244_;
  wire                _zz_1245_;
  wire                _zz_1246_;
  wire                _zz_1247_;
  wire                _zz_1248_;
  wire                _zz_1249_;
  wire                _zz_1250_;
  wire                _zz_1251_;
  wire                _zz_1252_;
  wire                _zz_1253_;
  wire                _zz_1254_;
  wire                _zz_1255_;
  wire                _zz_1256_;
  wire                _zz_1257_;
  wire                _zz_1258_;
  wire                _zz_1259_;
  wire                _zz_1260_;
  wire                _zz_1261_;
  wire                _zz_1262_;
  wire                _zz_1263_;
  wire       [31:0]   _zz_1264_;
  wire       [15:0]   _zz_1265_;
  wire       [15:0]   _zz_1266_;
  wire       [5:0]    _zz_1267_;
  wire       [63:0]   _zz_1268_;
  wire                _zz_1269_;
  wire                _zz_1270_;
  wire                _zz_1271_;
  wire                _zz_1272_;
  wire                _zz_1273_;
  wire                _zz_1274_;
  wire                _zz_1275_;
  wire                _zz_1276_;
  wire                _zz_1277_;
  wire                _zz_1278_;
  wire                _zz_1279_;
  wire                _zz_1280_;
  wire                _zz_1281_;
  wire                _zz_1282_;
  wire                _zz_1283_;
  wire                _zz_1284_;
  wire                _zz_1285_;
  wire                _zz_1286_;
  wire                _zz_1287_;
  wire                _zz_1288_;
  wire                _zz_1289_;
  wire                _zz_1290_;
  wire                _zz_1291_;
  wire                _zz_1292_;
  wire                _zz_1293_;
  wire                _zz_1294_;
  wire                _zz_1295_;
  wire                _zz_1296_;
  wire                _zz_1297_;
  wire                _zz_1298_;
  wire                _zz_1299_;
  wire                _zz_1300_;
  wire                _zz_1301_;
  wire                _zz_1302_;
  wire                _zz_1303_;
  wire                _zz_1304_;
  wire                _zz_1305_;
  wire                _zz_1306_;
  wire                _zz_1307_;
  wire                _zz_1308_;
  wire                _zz_1309_;
  wire                _zz_1310_;
  wire                _zz_1311_;
  wire                _zz_1312_;
  wire                _zz_1313_;
  wire                _zz_1314_;
  wire                _zz_1315_;
  wire                _zz_1316_;
  wire                _zz_1317_;
  wire                _zz_1318_;
  wire       [31:0]   _zz_1319_;
  wire       [15:0]   _zz_1320_;
  wire       [15:0]   _zz_1321_;
  wire       [5:0]    _zz_1322_;
  wire       [63:0]   _zz_1323_;
  wire                _zz_1324_;
  wire                _zz_1325_;
  wire                _zz_1326_;
  wire                _zz_1327_;
  wire                _zz_1328_;
  wire                _zz_1329_;
  wire                _zz_1330_;
  wire                _zz_1331_;
  wire                _zz_1332_;
  wire                _zz_1333_;
  wire                _zz_1334_;
  wire                _zz_1335_;
  wire                _zz_1336_;
  wire                _zz_1337_;
  wire                _zz_1338_;
  wire                _zz_1339_;
  wire                _zz_1340_;
  wire                _zz_1341_;
  wire                _zz_1342_;
  wire                _zz_1343_;
  wire                _zz_1344_;
  wire                _zz_1345_;
  wire                _zz_1346_;
  wire                _zz_1347_;
  wire                _zz_1348_;
  wire                _zz_1349_;
  wire                _zz_1350_;
  wire                _zz_1351_;
  wire                _zz_1352_;
  wire                _zz_1353_;
  wire                _zz_1354_;
  wire                _zz_1355_;
  wire                _zz_1356_;
  wire                _zz_1357_;
  wire                _zz_1358_;
  wire                _zz_1359_;
  wire                _zz_1360_;
  wire                _zz_1361_;
  wire                _zz_1362_;
  wire                _zz_1363_;
  wire                _zz_1364_;
  wire                _zz_1365_;
  wire                _zz_1366_;
  wire                _zz_1367_;
  wire                _zz_1368_;
  wire                _zz_1369_;
  wire                _zz_1370_;
  wire                _zz_1371_;
  wire                _zz_1372_;
  wire                _zz_1373_;
  wire       [31:0]   _zz_1374_;
  wire       [15:0]   _zz_1375_;
  wire       [15:0]   _zz_1376_;
  wire       [5:0]    _zz_1377_;
  wire       [63:0]   _zz_1378_;
  wire                _zz_1379_;
  wire                _zz_1380_;
  wire                _zz_1381_;
  wire                _zz_1382_;
  wire                _zz_1383_;
  wire                _zz_1384_;
  wire                _zz_1385_;
  wire                _zz_1386_;
  wire                _zz_1387_;
  wire                _zz_1388_;
  wire                _zz_1389_;
  wire                _zz_1390_;
  wire                _zz_1391_;
  wire                _zz_1392_;
  wire                _zz_1393_;
  wire                _zz_1394_;
  wire                _zz_1395_;
  wire                _zz_1396_;
  wire                _zz_1397_;
  wire                _zz_1398_;
  wire                _zz_1399_;
  wire                _zz_1400_;
  wire                _zz_1401_;
  wire                _zz_1402_;
  wire                _zz_1403_;
  wire                _zz_1404_;
  wire                _zz_1405_;
  wire                _zz_1406_;
  wire                _zz_1407_;
  wire                _zz_1408_;
  wire                _zz_1409_;
  wire                _zz_1410_;
  wire                _zz_1411_;
  wire                _zz_1412_;
  wire                _zz_1413_;
  wire                _zz_1414_;
  wire                _zz_1415_;
  wire                _zz_1416_;
  wire                _zz_1417_;
  wire                _zz_1418_;
  wire                _zz_1419_;
  wire                _zz_1420_;
  wire                _zz_1421_;
  wire                _zz_1422_;
  wire                _zz_1423_;
  wire                _zz_1424_;
  wire                _zz_1425_;
  wire                _zz_1426_;
  wire                _zz_1427_;
  wire                _zz_1428_;
  wire       [31:0]   _zz_1429_;
  wire       [15:0]   _zz_1430_;
  wire       [15:0]   _zz_1431_;
  wire       [5:0]    _zz_1432_;
  wire       [63:0]   _zz_1433_;
  wire                _zz_1434_;
  wire                _zz_1435_;
  wire                _zz_1436_;
  wire                _zz_1437_;
  wire                _zz_1438_;
  wire                _zz_1439_;
  wire                _zz_1440_;
  wire                _zz_1441_;
  wire                _zz_1442_;
  wire                _zz_1443_;
  wire                _zz_1444_;
  wire                _zz_1445_;
  wire                _zz_1446_;
  wire                _zz_1447_;
  wire                _zz_1448_;
  wire                _zz_1449_;
  wire                _zz_1450_;
  wire                _zz_1451_;
  wire                _zz_1452_;
  wire                _zz_1453_;
  wire                _zz_1454_;
  wire                _zz_1455_;
  wire                _zz_1456_;
  wire                _zz_1457_;
  wire                _zz_1458_;
  wire                _zz_1459_;
  wire                _zz_1460_;
  wire                _zz_1461_;
  wire                _zz_1462_;
  wire                _zz_1463_;
  wire                _zz_1464_;
  wire                _zz_1465_;
  wire                _zz_1466_;
  wire                _zz_1467_;
  wire                _zz_1468_;
  wire                _zz_1469_;
  wire                _zz_1470_;
  wire                _zz_1471_;
  wire                _zz_1472_;
  wire                _zz_1473_;
  wire                _zz_1474_;
  wire                _zz_1475_;
  wire                _zz_1476_;
  wire                _zz_1477_;
  wire                _zz_1478_;
  wire                _zz_1479_;
  wire                _zz_1480_;
  wire                _zz_1481_;
  wire                _zz_1482_;
  wire                _zz_1483_;
  wire       [31:0]   _zz_1484_;
  wire       [15:0]   _zz_1485_;
  wire       [15:0]   _zz_1486_;
  wire       [5:0]    _zz_1487_;
  wire       [63:0]   _zz_1488_;
  wire                _zz_1489_;
  wire                _zz_1490_;
  wire                _zz_1491_;
  wire                _zz_1492_;
  wire                _zz_1493_;
  wire                _zz_1494_;
  wire                _zz_1495_;
  wire                _zz_1496_;
  wire                _zz_1497_;
  wire                _zz_1498_;
  wire                _zz_1499_;
  wire                _zz_1500_;
  wire                _zz_1501_;
  wire                _zz_1502_;
  wire                _zz_1503_;
  wire                _zz_1504_;
  wire                _zz_1505_;
  wire                _zz_1506_;
  wire                _zz_1507_;
  wire                _zz_1508_;
  wire                _zz_1509_;
  wire                _zz_1510_;
  wire                _zz_1511_;
  wire                _zz_1512_;
  wire                _zz_1513_;
  wire                _zz_1514_;
  wire                _zz_1515_;
  wire                _zz_1516_;
  wire                _zz_1517_;
  wire                _zz_1518_;
  wire                _zz_1519_;
  wire                _zz_1520_;
  wire                _zz_1521_;
  wire                _zz_1522_;
  wire                _zz_1523_;
  wire                _zz_1524_;
  wire                _zz_1525_;
  wire                _zz_1526_;
  wire                _zz_1527_;
  wire                _zz_1528_;
  wire                _zz_1529_;
  wire                _zz_1530_;
  wire                _zz_1531_;
  wire                _zz_1532_;
  wire                _zz_1533_;
  wire                _zz_1534_;
  wire                _zz_1535_;
  wire                _zz_1536_;
  wire                _zz_1537_;
  wire                _zz_1538_;
  wire       [31:0]   _zz_1539_;
  wire       [15:0]   _zz_1540_;
  wire       [15:0]   _zz_1541_;
  wire       [5:0]    _zz_1542_;
  wire       [63:0]   _zz_1543_;
  wire                _zz_1544_;
  wire                _zz_1545_;
  wire                _zz_1546_;
  wire                _zz_1547_;
  wire                _zz_1548_;
  wire                _zz_1549_;
  wire                _zz_1550_;
  wire                _zz_1551_;
  wire                _zz_1552_;
  wire                _zz_1553_;
  wire                _zz_1554_;
  wire                _zz_1555_;
  wire                _zz_1556_;
  wire                _zz_1557_;
  wire                _zz_1558_;
  wire                _zz_1559_;
  wire                _zz_1560_;
  wire                _zz_1561_;
  wire                _zz_1562_;
  wire                _zz_1563_;
  wire                _zz_1564_;
  wire                _zz_1565_;
  wire                _zz_1566_;
  wire                _zz_1567_;
  wire                _zz_1568_;
  wire                _zz_1569_;
  wire                _zz_1570_;
  wire                _zz_1571_;
  wire                _zz_1572_;
  wire                _zz_1573_;
  wire                _zz_1574_;
  wire                _zz_1575_;
  wire                _zz_1576_;
  wire                _zz_1577_;
  wire                _zz_1578_;
  wire                _zz_1579_;
  wire                _zz_1580_;
  wire                _zz_1581_;
  wire                _zz_1582_;
  wire                _zz_1583_;
  wire                _zz_1584_;
  wire                _zz_1585_;
  wire                _zz_1586_;
  wire                _zz_1587_;
  wire                _zz_1588_;
  wire                _zz_1589_;
  wire                _zz_1590_;
  wire                _zz_1591_;
  wire                _zz_1592_;
  wire                _zz_1593_;
  wire       [31:0]   _zz_1594_;
  wire       [15:0]   _zz_1595_;
  wire       [15:0]   _zz_1596_;
  wire       [5:0]    _zz_1597_;
  wire       [63:0]   _zz_1598_;
  wire                _zz_1599_;
  wire                _zz_1600_;
  wire                _zz_1601_;
  wire                _zz_1602_;
  wire                _zz_1603_;
  wire                _zz_1604_;
  wire                _zz_1605_;
  wire                _zz_1606_;
  wire                _zz_1607_;
  wire                _zz_1608_;
  wire                _zz_1609_;
  wire                _zz_1610_;
  wire                _zz_1611_;
  wire                _zz_1612_;
  wire                _zz_1613_;
  wire                _zz_1614_;
  wire                _zz_1615_;
  wire                _zz_1616_;
  wire                _zz_1617_;
  wire                _zz_1618_;
  wire                _zz_1619_;
  wire                _zz_1620_;
  wire                _zz_1621_;
  wire                _zz_1622_;
  wire                _zz_1623_;
  wire                _zz_1624_;
  wire                _zz_1625_;
  wire                _zz_1626_;
  wire                _zz_1627_;
  wire                _zz_1628_;
  wire                _zz_1629_;
  wire                _zz_1630_;
  wire                _zz_1631_;
  wire                _zz_1632_;
  wire                _zz_1633_;
  wire                _zz_1634_;
  wire                _zz_1635_;
  wire                _zz_1636_;
  wire                _zz_1637_;
  wire                _zz_1638_;
  wire                _zz_1639_;
  wire                _zz_1640_;
  wire                _zz_1641_;
  wire                _zz_1642_;
  wire                _zz_1643_;
  wire                _zz_1644_;
  wire                _zz_1645_;
  wire                _zz_1646_;
  wire                _zz_1647_;
  wire                _zz_1648_;
  wire       [31:0]   _zz_1649_;
  wire       [15:0]   _zz_1650_;
  wire       [15:0]   _zz_1651_;
  wire       [5:0]    _zz_1652_;
  wire       [63:0]   _zz_1653_;
  wire                _zz_1654_;
  wire                _zz_1655_;
  wire                _zz_1656_;
  wire                _zz_1657_;
  wire                _zz_1658_;
  wire                _zz_1659_;
  wire                _zz_1660_;
  wire                _zz_1661_;
  wire                _zz_1662_;
  wire                _zz_1663_;
  wire                _zz_1664_;
  wire                _zz_1665_;
  wire                _zz_1666_;
  wire                _zz_1667_;
  wire                _zz_1668_;
  wire                _zz_1669_;
  wire                _zz_1670_;
  wire                _zz_1671_;
  wire                _zz_1672_;
  wire                _zz_1673_;
  wire                _zz_1674_;
  wire                _zz_1675_;
  wire                _zz_1676_;
  wire                _zz_1677_;
  wire                _zz_1678_;
  wire                _zz_1679_;
  wire                _zz_1680_;
  wire                _zz_1681_;
  wire                _zz_1682_;
  wire                _zz_1683_;
  wire                _zz_1684_;
  wire                _zz_1685_;
  wire                _zz_1686_;
  wire                _zz_1687_;
  wire                _zz_1688_;
  wire                _zz_1689_;
  wire                _zz_1690_;
  wire                _zz_1691_;
  wire                _zz_1692_;
  wire                _zz_1693_;
  wire                _zz_1694_;
  wire                _zz_1695_;
  wire                _zz_1696_;
  wire                _zz_1697_;
  wire                _zz_1698_;
  wire                _zz_1699_;
  wire                _zz_1700_;
  wire                _zz_1701_;
  wire                _zz_1702_;
  wire                _zz_1703_;
  wire       [31:0]   _zz_1704_;
  wire       [15:0]   _zz_1705_;
  wire       [15:0]   _zz_1706_;
  wire       [5:0]    _zz_1707_;
  wire       [63:0]   _zz_1708_;
  wire                _zz_1709_;
  wire                _zz_1710_;
  wire                _zz_1711_;
  wire                _zz_1712_;
  wire                _zz_1713_;
  wire                _zz_1714_;
  wire                _zz_1715_;
  wire                _zz_1716_;
  wire                _zz_1717_;
  wire                _zz_1718_;
  wire                _zz_1719_;
  wire                _zz_1720_;
  wire                _zz_1721_;
  wire                _zz_1722_;
  wire                _zz_1723_;
  wire                _zz_1724_;
  wire                _zz_1725_;
  wire                _zz_1726_;
  wire                _zz_1727_;
  wire                _zz_1728_;
  wire                _zz_1729_;
  wire                _zz_1730_;
  wire                _zz_1731_;
  wire                _zz_1732_;
  wire                _zz_1733_;
  wire                _zz_1734_;
  wire                _zz_1735_;
  wire                _zz_1736_;
  wire                _zz_1737_;
  wire                _zz_1738_;
  wire                _zz_1739_;
  wire                _zz_1740_;
  wire                _zz_1741_;
  wire                _zz_1742_;
  wire                _zz_1743_;
  wire                _zz_1744_;
  wire                _zz_1745_;
  wire                _zz_1746_;
  wire                _zz_1747_;
  wire                _zz_1748_;
  wire                _zz_1749_;
  wire                _zz_1750_;
  wire                _zz_1751_;
  wire                _zz_1752_;
  wire                _zz_1753_;
  wire                _zz_1754_;
  wire                _zz_1755_;
  wire                _zz_1756_;
  wire                _zz_1757_;
  wire                _zz_1758_;
  wire       [31:0]   _zz_1759_;
  wire       [15:0]   _zz_1760_;
  wire       [15:0]   _zz_1761_;
  wire       [5:0]    _zz_1762_;
  wire       [63:0]   _zz_1763_;
  wire                _zz_1764_;
  wire                _zz_1765_;
  wire                _zz_1766_;
  wire                _zz_1767_;
  wire                _zz_1768_;
  wire                _zz_1769_;
  wire                _zz_1770_;
  wire                _zz_1771_;
  wire                _zz_1772_;
  wire                _zz_1773_;
  wire                _zz_1774_;
  wire                _zz_1775_;
  wire                _zz_1776_;
  wire                _zz_1777_;
  wire                _zz_1778_;
  wire                _zz_1779_;
  wire                _zz_1780_;
  wire                _zz_1781_;
  wire                _zz_1782_;
  wire                _zz_1783_;
  wire                _zz_1784_;
  wire                _zz_1785_;
  wire                _zz_1786_;
  wire                _zz_1787_;
  wire                _zz_1788_;
  wire                _zz_1789_;
  wire                _zz_1790_;
  wire                _zz_1791_;
  wire                _zz_1792_;
  wire                _zz_1793_;
  wire                _zz_1794_;
  wire                _zz_1795_;
  wire                _zz_1796_;
  wire                _zz_1797_;
  wire                _zz_1798_;
  wire                _zz_1799_;
  wire                _zz_1800_;
  wire                _zz_1801_;
  wire                _zz_1802_;
  wire                _zz_1803_;
  wire                _zz_1804_;
  wire                _zz_1805_;
  wire                _zz_1806_;
  wire                _zz_1807_;
  wire                _zz_1808_;
  wire                _zz_1809_;
  wire                _zz_1810_;
  wire                _zz_1811_;
  wire                _zz_1812_;
  wire                _zz_1813_;
  wire       [31:0]   _zz_1814_;
  wire       [15:0]   _zz_1815_;
  wire       [15:0]   _zz_1816_;
  wire       [5:0]    _zz_1817_;
  wire       [63:0]   _zz_1818_;
  wire                _zz_1819_;
  wire                _zz_1820_;
  wire                _zz_1821_;
  wire                _zz_1822_;
  wire                _zz_1823_;
  wire                _zz_1824_;
  wire                _zz_1825_;
  wire                _zz_1826_;
  wire                _zz_1827_;
  wire                _zz_1828_;
  wire                _zz_1829_;
  wire                _zz_1830_;
  wire                _zz_1831_;
  wire                _zz_1832_;
  wire                _zz_1833_;
  wire                _zz_1834_;
  wire                _zz_1835_;
  wire                _zz_1836_;
  wire                _zz_1837_;
  wire                _zz_1838_;
  wire                _zz_1839_;
  wire                _zz_1840_;
  wire                _zz_1841_;
  wire                _zz_1842_;
  wire                _zz_1843_;
  wire                _zz_1844_;
  wire                _zz_1845_;
  wire                _zz_1846_;
  wire                _zz_1847_;
  wire                _zz_1848_;
  wire                _zz_1849_;
  wire                _zz_1850_;
  wire                _zz_1851_;
  wire                _zz_1852_;
  wire                _zz_1853_;
  wire                _zz_1854_;
  wire                _zz_1855_;
  wire                _zz_1856_;
  wire                _zz_1857_;
  wire                _zz_1858_;
  wire                _zz_1859_;
  wire                _zz_1860_;
  wire                _zz_1861_;
  wire                _zz_1862_;
  wire                _zz_1863_;
  wire                _zz_1864_;
  wire                _zz_1865_;
  wire                _zz_1866_;
  wire                _zz_1867_;
  wire                _zz_1868_;
  wire       [31:0]   _zz_1869_;
  wire       [15:0]   _zz_1870_;
  wire       [15:0]   _zz_1871_;
  wire       [5:0]    _zz_1872_;
  wire       [63:0]   _zz_1873_;
  wire                _zz_1874_;
  wire                _zz_1875_;
  wire                _zz_1876_;
  wire                _zz_1877_;
  wire                _zz_1878_;
  wire                _zz_1879_;
  wire                _zz_1880_;
  wire                _zz_1881_;
  wire                _zz_1882_;
  wire                _zz_1883_;
  wire                _zz_1884_;
  wire                _zz_1885_;
  wire                _zz_1886_;
  wire                _zz_1887_;
  wire                _zz_1888_;
  wire                _zz_1889_;
  wire                _zz_1890_;
  wire                _zz_1891_;
  wire                _zz_1892_;
  wire                _zz_1893_;
  wire                _zz_1894_;
  wire                _zz_1895_;
  wire                _zz_1896_;
  wire                _zz_1897_;
  wire                _zz_1898_;
  wire                _zz_1899_;
  wire                _zz_1900_;
  wire                _zz_1901_;
  wire                _zz_1902_;
  wire                _zz_1903_;
  wire                _zz_1904_;
  wire                _zz_1905_;
  wire                _zz_1906_;
  wire                _zz_1907_;
  wire                _zz_1908_;
  wire                _zz_1909_;
  wire                _zz_1910_;
  wire                _zz_1911_;
  wire                _zz_1912_;
  wire                _zz_1913_;
  wire                _zz_1914_;
  wire                _zz_1915_;
  wire                _zz_1916_;
  wire                _zz_1917_;
  wire                _zz_1918_;
  wire                _zz_1919_;
  wire                _zz_1920_;
  wire                _zz_1921_;
  wire                _zz_1922_;
  wire                _zz_1923_;
  wire       [31:0]   _zz_1924_;
  wire       [15:0]   _zz_1925_;
  wire       [15:0]   _zz_1926_;
  wire       [5:0]    _zz_1927_;
  wire       [63:0]   _zz_1928_;
  wire                _zz_1929_;
  wire                _zz_1930_;
  wire                _zz_1931_;
  wire                _zz_1932_;
  wire                _zz_1933_;
  wire                _zz_1934_;
  wire                _zz_1935_;
  wire                _zz_1936_;
  wire                _zz_1937_;
  wire                _zz_1938_;
  wire                _zz_1939_;
  wire                _zz_1940_;
  wire                _zz_1941_;
  wire                _zz_1942_;
  wire                _zz_1943_;
  wire                _zz_1944_;
  wire                _zz_1945_;
  wire                _zz_1946_;
  wire                _zz_1947_;
  wire                _zz_1948_;
  wire                _zz_1949_;
  wire                _zz_1950_;
  wire                _zz_1951_;
  wire                _zz_1952_;
  wire                _zz_1953_;
  wire                _zz_1954_;
  wire                _zz_1955_;
  wire                _zz_1956_;
  wire                _zz_1957_;
  wire                _zz_1958_;
  wire                _zz_1959_;
  wire                _zz_1960_;
  wire                _zz_1961_;
  wire                _zz_1962_;
  wire                _zz_1963_;
  wire                _zz_1964_;
  wire                _zz_1965_;
  wire                _zz_1966_;
  wire                _zz_1967_;
  wire                _zz_1968_;
  wire                _zz_1969_;
  wire                _zz_1970_;
  wire                _zz_1971_;
  wire                _zz_1972_;
  wire                _zz_1973_;
  wire                _zz_1974_;
  wire                _zz_1975_;
  wire                _zz_1976_;
  wire                _zz_1977_;
  wire                _zz_1978_;
  wire       [31:0]   _zz_1979_;
  wire       [15:0]   _zz_1980_;
  wire       [15:0]   _zz_1981_;
  wire       [5:0]    _zz_1982_;
  wire       [63:0]   _zz_1983_;
  wire                _zz_1984_;
  wire                _zz_1985_;
  wire                _zz_1986_;
  wire                _zz_1987_;
  wire                _zz_1988_;
  wire                _zz_1989_;
  wire                _zz_1990_;
  wire                _zz_1991_;
  wire                _zz_1992_;
  wire                _zz_1993_;
  wire                _zz_1994_;
  wire                _zz_1995_;
  wire                _zz_1996_;
  wire                _zz_1997_;
  wire                _zz_1998_;
  wire                _zz_1999_;
  wire                _zz_2000_;
  wire                _zz_2001_;
  wire                _zz_2002_;
  wire                _zz_2003_;
  wire                _zz_2004_;
  wire                _zz_2005_;
  wire                _zz_2006_;
  wire                _zz_2007_;
  wire                _zz_2008_;
  wire                _zz_2009_;
  wire                _zz_2010_;
  wire                _zz_2011_;
  wire                _zz_2012_;
  wire                _zz_2013_;
  wire                _zz_2014_;
  wire                _zz_2015_;
  wire                _zz_2016_;
  wire                _zz_2017_;
  wire                _zz_2018_;
  wire                _zz_2019_;
  wire                _zz_2020_;
  wire                _zz_2021_;
  wire                _zz_2022_;
  wire                _zz_2023_;
  wire                _zz_2024_;
  wire                _zz_2025_;
  wire                _zz_2026_;
  wire                _zz_2027_;
  wire                _zz_2028_;
  wire                _zz_2029_;
  wire                _zz_2030_;
  wire                _zz_2031_;
  wire                _zz_2032_;
  wire                _zz_2033_;
  wire       [31:0]   _zz_2034_;
  wire       [15:0]   _zz_2035_;
  wire       [15:0]   _zz_2036_;
  wire       [5:0]    _zz_2037_;
  wire       [63:0]   _zz_2038_;
  wire                _zz_2039_;
  wire                _zz_2040_;
  wire                _zz_2041_;
  wire                _zz_2042_;
  wire                _zz_2043_;
  wire                _zz_2044_;
  wire                _zz_2045_;
  wire                _zz_2046_;
  wire                _zz_2047_;
  wire                _zz_2048_;
  wire                _zz_2049_;
  wire                _zz_2050_;
  wire                _zz_2051_;
  wire                _zz_2052_;
  wire                _zz_2053_;
  wire                _zz_2054_;
  wire                _zz_2055_;
  wire                _zz_2056_;
  wire                _zz_2057_;
  wire                _zz_2058_;
  wire                _zz_2059_;
  wire                _zz_2060_;
  wire                _zz_2061_;
  wire                _zz_2062_;
  wire                _zz_2063_;
  wire                _zz_2064_;
  wire                _zz_2065_;
  wire                _zz_2066_;
  wire                _zz_2067_;
  wire                _zz_2068_;
  wire                _zz_2069_;
  wire                _zz_2070_;
  wire                _zz_2071_;
  wire                _zz_2072_;
  wire                _zz_2073_;
  wire                _zz_2074_;
  wire                _zz_2075_;
  wire                _zz_2076_;
  wire                _zz_2077_;
  wire                _zz_2078_;
  wire                _zz_2079_;
  wire                _zz_2080_;
  wire                _zz_2081_;
  wire                _zz_2082_;
  wire                _zz_2083_;
  wire                _zz_2084_;
  wire                _zz_2085_;
  wire                _zz_2086_;
  wire                _zz_2087_;
  wire                _zz_2088_;
  wire       [31:0]   _zz_2089_;
  wire       [15:0]   _zz_2090_;
  wire       [15:0]   _zz_2091_;
  wire       [5:0]    _zz_2092_;
  wire       [63:0]   _zz_2093_;
  wire                _zz_2094_;
  wire                _zz_2095_;
  wire                _zz_2096_;
  wire                _zz_2097_;
  wire                _zz_2098_;
  wire                _zz_2099_;
  wire                _zz_2100_;
  wire                _zz_2101_;
  wire                _zz_2102_;
  wire                _zz_2103_;
  wire                _zz_2104_;
  wire                _zz_2105_;
  wire                _zz_2106_;
  wire                _zz_2107_;
  wire                _zz_2108_;
  wire                _zz_2109_;
  wire                _zz_2110_;
  wire                _zz_2111_;
  wire                _zz_2112_;
  wire                _zz_2113_;
  wire                _zz_2114_;
  wire                _zz_2115_;
  wire                _zz_2116_;
  wire                _zz_2117_;
  wire                _zz_2118_;
  wire                _zz_2119_;
  wire                _zz_2120_;
  wire                _zz_2121_;
  wire                _zz_2122_;
  wire                _zz_2123_;
  wire                _zz_2124_;
  wire                _zz_2125_;
  wire                _zz_2126_;
  wire                _zz_2127_;
  wire                _zz_2128_;
  wire                _zz_2129_;
  wire                _zz_2130_;
  wire                _zz_2131_;
  wire                _zz_2132_;
  wire                _zz_2133_;
  wire                _zz_2134_;
  wire                _zz_2135_;
  wire                _zz_2136_;
  wire                _zz_2137_;
  wire                _zz_2138_;
  wire                _zz_2139_;
  wire                _zz_2140_;
  wire                _zz_2141_;
  wire                _zz_2142_;
  wire                _zz_2143_;
  wire       [31:0]   _zz_2144_;
  wire       [15:0]   _zz_2145_;
  wire       [15:0]   _zz_2146_;
  wire       [5:0]    _zz_2147_;
  wire       [63:0]   _zz_2148_;
  wire                _zz_2149_;
  wire                _zz_2150_;
  wire                _zz_2151_;
  wire                _zz_2152_;
  wire                _zz_2153_;
  wire                _zz_2154_;
  wire                _zz_2155_;
  wire                _zz_2156_;
  wire                _zz_2157_;
  wire                _zz_2158_;
  wire                _zz_2159_;
  wire                _zz_2160_;
  wire                _zz_2161_;
  wire                _zz_2162_;
  wire                _zz_2163_;
  wire                _zz_2164_;
  wire                _zz_2165_;
  wire                _zz_2166_;
  wire                _zz_2167_;
  wire                _zz_2168_;
  wire                _zz_2169_;
  wire                _zz_2170_;
  wire                _zz_2171_;
  wire                _zz_2172_;
  wire                _zz_2173_;
  wire                _zz_2174_;
  wire                _zz_2175_;
  wire                _zz_2176_;
  wire                _zz_2177_;
  wire                _zz_2178_;
  wire                _zz_2179_;
  wire                _zz_2180_;
  wire                _zz_2181_;
  wire                _zz_2182_;
  wire                _zz_2183_;
  wire                _zz_2184_;
  wire                _zz_2185_;
  wire                _zz_2186_;
  wire                _zz_2187_;
  wire                _zz_2188_;
  wire                _zz_2189_;
  wire                _zz_2190_;
  wire                _zz_2191_;
  wire                _zz_2192_;
  wire                _zz_2193_;
  wire                _zz_2194_;
  wire                _zz_2195_;
  wire                _zz_2196_;
  wire                _zz_2197_;
  wire                _zz_2198_;
  wire       [31:0]   _zz_2199_;
  wire       [15:0]   _zz_2200_;
  wire       [15:0]   _zz_2201_;
  wire       [5:0]    _zz_2202_;
  wire       [63:0]   _zz_2203_;
  wire                _zz_2204_;
  wire                _zz_2205_;
  wire                _zz_2206_;
  wire                _zz_2207_;
  wire                _zz_2208_;
  wire                _zz_2209_;
  wire                _zz_2210_;
  wire                _zz_2211_;
  wire                _zz_2212_;
  wire                _zz_2213_;
  wire                _zz_2214_;
  wire                _zz_2215_;
  wire                _zz_2216_;
  wire                _zz_2217_;
  wire                _zz_2218_;
  wire                _zz_2219_;
  wire                _zz_2220_;
  wire                _zz_2221_;
  wire                _zz_2222_;
  wire                _zz_2223_;
  wire                _zz_2224_;
  wire                _zz_2225_;
  wire                _zz_2226_;
  wire                _zz_2227_;
  wire                _zz_2228_;
  wire                _zz_2229_;
  wire                _zz_2230_;
  wire                _zz_2231_;
  wire                _zz_2232_;
  wire                _zz_2233_;
  wire                _zz_2234_;
  wire                _zz_2235_;
  wire                _zz_2236_;
  wire                _zz_2237_;
  wire                _zz_2238_;
  wire                _zz_2239_;
  wire                _zz_2240_;
  wire                _zz_2241_;
  wire                _zz_2242_;
  wire                _zz_2243_;
  wire                _zz_2244_;
  wire                _zz_2245_;
  wire                _zz_2246_;
  wire                _zz_2247_;
  wire                _zz_2248_;
  wire                _zz_2249_;
  wire                _zz_2250_;
  wire                _zz_2251_;
  wire                _zz_2252_;
  wire                _zz_2253_;
  wire       [31:0]   _zz_2254_;
  wire       [15:0]   _zz_2255_;
  wire       [15:0]   _zz_2256_;
  wire       [5:0]    _zz_2257_;
  wire       [63:0]   _zz_2258_;
  wire                _zz_2259_;
  wire                _zz_2260_;
  wire                _zz_2261_;
  wire                _zz_2262_;
  wire                _zz_2263_;
  wire                _zz_2264_;
  wire                _zz_2265_;
  wire                _zz_2266_;
  wire                _zz_2267_;
  wire                _zz_2268_;
  wire                _zz_2269_;
  wire                _zz_2270_;
  wire                _zz_2271_;
  wire                _zz_2272_;
  wire                _zz_2273_;
  wire                _zz_2274_;
  wire                _zz_2275_;
  wire                _zz_2276_;
  wire                _zz_2277_;
  wire                _zz_2278_;
  wire                _zz_2279_;
  wire                _zz_2280_;
  wire                _zz_2281_;
  wire                _zz_2282_;
  wire                _zz_2283_;
  wire                _zz_2284_;
  wire                _zz_2285_;
  wire                _zz_2286_;
  wire                _zz_2287_;
  wire                _zz_2288_;
  wire                _zz_2289_;
  wire                _zz_2290_;
  wire                _zz_2291_;
  wire                _zz_2292_;
  wire                _zz_2293_;
  wire                _zz_2294_;
  wire                _zz_2295_;
  wire                _zz_2296_;
  wire                _zz_2297_;
  wire                _zz_2298_;
  wire                _zz_2299_;
  wire                _zz_2300_;
  wire                _zz_2301_;
  wire                _zz_2302_;
  wire                _zz_2303_;
  wire                _zz_2304_;
  wire                _zz_2305_;
  wire                _zz_2306_;
  wire                _zz_2307_;
  wire                _zz_2308_;
  wire       [31:0]   _zz_2309_;
  wire       [15:0]   _zz_2310_;
  wire       [15:0]   _zz_2311_;
  wire       [5:0]    _zz_2312_;
  wire       [63:0]   _zz_2313_;
  wire                _zz_2314_;
  wire                _zz_2315_;
  wire                _zz_2316_;
  wire                _zz_2317_;
  wire                _zz_2318_;
  wire                _zz_2319_;
  wire                _zz_2320_;
  wire                _zz_2321_;
  wire                _zz_2322_;
  wire                _zz_2323_;
  wire                _zz_2324_;
  wire                _zz_2325_;
  wire                _zz_2326_;
  wire                _zz_2327_;
  wire                _zz_2328_;
  wire                _zz_2329_;
  wire                _zz_2330_;
  wire                _zz_2331_;
  wire                _zz_2332_;
  wire                _zz_2333_;
  wire                _zz_2334_;
  wire                _zz_2335_;
  wire                _zz_2336_;
  wire                _zz_2337_;
  wire                _zz_2338_;
  wire                _zz_2339_;
  wire                _zz_2340_;
  wire                _zz_2341_;
  wire                _zz_2342_;
  wire                _zz_2343_;
  wire                _zz_2344_;
  wire                _zz_2345_;
  wire                _zz_2346_;
  wire                _zz_2347_;
  wire                _zz_2348_;
  wire                _zz_2349_;
  wire                _zz_2350_;
  wire                _zz_2351_;
  wire                _zz_2352_;
  wire                _zz_2353_;
  wire                _zz_2354_;
  wire                _zz_2355_;
  wire                _zz_2356_;
  wire                _zz_2357_;
  wire                _zz_2358_;
  wire                _zz_2359_;
  wire                _zz_2360_;
  wire                _zz_2361_;
  wire                _zz_2362_;
  wire                _zz_2363_;
  wire       [31:0]   _zz_2364_;
  wire       [15:0]   _zz_2365_;
  wire       [15:0]   _zz_2366_;
  wire       [5:0]    _zz_2367_;
  wire       [63:0]   _zz_2368_;
  wire                _zz_2369_;
  wire                _zz_2370_;
  wire                _zz_2371_;
  wire                _zz_2372_;
  wire                _zz_2373_;
  wire                _zz_2374_;
  wire                _zz_2375_;
  wire                _zz_2376_;
  wire                _zz_2377_;
  wire                _zz_2378_;
  wire                _zz_2379_;
  wire                _zz_2380_;
  wire                _zz_2381_;
  wire                _zz_2382_;
  wire                _zz_2383_;
  wire                _zz_2384_;
  wire                _zz_2385_;
  wire                _zz_2386_;
  wire                _zz_2387_;
  wire                _zz_2388_;
  wire                _zz_2389_;
  wire                _zz_2390_;
  wire                _zz_2391_;
  wire                _zz_2392_;
  wire                _zz_2393_;
  wire                _zz_2394_;
  wire                _zz_2395_;
  wire                _zz_2396_;
  wire                _zz_2397_;
  wire                _zz_2398_;
  wire                _zz_2399_;
  wire                _zz_2400_;
  wire                _zz_2401_;
  wire                _zz_2402_;
  wire                _zz_2403_;
  wire                _zz_2404_;
  wire                _zz_2405_;
  wire                _zz_2406_;
  wire                _zz_2407_;
  wire                _zz_2408_;
  wire                _zz_2409_;
  wire                _zz_2410_;
  wire                _zz_2411_;
  wire                _zz_2412_;
  wire                _zz_2413_;
  wire                _zz_2414_;
  wire                _zz_2415_;
  wire                _zz_2416_;
  wire                _zz_2417_;
  wire                _zz_2418_;
  wire       [31:0]   _zz_2419_;
  wire       [15:0]   _zz_2420_;
  wire       [15:0]   _zz_2421_;
  wire       [5:0]    _zz_2422_;
  wire       [63:0]   _zz_2423_;
  wire                _zz_2424_;
  wire                _zz_2425_;
  wire                _zz_2426_;
  wire                _zz_2427_;
  wire                _zz_2428_;
  wire                _zz_2429_;
  wire                _zz_2430_;
  wire                _zz_2431_;
  wire                _zz_2432_;
  wire                _zz_2433_;
  wire                _zz_2434_;
  wire                _zz_2435_;
  wire                _zz_2436_;
  wire                _zz_2437_;
  wire                _zz_2438_;
  wire                _zz_2439_;
  wire                _zz_2440_;
  wire                _zz_2441_;
  wire                _zz_2442_;
  wire                _zz_2443_;
  wire                _zz_2444_;
  wire                _zz_2445_;
  wire                _zz_2446_;
  wire                _zz_2447_;
  wire                _zz_2448_;
  wire                _zz_2449_;
  wire                _zz_2450_;
  wire                _zz_2451_;
  wire                _zz_2452_;
  wire                _zz_2453_;
  wire                _zz_2454_;
  wire                _zz_2455_;
  wire                _zz_2456_;
  wire                _zz_2457_;
  wire                _zz_2458_;
  wire                _zz_2459_;
  wire                _zz_2460_;
  wire                _zz_2461_;
  wire                _zz_2462_;
  wire                _zz_2463_;
  wire                _zz_2464_;
  wire                _zz_2465_;
  wire                _zz_2466_;
  wire                _zz_2467_;
  wire                _zz_2468_;
  wire                _zz_2469_;
  wire                _zz_2470_;
  wire                _zz_2471_;
  wire                _zz_2472_;
  wire                _zz_2473_;
  wire       [31:0]   _zz_2474_;
  wire       [15:0]   _zz_2475_;
  wire       [15:0]   _zz_2476_;
  wire       [5:0]    _zz_2477_;
  wire       [63:0]   _zz_2478_;
  wire                _zz_2479_;
  wire                _zz_2480_;
  wire                _zz_2481_;
  wire                _zz_2482_;
  wire                _zz_2483_;
  wire                _zz_2484_;
  wire                _zz_2485_;
  wire                _zz_2486_;
  wire                _zz_2487_;
  wire                _zz_2488_;
  wire                _zz_2489_;
  wire                _zz_2490_;
  wire                _zz_2491_;
  wire                _zz_2492_;
  wire                _zz_2493_;
  wire                _zz_2494_;
  wire                _zz_2495_;
  wire                _zz_2496_;
  wire                _zz_2497_;
  wire                _zz_2498_;
  wire                _zz_2499_;
  wire                _zz_2500_;
  wire                _zz_2501_;
  wire                _zz_2502_;
  wire                _zz_2503_;
  wire                _zz_2504_;
  wire                _zz_2505_;
  wire                _zz_2506_;
  wire                _zz_2507_;
  wire                _zz_2508_;
  wire                _zz_2509_;
  wire                _zz_2510_;
  wire                _zz_2511_;
  wire                _zz_2512_;
  wire                _zz_2513_;
  wire                _zz_2514_;
  wire                _zz_2515_;
  wire                _zz_2516_;
  wire                _zz_2517_;
  wire                _zz_2518_;
  wire                _zz_2519_;
  wire                _zz_2520_;
  wire                _zz_2521_;
  wire                _zz_2522_;
  wire                _zz_2523_;
  wire                _zz_2524_;
  wire                _zz_2525_;
  wire                _zz_2526_;
  wire                _zz_2527_;
  wire                _zz_2528_;
  wire       [31:0]   _zz_2529_;
  wire       [15:0]   _zz_2530_;
  wire       [15:0]   _zz_2531_;
  wire       [5:0]    _zz_2532_;
  wire       [63:0]   _zz_2533_;
  wire                _zz_2534_;
  wire                _zz_2535_;
  wire                _zz_2536_;
  wire                _zz_2537_;
  wire                _zz_2538_;
  wire                _zz_2539_;
  wire                _zz_2540_;
  wire                _zz_2541_;
  wire                _zz_2542_;
  wire                _zz_2543_;
  wire                _zz_2544_;
  wire                _zz_2545_;
  wire                _zz_2546_;
  wire                _zz_2547_;
  wire                _zz_2548_;
  wire                _zz_2549_;
  wire                _zz_2550_;
  wire                _zz_2551_;
  wire                _zz_2552_;
  wire                _zz_2553_;
  wire                _zz_2554_;
  wire                _zz_2555_;
  wire                _zz_2556_;
  wire                _zz_2557_;
  wire                _zz_2558_;
  wire                _zz_2559_;
  wire                _zz_2560_;
  wire                _zz_2561_;
  wire                _zz_2562_;
  wire                _zz_2563_;
  wire                _zz_2564_;
  wire                _zz_2565_;
  wire                _zz_2566_;
  wire                _zz_2567_;
  wire                _zz_2568_;
  wire                _zz_2569_;
  wire                _zz_2570_;
  wire                _zz_2571_;
  wire                _zz_2572_;
  wire                _zz_2573_;
  wire                _zz_2574_;
  wire                _zz_2575_;
  wire                _zz_2576_;
  wire                _zz_2577_;
  wire                _zz_2578_;
  wire                _zz_2579_;
  wire                _zz_2580_;
  wire                _zz_2581_;
  wire                _zz_2582_;
  wire                _zz_2583_;
  wire       [31:0]   _zz_2584_;
  wire       [15:0]   _zz_2585_;
  wire       [15:0]   _zz_2586_;
  wire       [5:0]    _zz_2587_;
  wire       [63:0]   _zz_2588_;
  wire                _zz_2589_;
  wire                _zz_2590_;
  wire                _zz_2591_;
  wire                _zz_2592_;
  wire                _zz_2593_;
  wire                _zz_2594_;
  wire                _zz_2595_;
  wire                _zz_2596_;
  wire                _zz_2597_;
  wire                _zz_2598_;
  wire                _zz_2599_;
  wire                _zz_2600_;
  wire                _zz_2601_;
  wire                _zz_2602_;
  wire                _zz_2603_;
  wire                _zz_2604_;
  wire                _zz_2605_;
  wire                _zz_2606_;
  wire                _zz_2607_;
  wire                _zz_2608_;
  wire                _zz_2609_;
  wire                _zz_2610_;
  wire                _zz_2611_;
  wire                _zz_2612_;
  wire                _zz_2613_;
  wire                _zz_2614_;
  wire                _zz_2615_;
  wire                _zz_2616_;
  wire                _zz_2617_;
  wire                _zz_2618_;
  wire                _zz_2619_;
  wire                _zz_2620_;
  wire                _zz_2621_;
  wire                _zz_2622_;
  wire                _zz_2623_;
  wire                _zz_2624_;
  wire                _zz_2625_;
  wire                _zz_2626_;
  wire                _zz_2627_;
  wire                _zz_2628_;
  wire                _zz_2629_;
  wire                _zz_2630_;
  wire                _zz_2631_;
  wire                _zz_2632_;
  wire                _zz_2633_;
  wire                _zz_2634_;
  wire                _zz_2635_;
  wire                _zz_2636_;
  wire                _zz_2637_;
  wire                _zz_2638_;
  wire       [31:0]   _zz_2639_;
  wire       [15:0]   _zz_2640_;
  wire       [15:0]   _zz_2641_;
  wire       [5:0]    _zz_2642_;
  wire       [63:0]   _zz_2643_;
  wire                _zz_2644_;
  wire                _zz_2645_;
  wire                _zz_2646_;
  wire                _zz_2647_;
  wire                _zz_2648_;
  wire                _zz_2649_;
  wire                _zz_2650_;
  wire                _zz_2651_;
  wire                _zz_2652_;
  wire                _zz_2653_;
  wire                _zz_2654_;
  wire                _zz_2655_;
  wire                _zz_2656_;
  wire                _zz_2657_;
  wire                _zz_2658_;
  wire                _zz_2659_;
  wire                _zz_2660_;
  wire                _zz_2661_;
  wire                _zz_2662_;
  wire                _zz_2663_;
  wire                _zz_2664_;
  wire                _zz_2665_;
  wire                _zz_2666_;
  wire                _zz_2667_;
  wire                _zz_2668_;
  wire                _zz_2669_;
  wire                _zz_2670_;
  wire                _zz_2671_;
  wire                _zz_2672_;
  wire                _zz_2673_;
  wire                _zz_2674_;
  wire                _zz_2675_;
  wire                _zz_2676_;
  wire                _zz_2677_;
  wire                _zz_2678_;
  wire                _zz_2679_;
  wire                _zz_2680_;
  wire                _zz_2681_;
  wire                _zz_2682_;
  wire                _zz_2683_;
  wire                _zz_2684_;
  wire                _zz_2685_;
  wire                _zz_2686_;
  wire                _zz_2687_;
  wire                _zz_2688_;
  wire                _zz_2689_;
  wire                _zz_2690_;
  wire                _zz_2691_;
  wire                _zz_2692_;
  wire                _zz_2693_;
  wire       [31:0]   _zz_2694_;
  wire       [15:0]   _zz_2695_;
  wire       [15:0]   _zz_2696_;
  wire       [5:0]    _zz_2697_;
  wire       [63:0]   _zz_2698_;
  wire                _zz_2699_;
  wire                _zz_2700_;
  wire                _zz_2701_;
  wire                _zz_2702_;
  wire                _zz_2703_;
  wire                _zz_2704_;
  wire                _zz_2705_;
  wire                _zz_2706_;
  wire                _zz_2707_;
  wire                _zz_2708_;
  wire                _zz_2709_;
  wire                _zz_2710_;
  wire                _zz_2711_;
  wire                _zz_2712_;
  wire                _zz_2713_;
  wire                _zz_2714_;
  wire                _zz_2715_;
  wire                _zz_2716_;
  wire                _zz_2717_;
  wire                _zz_2718_;
  wire                _zz_2719_;
  wire                _zz_2720_;
  wire                _zz_2721_;
  wire                _zz_2722_;
  wire                _zz_2723_;
  wire                _zz_2724_;
  wire                _zz_2725_;
  wire                _zz_2726_;
  wire                _zz_2727_;
  wire                _zz_2728_;
  wire                _zz_2729_;
  wire                _zz_2730_;
  wire                _zz_2731_;
  wire                _zz_2732_;
  wire                _zz_2733_;
  wire                _zz_2734_;
  wire                _zz_2735_;
  wire                _zz_2736_;
  wire                _zz_2737_;
  wire                _zz_2738_;
  wire                _zz_2739_;
  wire                _zz_2740_;
  wire                _zz_2741_;
  wire                _zz_2742_;
  wire                _zz_2743_;
  wire                _zz_2744_;
  wire                _zz_2745_;
  wire                _zz_2746_;
  wire                _zz_2747_;
  wire                _zz_2748_;
  wire       [31:0]   _zz_2749_;
  wire       [15:0]   _zz_2750_;
  wire       [15:0]   _zz_2751_;

  assign _zz_2853_ = aw_area_awaddr_r[11 : 0];
  assign _zz_2854_ = _zz_2853_;
  assign _zz_2855_ = {11'd0, Axi4Incr_sizeValue};
  assign _zz_2856_ = transfer_done;
  assign _zz_2857_ = (load_data_area_current_addr - 32'h00000064);
  assign _zz_2858_ = (load_data_area_current_addr - 32'h0000028a);
  assign _zz_2859_ = (load_data_area_current_addr - 32'h000002bc);
  assign _zz_2860_ = (load_data_area_current_addr - 32'h000003b6);
  assign _zz_2861_ = (load_data_area_current_addr - 32'h00000672);
  assign _zz_2862_ = (load_data_area_current_addr - 32'h00000352);
  assign _zz_2863_ = (load_data_area_current_addr - 32'h00000320);
  assign _zz_2864_ = (load_data_area_current_addr - 32'h00000226);
  assign _zz_2865_ = (load_data_area_current_addr - 32'h000001f4);
  assign _zz_2866_ = (load_data_area_current_addr - 32'h0000073a);
  assign _zz_2867_ = (load_data_area_current_addr - 32'h0000047e);
  assign _zz_2868_ = (load_data_area_current_addr - 32'h0000041a);
  assign _zz_2869_ = (load_data_area_current_addr - 32'h000008ca);
  assign _zz_2870_ = (load_data_area_current_addr - 32'h00000898);
  assign _zz_2871_ = (load_data_area_current_addr - 32'h000004b0);
  assign _zz_2872_ = (load_data_area_current_addr - 32'h00000834);
  assign _zz_2873_ = (load_data_area_current_addr - 32'h000005dc);
  assign _zz_2874_ = (load_data_area_current_addr - 32'h00000640);
  assign _zz_2875_ = (load_data_area_current_addr - 32'h00000546);
  assign _zz_2876_ = (load_data_area_current_addr - 32'h000004e2);
  assign _zz_2877_ = (load_data_area_current_addr - 32'h00000258);
  assign _zz_2878_ = (load_data_area_current_addr - 32'h00000992);
  assign _zz_2879_ = (load_data_area_current_addr - 32'h000003e8);
  assign _zz_2880_ = (load_data_area_current_addr - 32'h000005aa);
  assign _zz_2881_ = (load_data_area_current_addr - 32'h00000802);
  assign _zz_2882_ = (load_data_area_current_addr - 32'h0000076c);
  assign _zz_2883_ = (load_data_area_current_addr - 32'h00000096);
  assign _zz_2884_ = (load_data_area_current_addr - 32'h000006a4);
  assign _zz_2885_ = (load_data_area_current_addr - 32'h0000015e);
  assign _zz_2886_ = (load_data_area_current_addr - 32'h000001c2);
  assign _zz_2887_ = (load_data_area_current_addr - 32'h00000190);
  assign _zz_2888_ = (load_data_area_current_addr - 32'h00000384);
  assign _zz_2889_ = (load_data_area_current_addr - 32'h00000866);
  assign _zz_2890_ = (load_data_area_current_addr - 32'h00000960);
  assign _zz_2891_ = (load_data_area_current_addr - 32'h00000578);
  assign _zz_2892_ = (load_data_area_current_addr - 32'h000006d6);
  assign _zz_2893_ = (load_data_area_current_addr - 32'h000000c8);
  assign _zz_2894_ = (load_data_area_current_addr - 32'h00000032);
  assign _zz_2895_ = (load_data_area_current_addr - 32'h000002ee);
  assign _zz_2896_ = (load_data_area_current_addr - 32'h000008fc);
  assign _zz_2897_ = (load_data_area_current_addr - 32'h0);
  assign _zz_2898_ = (load_data_area_current_addr - 32'h0000044c);
  assign _zz_2899_ = (load_data_area_current_addr - 32'h00000514);
  assign _zz_2900_ = (load_data_area_current_addr - 32'h0000092e);
  assign _zz_2901_ = (load_data_area_current_addr - 32'h00000708);
  assign _zz_2902_ = (load_data_area_current_addr - 32'h0000060e);
  assign _zz_2903_ = (load_data_area_current_addr - 32'h000000fa);
  assign _zz_2904_ = (load_data_area_current_addr - 32'h000007d0);
  assign _zz_2905_ = (load_data_area_current_addr - 32'h0000079e);
  assign _zz_2906_ = (load_data_area_current_addr - 32'h0000012c);
  always @(*) begin
    case(Axi4Incr_wrapCase)
      2'b00 : begin
        _zz_2752_ = {Axi4Incr_base[11 : 1],Axi4Incr_baseIncr[0 : 0]};
      end
      2'b01 : begin
        _zz_2752_ = {Axi4Incr_base[11 : 2],Axi4Incr_baseIncr[1 : 0]};
      end
      2'b10 : begin
        _zz_2752_ = {Axi4Incr_base[11 : 3],Axi4Incr_baseIncr[2 : 0]};
      end
      default : begin
        _zz_2752_ = {Axi4Incr_base[11 : 4],Axi4Incr_baseIncr[3 : 0]};
      end
    endcase
  end

  always @(*) begin
    case(_zz_2_)
      6'b000000 : begin
        _zz_2753_ = int_reg_array_0_0_imag;
        _zz_2754_ = int_reg_array_0_0_real;
      end
      6'b000001 : begin
        _zz_2753_ = int_reg_array_0_1_imag;
        _zz_2754_ = int_reg_array_0_1_real;
      end
      6'b000010 : begin
        _zz_2753_ = int_reg_array_0_2_imag;
        _zz_2754_ = int_reg_array_0_2_real;
      end
      6'b000011 : begin
        _zz_2753_ = int_reg_array_0_3_imag;
        _zz_2754_ = int_reg_array_0_3_real;
      end
      6'b000100 : begin
        _zz_2753_ = int_reg_array_0_4_imag;
        _zz_2754_ = int_reg_array_0_4_real;
      end
      6'b000101 : begin
        _zz_2753_ = int_reg_array_0_5_imag;
        _zz_2754_ = int_reg_array_0_5_real;
      end
      6'b000110 : begin
        _zz_2753_ = int_reg_array_0_6_imag;
        _zz_2754_ = int_reg_array_0_6_real;
      end
      6'b000111 : begin
        _zz_2753_ = int_reg_array_0_7_imag;
        _zz_2754_ = int_reg_array_0_7_real;
      end
      6'b001000 : begin
        _zz_2753_ = int_reg_array_0_8_imag;
        _zz_2754_ = int_reg_array_0_8_real;
      end
      6'b001001 : begin
        _zz_2753_ = int_reg_array_0_9_imag;
        _zz_2754_ = int_reg_array_0_9_real;
      end
      6'b001010 : begin
        _zz_2753_ = int_reg_array_0_10_imag;
        _zz_2754_ = int_reg_array_0_10_real;
      end
      6'b001011 : begin
        _zz_2753_ = int_reg_array_0_11_imag;
        _zz_2754_ = int_reg_array_0_11_real;
      end
      6'b001100 : begin
        _zz_2753_ = int_reg_array_0_12_imag;
        _zz_2754_ = int_reg_array_0_12_real;
      end
      6'b001101 : begin
        _zz_2753_ = int_reg_array_0_13_imag;
        _zz_2754_ = int_reg_array_0_13_real;
      end
      6'b001110 : begin
        _zz_2753_ = int_reg_array_0_14_imag;
        _zz_2754_ = int_reg_array_0_14_real;
      end
      6'b001111 : begin
        _zz_2753_ = int_reg_array_0_15_imag;
        _zz_2754_ = int_reg_array_0_15_real;
      end
      6'b010000 : begin
        _zz_2753_ = int_reg_array_0_16_imag;
        _zz_2754_ = int_reg_array_0_16_real;
      end
      6'b010001 : begin
        _zz_2753_ = int_reg_array_0_17_imag;
        _zz_2754_ = int_reg_array_0_17_real;
      end
      6'b010010 : begin
        _zz_2753_ = int_reg_array_0_18_imag;
        _zz_2754_ = int_reg_array_0_18_real;
      end
      6'b010011 : begin
        _zz_2753_ = int_reg_array_0_19_imag;
        _zz_2754_ = int_reg_array_0_19_real;
      end
      6'b010100 : begin
        _zz_2753_ = int_reg_array_0_20_imag;
        _zz_2754_ = int_reg_array_0_20_real;
      end
      6'b010101 : begin
        _zz_2753_ = int_reg_array_0_21_imag;
        _zz_2754_ = int_reg_array_0_21_real;
      end
      6'b010110 : begin
        _zz_2753_ = int_reg_array_0_22_imag;
        _zz_2754_ = int_reg_array_0_22_real;
      end
      6'b010111 : begin
        _zz_2753_ = int_reg_array_0_23_imag;
        _zz_2754_ = int_reg_array_0_23_real;
      end
      6'b011000 : begin
        _zz_2753_ = int_reg_array_0_24_imag;
        _zz_2754_ = int_reg_array_0_24_real;
      end
      6'b011001 : begin
        _zz_2753_ = int_reg_array_0_25_imag;
        _zz_2754_ = int_reg_array_0_25_real;
      end
      6'b011010 : begin
        _zz_2753_ = int_reg_array_0_26_imag;
        _zz_2754_ = int_reg_array_0_26_real;
      end
      6'b011011 : begin
        _zz_2753_ = int_reg_array_0_27_imag;
        _zz_2754_ = int_reg_array_0_27_real;
      end
      6'b011100 : begin
        _zz_2753_ = int_reg_array_0_28_imag;
        _zz_2754_ = int_reg_array_0_28_real;
      end
      6'b011101 : begin
        _zz_2753_ = int_reg_array_0_29_imag;
        _zz_2754_ = int_reg_array_0_29_real;
      end
      6'b011110 : begin
        _zz_2753_ = int_reg_array_0_30_imag;
        _zz_2754_ = int_reg_array_0_30_real;
      end
      6'b011111 : begin
        _zz_2753_ = int_reg_array_0_31_imag;
        _zz_2754_ = int_reg_array_0_31_real;
      end
      6'b100000 : begin
        _zz_2753_ = int_reg_array_0_32_imag;
        _zz_2754_ = int_reg_array_0_32_real;
      end
      6'b100001 : begin
        _zz_2753_ = int_reg_array_0_33_imag;
        _zz_2754_ = int_reg_array_0_33_real;
      end
      6'b100010 : begin
        _zz_2753_ = int_reg_array_0_34_imag;
        _zz_2754_ = int_reg_array_0_34_real;
      end
      6'b100011 : begin
        _zz_2753_ = int_reg_array_0_35_imag;
        _zz_2754_ = int_reg_array_0_35_real;
      end
      6'b100100 : begin
        _zz_2753_ = int_reg_array_0_36_imag;
        _zz_2754_ = int_reg_array_0_36_real;
      end
      6'b100101 : begin
        _zz_2753_ = int_reg_array_0_37_imag;
        _zz_2754_ = int_reg_array_0_37_real;
      end
      6'b100110 : begin
        _zz_2753_ = int_reg_array_0_38_imag;
        _zz_2754_ = int_reg_array_0_38_real;
      end
      6'b100111 : begin
        _zz_2753_ = int_reg_array_0_39_imag;
        _zz_2754_ = int_reg_array_0_39_real;
      end
      6'b101000 : begin
        _zz_2753_ = int_reg_array_0_40_imag;
        _zz_2754_ = int_reg_array_0_40_real;
      end
      6'b101001 : begin
        _zz_2753_ = int_reg_array_0_41_imag;
        _zz_2754_ = int_reg_array_0_41_real;
      end
      6'b101010 : begin
        _zz_2753_ = int_reg_array_0_42_imag;
        _zz_2754_ = int_reg_array_0_42_real;
      end
      6'b101011 : begin
        _zz_2753_ = int_reg_array_0_43_imag;
        _zz_2754_ = int_reg_array_0_43_real;
      end
      6'b101100 : begin
        _zz_2753_ = int_reg_array_0_44_imag;
        _zz_2754_ = int_reg_array_0_44_real;
      end
      6'b101101 : begin
        _zz_2753_ = int_reg_array_0_45_imag;
        _zz_2754_ = int_reg_array_0_45_real;
      end
      6'b101110 : begin
        _zz_2753_ = int_reg_array_0_46_imag;
        _zz_2754_ = int_reg_array_0_46_real;
      end
      6'b101111 : begin
        _zz_2753_ = int_reg_array_0_47_imag;
        _zz_2754_ = int_reg_array_0_47_real;
      end
      6'b110000 : begin
        _zz_2753_ = int_reg_array_0_48_imag;
        _zz_2754_ = int_reg_array_0_48_real;
      end
      default : begin
        _zz_2753_ = int_reg_array_0_49_imag;
        _zz_2754_ = int_reg_array_0_49_real;
      end
    endcase
  end

  always @(*) begin
    case(_zz_57_)
      6'b000000 : begin
        _zz_2755_ = int_reg_array_1_0_imag;
        _zz_2756_ = int_reg_array_1_0_real;
      end
      6'b000001 : begin
        _zz_2755_ = int_reg_array_1_1_imag;
        _zz_2756_ = int_reg_array_1_1_real;
      end
      6'b000010 : begin
        _zz_2755_ = int_reg_array_1_2_imag;
        _zz_2756_ = int_reg_array_1_2_real;
      end
      6'b000011 : begin
        _zz_2755_ = int_reg_array_1_3_imag;
        _zz_2756_ = int_reg_array_1_3_real;
      end
      6'b000100 : begin
        _zz_2755_ = int_reg_array_1_4_imag;
        _zz_2756_ = int_reg_array_1_4_real;
      end
      6'b000101 : begin
        _zz_2755_ = int_reg_array_1_5_imag;
        _zz_2756_ = int_reg_array_1_5_real;
      end
      6'b000110 : begin
        _zz_2755_ = int_reg_array_1_6_imag;
        _zz_2756_ = int_reg_array_1_6_real;
      end
      6'b000111 : begin
        _zz_2755_ = int_reg_array_1_7_imag;
        _zz_2756_ = int_reg_array_1_7_real;
      end
      6'b001000 : begin
        _zz_2755_ = int_reg_array_1_8_imag;
        _zz_2756_ = int_reg_array_1_8_real;
      end
      6'b001001 : begin
        _zz_2755_ = int_reg_array_1_9_imag;
        _zz_2756_ = int_reg_array_1_9_real;
      end
      6'b001010 : begin
        _zz_2755_ = int_reg_array_1_10_imag;
        _zz_2756_ = int_reg_array_1_10_real;
      end
      6'b001011 : begin
        _zz_2755_ = int_reg_array_1_11_imag;
        _zz_2756_ = int_reg_array_1_11_real;
      end
      6'b001100 : begin
        _zz_2755_ = int_reg_array_1_12_imag;
        _zz_2756_ = int_reg_array_1_12_real;
      end
      6'b001101 : begin
        _zz_2755_ = int_reg_array_1_13_imag;
        _zz_2756_ = int_reg_array_1_13_real;
      end
      6'b001110 : begin
        _zz_2755_ = int_reg_array_1_14_imag;
        _zz_2756_ = int_reg_array_1_14_real;
      end
      6'b001111 : begin
        _zz_2755_ = int_reg_array_1_15_imag;
        _zz_2756_ = int_reg_array_1_15_real;
      end
      6'b010000 : begin
        _zz_2755_ = int_reg_array_1_16_imag;
        _zz_2756_ = int_reg_array_1_16_real;
      end
      6'b010001 : begin
        _zz_2755_ = int_reg_array_1_17_imag;
        _zz_2756_ = int_reg_array_1_17_real;
      end
      6'b010010 : begin
        _zz_2755_ = int_reg_array_1_18_imag;
        _zz_2756_ = int_reg_array_1_18_real;
      end
      6'b010011 : begin
        _zz_2755_ = int_reg_array_1_19_imag;
        _zz_2756_ = int_reg_array_1_19_real;
      end
      6'b010100 : begin
        _zz_2755_ = int_reg_array_1_20_imag;
        _zz_2756_ = int_reg_array_1_20_real;
      end
      6'b010101 : begin
        _zz_2755_ = int_reg_array_1_21_imag;
        _zz_2756_ = int_reg_array_1_21_real;
      end
      6'b010110 : begin
        _zz_2755_ = int_reg_array_1_22_imag;
        _zz_2756_ = int_reg_array_1_22_real;
      end
      6'b010111 : begin
        _zz_2755_ = int_reg_array_1_23_imag;
        _zz_2756_ = int_reg_array_1_23_real;
      end
      6'b011000 : begin
        _zz_2755_ = int_reg_array_1_24_imag;
        _zz_2756_ = int_reg_array_1_24_real;
      end
      6'b011001 : begin
        _zz_2755_ = int_reg_array_1_25_imag;
        _zz_2756_ = int_reg_array_1_25_real;
      end
      6'b011010 : begin
        _zz_2755_ = int_reg_array_1_26_imag;
        _zz_2756_ = int_reg_array_1_26_real;
      end
      6'b011011 : begin
        _zz_2755_ = int_reg_array_1_27_imag;
        _zz_2756_ = int_reg_array_1_27_real;
      end
      6'b011100 : begin
        _zz_2755_ = int_reg_array_1_28_imag;
        _zz_2756_ = int_reg_array_1_28_real;
      end
      6'b011101 : begin
        _zz_2755_ = int_reg_array_1_29_imag;
        _zz_2756_ = int_reg_array_1_29_real;
      end
      6'b011110 : begin
        _zz_2755_ = int_reg_array_1_30_imag;
        _zz_2756_ = int_reg_array_1_30_real;
      end
      6'b011111 : begin
        _zz_2755_ = int_reg_array_1_31_imag;
        _zz_2756_ = int_reg_array_1_31_real;
      end
      6'b100000 : begin
        _zz_2755_ = int_reg_array_1_32_imag;
        _zz_2756_ = int_reg_array_1_32_real;
      end
      6'b100001 : begin
        _zz_2755_ = int_reg_array_1_33_imag;
        _zz_2756_ = int_reg_array_1_33_real;
      end
      6'b100010 : begin
        _zz_2755_ = int_reg_array_1_34_imag;
        _zz_2756_ = int_reg_array_1_34_real;
      end
      6'b100011 : begin
        _zz_2755_ = int_reg_array_1_35_imag;
        _zz_2756_ = int_reg_array_1_35_real;
      end
      6'b100100 : begin
        _zz_2755_ = int_reg_array_1_36_imag;
        _zz_2756_ = int_reg_array_1_36_real;
      end
      6'b100101 : begin
        _zz_2755_ = int_reg_array_1_37_imag;
        _zz_2756_ = int_reg_array_1_37_real;
      end
      6'b100110 : begin
        _zz_2755_ = int_reg_array_1_38_imag;
        _zz_2756_ = int_reg_array_1_38_real;
      end
      6'b100111 : begin
        _zz_2755_ = int_reg_array_1_39_imag;
        _zz_2756_ = int_reg_array_1_39_real;
      end
      6'b101000 : begin
        _zz_2755_ = int_reg_array_1_40_imag;
        _zz_2756_ = int_reg_array_1_40_real;
      end
      6'b101001 : begin
        _zz_2755_ = int_reg_array_1_41_imag;
        _zz_2756_ = int_reg_array_1_41_real;
      end
      6'b101010 : begin
        _zz_2755_ = int_reg_array_1_42_imag;
        _zz_2756_ = int_reg_array_1_42_real;
      end
      6'b101011 : begin
        _zz_2755_ = int_reg_array_1_43_imag;
        _zz_2756_ = int_reg_array_1_43_real;
      end
      6'b101100 : begin
        _zz_2755_ = int_reg_array_1_44_imag;
        _zz_2756_ = int_reg_array_1_44_real;
      end
      6'b101101 : begin
        _zz_2755_ = int_reg_array_1_45_imag;
        _zz_2756_ = int_reg_array_1_45_real;
      end
      6'b101110 : begin
        _zz_2755_ = int_reg_array_1_46_imag;
        _zz_2756_ = int_reg_array_1_46_real;
      end
      6'b101111 : begin
        _zz_2755_ = int_reg_array_1_47_imag;
        _zz_2756_ = int_reg_array_1_47_real;
      end
      6'b110000 : begin
        _zz_2755_ = int_reg_array_1_48_imag;
        _zz_2756_ = int_reg_array_1_48_real;
      end
      default : begin
        _zz_2755_ = int_reg_array_1_49_imag;
        _zz_2756_ = int_reg_array_1_49_real;
      end
    endcase
  end

  always @(*) begin
    case(_zz_112_)
      6'b000000 : begin
        _zz_2757_ = int_reg_array_2_0_imag;
        _zz_2758_ = int_reg_array_2_0_real;
      end
      6'b000001 : begin
        _zz_2757_ = int_reg_array_2_1_imag;
        _zz_2758_ = int_reg_array_2_1_real;
      end
      6'b000010 : begin
        _zz_2757_ = int_reg_array_2_2_imag;
        _zz_2758_ = int_reg_array_2_2_real;
      end
      6'b000011 : begin
        _zz_2757_ = int_reg_array_2_3_imag;
        _zz_2758_ = int_reg_array_2_3_real;
      end
      6'b000100 : begin
        _zz_2757_ = int_reg_array_2_4_imag;
        _zz_2758_ = int_reg_array_2_4_real;
      end
      6'b000101 : begin
        _zz_2757_ = int_reg_array_2_5_imag;
        _zz_2758_ = int_reg_array_2_5_real;
      end
      6'b000110 : begin
        _zz_2757_ = int_reg_array_2_6_imag;
        _zz_2758_ = int_reg_array_2_6_real;
      end
      6'b000111 : begin
        _zz_2757_ = int_reg_array_2_7_imag;
        _zz_2758_ = int_reg_array_2_7_real;
      end
      6'b001000 : begin
        _zz_2757_ = int_reg_array_2_8_imag;
        _zz_2758_ = int_reg_array_2_8_real;
      end
      6'b001001 : begin
        _zz_2757_ = int_reg_array_2_9_imag;
        _zz_2758_ = int_reg_array_2_9_real;
      end
      6'b001010 : begin
        _zz_2757_ = int_reg_array_2_10_imag;
        _zz_2758_ = int_reg_array_2_10_real;
      end
      6'b001011 : begin
        _zz_2757_ = int_reg_array_2_11_imag;
        _zz_2758_ = int_reg_array_2_11_real;
      end
      6'b001100 : begin
        _zz_2757_ = int_reg_array_2_12_imag;
        _zz_2758_ = int_reg_array_2_12_real;
      end
      6'b001101 : begin
        _zz_2757_ = int_reg_array_2_13_imag;
        _zz_2758_ = int_reg_array_2_13_real;
      end
      6'b001110 : begin
        _zz_2757_ = int_reg_array_2_14_imag;
        _zz_2758_ = int_reg_array_2_14_real;
      end
      6'b001111 : begin
        _zz_2757_ = int_reg_array_2_15_imag;
        _zz_2758_ = int_reg_array_2_15_real;
      end
      6'b010000 : begin
        _zz_2757_ = int_reg_array_2_16_imag;
        _zz_2758_ = int_reg_array_2_16_real;
      end
      6'b010001 : begin
        _zz_2757_ = int_reg_array_2_17_imag;
        _zz_2758_ = int_reg_array_2_17_real;
      end
      6'b010010 : begin
        _zz_2757_ = int_reg_array_2_18_imag;
        _zz_2758_ = int_reg_array_2_18_real;
      end
      6'b010011 : begin
        _zz_2757_ = int_reg_array_2_19_imag;
        _zz_2758_ = int_reg_array_2_19_real;
      end
      6'b010100 : begin
        _zz_2757_ = int_reg_array_2_20_imag;
        _zz_2758_ = int_reg_array_2_20_real;
      end
      6'b010101 : begin
        _zz_2757_ = int_reg_array_2_21_imag;
        _zz_2758_ = int_reg_array_2_21_real;
      end
      6'b010110 : begin
        _zz_2757_ = int_reg_array_2_22_imag;
        _zz_2758_ = int_reg_array_2_22_real;
      end
      6'b010111 : begin
        _zz_2757_ = int_reg_array_2_23_imag;
        _zz_2758_ = int_reg_array_2_23_real;
      end
      6'b011000 : begin
        _zz_2757_ = int_reg_array_2_24_imag;
        _zz_2758_ = int_reg_array_2_24_real;
      end
      6'b011001 : begin
        _zz_2757_ = int_reg_array_2_25_imag;
        _zz_2758_ = int_reg_array_2_25_real;
      end
      6'b011010 : begin
        _zz_2757_ = int_reg_array_2_26_imag;
        _zz_2758_ = int_reg_array_2_26_real;
      end
      6'b011011 : begin
        _zz_2757_ = int_reg_array_2_27_imag;
        _zz_2758_ = int_reg_array_2_27_real;
      end
      6'b011100 : begin
        _zz_2757_ = int_reg_array_2_28_imag;
        _zz_2758_ = int_reg_array_2_28_real;
      end
      6'b011101 : begin
        _zz_2757_ = int_reg_array_2_29_imag;
        _zz_2758_ = int_reg_array_2_29_real;
      end
      6'b011110 : begin
        _zz_2757_ = int_reg_array_2_30_imag;
        _zz_2758_ = int_reg_array_2_30_real;
      end
      6'b011111 : begin
        _zz_2757_ = int_reg_array_2_31_imag;
        _zz_2758_ = int_reg_array_2_31_real;
      end
      6'b100000 : begin
        _zz_2757_ = int_reg_array_2_32_imag;
        _zz_2758_ = int_reg_array_2_32_real;
      end
      6'b100001 : begin
        _zz_2757_ = int_reg_array_2_33_imag;
        _zz_2758_ = int_reg_array_2_33_real;
      end
      6'b100010 : begin
        _zz_2757_ = int_reg_array_2_34_imag;
        _zz_2758_ = int_reg_array_2_34_real;
      end
      6'b100011 : begin
        _zz_2757_ = int_reg_array_2_35_imag;
        _zz_2758_ = int_reg_array_2_35_real;
      end
      6'b100100 : begin
        _zz_2757_ = int_reg_array_2_36_imag;
        _zz_2758_ = int_reg_array_2_36_real;
      end
      6'b100101 : begin
        _zz_2757_ = int_reg_array_2_37_imag;
        _zz_2758_ = int_reg_array_2_37_real;
      end
      6'b100110 : begin
        _zz_2757_ = int_reg_array_2_38_imag;
        _zz_2758_ = int_reg_array_2_38_real;
      end
      6'b100111 : begin
        _zz_2757_ = int_reg_array_2_39_imag;
        _zz_2758_ = int_reg_array_2_39_real;
      end
      6'b101000 : begin
        _zz_2757_ = int_reg_array_2_40_imag;
        _zz_2758_ = int_reg_array_2_40_real;
      end
      6'b101001 : begin
        _zz_2757_ = int_reg_array_2_41_imag;
        _zz_2758_ = int_reg_array_2_41_real;
      end
      6'b101010 : begin
        _zz_2757_ = int_reg_array_2_42_imag;
        _zz_2758_ = int_reg_array_2_42_real;
      end
      6'b101011 : begin
        _zz_2757_ = int_reg_array_2_43_imag;
        _zz_2758_ = int_reg_array_2_43_real;
      end
      6'b101100 : begin
        _zz_2757_ = int_reg_array_2_44_imag;
        _zz_2758_ = int_reg_array_2_44_real;
      end
      6'b101101 : begin
        _zz_2757_ = int_reg_array_2_45_imag;
        _zz_2758_ = int_reg_array_2_45_real;
      end
      6'b101110 : begin
        _zz_2757_ = int_reg_array_2_46_imag;
        _zz_2758_ = int_reg_array_2_46_real;
      end
      6'b101111 : begin
        _zz_2757_ = int_reg_array_2_47_imag;
        _zz_2758_ = int_reg_array_2_47_real;
      end
      6'b110000 : begin
        _zz_2757_ = int_reg_array_2_48_imag;
        _zz_2758_ = int_reg_array_2_48_real;
      end
      default : begin
        _zz_2757_ = int_reg_array_2_49_imag;
        _zz_2758_ = int_reg_array_2_49_real;
      end
    endcase
  end

  always @(*) begin
    case(_zz_167_)
      6'b000000 : begin
        _zz_2759_ = int_reg_array_3_0_imag;
        _zz_2760_ = int_reg_array_3_0_real;
      end
      6'b000001 : begin
        _zz_2759_ = int_reg_array_3_1_imag;
        _zz_2760_ = int_reg_array_3_1_real;
      end
      6'b000010 : begin
        _zz_2759_ = int_reg_array_3_2_imag;
        _zz_2760_ = int_reg_array_3_2_real;
      end
      6'b000011 : begin
        _zz_2759_ = int_reg_array_3_3_imag;
        _zz_2760_ = int_reg_array_3_3_real;
      end
      6'b000100 : begin
        _zz_2759_ = int_reg_array_3_4_imag;
        _zz_2760_ = int_reg_array_3_4_real;
      end
      6'b000101 : begin
        _zz_2759_ = int_reg_array_3_5_imag;
        _zz_2760_ = int_reg_array_3_5_real;
      end
      6'b000110 : begin
        _zz_2759_ = int_reg_array_3_6_imag;
        _zz_2760_ = int_reg_array_3_6_real;
      end
      6'b000111 : begin
        _zz_2759_ = int_reg_array_3_7_imag;
        _zz_2760_ = int_reg_array_3_7_real;
      end
      6'b001000 : begin
        _zz_2759_ = int_reg_array_3_8_imag;
        _zz_2760_ = int_reg_array_3_8_real;
      end
      6'b001001 : begin
        _zz_2759_ = int_reg_array_3_9_imag;
        _zz_2760_ = int_reg_array_3_9_real;
      end
      6'b001010 : begin
        _zz_2759_ = int_reg_array_3_10_imag;
        _zz_2760_ = int_reg_array_3_10_real;
      end
      6'b001011 : begin
        _zz_2759_ = int_reg_array_3_11_imag;
        _zz_2760_ = int_reg_array_3_11_real;
      end
      6'b001100 : begin
        _zz_2759_ = int_reg_array_3_12_imag;
        _zz_2760_ = int_reg_array_3_12_real;
      end
      6'b001101 : begin
        _zz_2759_ = int_reg_array_3_13_imag;
        _zz_2760_ = int_reg_array_3_13_real;
      end
      6'b001110 : begin
        _zz_2759_ = int_reg_array_3_14_imag;
        _zz_2760_ = int_reg_array_3_14_real;
      end
      6'b001111 : begin
        _zz_2759_ = int_reg_array_3_15_imag;
        _zz_2760_ = int_reg_array_3_15_real;
      end
      6'b010000 : begin
        _zz_2759_ = int_reg_array_3_16_imag;
        _zz_2760_ = int_reg_array_3_16_real;
      end
      6'b010001 : begin
        _zz_2759_ = int_reg_array_3_17_imag;
        _zz_2760_ = int_reg_array_3_17_real;
      end
      6'b010010 : begin
        _zz_2759_ = int_reg_array_3_18_imag;
        _zz_2760_ = int_reg_array_3_18_real;
      end
      6'b010011 : begin
        _zz_2759_ = int_reg_array_3_19_imag;
        _zz_2760_ = int_reg_array_3_19_real;
      end
      6'b010100 : begin
        _zz_2759_ = int_reg_array_3_20_imag;
        _zz_2760_ = int_reg_array_3_20_real;
      end
      6'b010101 : begin
        _zz_2759_ = int_reg_array_3_21_imag;
        _zz_2760_ = int_reg_array_3_21_real;
      end
      6'b010110 : begin
        _zz_2759_ = int_reg_array_3_22_imag;
        _zz_2760_ = int_reg_array_3_22_real;
      end
      6'b010111 : begin
        _zz_2759_ = int_reg_array_3_23_imag;
        _zz_2760_ = int_reg_array_3_23_real;
      end
      6'b011000 : begin
        _zz_2759_ = int_reg_array_3_24_imag;
        _zz_2760_ = int_reg_array_3_24_real;
      end
      6'b011001 : begin
        _zz_2759_ = int_reg_array_3_25_imag;
        _zz_2760_ = int_reg_array_3_25_real;
      end
      6'b011010 : begin
        _zz_2759_ = int_reg_array_3_26_imag;
        _zz_2760_ = int_reg_array_3_26_real;
      end
      6'b011011 : begin
        _zz_2759_ = int_reg_array_3_27_imag;
        _zz_2760_ = int_reg_array_3_27_real;
      end
      6'b011100 : begin
        _zz_2759_ = int_reg_array_3_28_imag;
        _zz_2760_ = int_reg_array_3_28_real;
      end
      6'b011101 : begin
        _zz_2759_ = int_reg_array_3_29_imag;
        _zz_2760_ = int_reg_array_3_29_real;
      end
      6'b011110 : begin
        _zz_2759_ = int_reg_array_3_30_imag;
        _zz_2760_ = int_reg_array_3_30_real;
      end
      6'b011111 : begin
        _zz_2759_ = int_reg_array_3_31_imag;
        _zz_2760_ = int_reg_array_3_31_real;
      end
      6'b100000 : begin
        _zz_2759_ = int_reg_array_3_32_imag;
        _zz_2760_ = int_reg_array_3_32_real;
      end
      6'b100001 : begin
        _zz_2759_ = int_reg_array_3_33_imag;
        _zz_2760_ = int_reg_array_3_33_real;
      end
      6'b100010 : begin
        _zz_2759_ = int_reg_array_3_34_imag;
        _zz_2760_ = int_reg_array_3_34_real;
      end
      6'b100011 : begin
        _zz_2759_ = int_reg_array_3_35_imag;
        _zz_2760_ = int_reg_array_3_35_real;
      end
      6'b100100 : begin
        _zz_2759_ = int_reg_array_3_36_imag;
        _zz_2760_ = int_reg_array_3_36_real;
      end
      6'b100101 : begin
        _zz_2759_ = int_reg_array_3_37_imag;
        _zz_2760_ = int_reg_array_3_37_real;
      end
      6'b100110 : begin
        _zz_2759_ = int_reg_array_3_38_imag;
        _zz_2760_ = int_reg_array_3_38_real;
      end
      6'b100111 : begin
        _zz_2759_ = int_reg_array_3_39_imag;
        _zz_2760_ = int_reg_array_3_39_real;
      end
      6'b101000 : begin
        _zz_2759_ = int_reg_array_3_40_imag;
        _zz_2760_ = int_reg_array_3_40_real;
      end
      6'b101001 : begin
        _zz_2759_ = int_reg_array_3_41_imag;
        _zz_2760_ = int_reg_array_3_41_real;
      end
      6'b101010 : begin
        _zz_2759_ = int_reg_array_3_42_imag;
        _zz_2760_ = int_reg_array_3_42_real;
      end
      6'b101011 : begin
        _zz_2759_ = int_reg_array_3_43_imag;
        _zz_2760_ = int_reg_array_3_43_real;
      end
      6'b101100 : begin
        _zz_2759_ = int_reg_array_3_44_imag;
        _zz_2760_ = int_reg_array_3_44_real;
      end
      6'b101101 : begin
        _zz_2759_ = int_reg_array_3_45_imag;
        _zz_2760_ = int_reg_array_3_45_real;
      end
      6'b101110 : begin
        _zz_2759_ = int_reg_array_3_46_imag;
        _zz_2760_ = int_reg_array_3_46_real;
      end
      6'b101111 : begin
        _zz_2759_ = int_reg_array_3_47_imag;
        _zz_2760_ = int_reg_array_3_47_real;
      end
      6'b110000 : begin
        _zz_2759_ = int_reg_array_3_48_imag;
        _zz_2760_ = int_reg_array_3_48_real;
      end
      default : begin
        _zz_2759_ = int_reg_array_3_49_imag;
        _zz_2760_ = int_reg_array_3_49_real;
      end
    endcase
  end

  always @(*) begin
    case(_zz_222_)
      6'b000000 : begin
        _zz_2761_ = int_reg_array_4_0_imag;
        _zz_2762_ = int_reg_array_4_0_real;
      end
      6'b000001 : begin
        _zz_2761_ = int_reg_array_4_1_imag;
        _zz_2762_ = int_reg_array_4_1_real;
      end
      6'b000010 : begin
        _zz_2761_ = int_reg_array_4_2_imag;
        _zz_2762_ = int_reg_array_4_2_real;
      end
      6'b000011 : begin
        _zz_2761_ = int_reg_array_4_3_imag;
        _zz_2762_ = int_reg_array_4_3_real;
      end
      6'b000100 : begin
        _zz_2761_ = int_reg_array_4_4_imag;
        _zz_2762_ = int_reg_array_4_4_real;
      end
      6'b000101 : begin
        _zz_2761_ = int_reg_array_4_5_imag;
        _zz_2762_ = int_reg_array_4_5_real;
      end
      6'b000110 : begin
        _zz_2761_ = int_reg_array_4_6_imag;
        _zz_2762_ = int_reg_array_4_6_real;
      end
      6'b000111 : begin
        _zz_2761_ = int_reg_array_4_7_imag;
        _zz_2762_ = int_reg_array_4_7_real;
      end
      6'b001000 : begin
        _zz_2761_ = int_reg_array_4_8_imag;
        _zz_2762_ = int_reg_array_4_8_real;
      end
      6'b001001 : begin
        _zz_2761_ = int_reg_array_4_9_imag;
        _zz_2762_ = int_reg_array_4_9_real;
      end
      6'b001010 : begin
        _zz_2761_ = int_reg_array_4_10_imag;
        _zz_2762_ = int_reg_array_4_10_real;
      end
      6'b001011 : begin
        _zz_2761_ = int_reg_array_4_11_imag;
        _zz_2762_ = int_reg_array_4_11_real;
      end
      6'b001100 : begin
        _zz_2761_ = int_reg_array_4_12_imag;
        _zz_2762_ = int_reg_array_4_12_real;
      end
      6'b001101 : begin
        _zz_2761_ = int_reg_array_4_13_imag;
        _zz_2762_ = int_reg_array_4_13_real;
      end
      6'b001110 : begin
        _zz_2761_ = int_reg_array_4_14_imag;
        _zz_2762_ = int_reg_array_4_14_real;
      end
      6'b001111 : begin
        _zz_2761_ = int_reg_array_4_15_imag;
        _zz_2762_ = int_reg_array_4_15_real;
      end
      6'b010000 : begin
        _zz_2761_ = int_reg_array_4_16_imag;
        _zz_2762_ = int_reg_array_4_16_real;
      end
      6'b010001 : begin
        _zz_2761_ = int_reg_array_4_17_imag;
        _zz_2762_ = int_reg_array_4_17_real;
      end
      6'b010010 : begin
        _zz_2761_ = int_reg_array_4_18_imag;
        _zz_2762_ = int_reg_array_4_18_real;
      end
      6'b010011 : begin
        _zz_2761_ = int_reg_array_4_19_imag;
        _zz_2762_ = int_reg_array_4_19_real;
      end
      6'b010100 : begin
        _zz_2761_ = int_reg_array_4_20_imag;
        _zz_2762_ = int_reg_array_4_20_real;
      end
      6'b010101 : begin
        _zz_2761_ = int_reg_array_4_21_imag;
        _zz_2762_ = int_reg_array_4_21_real;
      end
      6'b010110 : begin
        _zz_2761_ = int_reg_array_4_22_imag;
        _zz_2762_ = int_reg_array_4_22_real;
      end
      6'b010111 : begin
        _zz_2761_ = int_reg_array_4_23_imag;
        _zz_2762_ = int_reg_array_4_23_real;
      end
      6'b011000 : begin
        _zz_2761_ = int_reg_array_4_24_imag;
        _zz_2762_ = int_reg_array_4_24_real;
      end
      6'b011001 : begin
        _zz_2761_ = int_reg_array_4_25_imag;
        _zz_2762_ = int_reg_array_4_25_real;
      end
      6'b011010 : begin
        _zz_2761_ = int_reg_array_4_26_imag;
        _zz_2762_ = int_reg_array_4_26_real;
      end
      6'b011011 : begin
        _zz_2761_ = int_reg_array_4_27_imag;
        _zz_2762_ = int_reg_array_4_27_real;
      end
      6'b011100 : begin
        _zz_2761_ = int_reg_array_4_28_imag;
        _zz_2762_ = int_reg_array_4_28_real;
      end
      6'b011101 : begin
        _zz_2761_ = int_reg_array_4_29_imag;
        _zz_2762_ = int_reg_array_4_29_real;
      end
      6'b011110 : begin
        _zz_2761_ = int_reg_array_4_30_imag;
        _zz_2762_ = int_reg_array_4_30_real;
      end
      6'b011111 : begin
        _zz_2761_ = int_reg_array_4_31_imag;
        _zz_2762_ = int_reg_array_4_31_real;
      end
      6'b100000 : begin
        _zz_2761_ = int_reg_array_4_32_imag;
        _zz_2762_ = int_reg_array_4_32_real;
      end
      6'b100001 : begin
        _zz_2761_ = int_reg_array_4_33_imag;
        _zz_2762_ = int_reg_array_4_33_real;
      end
      6'b100010 : begin
        _zz_2761_ = int_reg_array_4_34_imag;
        _zz_2762_ = int_reg_array_4_34_real;
      end
      6'b100011 : begin
        _zz_2761_ = int_reg_array_4_35_imag;
        _zz_2762_ = int_reg_array_4_35_real;
      end
      6'b100100 : begin
        _zz_2761_ = int_reg_array_4_36_imag;
        _zz_2762_ = int_reg_array_4_36_real;
      end
      6'b100101 : begin
        _zz_2761_ = int_reg_array_4_37_imag;
        _zz_2762_ = int_reg_array_4_37_real;
      end
      6'b100110 : begin
        _zz_2761_ = int_reg_array_4_38_imag;
        _zz_2762_ = int_reg_array_4_38_real;
      end
      6'b100111 : begin
        _zz_2761_ = int_reg_array_4_39_imag;
        _zz_2762_ = int_reg_array_4_39_real;
      end
      6'b101000 : begin
        _zz_2761_ = int_reg_array_4_40_imag;
        _zz_2762_ = int_reg_array_4_40_real;
      end
      6'b101001 : begin
        _zz_2761_ = int_reg_array_4_41_imag;
        _zz_2762_ = int_reg_array_4_41_real;
      end
      6'b101010 : begin
        _zz_2761_ = int_reg_array_4_42_imag;
        _zz_2762_ = int_reg_array_4_42_real;
      end
      6'b101011 : begin
        _zz_2761_ = int_reg_array_4_43_imag;
        _zz_2762_ = int_reg_array_4_43_real;
      end
      6'b101100 : begin
        _zz_2761_ = int_reg_array_4_44_imag;
        _zz_2762_ = int_reg_array_4_44_real;
      end
      6'b101101 : begin
        _zz_2761_ = int_reg_array_4_45_imag;
        _zz_2762_ = int_reg_array_4_45_real;
      end
      6'b101110 : begin
        _zz_2761_ = int_reg_array_4_46_imag;
        _zz_2762_ = int_reg_array_4_46_real;
      end
      6'b101111 : begin
        _zz_2761_ = int_reg_array_4_47_imag;
        _zz_2762_ = int_reg_array_4_47_real;
      end
      6'b110000 : begin
        _zz_2761_ = int_reg_array_4_48_imag;
        _zz_2762_ = int_reg_array_4_48_real;
      end
      default : begin
        _zz_2761_ = int_reg_array_4_49_imag;
        _zz_2762_ = int_reg_array_4_49_real;
      end
    endcase
  end

  always @(*) begin
    case(_zz_277_)
      6'b000000 : begin
        _zz_2763_ = int_reg_array_5_0_imag;
        _zz_2764_ = int_reg_array_5_0_real;
      end
      6'b000001 : begin
        _zz_2763_ = int_reg_array_5_1_imag;
        _zz_2764_ = int_reg_array_5_1_real;
      end
      6'b000010 : begin
        _zz_2763_ = int_reg_array_5_2_imag;
        _zz_2764_ = int_reg_array_5_2_real;
      end
      6'b000011 : begin
        _zz_2763_ = int_reg_array_5_3_imag;
        _zz_2764_ = int_reg_array_5_3_real;
      end
      6'b000100 : begin
        _zz_2763_ = int_reg_array_5_4_imag;
        _zz_2764_ = int_reg_array_5_4_real;
      end
      6'b000101 : begin
        _zz_2763_ = int_reg_array_5_5_imag;
        _zz_2764_ = int_reg_array_5_5_real;
      end
      6'b000110 : begin
        _zz_2763_ = int_reg_array_5_6_imag;
        _zz_2764_ = int_reg_array_5_6_real;
      end
      6'b000111 : begin
        _zz_2763_ = int_reg_array_5_7_imag;
        _zz_2764_ = int_reg_array_5_7_real;
      end
      6'b001000 : begin
        _zz_2763_ = int_reg_array_5_8_imag;
        _zz_2764_ = int_reg_array_5_8_real;
      end
      6'b001001 : begin
        _zz_2763_ = int_reg_array_5_9_imag;
        _zz_2764_ = int_reg_array_5_9_real;
      end
      6'b001010 : begin
        _zz_2763_ = int_reg_array_5_10_imag;
        _zz_2764_ = int_reg_array_5_10_real;
      end
      6'b001011 : begin
        _zz_2763_ = int_reg_array_5_11_imag;
        _zz_2764_ = int_reg_array_5_11_real;
      end
      6'b001100 : begin
        _zz_2763_ = int_reg_array_5_12_imag;
        _zz_2764_ = int_reg_array_5_12_real;
      end
      6'b001101 : begin
        _zz_2763_ = int_reg_array_5_13_imag;
        _zz_2764_ = int_reg_array_5_13_real;
      end
      6'b001110 : begin
        _zz_2763_ = int_reg_array_5_14_imag;
        _zz_2764_ = int_reg_array_5_14_real;
      end
      6'b001111 : begin
        _zz_2763_ = int_reg_array_5_15_imag;
        _zz_2764_ = int_reg_array_5_15_real;
      end
      6'b010000 : begin
        _zz_2763_ = int_reg_array_5_16_imag;
        _zz_2764_ = int_reg_array_5_16_real;
      end
      6'b010001 : begin
        _zz_2763_ = int_reg_array_5_17_imag;
        _zz_2764_ = int_reg_array_5_17_real;
      end
      6'b010010 : begin
        _zz_2763_ = int_reg_array_5_18_imag;
        _zz_2764_ = int_reg_array_5_18_real;
      end
      6'b010011 : begin
        _zz_2763_ = int_reg_array_5_19_imag;
        _zz_2764_ = int_reg_array_5_19_real;
      end
      6'b010100 : begin
        _zz_2763_ = int_reg_array_5_20_imag;
        _zz_2764_ = int_reg_array_5_20_real;
      end
      6'b010101 : begin
        _zz_2763_ = int_reg_array_5_21_imag;
        _zz_2764_ = int_reg_array_5_21_real;
      end
      6'b010110 : begin
        _zz_2763_ = int_reg_array_5_22_imag;
        _zz_2764_ = int_reg_array_5_22_real;
      end
      6'b010111 : begin
        _zz_2763_ = int_reg_array_5_23_imag;
        _zz_2764_ = int_reg_array_5_23_real;
      end
      6'b011000 : begin
        _zz_2763_ = int_reg_array_5_24_imag;
        _zz_2764_ = int_reg_array_5_24_real;
      end
      6'b011001 : begin
        _zz_2763_ = int_reg_array_5_25_imag;
        _zz_2764_ = int_reg_array_5_25_real;
      end
      6'b011010 : begin
        _zz_2763_ = int_reg_array_5_26_imag;
        _zz_2764_ = int_reg_array_5_26_real;
      end
      6'b011011 : begin
        _zz_2763_ = int_reg_array_5_27_imag;
        _zz_2764_ = int_reg_array_5_27_real;
      end
      6'b011100 : begin
        _zz_2763_ = int_reg_array_5_28_imag;
        _zz_2764_ = int_reg_array_5_28_real;
      end
      6'b011101 : begin
        _zz_2763_ = int_reg_array_5_29_imag;
        _zz_2764_ = int_reg_array_5_29_real;
      end
      6'b011110 : begin
        _zz_2763_ = int_reg_array_5_30_imag;
        _zz_2764_ = int_reg_array_5_30_real;
      end
      6'b011111 : begin
        _zz_2763_ = int_reg_array_5_31_imag;
        _zz_2764_ = int_reg_array_5_31_real;
      end
      6'b100000 : begin
        _zz_2763_ = int_reg_array_5_32_imag;
        _zz_2764_ = int_reg_array_5_32_real;
      end
      6'b100001 : begin
        _zz_2763_ = int_reg_array_5_33_imag;
        _zz_2764_ = int_reg_array_5_33_real;
      end
      6'b100010 : begin
        _zz_2763_ = int_reg_array_5_34_imag;
        _zz_2764_ = int_reg_array_5_34_real;
      end
      6'b100011 : begin
        _zz_2763_ = int_reg_array_5_35_imag;
        _zz_2764_ = int_reg_array_5_35_real;
      end
      6'b100100 : begin
        _zz_2763_ = int_reg_array_5_36_imag;
        _zz_2764_ = int_reg_array_5_36_real;
      end
      6'b100101 : begin
        _zz_2763_ = int_reg_array_5_37_imag;
        _zz_2764_ = int_reg_array_5_37_real;
      end
      6'b100110 : begin
        _zz_2763_ = int_reg_array_5_38_imag;
        _zz_2764_ = int_reg_array_5_38_real;
      end
      6'b100111 : begin
        _zz_2763_ = int_reg_array_5_39_imag;
        _zz_2764_ = int_reg_array_5_39_real;
      end
      6'b101000 : begin
        _zz_2763_ = int_reg_array_5_40_imag;
        _zz_2764_ = int_reg_array_5_40_real;
      end
      6'b101001 : begin
        _zz_2763_ = int_reg_array_5_41_imag;
        _zz_2764_ = int_reg_array_5_41_real;
      end
      6'b101010 : begin
        _zz_2763_ = int_reg_array_5_42_imag;
        _zz_2764_ = int_reg_array_5_42_real;
      end
      6'b101011 : begin
        _zz_2763_ = int_reg_array_5_43_imag;
        _zz_2764_ = int_reg_array_5_43_real;
      end
      6'b101100 : begin
        _zz_2763_ = int_reg_array_5_44_imag;
        _zz_2764_ = int_reg_array_5_44_real;
      end
      6'b101101 : begin
        _zz_2763_ = int_reg_array_5_45_imag;
        _zz_2764_ = int_reg_array_5_45_real;
      end
      6'b101110 : begin
        _zz_2763_ = int_reg_array_5_46_imag;
        _zz_2764_ = int_reg_array_5_46_real;
      end
      6'b101111 : begin
        _zz_2763_ = int_reg_array_5_47_imag;
        _zz_2764_ = int_reg_array_5_47_real;
      end
      6'b110000 : begin
        _zz_2763_ = int_reg_array_5_48_imag;
        _zz_2764_ = int_reg_array_5_48_real;
      end
      default : begin
        _zz_2763_ = int_reg_array_5_49_imag;
        _zz_2764_ = int_reg_array_5_49_real;
      end
    endcase
  end

  always @(*) begin
    case(_zz_332_)
      6'b000000 : begin
        _zz_2765_ = int_reg_array_6_0_imag;
        _zz_2766_ = int_reg_array_6_0_real;
      end
      6'b000001 : begin
        _zz_2765_ = int_reg_array_6_1_imag;
        _zz_2766_ = int_reg_array_6_1_real;
      end
      6'b000010 : begin
        _zz_2765_ = int_reg_array_6_2_imag;
        _zz_2766_ = int_reg_array_6_2_real;
      end
      6'b000011 : begin
        _zz_2765_ = int_reg_array_6_3_imag;
        _zz_2766_ = int_reg_array_6_3_real;
      end
      6'b000100 : begin
        _zz_2765_ = int_reg_array_6_4_imag;
        _zz_2766_ = int_reg_array_6_4_real;
      end
      6'b000101 : begin
        _zz_2765_ = int_reg_array_6_5_imag;
        _zz_2766_ = int_reg_array_6_5_real;
      end
      6'b000110 : begin
        _zz_2765_ = int_reg_array_6_6_imag;
        _zz_2766_ = int_reg_array_6_6_real;
      end
      6'b000111 : begin
        _zz_2765_ = int_reg_array_6_7_imag;
        _zz_2766_ = int_reg_array_6_7_real;
      end
      6'b001000 : begin
        _zz_2765_ = int_reg_array_6_8_imag;
        _zz_2766_ = int_reg_array_6_8_real;
      end
      6'b001001 : begin
        _zz_2765_ = int_reg_array_6_9_imag;
        _zz_2766_ = int_reg_array_6_9_real;
      end
      6'b001010 : begin
        _zz_2765_ = int_reg_array_6_10_imag;
        _zz_2766_ = int_reg_array_6_10_real;
      end
      6'b001011 : begin
        _zz_2765_ = int_reg_array_6_11_imag;
        _zz_2766_ = int_reg_array_6_11_real;
      end
      6'b001100 : begin
        _zz_2765_ = int_reg_array_6_12_imag;
        _zz_2766_ = int_reg_array_6_12_real;
      end
      6'b001101 : begin
        _zz_2765_ = int_reg_array_6_13_imag;
        _zz_2766_ = int_reg_array_6_13_real;
      end
      6'b001110 : begin
        _zz_2765_ = int_reg_array_6_14_imag;
        _zz_2766_ = int_reg_array_6_14_real;
      end
      6'b001111 : begin
        _zz_2765_ = int_reg_array_6_15_imag;
        _zz_2766_ = int_reg_array_6_15_real;
      end
      6'b010000 : begin
        _zz_2765_ = int_reg_array_6_16_imag;
        _zz_2766_ = int_reg_array_6_16_real;
      end
      6'b010001 : begin
        _zz_2765_ = int_reg_array_6_17_imag;
        _zz_2766_ = int_reg_array_6_17_real;
      end
      6'b010010 : begin
        _zz_2765_ = int_reg_array_6_18_imag;
        _zz_2766_ = int_reg_array_6_18_real;
      end
      6'b010011 : begin
        _zz_2765_ = int_reg_array_6_19_imag;
        _zz_2766_ = int_reg_array_6_19_real;
      end
      6'b010100 : begin
        _zz_2765_ = int_reg_array_6_20_imag;
        _zz_2766_ = int_reg_array_6_20_real;
      end
      6'b010101 : begin
        _zz_2765_ = int_reg_array_6_21_imag;
        _zz_2766_ = int_reg_array_6_21_real;
      end
      6'b010110 : begin
        _zz_2765_ = int_reg_array_6_22_imag;
        _zz_2766_ = int_reg_array_6_22_real;
      end
      6'b010111 : begin
        _zz_2765_ = int_reg_array_6_23_imag;
        _zz_2766_ = int_reg_array_6_23_real;
      end
      6'b011000 : begin
        _zz_2765_ = int_reg_array_6_24_imag;
        _zz_2766_ = int_reg_array_6_24_real;
      end
      6'b011001 : begin
        _zz_2765_ = int_reg_array_6_25_imag;
        _zz_2766_ = int_reg_array_6_25_real;
      end
      6'b011010 : begin
        _zz_2765_ = int_reg_array_6_26_imag;
        _zz_2766_ = int_reg_array_6_26_real;
      end
      6'b011011 : begin
        _zz_2765_ = int_reg_array_6_27_imag;
        _zz_2766_ = int_reg_array_6_27_real;
      end
      6'b011100 : begin
        _zz_2765_ = int_reg_array_6_28_imag;
        _zz_2766_ = int_reg_array_6_28_real;
      end
      6'b011101 : begin
        _zz_2765_ = int_reg_array_6_29_imag;
        _zz_2766_ = int_reg_array_6_29_real;
      end
      6'b011110 : begin
        _zz_2765_ = int_reg_array_6_30_imag;
        _zz_2766_ = int_reg_array_6_30_real;
      end
      6'b011111 : begin
        _zz_2765_ = int_reg_array_6_31_imag;
        _zz_2766_ = int_reg_array_6_31_real;
      end
      6'b100000 : begin
        _zz_2765_ = int_reg_array_6_32_imag;
        _zz_2766_ = int_reg_array_6_32_real;
      end
      6'b100001 : begin
        _zz_2765_ = int_reg_array_6_33_imag;
        _zz_2766_ = int_reg_array_6_33_real;
      end
      6'b100010 : begin
        _zz_2765_ = int_reg_array_6_34_imag;
        _zz_2766_ = int_reg_array_6_34_real;
      end
      6'b100011 : begin
        _zz_2765_ = int_reg_array_6_35_imag;
        _zz_2766_ = int_reg_array_6_35_real;
      end
      6'b100100 : begin
        _zz_2765_ = int_reg_array_6_36_imag;
        _zz_2766_ = int_reg_array_6_36_real;
      end
      6'b100101 : begin
        _zz_2765_ = int_reg_array_6_37_imag;
        _zz_2766_ = int_reg_array_6_37_real;
      end
      6'b100110 : begin
        _zz_2765_ = int_reg_array_6_38_imag;
        _zz_2766_ = int_reg_array_6_38_real;
      end
      6'b100111 : begin
        _zz_2765_ = int_reg_array_6_39_imag;
        _zz_2766_ = int_reg_array_6_39_real;
      end
      6'b101000 : begin
        _zz_2765_ = int_reg_array_6_40_imag;
        _zz_2766_ = int_reg_array_6_40_real;
      end
      6'b101001 : begin
        _zz_2765_ = int_reg_array_6_41_imag;
        _zz_2766_ = int_reg_array_6_41_real;
      end
      6'b101010 : begin
        _zz_2765_ = int_reg_array_6_42_imag;
        _zz_2766_ = int_reg_array_6_42_real;
      end
      6'b101011 : begin
        _zz_2765_ = int_reg_array_6_43_imag;
        _zz_2766_ = int_reg_array_6_43_real;
      end
      6'b101100 : begin
        _zz_2765_ = int_reg_array_6_44_imag;
        _zz_2766_ = int_reg_array_6_44_real;
      end
      6'b101101 : begin
        _zz_2765_ = int_reg_array_6_45_imag;
        _zz_2766_ = int_reg_array_6_45_real;
      end
      6'b101110 : begin
        _zz_2765_ = int_reg_array_6_46_imag;
        _zz_2766_ = int_reg_array_6_46_real;
      end
      6'b101111 : begin
        _zz_2765_ = int_reg_array_6_47_imag;
        _zz_2766_ = int_reg_array_6_47_real;
      end
      6'b110000 : begin
        _zz_2765_ = int_reg_array_6_48_imag;
        _zz_2766_ = int_reg_array_6_48_real;
      end
      default : begin
        _zz_2765_ = int_reg_array_6_49_imag;
        _zz_2766_ = int_reg_array_6_49_real;
      end
    endcase
  end

  always @(*) begin
    case(_zz_387_)
      6'b000000 : begin
        _zz_2767_ = int_reg_array_7_0_imag;
        _zz_2768_ = int_reg_array_7_0_real;
      end
      6'b000001 : begin
        _zz_2767_ = int_reg_array_7_1_imag;
        _zz_2768_ = int_reg_array_7_1_real;
      end
      6'b000010 : begin
        _zz_2767_ = int_reg_array_7_2_imag;
        _zz_2768_ = int_reg_array_7_2_real;
      end
      6'b000011 : begin
        _zz_2767_ = int_reg_array_7_3_imag;
        _zz_2768_ = int_reg_array_7_3_real;
      end
      6'b000100 : begin
        _zz_2767_ = int_reg_array_7_4_imag;
        _zz_2768_ = int_reg_array_7_4_real;
      end
      6'b000101 : begin
        _zz_2767_ = int_reg_array_7_5_imag;
        _zz_2768_ = int_reg_array_7_5_real;
      end
      6'b000110 : begin
        _zz_2767_ = int_reg_array_7_6_imag;
        _zz_2768_ = int_reg_array_7_6_real;
      end
      6'b000111 : begin
        _zz_2767_ = int_reg_array_7_7_imag;
        _zz_2768_ = int_reg_array_7_7_real;
      end
      6'b001000 : begin
        _zz_2767_ = int_reg_array_7_8_imag;
        _zz_2768_ = int_reg_array_7_8_real;
      end
      6'b001001 : begin
        _zz_2767_ = int_reg_array_7_9_imag;
        _zz_2768_ = int_reg_array_7_9_real;
      end
      6'b001010 : begin
        _zz_2767_ = int_reg_array_7_10_imag;
        _zz_2768_ = int_reg_array_7_10_real;
      end
      6'b001011 : begin
        _zz_2767_ = int_reg_array_7_11_imag;
        _zz_2768_ = int_reg_array_7_11_real;
      end
      6'b001100 : begin
        _zz_2767_ = int_reg_array_7_12_imag;
        _zz_2768_ = int_reg_array_7_12_real;
      end
      6'b001101 : begin
        _zz_2767_ = int_reg_array_7_13_imag;
        _zz_2768_ = int_reg_array_7_13_real;
      end
      6'b001110 : begin
        _zz_2767_ = int_reg_array_7_14_imag;
        _zz_2768_ = int_reg_array_7_14_real;
      end
      6'b001111 : begin
        _zz_2767_ = int_reg_array_7_15_imag;
        _zz_2768_ = int_reg_array_7_15_real;
      end
      6'b010000 : begin
        _zz_2767_ = int_reg_array_7_16_imag;
        _zz_2768_ = int_reg_array_7_16_real;
      end
      6'b010001 : begin
        _zz_2767_ = int_reg_array_7_17_imag;
        _zz_2768_ = int_reg_array_7_17_real;
      end
      6'b010010 : begin
        _zz_2767_ = int_reg_array_7_18_imag;
        _zz_2768_ = int_reg_array_7_18_real;
      end
      6'b010011 : begin
        _zz_2767_ = int_reg_array_7_19_imag;
        _zz_2768_ = int_reg_array_7_19_real;
      end
      6'b010100 : begin
        _zz_2767_ = int_reg_array_7_20_imag;
        _zz_2768_ = int_reg_array_7_20_real;
      end
      6'b010101 : begin
        _zz_2767_ = int_reg_array_7_21_imag;
        _zz_2768_ = int_reg_array_7_21_real;
      end
      6'b010110 : begin
        _zz_2767_ = int_reg_array_7_22_imag;
        _zz_2768_ = int_reg_array_7_22_real;
      end
      6'b010111 : begin
        _zz_2767_ = int_reg_array_7_23_imag;
        _zz_2768_ = int_reg_array_7_23_real;
      end
      6'b011000 : begin
        _zz_2767_ = int_reg_array_7_24_imag;
        _zz_2768_ = int_reg_array_7_24_real;
      end
      6'b011001 : begin
        _zz_2767_ = int_reg_array_7_25_imag;
        _zz_2768_ = int_reg_array_7_25_real;
      end
      6'b011010 : begin
        _zz_2767_ = int_reg_array_7_26_imag;
        _zz_2768_ = int_reg_array_7_26_real;
      end
      6'b011011 : begin
        _zz_2767_ = int_reg_array_7_27_imag;
        _zz_2768_ = int_reg_array_7_27_real;
      end
      6'b011100 : begin
        _zz_2767_ = int_reg_array_7_28_imag;
        _zz_2768_ = int_reg_array_7_28_real;
      end
      6'b011101 : begin
        _zz_2767_ = int_reg_array_7_29_imag;
        _zz_2768_ = int_reg_array_7_29_real;
      end
      6'b011110 : begin
        _zz_2767_ = int_reg_array_7_30_imag;
        _zz_2768_ = int_reg_array_7_30_real;
      end
      6'b011111 : begin
        _zz_2767_ = int_reg_array_7_31_imag;
        _zz_2768_ = int_reg_array_7_31_real;
      end
      6'b100000 : begin
        _zz_2767_ = int_reg_array_7_32_imag;
        _zz_2768_ = int_reg_array_7_32_real;
      end
      6'b100001 : begin
        _zz_2767_ = int_reg_array_7_33_imag;
        _zz_2768_ = int_reg_array_7_33_real;
      end
      6'b100010 : begin
        _zz_2767_ = int_reg_array_7_34_imag;
        _zz_2768_ = int_reg_array_7_34_real;
      end
      6'b100011 : begin
        _zz_2767_ = int_reg_array_7_35_imag;
        _zz_2768_ = int_reg_array_7_35_real;
      end
      6'b100100 : begin
        _zz_2767_ = int_reg_array_7_36_imag;
        _zz_2768_ = int_reg_array_7_36_real;
      end
      6'b100101 : begin
        _zz_2767_ = int_reg_array_7_37_imag;
        _zz_2768_ = int_reg_array_7_37_real;
      end
      6'b100110 : begin
        _zz_2767_ = int_reg_array_7_38_imag;
        _zz_2768_ = int_reg_array_7_38_real;
      end
      6'b100111 : begin
        _zz_2767_ = int_reg_array_7_39_imag;
        _zz_2768_ = int_reg_array_7_39_real;
      end
      6'b101000 : begin
        _zz_2767_ = int_reg_array_7_40_imag;
        _zz_2768_ = int_reg_array_7_40_real;
      end
      6'b101001 : begin
        _zz_2767_ = int_reg_array_7_41_imag;
        _zz_2768_ = int_reg_array_7_41_real;
      end
      6'b101010 : begin
        _zz_2767_ = int_reg_array_7_42_imag;
        _zz_2768_ = int_reg_array_7_42_real;
      end
      6'b101011 : begin
        _zz_2767_ = int_reg_array_7_43_imag;
        _zz_2768_ = int_reg_array_7_43_real;
      end
      6'b101100 : begin
        _zz_2767_ = int_reg_array_7_44_imag;
        _zz_2768_ = int_reg_array_7_44_real;
      end
      6'b101101 : begin
        _zz_2767_ = int_reg_array_7_45_imag;
        _zz_2768_ = int_reg_array_7_45_real;
      end
      6'b101110 : begin
        _zz_2767_ = int_reg_array_7_46_imag;
        _zz_2768_ = int_reg_array_7_46_real;
      end
      6'b101111 : begin
        _zz_2767_ = int_reg_array_7_47_imag;
        _zz_2768_ = int_reg_array_7_47_real;
      end
      6'b110000 : begin
        _zz_2767_ = int_reg_array_7_48_imag;
        _zz_2768_ = int_reg_array_7_48_real;
      end
      default : begin
        _zz_2767_ = int_reg_array_7_49_imag;
        _zz_2768_ = int_reg_array_7_49_real;
      end
    endcase
  end

  always @(*) begin
    case(_zz_442_)
      6'b000000 : begin
        _zz_2769_ = int_reg_array_8_0_imag;
        _zz_2770_ = int_reg_array_8_0_real;
      end
      6'b000001 : begin
        _zz_2769_ = int_reg_array_8_1_imag;
        _zz_2770_ = int_reg_array_8_1_real;
      end
      6'b000010 : begin
        _zz_2769_ = int_reg_array_8_2_imag;
        _zz_2770_ = int_reg_array_8_2_real;
      end
      6'b000011 : begin
        _zz_2769_ = int_reg_array_8_3_imag;
        _zz_2770_ = int_reg_array_8_3_real;
      end
      6'b000100 : begin
        _zz_2769_ = int_reg_array_8_4_imag;
        _zz_2770_ = int_reg_array_8_4_real;
      end
      6'b000101 : begin
        _zz_2769_ = int_reg_array_8_5_imag;
        _zz_2770_ = int_reg_array_8_5_real;
      end
      6'b000110 : begin
        _zz_2769_ = int_reg_array_8_6_imag;
        _zz_2770_ = int_reg_array_8_6_real;
      end
      6'b000111 : begin
        _zz_2769_ = int_reg_array_8_7_imag;
        _zz_2770_ = int_reg_array_8_7_real;
      end
      6'b001000 : begin
        _zz_2769_ = int_reg_array_8_8_imag;
        _zz_2770_ = int_reg_array_8_8_real;
      end
      6'b001001 : begin
        _zz_2769_ = int_reg_array_8_9_imag;
        _zz_2770_ = int_reg_array_8_9_real;
      end
      6'b001010 : begin
        _zz_2769_ = int_reg_array_8_10_imag;
        _zz_2770_ = int_reg_array_8_10_real;
      end
      6'b001011 : begin
        _zz_2769_ = int_reg_array_8_11_imag;
        _zz_2770_ = int_reg_array_8_11_real;
      end
      6'b001100 : begin
        _zz_2769_ = int_reg_array_8_12_imag;
        _zz_2770_ = int_reg_array_8_12_real;
      end
      6'b001101 : begin
        _zz_2769_ = int_reg_array_8_13_imag;
        _zz_2770_ = int_reg_array_8_13_real;
      end
      6'b001110 : begin
        _zz_2769_ = int_reg_array_8_14_imag;
        _zz_2770_ = int_reg_array_8_14_real;
      end
      6'b001111 : begin
        _zz_2769_ = int_reg_array_8_15_imag;
        _zz_2770_ = int_reg_array_8_15_real;
      end
      6'b010000 : begin
        _zz_2769_ = int_reg_array_8_16_imag;
        _zz_2770_ = int_reg_array_8_16_real;
      end
      6'b010001 : begin
        _zz_2769_ = int_reg_array_8_17_imag;
        _zz_2770_ = int_reg_array_8_17_real;
      end
      6'b010010 : begin
        _zz_2769_ = int_reg_array_8_18_imag;
        _zz_2770_ = int_reg_array_8_18_real;
      end
      6'b010011 : begin
        _zz_2769_ = int_reg_array_8_19_imag;
        _zz_2770_ = int_reg_array_8_19_real;
      end
      6'b010100 : begin
        _zz_2769_ = int_reg_array_8_20_imag;
        _zz_2770_ = int_reg_array_8_20_real;
      end
      6'b010101 : begin
        _zz_2769_ = int_reg_array_8_21_imag;
        _zz_2770_ = int_reg_array_8_21_real;
      end
      6'b010110 : begin
        _zz_2769_ = int_reg_array_8_22_imag;
        _zz_2770_ = int_reg_array_8_22_real;
      end
      6'b010111 : begin
        _zz_2769_ = int_reg_array_8_23_imag;
        _zz_2770_ = int_reg_array_8_23_real;
      end
      6'b011000 : begin
        _zz_2769_ = int_reg_array_8_24_imag;
        _zz_2770_ = int_reg_array_8_24_real;
      end
      6'b011001 : begin
        _zz_2769_ = int_reg_array_8_25_imag;
        _zz_2770_ = int_reg_array_8_25_real;
      end
      6'b011010 : begin
        _zz_2769_ = int_reg_array_8_26_imag;
        _zz_2770_ = int_reg_array_8_26_real;
      end
      6'b011011 : begin
        _zz_2769_ = int_reg_array_8_27_imag;
        _zz_2770_ = int_reg_array_8_27_real;
      end
      6'b011100 : begin
        _zz_2769_ = int_reg_array_8_28_imag;
        _zz_2770_ = int_reg_array_8_28_real;
      end
      6'b011101 : begin
        _zz_2769_ = int_reg_array_8_29_imag;
        _zz_2770_ = int_reg_array_8_29_real;
      end
      6'b011110 : begin
        _zz_2769_ = int_reg_array_8_30_imag;
        _zz_2770_ = int_reg_array_8_30_real;
      end
      6'b011111 : begin
        _zz_2769_ = int_reg_array_8_31_imag;
        _zz_2770_ = int_reg_array_8_31_real;
      end
      6'b100000 : begin
        _zz_2769_ = int_reg_array_8_32_imag;
        _zz_2770_ = int_reg_array_8_32_real;
      end
      6'b100001 : begin
        _zz_2769_ = int_reg_array_8_33_imag;
        _zz_2770_ = int_reg_array_8_33_real;
      end
      6'b100010 : begin
        _zz_2769_ = int_reg_array_8_34_imag;
        _zz_2770_ = int_reg_array_8_34_real;
      end
      6'b100011 : begin
        _zz_2769_ = int_reg_array_8_35_imag;
        _zz_2770_ = int_reg_array_8_35_real;
      end
      6'b100100 : begin
        _zz_2769_ = int_reg_array_8_36_imag;
        _zz_2770_ = int_reg_array_8_36_real;
      end
      6'b100101 : begin
        _zz_2769_ = int_reg_array_8_37_imag;
        _zz_2770_ = int_reg_array_8_37_real;
      end
      6'b100110 : begin
        _zz_2769_ = int_reg_array_8_38_imag;
        _zz_2770_ = int_reg_array_8_38_real;
      end
      6'b100111 : begin
        _zz_2769_ = int_reg_array_8_39_imag;
        _zz_2770_ = int_reg_array_8_39_real;
      end
      6'b101000 : begin
        _zz_2769_ = int_reg_array_8_40_imag;
        _zz_2770_ = int_reg_array_8_40_real;
      end
      6'b101001 : begin
        _zz_2769_ = int_reg_array_8_41_imag;
        _zz_2770_ = int_reg_array_8_41_real;
      end
      6'b101010 : begin
        _zz_2769_ = int_reg_array_8_42_imag;
        _zz_2770_ = int_reg_array_8_42_real;
      end
      6'b101011 : begin
        _zz_2769_ = int_reg_array_8_43_imag;
        _zz_2770_ = int_reg_array_8_43_real;
      end
      6'b101100 : begin
        _zz_2769_ = int_reg_array_8_44_imag;
        _zz_2770_ = int_reg_array_8_44_real;
      end
      6'b101101 : begin
        _zz_2769_ = int_reg_array_8_45_imag;
        _zz_2770_ = int_reg_array_8_45_real;
      end
      6'b101110 : begin
        _zz_2769_ = int_reg_array_8_46_imag;
        _zz_2770_ = int_reg_array_8_46_real;
      end
      6'b101111 : begin
        _zz_2769_ = int_reg_array_8_47_imag;
        _zz_2770_ = int_reg_array_8_47_real;
      end
      6'b110000 : begin
        _zz_2769_ = int_reg_array_8_48_imag;
        _zz_2770_ = int_reg_array_8_48_real;
      end
      default : begin
        _zz_2769_ = int_reg_array_8_49_imag;
        _zz_2770_ = int_reg_array_8_49_real;
      end
    endcase
  end

  always @(*) begin
    case(_zz_497_)
      6'b000000 : begin
        _zz_2771_ = int_reg_array_9_0_imag;
        _zz_2772_ = int_reg_array_9_0_real;
      end
      6'b000001 : begin
        _zz_2771_ = int_reg_array_9_1_imag;
        _zz_2772_ = int_reg_array_9_1_real;
      end
      6'b000010 : begin
        _zz_2771_ = int_reg_array_9_2_imag;
        _zz_2772_ = int_reg_array_9_2_real;
      end
      6'b000011 : begin
        _zz_2771_ = int_reg_array_9_3_imag;
        _zz_2772_ = int_reg_array_9_3_real;
      end
      6'b000100 : begin
        _zz_2771_ = int_reg_array_9_4_imag;
        _zz_2772_ = int_reg_array_9_4_real;
      end
      6'b000101 : begin
        _zz_2771_ = int_reg_array_9_5_imag;
        _zz_2772_ = int_reg_array_9_5_real;
      end
      6'b000110 : begin
        _zz_2771_ = int_reg_array_9_6_imag;
        _zz_2772_ = int_reg_array_9_6_real;
      end
      6'b000111 : begin
        _zz_2771_ = int_reg_array_9_7_imag;
        _zz_2772_ = int_reg_array_9_7_real;
      end
      6'b001000 : begin
        _zz_2771_ = int_reg_array_9_8_imag;
        _zz_2772_ = int_reg_array_9_8_real;
      end
      6'b001001 : begin
        _zz_2771_ = int_reg_array_9_9_imag;
        _zz_2772_ = int_reg_array_9_9_real;
      end
      6'b001010 : begin
        _zz_2771_ = int_reg_array_9_10_imag;
        _zz_2772_ = int_reg_array_9_10_real;
      end
      6'b001011 : begin
        _zz_2771_ = int_reg_array_9_11_imag;
        _zz_2772_ = int_reg_array_9_11_real;
      end
      6'b001100 : begin
        _zz_2771_ = int_reg_array_9_12_imag;
        _zz_2772_ = int_reg_array_9_12_real;
      end
      6'b001101 : begin
        _zz_2771_ = int_reg_array_9_13_imag;
        _zz_2772_ = int_reg_array_9_13_real;
      end
      6'b001110 : begin
        _zz_2771_ = int_reg_array_9_14_imag;
        _zz_2772_ = int_reg_array_9_14_real;
      end
      6'b001111 : begin
        _zz_2771_ = int_reg_array_9_15_imag;
        _zz_2772_ = int_reg_array_9_15_real;
      end
      6'b010000 : begin
        _zz_2771_ = int_reg_array_9_16_imag;
        _zz_2772_ = int_reg_array_9_16_real;
      end
      6'b010001 : begin
        _zz_2771_ = int_reg_array_9_17_imag;
        _zz_2772_ = int_reg_array_9_17_real;
      end
      6'b010010 : begin
        _zz_2771_ = int_reg_array_9_18_imag;
        _zz_2772_ = int_reg_array_9_18_real;
      end
      6'b010011 : begin
        _zz_2771_ = int_reg_array_9_19_imag;
        _zz_2772_ = int_reg_array_9_19_real;
      end
      6'b010100 : begin
        _zz_2771_ = int_reg_array_9_20_imag;
        _zz_2772_ = int_reg_array_9_20_real;
      end
      6'b010101 : begin
        _zz_2771_ = int_reg_array_9_21_imag;
        _zz_2772_ = int_reg_array_9_21_real;
      end
      6'b010110 : begin
        _zz_2771_ = int_reg_array_9_22_imag;
        _zz_2772_ = int_reg_array_9_22_real;
      end
      6'b010111 : begin
        _zz_2771_ = int_reg_array_9_23_imag;
        _zz_2772_ = int_reg_array_9_23_real;
      end
      6'b011000 : begin
        _zz_2771_ = int_reg_array_9_24_imag;
        _zz_2772_ = int_reg_array_9_24_real;
      end
      6'b011001 : begin
        _zz_2771_ = int_reg_array_9_25_imag;
        _zz_2772_ = int_reg_array_9_25_real;
      end
      6'b011010 : begin
        _zz_2771_ = int_reg_array_9_26_imag;
        _zz_2772_ = int_reg_array_9_26_real;
      end
      6'b011011 : begin
        _zz_2771_ = int_reg_array_9_27_imag;
        _zz_2772_ = int_reg_array_9_27_real;
      end
      6'b011100 : begin
        _zz_2771_ = int_reg_array_9_28_imag;
        _zz_2772_ = int_reg_array_9_28_real;
      end
      6'b011101 : begin
        _zz_2771_ = int_reg_array_9_29_imag;
        _zz_2772_ = int_reg_array_9_29_real;
      end
      6'b011110 : begin
        _zz_2771_ = int_reg_array_9_30_imag;
        _zz_2772_ = int_reg_array_9_30_real;
      end
      6'b011111 : begin
        _zz_2771_ = int_reg_array_9_31_imag;
        _zz_2772_ = int_reg_array_9_31_real;
      end
      6'b100000 : begin
        _zz_2771_ = int_reg_array_9_32_imag;
        _zz_2772_ = int_reg_array_9_32_real;
      end
      6'b100001 : begin
        _zz_2771_ = int_reg_array_9_33_imag;
        _zz_2772_ = int_reg_array_9_33_real;
      end
      6'b100010 : begin
        _zz_2771_ = int_reg_array_9_34_imag;
        _zz_2772_ = int_reg_array_9_34_real;
      end
      6'b100011 : begin
        _zz_2771_ = int_reg_array_9_35_imag;
        _zz_2772_ = int_reg_array_9_35_real;
      end
      6'b100100 : begin
        _zz_2771_ = int_reg_array_9_36_imag;
        _zz_2772_ = int_reg_array_9_36_real;
      end
      6'b100101 : begin
        _zz_2771_ = int_reg_array_9_37_imag;
        _zz_2772_ = int_reg_array_9_37_real;
      end
      6'b100110 : begin
        _zz_2771_ = int_reg_array_9_38_imag;
        _zz_2772_ = int_reg_array_9_38_real;
      end
      6'b100111 : begin
        _zz_2771_ = int_reg_array_9_39_imag;
        _zz_2772_ = int_reg_array_9_39_real;
      end
      6'b101000 : begin
        _zz_2771_ = int_reg_array_9_40_imag;
        _zz_2772_ = int_reg_array_9_40_real;
      end
      6'b101001 : begin
        _zz_2771_ = int_reg_array_9_41_imag;
        _zz_2772_ = int_reg_array_9_41_real;
      end
      6'b101010 : begin
        _zz_2771_ = int_reg_array_9_42_imag;
        _zz_2772_ = int_reg_array_9_42_real;
      end
      6'b101011 : begin
        _zz_2771_ = int_reg_array_9_43_imag;
        _zz_2772_ = int_reg_array_9_43_real;
      end
      6'b101100 : begin
        _zz_2771_ = int_reg_array_9_44_imag;
        _zz_2772_ = int_reg_array_9_44_real;
      end
      6'b101101 : begin
        _zz_2771_ = int_reg_array_9_45_imag;
        _zz_2772_ = int_reg_array_9_45_real;
      end
      6'b101110 : begin
        _zz_2771_ = int_reg_array_9_46_imag;
        _zz_2772_ = int_reg_array_9_46_real;
      end
      6'b101111 : begin
        _zz_2771_ = int_reg_array_9_47_imag;
        _zz_2772_ = int_reg_array_9_47_real;
      end
      6'b110000 : begin
        _zz_2771_ = int_reg_array_9_48_imag;
        _zz_2772_ = int_reg_array_9_48_real;
      end
      default : begin
        _zz_2771_ = int_reg_array_9_49_imag;
        _zz_2772_ = int_reg_array_9_49_real;
      end
    endcase
  end

  always @(*) begin
    case(_zz_552_)
      6'b000000 : begin
        _zz_2773_ = int_reg_array_10_0_imag;
        _zz_2774_ = int_reg_array_10_0_real;
      end
      6'b000001 : begin
        _zz_2773_ = int_reg_array_10_1_imag;
        _zz_2774_ = int_reg_array_10_1_real;
      end
      6'b000010 : begin
        _zz_2773_ = int_reg_array_10_2_imag;
        _zz_2774_ = int_reg_array_10_2_real;
      end
      6'b000011 : begin
        _zz_2773_ = int_reg_array_10_3_imag;
        _zz_2774_ = int_reg_array_10_3_real;
      end
      6'b000100 : begin
        _zz_2773_ = int_reg_array_10_4_imag;
        _zz_2774_ = int_reg_array_10_4_real;
      end
      6'b000101 : begin
        _zz_2773_ = int_reg_array_10_5_imag;
        _zz_2774_ = int_reg_array_10_5_real;
      end
      6'b000110 : begin
        _zz_2773_ = int_reg_array_10_6_imag;
        _zz_2774_ = int_reg_array_10_6_real;
      end
      6'b000111 : begin
        _zz_2773_ = int_reg_array_10_7_imag;
        _zz_2774_ = int_reg_array_10_7_real;
      end
      6'b001000 : begin
        _zz_2773_ = int_reg_array_10_8_imag;
        _zz_2774_ = int_reg_array_10_8_real;
      end
      6'b001001 : begin
        _zz_2773_ = int_reg_array_10_9_imag;
        _zz_2774_ = int_reg_array_10_9_real;
      end
      6'b001010 : begin
        _zz_2773_ = int_reg_array_10_10_imag;
        _zz_2774_ = int_reg_array_10_10_real;
      end
      6'b001011 : begin
        _zz_2773_ = int_reg_array_10_11_imag;
        _zz_2774_ = int_reg_array_10_11_real;
      end
      6'b001100 : begin
        _zz_2773_ = int_reg_array_10_12_imag;
        _zz_2774_ = int_reg_array_10_12_real;
      end
      6'b001101 : begin
        _zz_2773_ = int_reg_array_10_13_imag;
        _zz_2774_ = int_reg_array_10_13_real;
      end
      6'b001110 : begin
        _zz_2773_ = int_reg_array_10_14_imag;
        _zz_2774_ = int_reg_array_10_14_real;
      end
      6'b001111 : begin
        _zz_2773_ = int_reg_array_10_15_imag;
        _zz_2774_ = int_reg_array_10_15_real;
      end
      6'b010000 : begin
        _zz_2773_ = int_reg_array_10_16_imag;
        _zz_2774_ = int_reg_array_10_16_real;
      end
      6'b010001 : begin
        _zz_2773_ = int_reg_array_10_17_imag;
        _zz_2774_ = int_reg_array_10_17_real;
      end
      6'b010010 : begin
        _zz_2773_ = int_reg_array_10_18_imag;
        _zz_2774_ = int_reg_array_10_18_real;
      end
      6'b010011 : begin
        _zz_2773_ = int_reg_array_10_19_imag;
        _zz_2774_ = int_reg_array_10_19_real;
      end
      6'b010100 : begin
        _zz_2773_ = int_reg_array_10_20_imag;
        _zz_2774_ = int_reg_array_10_20_real;
      end
      6'b010101 : begin
        _zz_2773_ = int_reg_array_10_21_imag;
        _zz_2774_ = int_reg_array_10_21_real;
      end
      6'b010110 : begin
        _zz_2773_ = int_reg_array_10_22_imag;
        _zz_2774_ = int_reg_array_10_22_real;
      end
      6'b010111 : begin
        _zz_2773_ = int_reg_array_10_23_imag;
        _zz_2774_ = int_reg_array_10_23_real;
      end
      6'b011000 : begin
        _zz_2773_ = int_reg_array_10_24_imag;
        _zz_2774_ = int_reg_array_10_24_real;
      end
      6'b011001 : begin
        _zz_2773_ = int_reg_array_10_25_imag;
        _zz_2774_ = int_reg_array_10_25_real;
      end
      6'b011010 : begin
        _zz_2773_ = int_reg_array_10_26_imag;
        _zz_2774_ = int_reg_array_10_26_real;
      end
      6'b011011 : begin
        _zz_2773_ = int_reg_array_10_27_imag;
        _zz_2774_ = int_reg_array_10_27_real;
      end
      6'b011100 : begin
        _zz_2773_ = int_reg_array_10_28_imag;
        _zz_2774_ = int_reg_array_10_28_real;
      end
      6'b011101 : begin
        _zz_2773_ = int_reg_array_10_29_imag;
        _zz_2774_ = int_reg_array_10_29_real;
      end
      6'b011110 : begin
        _zz_2773_ = int_reg_array_10_30_imag;
        _zz_2774_ = int_reg_array_10_30_real;
      end
      6'b011111 : begin
        _zz_2773_ = int_reg_array_10_31_imag;
        _zz_2774_ = int_reg_array_10_31_real;
      end
      6'b100000 : begin
        _zz_2773_ = int_reg_array_10_32_imag;
        _zz_2774_ = int_reg_array_10_32_real;
      end
      6'b100001 : begin
        _zz_2773_ = int_reg_array_10_33_imag;
        _zz_2774_ = int_reg_array_10_33_real;
      end
      6'b100010 : begin
        _zz_2773_ = int_reg_array_10_34_imag;
        _zz_2774_ = int_reg_array_10_34_real;
      end
      6'b100011 : begin
        _zz_2773_ = int_reg_array_10_35_imag;
        _zz_2774_ = int_reg_array_10_35_real;
      end
      6'b100100 : begin
        _zz_2773_ = int_reg_array_10_36_imag;
        _zz_2774_ = int_reg_array_10_36_real;
      end
      6'b100101 : begin
        _zz_2773_ = int_reg_array_10_37_imag;
        _zz_2774_ = int_reg_array_10_37_real;
      end
      6'b100110 : begin
        _zz_2773_ = int_reg_array_10_38_imag;
        _zz_2774_ = int_reg_array_10_38_real;
      end
      6'b100111 : begin
        _zz_2773_ = int_reg_array_10_39_imag;
        _zz_2774_ = int_reg_array_10_39_real;
      end
      6'b101000 : begin
        _zz_2773_ = int_reg_array_10_40_imag;
        _zz_2774_ = int_reg_array_10_40_real;
      end
      6'b101001 : begin
        _zz_2773_ = int_reg_array_10_41_imag;
        _zz_2774_ = int_reg_array_10_41_real;
      end
      6'b101010 : begin
        _zz_2773_ = int_reg_array_10_42_imag;
        _zz_2774_ = int_reg_array_10_42_real;
      end
      6'b101011 : begin
        _zz_2773_ = int_reg_array_10_43_imag;
        _zz_2774_ = int_reg_array_10_43_real;
      end
      6'b101100 : begin
        _zz_2773_ = int_reg_array_10_44_imag;
        _zz_2774_ = int_reg_array_10_44_real;
      end
      6'b101101 : begin
        _zz_2773_ = int_reg_array_10_45_imag;
        _zz_2774_ = int_reg_array_10_45_real;
      end
      6'b101110 : begin
        _zz_2773_ = int_reg_array_10_46_imag;
        _zz_2774_ = int_reg_array_10_46_real;
      end
      6'b101111 : begin
        _zz_2773_ = int_reg_array_10_47_imag;
        _zz_2774_ = int_reg_array_10_47_real;
      end
      6'b110000 : begin
        _zz_2773_ = int_reg_array_10_48_imag;
        _zz_2774_ = int_reg_array_10_48_real;
      end
      default : begin
        _zz_2773_ = int_reg_array_10_49_imag;
        _zz_2774_ = int_reg_array_10_49_real;
      end
    endcase
  end

  always @(*) begin
    case(_zz_607_)
      6'b000000 : begin
        _zz_2775_ = int_reg_array_11_0_imag;
        _zz_2776_ = int_reg_array_11_0_real;
      end
      6'b000001 : begin
        _zz_2775_ = int_reg_array_11_1_imag;
        _zz_2776_ = int_reg_array_11_1_real;
      end
      6'b000010 : begin
        _zz_2775_ = int_reg_array_11_2_imag;
        _zz_2776_ = int_reg_array_11_2_real;
      end
      6'b000011 : begin
        _zz_2775_ = int_reg_array_11_3_imag;
        _zz_2776_ = int_reg_array_11_3_real;
      end
      6'b000100 : begin
        _zz_2775_ = int_reg_array_11_4_imag;
        _zz_2776_ = int_reg_array_11_4_real;
      end
      6'b000101 : begin
        _zz_2775_ = int_reg_array_11_5_imag;
        _zz_2776_ = int_reg_array_11_5_real;
      end
      6'b000110 : begin
        _zz_2775_ = int_reg_array_11_6_imag;
        _zz_2776_ = int_reg_array_11_6_real;
      end
      6'b000111 : begin
        _zz_2775_ = int_reg_array_11_7_imag;
        _zz_2776_ = int_reg_array_11_7_real;
      end
      6'b001000 : begin
        _zz_2775_ = int_reg_array_11_8_imag;
        _zz_2776_ = int_reg_array_11_8_real;
      end
      6'b001001 : begin
        _zz_2775_ = int_reg_array_11_9_imag;
        _zz_2776_ = int_reg_array_11_9_real;
      end
      6'b001010 : begin
        _zz_2775_ = int_reg_array_11_10_imag;
        _zz_2776_ = int_reg_array_11_10_real;
      end
      6'b001011 : begin
        _zz_2775_ = int_reg_array_11_11_imag;
        _zz_2776_ = int_reg_array_11_11_real;
      end
      6'b001100 : begin
        _zz_2775_ = int_reg_array_11_12_imag;
        _zz_2776_ = int_reg_array_11_12_real;
      end
      6'b001101 : begin
        _zz_2775_ = int_reg_array_11_13_imag;
        _zz_2776_ = int_reg_array_11_13_real;
      end
      6'b001110 : begin
        _zz_2775_ = int_reg_array_11_14_imag;
        _zz_2776_ = int_reg_array_11_14_real;
      end
      6'b001111 : begin
        _zz_2775_ = int_reg_array_11_15_imag;
        _zz_2776_ = int_reg_array_11_15_real;
      end
      6'b010000 : begin
        _zz_2775_ = int_reg_array_11_16_imag;
        _zz_2776_ = int_reg_array_11_16_real;
      end
      6'b010001 : begin
        _zz_2775_ = int_reg_array_11_17_imag;
        _zz_2776_ = int_reg_array_11_17_real;
      end
      6'b010010 : begin
        _zz_2775_ = int_reg_array_11_18_imag;
        _zz_2776_ = int_reg_array_11_18_real;
      end
      6'b010011 : begin
        _zz_2775_ = int_reg_array_11_19_imag;
        _zz_2776_ = int_reg_array_11_19_real;
      end
      6'b010100 : begin
        _zz_2775_ = int_reg_array_11_20_imag;
        _zz_2776_ = int_reg_array_11_20_real;
      end
      6'b010101 : begin
        _zz_2775_ = int_reg_array_11_21_imag;
        _zz_2776_ = int_reg_array_11_21_real;
      end
      6'b010110 : begin
        _zz_2775_ = int_reg_array_11_22_imag;
        _zz_2776_ = int_reg_array_11_22_real;
      end
      6'b010111 : begin
        _zz_2775_ = int_reg_array_11_23_imag;
        _zz_2776_ = int_reg_array_11_23_real;
      end
      6'b011000 : begin
        _zz_2775_ = int_reg_array_11_24_imag;
        _zz_2776_ = int_reg_array_11_24_real;
      end
      6'b011001 : begin
        _zz_2775_ = int_reg_array_11_25_imag;
        _zz_2776_ = int_reg_array_11_25_real;
      end
      6'b011010 : begin
        _zz_2775_ = int_reg_array_11_26_imag;
        _zz_2776_ = int_reg_array_11_26_real;
      end
      6'b011011 : begin
        _zz_2775_ = int_reg_array_11_27_imag;
        _zz_2776_ = int_reg_array_11_27_real;
      end
      6'b011100 : begin
        _zz_2775_ = int_reg_array_11_28_imag;
        _zz_2776_ = int_reg_array_11_28_real;
      end
      6'b011101 : begin
        _zz_2775_ = int_reg_array_11_29_imag;
        _zz_2776_ = int_reg_array_11_29_real;
      end
      6'b011110 : begin
        _zz_2775_ = int_reg_array_11_30_imag;
        _zz_2776_ = int_reg_array_11_30_real;
      end
      6'b011111 : begin
        _zz_2775_ = int_reg_array_11_31_imag;
        _zz_2776_ = int_reg_array_11_31_real;
      end
      6'b100000 : begin
        _zz_2775_ = int_reg_array_11_32_imag;
        _zz_2776_ = int_reg_array_11_32_real;
      end
      6'b100001 : begin
        _zz_2775_ = int_reg_array_11_33_imag;
        _zz_2776_ = int_reg_array_11_33_real;
      end
      6'b100010 : begin
        _zz_2775_ = int_reg_array_11_34_imag;
        _zz_2776_ = int_reg_array_11_34_real;
      end
      6'b100011 : begin
        _zz_2775_ = int_reg_array_11_35_imag;
        _zz_2776_ = int_reg_array_11_35_real;
      end
      6'b100100 : begin
        _zz_2775_ = int_reg_array_11_36_imag;
        _zz_2776_ = int_reg_array_11_36_real;
      end
      6'b100101 : begin
        _zz_2775_ = int_reg_array_11_37_imag;
        _zz_2776_ = int_reg_array_11_37_real;
      end
      6'b100110 : begin
        _zz_2775_ = int_reg_array_11_38_imag;
        _zz_2776_ = int_reg_array_11_38_real;
      end
      6'b100111 : begin
        _zz_2775_ = int_reg_array_11_39_imag;
        _zz_2776_ = int_reg_array_11_39_real;
      end
      6'b101000 : begin
        _zz_2775_ = int_reg_array_11_40_imag;
        _zz_2776_ = int_reg_array_11_40_real;
      end
      6'b101001 : begin
        _zz_2775_ = int_reg_array_11_41_imag;
        _zz_2776_ = int_reg_array_11_41_real;
      end
      6'b101010 : begin
        _zz_2775_ = int_reg_array_11_42_imag;
        _zz_2776_ = int_reg_array_11_42_real;
      end
      6'b101011 : begin
        _zz_2775_ = int_reg_array_11_43_imag;
        _zz_2776_ = int_reg_array_11_43_real;
      end
      6'b101100 : begin
        _zz_2775_ = int_reg_array_11_44_imag;
        _zz_2776_ = int_reg_array_11_44_real;
      end
      6'b101101 : begin
        _zz_2775_ = int_reg_array_11_45_imag;
        _zz_2776_ = int_reg_array_11_45_real;
      end
      6'b101110 : begin
        _zz_2775_ = int_reg_array_11_46_imag;
        _zz_2776_ = int_reg_array_11_46_real;
      end
      6'b101111 : begin
        _zz_2775_ = int_reg_array_11_47_imag;
        _zz_2776_ = int_reg_array_11_47_real;
      end
      6'b110000 : begin
        _zz_2775_ = int_reg_array_11_48_imag;
        _zz_2776_ = int_reg_array_11_48_real;
      end
      default : begin
        _zz_2775_ = int_reg_array_11_49_imag;
        _zz_2776_ = int_reg_array_11_49_real;
      end
    endcase
  end

  always @(*) begin
    case(_zz_662_)
      6'b000000 : begin
        _zz_2777_ = int_reg_array_12_0_imag;
        _zz_2778_ = int_reg_array_12_0_real;
      end
      6'b000001 : begin
        _zz_2777_ = int_reg_array_12_1_imag;
        _zz_2778_ = int_reg_array_12_1_real;
      end
      6'b000010 : begin
        _zz_2777_ = int_reg_array_12_2_imag;
        _zz_2778_ = int_reg_array_12_2_real;
      end
      6'b000011 : begin
        _zz_2777_ = int_reg_array_12_3_imag;
        _zz_2778_ = int_reg_array_12_3_real;
      end
      6'b000100 : begin
        _zz_2777_ = int_reg_array_12_4_imag;
        _zz_2778_ = int_reg_array_12_4_real;
      end
      6'b000101 : begin
        _zz_2777_ = int_reg_array_12_5_imag;
        _zz_2778_ = int_reg_array_12_5_real;
      end
      6'b000110 : begin
        _zz_2777_ = int_reg_array_12_6_imag;
        _zz_2778_ = int_reg_array_12_6_real;
      end
      6'b000111 : begin
        _zz_2777_ = int_reg_array_12_7_imag;
        _zz_2778_ = int_reg_array_12_7_real;
      end
      6'b001000 : begin
        _zz_2777_ = int_reg_array_12_8_imag;
        _zz_2778_ = int_reg_array_12_8_real;
      end
      6'b001001 : begin
        _zz_2777_ = int_reg_array_12_9_imag;
        _zz_2778_ = int_reg_array_12_9_real;
      end
      6'b001010 : begin
        _zz_2777_ = int_reg_array_12_10_imag;
        _zz_2778_ = int_reg_array_12_10_real;
      end
      6'b001011 : begin
        _zz_2777_ = int_reg_array_12_11_imag;
        _zz_2778_ = int_reg_array_12_11_real;
      end
      6'b001100 : begin
        _zz_2777_ = int_reg_array_12_12_imag;
        _zz_2778_ = int_reg_array_12_12_real;
      end
      6'b001101 : begin
        _zz_2777_ = int_reg_array_12_13_imag;
        _zz_2778_ = int_reg_array_12_13_real;
      end
      6'b001110 : begin
        _zz_2777_ = int_reg_array_12_14_imag;
        _zz_2778_ = int_reg_array_12_14_real;
      end
      6'b001111 : begin
        _zz_2777_ = int_reg_array_12_15_imag;
        _zz_2778_ = int_reg_array_12_15_real;
      end
      6'b010000 : begin
        _zz_2777_ = int_reg_array_12_16_imag;
        _zz_2778_ = int_reg_array_12_16_real;
      end
      6'b010001 : begin
        _zz_2777_ = int_reg_array_12_17_imag;
        _zz_2778_ = int_reg_array_12_17_real;
      end
      6'b010010 : begin
        _zz_2777_ = int_reg_array_12_18_imag;
        _zz_2778_ = int_reg_array_12_18_real;
      end
      6'b010011 : begin
        _zz_2777_ = int_reg_array_12_19_imag;
        _zz_2778_ = int_reg_array_12_19_real;
      end
      6'b010100 : begin
        _zz_2777_ = int_reg_array_12_20_imag;
        _zz_2778_ = int_reg_array_12_20_real;
      end
      6'b010101 : begin
        _zz_2777_ = int_reg_array_12_21_imag;
        _zz_2778_ = int_reg_array_12_21_real;
      end
      6'b010110 : begin
        _zz_2777_ = int_reg_array_12_22_imag;
        _zz_2778_ = int_reg_array_12_22_real;
      end
      6'b010111 : begin
        _zz_2777_ = int_reg_array_12_23_imag;
        _zz_2778_ = int_reg_array_12_23_real;
      end
      6'b011000 : begin
        _zz_2777_ = int_reg_array_12_24_imag;
        _zz_2778_ = int_reg_array_12_24_real;
      end
      6'b011001 : begin
        _zz_2777_ = int_reg_array_12_25_imag;
        _zz_2778_ = int_reg_array_12_25_real;
      end
      6'b011010 : begin
        _zz_2777_ = int_reg_array_12_26_imag;
        _zz_2778_ = int_reg_array_12_26_real;
      end
      6'b011011 : begin
        _zz_2777_ = int_reg_array_12_27_imag;
        _zz_2778_ = int_reg_array_12_27_real;
      end
      6'b011100 : begin
        _zz_2777_ = int_reg_array_12_28_imag;
        _zz_2778_ = int_reg_array_12_28_real;
      end
      6'b011101 : begin
        _zz_2777_ = int_reg_array_12_29_imag;
        _zz_2778_ = int_reg_array_12_29_real;
      end
      6'b011110 : begin
        _zz_2777_ = int_reg_array_12_30_imag;
        _zz_2778_ = int_reg_array_12_30_real;
      end
      6'b011111 : begin
        _zz_2777_ = int_reg_array_12_31_imag;
        _zz_2778_ = int_reg_array_12_31_real;
      end
      6'b100000 : begin
        _zz_2777_ = int_reg_array_12_32_imag;
        _zz_2778_ = int_reg_array_12_32_real;
      end
      6'b100001 : begin
        _zz_2777_ = int_reg_array_12_33_imag;
        _zz_2778_ = int_reg_array_12_33_real;
      end
      6'b100010 : begin
        _zz_2777_ = int_reg_array_12_34_imag;
        _zz_2778_ = int_reg_array_12_34_real;
      end
      6'b100011 : begin
        _zz_2777_ = int_reg_array_12_35_imag;
        _zz_2778_ = int_reg_array_12_35_real;
      end
      6'b100100 : begin
        _zz_2777_ = int_reg_array_12_36_imag;
        _zz_2778_ = int_reg_array_12_36_real;
      end
      6'b100101 : begin
        _zz_2777_ = int_reg_array_12_37_imag;
        _zz_2778_ = int_reg_array_12_37_real;
      end
      6'b100110 : begin
        _zz_2777_ = int_reg_array_12_38_imag;
        _zz_2778_ = int_reg_array_12_38_real;
      end
      6'b100111 : begin
        _zz_2777_ = int_reg_array_12_39_imag;
        _zz_2778_ = int_reg_array_12_39_real;
      end
      6'b101000 : begin
        _zz_2777_ = int_reg_array_12_40_imag;
        _zz_2778_ = int_reg_array_12_40_real;
      end
      6'b101001 : begin
        _zz_2777_ = int_reg_array_12_41_imag;
        _zz_2778_ = int_reg_array_12_41_real;
      end
      6'b101010 : begin
        _zz_2777_ = int_reg_array_12_42_imag;
        _zz_2778_ = int_reg_array_12_42_real;
      end
      6'b101011 : begin
        _zz_2777_ = int_reg_array_12_43_imag;
        _zz_2778_ = int_reg_array_12_43_real;
      end
      6'b101100 : begin
        _zz_2777_ = int_reg_array_12_44_imag;
        _zz_2778_ = int_reg_array_12_44_real;
      end
      6'b101101 : begin
        _zz_2777_ = int_reg_array_12_45_imag;
        _zz_2778_ = int_reg_array_12_45_real;
      end
      6'b101110 : begin
        _zz_2777_ = int_reg_array_12_46_imag;
        _zz_2778_ = int_reg_array_12_46_real;
      end
      6'b101111 : begin
        _zz_2777_ = int_reg_array_12_47_imag;
        _zz_2778_ = int_reg_array_12_47_real;
      end
      6'b110000 : begin
        _zz_2777_ = int_reg_array_12_48_imag;
        _zz_2778_ = int_reg_array_12_48_real;
      end
      default : begin
        _zz_2777_ = int_reg_array_12_49_imag;
        _zz_2778_ = int_reg_array_12_49_real;
      end
    endcase
  end

  always @(*) begin
    case(_zz_717_)
      6'b000000 : begin
        _zz_2779_ = int_reg_array_13_0_imag;
        _zz_2780_ = int_reg_array_13_0_real;
      end
      6'b000001 : begin
        _zz_2779_ = int_reg_array_13_1_imag;
        _zz_2780_ = int_reg_array_13_1_real;
      end
      6'b000010 : begin
        _zz_2779_ = int_reg_array_13_2_imag;
        _zz_2780_ = int_reg_array_13_2_real;
      end
      6'b000011 : begin
        _zz_2779_ = int_reg_array_13_3_imag;
        _zz_2780_ = int_reg_array_13_3_real;
      end
      6'b000100 : begin
        _zz_2779_ = int_reg_array_13_4_imag;
        _zz_2780_ = int_reg_array_13_4_real;
      end
      6'b000101 : begin
        _zz_2779_ = int_reg_array_13_5_imag;
        _zz_2780_ = int_reg_array_13_5_real;
      end
      6'b000110 : begin
        _zz_2779_ = int_reg_array_13_6_imag;
        _zz_2780_ = int_reg_array_13_6_real;
      end
      6'b000111 : begin
        _zz_2779_ = int_reg_array_13_7_imag;
        _zz_2780_ = int_reg_array_13_7_real;
      end
      6'b001000 : begin
        _zz_2779_ = int_reg_array_13_8_imag;
        _zz_2780_ = int_reg_array_13_8_real;
      end
      6'b001001 : begin
        _zz_2779_ = int_reg_array_13_9_imag;
        _zz_2780_ = int_reg_array_13_9_real;
      end
      6'b001010 : begin
        _zz_2779_ = int_reg_array_13_10_imag;
        _zz_2780_ = int_reg_array_13_10_real;
      end
      6'b001011 : begin
        _zz_2779_ = int_reg_array_13_11_imag;
        _zz_2780_ = int_reg_array_13_11_real;
      end
      6'b001100 : begin
        _zz_2779_ = int_reg_array_13_12_imag;
        _zz_2780_ = int_reg_array_13_12_real;
      end
      6'b001101 : begin
        _zz_2779_ = int_reg_array_13_13_imag;
        _zz_2780_ = int_reg_array_13_13_real;
      end
      6'b001110 : begin
        _zz_2779_ = int_reg_array_13_14_imag;
        _zz_2780_ = int_reg_array_13_14_real;
      end
      6'b001111 : begin
        _zz_2779_ = int_reg_array_13_15_imag;
        _zz_2780_ = int_reg_array_13_15_real;
      end
      6'b010000 : begin
        _zz_2779_ = int_reg_array_13_16_imag;
        _zz_2780_ = int_reg_array_13_16_real;
      end
      6'b010001 : begin
        _zz_2779_ = int_reg_array_13_17_imag;
        _zz_2780_ = int_reg_array_13_17_real;
      end
      6'b010010 : begin
        _zz_2779_ = int_reg_array_13_18_imag;
        _zz_2780_ = int_reg_array_13_18_real;
      end
      6'b010011 : begin
        _zz_2779_ = int_reg_array_13_19_imag;
        _zz_2780_ = int_reg_array_13_19_real;
      end
      6'b010100 : begin
        _zz_2779_ = int_reg_array_13_20_imag;
        _zz_2780_ = int_reg_array_13_20_real;
      end
      6'b010101 : begin
        _zz_2779_ = int_reg_array_13_21_imag;
        _zz_2780_ = int_reg_array_13_21_real;
      end
      6'b010110 : begin
        _zz_2779_ = int_reg_array_13_22_imag;
        _zz_2780_ = int_reg_array_13_22_real;
      end
      6'b010111 : begin
        _zz_2779_ = int_reg_array_13_23_imag;
        _zz_2780_ = int_reg_array_13_23_real;
      end
      6'b011000 : begin
        _zz_2779_ = int_reg_array_13_24_imag;
        _zz_2780_ = int_reg_array_13_24_real;
      end
      6'b011001 : begin
        _zz_2779_ = int_reg_array_13_25_imag;
        _zz_2780_ = int_reg_array_13_25_real;
      end
      6'b011010 : begin
        _zz_2779_ = int_reg_array_13_26_imag;
        _zz_2780_ = int_reg_array_13_26_real;
      end
      6'b011011 : begin
        _zz_2779_ = int_reg_array_13_27_imag;
        _zz_2780_ = int_reg_array_13_27_real;
      end
      6'b011100 : begin
        _zz_2779_ = int_reg_array_13_28_imag;
        _zz_2780_ = int_reg_array_13_28_real;
      end
      6'b011101 : begin
        _zz_2779_ = int_reg_array_13_29_imag;
        _zz_2780_ = int_reg_array_13_29_real;
      end
      6'b011110 : begin
        _zz_2779_ = int_reg_array_13_30_imag;
        _zz_2780_ = int_reg_array_13_30_real;
      end
      6'b011111 : begin
        _zz_2779_ = int_reg_array_13_31_imag;
        _zz_2780_ = int_reg_array_13_31_real;
      end
      6'b100000 : begin
        _zz_2779_ = int_reg_array_13_32_imag;
        _zz_2780_ = int_reg_array_13_32_real;
      end
      6'b100001 : begin
        _zz_2779_ = int_reg_array_13_33_imag;
        _zz_2780_ = int_reg_array_13_33_real;
      end
      6'b100010 : begin
        _zz_2779_ = int_reg_array_13_34_imag;
        _zz_2780_ = int_reg_array_13_34_real;
      end
      6'b100011 : begin
        _zz_2779_ = int_reg_array_13_35_imag;
        _zz_2780_ = int_reg_array_13_35_real;
      end
      6'b100100 : begin
        _zz_2779_ = int_reg_array_13_36_imag;
        _zz_2780_ = int_reg_array_13_36_real;
      end
      6'b100101 : begin
        _zz_2779_ = int_reg_array_13_37_imag;
        _zz_2780_ = int_reg_array_13_37_real;
      end
      6'b100110 : begin
        _zz_2779_ = int_reg_array_13_38_imag;
        _zz_2780_ = int_reg_array_13_38_real;
      end
      6'b100111 : begin
        _zz_2779_ = int_reg_array_13_39_imag;
        _zz_2780_ = int_reg_array_13_39_real;
      end
      6'b101000 : begin
        _zz_2779_ = int_reg_array_13_40_imag;
        _zz_2780_ = int_reg_array_13_40_real;
      end
      6'b101001 : begin
        _zz_2779_ = int_reg_array_13_41_imag;
        _zz_2780_ = int_reg_array_13_41_real;
      end
      6'b101010 : begin
        _zz_2779_ = int_reg_array_13_42_imag;
        _zz_2780_ = int_reg_array_13_42_real;
      end
      6'b101011 : begin
        _zz_2779_ = int_reg_array_13_43_imag;
        _zz_2780_ = int_reg_array_13_43_real;
      end
      6'b101100 : begin
        _zz_2779_ = int_reg_array_13_44_imag;
        _zz_2780_ = int_reg_array_13_44_real;
      end
      6'b101101 : begin
        _zz_2779_ = int_reg_array_13_45_imag;
        _zz_2780_ = int_reg_array_13_45_real;
      end
      6'b101110 : begin
        _zz_2779_ = int_reg_array_13_46_imag;
        _zz_2780_ = int_reg_array_13_46_real;
      end
      6'b101111 : begin
        _zz_2779_ = int_reg_array_13_47_imag;
        _zz_2780_ = int_reg_array_13_47_real;
      end
      6'b110000 : begin
        _zz_2779_ = int_reg_array_13_48_imag;
        _zz_2780_ = int_reg_array_13_48_real;
      end
      default : begin
        _zz_2779_ = int_reg_array_13_49_imag;
        _zz_2780_ = int_reg_array_13_49_real;
      end
    endcase
  end

  always @(*) begin
    case(_zz_772_)
      6'b000000 : begin
        _zz_2781_ = int_reg_array_14_0_imag;
        _zz_2782_ = int_reg_array_14_0_real;
      end
      6'b000001 : begin
        _zz_2781_ = int_reg_array_14_1_imag;
        _zz_2782_ = int_reg_array_14_1_real;
      end
      6'b000010 : begin
        _zz_2781_ = int_reg_array_14_2_imag;
        _zz_2782_ = int_reg_array_14_2_real;
      end
      6'b000011 : begin
        _zz_2781_ = int_reg_array_14_3_imag;
        _zz_2782_ = int_reg_array_14_3_real;
      end
      6'b000100 : begin
        _zz_2781_ = int_reg_array_14_4_imag;
        _zz_2782_ = int_reg_array_14_4_real;
      end
      6'b000101 : begin
        _zz_2781_ = int_reg_array_14_5_imag;
        _zz_2782_ = int_reg_array_14_5_real;
      end
      6'b000110 : begin
        _zz_2781_ = int_reg_array_14_6_imag;
        _zz_2782_ = int_reg_array_14_6_real;
      end
      6'b000111 : begin
        _zz_2781_ = int_reg_array_14_7_imag;
        _zz_2782_ = int_reg_array_14_7_real;
      end
      6'b001000 : begin
        _zz_2781_ = int_reg_array_14_8_imag;
        _zz_2782_ = int_reg_array_14_8_real;
      end
      6'b001001 : begin
        _zz_2781_ = int_reg_array_14_9_imag;
        _zz_2782_ = int_reg_array_14_9_real;
      end
      6'b001010 : begin
        _zz_2781_ = int_reg_array_14_10_imag;
        _zz_2782_ = int_reg_array_14_10_real;
      end
      6'b001011 : begin
        _zz_2781_ = int_reg_array_14_11_imag;
        _zz_2782_ = int_reg_array_14_11_real;
      end
      6'b001100 : begin
        _zz_2781_ = int_reg_array_14_12_imag;
        _zz_2782_ = int_reg_array_14_12_real;
      end
      6'b001101 : begin
        _zz_2781_ = int_reg_array_14_13_imag;
        _zz_2782_ = int_reg_array_14_13_real;
      end
      6'b001110 : begin
        _zz_2781_ = int_reg_array_14_14_imag;
        _zz_2782_ = int_reg_array_14_14_real;
      end
      6'b001111 : begin
        _zz_2781_ = int_reg_array_14_15_imag;
        _zz_2782_ = int_reg_array_14_15_real;
      end
      6'b010000 : begin
        _zz_2781_ = int_reg_array_14_16_imag;
        _zz_2782_ = int_reg_array_14_16_real;
      end
      6'b010001 : begin
        _zz_2781_ = int_reg_array_14_17_imag;
        _zz_2782_ = int_reg_array_14_17_real;
      end
      6'b010010 : begin
        _zz_2781_ = int_reg_array_14_18_imag;
        _zz_2782_ = int_reg_array_14_18_real;
      end
      6'b010011 : begin
        _zz_2781_ = int_reg_array_14_19_imag;
        _zz_2782_ = int_reg_array_14_19_real;
      end
      6'b010100 : begin
        _zz_2781_ = int_reg_array_14_20_imag;
        _zz_2782_ = int_reg_array_14_20_real;
      end
      6'b010101 : begin
        _zz_2781_ = int_reg_array_14_21_imag;
        _zz_2782_ = int_reg_array_14_21_real;
      end
      6'b010110 : begin
        _zz_2781_ = int_reg_array_14_22_imag;
        _zz_2782_ = int_reg_array_14_22_real;
      end
      6'b010111 : begin
        _zz_2781_ = int_reg_array_14_23_imag;
        _zz_2782_ = int_reg_array_14_23_real;
      end
      6'b011000 : begin
        _zz_2781_ = int_reg_array_14_24_imag;
        _zz_2782_ = int_reg_array_14_24_real;
      end
      6'b011001 : begin
        _zz_2781_ = int_reg_array_14_25_imag;
        _zz_2782_ = int_reg_array_14_25_real;
      end
      6'b011010 : begin
        _zz_2781_ = int_reg_array_14_26_imag;
        _zz_2782_ = int_reg_array_14_26_real;
      end
      6'b011011 : begin
        _zz_2781_ = int_reg_array_14_27_imag;
        _zz_2782_ = int_reg_array_14_27_real;
      end
      6'b011100 : begin
        _zz_2781_ = int_reg_array_14_28_imag;
        _zz_2782_ = int_reg_array_14_28_real;
      end
      6'b011101 : begin
        _zz_2781_ = int_reg_array_14_29_imag;
        _zz_2782_ = int_reg_array_14_29_real;
      end
      6'b011110 : begin
        _zz_2781_ = int_reg_array_14_30_imag;
        _zz_2782_ = int_reg_array_14_30_real;
      end
      6'b011111 : begin
        _zz_2781_ = int_reg_array_14_31_imag;
        _zz_2782_ = int_reg_array_14_31_real;
      end
      6'b100000 : begin
        _zz_2781_ = int_reg_array_14_32_imag;
        _zz_2782_ = int_reg_array_14_32_real;
      end
      6'b100001 : begin
        _zz_2781_ = int_reg_array_14_33_imag;
        _zz_2782_ = int_reg_array_14_33_real;
      end
      6'b100010 : begin
        _zz_2781_ = int_reg_array_14_34_imag;
        _zz_2782_ = int_reg_array_14_34_real;
      end
      6'b100011 : begin
        _zz_2781_ = int_reg_array_14_35_imag;
        _zz_2782_ = int_reg_array_14_35_real;
      end
      6'b100100 : begin
        _zz_2781_ = int_reg_array_14_36_imag;
        _zz_2782_ = int_reg_array_14_36_real;
      end
      6'b100101 : begin
        _zz_2781_ = int_reg_array_14_37_imag;
        _zz_2782_ = int_reg_array_14_37_real;
      end
      6'b100110 : begin
        _zz_2781_ = int_reg_array_14_38_imag;
        _zz_2782_ = int_reg_array_14_38_real;
      end
      6'b100111 : begin
        _zz_2781_ = int_reg_array_14_39_imag;
        _zz_2782_ = int_reg_array_14_39_real;
      end
      6'b101000 : begin
        _zz_2781_ = int_reg_array_14_40_imag;
        _zz_2782_ = int_reg_array_14_40_real;
      end
      6'b101001 : begin
        _zz_2781_ = int_reg_array_14_41_imag;
        _zz_2782_ = int_reg_array_14_41_real;
      end
      6'b101010 : begin
        _zz_2781_ = int_reg_array_14_42_imag;
        _zz_2782_ = int_reg_array_14_42_real;
      end
      6'b101011 : begin
        _zz_2781_ = int_reg_array_14_43_imag;
        _zz_2782_ = int_reg_array_14_43_real;
      end
      6'b101100 : begin
        _zz_2781_ = int_reg_array_14_44_imag;
        _zz_2782_ = int_reg_array_14_44_real;
      end
      6'b101101 : begin
        _zz_2781_ = int_reg_array_14_45_imag;
        _zz_2782_ = int_reg_array_14_45_real;
      end
      6'b101110 : begin
        _zz_2781_ = int_reg_array_14_46_imag;
        _zz_2782_ = int_reg_array_14_46_real;
      end
      6'b101111 : begin
        _zz_2781_ = int_reg_array_14_47_imag;
        _zz_2782_ = int_reg_array_14_47_real;
      end
      6'b110000 : begin
        _zz_2781_ = int_reg_array_14_48_imag;
        _zz_2782_ = int_reg_array_14_48_real;
      end
      default : begin
        _zz_2781_ = int_reg_array_14_49_imag;
        _zz_2782_ = int_reg_array_14_49_real;
      end
    endcase
  end

  always @(*) begin
    case(_zz_827_)
      6'b000000 : begin
        _zz_2783_ = int_reg_array_15_0_imag;
        _zz_2784_ = int_reg_array_15_0_real;
      end
      6'b000001 : begin
        _zz_2783_ = int_reg_array_15_1_imag;
        _zz_2784_ = int_reg_array_15_1_real;
      end
      6'b000010 : begin
        _zz_2783_ = int_reg_array_15_2_imag;
        _zz_2784_ = int_reg_array_15_2_real;
      end
      6'b000011 : begin
        _zz_2783_ = int_reg_array_15_3_imag;
        _zz_2784_ = int_reg_array_15_3_real;
      end
      6'b000100 : begin
        _zz_2783_ = int_reg_array_15_4_imag;
        _zz_2784_ = int_reg_array_15_4_real;
      end
      6'b000101 : begin
        _zz_2783_ = int_reg_array_15_5_imag;
        _zz_2784_ = int_reg_array_15_5_real;
      end
      6'b000110 : begin
        _zz_2783_ = int_reg_array_15_6_imag;
        _zz_2784_ = int_reg_array_15_6_real;
      end
      6'b000111 : begin
        _zz_2783_ = int_reg_array_15_7_imag;
        _zz_2784_ = int_reg_array_15_7_real;
      end
      6'b001000 : begin
        _zz_2783_ = int_reg_array_15_8_imag;
        _zz_2784_ = int_reg_array_15_8_real;
      end
      6'b001001 : begin
        _zz_2783_ = int_reg_array_15_9_imag;
        _zz_2784_ = int_reg_array_15_9_real;
      end
      6'b001010 : begin
        _zz_2783_ = int_reg_array_15_10_imag;
        _zz_2784_ = int_reg_array_15_10_real;
      end
      6'b001011 : begin
        _zz_2783_ = int_reg_array_15_11_imag;
        _zz_2784_ = int_reg_array_15_11_real;
      end
      6'b001100 : begin
        _zz_2783_ = int_reg_array_15_12_imag;
        _zz_2784_ = int_reg_array_15_12_real;
      end
      6'b001101 : begin
        _zz_2783_ = int_reg_array_15_13_imag;
        _zz_2784_ = int_reg_array_15_13_real;
      end
      6'b001110 : begin
        _zz_2783_ = int_reg_array_15_14_imag;
        _zz_2784_ = int_reg_array_15_14_real;
      end
      6'b001111 : begin
        _zz_2783_ = int_reg_array_15_15_imag;
        _zz_2784_ = int_reg_array_15_15_real;
      end
      6'b010000 : begin
        _zz_2783_ = int_reg_array_15_16_imag;
        _zz_2784_ = int_reg_array_15_16_real;
      end
      6'b010001 : begin
        _zz_2783_ = int_reg_array_15_17_imag;
        _zz_2784_ = int_reg_array_15_17_real;
      end
      6'b010010 : begin
        _zz_2783_ = int_reg_array_15_18_imag;
        _zz_2784_ = int_reg_array_15_18_real;
      end
      6'b010011 : begin
        _zz_2783_ = int_reg_array_15_19_imag;
        _zz_2784_ = int_reg_array_15_19_real;
      end
      6'b010100 : begin
        _zz_2783_ = int_reg_array_15_20_imag;
        _zz_2784_ = int_reg_array_15_20_real;
      end
      6'b010101 : begin
        _zz_2783_ = int_reg_array_15_21_imag;
        _zz_2784_ = int_reg_array_15_21_real;
      end
      6'b010110 : begin
        _zz_2783_ = int_reg_array_15_22_imag;
        _zz_2784_ = int_reg_array_15_22_real;
      end
      6'b010111 : begin
        _zz_2783_ = int_reg_array_15_23_imag;
        _zz_2784_ = int_reg_array_15_23_real;
      end
      6'b011000 : begin
        _zz_2783_ = int_reg_array_15_24_imag;
        _zz_2784_ = int_reg_array_15_24_real;
      end
      6'b011001 : begin
        _zz_2783_ = int_reg_array_15_25_imag;
        _zz_2784_ = int_reg_array_15_25_real;
      end
      6'b011010 : begin
        _zz_2783_ = int_reg_array_15_26_imag;
        _zz_2784_ = int_reg_array_15_26_real;
      end
      6'b011011 : begin
        _zz_2783_ = int_reg_array_15_27_imag;
        _zz_2784_ = int_reg_array_15_27_real;
      end
      6'b011100 : begin
        _zz_2783_ = int_reg_array_15_28_imag;
        _zz_2784_ = int_reg_array_15_28_real;
      end
      6'b011101 : begin
        _zz_2783_ = int_reg_array_15_29_imag;
        _zz_2784_ = int_reg_array_15_29_real;
      end
      6'b011110 : begin
        _zz_2783_ = int_reg_array_15_30_imag;
        _zz_2784_ = int_reg_array_15_30_real;
      end
      6'b011111 : begin
        _zz_2783_ = int_reg_array_15_31_imag;
        _zz_2784_ = int_reg_array_15_31_real;
      end
      6'b100000 : begin
        _zz_2783_ = int_reg_array_15_32_imag;
        _zz_2784_ = int_reg_array_15_32_real;
      end
      6'b100001 : begin
        _zz_2783_ = int_reg_array_15_33_imag;
        _zz_2784_ = int_reg_array_15_33_real;
      end
      6'b100010 : begin
        _zz_2783_ = int_reg_array_15_34_imag;
        _zz_2784_ = int_reg_array_15_34_real;
      end
      6'b100011 : begin
        _zz_2783_ = int_reg_array_15_35_imag;
        _zz_2784_ = int_reg_array_15_35_real;
      end
      6'b100100 : begin
        _zz_2783_ = int_reg_array_15_36_imag;
        _zz_2784_ = int_reg_array_15_36_real;
      end
      6'b100101 : begin
        _zz_2783_ = int_reg_array_15_37_imag;
        _zz_2784_ = int_reg_array_15_37_real;
      end
      6'b100110 : begin
        _zz_2783_ = int_reg_array_15_38_imag;
        _zz_2784_ = int_reg_array_15_38_real;
      end
      6'b100111 : begin
        _zz_2783_ = int_reg_array_15_39_imag;
        _zz_2784_ = int_reg_array_15_39_real;
      end
      6'b101000 : begin
        _zz_2783_ = int_reg_array_15_40_imag;
        _zz_2784_ = int_reg_array_15_40_real;
      end
      6'b101001 : begin
        _zz_2783_ = int_reg_array_15_41_imag;
        _zz_2784_ = int_reg_array_15_41_real;
      end
      6'b101010 : begin
        _zz_2783_ = int_reg_array_15_42_imag;
        _zz_2784_ = int_reg_array_15_42_real;
      end
      6'b101011 : begin
        _zz_2783_ = int_reg_array_15_43_imag;
        _zz_2784_ = int_reg_array_15_43_real;
      end
      6'b101100 : begin
        _zz_2783_ = int_reg_array_15_44_imag;
        _zz_2784_ = int_reg_array_15_44_real;
      end
      6'b101101 : begin
        _zz_2783_ = int_reg_array_15_45_imag;
        _zz_2784_ = int_reg_array_15_45_real;
      end
      6'b101110 : begin
        _zz_2783_ = int_reg_array_15_46_imag;
        _zz_2784_ = int_reg_array_15_46_real;
      end
      6'b101111 : begin
        _zz_2783_ = int_reg_array_15_47_imag;
        _zz_2784_ = int_reg_array_15_47_real;
      end
      6'b110000 : begin
        _zz_2783_ = int_reg_array_15_48_imag;
        _zz_2784_ = int_reg_array_15_48_real;
      end
      default : begin
        _zz_2783_ = int_reg_array_15_49_imag;
        _zz_2784_ = int_reg_array_15_49_real;
      end
    endcase
  end

  always @(*) begin
    case(_zz_882_)
      6'b000000 : begin
        _zz_2785_ = int_reg_array_16_0_imag;
        _zz_2786_ = int_reg_array_16_0_real;
      end
      6'b000001 : begin
        _zz_2785_ = int_reg_array_16_1_imag;
        _zz_2786_ = int_reg_array_16_1_real;
      end
      6'b000010 : begin
        _zz_2785_ = int_reg_array_16_2_imag;
        _zz_2786_ = int_reg_array_16_2_real;
      end
      6'b000011 : begin
        _zz_2785_ = int_reg_array_16_3_imag;
        _zz_2786_ = int_reg_array_16_3_real;
      end
      6'b000100 : begin
        _zz_2785_ = int_reg_array_16_4_imag;
        _zz_2786_ = int_reg_array_16_4_real;
      end
      6'b000101 : begin
        _zz_2785_ = int_reg_array_16_5_imag;
        _zz_2786_ = int_reg_array_16_5_real;
      end
      6'b000110 : begin
        _zz_2785_ = int_reg_array_16_6_imag;
        _zz_2786_ = int_reg_array_16_6_real;
      end
      6'b000111 : begin
        _zz_2785_ = int_reg_array_16_7_imag;
        _zz_2786_ = int_reg_array_16_7_real;
      end
      6'b001000 : begin
        _zz_2785_ = int_reg_array_16_8_imag;
        _zz_2786_ = int_reg_array_16_8_real;
      end
      6'b001001 : begin
        _zz_2785_ = int_reg_array_16_9_imag;
        _zz_2786_ = int_reg_array_16_9_real;
      end
      6'b001010 : begin
        _zz_2785_ = int_reg_array_16_10_imag;
        _zz_2786_ = int_reg_array_16_10_real;
      end
      6'b001011 : begin
        _zz_2785_ = int_reg_array_16_11_imag;
        _zz_2786_ = int_reg_array_16_11_real;
      end
      6'b001100 : begin
        _zz_2785_ = int_reg_array_16_12_imag;
        _zz_2786_ = int_reg_array_16_12_real;
      end
      6'b001101 : begin
        _zz_2785_ = int_reg_array_16_13_imag;
        _zz_2786_ = int_reg_array_16_13_real;
      end
      6'b001110 : begin
        _zz_2785_ = int_reg_array_16_14_imag;
        _zz_2786_ = int_reg_array_16_14_real;
      end
      6'b001111 : begin
        _zz_2785_ = int_reg_array_16_15_imag;
        _zz_2786_ = int_reg_array_16_15_real;
      end
      6'b010000 : begin
        _zz_2785_ = int_reg_array_16_16_imag;
        _zz_2786_ = int_reg_array_16_16_real;
      end
      6'b010001 : begin
        _zz_2785_ = int_reg_array_16_17_imag;
        _zz_2786_ = int_reg_array_16_17_real;
      end
      6'b010010 : begin
        _zz_2785_ = int_reg_array_16_18_imag;
        _zz_2786_ = int_reg_array_16_18_real;
      end
      6'b010011 : begin
        _zz_2785_ = int_reg_array_16_19_imag;
        _zz_2786_ = int_reg_array_16_19_real;
      end
      6'b010100 : begin
        _zz_2785_ = int_reg_array_16_20_imag;
        _zz_2786_ = int_reg_array_16_20_real;
      end
      6'b010101 : begin
        _zz_2785_ = int_reg_array_16_21_imag;
        _zz_2786_ = int_reg_array_16_21_real;
      end
      6'b010110 : begin
        _zz_2785_ = int_reg_array_16_22_imag;
        _zz_2786_ = int_reg_array_16_22_real;
      end
      6'b010111 : begin
        _zz_2785_ = int_reg_array_16_23_imag;
        _zz_2786_ = int_reg_array_16_23_real;
      end
      6'b011000 : begin
        _zz_2785_ = int_reg_array_16_24_imag;
        _zz_2786_ = int_reg_array_16_24_real;
      end
      6'b011001 : begin
        _zz_2785_ = int_reg_array_16_25_imag;
        _zz_2786_ = int_reg_array_16_25_real;
      end
      6'b011010 : begin
        _zz_2785_ = int_reg_array_16_26_imag;
        _zz_2786_ = int_reg_array_16_26_real;
      end
      6'b011011 : begin
        _zz_2785_ = int_reg_array_16_27_imag;
        _zz_2786_ = int_reg_array_16_27_real;
      end
      6'b011100 : begin
        _zz_2785_ = int_reg_array_16_28_imag;
        _zz_2786_ = int_reg_array_16_28_real;
      end
      6'b011101 : begin
        _zz_2785_ = int_reg_array_16_29_imag;
        _zz_2786_ = int_reg_array_16_29_real;
      end
      6'b011110 : begin
        _zz_2785_ = int_reg_array_16_30_imag;
        _zz_2786_ = int_reg_array_16_30_real;
      end
      6'b011111 : begin
        _zz_2785_ = int_reg_array_16_31_imag;
        _zz_2786_ = int_reg_array_16_31_real;
      end
      6'b100000 : begin
        _zz_2785_ = int_reg_array_16_32_imag;
        _zz_2786_ = int_reg_array_16_32_real;
      end
      6'b100001 : begin
        _zz_2785_ = int_reg_array_16_33_imag;
        _zz_2786_ = int_reg_array_16_33_real;
      end
      6'b100010 : begin
        _zz_2785_ = int_reg_array_16_34_imag;
        _zz_2786_ = int_reg_array_16_34_real;
      end
      6'b100011 : begin
        _zz_2785_ = int_reg_array_16_35_imag;
        _zz_2786_ = int_reg_array_16_35_real;
      end
      6'b100100 : begin
        _zz_2785_ = int_reg_array_16_36_imag;
        _zz_2786_ = int_reg_array_16_36_real;
      end
      6'b100101 : begin
        _zz_2785_ = int_reg_array_16_37_imag;
        _zz_2786_ = int_reg_array_16_37_real;
      end
      6'b100110 : begin
        _zz_2785_ = int_reg_array_16_38_imag;
        _zz_2786_ = int_reg_array_16_38_real;
      end
      6'b100111 : begin
        _zz_2785_ = int_reg_array_16_39_imag;
        _zz_2786_ = int_reg_array_16_39_real;
      end
      6'b101000 : begin
        _zz_2785_ = int_reg_array_16_40_imag;
        _zz_2786_ = int_reg_array_16_40_real;
      end
      6'b101001 : begin
        _zz_2785_ = int_reg_array_16_41_imag;
        _zz_2786_ = int_reg_array_16_41_real;
      end
      6'b101010 : begin
        _zz_2785_ = int_reg_array_16_42_imag;
        _zz_2786_ = int_reg_array_16_42_real;
      end
      6'b101011 : begin
        _zz_2785_ = int_reg_array_16_43_imag;
        _zz_2786_ = int_reg_array_16_43_real;
      end
      6'b101100 : begin
        _zz_2785_ = int_reg_array_16_44_imag;
        _zz_2786_ = int_reg_array_16_44_real;
      end
      6'b101101 : begin
        _zz_2785_ = int_reg_array_16_45_imag;
        _zz_2786_ = int_reg_array_16_45_real;
      end
      6'b101110 : begin
        _zz_2785_ = int_reg_array_16_46_imag;
        _zz_2786_ = int_reg_array_16_46_real;
      end
      6'b101111 : begin
        _zz_2785_ = int_reg_array_16_47_imag;
        _zz_2786_ = int_reg_array_16_47_real;
      end
      6'b110000 : begin
        _zz_2785_ = int_reg_array_16_48_imag;
        _zz_2786_ = int_reg_array_16_48_real;
      end
      default : begin
        _zz_2785_ = int_reg_array_16_49_imag;
        _zz_2786_ = int_reg_array_16_49_real;
      end
    endcase
  end

  always @(*) begin
    case(_zz_937_)
      6'b000000 : begin
        _zz_2787_ = int_reg_array_17_0_imag;
        _zz_2788_ = int_reg_array_17_0_real;
      end
      6'b000001 : begin
        _zz_2787_ = int_reg_array_17_1_imag;
        _zz_2788_ = int_reg_array_17_1_real;
      end
      6'b000010 : begin
        _zz_2787_ = int_reg_array_17_2_imag;
        _zz_2788_ = int_reg_array_17_2_real;
      end
      6'b000011 : begin
        _zz_2787_ = int_reg_array_17_3_imag;
        _zz_2788_ = int_reg_array_17_3_real;
      end
      6'b000100 : begin
        _zz_2787_ = int_reg_array_17_4_imag;
        _zz_2788_ = int_reg_array_17_4_real;
      end
      6'b000101 : begin
        _zz_2787_ = int_reg_array_17_5_imag;
        _zz_2788_ = int_reg_array_17_5_real;
      end
      6'b000110 : begin
        _zz_2787_ = int_reg_array_17_6_imag;
        _zz_2788_ = int_reg_array_17_6_real;
      end
      6'b000111 : begin
        _zz_2787_ = int_reg_array_17_7_imag;
        _zz_2788_ = int_reg_array_17_7_real;
      end
      6'b001000 : begin
        _zz_2787_ = int_reg_array_17_8_imag;
        _zz_2788_ = int_reg_array_17_8_real;
      end
      6'b001001 : begin
        _zz_2787_ = int_reg_array_17_9_imag;
        _zz_2788_ = int_reg_array_17_9_real;
      end
      6'b001010 : begin
        _zz_2787_ = int_reg_array_17_10_imag;
        _zz_2788_ = int_reg_array_17_10_real;
      end
      6'b001011 : begin
        _zz_2787_ = int_reg_array_17_11_imag;
        _zz_2788_ = int_reg_array_17_11_real;
      end
      6'b001100 : begin
        _zz_2787_ = int_reg_array_17_12_imag;
        _zz_2788_ = int_reg_array_17_12_real;
      end
      6'b001101 : begin
        _zz_2787_ = int_reg_array_17_13_imag;
        _zz_2788_ = int_reg_array_17_13_real;
      end
      6'b001110 : begin
        _zz_2787_ = int_reg_array_17_14_imag;
        _zz_2788_ = int_reg_array_17_14_real;
      end
      6'b001111 : begin
        _zz_2787_ = int_reg_array_17_15_imag;
        _zz_2788_ = int_reg_array_17_15_real;
      end
      6'b010000 : begin
        _zz_2787_ = int_reg_array_17_16_imag;
        _zz_2788_ = int_reg_array_17_16_real;
      end
      6'b010001 : begin
        _zz_2787_ = int_reg_array_17_17_imag;
        _zz_2788_ = int_reg_array_17_17_real;
      end
      6'b010010 : begin
        _zz_2787_ = int_reg_array_17_18_imag;
        _zz_2788_ = int_reg_array_17_18_real;
      end
      6'b010011 : begin
        _zz_2787_ = int_reg_array_17_19_imag;
        _zz_2788_ = int_reg_array_17_19_real;
      end
      6'b010100 : begin
        _zz_2787_ = int_reg_array_17_20_imag;
        _zz_2788_ = int_reg_array_17_20_real;
      end
      6'b010101 : begin
        _zz_2787_ = int_reg_array_17_21_imag;
        _zz_2788_ = int_reg_array_17_21_real;
      end
      6'b010110 : begin
        _zz_2787_ = int_reg_array_17_22_imag;
        _zz_2788_ = int_reg_array_17_22_real;
      end
      6'b010111 : begin
        _zz_2787_ = int_reg_array_17_23_imag;
        _zz_2788_ = int_reg_array_17_23_real;
      end
      6'b011000 : begin
        _zz_2787_ = int_reg_array_17_24_imag;
        _zz_2788_ = int_reg_array_17_24_real;
      end
      6'b011001 : begin
        _zz_2787_ = int_reg_array_17_25_imag;
        _zz_2788_ = int_reg_array_17_25_real;
      end
      6'b011010 : begin
        _zz_2787_ = int_reg_array_17_26_imag;
        _zz_2788_ = int_reg_array_17_26_real;
      end
      6'b011011 : begin
        _zz_2787_ = int_reg_array_17_27_imag;
        _zz_2788_ = int_reg_array_17_27_real;
      end
      6'b011100 : begin
        _zz_2787_ = int_reg_array_17_28_imag;
        _zz_2788_ = int_reg_array_17_28_real;
      end
      6'b011101 : begin
        _zz_2787_ = int_reg_array_17_29_imag;
        _zz_2788_ = int_reg_array_17_29_real;
      end
      6'b011110 : begin
        _zz_2787_ = int_reg_array_17_30_imag;
        _zz_2788_ = int_reg_array_17_30_real;
      end
      6'b011111 : begin
        _zz_2787_ = int_reg_array_17_31_imag;
        _zz_2788_ = int_reg_array_17_31_real;
      end
      6'b100000 : begin
        _zz_2787_ = int_reg_array_17_32_imag;
        _zz_2788_ = int_reg_array_17_32_real;
      end
      6'b100001 : begin
        _zz_2787_ = int_reg_array_17_33_imag;
        _zz_2788_ = int_reg_array_17_33_real;
      end
      6'b100010 : begin
        _zz_2787_ = int_reg_array_17_34_imag;
        _zz_2788_ = int_reg_array_17_34_real;
      end
      6'b100011 : begin
        _zz_2787_ = int_reg_array_17_35_imag;
        _zz_2788_ = int_reg_array_17_35_real;
      end
      6'b100100 : begin
        _zz_2787_ = int_reg_array_17_36_imag;
        _zz_2788_ = int_reg_array_17_36_real;
      end
      6'b100101 : begin
        _zz_2787_ = int_reg_array_17_37_imag;
        _zz_2788_ = int_reg_array_17_37_real;
      end
      6'b100110 : begin
        _zz_2787_ = int_reg_array_17_38_imag;
        _zz_2788_ = int_reg_array_17_38_real;
      end
      6'b100111 : begin
        _zz_2787_ = int_reg_array_17_39_imag;
        _zz_2788_ = int_reg_array_17_39_real;
      end
      6'b101000 : begin
        _zz_2787_ = int_reg_array_17_40_imag;
        _zz_2788_ = int_reg_array_17_40_real;
      end
      6'b101001 : begin
        _zz_2787_ = int_reg_array_17_41_imag;
        _zz_2788_ = int_reg_array_17_41_real;
      end
      6'b101010 : begin
        _zz_2787_ = int_reg_array_17_42_imag;
        _zz_2788_ = int_reg_array_17_42_real;
      end
      6'b101011 : begin
        _zz_2787_ = int_reg_array_17_43_imag;
        _zz_2788_ = int_reg_array_17_43_real;
      end
      6'b101100 : begin
        _zz_2787_ = int_reg_array_17_44_imag;
        _zz_2788_ = int_reg_array_17_44_real;
      end
      6'b101101 : begin
        _zz_2787_ = int_reg_array_17_45_imag;
        _zz_2788_ = int_reg_array_17_45_real;
      end
      6'b101110 : begin
        _zz_2787_ = int_reg_array_17_46_imag;
        _zz_2788_ = int_reg_array_17_46_real;
      end
      6'b101111 : begin
        _zz_2787_ = int_reg_array_17_47_imag;
        _zz_2788_ = int_reg_array_17_47_real;
      end
      6'b110000 : begin
        _zz_2787_ = int_reg_array_17_48_imag;
        _zz_2788_ = int_reg_array_17_48_real;
      end
      default : begin
        _zz_2787_ = int_reg_array_17_49_imag;
        _zz_2788_ = int_reg_array_17_49_real;
      end
    endcase
  end

  always @(*) begin
    case(_zz_992_)
      6'b000000 : begin
        _zz_2789_ = int_reg_array_18_0_imag;
        _zz_2790_ = int_reg_array_18_0_real;
      end
      6'b000001 : begin
        _zz_2789_ = int_reg_array_18_1_imag;
        _zz_2790_ = int_reg_array_18_1_real;
      end
      6'b000010 : begin
        _zz_2789_ = int_reg_array_18_2_imag;
        _zz_2790_ = int_reg_array_18_2_real;
      end
      6'b000011 : begin
        _zz_2789_ = int_reg_array_18_3_imag;
        _zz_2790_ = int_reg_array_18_3_real;
      end
      6'b000100 : begin
        _zz_2789_ = int_reg_array_18_4_imag;
        _zz_2790_ = int_reg_array_18_4_real;
      end
      6'b000101 : begin
        _zz_2789_ = int_reg_array_18_5_imag;
        _zz_2790_ = int_reg_array_18_5_real;
      end
      6'b000110 : begin
        _zz_2789_ = int_reg_array_18_6_imag;
        _zz_2790_ = int_reg_array_18_6_real;
      end
      6'b000111 : begin
        _zz_2789_ = int_reg_array_18_7_imag;
        _zz_2790_ = int_reg_array_18_7_real;
      end
      6'b001000 : begin
        _zz_2789_ = int_reg_array_18_8_imag;
        _zz_2790_ = int_reg_array_18_8_real;
      end
      6'b001001 : begin
        _zz_2789_ = int_reg_array_18_9_imag;
        _zz_2790_ = int_reg_array_18_9_real;
      end
      6'b001010 : begin
        _zz_2789_ = int_reg_array_18_10_imag;
        _zz_2790_ = int_reg_array_18_10_real;
      end
      6'b001011 : begin
        _zz_2789_ = int_reg_array_18_11_imag;
        _zz_2790_ = int_reg_array_18_11_real;
      end
      6'b001100 : begin
        _zz_2789_ = int_reg_array_18_12_imag;
        _zz_2790_ = int_reg_array_18_12_real;
      end
      6'b001101 : begin
        _zz_2789_ = int_reg_array_18_13_imag;
        _zz_2790_ = int_reg_array_18_13_real;
      end
      6'b001110 : begin
        _zz_2789_ = int_reg_array_18_14_imag;
        _zz_2790_ = int_reg_array_18_14_real;
      end
      6'b001111 : begin
        _zz_2789_ = int_reg_array_18_15_imag;
        _zz_2790_ = int_reg_array_18_15_real;
      end
      6'b010000 : begin
        _zz_2789_ = int_reg_array_18_16_imag;
        _zz_2790_ = int_reg_array_18_16_real;
      end
      6'b010001 : begin
        _zz_2789_ = int_reg_array_18_17_imag;
        _zz_2790_ = int_reg_array_18_17_real;
      end
      6'b010010 : begin
        _zz_2789_ = int_reg_array_18_18_imag;
        _zz_2790_ = int_reg_array_18_18_real;
      end
      6'b010011 : begin
        _zz_2789_ = int_reg_array_18_19_imag;
        _zz_2790_ = int_reg_array_18_19_real;
      end
      6'b010100 : begin
        _zz_2789_ = int_reg_array_18_20_imag;
        _zz_2790_ = int_reg_array_18_20_real;
      end
      6'b010101 : begin
        _zz_2789_ = int_reg_array_18_21_imag;
        _zz_2790_ = int_reg_array_18_21_real;
      end
      6'b010110 : begin
        _zz_2789_ = int_reg_array_18_22_imag;
        _zz_2790_ = int_reg_array_18_22_real;
      end
      6'b010111 : begin
        _zz_2789_ = int_reg_array_18_23_imag;
        _zz_2790_ = int_reg_array_18_23_real;
      end
      6'b011000 : begin
        _zz_2789_ = int_reg_array_18_24_imag;
        _zz_2790_ = int_reg_array_18_24_real;
      end
      6'b011001 : begin
        _zz_2789_ = int_reg_array_18_25_imag;
        _zz_2790_ = int_reg_array_18_25_real;
      end
      6'b011010 : begin
        _zz_2789_ = int_reg_array_18_26_imag;
        _zz_2790_ = int_reg_array_18_26_real;
      end
      6'b011011 : begin
        _zz_2789_ = int_reg_array_18_27_imag;
        _zz_2790_ = int_reg_array_18_27_real;
      end
      6'b011100 : begin
        _zz_2789_ = int_reg_array_18_28_imag;
        _zz_2790_ = int_reg_array_18_28_real;
      end
      6'b011101 : begin
        _zz_2789_ = int_reg_array_18_29_imag;
        _zz_2790_ = int_reg_array_18_29_real;
      end
      6'b011110 : begin
        _zz_2789_ = int_reg_array_18_30_imag;
        _zz_2790_ = int_reg_array_18_30_real;
      end
      6'b011111 : begin
        _zz_2789_ = int_reg_array_18_31_imag;
        _zz_2790_ = int_reg_array_18_31_real;
      end
      6'b100000 : begin
        _zz_2789_ = int_reg_array_18_32_imag;
        _zz_2790_ = int_reg_array_18_32_real;
      end
      6'b100001 : begin
        _zz_2789_ = int_reg_array_18_33_imag;
        _zz_2790_ = int_reg_array_18_33_real;
      end
      6'b100010 : begin
        _zz_2789_ = int_reg_array_18_34_imag;
        _zz_2790_ = int_reg_array_18_34_real;
      end
      6'b100011 : begin
        _zz_2789_ = int_reg_array_18_35_imag;
        _zz_2790_ = int_reg_array_18_35_real;
      end
      6'b100100 : begin
        _zz_2789_ = int_reg_array_18_36_imag;
        _zz_2790_ = int_reg_array_18_36_real;
      end
      6'b100101 : begin
        _zz_2789_ = int_reg_array_18_37_imag;
        _zz_2790_ = int_reg_array_18_37_real;
      end
      6'b100110 : begin
        _zz_2789_ = int_reg_array_18_38_imag;
        _zz_2790_ = int_reg_array_18_38_real;
      end
      6'b100111 : begin
        _zz_2789_ = int_reg_array_18_39_imag;
        _zz_2790_ = int_reg_array_18_39_real;
      end
      6'b101000 : begin
        _zz_2789_ = int_reg_array_18_40_imag;
        _zz_2790_ = int_reg_array_18_40_real;
      end
      6'b101001 : begin
        _zz_2789_ = int_reg_array_18_41_imag;
        _zz_2790_ = int_reg_array_18_41_real;
      end
      6'b101010 : begin
        _zz_2789_ = int_reg_array_18_42_imag;
        _zz_2790_ = int_reg_array_18_42_real;
      end
      6'b101011 : begin
        _zz_2789_ = int_reg_array_18_43_imag;
        _zz_2790_ = int_reg_array_18_43_real;
      end
      6'b101100 : begin
        _zz_2789_ = int_reg_array_18_44_imag;
        _zz_2790_ = int_reg_array_18_44_real;
      end
      6'b101101 : begin
        _zz_2789_ = int_reg_array_18_45_imag;
        _zz_2790_ = int_reg_array_18_45_real;
      end
      6'b101110 : begin
        _zz_2789_ = int_reg_array_18_46_imag;
        _zz_2790_ = int_reg_array_18_46_real;
      end
      6'b101111 : begin
        _zz_2789_ = int_reg_array_18_47_imag;
        _zz_2790_ = int_reg_array_18_47_real;
      end
      6'b110000 : begin
        _zz_2789_ = int_reg_array_18_48_imag;
        _zz_2790_ = int_reg_array_18_48_real;
      end
      default : begin
        _zz_2789_ = int_reg_array_18_49_imag;
        _zz_2790_ = int_reg_array_18_49_real;
      end
    endcase
  end

  always @(*) begin
    case(_zz_1047_)
      6'b000000 : begin
        _zz_2791_ = int_reg_array_19_0_imag;
        _zz_2792_ = int_reg_array_19_0_real;
      end
      6'b000001 : begin
        _zz_2791_ = int_reg_array_19_1_imag;
        _zz_2792_ = int_reg_array_19_1_real;
      end
      6'b000010 : begin
        _zz_2791_ = int_reg_array_19_2_imag;
        _zz_2792_ = int_reg_array_19_2_real;
      end
      6'b000011 : begin
        _zz_2791_ = int_reg_array_19_3_imag;
        _zz_2792_ = int_reg_array_19_3_real;
      end
      6'b000100 : begin
        _zz_2791_ = int_reg_array_19_4_imag;
        _zz_2792_ = int_reg_array_19_4_real;
      end
      6'b000101 : begin
        _zz_2791_ = int_reg_array_19_5_imag;
        _zz_2792_ = int_reg_array_19_5_real;
      end
      6'b000110 : begin
        _zz_2791_ = int_reg_array_19_6_imag;
        _zz_2792_ = int_reg_array_19_6_real;
      end
      6'b000111 : begin
        _zz_2791_ = int_reg_array_19_7_imag;
        _zz_2792_ = int_reg_array_19_7_real;
      end
      6'b001000 : begin
        _zz_2791_ = int_reg_array_19_8_imag;
        _zz_2792_ = int_reg_array_19_8_real;
      end
      6'b001001 : begin
        _zz_2791_ = int_reg_array_19_9_imag;
        _zz_2792_ = int_reg_array_19_9_real;
      end
      6'b001010 : begin
        _zz_2791_ = int_reg_array_19_10_imag;
        _zz_2792_ = int_reg_array_19_10_real;
      end
      6'b001011 : begin
        _zz_2791_ = int_reg_array_19_11_imag;
        _zz_2792_ = int_reg_array_19_11_real;
      end
      6'b001100 : begin
        _zz_2791_ = int_reg_array_19_12_imag;
        _zz_2792_ = int_reg_array_19_12_real;
      end
      6'b001101 : begin
        _zz_2791_ = int_reg_array_19_13_imag;
        _zz_2792_ = int_reg_array_19_13_real;
      end
      6'b001110 : begin
        _zz_2791_ = int_reg_array_19_14_imag;
        _zz_2792_ = int_reg_array_19_14_real;
      end
      6'b001111 : begin
        _zz_2791_ = int_reg_array_19_15_imag;
        _zz_2792_ = int_reg_array_19_15_real;
      end
      6'b010000 : begin
        _zz_2791_ = int_reg_array_19_16_imag;
        _zz_2792_ = int_reg_array_19_16_real;
      end
      6'b010001 : begin
        _zz_2791_ = int_reg_array_19_17_imag;
        _zz_2792_ = int_reg_array_19_17_real;
      end
      6'b010010 : begin
        _zz_2791_ = int_reg_array_19_18_imag;
        _zz_2792_ = int_reg_array_19_18_real;
      end
      6'b010011 : begin
        _zz_2791_ = int_reg_array_19_19_imag;
        _zz_2792_ = int_reg_array_19_19_real;
      end
      6'b010100 : begin
        _zz_2791_ = int_reg_array_19_20_imag;
        _zz_2792_ = int_reg_array_19_20_real;
      end
      6'b010101 : begin
        _zz_2791_ = int_reg_array_19_21_imag;
        _zz_2792_ = int_reg_array_19_21_real;
      end
      6'b010110 : begin
        _zz_2791_ = int_reg_array_19_22_imag;
        _zz_2792_ = int_reg_array_19_22_real;
      end
      6'b010111 : begin
        _zz_2791_ = int_reg_array_19_23_imag;
        _zz_2792_ = int_reg_array_19_23_real;
      end
      6'b011000 : begin
        _zz_2791_ = int_reg_array_19_24_imag;
        _zz_2792_ = int_reg_array_19_24_real;
      end
      6'b011001 : begin
        _zz_2791_ = int_reg_array_19_25_imag;
        _zz_2792_ = int_reg_array_19_25_real;
      end
      6'b011010 : begin
        _zz_2791_ = int_reg_array_19_26_imag;
        _zz_2792_ = int_reg_array_19_26_real;
      end
      6'b011011 : begin
        _zz_2791_ = int_reg_array_19_27_imag;
        _zz_2792_ = int_reg_array_19_27_real;
      end
      6'b011100 : begin
        _zz_2791_ = int_reg_array_19_28_imag;
        _zz_2792_ = int_reg_array_19_28_real;
      end
      6'b011101 : begin
        _zz_2791_ = int_reg_array_19_29_imag;
        _zz_2792_ = int_reg_array_19_29_real;
      end
      6'b011110 : begin
        _zz_2791_ = int_reg_array_19_30_imag;
        _zz_2792_ = int_reg_array_19_30_real;
      end
      6'b011111 : begin
        _zz_2791_ = int_reg_array_19_31_imag;
        _zz_2792_ = int_reg_array_19_31_real;
      end
      6'b100000 : begin
        _zz_2791_ = int_reg_array_19_32_imag;
        _zz_2792_ = int_reg_array_19_32_real;
      end
      6'b100001 : begin
        _zz_2791_ = int_reg_array_19_33_imag;
        _zz_2792_ = int_reg_array_19_33_real;
      end
      6'b100010 : begin
        _zz_2791_ = int_reg_array_19_34_imag;
        _zz_2792_ = int_reg_array_19_34_real;
      end
      6'b100011 : begin
        _zz_2791_ = int_reg_array_19_35_imag;
        _zz_2792_ = int_reg_array_19_35_real;
      end
      6'b100100 : begin
        _zz_2791_ = int_reg_array_19_36_imag;
        _zz_2792_ = int_reg_array_19_36_real;
      end
      6'b100101 : begin
        _zz_2791_ = int_reg_array_19_37_imag;
        _zz_2792_ = int_reg_array_19_37_real;
      end
      6'b100110 : begin
        _zz_2791_ = int_reg_array_19_38_imag;
        _zz_2792_ = int_reg_array_19_38_real;
      end
      6'b100111 : begin
        _zz_2791_ = int_reg_array_19_39_imag;
        _zz_2792_ = int_reg_array_19_39_real;
      end
      6'b101000 : begin
        _zz_2791_ = int_reg_array_19_40_imag;
        _zz_2792_ = int_reg_array_19_40_real;
      end
      6'b101001 : begin
        _zz_2791_ = int_reg_array_19_41_imag;
        _zz_2792_ = int_reg_array_19_41_real;
      end
      6'b101010 : begin
        _zz_2791_ = int_reg_array_19_42_imag;
        _zz_2792_ = int_reg_array_19_42_real;
      end
      6'b101011 : begin
        _zz_2791_ = int_reg_array_19_43_imag;
        _zz_2792_ = int_reg_array_19_43_real;
      end
      6'b101100 : begin
        _zz_2791_ = int_reg_array_19_44_imag;
        _zz_2792_ = int_reg_array_19_44_real;
      end
      6'b101101 : begin
        _zz_2791_ = int_reg_array_19_45_imag;
        _zz_2792_ = int_reg_array_19_45_real;
      end
      6'b101110 : begin
        _zz_2791_ = int_reg_array_19_46_imag;
        _zz_2792_ = int_reg_array_19_46_real;
      end
      6'b101111 : begin
        _zz_2791_ = int_reg_array_19_47_imag;
        _zz_2792_ = int_reg_array_19_47_real;
      end
      6'b110000 : begin
        _zz_2791_ = int_reg_array_19_48_imag;
        _zz_2792_ = int_reg_array_19_48_real;
      end
      default : begin
        _zz_2791_ = int_reg_array_19_49_imag;
        _zz_2792_ = int_reg_array_19_49_real;
      end
    endcase
  end

  always @(*) begin
    case(_zz_1102_)
      6'b000000 : begin
        _zz_2793_ = int_reg_array_20_0_imag;
        _zz_2794_ = int_reg_array_20_0_real;
      end
      6'b000001 : begin
        _zz_2793_ = int_reg_array_20_1_imag;
        _zz_2794_ = int_reg_array_20_1_real;
      end
      6'b000010 : begin
        _zz_2793_ = int_reg_array_20_2_imag;
        _zz_2794_ = int_reg_array_20_2_real;
      end
      6'b000011 : begin
        _zz_2793_ = int_reg_array_20_3_imag;
        _zz_2794_ = int_reg_array_20_3_real;
      end
      6'b000100 : begin
        _zz_2793_ = int_reg_array_20_4_imag;
        _zz_2794_ = int_reg_array_20_4_real;
      end
      6'b000101 : begin
        _zz_2793_ = int_reg_array_20_5_imag;
        _zz_2794_ = int_reg_array_20_5_real;
      end
      6'b000110 : begin
        _zz_2793_ = int_reg_array_20_6_imag;
        _zz_2794_ = int_reg_array_20_6_real;
      end
      6'b000111 : begin
        _zz_2793_ = int_reg_array_20_7_imag;
        _zz_2794_ = int_reg_array_20_7_real;
      end
      6'b001000 : begin
        _zz_2793_ = int_reg_array_20_8_imag;
        _zz_2794_ = int_reg_array_20_8_real;
      end
      6'b001001 : begin
        _zz_2793_ = int_reg_array_20_9_imag;
        _zz_2794_ = int_reg_array_20_9_real;
      end
      6'b001010 : begin
        _zz_2793_ = int_reg_array_20_10_imag;
        _zz_2794_ = int_reg_array_20_10_real;
      end
      6'b001011 : begin
        _zz_2793_ = int_reg_array_20_11_imag;
        _zz_2794_ = int_reg_array_20_11_real;
      end
      6'b001100 : begin
        _zz_2793_ = int_reg_array_20_12_imag;
        _zz_2794_ = int_reg_array_20_12_real;
      end
      6'b001101 : begin
        _zz_2793_ = int_reg_array_20_13_imag;
        _zz_2794_ = int_reg_array_20_13_real;
      end
      6'b001110 : begin
        _zz_2793_ = int_reg_array_20_14_imag;
        _zz_2794_ = int_reg_array_20_14_real;
      end
      6'b001111 : begin
        _zz_2793_ = int_reg_array_20_15_imag;
        _zz_2794_ = int_reg_array_20_15_real;
      end
      6'b010000 : begin
        _zz_2793_ = int_reg_array_20_16_imag;
        _zz_2794_ = int_reg_array_20_16_real;
      end
      6'b010001 : begin
        _zz_2793_ = int_reg_array_20_17_imag;
        _zz_2794_ = int_reg_array_20_17_real;
      end
      6'b010010 : begin
        _zz_2793_ = int_reg_array_20_18_imag;
        _zz_2794_ = int_reg_array_20_18_real;
      end
      6'b010011 : begin
        _zz_2793_ = int_reg_array_20_19_imag;
        _zz_2794_ = int_reg_array_20_19_real;
      end
      6'b010100 : begin
        _zz_2793_ = int_reg_array_20_20_imag;
        _zz_2794_ = int_reg_array_20_20_real;
      end
      6'b010101 : begin
        _zz_2793_ = int_reg_array_20_21_imag;
        _zz_2794_ = int_reg_array_20_21_real;
      end
      6'b010110 : begin
        _zz_2793_ = int_reg_array_20_22_imag;
        _zz_2794_ = int_reg_array_20_22_real;
      end
      6'b010111 : begin
        _zz_2793_ = int_reg_array_20_23_imag;
        _zz_2794_ = int_reg_array_20_23_real;
      end
      6'b011000 : begin
        _zz_2793_ = int_reg_array_20_24_imag;
        _zz_2794_ = int_reg_array_20_24_real;
      end
      6'b011001 : begin
        _zz_2793_ = int_reg_array_20_25_imag;
        _zz_2794_ = int_reg_array_20_25_real;
      end
      6'b011010 : begin
        _zz_2793_ = int_reg_array_20_26_imag;
        _zz_2794_ = int_reg_array_20_26_real;
      end
      6'b011011 : begin
        _zz_2793_ = int_reg_array_20_27_imag;
        _zz_2794_ = int_reg_array_20_27_real;
      end
      6'b011100 : begin
        _zz_2793_ = int_reg_array_20_28_imag;
        _zz_2794_ = int_reg_array_20_28_real;
      end
      6'b011101 : begin
        _zz_2793_ = int_reg_array_20_29_imag;
        _zz_2794_ = int_reg_array_20_29_real;
      end
      6'b011110 : begin
        _zz_2793_ = int_reg_array_20_30_imag;
        _zz_2794_ = int_reg_array_20_30_real;
      end
      6'b011111 : begin
        _zz_2793_ = int_reg_array_20_31_imag;
        _zz_2794_ = int_reg_array_20_31_real;
      end
      6'b100000 : begin
        _zz_2793_ = int_reg_array_20_32_imag;
        _zz_2794_ = int_reg_array_20_32_real;
      end
      6'b100001 : begin
        _zz_2793_ = int_reg_array_20_33_imag;
        _zz_2794_ = int_reg_array_20_33_real;
      end
      6'b100010 : begin
        _zz_2793_ = int_reg_array_20_34_imag;
        _zz_2794_ = int_reg_array_20_34_real;
      end
      6'b100011 : begin
        _zz_2793_ = int_reg_array_20_35_imag;
        _zz_2794_ = int_reg_array_20_35_real;
      end
      6'b100100 : begin
        _zz_2793_ = int_reg_array_20_36_imag;
        _zz_2794_ = int_reg_array_20_36_real;
      end
      6'b100101 : begin
        _zz_2793_ = int_reg_array_20_37_imag;
        _zz_2794_ = int_reg_array_20_37_real;
      end
      6'b100110 : begin
        _zz_2793_ = int_reg_array_20_38_imag;
        _zz_2794_ = int_reg_array_20_38_real;
      end
      6'b100111 : begin
        _zz_2793_ = int_reg_array_20_39_imag;
        _zz_2794_ = int_reg_array_20_39_real;
      end
      6'b101000 : begin
        _zz_2793_ = int_reg_array_20_40_imag;
        _zz_2794_ = int_reg_array_20_40_real;
      end
      6'b101001 : begin
        _zz_2793_ = int_reg_array_20_41_imag;
        _zz_2794_ = int_reg_array_20_41_real;
      end
      6'b101010 : begin
        _zz_2793_ = int_reg_array_20_42_imag;
        _zz_2794_ = int_reg_array_20_42_real;
      end
      6'b101011 : begin
        _zz_2793_ = int_reg_array_20_43_imag;
        _zz_2794_ = int_reg_array_20_43_real;
      end
      6'b101100 : begin
        _zz_2793_ = int_reg_array_20_44_imag;
        _zz_2794_ = int_reg_array_20_44_real;
      end
      6'b101101 : begin
        _zz_2793_ = int_reg_array_20_45_imag;
        _zz_2794_ = int_reg_array_20_45_real;
      end
      6'b101110 : begin
        _zz_2793_ = int_reg_array_20_46_imag;
        _zz_2794_ = int_reg_array_20_46_real;
      end
      6'b101111 : begin
        _zz_2793_ = int_reg_array_20_47_imag;
        _zz_2794_ = int_reg_array_20_47_real;
      end
      6'b110000 : begin
        _zz_2793_ = int_reg_array_20_48_imag;
        _zz_2794_ = int_reg_array_20_48_real;
      end
      default : begin
        _zz_2793_ = int_reg_array_20_49_imag;
        _zz_2794_ = int_reg_array_20_49_real;
      end
    endcase
  end

  always @(*) begin
    case(_zz_1157_)
      6'b000000 : begin
        _zz_2795_ = int_reg_array_21_0_imag;
        _zz_2796_ = int_reg_array_21_0_real;
      end
      6'b000001 : begin
        _zz_2795_ = int_reg_array_21_1_imag;
        _zz_2796_ = int_reg_array_21_1_real;
      end
      6'b000010 : begin
        _zz_2795_ = int_reg_array_21_2_imag;
        _zz_2796_ = int_reg_array_21_2_real;
      end
      6'b000011 : begin
        _zz_2795_ = int_reg_array_21_3_imag;
        _zz_2796_ = int_reg_array_21_3_real;
      end
      6'b000100 : begin
        _zz_2795_ = int_reg_array_21_4_imag;
        _zz_2796_ = int_reg_array_21_4_real;
      end
      6'b000101 : begin
        _zz_2795_ = int_reg_array_21_5_imag;
        _zz_2796_ = int_reg_array_21_5_real;
      end
      6'b000110 : begin
        _zz_2795_ = int_reg_array_21_6_imag;
        _zz_2796_ = int_reg_array_21_6_real;
      end
      6'b000111 : begin
        _zz_2795_ = int_reg_array_21_7_imag;
        _zz_2796_ = int_reg_array_21_7_real;
      end
      6'b001000 : begin
        _zz_2795_ = int_reg_array_21_8_imag;
        _zz_2796_ = int_reg_array_21_8_real;
      end
      6'b001001 : begin
        _zz_2795_ = int_reg_array_21_9_imag;
        _zz_2796_ = int_reg_array_21_9_real;
      end
      6'b001010 : begin
        _zz_2795_ = int_reg_array_21_10_imag;
        _zz_2796_ = int_reg_array_21_10_real;
      end
      6'b001011 : begin
        _zz_2795_ = int_reg_array_21_11_imag;
        _zz_2796_ = int_reg_array_21_11_real;
      end
      6'b001100 : begin
        _zz_2795_ = int_reg_array_21_12_imag;
        _zz_2796_ = int_reg_array_21_12_real;
      end
      6'b001101 : begin
        _zz_2795_ = int_reg_array_21_13_imag;
        _zz_2796_ = int_reg_array_21_13_real;
      end
      6'b001110 : begin
        _zz_2795_ = int_reg_array_21_14_imag;
        _zz_2796_ = int_reg_array_21_14_real;
      end
      6'b001111 : begin
        _zz_2795_ = int_reg_array_21_15_imag;
        _zz_2796_ = int_reg_array_21_15_real;
      end
      6'b010000 : begin
        _zz_2795_ = int_reg_array_21_16_imag;
        _zz_2796_ = int_reg_array_21_16_real;
      end
      6'b010001 : begin
        _zz_2795_ = int_reg_array_21_17_imag;
        _zz_2796_ = int_reg_array_21_17_real;
      end
      6'b010010 : begin
        _zz_2795_ = int_reg_array_21_18_imag;
        _zz_2796_ = int_reg_array_21_18_real;
      end
      6'b010011 : begin
        _zz_2795_ = int_reg_array_21_19_imag;
        _zz_2796_ = int_reg_array_21_19_real;
      end
      6'b010100 : begin
        _zz_2795_ = int_reg_array_21_20_imag;
        _zz_2796_ = int_reg_array_21_20_real;
      end
      6'b010101 : begin
        _zz_2795_ = int_reg_array_21_21_imag;
        _zz_2796_ = int_reg_array_21_21_real;
      end
      6'b010110 : begin
        _zz_2795_ = int_reg_array_21_22_imag;
        _zz_2796_ = int_reg_array_21_22_real;
      end
      6'b010111 : begin
        _zz_2795_ = int_reg_array_21_23_imag;
        _zz_2796_ = int_reg_array_21_23_real;
      end
      6'b011000 : begin
        _zz_2795_ = int_reg_array_21_24_imag;
        _zz_2796_ = int_reg_array_21_24_real;
      end
      6'b011001 : begin
        _zz_2795_ = int_reg_array_21_25_imag;
        _zz_2796_ = int_reg_array_21_25_real;
      end
      6'b011010 : begin
        _zz_2795_ = int_reg_array_21_26_imag;
        _zz_2796_ = int_reg_array_21_26_real;
      end
      6'b011011 : begin
        _zz_2795_ = int_reg_array_21_27_imag;
        _zz_2796_ = int_reg_array_21_27_real;
      end
      6'b011100 : begin
        _zz_2795_ = int_reg_array_21_28_imag;
        _zz_2796_ = int_reg_array_21_28_real;
      end
      6'b011101 : begin
        _zz_2795_ = int_reg_array_21_29_imag;
        _zz_2796_ = int_reg_array_21_29_real;
      end
      6'b011110 : begin
        _zz_2795_ = int_reg_array_21_30_imag;
        _zz_2796_ = int_reg_array_21_30_real;
      end
      6'b011111 : begin
        _zz_2795_ = int_reg_array_21_31_imag;
        _zz_2796_ = int_reg_array_21_31_real;
      end
      6'b100000 : begin
        _zz_2795_ = int_reg_array_21_32_imag;
        _zz_2796_ = int_reg_array_21_32_real;
      end
      6'b100001 : begin
        _zz_2795_ = int_reg_array_21_33_imag;
        _zz_2796_ = int_reg_array_21_33_real;
      end
      6'b100010 : begin
        _zz_2795_ = int_reg_array_21_34_imag;
        _zz_2796_ = int_reg_array_21_34_real;
      end
      6'b100011 : begin
        _zz_2795_ = int_reg_array_21_35_imag;
        _zz_2796_ = int_reg_array_21_35_real;
      end
      6'b100100 : begin
        _zz_2795_ = int_reg_array_21_36_imag;
        _zz_2796_ = int_reg_array_21_36_real;
      end
      6'b100101 : begin
        _zz_2795_ = int_reg_array_21_37_imag;
        _zz_2796_ = int_reg_array_21_37_real;
      end
      6'b100110 : begin
        _zz_2795_ = int_reg_array_21_38_imag;
        _zz_2796_ = int_reg_array_21_38_real;
      end
      6'b100111 : begin
        _zz_2795_ = int_reg_array_21_39_imag;
        _zz_2796_ = int_reg_array_21_39_real;
      end
      6'b101000 : begin
        _zz_2795_ = int_reg_array_21_40_imag;
        _zz_2796_ = int_reg_array_21_40_real;
      end
      6'b101001 : begin
        _zz_2795_ = int_reg_array_21_41_imag;
        _zz_2796_ = int_reg_array_21_41_real;
      end
      6'b101010 : begin
        _zz_2795_ = int_reg_array_21_42_imag;
        _zz_2796_ = int_reg_array_21_42_real;
      end
      6'b101011 : begin
        _zz_2795_ = int_reg_array_21_43_imag;
        _zz_2796_ = int_reg_array_21_43_real;
      end
      6'b101100 : begin
        _zz_2795_ = int_reg_array_21_44_imag;
        _zz_2796_ = int_reg_array_21_44_real;
      end
      6'b101101 : begin
        _zz_2795_ = int_reg_array_21_45_imag;
        _zz_2796_ = int_reg_array_21_45_real;
      end
      6'b101110 : begin
        _zz_2795_ = int_reg_array_21_46_imag;
        _zz_2796_ = int_reg_array_21_46_real;
      end
      6'b101111 : begin
        _zz_2795_ = int_reg_array_21_47_imag;
        _zz_2796_ = int_reg_array_21_47_real;
      end
      6'b110000 : begin
        _zz_2795_ = int_reg_array_21_48_imag;
        _zz_2796_ = int_reg_array_21_48_real;
      end
      default : begin
        _zz_2795_ = int_reg_array_21_49_imag;
        _zz_2796_ = int_reg_array_21_49_real;
      end
    endcase
  end

  always @(*) begin
    case(_zz_1212_)
      6'b000000 : begin
        _zz_2797_ = int_reg_array_22_0_imag;
        _zz_2798_ = int_reg_array_22_0_real;
      end
      6'b000001 : begin
        _zz_2797_ = int_reg_array_22_1_imag;
        _zz_2798_ = int_reg_array_22_1_real;
      end
      6'b000010 : begin
        _zz_2797_ = int_reg_array_22_2_imag;
        _zz_2798_ = int_reg_array_22_2_real;
      end
      6'b000011 : begin
        _zz_2797_ = int_reg_array_22_3_imag;
        _zz_2798_ = int_reg_array_22_3_real;
      end
      6'b000100 : begin
        _zz_2797_ = int_reg_array_22_4_imag;
        _zz_2798_ = int_reg_array_22_4_real;
      end
      6'b000101 : begin
        _zz_2797_ = int_reg_array_22_5_imag;
        _zz_2798_ = int_reg_array_22_5_real;
      end
      6'b000110 : begin
        _zz_2797_ = int_reg_array_22_6_imag;
        _zz_2798_ = int_reg_array_22_6_real;
      end
      6'b000111 : begin
        _zz_2797_ = int_reg_array_22_7_imag;
        _zz_2798_ = int_reg_array_22_7_real;
      end
      6'b001000 : begin
        _zz_2797_ = int_reg_array_22_8_imag;
        _zz_2798_ = int_reg_array_22_8_real;
      end
      6'b001001 : begin
        _zz_2797_ = int_reg_array_22_9_imag;
        _zz_2798_ = int_reg_array_22_9_real;
      end
      6'b001010 : begin
        _zz_2797_ = int_reg_array_22_10_imag;
        _zz_2798_ = int_reg_array_22_10_real;
      end
      6'b001011 : begin
        _zz_2797_ = int_reg_array_22_11_imag;
        _zz_2798_ = int_reg_array_22_11_real;
      end
      6'b001100 : begin
        _zz_2797_ = int_reg_array_22_12_imag;
        _zz_2798_ = int_reg_array_22_12_real;
      end
      6'b001101 : begin
        _zz_2797_ = int_reg_array_22_13_imag;
        _zz_2798_ = int_reg_array_22_13_real;
      end
      6'b001110 : begin
        _zz_2797_ = int_reg_array_22_14_imag;
        _zz_2798_ = int_reg_array_22_14_real;
      end
      6'b001111 : begin
        _zz_2797_ = int_reg_array_22_15_imag;
        _zz_2798_ = int_reg_array_22_15_real;
      end
      6'b010000 : begin
        _zz_2797_ = int_reg_array_22_16_imag;
        _zz_2798_ = int_reg_array_22_16_real;
      end
      6'b010001 : begin
        _zz_2797_ = int_reg_array_22_17_imag;
        _zz_2798_ = int_reg_array_22_17_real;
      end
      6'b010010 : begin
        _zz_2797_ = int_reg_array_22_18_imag;
        _zz_2798_ = int_reg_array_22_18_real;
      end
      6'b010011 : begin
        _zz_2797_ = int_reg_array_22_19_imag;
        _zz_2798_ = int_reg_array_22_19_real;
      end
      6'b010100 : begin
        _zz_2797_ = int_reg_array_22_20_imag;
        _zz_2798_ = int_reg_array_22_20_real;
      end
      6'b010101 : begin
        _zz_2797_ = int_reg_array_22_21_imag;
        _zz_2798_ = int_reg_array_22_21_real;
      end
      6'b010110 : begin
        _zz_2797_ = int_reg_array_22_22_imag;
        _zz_2798_ = int_reg_array_22_22_real;
      end
      6'b010111 : begin
        _zz_2797_ = int_reg_array_22_23_imag;
        _zz_2798_ = int_reg_array_22_23_real;
      end
      6'b011000 : begin
        _zz_2797_ = int_reg_array_22_24_imag;
        _zz_2798_ = int_reg_array_22_24_real;
      end
      6'b011001 : begin
        _zz_2797_ = int_reg_array_22_25_imag;
        _zz_2798_ = int_reg_array_22_25_real;
      end
      6'b011010 : begin
        _zz_2797_ = int_reg_array_22_26_imag;
        _zz_2798_ = int_reg_array_22_26_real;
      end
      6'b011011 : begin
        _zz_2797_ = int_reg_array_22_27_imag;
        _zz_2798_ = int_reg_array_22_27_real;
      end
      6'b011100 : begin
        _zz_2797_ = int_reg_array_22_28_imag;
        _zz_2798_ = int_reg_array_22_28_real;
      end
      6'b011101 : begin
        _zz_2797_ = int_reg_array_22_29_imag;
        _zz_2798_ = int_reg_array_22_29_real;
      end
      6'b011110 : begin
        _zz_2797_ = int_reg_array_22_30_imag;
        _zz_2798_ = int_reg_array_22_30_real;
      end
      6'b011111 : begin
        _zz_2797_ = int_reg_array_22_31_imag;
        _zz_2798_ = int_reg_array_22_31_real;
      end
      6'b100000 : begin
        _zz_2797_ = int_reg_array_22_32_imag;
        _zz_2798_ = int_reg_array_22_32_real;
      end
      6'b100001 : begin
        _zz_2797_ = int_reg_array_22_33_imag;
        _zz_2798_ = int_reg_array_22_33_real;
      end
      6'b100010 : begin
        _zz_2797_ = int_reg_array_22_34_imag;
        _zz_2798_ = int_reg_array_22_34_real;
      end
      6'b100011 : begin
        _zz_2797_ = int_reg_array_22_35_imag;
        _zz_2798_ = int_reg_array_22_35_real;
      end
      6'b100100 : begin
        _zz_2797_ = int_reg_array_22_36_imag;
        _zz_2798_ = int_reg_array_22_36_real;
      end
      6'b100101 : begin
        _zz_2797_ = int_reg_array_22_37_imag;
        _zz_2798_ = int_reg_array_22_37_real;
      end
      6'b100110 : begin
        _zz_2797_ = int_reg_array_22_38_imag;
        _zz_2798_ = int_reg_array_22_38_real;
      end
      6'b100111 : begin
        _zz_2797_ = int_reg_array_22_39_imag;
        _zz_2798_ = int_reg_array_22_39_real;
      end
      6'b101000 : begin
        _zz_2797_ = int_reg_array_22_40_imag;
        _zz_2798_ = int_reg_array_22_40_real;
      end
      6'b101001 : begin
        _zz_2797_ = int_reg_array_22_41_imag;
        _zz_2798_ = int_reg_array_22_41_real;
      end
      6'b101010 : begin
        _zz_2797_ = int_reg_array_22_42_imag;
        _zz_2798_ = int_reg_array_22_42_real;
      end
      6'b101011 : begin
        _zz_2797_ = int_reg_array_22_43_imag;
        _zz_2798_ = int_reg_array_22_43_real;
      end
      6'b101100 : begin
        _zz_2797_ = int_reg_array_22_44_imag;
        _zz_2798_ = int_reg_array_22_44_real;
      end
      6'b101101 : begin
        _zz_2797_ = int_reg_array_22_45_imag;
        _zz_2798_ = int_reg_array_22_45_real;
      end
      6'b101110 : begin
        _zz_2797_ = int_reg_array_22_46_imag;
        _zz_2798_ = int_reg_array_22_46_real;
      end
      6'b101111 : begin
        _zz_2797_ = int_reg_array_22_47_imag;
        _zz_2798_ = int_reg_array_22_47_real;
      end
      6'b110000 : begin
        _zz_2797_ = int_reg_array_22_48_imag;
        _zz_2798_ = int_reg_array_22_48_real;
      end
      default : begin
        _zz_2797_ = int_reg_array_22_49_imag;
        _zz_2798_ = int_reg_array_22_49_real;
      end
    endcase
  end

  always @(*) begin
    case(_zz_1267_)
      6'b000000 : begin
        _zz_2799_ = int_reg_array_23_0_imag;
        _zz_2800_ = int_reg_array_23_0_real;
      end
      6'b000001 : begin
        _zz_2799_ = int_reg_array_23_1_imag;
        _zz_2800_ = int_reg_array_23_1_real;
      end
      6'b000010 : begin
        _zz_2799_ = int_reg_array_23_2_imag;
        _zz_2800_ = int_reg_array_23_2_real;
      end
      6'b000011 : begin
        _zz_2799_ = int_reg_array_23_3_imag;
        _zz_2800_ = int_reg_array_23_3_real;
      end
      6'b000100 : begin
        _zz_2799_ = int_reg_array_23_4_imag;
        _zz_2800_ = int_reg_array_23_4_real;
      end
      6'b000101 : begin
        _zz_2799_ = int_reg_array_23_5_imag;
        _zz_2800_ = int_reg_array_23_5_real;
      end
      6'b000110 : begin
        _zz_2799_ = int_reg_array_23_6_imag;
        _zz_2800_ = int_reg_array_23_6_real;
      end
      6'b000111 : begin
        _zz_2799_ = int_reg_array_23_7_imag;
        _zz_2800_ = int_reg_array_23_7_real;
      end
      6'b001000 : begin
        _zz_2799_ = int_reg_array_23_8_imag;
        _zz_2800_ = int_reg_array_23_8_real;
      end
      6'b001001 : begin
        _zz_2799_ = int_reg_array_23_9_imag;
        _zz_2800_ = int_reg_array_23_9_real;
      end
      6'b001010 : begin
        _zz_2799_ = int_reg_array_23_10_imag;
        _zz_2800_ = int_reg_array_23_10_real;
      end
      6'b001011 : begin
        _zz_2799_ = int_reg_array_23_11_imag;
        _zz_2800_ = int_reg_array_23_11_real;
      end
      6'b001100 : begin
        _zz_2799_ = int_reg_array_23_12_imag;
        _zz_2800_ = int_reg_array_23_12_real;
      end
      6'b001101 : begin
        _zz_2799_ = int_reg_array_23_13_imag;
        _zz_2800_ = int_reg_array_23_13_real;
      end
      6'b001110 : begin
        _zz_2799_ = int_reg_array_23_14_imag;
        _zz_2800_ = int_reg_array_23_14_real;
      end
      6'b001111 : begin
        _zz_2799_ = int_reg_array_23_15_imag;
        _zz_2800_ = int_reg_array_23_15_real;
      end
      6'b010000 : begin
        _zz_2799_ = int_reg_array_23_16_imag;
        _zz_2800_ = int_reg_array_23_16_real;
      end
      6'b010001 : begin
        _zz_2799_ = int_reg_array_23_17_imag;
        _zz_2800_ = int_reg_array_23_17_real;
      end
      6'b010010 : begin
        _zz_2799_ = int_reg_array_23_18_imag;
        _zz_2800_ = int_reg_array_23_18_real;
      end
      6'b010011 : begin
        _zz_2799_ = int_reg_array_23_19_imag;
        _zz_2800_ = int_reg_array_23_19_real;
      end
      6'b010100 : begin
        _zz_2799_ = int_reg_array_23_20_imag;
        _zz_2800_ = int_reg_array_23_20_real;
      end
      6'b010101 : begin
        _zz_2799_ = int_reg_array_23_21_imag;
        _zz_2800_ = int_reg_array_23_21_real;
      end
      6'b010110 : begin
        _zz_2799_ = int_reg_array_23_22_imag;
        _zz_2800_ = int_reg_array_23_22_real;
      end
      6'b010111 : begin
        _zz_2799_ = int_reg_array_23_23_imag;
        _zz_2800_ = int_reg_array_23_23_real;
      end
      6'b011000 : begin
        _zz_2799_ = int_reg_array_23_24_imag;
        _zz_2800_ = int_reg_array_23_24_real;
      end
      6'b011001 : begin
        _zz_2799_ = int_reg_array_23_25_imag;
        _zz_2800_ = int_reg_array_23_25_real;
      end
      6'b011010 : begin
        _zz_2799_ = int_reg_array_23_26_imag;
        _zz_2800_ = int_reg_array_23_26_real;
      end
      6'b011011 : begin
        _zz_2799_ = int_reg_array_23_27_imag;
        _zz_2800_ = int_reg_array_23_27_real;
      end
      6'b011100 : begin
        _zz_2799_ = int_reg_array_23_28_imag;
        _zz_2800_ = int_reg_array_23_28_real;
      end
      6'b011101 : begin
        _zz_2799_ = int_reg_array_23_29_imag;
        _zz_2800_ = int_reg_array_23_29_real;
      end
      6'b011110 : begin
        _zz_2799_ = int_reg_array_23_30_imag;
        _zz_2800_ = int_reg_array_23_30_real;
      end
      6'b011111 : begin
        _zz_2799_ = int_reg_array_23_31_imag;
        _zz_2800_ = int_reg_array_23_31_real;
      end
      6'b100000 : begin
        _zz_2799_ = int_reg_array_23_32_imag;
        _zz_2800_ = int_reg_array_23_32_real;
      end
      6'b100001 : begin
        _zz_2799_ = int_reg_array_23_33_imag;
        _zz_2800_ = int_reg_array_23_33_real;
      end
      6'b100010 : begin
        _zz_2799_ = int_reg_array_23_34_imag;
        _zz_2800_ = int_reg_array_23_34_real;
      end
      6'b100011 : begin
        _zz_2799_ = int_reg_array_23_35_imag;
        _zz_2800_ = int_reg_array_23_35_real;
      end
      6'b100100 : begin
        _zz_2799_ = int_reg_array_23_36_imag;
        _zz_2800_ = int_reg_array_23_36_real;
      end
      6'b100101 : begin
        _zz_2799_ = int_reg_array_23_37_imag;
        _zz_2800_ = int_reg_array_23_37_real;
      end
      6'b100110 : begin
        _zz_2799_ = int_reg_array_23_38_imag;
        _zz_2800_ = int_reg_array_23_38_real;
      end
      6'b100111 : begin
        _zz_2799_ = int_reg_array_23_39_imag;
        _zz_2800_ = int_reg_array_23_39_real;
      end
      6'b101000 : begin
        _zz_2799_ = int_reg_array_23_40_imag;
        _zz_2800_ = int_reg_array_23_40_real;
      end
      6'b101001 : begin
        _zz_2799_ = int_reg_array_23_41_imag;
        _zz_2800_ = int_reg_array_23_41_real;
      end
      6'b101010 : begin
        _zz_2799_ = int_reg_array_23_42_imag;
        _zz_2800_ = int_reg_array_23_42_real;
      end
      6'b101011 : begin
        _zz_2799_ = int_reg_array_23_43_imag;
        _zz_2800_ = int_reg_array_23_43_real;
      end
      6'b101100 : begin
        _zz_2799_ = int_reg_array_23_44_imag;
        _zz_2800_ = int_reg_array_23_44_real;
      end
      6'b101101 : begin
        _zz_2799_ = int_reg_array_23_45_imag;
        _zz_2800_ = int_reg_array_23_45_real;
      end
      6'b101110 : begin
        _zz_2799_ = int_reg_array_23_46_imag;
        _zz_2800_ = int_reg_array_23_46_real;
      end
      6'b101111 : begin
        _zz_2799_ = int_reg_array_23_47_imag;
        _zz_2800_ = int_reg_array_23_47_real;
      end
      6'b110000 : begin
        _zz_2799_ = int_reg_array_23_48_imag;
        _zz_2800_ = int_reg_array_23_48_real;
      end
      default : begin
        _zz_2799_ = int_reg_array_23_49_imag;
        _zz_2800_ = int_reg_array_23_49_real;
      end
    endcase
  end

  always @(*) begin
    case(_zz_1322_)
      6'b000000 : begin
        _zz_2801_ = int_reg_array_24_0_imag;
        _zz_2802_ = int_reg_array_24_0_real;
      end
      6'b000001 : begin
        _zz_2801_ = int_reg_array_24_1_imag;
        _zz_2802_ = int_reg_array_24_1_real;
      end
      6'b000010 : begin
        _zz_2801_ = int_reg_array_24_2_imag;
        _zz_2802_ = int_reg_array_24_2_real;
      end
      6'b000011 : begin
        _zz_2801_ = int_reg_array_24_3_imag;
        _zz_2802_ = int_reg_array_24_3_real;
      end
      6'b000100 : begin
        _zz_2801_ = int_reg_array_24_4_imag;
        _zz_2802_ = int_reg_array_24_4_real;
      end
      6'b000101 : begin
        _zz_2801_ = int_reg_array_24_5_imag;
        _zz_2802_ = int_reg_array_24_5_real;
      end
      6'b000110 : begin
        _zz_2801_ = int_reg_array_24_6_imag;
        _zz_2802_ = int_reg_array_24_6_real;
      end
      6'b000111 : begin
        _zz_2801_ = int_reg_array_24_7_imag;
        _zz_2802_ = int_reg_array_24_7_real;
      end
      6'b001000 : begin
        _zz_2801_ = int_reg_array_24_8_imag;
        _zz_2802_ = int_reg_array_24_8_real;
      end
      6'b001001 : begin
        _zz_2801_ = int_reg_array_24_9_imag;
        _zz_2802_ = int_reg_array_24_9_real;
      end
      6'b001010 : begin
        _zz_2801_ = int_reg_array_24_10_imag;
        _zz_2802_ = int_reg_array_24_10_real;
      end
      6'b001011 : begin
        _zz_2801_ = int_reg_array_24_11_imag;
        _zz_2802_ = int_reg_array_24_11_real;
      end
      6'b001100 : begin
        _zz_2801_ = int_reg_array_24_12_imag;
        _zz_2802_ = int_reg_array_24_12_real;
      end
      6'b001101 : begin
        _zz_2801_ = int_reg_array_24_13_imag;
        _zz_2802_ = int_reg_array_24_13_real;
      end
      6'b001110 : begin
        _zz_2801_ = int_reg_array_24_14_imag;
        _zz_2802_ = int_reg_array_24_14_real;
      end
      6'b001111 : begin
        _zz_2801_ = int_reg_array_24_15_imag;
        _zz_2802_ = int_reg_array_24_15_real;
      end
      6'b010000 : begin
        _zz_2801_ = int_reg_array_24_16_imag;
        _zz_2802_ = int_reg_array_24_16_real;
      end
      6'b010001 : begin
        _zz_2801_ = int_reg_array_24_17_imag;
        _zz_2802_ = int_reg_array_24_17_real;
      end
      6'b010010 : begin
        _zz_2801_ = int_reg_array_24_18_imag;
        _zz_2802_ = int_reg_array_24_18_real;
      end
      6'b010011 : begin
        _zz_2801_ = int_reg_array_24_19_imag;
        _zz_2802_ = int_reg_array_24_19_real;
      end
      6'b010100 : begin
        _zz_2801_ = int_reg_array_24_20_imag;
        _zz_2802_ = int_reg_array_24_20_real;
      end
      6'b010101 : begin
        _zz_2801_ = int_reg_array_24_21_imag;
        _zz_2802_ = int_reg_array_24_21_real;
      end
      6'b010110 : begin
        _zz_2801_ = int_reg_array_24_22_imag;
        _zz_2802_ = int_reg_array_24_22_real;
      end
      6'b010111 : begin
        _zz_2801_ = int_reg_array_24_23_imag;
        _zz_2802_ = int_reg_array_24_23_real;
      end
      6'b011000 : begin
        _zz_2801_ = int_reg_array_24_24_imag;
        _zz_2802_ = int_reg_array_24_24_real;
      end
      6'b011001 : begin
        _zz_2801_ = int_reg_array_24_25_imag;
        _zz_2802_ = int_reg_array_24_25_real;
      end
      6'b011010 : begin
        _zz_2801_ = int_reg_array_24_26_imag;
        _zz_2802_ = int_reg_array_24_26_real;
      end
      6'b011011 : begin
        _zz_2801_ = int_reg_array_24_27_imag;
        _zz_2802_ = int_reg_array_24_27_real;
      end
      6'b011100 : begin
        _zz_2801_ = int_reg_array_24_28_imag;
        _zz_2802_ = int_reg_array_24_28_real;
      end
      6'b011101 : begin
        _zz_2801_ = int_reg_array_24_29_imag;
        _zz_2802_ = int_reg_array_24_29_real;
      end
      6'b011110 : begin
        _zz_2801_ = int_reg_array_24_30_imag;
        _zz_2802_ = int_reg_array_24_30_real;
      end
      6'b011111 : begin
        _zz_2801_ = int_reg_array_24_31_imag;
        _zz_2802_ = int_reg_array_24_31_real;
      end
      6'b100000 : begin
        _zz_2801_ = int_reg_array_24_32_imag;
        _zz_2802_ = int_reg_array_24_32_real;
      end
      6'b100001 : begin
        _zz_2801_ = int_reg_array_24_33_imag;
        _zz_2802_ = int_reg_array_24_33_real;
      end
      6'b100010 : begin
        _zz_2801_ = int_reg_array_24_34_imag;
        _zz_2802_ = int_reg_array_24_34_real;
      end
      6'b100011 : begin
        _zz_2801_ = int_reg_array_24_35_imag;
        _zz_2802_ = int_reg_array_24_35_real;
      end
      6'b100100 : begin
        _zz_2801_ = int_reg_array_24_36_imag;
        _zz_2802_ = int_reg_array_24_36_real;
      end
      6'b100101 : begin
        _zz_2801_ = int_reg_array_24_37_imag;
        _zz_2802_ = int_reg_array_24_37_real;
      end
      6'b100110 : begin
        _zz_2801_ = int_reg_array_24_38_imag;
        _zz_2802_ = int_reg_array_24_38_real;
      end
      6'b100111 : begin
        _zz_2801_ = int_reg_array_24_39_imag;
        _zz_2802_ = int_reg_array_24_39_real;
      end
      6'b101000 : begin
        _zz_2801_ = int_reg_array_24_40_imag;
        _zz_2802_ = int_reg_array_24_40_real;
      end
      6'b101001 : begin
        _zz_2801_ = int_reg_array_24_41_imag;
        _zz_2802_ = int_reg_array_24_41_real;
      end
      6'b101010 : begin
        _zz_2801_ = int_reg_array_24_42_imag;
        _zz_2802_ = int_reg_array_24_42_real;
      end
      6'b101011 : begin
        _zz_2801_ = int_reg_array_24_43_imag;
        _zz_2802_ = int_reg_array_24_43_real;
      end
      6'b101100 : begin
        _zz_2801_ = int_reg_array_24_44_imag;
        _zz_2802_ = int_reg_array_24_44_real;
      end
      6'b101101 : begin
        _zz_2801_ = int_reg_array_24_45_imag;
        _zz_2802_ = int_reg_array_24_45_real;
      end
      6'b101110 : begin
        _zz_2801_ = int_reg_array_24_46_imag;
        _zz_2802_ = int_reg_array_24_46_real;
      end
      6'b101111 : begin
        _zz_2801_ = int_reg_array_24_47_imag;
        _zz_2802_ = int_reg_array_24_47_real;
      end
      6'b110000 : begin
        _zz_2801_ = int_reg_array_24_48_imag;
        _zz_2802_ = int_reg_array_24_48_real;
      end
      default : begin
        _zz_2801_ = int_reg_array_24_49_imag;
        _zz_2802_ = int_reg_array_24_49_real;
      end
    endcase
  end

  always @(*) begin
    case(_zz_1377_)
      6'b000000 : begin
        _zz_2803_ = int_reg_array_25_0_imag;
        _zz_2804_ = int_reg_array_25_0_real;
      end
      6'b000001 : begin
        _zz_2803_ = int_reg_array_25_1_imag;
        _zz_2804_ = int_reg_array_25_1_real;
      end
      6'b000010 : begin
        _zz_2803_ = int_reg_array_25_2_imag;
        _zz_2804_ = int_reg_array_25_2_real;
      end
      6'b000011 : begin
        _zz_2803_ = int_reg_array_25_3_imag;
        _zz_2804_ = int_reg_array_25_3_real;
      end
      6'b000100 : begin
        _zz_2803_ = int_reg_array_25_4_imag;
        _zz_2804_ = int_reg_array_25_4_real;
      end
      6'b000101 : begin
        _zz_2803_ = int_reg_array_25_5_imag;
        _zz_2804_ = int_reg_array_25_5_real;
      end
      6'b000110 : begin
        _zz_2803_ = int_reg_array_25_6_imag;
        _zz_2804_ = int_reg_array_25_6_real;
      end
      6'b000111 : begin
        _zz_2803_ = int_reg_array_25_7_imag;
        _zz_2804_ = int_reg_array_25_7_real;
      end
      6'b001000 : begin
        _zz_2803_ = int_reg_array_25_8_imag;
        _zz_2804_ = int_reg_array_25_8_real;
      end
      6'b001001 : begin
        _zz_2803_ = int_reg_array_25_9_imag;
        _zz_2804_ = int_reg_array_25_9_real;
      end
      6'b001010 : begin
        _zz_2803_ = int_reg_array_25_10_imag;
        _zz_2804_ = int_reg_array_25_10_real;
      end
      6'b001011 : begin
        _zz_2803_ = int_reg_array_25_11_imag;
        _zz_2804_ = int_reg_array_25_11_real;
      end
      6'b001100 : begin
        _zz_2803_ = int_reg_array_25_12_imag;
        _zz_2804_ = int_reg_array_25_12_real;
      end
      6'b001101 : begin
        _zz_2803_ = int_reg_array_25_13_imag;
        _zz_2804_ = int_reg_array_25_13_real;
      end
      6'b001110 : begin
        _zz_2803_ = int_reg_array_25_14_imag;
        _zz_2804_ = int_reg_array_25_14_real;
      end
      6'b001111 : begin
        _zz_2803_ = int_reg_array_25_15_imag;
        _zz_2804_ = int_reg_array_25_15_real;
      end
      6'b010000 : begin
        _zz_2803_ = int_reg_array_25_16_imag;
        _zz_2804_ = int_reg_array_25_16_real;
      end
      6'b010001 : begin
        _zz_2803_ = int_reg_array_25_17_imag;
        _zz_2804_ = int_reg_array_25_17_real;
      end
      6'b010010 : begin
        _zz_2803_ = int_reg_array_25_18_imag;
        _zz_2804_ = int_reg_array_25_18_real;
      end
      6'b010011 : begin
        _zz_2803_ = int_reg_array_25_19_imag;
        _zz_2804_ = int_reg_array_25_19_real;
      end
      6'b010100 : begin
        _zz_2803_ = int_reg_array_25_20_imag;
        _zz_2804_ = int_reg_array_25_20_real;
      end
      6'b010101 : begin
        _zz_2803_ = int_reg_array_25_21_imag;
        _zz_2804_ = int_reg_array_25_21_real;
      end
      6'b010110 : begin
        _zz_2803_ = int_reg_array_25_22_imag;
        _zz_2804_ = int_reg_array_25_22_real;
      end
      6'b010111 : begin
        _zz_2803_ = int_reg_array_25_23_imag;
        _zz_2804_ = int_reg_array_25_23_real;
      end
      6'b011000 : begin
        _zz_2803_ = int_reg_array_25_24_imag;
        _zz_2804_ = int_reg_array_25_24_real;
      end
      6'b011001 : begin
        _zz_2803_ = int_reg_array_25_25_imag;
        _zz_2804_ = int_reg_array_25_25_real;
      end
      6'b011010 : begin
        _zz_2803_ = int_reg_array_25_26_imag;
        _zz_2804_ = int_reg_array_25_26_real;
      end
      6'b011011 : begin
        _zz_2803_ = int_reg_array_25_27_imag;
        _zz_2804_ = int_reg_array_25_27_real;
      end
      6'b011100 : begin
        _zz_2803_ = int_reg_array_25_28_imag;
        _zz_2804_ = int_reg_array_25_28_real;
      end
      6'b011101 : begin
        _zz_2803_ = int_reg_array_25_29_imag;
        _zz_2804_ = int_reg_array_25_29_real;
      end
      6'b011110 : begin
        _zz_2803_ = int_reg_array_25_30_imag;
        _zz_2804_ = int_reg_array_25_30_real;
      end
      6'b011111 : begin
        _zz_2803_ = int_reg_array_25_31_imag;
        _zz_2804_ = int_reg_array_25_31_real;
      end
      6'b100000 : begin
        _zz_2803_ = int_reg_array_25_32_imag;
        _zz_2804_ = int_reg_array_25_32_real;
      end
      6'b100001 : begin
        _zz_2803_ = int_reg_array_25_33_imag;
        _zz_2804_ = int_reg_array_25_33_real;
      end
      6'b100010 : begin
        _zz_2803_ = int_reg_array_25_34_imag;
        _zz_2804_ = int_reg_array_25_34_real;
      end
      6'b100011 : begin
        _zz_2803_ = int_reg_array_25_35_imag;
        _zz_2804_ = int_reg_array_25_35_real;
      end
      6'b100100 : begin
        _zz_2803_ = int_reg_array_25_36_imag;
        _zz_2804_ = int_reg_array_25_36_real;
      end
      6'b100101 : begin
        _zz_2803_ = int_reg_array_25_37_imag;
        _zz_2804_ = int_reg_array_25_37_real;
      end
      6'b100110 : begin
        _zz_2803_ = int_reg_array_25_38_imag;
        _zz_2804_ = int_reg_array_25_38_real;
      end
      6'b100111 : begin
        _zz_2803_ = int_reg_array_25_39_imag;
        _zz_2804_ = int_reg_array_25_39_real;
      end
      6'b101000 : begin
        _zz_2803_ = int_reg_array_25_40_imag;
        _zz_2804_ = int_reg_array_25_40_real;
      end
      6'b101001 : begin
        _zz_2803_ = int_reg_array_25_41_imag;
        _zz_2804_ = int_reg_array_25_41_real;
      end
      6'b101010 : begin
        _zz_2803_ = int_reg_array_25_42_imag;
        _zz_2804_ = int_reg_array_25_42_real;
      end
      6'b101011 : begin
        _zz_2803_ = int_reg_array_25_43_imag;
        _zz_2804_ = int_reg_array_25_43_real;
      end
      6'b101100 : begin
        _zz_2803_ = int_reg_array_25_44_imag;
        _zz_2804_ = int_reg_array_25_44_real;
      end
      6'b101101 : begin
        _zz_2803_ = int_reg_array_25_45_imag;
        _zz_2804_ = int_reg_array_25_45_real;
      end
      6'b101110 : begin
        _zz_2803_ = int_reg_array_25_46_imag;
        _zz_2804_ = int_reg_array_25_46_real;
      end
      6'b101111 : begin
        _zz_2803_ = int_reg_array_25_47_imag;
        _zz_2804_ = int_reg_array_25_47_real;
      end
      6'b110000 : begin
        _zz_2803_ = int_reg_array_25_48_imag;
        _zz_2804_ = int_reg_array_25_48_real;
      end
      default : begin
        _zz_2803_ = int_reg_array_25_49_imag;
        _zz_2804_ = int_reg_array_25_49_real;
      end
    endcase
  end

  always @(*) begin
    case(_zz_1432_)
      6'b000000 : begin
        _zz_2805_ = int_reg_array_26_0_imag;
        _zz_2806_ = int_reg_array_26_0_real;
      end
      6'b000001 : begin
        _zz_2805_ = int_reg_array_26_1_imag;
        _zz_2806_ = int_reg_array_26_1_real;
      end
      6'b000010 : begin
        _zz_2805_ = int_reg_array_26_2_imag;
        _zz_2806_ = int_reg_array_26_2_real;
      end
      6'b000011 : begin
        _zz_2805_ = int_reg_array_26_3_imag;
        _zz_2806_ = int_reg_array_26_3_real;
      end
      6'b000100 : begin
        _zz_2805_ = int_reg_array_26_4_imag;
        _zz_2806_ = int_reg_array_26_4_real;
      end
      6'b000101 : begin
        _zz_2805_ = int_reg_array_26_5_imag;
        _zz_2806_ = int_reg_array_26_5_real;
      end
      6'b000110 : begin
        _zz_2805_ = int_reg_array_26_6_imag;
        _zz_2806_ = int_reg_array_26_6_real;
      end
      6'b000111 : begin
        _zz_2805_ = int_reg_array_26_7_imag;
        _zz_2806_ = int_reg_array_26_7_real;
      end
      6'b001000 : begin
        _zz_2805_ = int_reg_array_26_8_imag;
        _zz_2806_ = int_reg_array_26_8_real;
      end
      6'b001001 : begin
        _zz_2805_ = int_reg_array_26_9_imag;
        _zz_2806_ = int_reg_array_26_9_real;
      end
      6'b001010 : begin
        _zz_2805_ = int_reg_array_26_10_imag;
        _zz_2806_ = int_reg_array_26_10_real;
      end
      6'b001011 : begin
        _zz_2805_ = int_reg_array_26_11_imag;
        _zz_2806_ = int_reg_array_26_11_real;
      end
      6'b001100 : begin
        _zz_2805_ = int_reg_array_26_12_imag;
        _zz_2806_ = int_reg_array_26_12_real;
      end
      6'b001101 : begin
        _zz_2805_ = int_reg_array_26_13_imag;
        _zz_2806_ = int_reg_array_26_13_real;
      end
      6'b001110 : begin
        _zz_2805_ = int_reg_array_26_14_imag;
        _zz_2806_ = int_reg_array_26_14_real;
      end
      6'b001111 : begin
        _zz_2805_ = int_reg_array_26_15_imag;
        _zz_2806_ = int_reg_array_26_15_real;
      end
      6'b010000 : begin
        _zz_2805_ = int_reg_array_26_16_imag;
        _zz_2806_ = int_reg_array_26_16_real;
      end
      6'b010001 : begin
        _zz_2805_ = int_reg_array_26_17_imag;
        _zz_2806_ = int_reg_array_26_17_real;
      end
      6'b010010 : begin
        _zz_2805_ = int_reg_array_26_18_imag;
        _zz_2806_ = int_reg_array_26_18_real;
      end
      6'b010011 : begin
        _zz_2805_ = int_reg_array_26_19_imag;
        _zz_2806_ = int_reg_array_26_19_real;
      end
      6'b010100 : begin
        _zz_2805_ = int_reg_array_26_20_imag;
        _zz_2806_ = int_reg_array_26_20_real;
      end
      6'b010101 : begin
        _zz_2805_ = int_reg_array_26_21_imag;
        _zz_2806_ = int_reg_array_26_21_real;
      end
      6'b010110 : begin
        _zz_2805_ = int_reg_array_26_22_imag;
        _zz_2806_ = int_reg_array_26_22_real;
      end
      6'b010111 : begin
        _zz_2805_ = int_reg_array_26_23_imag;
        _zz_2806_ = int_reg_array_26_23_real;
      end
      6'b011000 : begin
        _zz_2805_ = int_reg_array_26_24_imag;
        _zz_2806_ = int_reg_array_26_24_real;
      end
      6'b011001 : begin
        _zz_2805_ = int_reg_array_26_25_imag;
        _zz_2806_ = int_reg_array_26_25_real;
      end
      6'b011010 : begin
        _zz_2805_ = int_reg_array_26_26_imag;
        _zz_2806_ = int_reg_array_26_26_real;
      end
      6'b011011 : begin
        _zz_2805_ = int_reg_array_26_27_imag;
        _zz_2806_ = int_reg_array_26_27_real;
      end
      6'b011100 : begin
        _zz_2805_ = int_reg_array_26_28_imag;
        _zz_2806_ = int_reg_array_26_28_real;
      end
      6'b011101 : begin
        _zz_2805_ = int_reg_array_26_29_imag;
        _zz_2806_ = int_reg_array_26_29_real;
      end
      6'b011110 : begin
        _zz_2805_ = int_reg_array_26_30_imag;
        _zz_2806_ = int_reg_array_26_30_real;
      end
      6'b011111 : begin
        _zz_2805_ = int_reg_array_26_31_imag;
        _zz_2806_ = int_reg_array_26_31_real;
      end
      6'b100000 : begin
        _zz_2805_ = int_reg_array_26_32_imag;
        _zz_2806_ = int_reg_array_26_32_real;
      end
      6'b100001 : begin
        _zz_2805_ = int_reg_array_26_33_imag;
        _zz_2806_ = int_reg_array_26_33_real;
      end
      6'b100010 : begin
        _zz_2805_ = int_reg_array_26_34_imag;
        _zz_2806_ = int_reg_array_26_34_real;
      end
      6'b100011 : begin
        _zz_2805_ = int_reg_array_26_35_imag;
        _zz_2806_ = int_reg_array_26_35_real;
      end
      6'b100100 : begin
        _zz_2805_ = int_reg_array_26_36_imag;
        _zz_2806_ = int_reg_array_26_36_real;
      end
      6'b100101 : begin
        _zz_2805_ = int_reg_array_26_37_imag;
        _zz_2806_ = int_reg_array_26_37_real;
      end
      6'b100110 : begin
        _zz_2805_ = int_reg_array_26_38_imag;
        _zz_2806_ = int_reg_array_26_38_real;
      end
      6'b100111 : begin
        _zz_2805_ = int_reg_array_26_39_imag;
        _zz_2806_ = int_reg_array_26_39_real;
      end
      6'b101000 : begin
        _zz_2805_ = int_reg_array_26_40_imag;
        _zz_2806_ = int_reg_array_26_40_real;
      end
      6'b101001 : begin
        _zz_2805_ = int_reg_array_26_41_imag;
        _zz_2806_ = int_reg_array_26_41_real;
      end
      6'b101010 : begin
        _zz_2805_ = int_reg_array_26_42_imag;
        _zz_2806_ = int_reg_array_26_42_real;
      end
      6'b101011 : begin
        _zz_2805_ = int_reg_array_26_43_imag;
        _zz_2806_ = int_reg_array_26_43_real;
      end
      6'b101100 : begin
        _zz_2805_ = int_reg_array_26_44_imag;
        _zz_2806_ = int_reg_array_26_44_real;
      end
      6'b101101 : begin
        _zz_2805_ = int_reg_array_26_45_imag;
        _zz_2806_ = int_reg_array_26_45_real;
      end
      6'b101110 : begin
        _zz_2805_ = int_reg_array_26_46_imag;
        _zz_2806_ = int_reg_array_26_46_real;
      end
      6'b101111 : begin
        _zz_2805_ = int_reg_array_26_47_imag;
        _zz_2806_ = int_reg_array_26_47_real;
      end
      6'b110000 : begin
        _zz_2805_ = int_reg_array_26_48_imag;
        _zz_2806_ = int_reg_array_26_48_real;
      end
      default : begin
        _zz_2805_ = int_reg_array_26_49_imag;
        _zz_2806_ = int_reg_array_26_49_real;
      end
    endcase
  end

  always @(*) begin
    case(_zz_1487_)
      6'b000000 : begin
        _zz_2807_ = int_reg_array_27_0_imag;
        _zz_2808_ = int_reg_array_27_0_real;
      end
      6'b000001 : begin
        _zz_2807_ = int_reg_array_27_1_imag;
        _zz_2808_ = int_reg_array_27_1_real;
      end
      6'b000010 : begin
        _zz_2807_ = int_reg_array_27_2_imag;
        _zz_2808_ = int_reg_array_27_2_real;
      end
      6'b000011 : begin
        _zz_2807_ = int_reg_array_27_3_imag;
        _zz_2808_ = int_reg_array_27_3_real;
      end
      6'b000100 : begin
        _zz_2807_ = int_reg_array_27_4_imag;
        _zz_2808_ = int_reg_array_27_4_real;
      end
      6'b000101 : begin
        _zz_2807_ = int_reg_array_27_5_imag;
        _zz_2808_ = int_reg_array_27_5_real;
      end
      6'b000110 : begin
        _zz_2807_ = int_reg_array_27_6_imag;
        _zz_2808_ = int_reg_array_27_6_real;
      end
      6'b000111 : begin
        _zz_2807_ = int_reg_array_27_7_imag;
        _zz_2808_ = int_reg_array_27_7_real;
      end
      6'b001000 : begin
        _zz_2807_ = int_reg_array_27_8_imag;
        _zz_2808_ = int_reg_array_27_8_real;
      end
      6'b001001 : begin
        _zz_2807_ = int_reg_array_27_9_imag;
        _zz_2808_ = int_reg_array_27_9_real;
      end
      6'b001010 : begin
        _zz_2807_ = int_reg_array_27_10_imag;
        _zz_2808_ = int_reg_array_27_10_real;
      end
      6'b001011 : begin
        _zz_2807_ = int_reg_array_27_11_imag;
        _zz_2808_ = int_reg_array_27_11_real;
      end
      6'b001100 : begin
        _zz_2807_ = int_reg_array_27_12_imag;
        _zz_2808_ = int_reg_array_27_12_real;
      end
      6'b001101 : begin
        _zz_2807_ = int_reg_array_27_13_imag;
        _zz_2808_ = int_reg_array_27_13_real;
      end
      6'b001110 : begin
        _zz_2807_ = int_reg_array_27_14_imag;
        _zz_2808_ = int_reg_array_27_14_real;
      end
      6'b001111 : begin
        _zz_2807_ = int_reg_array_27_15_imag;
        _zz_2808_ = int_reg_array_27_15_real;
      end
      6'b010000 : begin
        _zz_2807_ = int_reg_array_27_16_imag;
        _zz_2808_ = int_reg_array_27_16_real;
      end
      6'b010001 : begin
        _zz_2807_ = int_reg_array_27_17_imag;
        _zz_2808_ = int_reg_array_27_17_real;
      end
      6'b010010 : begin
        _zz_2807_ = int_reg_array_27_18_imag;
        _zz_2808_ = int_reg_array_27_18_real;
      end
      6'b010011 : begin
        _zz_2807_ = int_reg_array_27_19_imag;
        _zz_2808_ = int_reg_array_27_19_real;
      end
      6'b010100 : begin
        _zz_2807_ = int_reg_array_27_20_imag;
        _zz_2808_ = int_reg_array_27_20_real;
      end
      6'b010101 : begin
        _zz_2807_ = int_reg_array_27_21_imag;
        _zz_2808_ = int_reg_array_27_21_real;
      end
      6'b010110 : begin
        _zz_2807_ = int_reg_array_27_22_imag;
        _zz_2808_ = int_reg_array_27_22_real;
      end
      6'b010111 : begin
        _zz_2807_ = int_reg_array_27_23_imag;
        _zz_2808_ = int_reg_array_27_23_real;
      end
      6'b011000 : begin
        _zz_2807_ = int_reg_array_27_24_imag;
        _zz_2808_ = int_reg_array_27_24_real;
      end
      6'b011001 : begin
        _zz_2807_ = int_reg_array_27_25_imag;
        _zz_2808_ = int_reg_array_27_25_real;
      end
      6'b011010 : begin
        _zz_2807_ = int_reg_array_27_26_imag;
        _zz_2808_ = int_reg_array_27_26_real;
      end
      6'b011011 : begin
        _zz_2807_ = int_reg_array_27_27_imag;
        _zz_2808_ = int_reg_array_27_27_real;
      end
      6'b011100 : begin
        _zz_2807_ = int_reg_array_27_28_imag;
        _zz_2808_ = int_reg_array_27_28_real;
      end
      6'b011101 : begin
        _zz_2807_ = int_reg_array_27_29_imag;
        _zz_2808_ = int_reg_array_27_29_real;
      end
      6'b011110 : begin
        _zz_2807_ = int_reg_array_27_30_imag;
        _zz_2808_ = int_reg_array_27_30_real;
      end
      6'b011111 : begin
        _zz_2807_ = int_reg_array_27_31_imag;
        _zz_2808_ = int_reg_array_27_31_real;
      end
      6'b100000 : begin
        _zz_2807_ = int_reg_array_27_32_imag;
        _zz_2808_ = int_reg_array_27_32_real;
      end
      6'b100001 : begin
        _zz_2807_ = int_reg_array_27_33_imag;
        _zz_2808_ = int_reg_array_27_33_real;
      end
      6'b100010 : begin
        _zz_2807_ = int_reg_array_27_34_imag;
        _zz_2808_ = int_reg_array_27_34_real;
      end
      6'b100011 : begin
        _zz_2807_ = int_reg_array_27_35_imag;
        _zz_2808_ = int_reg_array_27_35_real;
      end
      6'b100100 : begin
        _zz_2807_ = int_reg_array_27_36_imag;
        _zz_2808_ = int_reg_array_27_36_real;
      end
      6'b100101 : begin
        _zz_2807_ = int_reg_array_27_37_imag;
        _zz_2808_ = int_reg_array_27_37_real;
      end
      6'b100110 : begin
        _zz_2807_ = int_reg_array_27_38_imag;
        _zz_2808_ = int_reg_array_27_38_real;
      end
      6'b100111 : begin
        _zz_2807_ = int_reg_array_27_39_imag;
        _zz_2808_ = int_reg_array_27_39_real;
      end
      6'b101000 : begin
        _zz_2807_ = int_reg_array_27_40_imag;
        _zz_2808_ = int_reg_array_27_40_real;
      end
      6'b101001 : begin
        _zz_2807_ = int_reg_array_27_41_imag;
        _zz_2808_ = int_reg_array_27_41_real;
      end
      6'b101010 : begin
        _zz_2807_ = int_reg_array_27_42_imag;
        _zz_2808_ = int_reg_array_27_42_real;
      end
      6'b101011 : begin
        _zz_2807_ = int_reg_array_27_43_imag;
        _zz_2808_ = int_reg_array_27_43_real;
      end
      6'b101100 : begin
        _zz_2807_ = int_reg_array_27_44_imag;
        _zz_2808_ = int_reg_array_27_44_real;
      end
      6'b101101 : begin
        _zz_2807_ = int_reg_array_27_45_imag;
        _zz_2808_ = int_reg_array_27_45_real;
      end
      6'b101110 : begin
        _zz_2807_ = int_reg_array_27_46_imag;
        _zz_2808_ = int_reg_array_27_46_real;
      end
      6'b101111 : begin
        _zz_2807_ = int_reg_array_27_47_imag;
        _zz_2808_ = int_reg_array_27_47_real;
      end
      6'b110000 : begin
        _zz_2807_ = int_reg_array_27_48_imag;
        _zz_2808_ = int_reg_array_27_48_real;
      end
      default : begin
        _zz_2807_ = int_reg_array_27_49_imag;
        _zz_2808_ = int_reg_array_27_49_real;
      end
    endcase
  end

  always @(*) begin
    case(_zz_1542_)
      6'b000000 : begin
        _zz_2809_ = int_reg_array_28_0_imag;
        _zz_2810_ = int_reg_array_28_0_real;
      end
      6'b000001 : begin
        _zz_2809_ = int_reg_array_28_1_imag;
        _zz_2810_ = int_reg_array_28_1_real;
      end
      6'b000010 : begin
        _zz_2809_ = int_reg_array_28_2_imag;
        _zz_2810_ = int_reg_array_28_2_real;
      end
      6'b000011 : begin
        _zz_2809_ = int_reg_array_28_3_imag;
        _zz_2810_ = int_reg_array_28_3_real;
      end
      6'b000100 : begin
        _zz_2809_ = int_reg_array_28_4_imag;
        _zz_2810_ = int_reg_array_28_4_real;
      end
      6'b000101 : begin
        _zz_2809_ = int_reg_array_28_5_imag;
        _zz_2810_ = int_reg_array_28_5_real;
      end
      6'b000110 : begin
        _zz_2809_ = int_reg_array_28_6_imag;
        _zz_2810_ = int_reg_array_28_6_real;
      end
      6'b000111 : begin
        _zz_2809_ = int_reg_array_28_7_imag;
        _zz_2810_ = int_reg_array_28_7_real;
      end
      6'b001000 : begin
        _zz_2809_ = int_reg_array_28_8_imag;
        _zz_2810_ = int_reg_array_28_8_real;
      end
      6'b001001 : begin
        _zz_2809_ = int_reg_array_28_9_imag;
        _zz_2810_ = int_reg_array_28_9_real;
      end
      6'b001010 : begin
        _zz_2809_ = int_reg_array_28_10_imag;
        _zz_2810_ = int_reg_array_28_10_real;
      end
      6'b001011 : begin
        _zz_2809_ = int_reg_array_28_11_imag;
        _zz_2810_ = int_reg_array_28_11_real;
      end
      6'b001100 : begin
        _zz_2809_ = int_reg_array_28_12_imag;
        _zz_2810_ = int_reg_array_28_12_real;
      end
      6'b001101 : begin
        _zz_2809_ = int_reg_array_28_13_imag;
        _zz_2810_ = int_reg_array_28_13_real;
      end
      6'b001110 : begin
        _zz_2809_ = int_reg_array_28_14_imag;
        _zz_2810_ = int_reg_array_28_14_real;
      end
      6'b001111 : begin
        _zz_2809_ = int_reg_array_28_15_imag;
        _zz_2810_ = int_reg_array_28_15_real;
      end
      6'b010000 : begin
        _zz_2809_ = int_reg_array_28_16_imag;
        _zz_2810_ = int_reg_array_28_16_real;
      end
      6'b010001 : begin
        _zz_2809_ = int_reg_array_28_17_imag;
        _zz_2810_ = int_reg_array_28_17_real;
      end
      6'b010010 : begin
        _zz_2809_ = int_reg_array_28_18_imag;
        _zz_2810_ = int_reg_array_28_18_real;
      end
      6'b010011 : begin
        _zz_2809_ = int_reg_array_28_19_imag;
        _zz_2810_ = int_reg_array_28_19_real;
      end
      6'b010100 : begin
        _zz_2809_ = int_reg_array_28_20_imag;
        _zz_2810_ = int_reg_array_28_20_real;
      end
      6'b010101 : begin
        _zz_2809_ = int_reg_array_28_21_imag;
        _zz_2810_ = int_reg_array_28_21_real;
      end
      6'b010110 : begin
        _zz_2809_ = int_reg_array_28_22_imag;
        _zz_2810_ = int_reg_array_28_22_real;
      end
      6'b010111 : begin
        _zz_2809_ = int_reg_array_28_23_imag;
        _zz_2810_ = int_reg_array_28_23_real;
      end
      6'b011000 : begin
        _zz_2809_ = int_reg_array_28_24_imag;
        _zz_2810_ = int_reg_array_28_24_real;
      end
      6'b011001 : begin
        _zz_2809_ = int_reg_array_28_25_imag;
        _zz_2810_ = int_reg_array_28_25_real;
      end
      6'b011010 : begin
        _zz_2809_ = int_reg_array_28_26_imag;
        _zz_2810_ = int_reg_array_28_26_real;
      end
      6'b011011 : begin
        _zz_2809_ = int_reg_array_28_27_imag;
        _zz_2810_ = int_reg_array_28_27_real;
      end
      6'b011100 : begin
        _zz_2809_ = int_reg_array_28_28_imag;
        _zz_2810_ = int_reg_array_28_28_real;
      end
      6'b011101 : begin
        _zz_2809_ = int_reg_array_28_29_imag;
        _zz_2810_ = int_reg_array_28_29_real;
      end
      6'b011110 : begin
        _zz_2809_ = int_reg_array_28_30_imag;
        _zz_2810_ = int_reg_array_28_30_real;
      end
      6'b011111 : begin
        _zz_2809_ = int_reg_array_28_31_imag;
        _zz_2810_ = int_reg_array_28_31_real;
      end
      6'b100000 : begin
        _zz_2809_ = int_reg_array_28_32_imag;
        _zz_2810_ = int_reg_array_28_32_real;
      end
      6'b100001 : begin
        _zz_2809_ = int_reg_array_28_33_imag;
        _zz_2810_ = int_reg_array_28_33_real;
      end
      6'b100010 : begin
        _zz_2809_ = int_reg_array_28_34_imag;
        _zz_2810_ = int_reg_array_28_34_real;
      end
      6'b100011 : begin
        _zz_2809_ = int_reg_array_28_35_imag;
        _zz_2810_ = int_reg_array_28_35_real;
      end
      6'b100100 : begin
        _zz_2809_ = int_reg_array_28_36_imag;
        _zz_2810_ = int_reg_array_28_36_real;
      end
      6'b100101 : begin
        _zz_2809_ = int_reg_array_28_37_imag;
        _zz_2810_ = int_reg_array_28_37_real;
      end
      6'b100110 : begin
        _zz_2809_ = int_reg_array_28_38_imag;
        _zz_2810_ = int_reg_array_28_38_real;
      end
      6'b100111 : begin
        _zz_2809_ = int_reg_array_28_39_imag;
        _zz_2810_ = int_reg_array_28_39_real;
      end
      6'b101000 : begin
        _zz_2809_ = int_reg_array_28_40_imag;
        _zz_2810_ = int_reg_array_28_40_real;
      end
      6'b101001 : begin
        _zz_2809_ = int_reg_array_28_41_imag;
        _zz_2810_ = int_reg_array_28_41_real;
      end
      6'b101010 : begin
        _zz_2809_ = int_reg_array_28_42_imag;
        _zz_2810_ = int_reg_array_28_42_real;
      end
      6'b101011 : begin
        _zz_2809_ = int_reg_array_28_43_imag;
        _zz_2810_ = int_reg_array_28_43_real;
      end
      6'b101100 : begin
        _zz_2809_ = int_reg_array_28_44_imag;
        _zz_2810_ = int_reg_array_28_44_real;
      end
      6'b101101 : begin
        _zz_2809_ = int_reg_array_28_45_imag;
        _zz_2810_ = int_reg_array_28_45_real;
      end
      6'b101110 : begin
        _zz_2809_ = int_reg_array_28_46_imag;
        _zz_2810_ = int_reg_array_28_46_real;
      end
      6'b101111 : begin
        _zz_2809_ = int_reg_array_28_47_imag;
        _zz_2810_ = int_reg_array_28_47_real;
      end
      6'b110000 : begin
        _zz_2809_ = int_reg_array_28_48_imag;
        _zz_2810_ = int_reg_array_28_48_real;
      end
      default : begin
        _zz_2809_ = int_reg_array_28_49_imag;
        _zz_2810_ = int_reg_array_28_49_real;
      end
    endcase
  end

  always @(*) begin
    case(_zz_1597_)
      6'b000000 : begin
        _zz_2811_ = int_reg_array_29_0_imag;
        _zz_2812_ = int_reg_array_29_0_real;
      end
      6'b000001 : begin
        _zz_2811_ = int_reg_array_29_1_imag;
        _zz_2812_ = int_reg_array_29_1_real;
      end
      6'b000010 : begin
        _zz_2811_ = int_reg_array_29_2_imag;
        _zz_2812_ = int_reg_array_29_2_real;
      end
      6'b000011 : begin
        _zz_2811_ = int_reg_array_29_3_imag;
        _zz_2812_ = int_reg_array_29_3_real;
      end
      6'b000100 : begin
        _zz_2811_ = int_reg_array_29_4_imag;
        _zz_2812_ = int_reg_array_29_4_real;
      end
      6'b000101 : begin
        _zz_2811_ = int_reg_array_29_5_imag;
        _zz_2812_ = int_reg_array_29_5_real;
      end
      6'b000110 : begin
        _zz_2811_ = int_reg_array_29_6_imag;
        _zz_2812_ = int_reg_array_29_6_real;
      end
      6'b000111 : begin
        _zz_2811_ = int_reg_array_29_7_imag;
        _zz_2812_ = int_reg_array_29_7_real;
      end
      6'b001000 : begin
        _zz_2811_ = int_reg_array_29_8_imag;
        _zz_2812_ = int_reg_array_29_8_real;
      end
      6'b001001 : begin
        _zz_2811_ = int_reg_array_29_9_imag;
        _zz_2812_ = int_reg_array_29_9_real;
      end
      6'b001010 : begin
        _zz_2811_ = int_reg_array_29_10_imag;
        _zz_2812_ = int_reg_array_29_10_real;
      end
      6'b001011 : begin
        _zz_2811_ = int_reg_array_29_11_imag;
        _zz_2812_ = int_reg_array_29_11_real;
      end
      6'b001100 : begin
        _zz_2811_ = int_reg_array_29_12_imag;
        _zz_2812_ = int_reg_array_29_12_real;
      end
      6'b001101 : begin
        _zz_2811_ = int_reg_array_29_13_imag;
        _zz_2812_ = int_reg_array_29_13_real;
      end
      6'b001110 : begin
        _zz_2811_ = int_reg_array_29_14_imag;
        _zz_2812_ = int_reg_array_29_14_real;
      end
      6'b001111 : begin
        _zz_2811_ = int_reg_array_29_15_imag;
        _zz_2812_ = int_reg_array_29_15_real;
      end
      6'b010000 : begin
        _zz_2811_ = int_reg_array_29_16_imag;
        _zz_2812_ = int_reg_array_29_16_real;
      end
      6'b010001 : begin
        _zz_2811_ = int_reg_array_29_17_imag;
        _zz_2812_ = int_reg_array_29_17_real;
      end
      6'b010010 : begin
        _zz_2811_ = int_reg_array_29_18_imag;
        _zz_2812_ = int_reg_array_29_18_real;
      end
      6'b010011 : begin
        _zz_2811_ = int_reg_array_29_19_imag;
        _zz_2812_ = int_reg_array_29_19_real;
      end
      6'b010100 : begin
        _zz_2811_ = int_reg_array_29_20_imag;
        _zz_2812_ = int_reg_array_29_20_real;
      end
      6'b010101 : begin
        _zz_2811_ = int_reg_array_29_21_imag;
        _zz_2812_ = int_reg_array_29_21_real;
      end
      6'b010110 : begin
        _zz_2811_ = int_reg_array_29_22_imag;
        _zz_2812_ = int_reg_array_29_22_real;
      end
      6'b010111 : begin
        _zz_2811_ = int_reg_array_29_23_imag;
        _zz_2812_ = int_reg_array_29_23_real;
      end
      6'b011000 : begin
        _zz_2811_ = int_reg_array_29_24_imag;
        _zz_2812_ = int_reg_array_29_24_real;
      end
      6'b011001 : begin
        _zz_2811_ = int_reg_array_29_25_imag;
        _zz_2812_ = int_reg_array_29_25_real;
      end
      6'b011010 : begin
        _zz_2811_ = int_reg_array_29_26_imag;
        _zz_2812_ = int_reg_array_29_26_real;
      end
      6'b011011 : begin
        _zz_2811_ = int_reg_array_29_27_imag;
        _zz_2812_ = int_reg_array_29_27_real;
      end
      6'b011100 : begin
        _zz_2811_ = int_reg_array_29_28_imag;
        _zz_2812_ = int_reg_array_29_28_real;
      end
      6'b011101 : begin
        _zz_2811_ = int_reg_array_29_29_imag;
        _zz_2812_ = int_reg_array_29_29_real;
      end
      6'b011110 : begin
        _zz_2811_ = int_reg_array_29_30_imag;
        _zz_2812_ = int_reg_array_29_30_real;
      end
      6'b011111 : begin
        _zz_2811_ = int_reg_array_29_31_imag;
        _zz_2812_ = int_reg_array_29_31_real;
      end
      6'b100000 : begin
        _zz_2811_ = int_reg_array_29_32_imag;
        _zz_2812_ = int_reg_array_29_32_real;
      end
      6'b100001 : begin
        _zz_2811_ = int_reg_array_29_33_imag;
        _zz_2812_ = int_reg_array_29_33_real;
      end
      6'b100010 : begin
        _zz_2811_ = int_reg_array_29_34_imag;
        _zz_2812_ = int_reg_array_29_34_real;
      end
      6'b100011 : begin
        _zz_2811_ = int_reg_array_29_35_imag;
        _zz_2812_ = int_reg_array_29_35_real;
      end
      6'b100100 : begin
        _zz_2811_ = int_reg_array_29_36_imag;
        _zz_2812_ = int_reg_array_29_36_real;
      end
      6'b100101 : begin
        _zz_2811_ = int_reg_array_29_37_imag;
        _zz_2812_ = int_reg_array_29_37_real;
      end
      6'b100110 : begin
        _zz_2811_ = int_reg_array_29_38_imag;
        _zz_2812_ = int_reg_array_29_38_real;
      end
      6'b100111 : begin
        _zz_2811_ = int_reg_array_29_39_imag;
        _zz_2812_ = int_reg_array_29_39_real;
      end
      6'b101000 : begin
        _zz_2811_ = int_reg_array_29_40_imag;
        _zz_2812_ = int_reg_array_29_40_real;
      end
      6'b101001 : begin
        _zz_2811_ = int_reg_array_29_41_imag;
        _zz_2812_ = int_reg_array_29_41_real;
      end
      6'b101010 : begin
        _zz_2811_ = int_reg_array_29_42_imag;
        _zz_2812_ = int_reg_array_29_42_real;
      end
      6'b101011 : begin
        _zz_2811_ = int_reg_array_29_43_imag;
        _zz_2812_ = int_reg_array_29_43_real;
      end
      6'b101100 : begin
        _zz_2811_ = int_reg_array_29_44_imag;
        _zz_2812_ = int_reg_array_29_44_real;
      end
      6'b101101 : begin
        _zz_2811_ = int_reg_array_29_45_imag;
        _zz_2812_ = int_reg_array_29_45_real;
      end
      6'b101110 : begin
        _zz_2811_ = int_reg_array_29_46_imag;
        _zz_2812_ = int_reg_array_29_46_real;
      end
      6'b101111 : begin
        _zz_2811_ = int_reg_array_29_47_imag;
        _zz_2812_ = int_reg_array_29_47_real;
      end
      6'b110000 : begin
        _zz_2811_ = int_reg_array_29_48_imag;
        _zz_2812_ = int_reg_array_29_48_real;
      end
      default : begin
        _zz_2811_ = int_reg_array_29_49_imag;
        _zz_2812_ = int_reg_array_29_49_real;
      end
    endcase
  end

  always @(*) begin
    case(_zz_1652_)
      6'b000000 : begin
        _zz_2813_ = int_reg_array_30_0_imag;
        _zz_2814_ = int_reg_array_30_0_real;
      end
      6'b000001 : begin
        _zz_2813_ = int_reg_array_30_1_imag;
        _zz_2814_ = int_reg_array_30_1_real;
      end
      6'b000010 : begin
        _zz_2813_ = int_reg_array_30_2_imag;
        _zz_2814_ = int_reg_array_30_2_real;
      end
      6'b000011 : begin
        _zz_2813_ = int_reg_array_30_3_imag;
        _zz_2814_ = int_reg_array_30_3_real;
      end
      6'b000100 : begin
        _zz_2813_ = int_reg_array_30_4_imag;
        _zz_2814_ = int_reg_array_30_4_real;
      end
      6'b000101 : begin
        _zz_2813_ = int_reg_array_30_5_imag;
        _zz_2814_ = int_reg_array_30_5_real;
      end
      6'b000110 : begin
        _zz_2813_ = int_reg_array_30_6_imag;
        _zz_2814_ = int_reg_array_30_6_real;
      end
      6'b000111 : begin
        _zz_2813_ = int_reg_array_30_7_imag;
        _zz_2814_ = int_reg_array_30_7_real;
      end
      6'b001000 : begin
        _zz_2813_ = int_reg_array_30_8_imag;
        _zz_2814_ = int_reg_array_30_8_real;
      end
      6'b001001 : begin
        _zz_2813_ = int_reg_array_30_9_imag;
        _zz_2814_ = int_reg_array_30_9_real;
      end
      6'b001010 : begin
        _zz_2813_ = int_reg_array_30_10_imag;
        _zz_2814_ = int_reg_array_30_10_real;
      end
      6'b001011 : begin
        _zz_2813_ = int_reg_array_30_11_imag;
        _zz_2814_ = int_reg_array_30_11_real;
      end
      6'b001100 : begin
        _zz_2813_ = int_reg_array_30_12_imag;
        _zz_2814_ = int_reg_array_30_12_real;
      end
      6'b001101 : begin
        _zz_2813_ = int_reg_array_30_13_imag;
        _zz_2814_ = int_reg_array_30_13_real;
      end
      6'b001110 : begin
        _zz_2813_ = int_reg_array_30_14_imag;
        _zz_2814_ = int_reg_array_30_14_real;
      end
      6'b001111 : begin
        _zz_2813_ = int_reg_array_30_15_imag;
        _zz_2814_ = int_reg_array_30_15_real;
      end
      6'b010000 : begin
        _zz_2813_ = int_reg_array_30_16_imag;
        _zz_2814_ = int_reg_array_30_16_real;
      end
      6'b010001 : begin
        _zz_2813_ = int_reg_array_30_17_imag;
        _zz_2814_ = int_reg_array_30_17_real;
      end
      6'b010010 : begin
        _zz_2813_ = int_reg_array_30_18_imag;
        _zz_2814_ = int_reg_array_30_18_real;
      end
      6'b010011 : begin
        _zz_2813_ = int_reg_array_30_19_imag;
        _zz_2814_ = int_reg_array_30_19_real;
      end
      6'b010100 : begin
        _zz_2813_ = int_reg_array_30_20_imag;
        _zz_2814_ = int_reg_array_30_20_real;
      end
      6'b010101 : begin
        _zz_2813_ = int_reg_array_30_21_imag;
        _zz_2814_ = int_reg_array_30_21_real;
      end
      6'b010110 : begin
        _zz_2813_ = int_reg_array_30_22_imag;
        _zz_2814_ = int_reg_array_30_22_real;
      end
      6'b010111 : begin
        _zz_2813_ = int_reg_array_30_23_imag;
        _zz_2814_ = int_reg_array_30_23_real;
      end
      6'b011000 : begin
        _zz_2813_ = int_reg_array_30_24_imag;
        _zz_2814_ = int_reg_array_30_24_real;
      end
      6'b011001 : begin
        _zz_2813_ = int_reg_array_30_25_imag;
        _zz_2814_ = int_reg_array_30_25_real;
      end
      6'b011010 : begin
        _zz_2813_ = int_reg_array_30_26_imag;
        _zz_2814_ = int_reg_array_30_26_real;
      end
      6'b011011 : begin
        _zz_2813_ = int_reg_array_30_27_imag;
        _zz_2814_ = int_reg_array_30_27_real;
      end
      6'b011100 : begin
        _zz_2813_ = int_reg_array_30_28_imag;
        _zz_2814_ = int_reg_array_30_28_real;
      end
      6'b011101 : begin
        _zz_2813_ = int_reg_array_30_29_imag;
        _zz_2814_ = int_reg_array_30_29_real;
      end
      6'b011110 : begin
        _zz_2813_ = int_reg_array_30_30_imag;
        _zz_2814_ = int_reg_array_30_30_real;
      end
      6'b011111 : begin
        _zz_2813_ = int_reg_array_30_31_imag;
        _zz_2814_ = int_reg_array_30_31_real;
      end
      6'b100000 : begin
        _zz_2813_ = int_reg_array_30_32_imag;
        _zz_2814_ = int_reg_array_30_32_real;
      end
      6'b100001 : begin
        _zz_2813_ = int_reg_array_30_33_imag;
        _zz_2814_ = int_reg_array_30_33_real;
      end
      6'b100010 : begin
        _zz_2813_ = int_reg_array_30_34_imag;
        _zz_2814_ = int_reg_array_30_34_real;
      end
      6'b100011 : begin
        _zz_2813_ = int_reg_array_30_35_imag;
        _zz_2814_ = int_reg_array_30_35_real;
      end
      6'b100100 : begin
        _zz_2813_ = int_reg_array_30_36_imag;
        _zz_2814_ = int_reg_array_30_36_real;
      end
      6'b100101 : begin
        _zz_2813_ = int_reg_array_30_37_imag;
        _zz_2814_ = int_reg_array_30_37_real;
      end
      6'b100110 : begin
        _zz_2813_ = int_reg_array_30_38_imag;
        _zz_2814_ = int_reg_array_30_38_real;
      end
      6'b100111 : begin
        _zz_2813_ = int_reg_array_30_39_imag;
        _zz_2814_ = int_reg_array_30_39_real;
      end
      6'b101000 : begin
        _zz_2813_ = int_reg_array_30_40_imag;
        _zz_2814_ = int_reg_array_30_40_real;
      end
      6'b101001 : begin
        _zz_2813_ = int_reg_array_30_41_imag;
        _zz_2814_ = int_reg_array_30_41_real;
      end
      6'b101010 : begin
        _zz_2813_ = int_reg_array_30_42_imag;
        _zz_2814_ = int_reg_array_30_42_real;
      end
      6'b101011 : begin
        _zz_2813_ = int_reg_array_30_43_imag;
        _zz_2814_ = int_reg_array_30_43_real;
      end
      6'b101100 : begin
        _zz_2813_ = int_reg_array_30_44_imag;
        _zz_2814_ = int_reg_array_30_44_real;
      end
      6'b101101 : begin
        _zz_2813_ = int_reg_array_30_45_imag;
        _zz_2814_ = int_reg_array_30_45_real;
      end
      6'b101110 : begin
        _zz_2813_ = int_reg_array_30_46_imag;
        _zz_2814_ = int_reg_array_30_46_real;
      end
      6'b101111 : begin
        _zz_2813_ = int_reg_array_30_47_imag;
        _zz_2814_ = int_reg_array_30_47_real;
      end
      6'b110000 : begin
        _zz_2813_ = int_reg_array_30_48_imag;
        _zz_2814_ = int_reg_array_30_48_real;
      end
      default : begin
        _zz_2813_ = int_reg_array_30_49_imag;
        _zz_2814_ = int_reg_array_30_49_real;
      end
    endcase
  end

  always @(*) begin
    case(_zz_1707_)
      6'b000000 : begin
        _zz_2815_ = int_reg_array_31_0_imag;
        _zz_2816_ = int_reg_array_31_0_real;
      end
      6'b000001 : begin
        _zz_2815_ = int_reg_array_31_1_imag;
        _zz_2816_ = int_reg_array_31_1_real;
      end
      6'b000010 : begin
        _zz_2815_ = int_reg_array_31_2_imag;
        _zz_2816_ = int_reg_array_31_2_real;
      end
      6'b000011 : begin
        _zz_2815_ = int_reg_array_31_3_imag;
        _zz_2816_ = int_reg_array_31_3_real;
      end
      6'b000100 : begin
        _zz_2815_ = int_reg_array_31_4_imag;
        _zz_2816_ = int_reg_array_31_4_real;
      end
      6'b000101 : begin
        _zz_2815_ = int_reg_array_31_5_imag;
        _zz_2816_ = int_reg_array_31_5_real;
      end
      6'b000110 : begin
        _zz_2815_ = int_reg_array_31_6_imag;
        _zz_2816_ = int_reg_array_31_6_real;
      end
      6'b000111 : begin
        _zz_2815_ = int_reg_array_31_7_imag;
        _zz_2816_ = int_reg_array_31_7_real;
      end
      6'b001000 : begin
        _zz_2815_ = int_reg_array_31_8_imag;
        _zz_2816_ = int_reg_array_31_8_real;
      end
      6'b001001 : begin
        _zz_2815_ = int_reg_array_31_9_imag;
        _zz_2816_ = int_reg_array_31_9_real;
      end
      6'b001010 : begin
        _zz_2815_ = int_reg_array_31_10_imag;
        _zz_2816_ = int_reg_array_31_10_real;
      end
      6'b001011 : begin
        _zz_2815_ = int_reg_array_31_11_imag;
        _zz_2816_ = int_reg_array_31_11_real;
      end
      6'b001100 : begin
        _zz_2815_ = int_reg_array_31_12_imag;
        _zz_2816_ = int_reg_array_31_12_real;
      end
      6'b001101 : begin
        _zz_2815_ = int_reg_array_31_13_imag;
        _zz_2816_ = int_reg_array_31_13_real;
      end
      6'b001110 : begin
        _zz_2815_ = int_reg_array_31_14_imag;
        _zz_2816_ = int_reg_array_31_14_real;
      end
      6'b001111 : begin
        _zz_2815_ = int_reg_array_31_15_imag;
        _zz_2816_ = int_reg_array_31_15_real;
      end
      6'b010000 : begin
        _zz_2815_ = int_reg_array_31_16_imag;
        _zz_2816_ = int_reg_array_31_16_real;
      end
      6'b010001 : begin
        _zz_2815_ = int_reg_array_31_17_imag;
        _zz_2816_ = int_reg_array_31_17_real;
      end
      6'b010010 : begin
        _zz_2815_ = int_reg_array_31_18_imag;
        _zz_2816_ = int_reg_array_31_18_real;
      end
      6'b010011 : begin
        _zz_2815_ = int_reg_array_31_19_imag;
        _zz_2816_ = int_reg_array_31_19_real;
      end
      6'b010100 : begin
        _zz_2815_ = int_reg_array_31_20_imag;
        _zz_2816_ = int_reg_array_31_20_real;
      end
      6'b010101 : begin
        _zz_2815_ = int_reg_array_31_21_imag;
        _zz_2816_ = int_reg_array_31_21_real;
      end
      6'b010110 : begin
        _zz_2815_ = int_reg_array_31_22_imag;
        _zz_2816_ = int_reg_array_31_22_real;
      end
      6'b010111 : begin
        _zz_2815_ = int_reg_array_31_23_imag;
        _zz_2816_ = int_reg_array_31_23_real;
      end
      6'b011000 : begin
        _zz_2815_ = int_reg_array_31_24_imag;
        _zz_2816_ = int_reg_array_31_24_real;
      end
      6'b011001 : begin
        _zz_2815_ = int_reg_array_31_25_imag;
        _zz_2816_ = int_reg_array_31_25_real;
      end
      6'b011010 : begin
        _zz_2815_ = int_reg_array_31_26_imag;
        _zz_2816_ = int_reg_array_31_26_real;
      end
      6'b011011 : begin
        _zz_2815_ = int_reg_array_31_27_imag;
        _zz_2816_ = int_reg_array_31_27_real;
      end
      6'b011100 : begin
        _zz_2815_ = int_reg_array_31_28_imag;
        _zz_2816_ = int_reg_array_31_28_real;
      end
      6'b011101 : begin
        _zz_2815_ = int_reg_array_31_29_imag;
        _zz_2816_ = int_reg_array_31_29_real;
      end
      6'b011110 : begin
        _zz_2815_ = int_reg_array_31_30_imag;
        _zz_2816_ = int_reg_array_31_30_real;
      end
      6'b011111 : begin
        _zz_2815_ = int_reg_array_31_31_imag;
        _zz_2816_ = int_reg_array_31_31_real;
      end
      6'b100000 : begin
        _zz_2815_ = int_reg_array_31_32_imag;
        _zz_2816_ = int_reg_array_31_32_real;
      end
      6'b100001 : begin
        _zz_2815_ = int_reg_array_31_33_imag;
        _zz_2816_ = int_reg_array_31_33_real;
      end
      6'b100010 : begin
        _zz_2815_ = int_reg_array_31_34_imag;
        _zz_2816_ = int_reg_array_31_34_real;
      end
      6'b100011 : begin
        _zz_2815_ = int_reg_array_31_35_imag;
        _zz_2816_ = int_reg_array_31_35_real;
      end
      6'b100100 : begin
        _zz_2815_ = int_reg_array_31_36_imag;
        _zz_2816_ = int_reg_array_31_36_real;
      end
      6'b100101 : begin
        _zz_2815_ = int_reg_array_31_37_imag;
        _zz_2816_ = int_reg_array_31_37_real;
      end
      6'b100110 : begin
        _zz_2815_ = int_reg_array_31_38_imag;
        _zz_2816_ = int_reg_array_31_38_real;
      end
      6'b100111 : begin
        _zz_2815_ = int_reg_array_31_39_imag;
        _zz_2816_ = int_reg_array_31_39_real;
      end
      6'b101000 : begin
        _zz_2815_ = int_reg_array_31_40_imag;
        _zz_2816_ = int_reg_array_31_40_real;
      end
      6'b101001 : begin
        _zz_2815_ = int_reg_array_31_41_imag;
        _zz_2816_ = int_reg_array_31_41_real;
      end
      6'b101010 : begin
        _zz_2815_ = int_reg_array_31_42_imag;
        _zz_2816_ = int_reg_array_31_42_real;
      end
      6'b101011 : begin
        _zz_2815_ = int_reg_array_31_43_imag;
        _zz_2816_ = int_reg_array_31_43_real;
      end
      6'b101100 : begin
        _zz_2815_ = int_reg_array_31_44_imag;
        _zz_2816_ = int_reg_array_31_44_real;
      end
      6'b101101 : begin
        _zz_2815_ = int_reg_array_31_45_imag;
        _zz_2816_ = int_reg_array_31_45_real;
      end
      6'b101110 : begin
        _zz_2815_ = int_reg_array_31_46_imag;
        _zz_2816_ = int_reg_array_31_46_real;
      end
      6'b101111 : begin
        _zz_2815_ = int_reg_array_31_47_imag;
        _zz_2816_ = int_reg_array_31_47_real;
      end
      6'b110000 : begin
        _zz_2815_ = int_reg_array_31_48_imag;
        _zz_2816_ = int_reg_array_31_48_real;
      end
      default : begin
        _zz_2815_ = int_reg_array_31_49_imag;
        _zz_2816_ = int_reg_array_31_49_real;
      end
    endcase
  end

  always @(*) begin
    case(_zz_1762_)
      6'b000000 : begin
        _zz_2817_ = int_reg_array_32_0_imag;
        _zz_2818_ = int_reg_array_32_0_real;
      end
      6'b000001 : begin
        _zz_2817_ = int_reg_array_32_1_imag;
        _zz_2818_ = int_reg_array_32_1_real;
      end
      6'b000010 : begin
        _zz_2817_ = int_reg_array_32_2_imag;
        _zz_2818_ = int_reg_array_32_2_real;
      end
      6'b000011 : begin
        _zz_2817_ = int_reg_array_32_3_imag;
        _zz_2818_ = int_reg_array_32_3_real;
      end
      6'b000100 : begin
        _zz_2817_ = int_reg_array_32_4_imag;
        _zz_2818_ = int_reg_array_32_4_real;
      end
      6'b000101 : begin
        _zz_2817_ = int_reg_array_32_5_imag;
        _zz_2818_ = int_reg_array_32_5_real;
      end
      6'b000110 : begin
        _zz_2817_ = int_reg_array_32_6_imag;
        _zz_2818_ = int_reg_array_32_6_real;
      end
      6'b000111 : begin
        _zz_2817_ = int_reg_array_32_7_imag;
        _zz_2818_ = int_reg_array_32_7_real;
      end
      6'b001000 : begin
        _zz_2817_ = int_reg_array_32_8_imag;
        _zz_2818_ = int_reg_array_32_8_real;
      end
      6'b001001 : begin
        _zz_2817_ = int_reg_array_32_9_imag;
        _zz_2818_ = int_reg_array_32_9_real;
      end
      6'b001010 : begin
        _zz_2817_ = int_reg_array_32_10_imag;
        _zz_2818_ = int_reg_array_32_10_real;
      end
      6'b001011 : begin
        _zz_2817_ = int_reg_array_32_11_imag;
        _zz_2818_ = int_reg_array_32_11_real;
      end
      6'b001100 : begin
        _zz_2817_ = int_reg_array_32_12_imag;
        _zz_2818_ = int_reg_array_32_12_real;
      end
      6'b001101 : begin
        _zz_2817_ = int_reg_array_32_13_imag;
        _zz_2818_ = int_reg_array_32_13_real;
      end
      6'b001110 : begin
        _zz_2817_ = int_reg_array_32_14_imag;
        _zz_2818_ = int_reg_array_32_14_real;
      end
      6'b001111 : begin
        _zz_2817_ = int_reg_array_32_15_imag;
        _zz_2818_ = int_reg_array_32_15_real;
      end
      6'b010000 : begin
        _zz_2817_ = int_reg_array_32_16_imag;
        _zz_2818_ = int_reg_array_32_16_real;
      end
      6'b010001 : begin
        _zz_2817_ = int_reg_array_32_17_imag;
        _zz_2818_ = int_reg_array_32_17_real;
      end
      6'b010010 : begin
        _zz_2817_ = int_reg_array_32_18_imag;
        _zz_2818_ = int_reg_array_32_18_real;
      end
      6'b010011 : begin
        _zz_2817_ = int_reg_array_32_19_imag;
        _zz_2818_ = int_reg_array_32_19_real;
      end
      6'b010100 : begin
        _zz_2817_ = int_reg_array_32_20_imag;
        _zz_2818_ = int_reg_array_32_20_real;
      end
      6'b010101 : begin
        _zz_2817_ = int_reg_array_32_21_imag;
        _zz_2818_ = int_reg_array_32_21_real;
      end
      6'b010110 : begin
        _zz_2817_ = int_reg_array_32_22_imag;
        _zz_2818_ = int_reg_array_32_22_real;
      end
      6'b010111 : begin
        _zz_2817_ = int_reg_array_32_23_imag;
        _zz_2818_ = int_reg_array_32_23_real;
      end
      6'b011000 : begin
        _zz_2817_ = int_reg_array_32_24_imag;
        _zz_2818_ = int_reg_array_32_24_real;
      end
      6'b011001 : begin
        _zz_2817_ = int_reg_array_32_25_imag;
        _zz_2818_ = int_reg_array_32_25_real;
      end
      6'b011010 : begin
        _zz_2817_ = int_reg_array_32_26_imag;
        _zz_2818_ = int_reg_array_32_26_real;
      end
      6'b011011 : begin
        _zz_2817_ = int_reg_array_32_27_imag;
        _zz_2818_ = int_reg_array_32_27_real;
      end
      6'b011100 : begin
        _zz_2817_ = int_reg_array_32_28_imag;
        _zz_2818_ = int_reg_array_32_28_real;
      end
      6'b011101 : begin
        _zz_2817_ = int_reg_array_32_29_imag;
        _zz_2818_ = int_reg_array_32_29_real;
      end
      6'b011110 : begin
        _zz_2817_ = int_reg_array_32_30_imag;
        _zz_2818_ = int_reg_array_32_30_real;
      end
      6'b011111 : begin
        _zz_2817_ = int_reg_array_32_31_imag;
        _zz_2818_ = int_reg_array_32_31_real;
      end
      6'b100000 : begin
        _zz_2817_ = int_reg_array_32_32_imag;
        _zz_2818_ = int_reg_array_32_32_real;
      end
      6'b100001 : begin
        _zz_2817_ = int_reg_array_32_33_imag;
        _zz_2818_ = int_reg_array_32_33_real;
      end
      6'b100010 : begin
        _zz_2817_ = int_reg_array_32_34_imag;
        _zz_2818_ = int_reg_array_32_34_real;
      end
      6'b100011 : begin
        _zz_2817_ = int_reg_array_32_35_imag;
        _zz_2818_ = int_reg_array_32_35_real;
      end
      6'b100100 : begin
        _zz_2817_ = int_reg_array_32_36_imag;
        _zz_2818_ = int_reg_array_32_36_real;
      end
      6'b100101 : begin
        _zz_2817_ = int_reg_array_32_37_imag;
        _zz_2818_ = int_reg_array_32_37_real;
      end
      6'b100110 : begin
        _zz_2817_ = int_reg_array_32_38_imag;
        _zz_2818_ = int_reg_array_32_38_real;
      end
      6'b100111 : begin
        _zz_2817_ = int_reg_array_32_39_imag;
        _zz_2818_ = int_reg_array_32_39_real;
      end
      6'b101000 : begin
        _zz_2817_ = int_reg_array_32_40_imag;
        _zz_2818_ = int_reg_array_32_40_real;
      end
      6'b101001 : begin
        _zz_2817_ = int_reg_array_32_41_imag;
        _zz_2818_ = int_reg_array_32_41_real;
      end
      6'b101010 : begin
        _zz_2817_ = int_reg_array_32_42_imag;
        _zz_2818_ = int_reg_array_32_42_real;
      end
      6'b101011 : begin
        _zz_2817_ = int_reg_array_32_43_imag;
        _zz_2818_ = int_reg_array_32_43_real;
      end
      6'b101100 : begin
        _zz_2817_ = int_reg_array_32_44_imag;
        _zz_2818_ = int_reg_array_32_44_real;
      end
      6'b101101 : begin
        _zz_2817_ = int_reg_array_32_45_imag;
        _zz_2818_ = int_reg_array_32_45_real;
      end
      6'b101110 : begin
        _zz_2817_ = int_reg_array_32_46_imag;
        _zz_2818_ = int_reg_array_32_46_real;
      end
      6'b101111 : begin
        _zz_2817_ = int_reg_array_32_47_imag;
        _zz_2818_ = int_reg_array_32_47_real;
      end
      6'b110000 : begin
        _zz_2817_ = int_reg_array_32_48_imag;
        _zz_2818_ = int_reg_array_32_48_real;
      end
      default : begin
        _zz_2817_ = int_reg_array_32_49_imag;
        _zz_2818_ = int_reg_array_32_49_real;
      end
    endcase
  end

  always @(*) begin
    case(_zz_1817_)
      6'b000000 : begin
        _zz_2819_ = int_reg_array_33_0_imag;
        _zz_2820_ = int_reg_array_33_0_real;
      end
      6'b000001 : begin
        _zz_2819_ = int_reg_array_33_1_imag;
        _zz_2820_ = int_reg_array_33_1_real;
      end
      6'b000010 : begin
        _zz_2819_ = int_reg_array_33_2_imag;
        _zz_2820_ = int_reg_array_33_2_real;
      end
      6'b000011 : begin
        _zz_2819_ = int_reg_array_33_3_imag;
        _zz_2820_ = int_reg_array_33_3_real;
      end
      6'b000100 : begin
        _zz_2819_ = int_reg_array_33_4_imag;
        _zz_2820_ = int_reg_array_33_4_real;
      end
      6'b000101 : begin
        _zz_2819_ = int_reg_array_33_5_imag;
        _zz_2820_ = int_reg_array_33_5_real;
      end
      6'b000110 : begin
        _zz_2819_ = int_reg_array_33_6_imag;
        _zz_2820_ = int_reg_array_33_6_real;
      end
      6'b000111 : begin
        _zz_2819_ = int_reg_array_33_7_imag;
        _zz_2820_ = int_reg_array_33_7_real;
      end
      6'b001000 : begin
        _zz_2819_ = int_reg_array_33_8_imag;
        _zz_2820_ = int_reg_array_33_8_real;
      end
      6'b001001 : begin
        _zz_2819_ = int_reg_array_33_9_imag;
        _zz_2820_ = int_reg_array_33_9_real;
      end
      6'b001010 : begin
        _zz_2819_ = int_reg_array_33_10_imag;
        _zz_2820_ = int_reg_array_33_10_real;
      end
      6'b001011 : begin
        _zz_2819_ = int_reg_array_33_11_imag;
        _zz_2820_ = int_reg_array_33_11_real;
      end
      6'b001100 : begin
        _zz_2819_ = int_reg_array_33_12_imag;
        _zz_2820_ = int_reg_array_33_12_real;
      end
      6'b001101 : begin
        _zz_2819_ = int_reg_array_33_13_imag;
        _zz_2820_ = int_reg_array_33_13_real;
      end
      6'b001110 : begin
        _zz_2819_ = int_reg_array_33_14_imag;
        _zz_2820_ = int_reg_array_33_14_real;
      end
      6'b001111 : begin
        _zz_2819_ = int_reg_array_33_15_imag;
        _zz_2820_ = int_reg_array_33_15_real;
      end
      6'b010000 : begin
        _zz_2819_ = int_reg_array_33_16_imag;
        _zz_2820_ = int_reg_array_33_16_real;
      end
      6'b010001 : begin
        _zz_2819_ = int_reg_array_33_17_imag;
        _zz_2820_ = int_reg_array_33_17_real;
      end
      6'b010010 : begin
        _zz_2819_ = int_reg_array_33_18_imag;
        _zz_2820_ = int_reg_array_33_18_real;
      end
      6'b010011 : begin
        _zz_2819_ = int_reg_array_33_19_imag;
        _zz_2820_ = int_reg_array_33_19_real;
      end
      6'b010100 : begin
        _zz_2819_ = int_reg_array_33_20_imag;
        _zz_2820_ = int_reg_array_33_20_real;
      end
      6'b010101 : begin
        _zz_2819_ = int_reg_array_33_21_imag;
        _zz_2820_ = int_reg_array_33_21_real;
      end
      6'b010110 : begin
        _zz_2819_ = int_reg_array_33_22_imag;
        _zz_2820_ = int_reg_array_33_22_real;
      end
      6'b010111 : begin
        _zz_2819_ = int_reg_array_33_23_imag;
        _zz_2820_ = int_reg_array_33_23_real;
      end
      6'b011000 : begin
        _zz_2819_ = int_reg_array_33_24_imag;
        _zz_2820_ = int_reg_array_33_24_real;
      end
      6'b011001 : begin
        _zz_2819_ = int_reg_array_33_25_imag;
        _zz_2820_ = int_reg_array_33_25_real;
      end
      6'b011010 : begin
        _zz_2819_ = int_reg_array_33_26_imag;
        _zz_2820_ = int_reg_array_33_26_real;
      end
      6'b011011 : begin
        _zz_2819_ = int_reg_array_33_27_imag;
        _zz_2820_ = int_reg_array_33_27_real;
      end
      6'b011100 : begin
        _zz_2819_ = int_reg_array_33_28_imag;
        _zz_2820_ = int_reg_array_33_28_real;
      end
      6'b011101 : begin
        _zz_2819_ = int_reg_array_33_29_imag;
        _zz_2820_ = int_reg_array_33_29_real;
      end
      6'b011110 : begin
        _zz_2819_ = int_reg_array_33_30_imag;
        _zz_2820_ = int_reg_array_33_30_real;
      end
      6'b011111 : begin
        _zz_2819_ = int_reg_array_33_31_imag;
        _zz_2820_ = int_reg_array_33_31_real;
      end
      6'b100000 : begin
        _zz_2819_ = int_reg_array_33_32_imag;
        _zz_2820_ = int_reg_array_33_32_real;
      end
      6'b100001 : begin
        _zz_2819_ = int_reg_array_33_33_imag;
        _zz_2820_ = int_reg_array_33_33_real;
      end
      6'b100010 : begin
        _zz_2819_ = int_reg_array_33_34_imag;
        _zz_2820_ = int_reg_array_33_34_real;
      end
      6'b100011 : begin
        _zz_2819_ = int_reg_array_33_35_imag;
        _zz_2820_ = int_reg_array_33_35_real;
      end
      6'b100100 : begin
        _zz_2819_ = int_reg_array_33_36_imag;
        _zz_2820_ = int_reg_array_33_36_real;
      end
      6'b100101 : begin
        _zz_2819_ = int_reg_array_33_37_imag;
        _zz_2820_ = int_reg_array_33_37_real;
      end
      6'b100110 : begin
        _zz_2819_ = int_reg_array_33_38_imag;
        _zz_2820_ = int_reg_array_33_38_real;
      end
      6'b100111 : begin
        _zz_2819_ = int_reg_array_33_39_imag;
        _zz_2820_ = int_reg_array_33_39_real;
      end
      6'b101000 : begin
        _zz_2819_ = int_reg_array_33_40_imag;
        _zz_2820_ = int_reg_array_33_40_real;
      end
      6'b101001 : begin
        _zz_2819_ = int_reg_array_33_41_imag;
        _zz_2820_ = int_reg_array_33_41_real;
      end
      6'b101010 : begin
        _zz_2819_ = int_reg_array_33_42_imag;
        _zz_2820_ = int_reg_array_33_42_real;
      end
      6'b101011 : begin
        _zz_2819_ = int_reg_array_33_43_imag;
        _zz_2820_ = int_reg_array_33_43_real;
      end
      6'b101100 : begin
        _zz_2819_ = int_reg_array_33_44_imag;
        _zz_2820_ = int_reg_array_33_44_real;
      end
      6'b101101 : begin
        _zz_2819_ = int_reg_array_33_45_imag;
        _zz_2820_ = int_reg_array_33_45_real;
      end
      6'b101110 : begin
        _zz_2819_ = int_reg_array_33_46_imag;
        _zz_2820_ = int_reg_array_33_46_real;
      end
      6'b101111 : begin
        _zz_2819_ = int_reg_array_33_47_imag;
        _zz_2820_ = int_reg_array_33_47_real;
      end
      6'b110000 : begin
        _zz_2819_ = int_reg_array_33_48_imag;
        _zz_2820_ = int_reg_array_33_48_real;
      end
      default : begin
        _zz_2819_ = int_reg_array_33_49_imag;
        _zz_2820_ = int_reg_array_33_49_real;
      end
    endcase
  end

  always @(*) begin
    case(_zz_1872_)
      6'b000000 : begin
        _zz_2821_ = int_reg_array_34_0_imag;
        _zz_2822_ = int_reg_array_34_0_real;
      end
      6'b000001 : begin
        _zz_2821_ = int_reg_array_34_1_imag;
        _zz_2822_ = int_reg_array_34_1_real;
      end
      6'b000010 : begin
        _zz_2821_ = int_reg_array_34_2_imag;
        _zz_2822_ = int_reg_array_34_2_real;
      end
      6'b000011 : begin
        _zz_2821_ = int_reg_array_34_3_imag;
        _zz_2822_ = int_reg_array_34_3_real;
      end
      6'b000100 : begin
        _zz_2821_ = int_reg_array_34_4_imag;
        _zz_2822_ = int_reg_array_34_4_real;
      end
      6'b000101 : begin
        _zz_2821_ = int_reg_array_34_5_imag;
        _zz_2822_ = int_reg_array_34_5_real;
      end
      6'b000110 : begin
        _zz_2821_ = int_reg_array_34_6_imag;
        _zz_2822_ = int_reg_array_34_6_real;
      end
      6'b000111 : begin
        _zz_2821_ = int_reg_array_34_7_imag;
        _zz_2822_ = int_reg_array_34_7_real;
      end
      6'b001000 : begin
        _zz_2821_ = int_reg_array_34_8_imag;
        _zz_2822_ = int_reg_array_34_8_real;
      end
      6'b001001 : begin
        _zz_2821_ = int_reg_array_34_9_imag;
        _zz_2822_ = int_reg_array_34_9_real;
      end
      6'b001010 : begin
        _zz_2821_ = int_reg_array_34_10_imag;
        _zz_2822_ = int_reg_array_34_10_real;
      end
      6'b001011 : begin
        _zz_2821_ = int_reg_array_34_11_imag;
        _zz_2822_ = int_reg_array_34_11_real;
      end
      6'b001100 : begin
        _zz_2821_ = int_reg_array_34_12_imag;
        _zz_2822_ = int_reg_array_34_12_real;
      end
      6'b001101 : begin
        _zz_2821_ = int_reg_array_34_13_imag;
        _zz_2822_ = int_reg_array_34_13_real;
      end
      6'b001110 : begin
        _zz_2821_ = int_reg_array_34_14_imag;
        _zz_2822_ = int_reg_array_34_14_real;
      end
      6'b001111 : begin
        _zz_2821_ = int_reg_array_34_15_imag;
        _zz_2822_ = int_reg_array_34_15_real;
      end
      6'b010000 : begin
        _zz_2821_ = int_reg_array_34_16_imag;
        _zz_2822_ = int_reg_array_34_16_real;
      end
      6'b010001 : begin
        _zz_2821_ = int_reg_array_34_17_imag;
        _zz_2822_ = int_reg_array_34_17_real;
      end
      6'b010010 : begin
        _zz_2821_ = int_reg_array_34_18_imag;
        _zz_2822_ = int_reg_array_34_18_real;
      end
      6'b010011 : begin
        _zz_2821_ = int_reg_array_34_19_imag;
        _zz_2822_ = int_reg_array_34_19_real;
      end
      6'b010100 : begin
        _zz_2821_ = int_reg_array_34_20_imag;
        _zz_2822_ = int_reg_array_34_20_real;
      end
      6'b010101 : begin
        _zz_2821_ = int_reg_array_34_21_imag;
        _zz_2822_ = int_reg_array_34_21_real;
      end
      6'b010110 : begin
        _zz_2821_ = int_reg_array_34_22_imag;
        _zz_2822_ = int_reg_array_34_22_real;
      end
      6'b010111 : begin
        _zz_2821_ = int_reg_array_34_23_imag;
        _zz_2822_ = int_reg_array_34_23_real;
      end
      6'b011000 : begin
        _zz_2821_ = int_reg_array_34_24_imag;
        _zz_2822_ = int_reg_array_34_24_real;
      end
      6'b011001 : begin
        _zz_2821_ = int_reg_array_34_25_imag;
        _zz_2822_ = int_reg_array_34_25_real;
      end
      6'b011010 : begin
        _zz_2821_ = int_reg_array_34_26_imag;
        _zz_2822_ = int_reg_array_34_26_real;
      end
      6'b011011 : begin
        _zz_2821_ = int_reg_array_34_27_imag;
        _zz_2822_ = int_reg_array_34_27_real;
      end
      6'b011100 : begin
        _zz_2821_ = int_reg_array_34_28_imag;
        _zz_2822_ = int_reg_array_34_28_real;
      end
      6'b011101 : begin
        _zz_2821_ = int_reg_array_34_29_imag;
        _zz_2822_ = int_reg_array_34_29_real;
      end
      6'b011110 : begin
        _zz_2821_ = int_reg_array_34_30_imag;
        _zz_2822_ = int_reg_array_34_30_real;
      end
      6'b011111 : begin
        _zz_2821_ = int_reg_array_34_31_imag;
        _zz_2822_ = int_reg_array_34_31_real;
      end
      6'b100000 : begin
        _zz_2821_ = int_reg_array_34_32_imag;
        _zz_2822_ = int_reg_array_34_32_real;
      end
      6'b100001 : begin
        _zz_2821_ = int_reg_array_34_33_imag;
        _zz_2822_ = int_reg_array_34_33_real;
      end
      6'b100010 : begin
        _zz_2821_ = int_reg_array_34_34_imag;
        _zz_2822_ = int_reg_array_34_34_real;
      end
      6'b100011 : begin
        _zz_2821_ = int_reg_array_34_35_imag;
        _zz_2822_ = int_reg_array_34_35_real;
      end
      6'b100100 : begin
        _zz_2821_ = int_reg_array_34_36_imag;
        _zz_2822_ = int_reg_array_34_36_real;
      end
      6'b100101 : begin
        _zz_2821_ = int_reg_array_34_37_imag;
        _zz_2822_ = int_reg_array_34_37_real;
      end
      6'b100110 : begin
        _zz_2821_ = int_reg_array_34_38_imag;
        _zz_2822_ = int_reg_array_34_38_real;
      end
      6'b100111 : begin
        _zz_2821_ = int_reg_array_34_39_imag;
        _zz_2822_ = int_reg_array_34_39_real;
      end
      6'b101000 : begin
        _zz_2821_ = int_reg_array_34_40_imag;
        _zz_2822_ = int_reg_array_34_40_real;
      end
      6'b101001 : begin
        _zz_2821_ = int_reg_array_34_41_imag;
        _zz_2822_ = int_reg_array_34_41_real;
      end
      6'b101010 : begin
        _zz_2821_ = int_reg_array_34_42_imag;
        _zz_2822_ = int_reg_array_34_42_real;
      end
      6'b101011 : begin
        _zz_2821_ = int_reg_array_34_43_imag;
        _zz_2822_ = int_reg_array_34_43_real;
      end
      6'b101100 : begin
        _zz_2821_ = int_reg_array_34_44_imag;
        _zz_2822_ = int_reg_array_34_44_real;
      end
      6'b101101 : begin
        _zz_2821_ = int_reg_array_34_45_imag;
        _zz_2822_ = int_reg_array_34_45_real;
      end
      6'b101110 : begin
        _zz_2821_ = int_reg_array_34_46_imag;
        _zz_2822_ = int_reg_array_34_46_real;
      end
      6'b101111 : begin
        _zz_2821_ = int_reg_array_34_47_imag;
        _zz_2822_ = int_reg_array_34_47_real;
      end
      6'b110000 : begin
        _zz_2821_ = int_reg_array_34_48_imag;
        _zz_2822_ = int_reg_array_34_48_real;
      end
      default : begin
        _zz_2821_ = int_reg_array_34_49_imag;
        _zz_2822_ = int_reg_array_34_49_real;
      end
    endcase
  end

  always @(*) begin
    case(_zz_1927_)
      6'b000000 : begin
        _zz_2823_ = int_reg_array_35_0_imag;
        _zz_2824_ = int_reg_array_35_0_real;
      end
      6'b000001 : begin
        _zz_2823_ = int_reg_array_35_1_imag;
        _zz_2824_ = int_reg_array_35_1_real;
      end
      6'b000010 : begin
        _zz_2823_ = int_reg_array_35_2_imag;
        _zz_2824_ = int_reg_array_35_2_real;
      end
      6'b000011 : begin
        _zz_2823_ = int_reg_array_35_3_imag;
        _zz_2824_ = int_reg_array_35_3_real;
      end
      6'b000100 : begin
        _zz_2823_ = int_reg_array_35_4_imag;
        _zz_2824_ = int_reg_array_35_4_real;
      end
      6'b000101 : begin
        _zz_2823_ = int_reg_array_35_5_imag;
        _zz_2824_ = int_reg_array_35_5_real;
      end
      6'b000110 : begin
        _zz_2823_ = int_reg_array_35_6_imag;
        _zz_2824_ = int_reg_array_35_6_real;
      end
      6'b000111 : begin
        _zz_2823_ = int_reg_array_35_7_imag;
        _zz_2824_ = int_reg_array_35_7_real;
      end
      6'b001000 : begin
        _zz_2823_ = int_reg_array_35_8_imag;
        _zz_2824_ = int_reg_array_35_8_real;
      end
      6'b001001 : begin
        _zz_2823_ = int_reg_array_35_9_imag;
        _zz_2824_ = int_reg_array_35_9_real;
      end
      6'b001010 : begin
        _zz_2823_ = int_reg_array_35_10_imag;
        _zz_2824_ = int_reg_array_35_10_real;
      end
      6'b001011 : begin
        _zz_2823_ = int_reg_array_35_11_imag;
        _zz_2824_ = int_reg_array_35_11_real;
      end
      6'b001100 : begin
        _zz_2823_ = int_reg_array_35_12_imag;
        _zz_2824_ = int_reg_array_35_12_real;
      end
      6'b001101 : begin
        _zz_2823_ = int_reg_array_35_13_imag;
        _zz_2824_ = int_reg_array_35_13_real;
      end
      6'b001110 : begin
        _zz_2823_ = int_reg_array_35_14_imag;
        _zz_2824_ = int_reg_array_35_14_real;
      end
      6'b001111 : begin
        _zz_2823_ = int_reg_array_35_15_imag;
        _zz_2824_ = int_reg_array_35_15_real;
      end
      6'b010000 : begin
        _zz_2823_ = int_reg_array_35_16_imag;
        _zz_2824_ = int_reg_array_35_16_real;
      end
      6'b010001 : begin
        _zz_2823_ = int_reg_array_35_17_imag;
        _zz_2824_ = int_reg_array_35_17_real;
      end
      6'b010010 : begin
        _zz_2823_ = int_reg_array_35_18_imag;
        _zz_2824_ = int_reg_array_35_18_real;
      end
      6'b010011 : begin
        _zz_2823_ = int_reg_array_35_19_imag;
        _zz_2824_ = int_reg_array_35_19_real;
      end
      6'b010100 : begin
        _zz_2823_ = int_reg_array_35_20_imag;
        _zz_2824_ = int_reg_array_35_20_real;
      end
      6'b010101 : begin
        _zz_2823_ = int_reg_array_35_21_imag;
        _zz_2824_ = int_reg_array_35_21_real;
      end
      6'b010110 : begin
        _zz_2823_ = int_reg_array_35_22_imag;
        _zz_2824_ = int_reg_array_35_22_real;
      end
      6'b010111 : begin
        _zz_2823_ = int_reg_array_35_23_imag;
        _zz_2824_ = int_reg_array_35_23_real;
      end
      6'b011000 : begin
        _zz_2823_ = int_reg_array_35_24_imag;
        _zz_2824_ = int_reg_array_35_24_real;
      end
      6'b011001 : begin
        _zz_2823_ = int_reg_array_35_25_imag;
        _zz_2824_ = int_reg_array_35_25_real;
      end
      6'b011010 : begin
        _zz_2823_ = int_reg_array_35_26_imag;
        _zz_2824_ = int_reg_array_35_26_real;
      end
      6'b011011 : begin
        _zz_2823_ = int_reg_array_35_27_imag;
        _zz_2824_ = int_reg_array_35_27_real;
      end
      6'b011100 : begin
        _zz_2823_ = int_reg_array_35_28_imag;
        _zz_2824_ = int_reg_array_35_28_real;
      end
      6'b011101 : begin
        _zz_2823_ = int_reg_array_35_29_imag;
        _zz_2824_ = int_reg_array_35_29_real;
      end
      6'b011110 : begin
        _zz_2823_ = int_reg_array_35_30_imag;
        _zz_2824_ = int_reg_array_35_30_real;
      end
      6'b011111 : begin
        _zz_2823_ = int_reg_array_35_31_imag;
        _zz_2824_ = int_reg_array_35_31_real;
      end
      6'b100000 : begin
        _zz_2823_ = int_reg_array_35_32_imag;
        _zz_2824_ = int_reg_array_35_32_real;
      end
      6'b100001 : begin
        _zz_2823_ = int_reg_array_35_33_imag;
        _zz_2824_ = int_reg_array_35_33_real;
      end
      6'b100010 : begin
        _zz_2823_ = int_reg_array_35_34_imag;
        _zz_2824_ = int_reg_array_35_34_real;
      end
      6'b100011 : begin
        _zz_2823_ = int_reg_array_35_35_imag;
        _zz_2824_ = int_reg_array_35_35_real;
      end
      6'b100100 : begin
        _zz_2823_ = int_reg_array_35_36_imag;
        _zz_2824_ = int_reg_array_35_36_real;
      end
      6'b100101 : begin
        _zz_2823_ = int_reg_array_35_37_imag;
        _zz_2824_ = int_reg_array_35_37_real;
      end
      6'b100110 : begin
        _zz_2823_ = int_reg_array_35_38_imag;
        _zz_2824_ = int_reg_array_35_38_real;
      end
      6'b100111 : begin
        _zz_2823_ = int_reg_array_35_39_imag;
        _zz_2824_ = int_reg_array_35_39_real;
      end
      6'b101000 : begin
        _zz_2823_ = int_reg_array_35_40_imag;
        _zz_2824_ = int_reg_array_35_40_real;
      end
      6'b101001 : begin
        _zz_2823_ = int_reg_array_35_41_imag;
        _zz_2824_ = int_reg_array_35_41_real;
      end
      6'b101010 : begin
        _zz_2823_ = int_reg_array_35_42_imag;
        _zz_2824_ = int_reg_array_35_42_real;
      end
      6'b101011 : begin
        _zz_2823_ = int_reg_array_35_43_imag;
        _zz_2824_ = int_reg_array_35_43_real;
      end
      6'b101100 : begin
        _zz_2823_ = int_reg_array_35_44_imag;
        _zz_2824_ = int_reg_array_35_44_real;
      end
      6'b101101 : begin
        _zz_2823_ = int_reg_array_35_45_imag;
        _zz_2824_ = int_reg_array_35_45_real;
      end
      6'b101110 : begin
        _zz_2823_ = int_reg_array_35_46_imag;
        _zz_2824_ = int_reg_array_35_46_real;
      end
      6'b101111 : begin
        _zz_2823_ = int_reg_array_35_47_imag;
        _zz_2824_ = int_reg_array_35_47_real;
      end
      6'b110000 : begin
        _zz_2823_ = int_reg_array_35_48_imag;
        _zz_2824_ = int_reg_array_35_48_real;
      end
      default : begin
        _zz_2823_ = int_reg_array_35_49_imag;
        _zz_2824_ = int_reg_array_35_49_real;
      end
    endcase
  end

  always @(*) begin
    case(_zz_1982_)
      6'b000000 : begin
        _zz_2825_ = int_reg_array_36_0_imag;
        _zz_2826_ = int_reg_array_36_0_real;
      end
      6'b000001 : begin
        _zz_2825_ = int_reg_array_36_1_imag;
        _zz_2826_ = int_reg_array_36_1_real;
      end
      6'b000010 : begin
        _zz_2825_ = int_reg_array_36_2_imag;
        _zz_2826_ = int_reg_array_36_2_real;
      end
      6'b000011 : begin
        _zz_2825_ = int_reg_array_36_3_imag;
        _zz_2826_ = int_reg_array_36_3_real;
      end
      6'b000100 : begin
        _zz_2825_ = int_reg_array_36_4_imag;
        _zz_2826_ = int_reg_array_36_4_real;
      end
      6'b000101 : begin
        _zz_2825_ = int_reg_array_36_5_imag;
        _zz_2826_ = int_reg_array_36_5_real;
      end
      6'b000110 : begin
        _zz_2825_ = int_reg_array_36_6_imag;
        _zz_2826_ = int_reg_array_36_6_real;
      end
      6'b000111 : begin
        _zz_2825_ = int_reg_array_36_7_imag;
        _zz_2826_ = int_reg_array_36_7_real;
      end
      6'b001000 : begin
        _zz_2825_ = int_reg_array_36_8_imag;
        _zz_2826_ = int_reg_array_36_8_real;
      end
      6'b001001 : begin
        _zz_2825_ = int_reg_array_36_9_imag;
        _zz_2826_ = int_reg_array_36_9_real;
      end
      6'b001010 : begin
        _zz_2825_ = int_reg_array_36_10_imag;
        _zz_2826_ = int_reg_array_36_10_real;
      end
      6'b001011 : begin
        _zz_2825_ = int_reg_array_36_11_imag;
        _zz_2826_ = int_reg_array_36_11_real;
      end
      6'b001100 : begin
        _zz_2825_ = int_reg_array_36_12_imag;
        _zz_2826_ = int_reg_array_36_12_real;
      end
      6'b001101 : begin
        _zz_2825_ = int_reg_array_36_13_imag;
        _zz_2826_ = int_reg_array_36_13_real;
      end
      6'b001110 : begin
        _zz_2825_ = int_reg_array_36_14_imag;
        _zz_2826_ = int_reg_array_36_14_real;
      end
      6'b001111 : begin
        _zz_2825_ = int_reg_array_36_15_imag;
        _zz_2826_ = int_reg_array_36_15_real;
      end
      6'b010000 : begin
        _zz_2825_ = int_reg_array_36_16_imag;
        _zz_2826_ = int_reg_array_36_16_real;
      end
      6'b010001 : begin
        _zz_2825_ = int_reg_array_36_17_imag;
        _zz_2826_ = int_reg_array_36_17_real;
      end
      6'b010010 : begin
        _zz_2825_ = int_reg_array_36_18_imag;
        _zz_2826_ = int_reg_array_36_18_real;
      end
      6'b010011 : begin
        _zz_2825_ = int_reg_array_36_19_imag;
        _zz_2826_ = int_reg_array_36_19_real;
      end
      6'b010100 : begin
        _zz_2825_ = int_reg_array_36_20_imag;
        _zz_2826_ = int_reg_array_36_20_real;
      end
      6'b010101 : begin
        _zz_2825_ = int_reg_array_36_21_imag;
        _zz_2826_ = int_reg_array_36_21_real;
      end
      6'b010110 : begin
        _zz_2825_ = int_reg_array_36_22_imag;
        _zz_2826_ = int_reg_array_36_22_real;
      end
      6'b010111 : begin
        _zz_2825_ = int_reg_array_36_23_imag;
        _zz_2826_ = int_reg_array_36_23_real;
      end
      6'b011000 : begin
        _zz_2825_ = int_reg_array_36_24_imag;
        _zz_2826_ = int_reg_array_36_24_real;
      end
      6'b011001 : begin
        _zz_2825_ = int_reg_array_36_25_imag;
        _zz_2826_ = int_reg_array_36_25_real;
      end
      6'b011010 : begin
        _zz_2825_ = int_reg_array_36_26_imag;
        _zz_2826_ = int_reg_array_36_26_real;
      end
      6'b011011 : begin
        _zz_2825_ = int_reg_array_36_27_imag;
        _zz_2826_ = int_reg_array_36_27_real;
      end
      6'b011100 : begin
        _zz_2825_ = int_reg_array_36_28_imag;
        _zz_2826_ = int_reg_array_36_28_real;
      end
      6'b011101 : begin
        _zz_2825_ = int_reg_array_36_29_imag;
        _zz_2826_ = int_reg_array_36_29_real;
      end
      6'b011110 : begin
        _zz_2825_ = int_reg_array_36_30_imag;
        _zz_2826_ = int_reg_array_36_30_real;
      end
      6'b011111 : begin
        _zz_2825_ = int_reg_array_36_31_imag;
        _zz_2826_ = int_reg_array_36_31_real;
      end
      6'b100000 : begin
        _zz_2825_ = int_reg_array_36_32_imag;
        _zz_2826_ = int_reg_array_36_32_real;
      end
      6'b100001 : begin
        _zz_2825_ = int_reg_array_36_33_imag;
        _zz_2826_ = int_reg_array_36_33_real;
      end
      6'b100010 : begin
        _zz_2825_ = int_reg_array_36_34_imag;
        _zz_2826_ = int_reg_array_36_34_real;
      end
      6'b100011 : begin
        _zz_2825_ = int_reg_array_36_35_imag;
        _zz_2826_ = int_reg_array_36_35_real;
      end
      6'b100100 : begin
        _zz_2825_ = int_reg_array_36_36_imag;
        _zz_2826_ = int_reg_array_36_36_real;
      end
      6'b100101 : begin
        _zz_2825_ = int_reg_array_36_37_imag;
        _zz_2826_ = int_reg_array_36_37_real;
      end
      6'b100110 : begin
        _zz_2825_ = int_reg_array_36_38_imag;
        _zz_2826_ = int_reg_array_36_38_real;
      end
      6'b100111 : begin
        _zz_2825_ = int_reg_array_36_39_imag;
        _zz_2826_ = int_reg_array_36_39_real;
      end
      6'b101000 : begin
        _zz_2825_ = int_reg_array_36_40_imag;
        _zz_2826_ = int_reg_array_36_40_real;
      end
      6'b101001 : begin
        _zz_2825_ = int_reg_array_36_41_imag;
        _zz_2826_ = int_reg_array_36_41_real;
      end
      6'b101010 : begin
        _zz_2825_ = int_reg_array_36_42_imag;
        _zz_2826_ = int_reg_array_36_42_real;
      end
      6'b101011 : begin
        _zz_2825_ = int_reg_array_36_43_imag;
        _zz_2826_ = int_reg_array_36_43_real;
      end
      6'b101100 : begin
        _zz_2825_ = int_reg_array_36_44_imag;
        _zz_2826_ = int_reg_array_36_44_real;
      end
      6'b101101 : begin
        _zz_2825_ = int_reg_array_36_45_imag;
        _zz_2826_ = int_reg_array_36_45_real;
      end
      6'b101110 : begin
        _zz_2825_ = int_reg_array_36_46_imag;
        _zz_2826_ = int_reg_array_36_46_real;
      end
      6'b101111 : begin
        _zz_2825_ = int_reg_array_36_47_imag;
        _zz_2826_ = int_reg_array_36_47_real;
      end
      6'b110000 : begin
        _zz_2825_ = int_reg_array_36_48_imag;
        _zz_2826_ = int_reg_array_36_48_real;
      end
      default : begin
        _zz_2825_ = int_reg_array_36_49_imag;
        _zz_2826_ = int_reg_array_36_49_real;
      end
    endcase
  end

  always @(*) begin
    case(_zz_2037_)
      6'b000000 : begin
        _zz_2827_ = int_reg_array_37_0_imag;
        _zz_2828_ = int_reg_array_37_0_real;
      end
      6'b000001 : begin
        _zz_2827_ = int_reg_array_37_1_imag;
        _zz_2828_ = int_reg_array_37_1_real;
      end
      6'b000010 : begin
        _zz_2827_ = int_reg_array_37_2_imag;
        _zz_2828_ = int_reg_array_37_2_real;
      end
      6'b000011 : begin
        _zz_2827_ = int_reg_array_37_3_imag;
        _zz_2828_ = int_reg_array_37_3_real;
      end
      6'b000100 : begin
        _zz_2827_ = int_reg_array_37_4_imag;
        _zz_2828_ = int_reg_array_37_4_real;
      end
      6'b000101 : begin
        _zz_2827_ = int_reg_array_37_5_imag;
        _zz_2828_ = int_reg_array_37_5_real;
      end
      6'b000110 : begin
        _zz_2827_ = int_reg_array_37_6_imag;
        _zz_2828_ = int_reg_array_37_6_real;
      end
      6'b000111 : begin
        _zz_2827_ = int_reg_array_37_7_imag;
        _zz_2828_ = int_reg_array_37_7_real;
      end
      6'b001000 : begin
        _zz_2827_ = int_reg_array_37_8_imag;
        _zz_2828_ = int_reg_array_37_8_real;
      end
      6'b001001 : begin
        _zz_2827_ = int_reg_array_37_9_imag;
        _zz_2828_ = int_reg_array_37_9_real;
      end
      6'b001010 : begin
        _zz_2827_ = int_reg_array_37_10_imag;
        _zz_2828_ = int_reg_array_37_10_real;
      end
      6'b001011 : begin
        _zz_2827_ = int_reg_array_37_11_imag;
        _zz_2828_ = int_reg_array_37_11_real;
      end
      6'b001100 : begin
        _zz_2827_ = int_reg_array_37_12_imag;
        _zz_2828_ = int_reg_array_37_12_real;
      end
      6'b001101 : begin
        _zz_2827_ = int_reg_array_37_13_imag;
        _zz_2828_ = int_reg_array_37_13_real;
      end
      6'b001110 : begin
        _zz_2827_ = int_reg_array_37_14_imag;
        _zz_2828_ = int_reg_array_37_14_real;
      end
      6'b001111 : begin
        _zz_2827_ = int_reg_array_37_15_imag;
        _zz_2828_ = int_reg_array_37_15_real;
      end
      6'b010000 : begin
        _zz_2827_ = int_reg_array_37_16_imag;
        _zz_2828_ = int_reg_array_37_16_real;
      end
      6'b010001 : begin
        _zz_2827_ = int_reg_array_37_17_imag;
        _zz_2828_ = int_reg_array_37_17_real;
      end
      6'b010010 : begin
        _zz_2827_ = int_reg_array_37_18_imag;
        _zz_2828_ = int_reg_array_37_18_real;
      end
      6'b010011 : begin
        _zz_2827_ = int_reg_array_37_19_imag;
        _zz_2828_ = int_reg_array_37_19_real;
      end
      6'b010100 : begin
        _zz_2827_ = int_reg_array_37_20_imag;
        _zz_2828_ = int_reg_array_37_20_real;
      end
      6'b010101 : begin
        _zz_2827_ = int_reg_array_37_21_imag;
        _zz_2828_ = int_reg_array_37_21_real;
      end
      6'b010110 : begin
        _zz_2827_ = int_reg_array_37_22_imag;
        _zz_2828_ = int_reg_array_37_22_real;
      end
      6'b010111 : begin
        _zz_2827_ = int_reg_array_37_23_imag;
        _zz_2828_ = int_reg_array_37_23_real;
      end
      6'b011000 : begin
        _zz_2827_ = int_reg_array_37_24_imag;
        _zz_2828_ = int_reg_array_37_24_real;
      end
      6'b011001 : begin
        _zz_2827_ = int_reg_array_37_25_imag;
        _zz_2828_ = int_reg_array_37_25_real;
      end
      6'b011010 : begin
        _zz_2827_ = int_reg_array_37_26_imag;
        _zz_2828_ = int_reg_array_37_26_real;
      end
      6'b011011 : begin
        _zz_2827_ = int_reg_array_37_27_imag;
        _zz_2828_ = int_reg_array_37_27_real;
      end
      6'b011100 : begin
        _zz_2827_ = int_reg_array_37_28_imag;
        _zz_2828_ = int_reg_array_37_28_real;
      end
      6'b011101 : begin
        _zz_2827_ = int_reg_array_37_29_imag;
        _zz_2828_ = int_reg_array_37_29_real;
      end
      6'b011110 : begin
        _zz_2827_ = int_reg_array_37_30_imag;
        _zz_2828_ = int_reg_array_37_30_real;
      end
      6'b011111 : begin
        _zz_2827_ = int_reg_array_37_31_imag;
        _zz_2828_ = int_reg_array_37_31_real;
      end
      6'b100000 : begin
        _zz_2827_ = int_reg_array_37_32_imag;
        _zz_2828_ = int_reg_array_37_32_real;
      end
      6'b100001 : begin
        _zz_2827_ = int_reg_array_37_33_imag;
        _zz_2828_ = int_reg_array_37_33_real;
      end
      6'b100010 : begin
        _zz_2827_ = int_reg_array_37_34_imag;
        _zz_2828_ = int_reg_array_37_34_real;
      end
      6'b100011 : begin
        _zz_2827_ = int_reg_array_37_35_imag;
        _zz_2828_ = int_reg_array_37_35_real;
      end
      6'b100100 : begin
        _zz_2827_ = int_reg_array_37_36_imag;
        _zz_2828_ = int_reg_array_37_36_real;
      end
      6'b100101 : begin
        _zz_2827_ = int_reg_array_37_37_imag;
        _zz_2828_ = int_reg_array_37_37_real;
      end
      6'b100110 : begin
        _zz_2827_ = int_reg_array_37_38_imag;
        _zz_2828_ = int_reg_array_37_38_real;
      end
      6'b100111 : begin
        _zz_2827_ = int_reg_array_37_39_imag;
        _zz_2828_ = int_reg_array_37_39_real;
      end
      6'b101000 : begin
        _zz_2827_ = int_reg_array_37_40_imag;
        _zz_2828_ = int_reg_array_37_40_real;
      end
      6'b101001 : begin
        _zz_2827_ = int_reg_array_37_41_imag;
        _zz_2828_ = int_reg_array_37_41_real;
      end
      6'b101010 : begin
        _zz_2827_ = int_reg_array_37_42_imag;
        _zz_2828_ = int_reg_array_37_42_real;
      end
      6'b101011 : begin
        _zz_2827_ = int_reg_array_37_43_imag;
        _zz_2828_ = int_reg_array_37_43_real;
      end
      6'b101100 : begin
        _zz_2827_ = int_reg_array_37_44_imag;
        _zz_2828_ = int_reg_array_37_44_real;
      end
      6'b101101 : begin
        _zz_2827_ = int_reg_array_37_45_imag;
        _zz_2828_ = int_reg_array_37_45_real;
      end
      6'b101110 : begin
        _zz_2827_ = int_reg_array_37_46_imag;
        _zz_2828_ = int_reg_array_37_46_real;
      end
      6'b101111 : begin
        _zz_2827_ = int_reg_array_37_47_imag;
        _zz_2828_ = int_reg_array_37_47_real;
      end
      6'b110000 : begin
        _zz_2827_ = int_reg_array_37_48_imag;
        _zz_2828_ = int_reg_array_37_48_real;
      end
      default : begin
        _zz_2827_ = int_reg_array_37_49_imag;
        _zz_2828_ = int_reg_array_37_49_real;
      end
    endcase
  end

  always @(*) begin
    case(_zz_2092_)
      6'b000000 : begin
        _zz_2829_ = int_reg_array_38_0_imag;
        _zz_2830_ = int_reg_array_38_0_real;
      end
      6'b000001 : begin
        _zz_2829_ = int_reg_array_38_1_imag;
        _zz_2830_ = int_reg_array_38_1_real;
      end
      6'b000010 : begin
        _zz_2829_ = int_reg_array_38_2_imag;
        _zz_2830_ = int_reg_array_38_2_real;
      end
      6'b000011 : begin
        _zz_2829_ = int_reg_array_38_3_imag;
        _zz_2830_ = int_reg_array_38_3_real;
      end
      6'b000100 : begin
        _zz_2829_ = int_reg_array_38_4_imag;
        _zz_2830_ = int_reg_array_38_4_real;
      end
      6'b000101 : begin
        _zz_2829_ = int_reg_array_38_5_imag;
        _zz_2830_ = int_reg_array_38_5_real;
      end
      6'b000110 : begin
        _zz_2829_ = int_reg_array_38_6_imag;
        _zz_2830_ = int_reg_array_38_6_real;
      end
      6'b000111 : begin
        _zz_2829_ = int_reg_array_38_7_imag;
        _zz_2830_ = int_reg_array_38_7_real;
      end
      6'b001000 : begin
        _zz_2829_ = int_reg_array_38_8_imag;
        _zz_2830_ = int_reg_array_38_8_real;
      end
      6'b001001 : begin
        _zz_2829_ = int_reg_array_38_9_imag;
        _zz_2830_ = int_reg_array_38_9_real;
      end
      6'b001010 : begin
        _zz_2829_ = int_reg_array_38_10_imag;
        _zz_2830_ = int_reg_array_38_10_real;
      end
      6'b001011 : begin
        _zz_2829_ = int_reg_array_38_11_imag;
        _zz_2830_ = int_reg_array_38_11_real;
      end
      6'b001100 : begin
        _zz_2829_ = int_reg_array_38_12_imag;
        _zz_2830_ = int_reg_array_38_12_real;
      end
      6'b001101 : begin
        _zz_2829_ = int_reg_array_38_13_imag;
        _zz_2830_ = int_reg_array_38_13_real;
      end
      6'b001110 : begin
        _zz_2829_ = int_reg_array_38_14_imag;
        _zz_2830_ = int_reg_array_38_14_real;
      end
      6'b001111 : begin
        _zz_2829_ = int_reg_array_38_15_imag;
        _zz_2830_ = int_reg_array_38_15_real;
      end
      6'b010000 : begin
        _zz_2829_ = int_reg_array_38_16_imag;
        _zz_2830_ = int_reg_array_38_16_real;
      end
      6'b010001 : begin
        _zz_2829_ = int_reg_array_38_17_imag;
        _zz_2830_ = int_reg_array_38_17_real;
      end
      6'b010010 : begin
        _zz_2829_ = int_reg_array_38_18_imag;
        _zz_2830_ = int_reg_array_38_18_real;
      end
      6'b010011 : begin
        _zz_2829_ = int_reg_array_38_19_imag;
        _zz_2830_ = int_reg_array_38_19_real;
      end
      6'b010100 : begin
        _zz_2829_ = int_reg_array_38_20_imag;
        _zz_2830_ = int_reg_array_38_20_real;
      end
      6'b010101 : begin
        _zz_2829_ = int_reg_array_38_21_imag;
        _zz_2830_ = int_reg_array_38_21_real;
      end
      6'b010110 : begin
        _zz_2829_ = int_reg_array_38_22_imag;
        _zz_2830_ = int_reg_array_38_22_real;
      end
      6'b010111 : begin
        _zz_2829_ = int_reg_array_38_23_imag;
        _zz_2830_ = int_reg_array_38_23_real;
      end
      6'b011000 : begin
        _zz_2829_ = int_reg_array_38_24_imag;
        _zz_2830_ = int_reg_array_38_24_real;
      end
      6'b011001 : begin
        _zz_2829_ = int_reg_array_38_25_imag;
        _zz_2830_ = int_reg_array_38_25_real;
      end
      6'b011010 : begin
        _zz_2829_ = int_reg_array_38_26_imag;
        _zz_2830_ = int_reg_array_38_26_real;
      end
      6'b011011 : begin
        _zz_2829_ = int_reg_array_38_27_imag;
        _zz_2830_ = int_reg_array_38_27_real;
      end
      6'b011100 : begin
        _zz_2829_ = int_reg_array_38_28_imag;
        _zz_2830_ = int_reg_array_38_28_real;
      end
      6'b011101 : begin
        _zz_2829_ = int_reg_array_38_29_imag;
        _zz_2830_ = int_reg_array_38_29_real;
      end
      6'b011110 : begin
        _zz_2829_ = int_reg_array_38_30_imag;
        _zz_2830_ = int_reg_array_38_30_real;
      end
      6'b011111 : begin
        _zz_2829_ = int_reg_array_38_31_imag;
        _zz_2830_ = int_reg_array_38_31_real;
      end
      6'b100000 : begin
        _zz_2829_ = int_reg_array_38_32_imag;
        _zz_2830_ = int_reg_array_38_32_real;
      end
      6'b100001 : begin
        _zz_2829_ = int_reg_array_38_33_imag;
        _zz_2830_ = int_reg_array_38_33_real;
      end
      6'b100010 : begin
        _zz_2829_ = int_reg_array_38_34_imag;
        _zz_2830_ = int_reg_array_38_34_real;
      end
      6'b100011 : begin
        _zz_2829_ = int_reg_array_38_35_imag;
        _zz_2830_ = int_reg_array_38_35_real;
      end
      6'b100100 : begin
        _zz_2829_ = int_reg_array_38_36_imag;
        _zz_2830_ = int_reg_array_38_36_real;
      end
      6'b100101 : begin
        _zz_2829_ = int_reg_array_38_37_imag;
        _zz_2830_ = int_reg_array_38_37_real;
      end
      6'b100110 : begin
        _zz_2829_ = int_reg_array_38_38_imag;
        _zz_2830_ = int_reg_array_38_38_real;
      end
      6'b100111 : begin
        _zz_2829_ = int_reg_array_38_39_imag;
        _zz_2830_ = int_reg_array_38_39_real;
      end
      6'b101000 : begin
        _zz_2829_ = int_reg_array_38_40_imag;
        _zz_2830_ = int_reg_array_38_40_real;
      end
      6'b101001 : begin
        _zz_2829_ = int_reg_array_38_41_imag;
        _zz_2830_ = int_reg_array_38_41_real;
      end
      6'b101010 : begin
        _zz_2829_ = int_reg_array_38_42_imag;
        _zz_2830_ = int_reg_array_38_42_real;
      end
      6'b101011 : begin
        _zz_2829_ = int_reg_array_38_43_imag;
        _zz_2830_ = int_reg_array_38_43_real;
      end
      6'b101100 : begin
        _zz_2829_ = int_reg_array_38_44_imag;
        _zz_2830_ = int_reg_array_38_44_real;
      end
      6'b101101 : begin
        _zz_2829_ = int_reg_array_38_45_imag;
        _zz_2830_ = int_reg_array_38_45_real;
      end
      6'b101110 : begin
        _zz_2829_ = int_reg_array_38_46_imag;
        _zz_2830_ = int_reg_array_38_46_real;
      end
      6'b101111 : begin
        _zz_2829_ = int_reg_array_38_47_imag;
        _zz_2830_ = int_reg_array_38_47_real;
      end
      6'b110000 : begin
        _zz_2829_ = int_reg_array_38_48_imag;
        _zz_2830_ = int_reg_array_38_48_real;
      end
      default : begin
        _zz_2829_ = int_reg_array_38_49_imag;
        _zz_2830_ = int_reg_array_38_49_real;
      end
    endcase
  end

  always @(*) begin
    case(_zz_2147_)
      6'b000000 : begin
        _zz_2831_ = int_reg_array_39_0_imag;
        _zz_2832_ = int_reg_array_39_0_real;
      end
      6'b000001 : begin
        _zz_2831_ = int_reg_array_39_1_imag;
        _zz_2832_ = int_reg_array_39_1_real;
      end
      6'b000010 : begin
        _zz_2831_ = int_reg_array_39_2_imag;
        _zz_2832_ = int_reg_array_39_2_real;
      end
      6'b000011 : begin
        _zz_2831_ = int_reg_array_39_3_imag;
        _zz_2832_ = int_reg_array_39_3_real;
      end
      6'b000100 : begin
        _zz_2831_ = int_reg_array_39_4_imag;
        _zz_2832_ = int_reg_array_39_4_real;
      end
      6'b000101 : begin
        _zz_2831_ = int_reg_array_39_5_imag;
        _zz_2832_ = int_reg_array_39_5_real;
      end
      6'b000110 : begin
        _zz_2831_ = int_reg_array_39_6_imag;
        _zz_2832_ = int_reg_array_39_6_real;
      end
      6'b000111 : begin
        _zz_2831_ = int_reg_array_39_7_imag;
        _zz_2832_ = int_reg_array_39_7_real;
      end
      6'b001000 : begin
        _zz_2831_ = int_reg_array_39_8_imag;
        _zz_2832_ = int_reg_array_39_8_real;
      end
      6'b001001 : begin
        _zz_2831_ = int_reg_array_39_9_imag;
        _zz_2832_ = int_reg_array_39_9_real;
      end
      6'b001010 : begin
        _zz_2831_ = int_reg_array_39_10_imag;
        _zz_2832_ = int_reg_array_39_10_real;
      end
      6'b001011 : begin
        _zz_2831_ = int_reg_array_39_11_imag;
        _zz_2832_ = int_reg_array_39_11_real;
      end
      6'b001100 : begin
        _zz_2831_ = int_reg_array_39_12_imag;
        _zz_2832_ = int_reg_array_39_12_real;
      end
      6'b001101 : begin
        _zz_2831_ = int_reg_array_39_13_imag;
        _zz_2832_ = int_reg_array_39_13_real;
      end
      6'b001110 : begin
        _zz_2831_ = int_reg_array_39_14_imag;
        _zz_2832_ = int_reg_array_39_14_real;
      end
      6'b001111 : begin
        _zz_2831_ = int_reg_array_39_15_imag;
        _zz_2832_ = int_reg_array_39_15_real;
      end
      6'b010000 : begin
        _zz_2831_ = int_reg_array_39_16_imag;
        _zz_2832_ = int_reg_array_39_16_real;
      end
      6'b010001 : begin
        _zz_2831_ = int_reg_array_39_17_imag;
        _zz_2832_ = int_reg_array_39_17_real;
      end
      6'b010010 : begin
        _zz_2831_ = int_reg_array_39_18_imag;
        _zz_2832_ = int_reg_array_39_18_real;
      end
      6'b010011 : begin
        _zz_2831_ = int_reg_array_39_19_imag;
        _zz_2832_ = int_reg_array_39_19_real;
      end
      6'b010100 : begin
        _zz_2831_ = int_reg_array_39_20_imag;
        _zz_2832_ = int_reg_array_39_20_real;
      end
      6'b010101 : begin
        _zz_2831_ = int_reg_array_39_21_imag;
        _zz_2832_ = int_reg_array_39_21_real;
      end
      6'b010110 : begin
        _zz_2831_ = int_reg_array_39_22_imag;
        _zz_2832_ = int_reg_array_39_22_real;
      end
      6'b010111 : begin
        _zz_2831_ = int_reg_array_39_23_imag;
        _zz_2832_ = int_reg_array_39_23_real;
      end
      6'b011000 : begin
        _zz_2831_ = int_reg_array_39_24_imag;
        _zz_2832_ = int_reg_array_39_24_real;
      end
      6'b011001 : begin
        _zz_2831_ = int_reg_array_39_25_imag;
        _zz_2832_ = int_reg_array_39_25_real;
      end
      6'b011010 : begin
        _zz_2831_ = int_reg_array_39_26_imag;
        _zz_2832_ = int_reg_array_39_26_real;
      end
      6'b011011 : begin
        _zz_2831_ = int_reg_array_39_27_imag;
        _zz_2832_ = int_reg_array_39_27_real;
      end
      6'b011100 : begin
        _zz_2831_ = int_reg_array_39_28_imag;
        _zz_2832_ = int_reg_array_39_28_real;
      end
      6'b011101 : begin
        _zz_2831_ = int_reg_array_39_29_imag;
        _zz_2832_ = int_reg_array_39_29_real;
      end
      6'b011110 : begin
        _zz_2831_ = int_reg_array_39_30_imag;
        _zz_2832_ = int_reg_array_39_30_real;
      end
      6'b011111 : begin
        _zz_2831_ = int_reg_array_39_31_imag;
        _zz_2832_ = int_reg_array_39_31_real;
      end
      6'b100000 : begin
        _zz_2831_ = int_reg_array_39_32_imag;
        _zz_2832_ = int_reg_array_39_32_real;
      end
      6'b100001 : begin
        _zz_2831_ = int_reg_array_39_33_imag;
        _zz_2832_ = int_reg_array_39_33_real;
      end
      6'b100010 : begin
        _zz_2831_ = int_reg_array_39_34_imag;
        _zz_2832_ = int_reg_array_39_34_real;
      end
      6'b100011 : begin
        _zz_2831_ = int_reg_array_39_35_imag;
        _zz_2832_ = int_reg_array_39_35_real;
      end
      6'b100100 : begin
        _zz_2831_ = int_reg_array_39_36_imag;
        _zz_2832_ = int_reg_array_39_36_real;
      end
      6'b100101 : begin
        _zz_2831_ = int_reg_array_39_37_imag;
        _zz_2832_ = int_reg_array_39_37_real;
      end
      6'b100110 : begin
        _zz_2831_ = int_reg_array_39_38_imag;
        _zz_2832_ = int_reg_array_39_38_real;
      end
      6'b100111 : begin
        _zz_2831_ = int_reg_array_39_39_imag;
        _zz_2832_ = int_reg_array_39_39_real;
      end
      6'b101000 : begin
        _zz_2831_ = int_reg_array_39_40_imag;
        _zz_2832_ = int_reg_array_39_40_real;
      end
      6'b101001 : begin
        _zz_2831_ = int_reg_array_39_41_imag;
        _zz_2832_ = int_reg_array_39_41_real;
      end
      6'b101010 : begin
        _zz_2831_ = int_reg_array_39_42_imag;
        _zz_2832_ = int_reg_array_39_42_real;
      end
      6'b101011 : begin
        _zz_2831_ = int_reg_array_39_43_imag;
        _zz_2832_ = int_reg_array_39_43_real;
      end
      6'b101100 : begin
        _zz_2831_ = int_reg_array_39_44_imag;
        _zz_2832_ = int_reg_array_39_44_real;
      end
      6'b101101 : begin
        _zz_2831_ = int_reg_array_39_45_imag;
        _zz_2832_ = int_reg_array_39_45_real;
      end
      6'b101110 : begin
        _zz_2831_ = int_reg_array_39_46_imag;
        _zz_2832_ = int_reg_array_39_46_real;
      end
      6'b101111 : begin
        _zz_2831_ = int_reg_array_39_47_imag;
        _zz_2832_ = int_reg_array_39_47_real;
      end
      6'b110000 : begin
        _zz_2831_ = int_reg_array_39_48_imag;
        _zz_2832_ = int_reg_array_39_48_real;
      end
      default : begin
        _zz_2831_ = int_reg_array_39_49_imag;
        _zz_2832_ = int_reg_array_39_49_real;
      end
    endcase
  end

  always @(*) begin
    case(_zz_2202_)
      6'b000000 : begin
        _zz_2833_ = int_reg_array_40_0_imag;
        _zz_2834_ = int_reg_array_40_0_real;
      end
      6'b000001 : begin
        _zz_2833_ = int_reg_array_40_1_imag;
        _zz_2834_ = int_reg_array_40_1_real;
      end
      6'b000010 : begin
        _zz_2833_ = int_reg_array_40_2_imag;
        _zz_2834_ = int_reg_array_40_2_real;
      end
      6'b000011 : begin
        _zz_2833_ = int_reg_array_40_3_imag;
        _zz_2834_ = int_reg_array_40_3_real;
      end
      6'b000100 : begin
        _zz_2833_ = int_reg_array_40_4_imag;
        _zz_2834_ = int_reg_array_40_4_real;
      end
      6'b000101 : begin
        _zz_2833_ = int_reg_array_40_5_imag;
        _zz_2834_ = int_reg_array_40_5_real;
      end
      6'b000110 : begin
        _zz_2833_ = int_reg_array_40_6_imag;
        _zz_2834_ = int_reg_array_40_6_real;
      end
      6'b000111 : begin
        _zz_2833_ = int_reg_array_40_7_imag;
        _zz_2834_ = int_reg_array_40_7_real;
      end
      6'b001000 : begin
        _zz_2833_ = int_reg_array_40_8_imag;
        _zz_2834_ = int_reg_array_40_8_real;
      end
      6'b001001 : begin
        _zz_2833_ = int_reg_array_40_9_imag;
        _zz_2834_ = int_reg_array_40_9_real;
      end
      6'b001010 : begin
        _zz_2833_ = int_reg_array_40_10_imag;
        _zz_2834_ = int_reg_array_40_10_real;
      end
      6'b001011 : begin
        _zz_2833_ = int_reg_array_40_11_imag;
        _zz_2834_ = int_reg_array_40_11_real;
      end
      6'b001100 : begin
        _zz_2833_ = int_reg_array_40_12_imag;
        _zz_2834_ = int_reg_array_40_12_real;
      end
      6'b001101 : begin
        _zz_2833_ = int_reg_array_40_13_imag;
        _zz_2834_ = int_reg_array_40_13_real;
      end
      6'b001110 : begin
        _zz_2833_ = int_reg_array_40_14_imag;
        _zz_2834_ = int_reg_array_40_14_real;
      end
      6'b001111 : begin
        _zz_2833_ = int_reg_array_40_15_imag;
        _zz_2834_ = int_reg_array_40_15_real;
      end
      6'b010000 : begin
        _zz_2833_ = int_reg_array_40_16_imag;
        _zz_2834_ = int_reg_array_40_16_real;
      end
      6'b010001 : begin
        _zz_2833_ = int_reg_array_40_17_imag;
        _zz_2834_ = int_reg_array_40_17_real;
      end
      6'b010010 : begin
        _zz_2833_ = int_reg_array_40_18_imag;
        _zz_2834_ = int_reg_array_40_18_real;
      end
      6'b010011 : begin
        _zz_2833_ = int_reg_array_40_19_imag;
        _zz_2834_ = int_reg_array_40_19_real;
      end
      6'b010100 : begin
        _zz_2833_ = int_reg_array_40_20_imag;
        _zz_2834_ = int_reg_array_40_20_real;
      end
      6'b010101 : begin
        _zz_2833_ = int_reg_array_40_21_imag;
        _zz_2834_ = int_reg_array_40_21_real;
      end
      6'b010110 : begin
        _zz_2833_ = int_reg_array_40_22_imag;
        _zz_2834_ = int_reg_array_40_22_real;
      end
      6'b010111 : begin
        _zz_2833_ = int_reg_array_40_23_imag;
        _zz_2834_ = int_reg_array_40_23_real;
      end
      6'b011000 : begin
        _zz_2833_ = int_reg_array_40_24_imag;
        _zz_2834_ = int_reg_array_40_24_real;
      end
      6'b011001 : begin
        _zz_2833_ = int_reg_array_40_25_imag;
        _zz_2834_ = int_reg_array_40_25_real;
      end
      6'b011010 : begin
        _zz_2833_ = int_reg_array_40_26_imag;
        _zz_2834_ = int_reg_array_40_26_real;
      end
      6'b011011 : begin
        _zz_2833_ = int_reg_array_40_27_imag;
        _zz_2834_ = int_reg_array_40_27_real;
      end
      6'b011100 : begin
        _zz_2833_ = int_reg_array_40_28_imag;
        _zz_2834_ = int_reg_array_40_28_real;
      end
      6'b011101 : begin
        _zz_2833_ = int_reg_array_40_29_imag;
        _zz_2834_ = int_reg_array_40_29_real;
      end
      6'b011110 : begin
        _zz_2833_ = int_reg_array_40_30_imag;
        _zz_2834_ = int_reg_array_40_30_real;
      end
      6'b011111 : begin
        _zz_2833_ = int_reg_array_40_31_imag;
        _zz_2834_ = int_reg_array_40_31_real;
      end
      6'b100000 : begin
        _zz_2833_ = int_reg_array_40_32_imag;
        _zz_2834_ = int_reg_array_40_32_real;
      end
      6'b100001 : begin
        _zz_2833_ = int_reg_array_40_33_imag;
        _zz_2834_ = int_reg_array_40_33_real;
      end
      6'b100010 : begin
        _zz_2833_ = int_reg_array_40_34_imag;
        _zz_2834_ = int_reg_array_40_34_real;
      end
      6'b100011 : begin
        _zz_2833_ = int_reg_array_40_35_imag;
        _zz_2834_ = int_reg_array_40_35_real;
      end
      6'b100100 : begin
        _zz_2833_ = int_reg_array_40_36_imag;
        _zz_2834_ = int_reg_array_40_36_real;
      end
      6'b100101 : begin
        _zz_2833_ = int_reg_array_40_37_imag;
        _zz_2834_ = int_reg_array_40_37_real;
      end
      6'b100110 : begin
        _zz_2833_ = int_reg_array_40_38_imag;
        _zz_2834_ = int_reg_array_40_38_real;
      end
      6'b100111 : begin
        _zz_2833_ = int_reg_array_40_39_imag;
        _zz_2834_ = int_reg_array_40_39_real;
      end
      6'b101000 : begin
        _zz_2833_ = int_reg_array_40_40_imag;
        _zz_2834_ = int_reg_array_40_40_real;
      end
      6'b101001 : begin
        _zz_2833_ = int_reg_array_40_41_imag;
        _zz_2834_ = int_reg_array_40_41_real;
      end
      6'b101010 : begin
        _zz_2833_ = int_reg_array_40_42_imag;
        _zz_2834_ = int_reg_array_40_42_real;
      end
      6'b101011 : begin
        _zz_2833_ = int_reg_array_40_43_imag;
        _zz_2834_ = int_reg_array_40_43_real;
      end
      6'b101100 : begin
        _zz_2833_ = int_reg_array_40_44_imag;
        _zz_2834_ = int_reg_array_40_44_real;
      end
      6'b101101 : begin
        _zz_2833_ = int_reg_array_40_45_imag;
        _zz_2834_ = int_reg_array_40_45_real;
      end
      6'b101110 : begin
        _zz_2833_ = int_reg_array_40_46_imag;
        _zz_2834_ = int_reg_array_40_46_real;
      end
      6'b101111 : begin
        _zz_2833_ = int_reg_array_40_47_imag;
        _zz_2834_ = int_reg_array_40_47_real;
      end
      6'b110000 : begin
        _zz_2833_ = int_reg_array_40_48_imag;
        _zz_2834_ = int_reg_array_40_48_real;
      end
      default : begin
        _zz_2833_ = int_reg_array_40_49_imag;
        _zz_2834_ = int_reg_array_40_49_real;
      end
    endcase
  end

  always @(*) begin
    case(_zz_2257_)
      6'b000000 : begin
        _zz_2835_ = int_reg_array_41_0_imag;
        _zz_2836_ = int_reg_array_41_0_real;
      end
      6'b000001 : begin
        _zz_2835_ = int_reg_array_41_1_imag;
        _zz_2836_ = int_reg_array_41_1_real;
      end
      6'b000010 : begin
        _zz_2835_ = int_reg_array_41_2_imag;
        _zz_2836_ = int_reg_array_41_2_real;
      end
      6'b000011 : begin
        _zz_2835_ = int_reg_array_41_3_imag;
        _zz_2836_ = int_reg_array_41_3_real;
      end
      6'b000100 : begin
        _zz_2835_ = int_reg_array_41_4_imag;
        _zz_2836_ = int_reg_array_41_4_real;
      end
      6'b000101 : begin
        _zz_2835_ = int_reg_array_41_5_imag;
        _zz_2836_ = int_reg_array_41_5_real;
      end
      6'b000110 : begin
        _zz_2835_ = int_reg_array_41_6_imag;
        _zz_2836_ = int_reg_array_41_6_real;
      end
      6'b000111 : begin
        _zz_2835_ = int_reg_array_41_7_imag;
        _zz_2836_ = int_reg_array_41_7_real;
      end
      6'b001000 : begin
        _zz_2835_ = int_reg_array_41_8_imag;
        _zz_2836_ = int_reg_array_41_8_real;
      end
      6'b001001 : begin
        _zz_2835_ = int_reg_array_41_9_imag;
        _zz_2836_ = int_reg_array_41_9_real;
      end
      6'b001010 : begin
        _zz_2835_ = int_reg_array_41_10_imag;
        _zz_2836_ = int_reg_array_41_10_real;
      end
      6'b001011 : begin
        _zz_2835_ = int_reg_array_41_11_imag;
        _zz_2836_ = int_reg_array_41_11_real;
      end
      6'b001100 : begin
        _zz_2835_ = int_reg_array_41_12_imag;
        _zz_2836_ = int_reg_array_41_12_real;
      end
      6'b001101 : begin
        _zz_2835_ = int_reg_array_41_13_imag;
        _zz_2836_ = int_reg_array_41_13_real;
      end
      6'b001110 : begin
        _zz_2835_ = int_reg_array_41_14_imag;
        _zz_2836_ = int_reg_array_41_14_real;
      end
      6'b001111 : begin
        _zz_2835_ = int_reg_array_41_15_imag;
        _zz_2836_ = int_reg_array_41_15_real;
      end
      6'b010000 : begin
        _zz_2835_ = int_reg_array_41_16_imag;
        _zz_2836_ = int_reg_array_41_16_real;
      end
      6'b010001 : begin
        _zz_2835_ = int_reg_array_41_17_imag;
        _zz_2836_ = int_reg_array_41_17_real;
      end
      6'b010010 : begin
        _zz_2835_ = int_reg_array_41_18_imag;
        _zz_2836_ = int_reg_array_41_18_real;
      end
      6'b010011 : begin
        _zz_2835_ = int_reg_array_41_19_imag;
        _zz_2836_ = int_reg_array_41_19_real;
      end
      6'b010100 : begin
        _zz_2835_ = int_reg_array_41_20_imag;
        _zz_2836_ = int_reg_array_41_20_real;
      end
      6'b010101 : begin
        _zz_2835_ = int_reg_array_41_21_imag;
        _zz_2836_ = int_reg_array_41_21_real;
      end
      6'b010110 : begin
        _zz_2835_ = int_reg_array_41_22_imag;
        _zz_2836_ = int_reg_array_41_22_real;
      end
      6'b010111 : begin
        _zz_2835_ = int_reg_array_41_23_imag;
        _zz_2836_ = int_reg_array_41_23_real;
      end
      6'b011000 : begin
        _zz_2835_ = int_reg_array_41_24_imag;
        _zz_2836_ = int_reg_array_41_24_real;
      end
      6'b011001 : begin
        _zz_2835_ = int_reg_array_41_25_imag;
        _zz_2836_ = int_reg_array_41_25_real;
      end
      6'b011010 : begin
        _zz_2835_ = int_reg_array_41_26_imag;
        _zz_2836_ = int_reg_array_41_26_real;
      end
      6'b011011 : begin
        _zz_2835_ = int_reg_array_41_27_imag;
        _zz_2836_ = int_reg_array_41_27_real;
      end
      6'b011100 : begin
        _zz_2835_ = int_reg_array_41_28_imag;
        _zz_2836_ = int_reg_array_41_28_real;
      end
      6'b011101 : begin
        _zz_2835_ = int_reg_array_41_29_imag;
        _zz_2836_ = int_reg_array_41_29_real;
      end
      6'b011110 : begin
        _zz_2835_ = int_reg_array_41_30_imag;
        _zz_2836_ = int_reg_array_41_30_real;
      end
      6'b011111 : begin
        _zz_2835_ = int_reg_array_41_31_imag;
        _zz_2836_ = int_reg_array_41_31_real;
      end
      6'b100000 : begin
        _zz_2835_ = int_reg_array_41_32_imag;
        _zz_2836_ = int_reg_array_41_32_real;
      end
      6'b100001 : begin
        _zz_2835_ = int_reg_array_41_33_imag;
        _zz_2836_ = int_reg_array_41_33_real;
      end
      6'b100010 : begin
        _zz_2835_ = int_reg_array_41_34_imag;
        _zz_2836_ = int_reg_array_41_34_real;
      end
      6'b100011 : begin
        _zz_2835_ = int_reg_array_41_35_imag;
        _zz_2836_ = int_reg_array_41_35_real;
      end
      6'b100100 : begin
        _zz_2835_ = int_reg_array_41_36_imag;
        _zz_2836_ = int_reg_array_41_36_real;
      end
      6'b100101 : begin
        _zz_2835_ = int_reg_array_41_37_imag;
        _zz_2836_ = int_reg_array_41_37_real;
      end
      6'b100110 : begin
        _zz_2835_ = int_reg_array_41_38_imag;
        _zz_2836_ = int_reg_array_41_38_real;
      end
      6'b100111 : begin
        _zz_2835_ = int_reg_array_41_39_imag;
        _zz_2836_ = int_reg_array_41_39_real;
      end
      6'b101000 : begin
        _zz_2835_ = int_reg_array_41_40_imag;
        _zz_2836_ = int_reg_array_41_40_real;
      end
      6'b101001 : begin
        _zz_2835_ = int_reg_array_41_41_imag;
        _zz_2836_ = int_reg_array_41_41_real;
      end
      6'b101010 : begin
        _zz_2835_ = int_reg_array_41_42_imag;
        _zz_2836_ = int_reg_array_41_42_real;
      end
      6'b101011 : begin
        _zz_2835_ = int_reg_array_41_43_imag;
        _zz_2836_ = int_reg_array_41_43_real;
      end
      6'b101100 : begin
        _zz_2835_ = int_reg_array_41_44_imag;
        _zz_2836_ = int_reg_array_41_44_real;
      end
      6'b101101 : begin
        _zz_2835_ = int_reg_array_41_45_imag;
        _zz_2836_ = int_reg_array_41_45_real;
      end
      6'b101110 : begin
        _zz_2835_ = int_reg_array_41_46_imag;
        _zz_2836_ = int_reg_array_41_46_real;
      end
      6'b101111 : begin
        _zz_2835_ = int_reg_array_41_47_imag;
        _zz_2836_ = int_reg_array_41_47_real;
      end
      6'b110000 : begin
        _zz_2835_ = int_reg_array_41_48_imag;
        _zz_2836_ = int_reg_array_41_48_real;
      end
      default : begin
        _zz_2835_ = int_reg_array_41_49_imag;
        _zz_2836_ = int_reg_array_41_49_real;
      end
    endcase
  end

  always @(*) begin
    case(_zz_2312_)
      6'b000000 : begin
        _zz_2837_ = int_reg_array_42_0_imag;
        _zz_2838_ = int_reg_array_42_0_real;
      end
      6'b000001 : begin
        _zz_2837_ = int_reg_array_42_1_imag;
        _zz_2838_ = int_reg_array_42_1_real;
      end
      6'b000010 : begin
        _zz_2837_ = int_reg_array_42_2_imag;
        _zz_2838_ = int_reg_array_42_2_real;
      end
      6'b000011 : begin
        _zz_2837_ = int_reg_array_42_3_imag;
        _zz_2838_ = int_reg_array_42_3_real;
      end
      6'b000100 : begin
        _zz_2837_ = int_reg_array_42_4_imag;
        _zz_2838_ = int_reg_array_42_4_real;
      end
      6'b000101 : begin
        _zz_2837_ = int_reg_array_42_5_imag;
        _zz_2838_ = int_reg_array_42_5_real;
      end
      6'b000110 : begin
        _zz_2837_ = int_reg_array_42_6_imag;
        _zz_2838_ = int_reg_array_42_6_real;
      end
      6'b000111 : begin
        _zz_2837_ = int_reg_array_42_7_imag;
        _zz_2838_ = int_reg_array_42_7_real;
      end
      6'b001000 : begin
        _zz_2837_ = int_reg_array_42_8_imag;
        _zz_2838_ = int_reg_array_42_8_real;
      end
      6'b001001 : begin
        _zz_2837_ = int_reg_array_42_9_imag;
        _zz_2838_ = int_reg_array_42_9_real;
      end
      6'b001010 : begin
        _zz_2837_ = int_reg_array_42_10_imag;
        _zz_2838_ = int_reg_array_42_10_real;
      end
      6'b001011 : begin
        _zz_2837_ = int_reg_array_42_11_imag;
        _zz_2838_ = int_reg_array_42_11_real;
      end
      6'b001100 : begin
        _zz_2837_ = int_reg_array_42_12_imag;
        _zz_2838_ = int_reg_array_42_12_real;
      end
      6'b001101 : begin
        _zz_2837_ = int_reg_array_42_13_imag;
        _zz_2838_ = int_reg_array_42_13_real;
      end
      6'b001110 : begin
        _zz_2837_ = int_reg_array_42_14_imag;
        _zz_2838_ = int_reg_array_42_14_real;
      end
      6'b001111 : begin
        _zz_2837_ = int_reg_array_42_15_imag;
        _zz_2838_ = int_reg_array_42_15_real;
      end
      6'b010000 : begin
        _zz_2837_ = int_reg_array_42_16_imag;
        _zz_2838_ = int_reg_array_42_16_real;
      end
      6'b010001 : begin
        _zz_2837_ = int_reg_array_42_17_imag;
        _zz_2838_ = int_reg_array_42_17_real;
      end
      6'b010010 : begin
        _zz_2837_ = int_reg_array_42_18_imag;
        _zz_2838_ = int_reg_array_42_18_real;
      end
      6'b010011 : begin
        _zz_2837_ = int_reg_array_42_19_imag;
        _zz_2838_ = int_reg_array_42_19_real;
      end
      6'b010100 : begin
        _zz_2837_ = int_reg_array_42_20_imag;
        _zz_2838_ = int_reg_array_42_20_real;
      end
      6'b010101 : begin
        _zz_2837_ = int_reg_array_42_21_imag;
        _zz_2838_ = int_reg_array_42_21_real;
      end
      6'b010110 : begin
        _zz_2837_ = int_reg_array_42_22_imag;
        _zz_2838_ = int_reg_array_42_22_real;
      end
      6'b010111 : begin
        _zz_2837_ = int_reg_array_42_23_imag;
        _zz_2838_ = int_reg_array_42_23_real;
      end
      6'b011000 : begin
        _zz_2837_ = int_reg_array_42_24_imag;
        _zz_2838_ = int_reg_array_42_24_real;
      end
      6'b011001 : begin
        _zz_2837_ = int_reg_array_42_25_imag;
        _zz_2838_ = int_reg_array_42_25_real;
      end
      6'b011010 : begin
        _zz_2837_ = int_reg_array_42_26_imag;
        _zz_2838_ = int_reg_array_42_26_real;
      end
      6'b011011 : begin
        _zz_2837_ = int_reg_array_42_27_imag;
        _zz_2838_ = int_reg_array_42_27_real;
      end
      6'b011100 : begin
        _zz_2837_ = int_reg_array_42_28_imag;
        _zz_2838_ = int_reg_array_42_28_real;
      end
      6'b011101 : begin
        _zz_2837_ = int_reg_array_42_29_imag;
        _zz_2838_ = int_reg_array_42_29_real;
      end
      6'b011110 : begin
        _zz_2837_ = int_reg_array_42_30_imag;
        _zz_2838_ = int_reg_array_42_30_real;
      end
      6'b011111 : begin
        _zz_2837_ = int_reg_array_42_31_imag;
        _zz_2838_ = int_reg_array_42_31_real;
      end
      6'b100000 : begin
        _zz_2837_ = int_reg_array_42_32_imag;
        _zz_2838_ = int_reg_array_42_32_real;
      end
      6'b100001 : begin
        _zz_2837_ = int_reg_array_42_33_imag;
        _zz_2838_ = int_reg_array_42_33_real;
      end
      6'b100010 : begin
        _zz_2837_ = int_reg_array_42_34_imag;
        _zz_2838_ = int_reg_array_42_34_real;
      end
      6'b100011 : begin
        _zz_2837_ = int_reg_array_42_35_imag;
        _zz_2838_ = int_reg_array_42_35_real;
      end
      6'b100100 : begin
        _zz_2837_ = int_reg_array_42_36_imag;
        _zz_2838_ = int_reg_array_42_36_real;
      end
      6'b100101 : begin
        _zz_2837_ = int_reg_array_42_37_imag;
        _zz_2838_ = int_reg_array_42_37_real;
      end
      6'b100110 : begin
        _zz_2837_ = int_reg_array_42_38_imag;
        _zz_2838_ = int_reg_array_42_38_real;
      end
      6'b100111 : begin
        _zz_2837_ = int_reg_array_42_39_imag;
        _zz_2838_ = int_reg_array_42_39_real;
      end
      6'b101000 : begin
        _zz_2837_ = int_reg_array_42_40_imag;
        _zz_2838_ = int_reg_array_42_40_real;
      end
      6'b101001 : begin
        _zz_2837_ = int_reg_array_42_41_imag;
        _zz_2838_ = int_reg_array_42_41_real;
      end
      6'b101010 : begin
        _zz_2837_ = int_reg_array_42_42_imag;
        _zz_2838_ = int_reg_array_42_42_real;
      end
      6'b101011 : begin
        _zz_2837_ = int_reg_array_42_43_imag;
        _zz_2838_ = int_reg_array_42_43_real;
      end
      6'b101100 : begin
        _zz_2837_ = int_reg_array_42_44_imag;
        _zz_2838_ = int_reg_array_42_44_real;
      end
      6'b101101 : begin
        _zz_2837_ = int_reg_array_42_45_imag;
        _zz_2838_ = int_reg_array_42_45_real;
      end
      6'b101110 : begin
        _zz_2837_ = int_reg_array_42_46_imag;
        _zz_2838_ = int_reg_array_42_46_real;
      end
      6'b101111 : begin
        _zz_2837_ = int_reg_array_42_47_imag;
        _zz_2838_ = int_reg_array_42_47_real;
      end
      6'b110000 : begin
        _zz_2837_ = int_reg_array_42_48_imag;
        _zz_2838_ = int_reg_array_42_48_real;
      end
      default : begin
        _zz_2837_ = int_reg_array_42_49_imag;
        _zz_2838_ = int_reg_array_42_49_real;
      end
    endcase
  end

  always @(*) begin
    case(_zz_2367_)
      6'b000000 : begin
        _zz_2839_ = int_reg_array_43_0_imag;
        _zz_2840_ = int_reg_array_43_0_real;
      end
      6'b000001 : begin
        _zz_2839_ = int_reg_array_43_1_imag;
        _zz_2840_ = int_reg_array_43_1_real;
      end
      6'b000010 : begin
        _zz_2839_ = int_reg_array_43_2_imag;
        _zz_2840_ = int_reg_array_43_2_real;
      end
      6'b000011 : begin
        _zz_2839_ = int_reg_array_43_3_imag;
        _zz_2840_ = int_reg_array_43_3_real;
      end
      6'b000100 : begin
        _zz_2839_ = int_reg_array_43_4_imag;
        _zz_2840_ = int_reg_array_43_4_real;
      end
      6'b000101 : begin
        _zz_2839_ = int_reg_array_43_5_imag;
        _zz_2840_ = int_reg_array_43_5_real;
      end
      6'b000110 : begin
        _zz_2839_ = int_reg_array_43_6_imag;
        _zz_2840_ = int_reg_array_43_6_real;
      end
      6'b000111 : begin
        _zz_2839_ = int_reg_array_43_7_imag;
        _zz_2840_ = int_reg_array_43_7_real;
      end
      6'b001000 : begin
        _zz_2839_ = int_reg_array_43_8_imag;
        _zz_2840_ = int_reg_array_43_8_real;
      end
      6'b001001 : begin
        _zz_2839_ = int_reg_array_43_9_imag;
        _zz_2840_ = int_reg_array_43_9_real;
      end
      6'b001010 : begin
        _zz_2839_ = int_reg_array_43_10_imag;
        _zz_2840_ = int_reg_array_43_10_real;
      end
      6'b001011 : begin
        _zz_2839_ = int_reg_array_43_11_imag;
        _zz_2840_ = int_reg_array_43_11_real;
      end
      6'b001100 : begin
        _zz_2839_ = int_reg_array_43_12_imag;
        _zz_2840_ = int_reg_array_43_12_real;
      end
      6'b001101 : begin
        _zz_2839_ = int_reg_array_43_13_imag;
        _zz_2840_ = int_reg_array_43_13_real;
      end
      6'b001110 : begin
        _zz_2839_ = int_reg_array_43_14_imag;
        _zz_2840_ = int_reg_array_43_14_real;
      end
      6'b001111 : begin
        _zz_2839_ = int_reg_array_43_15_imag;
        _zz_2840_ = int_reg_array_43_15_real;
      end
      6'b010000 : begin
        _zz_2839_ = int_reg_array_43_16_imag;
        _zz_2840_ = int_reg_array_43_16_real;
      end
      6'b010001 : begin
        _zz_2839_ = int_reg_array_43_17_imag;
        _zz_2840_ = int_reg_array_43_17_real;
      end
      6'b010010 : begin
        _zz_2839_ = int_reg_array_43_18_imag;
        _zz_2840_ = int_reg_array_43_18_real;
      end
      6'b010011 : begin
        _zz_2839_ = int_reg_array_43_19_imag;
        _zz_2840_ = int_reg_array_43_19_real;
      end
      6'b010100 : begin
        _zz_2839_ = int_reg_array_43_20_imag;
        _zz_2840_ = int_reg_array_43_20_real;
      end
      6'b010101 : begin
        _zz_2839_ = int_reg_array_43_21_imag;
        _zz_2840_ = int_reg_array_43_21_real;
      end
      6'b010110 : begin
        _zz_2839_ = int_reg_array_43_22_imag;
        _zz_2840_ = int_reg_array_43_22_real;
      end
      6'b010111 : begin
        _zz_2839_ = int_reg_array_43_23_imag;
        _zz_2840_ = int_reg_array_43_23_real;
      end
      6'b011000 : begin
        _zz_2839_ = int_reg_array_43_24_imag;
        _zz_2840_ = int_reg_array_43_24_real;
      end
      6'b011001 : begin
        _zz_2839_ = int_reg_array_43_25_imag;
        _zz_2840_ = int_reg_array_43_25_real;
      end
      6'b011010 : begin
        _zz_2839_ = int_reg_array_43_26_imag;
        _zz_2840_ = int_reg_array_43_26_real;
      end
      6'b011011 : begin
        _zz_2839_ = int_reg_array_43_27_imag;
        _zz_2840_ = int_reg_array_43_27_real;
      end
      6'b011100 : begin
        _zz_2839_ = int_reg_array_43_28_imag;
        _zz_2840_ = int_reg_array_43_28_real;
      end
      6'b011101 : begin
        _zz_2839_ = int_reg_array_43_29_imag;
        _zz_2840_ = int_reg_array_43_29_real;
      end
      6'b011110 : begin
        _zz_2839_ = int_reg_array_43_30_imag;
        _zz_2840_ = int_reg_array_43_30_real;
      end
      6'b011111 : begin
        _zz_2839_ = int_reg_array_43_31_imag;
        _zz_2840_ = int_reg_array_43_31_real;
      end
      6'b100000 : begin
        _zz_2839_ = int_reg_array_43_32_imag;
        _zz_2840_ = int_reg_array_43_32_real;
      end
      6'b100001 : begin
        _zz_2839_ = int_reg_array_43_33_imag;
        _zz_2840_ = int_reg_array_43_33_real;
      end
      6'b100010 : begin
        _zz_2839_ = int_reg_array_43_34_imag;
        _zz_2840_ = int_reg_array_43_34_real;
      end
      6'b100011 : begin
        _zz_2839_ = int_reg_array_43_35_imag;
        _zz_2840_ = int_reg_array_43_35_real;
      end
      6'b100100 : begin
        _zz_2839_ = int_reg_array_43_36_imag;
        _zz_2840_ = int_reg_array_43_36_real;
      end
      6'b100101 : begin
        _zz_2839_ = int_reg_array_43_37_imag;
        _zz_2840_ = int_reg_array_43_37_real;
      end
      6'b100110 : begin
        _zz_2839_ = int_reg_array_43_38_imag;
        _zz_2840_ = int_reg_array_43_38_real;
      end
      6'b100111 : begin
        _zz_2839_ = int_reg_array_43_39_imag;
        _zz_2840_ = int_reg_array_43_39_real;
      end
      6'b101000 : begin
        _zz_2839_ = int_reg_array_43_40_imag;
        _zz_2840_ = int_reg_array_43_40_real;
      end
      6'b101001 : begin
        _zz_2839_ = int_reg_array_43_41_imag;
        _zz_2840_ = int_reg_array_43_41_real;
      end
      6'b101010 : begin
        _zz_2839_ = int_reg_array_43_42_imag;
        _zz_2840_ = int_reg_array_43_42_real;
      end
      6'b101011 : begin
        _zz_2839_ = int_reg_array_43_43_imag;
        _zz_2840_ = int_reg_array_43_43_real;
      end
      6'b101100 : begin
        _zz_2839_ = int_reg_array_43_44_imag;
        _zz_2840_ = int_reg_array_43_44_real;
      end
      6'b101101 : begin
        _zz_2839_ = int_reg_array_43_45_imag;
        _zz_2840_ = int_reg_array_43_45_real;
      end
      6'b101110 : begin
        _zz_2839_ = int_reg_array_43_46_imag;
        _zz_2840_ = int_reg_array_43_46_real;
      end
      6'b101111 : begin
        _zz_2839_ = int_reg_array_43_47_imag;
        _zz_2840_ = int_reg_array_43_47_real;
      end
      6'b110000 : begin
        _zz_2839_ = int_reg_array_43_48_imag;
        _zz_2840_ = int_reg_array_43_48_real;
      end
      default : begin
        _zz_2839_ = int_reg_array_43_49_imag;
        _zz_2840_ = int_reg_array_43_49_real;
      end
    endcase
  end

  always @(*) begin
    case(_zz_2422_)
      6'b000000 : begin
        _zz_2841_ = int_reg_array_44_0_imag;
        _zz_2842_ = int_reg_array_44_0_real;
      end
      6'b000001 : begin
        _zz_2841_ = int_reg_array_44_1_imag;
        _zz_2842_ = int_reg_array_44_1_real;
      end
      6'b000010 : begin
        _zz_2841_ = int_reg_array_44_2_imag;
        _zz_2842_ = int_reg_array_44_2_real;
      end
      6'b000011 : begin
        _zz_2841_ = int_reg_array_44_3_imag;
        _zz_2842_ = int_reg_array_44_3_real;
      end
      6'b000100 : begin
        _zz_2841_ = int_reg_array_44_4_imag;
        _zz_2842_ = int_reg_array_44_4_real;
      end
      6'b000101 : begin
        _zz_2841_ = int_reg_array_44_5_imag;
        _zz_2842_ = int_reg_array_44_5_real;
      end
      6'b000110 : begin
        _zz_2841_ = int_reg_array_44_6_imag;
        _zz_2842_ = int_reg_array_44_6_real;
      end
      6'b000111 : begin
        _zz_2841_ = int_reg_array_44_7_imag;
        _zz_2842_ = int_reg_array_44_7_real;
      end
      6'b001000 : begin
        _zz_2841_ = int_reg_array_44_8_imag;
        _zz_2842_ = int_reg_array_44_8_real;
      end
      6'b001001 : begin
        _zz_2841_ = int_reg_array_44_9_imag;
        _zz_2842_ = int_reg_array_44_9_real;
      end
      6'b001010 : begin
        _zz_2841_ = int_reg_array_44_10_imag;
        _zz_2842_ = int_reg_array_44_10_real;
      end
      6'b001011 : begin
        _zz_2841_ = int_reg_array_44_11_imag;
        _zz_2842_ = int_reg_array_44_11_real;
      end
      6'b001100 : begin
        _zz_2841_ = int_reg_array_44_12_imag;
        _zz_2842_ = int_reg_array_44_12_real;
      end
      6'b001101 : begin
        _zz_2841_ = int_reg_array_44_13_imag;
        _zz_2842_ = int_reg_array_44_13_real;
      end
      6'b001110 : begin
        _zz_2841_ = int_reg_array_44_14_imag;
        _zz_2842_ = int_reg_array_44_14_real;
      end
      6'b001111 : begin
        _zz_2841_ = int_reg_array_44_15_imag;
        _zz_2842_ = int_reg_array_44_15_real;
      end
      6'b010000 : begin
        _zz_2841_ = int_reg_array_44_16_imag;
        _zz_2842_ = int_reg_array_44_16_real;
      end
      6'b010001 : begin
        _zz_2841_ = int_reg_array_44_17_imag;
        _zz_2842_ = int_reg_array_44_17_real;
      end
      6'b010010 : begin
        _zz_2841_ = int_reg_array_44_18_imag;
        _zz_2842_ = int_reg_array_44_18_real;
      end
      6'b010011 : begin
        _zz_2841_ = int_reg_array_44_19_imag;
        _zz_2842_ = int_reg_array_44_19_real;
      end
      6'b010100 : begin
        _zz_2841_ = int_reg_array_44_20_imag;
        _zz_2842_ = int_reg_array_44_20_real;
      end
      6'b010101 : begin
        _zz_2841_ = int_reg_array_44_21_imag;
        _zz_2842_ = int_reg_array_44_21_real;
      end
      6'b010110 : begin
        _zz_2841_ = int_reg_array_44_22_imag;
        _zz_2842_ = int_reg_array_44_22_real;
      end
      6'b010111 : begin
        _zz_2841_ = int_reg_array_44_23_imag;
        _zz_2842_ = int_reg_array_44_23_real;
      end
      6'b011000 : begin
        _zz_2841_ = int_reg_array_44_24_imag;
        _zz_2842_ = int_reg_array_44_24_real;
      end
      6'b011001 : begin
        _zz_2841_ = int_reg_array_44_25_imag;
        _zz_2842_ = int_reg_array_44_25_real;
      end
      6'b011010 : begin
        _zz_2841_ = int_reg_array_44_26_imag;
        _zz_2842_ = int_reg_array_44_26_real;
      end
      6'b011011 : begin
        _zz_2841_ = int_reg_array_44_27_imag;
        _zz_2842_ = int_reg_array_44_27_real;
      end
      6'b011100 : begin
        _zz_2841_ = int_reg_array_44_28_imag;
        _zz_2842_ = int_reg_array_44_28_real;
      end
      6'b011101 : begin
        _zz_2841_ = int_reg_array_44_29_imag;
        _zz_2842_ = int_reg_array_44_29_real;
      end
      6'b011110 : begin
        _zz_2841_ = int_reg_array_44_30_imag;
        _zz_2842_ = int_reg_array_44_30_real;
      end
      6'b011111 : begin
        _zz_2841_ = int_reg_array_44_31_imag;
        _zz_2842_ = int_reg_array_44_31_real;
      end
      6'b100000 : begin
        _zz_2841_ = int_reg_array_44_32_imag;
        _zz_2842_ = int_reg_array_44_32_real;
      end
      6'b100001 : begin
        _zz_2841_ = int_reg_array_44_33_imag;
        _zz_2842_ = int_reg_array_44_33_real;
      end
      6'b100010 : begin
        _zz_2841_ = int_reg_array_44_34_imag;
        _zz_2842_ = int_reg_array_44_34_real;
      end
      6'b100011 : begin
        _zz_2841_ = int_reg_array_44_35_imag;
        _zz_2842_ = int_reg_array_44_35_real;
      end
      6'b100100 : begin
        _zz_2841_ = int_reg_array_44_36_imag;
        _zz_2842_ = int_reg_array_44_36_real;
      end
      6'b100101 : begin
        _zz_2841_ = int_reg_array_44_37_imag;
        _zz_2842_ = int_reg_array_44_37_real;
      end
      6'b100110 : begin
        _zz_2841_ = int_reg_array_44_38_imag;
        _zz_2842_ = int_reg_array_44_38_real;
      end
      6'b100111 : begin
        _zz_2841_ = int_reg_array_44_39_imag;
        _zz_2842_ = int_reg_array_44_39_real;
      end
      6'b101000 : begin
        _zz_2841_ = int_reg_array_44_40_imag;
        _zz_2842_ = int_reg_array_44_40_real;
      end
      6'b101001 : begin
        _zz_2841_ = int_reg_array_44_41_imag;
        _zz_2842_ = int_reg_array_44_41_real;
      end
      6'b101010 : begin
        _zz_2841_ = int_reg_array_44_42_imag;
        _zz_2842_ = int_reg_array_44_42_real;
      end
      6'b101011 : begin
        _zz_2841_ = int_reg_array_44_43_imag;
        _zz_2842_ = int_reg_array_44_43_real;
      end
      6'b101100 : begin
        _zz_2841_ = int_reg_array_44_44_imag;
        _zz_2842_ = int_reg_array_44_44_real;
      end
      6'b101101 : begin
        _zz_2841_ = int_reg_array_44_45_imag;
        _zz_2842_ = int_reg_array_44_45_real;
      end
      6'b101110 : begin
        _zz_2841_ = int_reg_array_44_46_imag;
        _zz_2842_ = int_reg_array_44_46_real;
      end
      6'b101111 : begin
        _zz_2841_ = int_reg_array_44_47_imag;
        _zz_2842_ = int_reg_array_44_47_real;
      end
      6'b110000 : begin
        _zz_2841_ = int_reg_array_44_48_imag;
        _zz_2842_ = int_reg_array_44_48_real;
      end
      default : begin
        _zz_2841_ = int_reg_array_44_49_imag;
        _zz_2842_ = int_reg_array_44_49_real;
      end
    endcase
  end

  always @(*) begin
    case(_zz_2477_)
      6'b000000 : begin
        _zz_2843_ = int_reg_array_45_0_imag;
        _zz_2844_ = int_reg_array_45_0_real;
      end
      6'b000001 : begin
        _zz_2843_ = int_reg_array_45_1_imag;
        _zz_2844_ = int_reg_array_45_1_real;
      end
      6'b000010 : begin
        _zz_2843_ = int_reg_array_45_2_imag;
        _zz_2844_ = int_reg_array_45_2_real;
      end
      6'b000011 : begin
        _zz_2843_ = int_reg_array_45_3_imag;
        _zz_2844_ = int_reg_array_45_3_real;
      end
      6'b000100 : begin
        _zz_2843_ = int_reg_array_45_4_imag;
        _zz_2844_ = int_reg_array_45_4_real;
      end
      6'b000101 : begin
        _zz_2843_ = int_reg_array_45_5_imag;
        _zz_2844_ = int_reg_array_45_5_real;
      end
      6'b000110 : begin
        _zz_2843_ = int_reg_array_45_6_imag;
        _zz_2844_ = int_reg_array_45_6_real;
      end
      6'b000111 : begin
        _zz_2843_ = int_reg_array_45_7_imag;
        _zz_2844_ = int_reg_array_45_7_real;
      end
      6'b001000 : begin
        _zz_2843_ = int_reg_array_45_8_imag;
        _zz_2844_ = int_reg_array_45_8_real;
      end
      6'b001001 : begin
        _zz_2843_ = int_reg_array_45_9_imag;
        _zz_2844_ = int_reg_array_45_9_real;
      end
      6'b001010 : begin
        _zz_2843_ = int_reg_array_45_10_imag;
        _zz_2844_ = int_reg_array_45_10_real;
      end
      6'b001011 : begin
        _zz_2843_ = int_reg_array_45_11_imag;
        _zz_2844_ = int_reg_array_45_11_real;
      end
      6'b001100 : begin
        _zz_2843_ = int_reg_array_45_12_imag;
        _zz_2844_ = int_reg_array_45_12_real;
      end
      6'b001101 : begin
        _zz_2843_ = int_reg_array_45_13_imag;
        _zz_2844_ = int_reg_array_45_13_real;
      end
      6'b001110 : begin
        _zz_2843_ = int_reg_array_45_14_imag;
        _zz_2844_ = int_reg_array_45_14_real;
      end
      6'b001111 : begin
        _zz_2843_ = int_reg_array_45_15_imag;
        _zz_2844_ = int_reg_array_45_15_real;
      end
      6'b010000 : begin
        _zz_2843_ = int_reg_array_45_16_imag;
        _zz_2844_ = int_reg_array_45_16_real;
      end
      6'b010001 : begin
        _zz_2843_ = int_reg_array_45_17_imag;
        _zz_2844_ = int_reg_array_45_17_real;
      end
      6'b010010 : begin
        _zz_2843_ = int_reg_array_45_18_imag;
        _zz_2844_ = int_reg_array_45_18_real;
      end
      6'b010011 : begin
        _zz_2843_ = int_reg_array_45_19_imag;
        _zz_2844_ = int_reg_array_45_19_real;
      end
      6'b010100 : begin
        _zz_2843_ = int_reg_array_45_20_imag;
        _zz_2844_ = int_reg_array_45_20_real;
      end
      6'b010101 : begin
        _zz_2843_ = int_reg_array_45_21_imag;
        _zz_2844_ = int_reg_array_45_21_real;
      end
      6'b010110 : begin
        _zz_2843_ = int_reg_array_45_22_imag;
        _zz_2844_ = int_reg_array_45_22_real;
      end
      6'b010111 : begin
        _zz_2843_ = int_reg_array_45_23_imag;
        _zz_2844_ = int_reg_array_45_23_real;
      end
      6'b011000 : begin
        _zz_2843_ = int_reg_array_45_24_imag;
        _zz_2844_ = int_reg_array_45_24_real;
      end
      6'b011001 : begin
        _zz_2843_ = int_reg_array_45_25_imag;
        _zz_2844_ = int_reg_array_45_25_real;
      end
      6'b011010 : begin
        _zz_2843_ = int_reg_array_45_26_imag;
        _zz_2844_ = int_reg_array_45_26_real;
      end
      6'b011011 : begin
        _zz_2843_ = int_reg_array_45_27_imag;
        _zz_2844_ = int_reg_array_45_27_real;
      end
      6'b011100 : begin
        _zz_2843_ = int_reg_array_45_28_imag;
        _zz_2844_ = int_reg_array_45_28_real;
      end
      6'b011101 : begin
        _zz_2843_ = int_reg_array_45_29_imag;
        _zz_2844_ = int_reg_array_45_29_real;
      end
      6'b011110 : begin
        _zz_2843_ = int_reg_array_45_30_imag;
        _zz_2844_ = int_reg_array_45_30_real;
      end
      6'b011111 : begin
        _zz_2843_ = int_reg_array_45_31_imag;
        _zz_2844_ = int_reg_array_45_31_real;
      end
      6'b100000 : begin
        _zz_2843_ = int_reg_array_45_32_imag;
        _zz_2844_ = int_reg_array_45_32_real;
      end
      6'b100001 : begin
        _zz_2843_ = int_reg_array_45_33_imag;
        _zz_2844_ = int_reg_array_45_33_real;
      end
      6'b100010 : begin
        _zz_2843_ = int_reg_array_45_34_imag;
        _zz_2844_ = int_reg_array_45_34_real;
      end
      6'b100011 : begin
        _zz_2843_ = int_reg_array_45_35_imag;
        _zz_2844_ = int_reg_array_45_35_real;
      end
      6'b100100 : begin
        _zz_2843_ = int_reg_array_45_36_imag;
        _zz_2844_ = int_reg_array_45_36_real;
      end
      6'b100101 : begin
        _zz_2843_ = int_reg_array_45_37_imag;
        _zz_2844_ = int_reg_array_45_37_real;
      end
      6'b100110 : begin
        _zz_2843_ = int_reg_array_45_38_imag;
        _zz_2844_ = int_reg_array_45_38_real;
      end
      6'b100111 : begin
        _zz_2843_ = int_reg_array_45_39_imag;
        _zz_2844_ = int_reg_array_45_39_real;
      end
      6'b101000 : begin
        _zz_2843_ = int_reg_array_45_40_imag;
        _zz_2844_ = int_reg_array_45_40_real;
      end
      6'b101001 : begin
        _zz_2843_ = int_reg_array_45_41_imag;
        _zz_2844_ = int_reg_array_45_41_real;
      end
      6'b101010 : begin
        _zz_2843_ = int_reg_array_45_42_imag;
        _zz_2844_ = int_reg_array_45_42_real;
      end
      6'b101011 : begin
        _zz_2843_ = int_reg_array_45_43_imag;
        _zz_2844_ = int_reg_array_45_43_real;
      end
      6'b101100 : begin
        _zz_2843_ = int_reg_array_45_44_imag;
        _zz_2844_ = int_reg_array_45_44_real;
      end
      6'b101101 : begin
        _zz_2843_ = int_reg_array_45_45_imag;
        _zz_2844_ = int_reg_array_45_45_real;
      end
      6'b101110 : begin
        _zz_2843_ = int_reg_array_45_46_imag;
        _zz_2844_ = int_reg_array_45_46_real;
      end
      6'b101111 : begin
        _zz_2843_ = int_reg_array_45_47_imag;
        _zz_2844_ = int_reg_array_45_47_real;
      end
      6'b110000 : begin
        _zz_2843_ = int_reg_array_45_48_imag;
        _zz_2844_ = int_reg_array_45_48_real;
      end
      default : begin
        _zz_2843_ = int_reg_array_45_49_imag;
        _zz_2844_ = int_reg_array_45_49_real;
      end
    endcase
  end

  always @(*) begin
    case(_zz_2532_)
      6'b000000 : begin
        _zz_2845_ = int_reg_array_46_0_imag;
        _zz_2846_ = int_reg_array_46_0_real;
      end
      6'b000001 : begin
        _zz_2845_ = int_reg_array_46_1_imag;
        _zz_2846_ = int_reg_array_46_1_real;
      end
      6'b000010 : begin
        _zz_2845_ = int_reg_array_46_2_imag;
        _zz_2846_ = int_reg_array_46_2_real;
      end
      6'b000011 : begin
        _zz_2845_ = int_reg_array_46_3_imag;
        _zz_2846_ = int_reg_array_46_3_real;
      end
      6'b000100 : begin
        _zz_2845_ = int_reg_array_46_4_imag;
        _zz_2846_ = int_reg_array_46_4_real;
      end
      6'b000101 : begin
        _zz_2845_ = int_reg_array_46_5_imag;
        _zz_2846_ = int_reg_array_46_5_real;
      end
      6'b000110 : begin
        _zz_2845_ = int_reg_array_46_6_imag;
        _zz_2846_ = int_reg_array_46_6_real;
      end
      6'b000111 : begin
        _zz_2845_ = int_reg_array_46_7_imag;
        _zz_2846_ = int_reg_array_46_7_real;
      end
      6'b001000 : begin
        _zz_2845_ = int_reg_array_46_8_imag;
        _zz_2846_ = int_reg_array_46_8_real;
      end
      6'b001001 : begin
        _zz_2845_ = int_reg_array_46_9_imag;
        _zz_2846_ = int_reg_array_46_9_real;
      end
      6'b001010 : begin
        _zz_2845_ = int_reg_array_46_10_imag;
        _zz_2846_ = int_reg_array_46_10_real;
      end
      6'b001011 : begin
        _zz_2845_ = int_reg_array_46_11_imag;
        _zz_2846_ = int_reg_array_46_11_real;
      end
      6'b001100 : begin
        _zz_2845_ = int_reg_array_46_12_imag;
        _zz_2846_ = int_reg_array_46_12_real;
      end
      6'b001101 : begin
        _zz_2845_ = int_reg_array_46_13_imag;
        _zz_2846_ = int_reg_array_46_13_real;
      end
      6'b001110 : begin
        _zz_2845_ = int_reg_array_46_14_imag;
        _zz_2846_ = int_reg_array_46_14_real;
      end
      6'b001111 : begin
        _zz_2845_ = int_reg_array_46_15_imag;
        _zz_2846_ = int_reg_array_46_15_real;
      end
      6'b010000 : begin
        _zz_2845_ = int_reg_array_46_16_imag;
        _zz_2846_ = int_reg_array_46_16_real;
      end
      6'b010001 : begin
        _zz_2845_ = int_reg_array_46_17_imag;
        _zz_2846_ = int_reg_array_46_17_real;
      end
      6'b010010 : begin
        _zz_2845_ = int_reg_array_46_18_imag;
        _zz_2846_ = int_reg_array_46_18_real;
      end
      6'b010011 : begin
        _zz_2845_ = int_reg_array_46_19_imag;
        _zz_2846_ = int_reg_array_46_19_real;
      end
      6'b010100 : begin
        _zz_2845_ = int_reg_array_46_20_imag;
        _zz_2846_ = int_reg_array_46_20_real;
      end
      6'b010101 : begin
        _zz_2845_ = int_reg_array_46_21_imag;
        _zz_2846_ = int_reg_array_46_21_real;
      end
      6'b010110 : begin
        _zz_2845_ = int_reg_array_46_22_imag;
        _zz_2846_ = int_reg_array_46_22_real;
      end
      6'b010111 : begin
        _zz_2845_ = int_reg_array_46_23_imag;
        _zz_2846_ = int_reg_array_46_23_real;
      end
      6'b011000 : begin
        _zz_2845_ = int_reg_array_46_24_imag;
        _zz_2846_ = int_reg_array_46_24_real;
      end
      6'b011001 : begin
        _zz_2845_ = int_reg_array_46_25_imag;
        _zz_2846_ = int_reg_array_46_25_real;
      end
      6'b011010 : begin
        _zz_2845_ = int_reg_array_46_26_imag;
        _zz_2846_ = int_reg_array_46_26_real;
      end
      6'b011011 : begin
        _zz_2845_ = int_reg_array_46_27_imag;
        _zz_2846_ = int_reg_array_46_27_real;
      end
      6'b011100 : begin
        _zz_2845_ = int_reg_array_46_28_imag;
        _zz_2846_ = int_reg_array_46_28_real;
      end
      6'b011101 : begin
        _zz_2845_ = int_reg_array_46_29_imag;
        _zz_2846_ = int_reg_array_46_29_real;
      end
      6'b011110 : begin
        _zz_2845_ = int_reg_array_46_30_imag;
        _zz_2846_ = int_reg_array_46_30_real;
      end
      6'b011111 : begin
        _zz_2845_ = int_reg_array_46_31_imag;
        _zz_2846_ = int_reg_array_46_31_real;
      end
      6'b100000 : begin
        _zz_2845_ = int_reg_array_46_32_imag;
        _zz_2846_ = int_reg_array_46_32_real;
      end
      6'b100001 : begin
        _zz_2845_ = int_reg_array_46_33_imag;
        _zz_2846_ = int_reg_array_46_33_real;
      end
      6'b100010 : begin
        _zz_2845_ = int_reg_array_46_34_imag;
        _zz_2846_ = int_reg_array_46_34_real;
      end
      6'b100011 : begin
        _zz_2845_ = int_reg_array_46_35_imag;
        _zz_2846_ = int_reg_array_46_35_real;
      end
      6'b100100 : begin
        _zz_2845_ = int_reg_array_46_36_imag;
        _zz_2846_ = int_reg_array_46_36_real;
      end
      6'b100101 : begin
        _zz_2845_ = int_reg_array_46_37_imag;
        _zz_2846_ = int_reg_array_46_37_real;
      end
      6'b100110 : begin
        _zz_2845_ = int_reg_array_46_38_imag;
        _zz_2846_ = int_reg_array_46_38_real;
      end
      6'b100111 : begin
        _zz_2845_ = int_reg_array_46_39_imag;
        _zz_2846_ = int_reg_array_46_39_real;
      end
      6'b101000 : begin
        _zz_2845_ = int_reg_array_46_40_imag;
        _zz_2846_ = int_reg_array_46_40_real;
      end
      6'b101001 : begin
        _zz_2845_ = int_reg_array_46_41_imag;
        _zz_2846_ = int_reg_array_46_41_real;
      end
      6'b101010 : begin
        _zz_2845_ = int_reg_array_46_42_imag;
        _zz_2846_ = int_reg_array_46_42_real;
      end
      6'b101011 : begin
        _zz_2845_ = int_reg_array_46_43_imag;
        _zz_2846_ = int_reg_array_46_43_real;
      end
      6'b101100 : begin
        _zz_2845_ = int_reg_array_46_44_imag;
        _zz_2846_ = int_reg_array_46_44_real;
      end
      6'b101101 : begin
        _zz_2845_ = int_reg_array_46_45_imag;
        _zz_2846_ = int_reg_array_46_45_real;
      end
      6'b101110 : begin
        _zz_2845_ = int_reg_array_46_46_imag;
        _zz_2846_ = int_reg_array_46_46_real;
      end
      6'b101111 : begin
        _zz_2845_ = int_reg_array_46_47_imag;
        _zz_2846_ = int_reg_array_46_47_real;
      end
      6'b110000 : begin
        _zz_2845_ = int_reg_array_46_48_imag;
        _zz_2846_ = int_reg_array_46_48_real;
      end
      default : begin
        _zz_2845_ = int_reg_array_46_49_imag;
        _zz_2846_ = int_reg_array_46_49_real;
      end
    endcase
  end

  always @(*) begin
    case(_zz_2587_)
      6'b000000 : begin
        _zz_2847_ = int_reg_array_47_0_imag;
        _zz_2848_ = int_reg_array_47_0_real;
      end
      6'b000001 : begin
        _zz_2847_ = int_reg_array_47_1_imag;
        _zz_2848_ = int_reg_array_47_1_real;
      end
      6'b000010 : begin
        _zz_2847_ = int_reg_array_47_2_imag;
        _zz_2848_ = int_reg_array_47_2_real;
      end
      6'b000011 : begin
        _zz_2847_ = int_reg_array_47_3_imag;
        _zz_2848_ = int_reg_array_47_3_real;
      end
      6'b000100 : begin
        _zz_2847_ = int_reg_array_47_4_imag;
        _zz_2848_ = int_reg_array_47_4_real;
      end
      6'b000101 : begin
        _zz_2847_ = int_reg_array_47_5_imag;
        _zz_2848_ = int_reg_array_47_5_real;
      end
      6'b000110 : begin
        _zz_2847_ = int_reg_array_47_6_imag;
        _zz_2848_ = int_reg_array_47_6_real;
      end
      6'b000111 : begin
        _zz_2847_ = int_reg_array_47_7_imag;
        _zz_2848_ = int_reg_array_47_7_real;
      end
      6'b001000 : begin
        _zz_2847_ = int_reg_array_47_8_imag;
        _zz_2848_ = int_reg_array_47_8_real;
      end
      6'b001001 : begin
        _zz_2847_ = int_reg_array_47_9_imag;
        _zz_2848_ = int_reg_array_47_9_real;
      end
      6'b001010 : begin
        _zz_2847_ = int_reg_array_47_10_imag;
        _zz_2848_ = int_reg_array_47_10_real;
      end
      6'b001011 : begin
        _zz_2847_ = int_reg_array_47_11_imag;
        _zz_2848_ = int_reg_array_47_11_real;
      end
      6'b001100 : begin
        _zz_2847_ = int_reg_array_47_12_imag;
        _zz_2848_ = int_reg_array_47_12_real;
      end
      6'b001101 : begin
        _zz_2847_ = int_reg_array_47_13_imag;
        _zz_2848_ = int_reg_array_47_13_real;
      end
      6'b001110 : begin
        _zz_2847_ = int_reg_array_47_14_imag;
        _zz_2848_ = int_reg_array_47_14_real;
      end
      6'b001111 : begin
        _zz_2847_ = int_reg_array_47_15_imag;
        _zz_2848_ = int_reg_array_47_15_real;
      end
      6'b010000 : begin
        _zz_2847_ = int_reg_array_47_16_imag;
        _zz_2848_ = int_reg_array_47_16_real;
      end
      6'b010001 : begin
        _zz_2847_ = int_reg_array_47_17_imag;
        _zz_2848_ = int_reg_array_47_17_real;
      end
      6'b010010 : begin
        _zz_2847_ = int_reg_array_47_18_imag;
        _zz_2848_ = int_reg_array_47_18_real;
      end
      6'b010011 : begin
        _zz_2847_ = int_reg_array_47_19_imag;
        _zz_2848_ = int_reg_array_47_19_real;
      end
      6'b010100 : begin
        _zz_2847_ = int_reg_array_47_20_imag;
        _zz_2848_ = int_reg_array_47_20_real;
      end
      6'b010101 : begin
        _zz_2847_ = int_reg_array_47_21_imag;
        _zz_2848_ = int_reg_array_47_21_real;
      end
      6'b010110 : begin
        _zz_2847_ = int_reg_array_47_22_imag;
        _zz_2848_ = int_reg_array_47_22_real;
      end
      6'b010111 : begin
        _zz_2847_ = int_reg_array_47_23_imag;
        _zz_2848_ = int_reg_array_47_23_real;
      end
      6'b011000 : begin
        _zz_2847_ = int_reg_array_47_24_imag;
        _zz_2848_ = int_reg_array_47_24_real;
      end
      6'b011001 : begin
        _zz_2847_ = int_reg_array_47_25_imag;
        _zz_2848_ = int_reg_array_47_25_real;
      end
      6'b011010 : begin
        _zz_2847_ = int_reg_array_47_26_imag;
        _zz_2848_ = int_reg_array_47_26_real;
      end
      6'b011011 : begin
        _zz_2847_ = int_reg_array_47_27_imag;
        _zz_2848_ = int_reg_array_47_27_real;
      end
      6'b011100 : begin
        _zz_2847_ = int_reg_array_47_28_imag;
        _zz_2848_ = int_reg_array_47_28_real;
      end
      6'b011101 : begin
        _zz_2847_ = int_reg_array_47_29_imag;
        _zz_2848_ = int_reg_array_47_29_real;
      end
      6'b011110 : begin
        _zz_2847_ = int_reg_array_47_30_imag;
        _zz_2848_ = int_reg_array_47_30_real;
      end
      6'b011111 : begin
        _zz_2847_ = int_reg_array_47_31_imag;
        _zz_2848_ = int_reg_array_47_31_real;
      end
      6'b100000 : begin
        _zz_2847_ = int_reg_array_47_32_imag;
        _zz_2848_ = int_reg_array_47_32_real;
      end
      6'b100001 : begin
        _zz_2847_ = int_reg_array_47_33_imag;
        _zz_2848_ = int_reg_array_47_33_real;
      end
      6'b100010 : begin
        _zz_2847_ = int_reg_array_47_34_imag;
        _zz_2848_ = int_reg_array_47_34_real;
      end
      6'b100011 : begin
        _zz_2847_ = int_reg_array_47_35_imag;
        _zz_2848_ = int_reg_array_47_35_real;
      end
      6'b100100 : begin
        _zz_2847_ = int_reg_array_47_36_imag;
        _zz_2848_ = int_reg_array_47_36_real;
      end
      6'b100101 : begin
        _zz_2847_ = int_reg_array_47_37_imag;
        _zz_2848_ = int_reg_array_47_37_real;
      end
      6'b100110 : begin
        _zz_2847_ = int_reg_array_47_38_imag;
        _zz_2848_ = int_reg_array_47_38_real;
      end
      6'b100111 : begin
        _zz_2847_ = int_reg_array_47_39_imag;
        _zz_2848_ = int_reg_array_47_39_real;
      end
      6'b101000 : begin
        _zz_2847_ = int_reg_array_47_40_imag;
        _zz_2848_ = int_reg_array_47_40_real;
      end
      6'b101001 : begin
        _zz_2847_ = int_reg_array_47_41_imag;
        _zz_2848_ = int_reg_array_47_41_real;
      end
      6'b101010 : begin
        _zz_2847_ = int_reg_array_47_42_imag;
        _zz_2848_ = int_reg_array_47_42_real;
      end
      6'b101011 : begin
        _zz_2847_ = int_reg_array_47_43_imag;
        _zz_2848_ = int_reg_array_47_43_real;
      end
      6'b101100 : begin
        _zz_2847_ = int_reg_array_47_44_imag;
        _zz_2848_ = int_reg_array_47_44_real;
      end
      6'b101101 : begin
        _zz_2847_ = int_reg_array_47_45_imag;
        _zz_2848_ = int_reg_array_47_45_real;
      end
      6'b101110 : begin
        _zz_2847_ = int_reg_array_47_46_imag;
        _zz_2848_ = int_reg_array_47_46_real;
      end
      6'b101111 : begin
        _zz_2847_ = int_reg_array_47_47_imag;
        _zz_2848_ = int_reg_array_47_47_real;
      end
      6'b110000 : begin
        _zz_2847_ = int_reg_array_47_48_imag;
        _zz_2848_ = int_reg_array_47_48_real;
      end
      default : begin
        _zz_2847_ = int_reg_array_47_49_imag;
        _zz_2848_ = int_reg_array_47_49_real;
      end
    endcase
  end

  always @(*) begin
    case(_zz_2642_)
      6'b000000 : begin
        _zz_2849_ = int_reg_array_48_0_imag;
        _zz_2850_ = int_reg_array_48_0_real;
      end
      6'b000001 : begin
        _zz_2849_ = int_reg_array_48_1_imag;
        _zz_2850_ = int_reg_array_48_1_real;
      end
      6'b000010 : begin
        _zz_2849_ = int_reg_array_48_2_imag;
        _zz_2850_ = int_reg_array_48_2_real;
      end
      6'b000011 : begin
        _zz_2849_ = int_reg_array_48_3_imag;
        _zz_2850_ = int_reg_array_48_3_real;
      end
      6'b000100 : begin
        _zz_2849_ = int_reg_array_48_4_imag;
        _zz_2850_ = int_reg_array_48_4_real;
      end
      6'b000101 : begin
        _zz_2849_ = int_reg_array_48_5_imag;
        _zz_2850_ = int_reg_array_48_5_real;
      end
      6'b000110 : begin
        _zz_2849_ = int_reg_array_48_6_imag;
        _zz_2850_ = int_reg_array_48_6_real;
      end
      6'b000111 : begin
        _zz_2849_ = int_reg_array_48_7_imag;
        _zz_2850_ = int_reg_array_48_7_real;
      end
      6'b001000 : begin
        _zz_2849_ = int_reg_array_48_8_imag;
        _zz_2850_ = int_reg_array_48_8_real;
      end
      6'b001001 : begin
        _zz_2849_ = int_reg_array_48_9_imag;
        _zz_2850_ = int_reg_array_48_9_real;
      end
      6'b001010 : begin
        _zz_2849_ = int_reg_array_48_10_imag;
        _zz_2850_ = int_reg_array_48_10_real;
      end
      6'b001011 : begin
        _zz_2849_ = int_reg_array_48_11_imag;
        _zz_2850_ = int_reg_array_48_11_real;
      end
      6'b001100 : begin
        _zz_2849_ = int_reg_array_48_12_imag;
        _zz_2850_ = int_reg_array_48_12_real;
      end
      6'b001101 : begin
        _zz_2849_ = int_reg_array_48_13_imag;
        _zz_2850_ = int_reg_array_48_13_real;
      end
      6'b001110 : begin
        _zz_2849_ = int_reg_array_48_14_imag;
        _zz_2850_ = int_reg_array_48_14_real;
      end
      6'b001111 : begin
        _zz_2849_ = int_reg_array_48_15_imag;
        _zz_2850_ = int_reg_array_48_15_real;
      end
      6'b010000 : begin
        _zz_2849_ = int_reg_array_48_16_imag;
        _zz_2850_ = int_reg_array_48_16_real;
      end
      6'b010001 : begin
        _zz_2849_ = int_reg_array_48_17_imag;
        _zz_2850_ = int_reg_array_48_17_real;
      end
      6'b010010 : begin
        _zz_2849_ = int_reg_array_48_18_imag;
        _zz_2850_ = int_reg_array_48_18_real;
      end
      6'b010011 : begin
        _zz_2849_ = int_reg_array_48_19_imag;
        _zz_2850_ = int_reg_array_48_19_real;
      end
      6'b010100 : begin
        _zz_2849_ = int_reg_array_48_20_imag;
        _zz_2850_ = int_reg_array_48_20_real;
      end
      6'b010101 : begin
        _zz_2849_ = int_reg_array_48_21_imag;
        _zz_2850_ = int_reg_array_48_21_real;
      end
      6'b010110 : begin
        _zz_2849_ = int_reg_array_48_22_imag;
        _zz_2850_ = int_reg_array_48_22_real;
      end
      6'b010111 : begin
        _zz_2849_ = int_reg_array_48_23_imag;
        _zz_2850_ = int_reg_array_48_23_real;
      end
      6'b011000 : begin
        _zz_2849_ = int_reg_array_48_24_imag;
        _zz_2850_ = int_reg_array_48_24_real;
      end
      6'b011001 : begin
        _zz_2849_ = int_reg_array_48_25_imag;
        _zz_2850_ = int_reg_array_48_25_real;
      end
      6'b011010 : begin
        _zz_2849_ = int_reg_array_48_26_imag;
        _zz_2850_ = int_reg_array_48_26_real;
      end
      6'b011011 : begin
        _zz_2849_ = int_reg_array_48_27_imag;
        _zz_2850_ = int_reg_array_48_27_real;
      end
      6'b011100 : begin
        _zz_2849_ = int_reg_array_48_28_imag;
        _zz_2850_ = int_reg_array_48_28_real;
      end
      6'b011101 : begin
        _zz_2849_ = int_reg_array_48_29_imag;
        _zz_2850_ = int_reg_array_48_29_real;
      end
      6'b011110 : begin
        _zz_2849_ = int_reg_array_48_30_imag;
        _zz_2850_ = int_reg_array_48_30_real;
      end
      6'b011111 : begin
        _zz_2849_ = int_reg_array_48_31_imag;
        _zz_2850_ = int_reg_array_48_31_real;
      end
      6'b100000 : begin
        _zz_2849_ = int_reg_array_48_32_imag;
        _zz_2850_ = int_reg_array_48_32_real;
      end
      6'b100001 : begin
        _zz_2849_ = int_reg_array_48_33_imag;
        _zz_2850_ = int_reg_array_48_33_real;
      end
      6'b100010 : begin
        _zz_2849_ = int_reg_array_48_34_imag;
        _zz_2850_ = int_reg_array_48_34_real;
      end
      6'b100011 : begin
        _zz_2849_ = int_reg_array_48_35_imag;
        _zz_2850_ = int_reg_array_48_35_real;
      end
      6'b100100 : begin
        _zz_2849_ = int_reg_array_48_36_imag;
        _zz_2850_ = int_reg_array_48_36_real;
      end
      6'b100101 : begin
        _zz_2849_ = int_reg_array_48_37_imag;
        _zz_2850_ = int_reg_array_48_37_real;
      end
      6'b100110 : begin
        _zz_2849_ = int_reg_array_48_38_imag;
        _zz_2850_ = int_reg_array_48_38_real;
      end
      6'b100111 : begin
        _zz_2849_ = int_reg_array_48_39_imag;
        _zz_2850_ = int_reg_array_48_39_real;
      end
      6'b101000 : begin
        _zz_2849_ = int_reg_array_48_40_imag;
        _zz_2850_ = int_reg_array_48_40_real;
      end
      6'b101001 : begin
        _zz_2849_ = int_reg_array_48_41_imag;
        _zz_2850_ = int_reg_array_48_41_real;
      end
      6'b101010 : begin
        _zz_2849_ = int_reg_array_48_42_imag;
        _zz_2850_ = int_reg_array_48_42_real;
      end
      6'b101011 : begin
        _zz_2849_ = int_reg_array_48_43_imag;
        _zz_2850_ = int_reg_array_48_43_real;
      end
      6'b101100 : begin
        _zz_2849_ = int_reg_array_48_44_imag;
        _zz_2850_ = int_reg_array_48_44_real;
      end
      6'b101101 : begin
        _zz_2849_ = int_reg_array_48_45_imag;
        _zz_2850_ = int_reg_array_48_45_real;
      end
      6'b101110 : begin
        _zz_2849_ = int_reg_array_48_46_imag;
        _zz_2850_ = int_reg_array_48_46_real;
      end
      6'b101111 : begin
        _zz_2849_ = int_reg_array_48_47_imag;
        _zz_2850_ = int_reg_array_48_47_real;
      end
      6'b110000 : begin
        _zz_2849_ = int_reg_array_48_48_imag;
        _zz_2850_ = int_reg_array_48_48_real;
      end
      default : begin
        _zz_2849_ = int_reg_array_48_49_imag;
        _zz_2850_ = int_reg_array_48_49_real;
      end
    endcase
  end

  always @(*) begin
    case(_zz_2697_)
      6'b000000 : begin
        _zz_2851_ = int_reg_array_49_0_imag;
        _zz_2852_ = int_reg_array_49_0_real;
      end
      6'b000001 : begin
        _zz_2851_ = int_reg_array_49_1_imag;
        _zz_2852_ = int_reg_array_49_1_real;
      end
      6'b000010 : begin
        _zz_2851_ = int_reg_array_49_2_imag;
        _zz_2852_ = int_reg_array_49_2_real;
      end
      6'b000011 : begin
        _zz_2851_ = int_reg_array_49_3_imag;
        _zz_2852_ = int_reg_array_49_3_real;
      end
      6'b000100 : begin
        _zz_2851_ = int_reg_array_49_4_imag;
        _zz_2852_ = int_reg_array_49_4_real;
      end
      6'b000101 : begin
        _zz_2851_ = int_reg_array_49_5_imag;
        _zz_2852_ = int_reg_array_49_5_real;
      end
      6'b000110 : begin
        _zz_2851_ = int_reg_array_49_6_imag;
        _zz_2852_ = int_reg_array_49_6_real;
      end
      6'b000111 : begin
        _zz_2851_ = int_reg_array_49_7_imag;
        _zz_2852_ = int_reg_array_49_7_real;
      end
      6'b001000 : begin
        _zz_2851_ = int_reg_array_49_8_imag;
        _zz_2852_ = int_reg_array_49_8_real;
      end
      6'b001001 : begin
        _zz_2851_ = int_reg_array_49_9_imag;
        _zz_2852_ = int_reg_array_49_9_real;
      end
      6'b001010 : begin
        _zz_2851_ = int_reg_array_49_10_imag;
        _zz_2852_ = int_reg_array_49_10_real;
      end
      6'b001011 : begin
        _zz_2851_ = int_reg_array_49_11_imag;
        _zz_2852_ = int_reg_array_49_11_real;
      end
      6'b001100 : begin
        _zz_2851_ = int_reg_array_49_12_imag;
        _zz_2852_ = int_reg_array_49_12_real;
      end
      6'b001101 : begin
        _zz_2851_ = int_reg_array_49_13_imag;
        _zz_2852_ = int_reg_array_49_13_real;
      end
      6'b001110 : begin
        _zz_2851_ = int_reg_array_49_14_imag;
        _zz_2852_ = int_reg_array_49_14_real;
      end
      6'b001111 : begin
        _zz_2851_ = int_reg_array_49_15_imag;
        _zz_2852_ = int_reg_array_49_15_real;
      end
      6'b010000 : begin
        _zz_2851_ = int_reg_array_49_16_imag;
        _zz_2852_ = int_reg_array_49_16_real;
      end
      6'b010001 : begin
        _zz_2851_ = int_reg_array_49_17_imag;
        _zz_2852_ = int_reg_array_49_17_real;
      end
      6'b010010 : begin
        _zz_2851_ = int_reg_array_49_18_imag;
        _zz_2852_ = int_reg_array_49_18_real;
      end
      6'b010011 : begin
        _zz_2851_ = int_reg_array_49_19_imag;
        _zz_2852_ = int_reg_array_49_19_real;
      end
      6'b010100 : begin
        _zz_2851_ = int_reg_array_49_20_imag;
        _zz_2852_ = int_reg_array_49_20_real;
      end
      6'b010101 : begin
        _zz_2851_ = int_reg_array_49_21_imag;
        _zz_2852_ = int_reg_array_49_21_real;
      end
      6'b010110 : begin
        _zz_2851_ = int_reg_array_49_22_imag;
        _zz_2852_ = int_reg_array_49_22_real;
      end
      6'b010111 : begin
        _zz_2851_ = int_reg_array_49_23_imag;
        _zz_2852_ = int_reg_array_49_23_real;
      end
      6'b011000 : begin
        _zz_2851_ = int_reg_array_49_24_imag;
        _zz_2852_ = int_reg_array_49_24_real;
      end
      6'b011001 : begin
        _zz_2851_ = int_reg_array_49_25_imag;
        _zz_2852_ = int_reg_array_49_25_real;
      end
      6'b011010 : begin
        _zz_2851_ = int_reg_array_49_26_imag;
        _zz_2852_ = int_reg_array_49_26_real;
      end
      6'b011011 : begin
        _zz_2851_ = int_reg_array_49_27_imag;
        _zz_2852_ = int_reg_array_49_27_real;
      end
      6'b011100 : begin
        _zz_2851_ = int_reg_array_49_28_imag;
        _zz_2852_ = int_reg_array_49_28_real;
      end
      6'b011101 : begin
        _zz_2851_ = int_reg_array_49_29_imag;
        _zz_2852_ = int_reg_array_49_29_real;
      end
      6'b011110 : begin
        _zz_2851_ = int_reg_array_49_30_imag;
        _zz_2852_ = int_reg_array_49_30_real;
      end
      6'b011111 : begin
        _zz_2851_ = int_reg_array_49_31_imag;
        _zz_2852_ = int_reg_array_49_31_real;
      end
      6'b100000 : begin
        _zz_2851_ = int_reg_array_49_32_imag;
        _zz_2852_ = int_reg_array_49_32_real;
      end
      6'b100001 : begin
        _zz_2851_ = int_reg_array_49_33_imag;
        _zz_2852_ = int_reg_array_49_33_real;
      end
      6'b100010 : begin
        _zz_2851_ = int_reg_array_49_34_imag;
        _zz_2852_ = int_reg_array_49_34_real;
      end
      6'b100011 : begin
        _zz_2851_ = int_reg_array_49_35_imag;
        _zz_2852_ = int_reg_array_49_35_real;
      end
      6'b100100 : begin
        _zz_2851_ = int_reg_array_49_36_imag;
        _zz_2852_ = int_reg_array_49_36_real;
      end
      6'b100101 : begin
        _zz_2851_ = int_reg_array_49_37_imag;
        _zz_2852_ = int_reg_array_49_37_real;
      end
      6'b100110 : begin
        _zz_2851_ = int_reg_array_49_38_imag;
        _zz_2852_ = int_reg_array_49_38_real;
      end
      6'b100111 : begin
        _zz_2851_ = int_reg_array_49_39_imag;
        _zz_2852_ = int_reg_array_49_39_real;
      end
      6'b101000 : begin
        _zz_2851_ = int_reg_array_49_40_imag;
        _zz_2852_ = int_reg_array_49_40_real;
      end
      6'b101001 : begin
        _zz_2851_ = int_reg_array_49_41_imag;
        _zz_2852_ = int_reg_array_49_41_real;
      end
      6'b101010 : begin
        _zz_2851_ = int_reg_array_49_42_imag;
        _zz_2852_ = int_reg_array_49_42_real;
      end
      6'b101011 : begin
        _zz_2851_ = int_reg_array_49_43_imag;
        _zz_2852_ = int_reg_array_49_43_real;
      end
      6'b101100 : begin
        _zz_2851_ = int_reg_array_49_44_imag;
        _zz_2852_ = int_reg_array_49_44_real;
      end
      6'b101101 : begin
        _zz_2851_ = int_reg_array_49_45_imag;
        _zz_2852_ = int_reg_array_49_45_real;
      end
      6'b101110 : begin
        _zz_2851_ = int_reg_array_49_46_imag;
        _zz_2852_ = int_reg_array_49_46_real;
      end
      6'b101111 : begin
        _zz_2851_ = int_reg_array_49_47_imag;
        _zz_2852_ = int_reg_array_49_47_real;
      end
      6'b110000 : begin
        _zz_2851_ = int_reg_array_49_48_imag;
        _zz_2852_ = int_reg_array_49_48_real;
      end
      default : begin
        _zz_2851_ = int_reg_array_49_49_imag;
        _zz_2852_ = int_reg_array_49_49_real;
      end
    endcase
  end

  assign axi4_b_valid = axi4_w_valid;
  assign axi4_b_payload_id = aw_area_awid_r;
  assign axi4_b_payload_resp = (2'b00);
  assign axi4_aw_ready = 1'b1;
  assign axi4_w_ready = 1'b1;
  assign Axi4Incr_highCat = aw_area_awaddr_r[31 : 12];
  assign Axi4Incr_sizeValue = 1'b1;
  assign Axi4Incr_alignMask = 12'h0;
  assign Axi4Incr_base = (_zz_2854_ & (~ Axi4Incr_alignMask));
  assign Axi4Incr_baseIncr = (Axi4Incr_base + _zz_2855_);
  always @ (*) begin
    if((((aw_area_awlen_r & 8'h08) == 8'h08))) begin
        _zz_1_ = (2'b11);
    end else if((((aw_area_awlen_r & 8'h04) == 8'h04))) begin
        _zz_1_ = (2'b10);
    end else if((((aw_area_awlen_r & 8'h02) == 8'h02))) begin
        _zz_1_ = (2'b01);
    end else begin
        _zz_1_ = (2'b00);
    end
  end

  assign Axi4Incr_wrapCase = ((2'b00) + _zz_1_);
  always @ (*) begin
    case(axi4_aw_payload_burst)
      2'b00 : begin
        Axi4Incr_result = aw_area_awaddr_r;
      end
      2'b10 : begin
        Axi4Incr_result = {Axi4Incr_highCat,_zz_2752_};
      end
      default : begin
        Axi4Incr_result = {Axi4Incr_highCat,Axi4Incr_baseIncr};
      end
    endcase
  end

  assign _zz_2_ = _zz_2857_[5:0];
  assign _zz_3_ = ({63'd0,(1'b1)} <<< _zz_2_);
  assign _zz_4_ = _zz_3_[0];
  assign _zz_5_ = _zz_3_[1];
  assign _zz_6_ = _zz_3_[2];
  assign _zz_7_ = _zz_3_[3];
  assign _zz_8_ = _zz_3_[4];
  assign _zz_9_ = _zz_3_[5];
  assign _zz_10_ = _zz_3_[6];
  assign _zz_11_ = _zz_3_[7];
  assign _zz_12_ = _zz_3_[8];
  assign _zz_13_ = _zz_3_[9];
  assign _zz_14_ = _zz_3_[10];
  assign _zz_15_ = _zz_3_[11];
  assign _zz_16_ = _zz_3_[12];
  assign _zz_17_ = _zz_3_[13];
  assign _zz_18_ = _zz_3_[14];
  assign _zz_19_ = _zz_3_[15];
  assign _zz_20_ = _zz_3_[16];
  assign _zz_21_ = _zz_3_[17];
  assign _zz_22_ = _zz_3_[18];
  assign _zz_23_ = _zz_3_[19];
  assign _zz_24_ = _zz_3_[20];
  assign _zz_25_ = _zz_3_[21];
  assign _zz_26_ = _zz_3_[22];
  assign _zz_27_ = _zz_3_[23];
  assign _zz_28_ = _zz_3_[24];
  assign _zz_29_ = _zz_3_[25];
  assign _zz_30_ = _zz_3_[26];
  assign _zz_31_ = _zz_3_[27];
  assign _zz_32_ = _zz_3_[28];
  assign _zz_33_ = _zz_3_[29];
  assign _zz_34_ = _zz_3_[30];
  assign _zz_35_ = _zz_3_[31];
  assign _zz_36_ = _zz_3_[32];
  assign _zz_37_ = _zz_3_[33];
  assign _zz_38_ = _zz_3_[34];
  assign _zz_39_ = _zz_3_[35];
  assign _zz_40_ = _zz_3_[36];
  assign _zz_41_ = _zz_3_[37];
  assign _zz_42_ = _zz_3_[38];
  assign _zz_43_ = _zz_3_[39];
  assign _zz_44_ = _zz_3_[40];
  assign _zz_45_ = _zz_3_[41];
  assign _zz_46_ = _zz_3_[42];
  assign _zz_47_ = _zz_3_[43];
  assign _zz_48_ = _zz_3_[44];
  assign _zz_49_ = _zz_3_[45];
  assign _zz_50_ = _zz_3_[46];
  assign _zz_51_ = _zz_3_[47];
  assign _zz_52_ = _zz_3_[48];
  assign _zz_53_ = _zz_3_[49];
  assign _zz_54_ = (((32'h00000064 <= load_data_area_current_addr) && (load_data_area_current_addr < 32'h00000096)) ? axi4_w_payload_data_regNext : {_zz_2753_,_zz_2754_});
  assign _zz_55_ = _zz_54_[15 : 0];
  assign _zz_56_ = _zz_54_[31 : 16];
  assign _zz_57_ = _zz_2858_[5:0];
  assign _zz_58_ = ({63'd0,(1'b1)} <<< _zz_57_);
  assign _zz_59_ = _zz_58_[0];
  assign _zz_60_ = _zz_58_[1];
  assign _zz_61_ = _zz_58_[2];
  assign _zz_62_ = _zz_58_[3];
  assign _zz_63_ = _zz_58_[4];
  assign _zz_64_ = _zz_58_[5];
  assign _zz_65_ = _zz_58_[6];
  assign _zz_66_ = _zz_58_[7];
  assign _zz_67_ = _zz_58_[8];
  assign _zz_68_ = _zz_58_[9];
  assign _zz_69_ = _zz_58_[10];
  assign _zz_70_ = _zz_58_[11];
  assign _zz_71_ = _zz_58_[12];
  assign _zz_72_ = _zz_58_[13];
  assign _zz_73_ = _zz_58_[14];
  assign _zz_74_ = _zz_58_[15];
  assign _zz_75_ = _zz_58_[16];
  assign _zz_76_ = _zz_58_[17];
  assign _zz_77_ = _zz_58_[18];
  assign _zz_78_ = _zz_58_[19];
  assign _zz_79_ = _zz_58_[20];
  assign _zz_80_ = _zz_58_[21];
  assign _zz_81_ = _zz_58_[22];
  assign _zz_82_ = _zz_58_[23];
  assign _zz_83_ = _zz_58_[24];
  assign _zz_84_ = _zz_58_[25];
  assign _zz_85_ = _zz_58_[26];
  assign _zz_86_ = _zz_58_[27];
  assign _zz_87_ = _zz_58_[28];
  assign _zz_88_ = _zz_58_[29];
  assign _zz_89_ = _zz_58_[30];
  assign _zz_90_ = _zz_58_[31];
  assign _zz_91_ = _zz_58_[32];
  assign _zz_92_ = _zz_58_[33];
  assign _zz_93_ = _zz_58_[34];
  assign _zz_94_ = _zz_58_[35];
  assign _zz_95_ = _zz_58_[36];
  assign _zz_96_ = _zz_58_[37];
  assign _zz_97_ = _zz_58_[38];
  assign _zz_98_ = _zz_58_[39];
  assign _zz_99_ = _zz_58_[40];
  assign _zz_100_ = _zz_58_[41];
  assign _zz_101_ = _zz_58_[42];
  assign _zz_102_ = _zz_58_[43];
  assign _zz_103_ = _zz_58_[44];
  assign _zz_104_ = _zz_58_[45];
  assign _zz_105_ = _zz_58_[46];
  assign _zz_106_ = _zz_58_[47];
  assign _zz_107_ = _zz_58_[48];
  assign _zz_108_ = _zz_58_[49];
  assign _zz_109_ = (((32'h0000028a <= load_data_area_current_addr) && (load_data_area_current_addr < 32'h000002bc)) ? axi4_w_payload_data_regNext : {_zz_2755_,_zz_2756_});
  assign _zz_110_ = _zz_109_[15 : 0];
  assign _zz_111_ = _zz_109_[31 : 16];
  assign _zz_112_ = _zz_2859_[5:0];
  assign _zz_113_ = ({63'd0,(1'b1)} <<< _zz_112_);
  assign _zz_114_ = _zz_113_[0];
  assign _zz_115_ = _zz_113_[1];
  assign _zz_116_ = _zz_113_[2];
  assign _zz_117_ = _zz_113_[3];
  assign _zz_118_ = _zz_113_[4];
  assign _zz_119_ = _zz_113_[5];
  assign _zz_120_ = _zz_113_[6];
  assign _zz_121_ = _zz_113_[7];
  assign _zz_122_ = _zz_113_[8];
  assign _zz_123_ = _zz_113_[9];
  assign _zz_124_ = _zz_113_[10];
  assign _zz_125_ = _zz_113_[11];
  assign _zz_126_ = _zz_113_[12];
  assign _zz_127_ = _zz_113_[13];
  assign _zz_128_ = _zz_113_[14];
  assign _zz_129_ = _zz_113_[15];
  assign _zz_130_ = _zz_113_[16];
  assign _zz_131_ = _zz_113_[17];
  assign _zz_132_ = _zz_113_[18];
  assign _zz_133_ = _zz_113_[19];
  assign _zz_134_ = _zz_113_[20];
  assign _zz_135_ = _zz_113_[21];
  assign _zz_136_ = _zz_113_[22];
  assign _zz_137_ = _zz_113_[23];
  assign _zz_138_ = _zz_113_[24];
  assign _zz_139_ = _zz_113_[25];
  assign _zz_140_ = _zz_113_[26];
  assign _zz_141_ = _zz_113_[27];
  assign _zz_142_ = _zz_113_[28];
  assign _zz_143_ = _zz_113_[29];
  assign _zz_144_ = _zz_113_[30];
  assign _zz_145_ = _zz_113_[31];
  assign _zz_146_ = _zz_113_[32];
  assign _zz_147_ = _zz_113_[33];
  assign _zz_148_ = _zz_113_[34];
  assign _zz_149_ = _zz_113_[35];
  assign _zz_150_ = _zz_113_[36];
  assign _zz_151_ = _zz_113_[37];
  assign _zz_152_ = _zz_113_[38];
  assign _zz_153_ = _zz_113_[39];
  assign _zz_154_ = _zz_113_[40];
  assign _zz_155_ = _zz_113_[41];
  assign _zz_156_ = _zz_113_[42];
  assign _zz_157_ = _zz_113_[43];
  assign _zz_158_ = _zz_113_[44];
  assign _zz_159_ = _zz_113_[45];
  assign _zz_160_ = _zz_113_[46];
  assign _zz_161_ = _zz_113_[47];
  assign _zz_162_ = _zz_113_[48];
  assign _zz_163_ = _zz_113_[49];
  assign _zz_164_ = (((32'h000002bc <= load_data_area_current_addr) && (load_data_area_current_addr < 32'h000002ee)) ? axi4_w_payload_data_regNext : {_zz_2757_,_zz_2758_});
  assign _zz_165_ = _zz_164_[15 : 0];
  assign _zz_166_ = _zz_164_[31 : 16];
  assign _zz_167_ = _zz_2860_[5:0];
  assign _zz_168_ = ({63'd0,(1'b1)} <<< _zz_167_);
  assign _zz_169_ = _zz_168_[0];
  assign _zz_170_ = _zz_168_[1];
  assign _zz_171_ = _zz_168_[2];
  assign _zz_172_ = _zz_168_[3];
  assign _zz_173_ = _zz_168_[4];
  assign _zz_174_ = _zz_168_[5];
  assign _zz_175_ = _zz_168_[6];
  assign _zz_176_ = _zz_168_[7];
  assign _zz_177_ = _zz_168_[8];
  assign _zz_178_ = _zz_168_[9];
  assign _zz_179_ = _zz_168_[10];
  assign _zz_180_ = _zz_168_[11];
  assign _zz_181_ = _zz_168_[12];
  assign _zz_182_ = _zz_168_[13];
  assign _zz_183_ = _zz_168_[14];
  assign _zz_184_ = _zz_168_[15];
  assign _zz_185_ = _zz_168_[16];
  assign _zz_186_ = _zz_168_[17];
  assign _zz_187_ = _zz_168_[18];
  assign _zz_188_ = _zz_168_[19];
  assign _zz_189_ = _zz_168_[20];
  assign _zz_190_ = _zz_168_[21];
  assign _zz_191_ = _zz_168_[22];
  assign _zz_192_ = _zz_168_[23];
  assign _zz_193_ = _zz_168_[24];
  assign _zz_194_ = _zz_168_[25];
  assign _zz_195_ = _zz_168_[26];
  assign _zz_196_ = _zz_168_[27];
  assign _zz_197_ = _zz_168_[28];
  assign _zz_198_ = _zz_168_[29];
  assign _zz_199_ = _zz_168_[30];
  assign _zz_200_ = _zz_168_[31];
  assign _zz_201_ = _zz_168_[32];
  assign _zz_202_ = _zz_168_[33];
  assign _zz_203_ = _zz_168_[34];
  assign _zz_204_ = _zz_168_[35];
  assign _zz_205_ = _zz_168_[36];
  assign _zz_206_ = _zz_168_[37];
  assign _zz_207_ = _zz_168_[38];
  assign _zz_208_ = _zz_168_[39];
  assign _zz_209_ = _zz_168_[40];
  assign _zz_210_ = _zz_168_[41];
  assign _zz_211_ = _zz_168_[42];
  assign _zz_212_ = _zz_168_[43];
  assign _zz_213_ = _zz_168_[44];
  assign _zz_214_ = _zz_168_[45];
  assign _zz_215_ = _zz_168_[46];
  assign _zz_216_ = _zz_168_[47];
  assign _zz_217_ = _zz_168_[48];
  assign _zz_218_ = _zz_168_[49];
  assign _zz_219_ = (((32'h000003b6 <= load_data_area_current_addr) && (load_data_area_current_addr < 32'h000003e8)) ? axi4_w_payload_data_regNext : {_zz_2759_,_zz_2760_});
  assign _zz_220_ = _zz_219_[15 : 0];
  assign _zz_221_ = _zz_219_[31 : 16];
  assign _zz_222_ = _zz_2861_[5:0];
  assign _zz_223_ = ({63'd0,(1'b1)} <<< _zz_222_);
  assign _zz_224_ = _zz_223_[0];
  assign _zz_225_ = _zz_223_[1];
  assign _zz_226_ = _zz_223_[2];
  assign _zz_227_ = _zz_223_[3];
  assign _zz_228_ = _zz_223_[4];
  assign _zz_229_ = _zz_223_[5];
  assign _zz_230_ = _zz_223_[6];
  assign _zz_231_ = _zz_223_[7];
  assign _zz_232_ = _zz_223_[8];
  assign _zz_233_ = _zz_223_[9];
  assign _zz_234_ = _zz_223_[10];
  assign _zz_235_ = _zz_223_[11];
  assign _zz_236_ = _zz_223_[12];
  assign _zz_237_ = _zz_223_[13];
  assign _zz_238_ = _zz_223_[14];
  assign _zz_239_ = _zz_223_[15];
  assign _zz_240_ = _zz_223_[16];
  assign _zz_241_ = _zz_223_[17];
  assign _zz_242_ = _zz_223_[18];
  assign _zz_243_ = _zz_223_[19];
  assign _zz_244_ = _zz_223_[20];
  assign _zz_245_ = _zz_223_[21];
  assign _zz_246_ = _zz_223_[22];
  assign _zz_247_ = _zz_223_[23];
  assign _zz_248_ = _zz_223_[24];
  assign _zz_249_ = _zz_223_[25];
  assign _zz_250_ = _zz_223_[26];
  assign _zz_251_ = _zz_223_[27];
  assign _zz_252_ = _zz_223_[28];
  assign _zz_253_ = _zz_223_[29];
  assign _zz_254_ = _zz_223_[30];
  assign _zz_255_ = _zz_223_[31];
  assign _zz_256_ = _zz_223_[32];
  assign _zz_257_ = _zz_223_[33];
  assign _zz_258_ = _zz_223_[34];
  assign _zz_259_ = _zz_223_[35];
  assign _zz_260_ = _zz_223_[36];
  assign _zz_261_ = _zz_223_[37];
  assign _zz_262_ = _zz_223_[38];
  assign _zz_263_ = _zz_223_[39];
  assign _zz_264_ = _zz_223_[40];
  assign _zz_265_ = _zz_223_[41];
  assign _zz_266_ = _zz_223_[42];
  assign _zz_267_ = _zz_223_[43];
  assign _zz_268_ = _zz_223_[44];
  assign _zz_269_ = _zz_223_[45];
  assign _zz_270_ = _zz_223_[46];
  assign _zz_271_ = _zz_223_[47];
  assign _zz_272_ = _zz_223_[48];
  assign _zz_273_ = _zz_223_[49];
  assign _zz_274_ = (((32'h00000672 <= load_data_area_current_addr) && (load_data_area_current_addr < 32'h000006a4)) ? axi4_w_payload_data_regNext : {_zz_2761_,_zz_2762_});
  assign _zz_275_ = _zz_274_[15 : 0];
  assign _zz_276_ = _zz_274_[31 : 16];
  assign _zz_277_ = _zz_2862_[5:0];
  assign _zz_278_ = ({63'd0,(1'b1)} <<< _zz_277_);
  assign _zz_279_ = _zz_278_[0];
  assign _zz_280_ = _zz_278_[1];
  assign _zz_281_ = _zz_278_[2];
  assign _zz_282_ = _zz_278_[3];
  assign _zz_283_ = _zz_278_[4];
  assign _zz_284_ = _zz_278_[5];
  assign _zz_285_ = _zz_278_[6];
  assign _zz_286_ = _zz_278_[7];
  assign _zz_287_ = _zz_278_[8];
  assign _zz_288_ = _zz_278_[9];
  assign _zz_289_ = _zz_278_[10];
  assign _zz_290_ = _zz_278_[11];
  assign _zz_291_ = _zz_278_[12];
  assign _zz_292_ = _zz_278_[13];
  assign _zz_293_ = _zz_278_[14];
  assign _zz_294_ = _zz_278_[15];
  assign _zz_295_ = _zz_278_[16];
  assign _zz_296_ = _zz_278_[17];
  assign _zz_297_ = _zz_278_[18];
  assign _zz_298_ = _zz_278_[19];
  assign _zz_299_ = _zz_278_[20];
  assign _zz_300_ = _zz_278_[21];
  assign _zz_301_ = _zz_278_[22];
  assign _zz_302_ = _zz_278_[23];
  assign _zz_303_ = _zz_278_[24];
  assign _zz_304_ = _zz_278_[25];
  assign _zz_305_ = _zz_278_[26];
  assign _zz_306_ = _zz_278_[27];
  assign _zz_307_ = _zz_278_[28];
  assign _zz_308_ = _zz_278_[29];
  assign _zz_309_ = _zz_278_[30];
  assign _zz_310_ = _zz_278_[31];
  assign _zz_311_ = _zz_278_[32];
  assign _zz_312_ = _zz_278_[33];
  assign _zz_313_ = _zz_278_[34];
  assign _zz_314_ = _zz_278_[35];
  assign _zz_315_ = _zz_278_[36];
  assign _zz_316_ = _zz_278_[37];
  assign _zz_317_ = _zz_278_[38];
  assign _zz_318_ = _zz_278_[39];
  assign _zz_319_ = _zz_278_[40];
  assign _zz_320_ = _zz_278_[41];
  assign _zz_321_ = _zz_278_[42];
  assign _zz_322_ = _zz_278_[43];
  assign _zz_323_ = _zz_278_[44];
  assign _zz_324_ = _zz_278_[45];
  assign _zz_325_ = _zz_278_[46];
  assign _zz_326_ = _zz_278_[47];
  assign _zz_327_ = _zz_278_[48];
  assign _zz_328_ = _zz_278_[49];
  assign _zz_329_ = (((32'h00000352 <= load_data_area_current_addr) && (load_data_area_current_addr < 32'h00000384)) ? axi4_w_payload_data_regNext : {_zz_2763_,_zz_2764_});
  assign _zz_330_ = _zz_329_[15 : 0];
  assign _zz_331_ = _zz_329_[31 : 16];
  assign _zz_332_ = _zz_2863_[5:0];
  assign _zz_333_ = ({63'd0,(1'b1)} <<< _zz_332_);
  assign _zz_334_ = _zz_333_[0];
  assign _zz_335_ = _zz_333_[1];
  assign _zz_336_ = _zz_333_[2];
  assign _zz_337_ = _zz_333_[3];
  assign _zz_338_ = _zz_333_[4];
  assign _zz_339_ = _zz_333_[5];
  assign _zz_340_ = _zz_333_[6];
  assign _zz_341_ = _zz_333_[7];
  assign _zz_342_ = _zz_333_[8];
  assign _zz_343_ = _zz_333_[9];
  assign _zz_344_ = _zz_333_[10];
  assign _zz_345_ = _zz_333_[11];
  assign _zz_346_ = _zz_333_[12];
  assign _zz_347_ = _zz_333_[13];
  assign _zz_348_ = _zz_333_[14];
  assign _zz_349_ = _zz_333_[15];
  assign _zz_350_ = _zz_333_[16];
  assign _zz_351_ = _zz_333_[17];
  assign _zz_352_ = _zz_333_[18];
  assign _zz_353_ = _zz_333_[19];
  assign _zz_354_ = _zz_333_[20];
  assign _zz_355_ = _zz_333_[21];
  assign _zz_356_ = _zz_333_[22];
  assign _zz_357_ = _zz_333_[23];
  assign _zz_358_ = _zz_333_[24];
  assign _zz_359_ = _zz_333_[25];
  assign _zz_360_ = _zz_333_[26];
  assign _zz_361_ = _zz_333_[27];
  assign _zz_362_ = _zz_333_[28];
  assign _zz_363_ = _zz_333_[29];
  assign _zz_364_ = _zz_333_[30];
  assign _zz_365_ = _zz_333_[31];
  assign _zz_366_ = _zz_333_[32];
  assign _zz_367_ = _zz_333_[33];
  assign _zz_368_ = _zz_333_[34];
  assign _zz_369_ = _zz_333_[35];
  assign _zz_370_ = _zz_333_[36];
  assign _zz_371_ = _zz_333_[37];
  assign _zz_372_ = _zz_333_[38];
  assign _zz_373_ = _zz_333_[39];
  assign _zz_374_ = _zz_333_[40];
  assign _zz_375_ = _zz_333_[41];
  assign _zz_376_ = _zz_333_[42];
  assign _zz_377_ = _zz_333_[43];
  assign _zz_378_ = _zz_333_[44];
  assign _zz_379_ = _zz_333_[45];
  assign _zz_380_ = _zz_333_[46];
  assign _zz_381_ = _zz_333_[47];
  assign _zz_382_ = _zz_333_[48];
  assign _zz_383_ = _zz_333_[49];
  assign _zz_384_ = (((32'h00000320 <= load_data_area_current_addr) && (load_data_area_current_addr < 32'h00000352)) ? axi4_w_payload_data_regNext : {_zz_2765_,_zz_2766_});
  assign _zz_385_ = _zz_384_[15 : 0];
  assign _zz_386_ = _zz_384_[31 : 16];
  assign _zz_387_ = _zz_2864_[5:0];
  assign _zz_388_ = ({63'd0,(1'b1)} <<< _zz_387_);
  assign _zz_389_ = _zz_388_[0];
  assign _zz_390_ = _zz_388_[1];
  assign _zz_391_ = _zz_388_[2];
  assign _zz_392_ = _zz_388_[3];
  assign _zz_393_ = _zz_388_[4];
  assign _zz_394_ = _zz_388_[5];
  assign _zz_395_ = _zz_388_[6];
  assign _zz_396_ = _zz_388_[7];
  assign _zz_397_ = _zz_388_[8];
  assign _zz_398_ = _zz_388_[9];
  assign _zz_399_ = _zz_388_[10];
  assign _zz_400_ = _zz_388_[11];
  assign _zz_401_ = _zz_388_[12];
  assign _zz_402_ = _zz_388_[13];
  assign _zz_403_ = _zz_388_[14];
  assign _zz_404_ = _zz_388_[15];
  assign _zz_405_ = _zz_388_[16];
  assign _zz_406_ = _zz_388_[17];
  assign _zz_407_ = _zz_388_[18];
  assign _zz_408_ = _zz_388_[19];
  assign _zz_409_ = _zz_388_[20];
  assign _zz_410_ = _zz_388_[21];
  assign _zz_411_ = _zz_388_[22];
  assign _zz_412_ = _zz_388_[23];
  assign _zz_413_ = _zz_388_[24];
  assign _zz_414_ = _zz_388_[25];
  assign _zz_415_ = _zz_388_[26];
  assign _zz_416_ = _zz_388_[27];
  assign _zz_417_ = _zz_388_[28];
  assign _zz_418_ = _zz_388_[29];
  assign _zz_419_ = _zz_388_[30];
  assign _zz_420_ = _zz_388_[31];
  assign _zz_421_ = _zz_388_[32];
  assign _zz_422_ = _zz_388_[33];
  assign _zz_423_ = _zz_388_[34];
  assign _zz_424_ = _zz_388_[35];
  assign _zz_425_ = _zz_388_[36];
  assign _zz_426_ = _zz_388_[37];
  assign _zz_427_ = _zz_388_[38];
  assign _zz_428_ = _zz_388_[39];
  assign _zz_429_ = _zz_388_[40];
  assign _zz_430_ = _zz_388_[41];
  assign _zz_431_ = _zz_388_[42];
  assign _zz_432_ = _zz_388_[43];
  assign _zz_433_ = _zz_388_[44];
  assign _zz_434_ = _zz_388_[45];
  assign _zz_435_ = _zz_388_[46];
  assign _zz_436_ = _zz_388_[47];
  assign _zz_437_ = _zz_388_[48];
  assign _zz_438_ = _zz_388_[49];
  assign _zz_439_ = (((32'h00000226 <= load_data_area_current_addr) && (load_data_area_current_addr < 32'h00000258)) ? axi4_w_payload_data_regNext : {_zz_2767_,_zz_2768_});
  assign _zz_440_ = _zz_439_[15 : 0];
  assign _zz_441_ = _zz_439_[31 : 16];
  assign _zz_442_ = _zz_2865_[5:0];
  assign _zz_443_ = ({63'd0,(1'b1)} <<< _zz_442_);
  assign _zz_444_ = _zz_443_[0];
  assign _zz_445_ = _zz_443_[1];
  assign _zz_446_ = _zz_443_[2];
  assign _zz_447_ = _zz_443_[3];
  assign _zz_448_ = _zz_443_[4];
  assign _zz_449_ = _zz_443_[5];
  assign _zz_450_ = _zz_443_[6];
  assign _zz_451_ = _zz_443_[7];
  assign _zz_452_ = _zz_443_[8];
  assign _zz_453_ = _zz_443_[9];
  assign _zz_454_ = _zz_443_[10];
  assign _zz_455_ = _zz_443_[11];
  assign _zz_456_ = _zz_443_[12];
  assign _zz_457_ = _zz_443_[13];
  assign _zz_458_ = _zz_443_[14];
  assign _zz_459_ = _zz_443_[15];
  assign _zz_460_ = _zz_443_[16];
  assign _zz_461_ = _zz_443_[17];
  assign _zz_462_ = _zz_443_[18];
  assign _zz_463_ = _zz_443_[19];
  assign _zz_464_ = _zz_443_[20];
  assign _zz_465_ = _zz_443_[21];
  assign _zz_466_ = _zz_443_[22];
  assign _zz_467_ = _zz_443_[23];
  assign _zz_468_ = _zz_443_[24];
  assign _zz_469_ = _zz_443_[25];
  assign _zz_470_ = _zz_443_[26];
  assign _zz_471_ = _zz_443_[27];
  assign _zz_472_ = _zz_443_[28];
  assign _zz_473_ = _zz_443_[29];
  assign _zz_474_ = _zz_443_[30];
  assign _zz_475_ = _zz_443_[31];
  assign _zz_476_ = _zz_443_[32];
  assign _zz_477_ = _zz_443_[33];
  assign _zz_478_ = _zz_443_[34];
  assign _zz_479_ = _zz_443_[35];
  assign _zz_480_ = _zz_443_[36];
  assign _zz_481_ = _zz_443_[37];
  assign _zz_482_ = _zz_443_[38];
  assign _zz_483_ = _zz_443_[39];
  assign _zz_484_ = _zz_443_[40];
  assign _zz_485_ = _zz_443_[41];
  assign _zz_486_ = _zz_443_[42];
  assign _zz_487_ = _zz_443_[43];
  assign _zz_488_ = _zz_443_[44];
  assign _zz_489_ = _zz_443_[45];
  assign _zz_490_ = _zz_443_[46];
  assign _zz_491_ = _zz_443_[47];
  assign _zz_492_ = _zz_443_[48];
  assign _zz_493_ = _zz_443_[49];
  assign _zz_494_ = (((32'h000001f4 <= load_data_area_current_addr) && (load_data_area_current_addr < 32'h00000226)) ? axi4_w_payload_data_regNext : {_zz_2769_,_zz_2770_});
  assign _zz_495_ = _zz_494_[15 : 0];
  assign _zz_496_ = _zz_494_[31 : 16];
  assign _zz_497_ = _zz_2866_[5:0];
  assign _zz_498_ = ({63'd0,(1'b1)} <<< _zz_497_);
  assign _zz_499_ = _zz_498_[0];
  assign _zz_500_ = _zz_498_[1];
  assign _zz_501_ = _zz_498_[2];
  assign _zz_502_ = _zz_498_[3];
  assign _zz_503_ = _zz_498_[4];
  assign _zz_504_ = _zz_498_[5];
  assign _zz_505_ = _zz_498_[6];
  assign _zz_506_ = _zz_498_[7];
  assign _zz_507_ = _zz_498_[8];
  assign _zz_508_ = _zz_498_[9];
  assign _zz_509_ = _zz_498_[10];
  assign _zz_510_ = _zz_498_[11];
  assign _zz_511_ = _zz_498_[12];
  assign _zz_512_ = _zz_498_[13];
  assign _zz_513_ = _zz_498_[14];
  assign _zz_514_ = _zz_498_[15];
  assign _zz_515_ = _zz_498_[16];
  assign _zz_516_ = _zz_498_[17];
  assign _zz_517_ = _zz_498_[18];
  assign _zz_518_ = _zz_498_[19];
  assign _zz_519_ = _zz_498_[20];
  assign _zz_520_ = _zz_498_[21];
  assign _zz_521_ = _zz_498_[22];
  assign _zz_522_ = _zz_498_[23];
  assign _zz_523_ = _zz_498_[24];
  assign _zz_524_ = _zz_498_[25];
  assign _zz_525_ = _zz_498_[26];
  assign _zz_526_ = _zz_498_[27];
  assign _zz_527_ = _zz_498_[28];
  assign _zz_528_ = _zz_498_[29];
  assign _zz_529_ = _zz_498_[30];
  assign _zz_530_ = _zz_498_[31];
  assign _zz_531_ = _zz_498_[32];
  assign _zz_532_ = _zz_498_[33];
  assign _zz_533_ = _zz_498_[34];
  assign _zz_534_ = _zz_498_[35];
  assign _zz_535_ = _zz_498_[36];
  assign _zz_536_ = _zz_498_[37];
  assign _zz_537_ = _zz_498_[38];
  assign _zz_538_ = _zz_498_[39];
  assign _zz_539_ = _zz_498_[40];
  assign _zz_540_ = _zz_498_[41];
  assign _zz_541_ = _zz_498_[42];
  assign _zz_542_ = _zz_498_[43];
  assign _zz_543_ = _zz_498_[44];
  assign _zz_544_ = _zz_498_[45];
  assign _zz_545_ = _zz_498_[46];
  assign _zz_546_ = _zz_498_[47];
  assign _zz_547_ = _zz_498_[48];
  assign _zz_548_ = _zz_498_[49];
  assign _zz_549_ = (((32'h0000073a <= load_data_area_current_addr) && (load_data_area_current_addr < 32'h0000076c)) ? axi4_w_payload_data_regNext : {_zz_2771_,_zz_2772_});
  assign _zz_550_ = _zz_549_[15 : 0];
  assign _zz_551_ = _zz_549_[31 : 16];
  assign _zz_552_ = _zz_2867_[5:0];
  assign _zz_553_ = ({63'd0,(1'b1)} <<< _zz_552_);
  assign _zz_554_ = _zz_553_[0];
  assign _zz_555_ = _zz_553_[1];
  assign _zz_556_ = _zz_553_[2];
  assign _zz_557_ = _zz_553_[3];
  assign _zz_558_ = _zz_553_[4];
  assign _zz_559_ = _zz_553_[5];
  assign _zz_560_ = _zz_553_[6];
  assign _zz_561_ = _zz_553_[7];
  assign _zz_562_ = _zz_553_[8];
  assign _zz_563_ = _zz_553_[9];
  assign _zz_564_ = _zz_553_[10];
  assign _zz_565_ = _zz_553_[11];
  assign _zz_566_ = _zz_553_[12];
  assign _zz_567_ = _zz_553_[13];
  assign _zz_568_ = _zz_553_[14];
  assign _zz_569_ = _zz_553_[15];
  assign _zz_570_ = _zz_553_[16];
  assign _zz_571_ = _zz_553_[17];
  assign _zz_572_ = _zz_553_[18];
  assign _zz_573_ = _zz_553_[19];
  assign _zz_574_ = _zz_553_[20];
  assign _zz_575_ = _zz_553_[21];
  assign _zz_576_ = _zz_553_[22];
  assign _zz_577_ = _zz_553_[23];
  assign _zz_578_ = _zz_553_[24];
  assign _zz_579_ = _zz_553_[25];
  assign _zz_580_ = _zz_553_[26];
  assign _zz_581_ = _zz_553_[27];
  assign _zz_582_ = _zz_553_[28];
  assign _zz_583_ = _zz_553_[29];
  assign _zz_584_ = _zz_553_[30];
  assign _zz_585_ = _zz_553_[31];
  assign _zz_586_ = _zz_553_[32];
  assign _zz_587_ = _zz_553_[33];
  assign _zz_588_ = _zz_553_[34];
  assign _zz_589_ = _zz_553_[35];
  assign _zz_590_ = _zz_553_[36];
  assign _zz_591_ = _zz_553_[37];
  assign _zz_592_ = _zz_553_[38];
  assign _zz_593_ = _zz_553_[39];
  assign _zz_594_ = _zz_553_[40];
  assign _zz_595_ = _zz_553_[41];
  assign _zz_596_ = _zz_553_[42];
  assign _zz_597_ = _zz_553_[43];
  assign _zz_598_ = _zz_553_[44];
  assign _zz_599_ = _zz_553_[45];
  assign _zz_600_ = _zz_553_[46];
  assign _zz_601_ = _zz_553_[47];
  assign _zz_602_ = _zz_553_[48];
  assign _zz_603_ = _zz_553_[49];
  assign _zz_604_ = (((32'h0000047e <= load_data_area_current_addr) && (load_data_area_current_addr < 32'h000004b0)) ? axi4_w_payload_data_regNext : {_zz_2773_,_zz_2774_});
  assign _zz_605_ = _zz_604_[15 : 0];
  assign _zz_606_ = _zz_604_[31 : 16];
  assign _zz_607_ = _zz_2868_[5:0];
  assign _zz_608_ = ({63'd0,(1'b1)} <<< _zz_607_);
  assign _zz_609_ = _zz_608_[0];
  assign _zz_610_ = _zz_608_[1];
  assign _zz_611_ = _zz_608_[2];
  assign _zz_612_ = _zz_608_[3];
  assign _zz_613_ = _zz_608_[4];
  assign _zz_614_ = _zz_608_[5];
  assign _zz_615_ = _zz_608_[6];
  assign _zz_616_ = _zz_608_[7];
  assign _zz_617_ = _zz_608_[8];
  assign _zz_618_ = _zz_608_[9];
  assign _zz_619_ = _zz_608_[10];
  assign _zz_620_ = _zz_608_[11];
  assign _zz_621_ = _zz_608_[12];
  assign _zz_622_ = _zz_608_[13];
  assign _zz_623_ = _zz_608_[14];
  assign _zz_624_ = _zz_608_[15];
  assign _zz_625_ = _zz_608_[16];
  assign _zz_626_ = _zz_608_[17];
  assign _zz_627_ = _zz_608_[18];
  assign _zz_628_ = _zz_608_[19];
  assign _zz_629_ = _zz_608_[20];
  assign _zz_630_ = _zz_608_[21];
  assign _zz_631_ = _zz_608_[22];
  assign _zz_632_ = _zz_608_[23];
  assign _zz_633_ = _zz_608_[24];
  assign _zz_634_ = _zz_608_[25];
  assign _zz_635_ = _zz_608_[26];
  assign _zz_636_ = _zz_608_[27];
  assign _zz_637_ = _zz_608_[28];
  assign _zz_638_ = _zz_608_[29];
  assign _zz_639_ = _zz_608_[30];
  assign _zz_640_ = _zz_608_[31];
  assign _zz_641_ = _zz_608_[32];
  assign _zz_642_ = _zz_608_[33];
  assign _zz_643_ = _zz_608_[34];
  assign _zz_644_ = _zz_608_[35];
  assign _zz_645_ = _zz_608_[36];
  assign _zz_646_ = _zz_608_[37];
  assign _zz_647_ = _zz_608_[38];
  assign _zz_648_ = _zz_608_[39];
  assign _zz_649_ = _zz_608_[40];
  assign _zz_650_ = _zz_608_[41];
  assign _zz_651_ = _zz_608_[42];
  assign _zz_652_ = _zz_608_[43];
  assign _zz_653_ = _zz_608_[44];
  assign _zz_654_ = _zz_608_[45];
  assign _zz_655_ = _zz_608_[46];
  assign _zz_656_ = _zz_608_[47];
  assign _zz_657_ = _zz_608_[48];
  assign _zz_658_ = _zz_608_[49];
  assign _zz_659_ = (((32'h0000041a <= load_data_area_current_addr) && (load_data_area_current_addr < 32'h0000044c)) ? axi4_w_payload_data_regNext : {_zz_2775_,_zz_2776_});
  assign _zz_660_ = _zz_659_[15 : 0];
  assign _zz_661_ = _zz_659_[31 : 16];
  assign _zz_662_ = _zz_2869_[5:0];
  assign _zz_663_ = ({63'd0,(1'b1)} <<< _zz_662_);
  assign _zz_664_ = _zz_663_[0];
  assign _zz_665_ = _zz_663_[1];
  assign _zz_666_ = _zz_663_[2];
  assign _zz_667_ = _zz_663_[3];
  assign _zz_668_ = _zz_663_[4];
  assign _zz_669_ = _zz_663_[5];
  assign _zz_670_ = _zz_663_[6];
  assign _zz_671_ = _zz_663_[7];
  assign _zz_672_ = _zz_663_[8];
  assign _zz_673_ = _zz_663_[9];
  assign _zz_674_ = _zz_663_[10];
  assign _zz_675_ = _zz_663_[11];
  assign _zz_676_ = _zz_663_[12];
  assign _zz_677_ = _zz_663_[13];
  assign _zz_678_ = _zz_663_[14];
  assign _zz_679_ = _zz_663_[15];
  assign _zz_680_ = _zz_663_[16];
  assign _zz_681_ = _zz_663_[17];
  assign _zz_682_ = _zz_663_[18];
  assign _zz_683_ = _zz_663_[19];
  assign _zz_684_ = _zz_663_[20];
  assign _zz_685_ = _zz_663_[21];
  assign _zz_686_ = _zz_663_[22];
  assign _zz_687_ = _zz_663_[23];
  assign _zz_688_ = _zz_663_[24];
  assign _zz_689_ = _zz_663_[25];
  assign _zz_690_ = _zz_663_[26];
  assign _zz_691_ = _zz_663_[27];
  assign _zz_692_ = _zz_663_[28];
  assign _zz_693_ = _zz_663_[29];
  assign _zz_694_ = _zz_663_[30];
  assign _zz_695_ = _zz_663_[31];
  assign _zz_696_ = _zz_663_[32];
  assign _zz_697_ = _zz_663_[33];
  assign _zz_698_ = _zz_663_[34];
  assign _zz_699_ = _zz_663_[35];
  assign _zz_700_ = _zz_663_[36];
  assign _zz_701_ = _zz_663_[37];
  assign _zz_702_ = _zz_663_[38];
  assign _zz_703_ = _zz_663_[39];
  assign _zz_704_ = _zz_663_[40];
  assign _zz_705_ = _zz_663_[41];
  assign _zz_706_ = _zz_663_[42];
  assign _zz_707_ = _zz_663_[43];
  assign _zz_708_ = _zz_663_[44];
  assign _zz_709_ = _zz_663_[45];
  assign _zz_710_ = _zz_663_[46];
  assign _zz_711_ = _zz_663_[47];
  assign _zz_712_ = _zz_663_[48];
  assign _zz_713_ = _zz_663_[49];
  assign _zz_714_ = (((32'h000008ca <= load_data_area_current_addr) && (load_data_area_current_addr < 32'h000008fc)) ? axi4_w_payload_data_regNext : {_zz_2777_,_zz_2778_});
  assign _zz_715_ = _zz_714_[15 : 0];
  assign _zz_716_ = _zz_714_[31 : 16];
  assign _zz_717_ = _zz_2870_[5:0];
  assign _zz_718_ = ({63'd0,(1'b1)} <<< _zz_717_);
  assign _zz_719_ = _zz_718_[0];
  assign _zz_720_ = _zz_718_[1];
  assign _zz_721_ = _zz_718_[2];
  assign _zz_722_ = _zz_718_[3];
  assign _zz_723_ = _zz_718_[4];
  assign _zz_724_ = _zz_718_[5];
  assign _zz_725_ = _zz_718_[6];
  assign _zz_726_ = _zz_718_[7];
  assign _zz_727_ = _zz_718_[8];
  assign _zz_728_ = _zz_718_[9];
  assign _zz_729_ = _zz_718_[10];
  assign _zz_730_ = _zz_718_[11];
  assign _zz_731_ = _zz_718_[12];
  assign _zz_732_ = _zz_718_[13];
  assign _zz_733_ = _zz_718_[14];
  assign _zz_734_ = _zz_718_[15];
  assign _zz_735_ = _zz_718_[16];
  assign _zz_736_ = _zz_718_[17];
  assign _zz_737_ = _zz_718_[18];
  assign _zz_738_ = _zz_718_[19];
  assign _zz_739_ = _zz_718_[20];
  assign _zz_740_ = _zz_718_[21];
  assign _zz_741_ = _zz_718_[22];
  assign _zz_742_ = _zz_718_[23];
  assign _zz_743_ = _zz_718_[24];
  assign _zz_744_ = _zz_718_[25];
  assign _zz_745_ = _zz_718_[26];
  assign _zz_746_ = _zz_718_[27];
  assign _zz_747_ = _zz_718_[28];
  assign _zz_748_ = _zz_718_[29];
  assign _zz_749_ = _zz_718_[30];
  assign _zz_750_ = _zz_718_[31];
  assign _zz_751_ = _zz_718_[32];
  assign _zz_752_ = _zz_718_[33];
  assign _zz_753_ = _zz_718_[34];
  assign _zz_754_ = _zz_718_[35];
  assign _zz_755_ = _zz_718_[36];
  assign _zz_756_ = _zz_718_[37];
  assign _zz_757_ = _zz_718_[38];
  assign _zz_758_ = _zz_718_[39];
  assign _zz_759_ = _zz_718_[40];
  assign _zz_760_ = _zz_718_[41];
  assign _zz_761_ = _zz_718_[42];
  assign _zz_762_ = _zz_718_[43];
  assign _zz_763_ = _zz_718_[44];
  assign _zz_764_ = _zz_718_[45];
  assign _zz_765_ = _zz_718_[46];
  assign _zz_766_ = _zz_718_[47];
  assign _zz_767_ = _zz_718_[48];
  assign _zz_768_ = _zz_718_[49];
  assign _zz_769_ = (((32'h00000898 <= load_data_area_current_addr) && (load_data_area_current_addr < 32'h000008ca)) ? axi4_w_payload_data_regNext : {_zz_2779_,_zz_2780_});
  assign _zz_770_ = _zz_769_[15 : 0];
  assign _zz_771_ = _zz_769_[31 : 16];
  assign _zz_772_ = _zz_2871_[5:0];
  assign _zz_773_ = ({63'd0,(1'b1)} <<< _zz_772_);
  assign _zz_774_ = _zz_773_[0];
  assign _zz_775_ = _zz_773_[1];
  assign _zz_776_ = _zz_773_[2];
  assign _zz_777_ = _zz_773_[3];
  assign _zz_778_ = _zz_773_[4];
  assign _zz_779_ = _zz_773_[5];
  assign _zz_780_ = _zz_773_[6];
  assign _zz_781_ = _zz_773_[7];
  assign _zz_782_ = _zz_773_[8];
  assign _zz_783_ = _zz_773_[9];
  assign _zz_784_ = _zz_773_[10];
  assign _zz_785_ = _zz_773_[11];
  assign _zz_786_ = _zz_773_[12];
  assign _zz_787_ = _zz_773_[13];
  assign _zz_788_ = _zz_773_[14];
  assign _zz_789_ = _zz_773_[15];
  assign _zz_790_ = _zz_773_[16];
  assign _zz_791_ = _zz_773_[17];
  assign _zz_792_ = _zz_773_[18];
  assign _zz_793_ = _zz_773_[19];
  assign _zz_794_ = _zz_773_[20];
  assign _zz_795_ = _zz_773_[21];
  assign _zz_796_ = _zz_773_[22];
  assign _zz_797_ = _zz_773_[23];
  assign _zz_798_ = _zz_773_[24];
  assign _zz_799_ = _zz_773_[25];
  assign _zz_800_ = _zz_773_[26];
  assign _zz_801_ = _zz_773_[27];
  assign _zz_802_ = _zz_773_[28];
  assign _zz_803_ = _zz_773_[29];
  assign _zz_804_ = _zz_773_[30];
  assign _zz_805_ = _zz_773_[31];
  assign _zz_806_ = _zz_773_[32];
  assign _zz_807_ = _zz_773_[33];
  assign _zz_808_ = _zz_773_[34];
  assign _zz_809_ = _zz_773_[35];
  assign _zz_810_ = _zz_773_[36];
  assign _zz_811_ = _zz_773_[37];
  assign _zz_812_ = _zz_773_[38];
  assign _zz_813_ = _zz_773_[39];
  assign _zz_814_ = _zz_773_[40];
  assign _zz_815_ = _zz_773_[41];
  assign _zz_816_ = _zz_773_[42];
  assign _zz_817_ = _zz_773_[43];
  assign _zz_818_ = _zz_773_[44];
  assign _zz_819_ = _zz_773_[45];
  assign _zz_820_ = _zz_773_[46];
  assign _zz_821_ = _zz_773_[47];
  assign _zz_822_ = _zz_773_[48];
  assign _zz_823_ = _zz_773_[49];
  assign _zz_824_ = (((32'h000004b0 <= load_data_area_current_addr) && (load_data_area_current_addr < 32'h000004e2)) ? axi4_w_payload_data_regNext : {_zz_2781_,_zz_2782_});
  assign _zz_825_ = _zz_824_[15 : 0];
  assign _zz_826_ = _zz_824_[31 : 16];
  assign _zz_827_ = _zz_2872_[5:0];
  assign _zz_828_ = ({63'd0,(1'b1)} <<< _zz_827_);
  assign _zz_829_ = _zz_828_[0];
  assign _zz_830_ = _zz_828_[1];
  assign _zz_831_ = _zz_828_[2];
  assign _zz_832_ = _zz_828_[3];
  assign _zz_833_ = _zz_828_[4];
  assign _zz_834_ = _zz_828_[5];
  assign _zz_835_ = _zz_828_[6];
  assign _zz_836_ = _zz_828_[7];
  assign _zz_837_ = _zz_828_[8];
  assign _zz_838_ = _zz_828_[9];
  assign _zz_839_ = _zz_828_[10];
  assign _zz_840_ = _zz_828_[11];
  assign _zz_841_ = _zz_828_[12];
  assign _zz_842_ = _zz_828_[13];
  assign _zz_843_ = _zz_828_[14];
  assign _zz_844_ = _zz_828_[15];
  assign _zz_845_ = _zz_828_[16];
  assign _zz_846_ = _zz_828_[17];
  assign _zz_847_ = _zz_828_[18];
  assign _zz_848_ = _zz_828_[19];
  assign _zz_849_ = _zz_828_[20];
  assign _zz_850_ = _zz_828_[21];
  assign _zz_851_ = _zz_828_[22];
  assign _zz_852_ = _zz_828_[23];
  assign _zz_853_ = _zz_828_[24];
  assign _zz_854_ = _zz_828_[25];
  assign _zz_855_ = _zz_828_[26];
  assign _zz_856_ = _zz_828_[27];
  assign _zz_857_ = _zz_828_[28];
  assign _zz_858_ = _zz_828_[29];
  assign _zz_859_ = _zz_828_[30];
  assign _zz_860_ = _zz_828_[31];
  assign _zz_861_ = _zz_828_[32];
  assign _zz_862_ = _zz_828_[33];
  assign _zz_863_ = _zz_828_[34];
  assign _zz_864_ = _zz_828_[35];
  assign _zz_865_ = _zz_828_[36];
  assign _zz_866_ = _zz_828_[37];
  assign _zz_867_ = _zz_828_[38];
  assign _zz_868_ = _zz_828_[39];
  assign _zz_869_ = _zz_828_[40];
  assign _zz_870_ = _zz_828_[41];
  assign _zz_871_ = _zz_828_[42];
  assign _zz_872_ = _zz_828_[43];
  assign _zz_873_ = _zz_828_[44];
  assign _zz_874_ = _zz_828_[45];
  assign _zz_875_ = _zz_828_[46];
  assign _zz_876_ = _zz_828_[47];
  assign _zz_877_ = _zz_828_[48];
  assign _zz_878_ = _zz_828_[49];
  assign _zz_879_ = (((32'h00000834 <= load_data_area_current_addr) && (load_data_area_current_addr < 32'h00000866)) ? axi4_w_payload_data_regNext : {_zz_2783_,_zz_2784_});
  assign _zz_880_ = _zz_879_[15 : 0];
  assign _zz_881_ = _zz_879_[31 : 16];
  assign _zz_882_ = _zz_2873_[5:0];
  assign _zz_883_ = ({63'd0,(1'b1)} <<< _zz_882_);
  assign _zz_884_ = _zz_883_[0];
  assign _zz_885_ = _zz_883_[1];
  assign _zz_886_ = _zz_883_[2];
  assign _zz_887_ = _zz_883_[3];
  assign _zz_888_ = _zz_883_[4];
  assign _zz_889_ = _zz_883_[5];
  assign _zz_890_ = _zz_883_[6];
  assign _zz_891_ = _zz_883_[7];
  assign _zz_892_ = _zz_883_[8];
  assign _zz_893_ = _zz_883_[9];
  assign _zz_894_ = _zz_883_[10];
  assign _zz_895_ = _zz_883_[11];
  assign _zz_896_ = _zz_883_[12];
  assign _zz_897_ = _zz_883_[13];
  assign _zz_898_ = _zz_883_[14];
  assign _zz_899_ = _zz_883_[15];
  assign _zz_900_ = _zz_883_[16];
  assign _zz_901_ = _zz_883_[17];
  assign _zz_902_ = _zz_883_[18];
  assign _zz_903_ = _zz_883_[19];
  assign _zz_904_ = _zz_883_[20];
  assign _zz_905_ = _zz_883_[21];
  assign _zz_906_ = _zz_883_[22];
  assign _zz_907_ = _zz_883_[23];
  assign _zz_908_ = _zz_883_[24];
  assign _zz_909_ = _zz_883_[25];
  assign _zz_910_ = _zz_883_[26];
  assign _zz_911_ = _zz_883_[27];
  assign _zz_912_ = _zz_883_[28];
  assign _zz_913_ = _zz_883_[29];
  assign _zz_914_ = _zz_883_[30];
  assign _zz_915_ = _zz_883_[31];
  assign _zz_916_ = _zz_883_[32];
  assign _zz_917_ = _zz_883_[33];
  assign _zz_918_ = _zz_883_[34];
  assign _zz_919_ = _zz_883_[35];
  assign _zz_920_ = _zz_883_[36];
  assign _zz_921_ = _zz_883_[37];
  assign _zz_922_ = _zz_883_[38];
  assign _zz_923_ = _zz_883_[39];
  assign _zz_924_ = _zz_883_[40];
  assign _zz_925_ = _zz_883_[41];
  assign _zz_926_ = _zz_883_[42];
  assign _zz_927_ = _zz_883_[43];
  assign _zz_928_ = _zz_883_[44];
  assign _zz_929_ = _zz_883_[45];
  assign _zz_930_ = _zz_883_[46];
  assign _zz_931_ = _zz_883_[47];
  assign _zz_932_ = _zz_883_[48];
  assign _zz_933_ = _zz_883_[49];
  assign _zz_934_ = (((32'h000005dc <= load_data_area_current_addr) && (load_data_area_current_addr < 32'h0000060e)) ? axi4_w_payload_data_regNext : {_zz_2785_,_zz_2786_});
  assign _zz_935_ = _zz_934_[15 : 0];
  assign _zz_936_ = _zz_934_[31 : 16];
  assign _zz_937_ = _zz_2874_[5:0];
  assign _zz_938_ = ({63'd0,(1'b1)} <<< _zz_937_);
  assign _zz_939_ = _zz_938_[0];
  assign _zz_940_ = _zz_938_[1];
  assign _zz_941_ = _zz_938_[2];
  assign _zz_942_ = _zz_938_[3];
  assign _zz_943_ = _zz_938_[4];
  assign _zz_944_ = _zz_938_[5];
  assign _zz_945_ = _zz_938_[6];
  assign _zz_946_ = _zz_938_[7];
  assign _zz_947_ = _zz_938_[8];
  assign _zz_948_ = _zz_938_[9];
  assign _zz_949_ = _zz_938_[10];
  assign _zz_950_ = _zz_938_[11];
  assign _zz_951_ = _zz_938_[12];
  assign _zz_952_ = _zz_938_[13];
  assign _zz_953_ = _zz_938_[14];
  assign _zz_954_ = _zz_938_[15];
  assign _zz_955_ = _zz_938_[16];
  assign _zz_956_ = _zz_938_[17];
  assign _zz_957_ = _zz_938_[18];
  assign _zz_958_ = _zz_938_[19];
  assign _zz_959_ = _zz_938_[20];
  assign _zz_960_ = _zz_938_[21];
  assign _zz_961_ = _zz_938_[22];
  assign _zz_962_ = _zz_938_[23];
  assign _zz_963_ = _zz_938_[24];
  assign _zz_964_ = _zz_938_[25];
  assign _zz_965_ = _zz_938_[26];
  assign _zz_966_ = _zz_938_[27];
  assign _zz_967_ = _zz_938_[28];
  assign _zz_968_ = _zz_938_[29];
  assign _zz_969_ = _zz_938_[30];
  assign _zz_970_ = _zz_938_[31];
  assign _zz_971_ = _zz_938_[32];
  assign _zz_972_ = _zz_938_[33];
  assign _zz_973_ = _zz_938_[34];
  assign _zz_974_ = _zz_938_[35];
  assign _zz_975_ = _zz_938_[36];
  assign _zz_976_ = _zz_938_[37];
  assign _zz_977_ = _zz_938_[38];
  assign _zz_978_ = _zz_938_[39];
  assign _zz_979_ = _zz_938_[40];
  assign _zz_980_ = _zz_938_[41];
  assign _zz_981_ = _zz_938_[42];
  assign _zz_982_ = _zz_938_[43];
  assign _zz_983_ = _zz_938_[44];
  assign _zz_984_ = _zz_938_[45];
  assign _zz_985_ = _zz_938_[46];
  assign _zz_986_ = _zz_938_[47];
  assign _zz_987_ = _zz_938_[48];
  assign _zz_988_ = _zz_938_[49];
  assign _zz_989_ = (((32'h00000640 <= load_data_area_current_addr) && (load_data_area_current_addr < 32'h00000672)) ? axi4_w_payload_data_regNext : {_zz_2787_,_zz_2788_});
  assign _zz_990_ = _zz_989_[15 : 0];
  assign _zz_991_ = _zz_989_[31 : 16];
  assign _zz_992_ = _zz_2875_[5:0];
  assign _zz_993_ = ({63'd0,(1'b1)} <<< _zz_992_);
  assign _zz_994_ = _zz_993_[0];
  assign _zz_995_ = _zz_993_[1];
  assign _zz_996_ = _zz_993_[2];
  assign _zz_997_ = _zz_993_[3];
  assign _zz_998_ = _zz_993_[4];
  assign _zz_999_ = _zz_993_[5];
  assign _zz_1000_ = _zz_993_[6];
  assign _zz_1001_ = _zz_993_[7];
  assign _zz_1002_ = _zz_993_[8];
  assign _zz_1003_ = _zz_993_[9];
  assign _zz_1004_ = _zz_993_[10];
  assign _zz_1005_ = _zz_993_[11];
  assign _zz_1006_ = _zz_993_[12];
  assign _zz_1007_ = _zz_993_[13];
  assign _zz_1008_ = _zz_993_[14];
  assign _zz_1009_ = _zz_993_[15];
  assign _zz_1010_ = _zz_993_[16];
  assign _zz_1011_ = _zz_993_[17];
  assign _zz_1012_ = _zz_993_[18];
  assign _zz_1013_ = _zz_993_[19];
  assign _zz_1014_ = _zz_993_[20];
  assign _zz_1015_ = _zz_993_[21];
  assign _zz_1016_ = _zz_993_[22];
  assign _zz_1017_ = _zz_993_[23];
  assign _zz_1018_ = _zz_993_[24];
  assign _zz_1019_ = _zz_993_[25];
  assign _zz_1020_ = _zz_993_[26];
  assign _zz_1021_ = _zz_993_[27];
  assign _zz_1022_ = _zz_993_[28];
  assign _zz_1023_ = _zz_993_[29];
  assign _zz_1024_ = _zz_993_[30];
  assign _zz_1025_ = _zz_993_[31];
  assign _zz_1026_ = _zz_993_[32];
  assign _zz_1027_ = _zz_993_[33];
  assign _zz_1028_ = _zz_993_[34];
  assign _zz_1029_ = _zz_993_[35];
  assign _zz_1030_ = _zz_993_[36];
  assign _zz_1031_ = _zz_993_[37];
  assign _zz_1032_ = _zz_993_[38];
  assign _zz_1033_ = _zz_993_[39];
  assign _zz_1034_ = _zz_993_[40];
  assign _zz_1035_ = _zz_993_[41];
  assign _zz_1036_ = _zz_993_[42];
  assign _zz_1037_ = _zz_993_[43];
  assign _zz_1038_ = _zz_993_[44];
  assign _zz_1039_ = _zz_993_[45];
  assign _zz_1040_ = _zz_993_[46];
  assign _zz_1041_ = _zz_993_[47];
  assign _zz_1042_ = _zz_993_[48];
  assign _zz_1043_ = _zz_993_[49];
  assign _zz_1044_ = (((32'h00000546 <= load_data_area_current_addr) && (load_data_area_current_addr < 32'h00000578)) ? axi4_w_payload_data_regNext : {_zz_2789_,_zz_2790_});
  assign _zz_1045_ = _zz_1044_[15 : 0];
  assign _zz_1046_ = _zz_1044_[31 : 16];
  assign _zz_1047_ = _zz_2876_[5:0];
  assign _zz_1048_ = ({63'd0,(1'b1)} <<< _zz_1047_);
  assign _zz_1049_ = _zz_1048_[0];
  assign _zz_1050_ = _zz_1048_[1];
  assign _zz_1051_ = _zz_1048_[2];
  assign _zz_1052_ = _zz_1048_[3];
  assign _zz_1053_ = _zz_1048_[4];
  assign _zz_1054_ = _zz_1048_[5];
  assign _zz_1055_ = _zz_1048_[6];
  assign _zz_1056_ = _zz_1048_[7];
  assign _zz_1057_ = _zz_1048_[8];
  assign _zz_1058_ = _zz_1048_[9];
  assign _zz_1059_ = _zz_1048_[10];
  assign _zz_1060_ = _zz_1048_[11];
  assign _zz_1061_ = _zz_1048_[12];
  assign _zz_1062_ = _zz_1048_[13];
  assign _zz_1063_ = _zz_1048_[14];
  assign _zz_1064_ = _zz_1048_[15];
  assign _zz_1065_ = _zz_1048_[16];
  assign _zz_1066_ = _zz_1048_[17];
  assign _zz_1067_ = _zz_1048_[18];
  assign _zz_1068_ = _zz_1048_[19];
  assign _zz_1069_ = _zz_1048_[20];
  assign _zz_1070_ = _zz_1048_[21];
  assign _zz_1071_ = _zz_1048_[22];
  assign _zz_1072_ = _zz_1048_[23];
  assign _zz_1073_ = _zz_1048_[24];
  assign _zz_1074_ = _zz_1048_[25];
  assign _zz_1075_ = _zz_1048_[26];
  assign _zz_1076_ = _zz_1048_[27];
  assign _zz_1077_ = _zz_1048_[28];
  assign _zz_1078_ = _zz_1048_[29];
  assign _zz_1079_ = _zz_1048_[30];
  assign _zz_1080_ = _zz_1048_[31];
  assign _zz_1081_ = _zz_1048_[32];
  assign _zz_1082_ = _zz_1048_[33];
  assign _zz_1083_ = _zz_1048_[34];
  assign _zz_1084_ = _zz_1048_[35];
  assign _zz_1085_ = _zz_1048_[36];
  assign _zz_1086_ = _zz_1048_[37];
  assign _zz_1087_ = _zz_1048_[38];
  assign _zz_1088_ = _zz_1048_[39];
  assign _zz_1089_ = _zz_1048_[40];
  assign _zz_1090_ = _zz_1048_[41];
  assign _zz_1091_ = _zz_1048_[42];
  assign _zz_1092_ = _zz_1048_[43];
  assign _zz_1093_ = _zz_1048_[44];
  assign _zz_1094_ = _zz_1048_[45];
  assign _zz_1095_ = _zz_1048_[46];
  assign _zz_1096_ = _zz_1048_[47];
  assign _zz_1097_ = _zz_1048_[48];
  assign _zz_1098_ = _zz_1048_[49];
  assign _zz_1099_ = (((32'h000004e2 <= load_data_area_current_addr) && (load_data_area_current_addr < 32'h00000514)) ? axi4_w_payload_data_regNext : {_zz_2791_,_zz_2792_});
  assign _zz_1100_ = _zz_1099_[15 : 0];
  assign _zz_1101_ = _zz_1099_[31 : 16];
  assign _zz_1102_ = _zz_2877_[5:0];
  assign _zz_1103_ = ({63'd0,(1'b1)} <<< _zz_1102_);
  assign _zz_1104_ = _zz_1103_[0];
  assign _zz_1105_ = _zz_1103_[1];
  assign _zz_1106_ = _zz_1103_[2];
  assign _zz_1107_ = _zz_1103_[3];
  assign _zz_1108_ = _zz_1103_[4];
  assign _zz_1109_ = _zz_1103_[5];
  assign _zz_1110_ = _zz_1103_[6];
  assign _zz_1111_ = _zz_1103_[7];
  assign _zz_1112_ = _zz_1103_[8];
  assign _zz_1113_ = _zz_1103_[9];
  assign _zz_1114_ = _zz_1103_[10];
  assign _zz_1115_ = _zz_1103_[11];
  assign _zz_1116_ = _zz_1103_[12];
  assign _zz_1117_ = _zz_1103_[13];
  assign _zz_1118_ = _zz_1103_[14];
  assign _zz_1119_ = _zz_1103_[15];
  assign _zz_1120_ = _zz_1103_[16];
  assign _zz_1121_ = _zz_1103_[17];
  assign _zz_1122_ = _zz_1103_[18];
  assign _zz_1123_ = _zz_1103_[19];
  assign _zz_1124_ = _zz_1103_[20];
  assign _zz_1125_ = _zz_1103_[21];
  assign _zz_1126_ = _zz_1103_[22];
  assign _zz_1127_ = _zz_1103_[23];
  assign _zz_1128_ = _zz_1103_[24];
  assign _zz_1129_ = _zz_1103_[25];
  assign _zz_1130_ = _zz_1103_[26];
  assign _zz_1131_ = _zz_1103_[27];
  assign _zz_1132_ = _zz_1103_[28];
  assign _zz_1133_ = _zz_1103_[29];
  assign _zz_1134_ = _zz_1103_[30];
  assign _zz_1135_ = _zz_1103_[31];
  assign _zz_1136_ = _zz_1103_[32];
  assign _zz_1137_ = _zz_1103_[33];
  assign _zz_1138_ = _zz_1103_[34];
  assign _zz_1139_ = _zz_1103_[35];
  assign _zz_1140_ = _zz_1103_[36];
  assign _zz_1141_ = _zz_1103_[37];
  assign _zz_1142_ = _zz_1103_[38];
  assign _zz_1143_ = _zz_1103_[39];
  assign _zz_1144_ = _zz_1103_[40];
  assign _zz_1145_ = _zz_1103_[41];
  assign _zz_1146_ = _zz_1103_[42];
  assign _zz_1147_ = _zz_1103_[43];
  assign _zz_1148_ = _zz_1103_[44];
  assign _zz_1149_ = _zz_1103_[45];
  assign _zz_1150_ = _zz_1103_[46];
  assign _zz_1151_ = _zz_1103_[47];
  assign _zz_1152_ = _zz_1103_[48];
  assign _zz_1153_ = _zz_1103_[49];
  assign _zz_1154_ = (((32'h00000258 <= load_data_area_current_addr) && (load_data_area_current_addr < 32'h0000028a)) ? axi4_w_payload_data_regNext : {_zz_2793_,_zz_2794_});
  assign _zz_1155_ = _zz_1154_[15 : 0];
  assign _zz_1156_ = _zz_1154_[31 : 16];
  assign _zz_1157_ = _zz_2878_[5:0];
  assign _zz_1158_ = ({63'd0,(1'b1)} <<< _zz_1157_);
  assign _zz_1159_ = _zz_1158_[0];
  assign _zz_1160_ = _zz_1158_[1];
  assign _zz_1161_ = _zz_1158_[2];
  assign _zz_1162_ = _zz_1158_[3];
  assign _zz_1163_ = _zz_1158_[4];
  assign _zz_1164_ = _zz_1158_[5];
  assign _zz_1165_ = _zz_1158_[6];
  assign _zz_1166_ = _zz_1158_[7];
  assign _zz_1167_ = _zz_1158_[8];
  assign _zz_1168_ = _zz_1158_[9];
  assign _zz_1169_ = _zz_1158_[10];
  assign _zz_1170_ = _zz_1158_[11];
  assign _zz_1171_ = _zz_1158_[12];
  assign _zz_1172_ = _zz_1158_[13];
  assign _zz_1173_ = _zz_1158_[14];
  assign _zz_1174_ = _zz_1158_[15];
  assign _zz_1175_ = _zz_1158_[16];
  assign _zz_1176_ = _zz_1158_[17];
  assign _zz_1177_ = _zz_1158_[18];
  assign _zz_1178_ = _zz_1158_[19];
  assign _zz_1179_ = _zz_1158_[20];
  assign _zz_1180_ = _zz_1158_[21];
  assign _zz_1181_ = _zz_1158_[22];
  assign _zz_1182_ = _zz_1158_[23];
  assign _zz_1183_ = _zz_1158_[24];
  assign _zz_1184_ = _zz_1158_[25];
  assign _zz_1185_ = _zz_1158_[26];
  assign _zz_1186_ = _zz_1158_[27];
  assign _zz_1187_ = _zz_1158_[28];
  assign _zz_1188_ = _zz_1158_[29];
  assign _zz_1189_ = _zz_1158_[30];
  assign _zz_1190_ = _zz_1158_[31];
  assign _zz_1191_ = _zz_1158_[32];
  assign _zz_1192_ = _zz_1158_[33];
  assign _zz_1193_ = _zz_1158_[34];
  assign _zz_1194_ = _zz_1158_[35];
  assign _zz_1195_ = _zz_1158_[36];
  assign _zz_1196_ = _zz_1158_[37];
  assign _zz_1197_ = _zz_1158_[38];
  assign _zz_1198_ = _zz_1158_[39];
  assign _zz_1199_ = _zz_1158_[40];
  assign _zz_1200_ = _zz_1158_[41];
  assign _zz_1201_ = _zz_1158_[42];
  assign _zz_1202_ = _zz_1158_[43];
  assign _zz_1203_ = _zz_1158_[44];
  assign _zz_1204_ = _zz_1158_[45];
  assign _zz_1205_ = _zz_1158_[46];
  assign _zz_1206_ = _zz_1158_[47];
  assign _zz_1207_ = _zz_1158_[48];
  assign _zz_1208_ = _zz_1158_[49];
  assign _zz_1209_ = (((32'h00000992 <= load_data_area_current_addr) && (load_data_area_current_addr < 32'h000009c4)) ? axi4_w_payload_data_regNext : {_zz_2795_,_zz_2796_});
  assign _zz_1210_ = _zz_1209_[15 : 0];
  assign _zz_1211_ = _zz_1209_[31 : 16];
  assign _zz_1212_ = _zz_2879_[5:0];
  assign _zz_1213_ = ({63'd0,(1'b1)} <<< _zz_1212_);
  assign _zz_1214_ = _zz_1213_[0];
  assign _zz_1215_ = _zz_1213_[1];
  assign _zz_1216_ = _zz_1213_[2];
  assign _zz_1217_ = _zz_1213_[3];
  assign _zz_1218_ = _zz_1213_[4];
  assign _zz_1219_ = _zz_1213_[5];
  assign _zz_1220_ = _zz_1213_[6];
  assign _zz_1221_ = _zz_1213_[7];
  assign _zz_1222_ = _zz_1213_[8];
  assign _zz_1223_ = _zz_1213_[9];
  assign _zz_1224_ = _zz_1213_[10];
  assign _zz_1225_ = _zz_1213_[11];
  assign _zz_1226_ = _zz_1213_[12];
  assign _zz_1227_ = _zz_1213_[13];
  assign _zz_1228_ = _zz_1213_[14];
  assign _zz_1229_ = _zz_1213_[15];
  assign _zz_1230_ = _zz_1213_[16];
  assign _zz_1231_ = _zz_1213_[17];
  assign _zz_1232_ = _zz_1213_[18];
  assign _zz_1233_ = _zz_1213_[19];
  assign _zz_1234_ = _zz_1213_[20];
  assign _zz_1235_ = _zz_1213_[21];
  assign _zz_1236_ = _zz_1213_[22];
  assign _zz_1237_ = _zz_1213_[23];
  assign _zz_1238_ = _zz_1213_[24];
  assign _zz_1239_ = _zz_1213_[25];
  assign _zz_1240_ = _zz_1213_[26];
  assign _zz_1241_ = _zz_1213_[27];
  assign _zz_1242_ = _zz_1213_[28];
  assign _zz_1243_ = _zz_1213_[29];
  assign _zz_1244_ = _zz_1213_[30];
  assign _zz_1245_ = _zz_1213_[31];
  assign _zz_1246_ = _zz_1213_[32];
  assign _zz_1247_ = _zz_1213_[33];
  assign _zz_1248_ = _zz_1213_[34];
  assign _zz_1249_ = _zz_1213_[35];
  assign _zz_1250_ = _zz_1213_[36];
  assign _zz_1251_ = _zz_1213_[37];
  assign _zz_1252_ = _zz_1213_[38];
  assign _zz_1253_ = _zz_1213_[39];
  assign _zz_1254_ = _zz_1213_[40];
  assign _zz_1255_ = _zz_1213_[41];
  assign _zz_1256_ = _zz_1213_[42];
  assign _zz_1257_ = _zz_1213_[43];
  assign _zz_1258_ = _zz_1213_[44];
  assign _zz_1259_ = _zz_1213_[45];
  assign _zz_1260_ = _zz_1213_[46];
  assign _zz_1261_ = _zz_1213_[47];
  assign _zz_1262_ = _zz_1213_[48];
  assign _zz_1263_ = _zz_1213_[49];
  assign _zz_1264_ = (((32'h000003e8 <= load_data_area_current_addr) && (load_data_area_current_addr < 32'h0000041a)) ? axi4_w_payload_data_regNext : {_zz_2797_,_zz_2798_});
  assign _zz_1265_ = _zz_1264_[15 : 0];
  assign _zz_1266_ = _zz_1264_[31 : 16];
  assign _zz_1267_ = _zz_2880_[5:0];
  assign _zz_1268_ = ({63'd0,(1'b1)} <<< _zz_1267_);
  assign _zz_1269_ = _zz_1268_[0];
  assign _zz_1270_ = _zz_1268_[1];
  assign _zz_1271_ = _zz_1268_[2];
  assign _zz_1272_ = _zz_1268_[3];
  assign _zz_1273_ = _zz_1268_[4];
  assign _zz_1274_ = _zz_1268_[5];
  assign _zz_1275_ = _zz_1268_[6];
  assign _zz_1276_ = _zz_1268_[7];
  assign _zz_1277_ = _zz_1268_[8];
  assign _zz_1278_ = _zz_1268_[9];
  assign _zz_1279_ = _zz_1268_[10];
  assign _zz_1280_ = _zz_1268_[11];
  assign _zz_1281_ = _zz_1268_[12];
  assign _zz_1282_ = _zz_1268_[13];
  assign _zz_1283_ = _zz_1268_[14];
  assign _zz_1284_ = _zz_1268_[15];
  assign _zz_1285_ = _zz_1268_[16];
  assign _zz_1286_ = _zz_1268_[17];
  assign _zz_1287_ = _zz_1268_[18];
  assign _zz_1288_ = _zz_1268_[19];
  assign _zz_1289_ = _zz_1268_[20];
  assign _zz_1290_ = _zz_1268_[21];
  assign _zz_1291_ = _zz_1268_[22];
  assign _zz_1292_ = _zz_1268_[23];
  assign _zz_1293_ = _zz_1268_[24];
  assign _zz_1294_ = _zz_1268_[25];
  assign _zz_1295_ = _zz_1268_[26];
  assign _zz_1296_ = _zz_1268_[27];
  assign _zz_1297_ = _zz_1268_[28];
  assign _zz_1298_ = _zz_1268_[29];
  assign _zz_1299_ = _zz_1268_[30];
  assign _zz_1300_ = _zz_1268_[31];
  assign _zz_1301_ = _zz_1268_[32];
  assign _zz_1302_ = _zz_1268_[33];
  assign _zz_1303_ = _zz_1268_[34];
  assign _zz_1304_ = _zz_1268_[35];
  assign _zz_1305_ = _zz_1268_[36];
  assign _zz_1306_ = _zz_1268_[37];
  assign _zz_1307_ = _zz_1268_[38];
  assign _zz_1308_ = _zz_1268_[39];
  assign _zz_1309_ = _zz_1268_[40];
  assign _zz_1310_ = _zz_1268_[41];
  assign _zz_1311_ = _zz_1268_[42];
  assign _zz_1312_ = _zz_1268_[43];
  assign _zz_1313_ = _zz_1268_[44];
  assign _zz_1314_ = _zz_1268_[45];
  assign _zz_1315_ = _zz_1268_[46];
  assign _zz_1316_ = _zz_1268_[47];
  assign _zz_1317_ = _zz_1268_[48];
  assign _zz_1318_ = _zz_1268_[49];
  assign _zz_1319_ = (((32'h000005aa <= load_data_area_current_addr) && (load_data_area_current_addr < 32'h000005dc)) ? axi4_w_payload_data_regNext : {_zz_2799_,_zz_2800_});
  assign _zz_1320_ = _zz_1319_[15 : 0];
  assign _zz_1321_ = _zz_1319_[31 : 16];
  assign _zz_1322_ = _zz_2881_[5:0];
  assign _zz_1323_ = ({63'd0,(1'b1)} <<< _zz_1322_);
  assign _zz_1324_ = _zz_1323_[0];
  assign _zz_1325_ = _zz_1323_[1];
  assign _zz_1326_ = _zz_1323_[2];
  assign _zz_1327_ = _zz_1323_[3];
  assign _zz_1328_ = _zz_1323_[4];
  assign _zz_1329_ = _zz_1323_[5];
  assign _zz_1330_ = _zz_1323_[6];
  assign _zz_1331_ = _zz_1323_[7];
  assign _zz_1332_ = _zz_1323_[8];
  assign _zz_1333_ = _zz_1323_[9];
  assign _zz_1334_ = _zz_1323_[10];
  assign _zz_1335_ = _zz_1323_[11];
  assign _zz_1336_ = _zz_1323_[12];
  assign _zz_1337_ = _zz_1323_[13];
  assign _zz_1338_ = _zz_1323_[14];
  assign _zz_1339_ = _zz_1323_[15];
  assign _zz_1340_ = _zz_1323_[16];
  assign _zz_1341_ = _zz_1323_[17];
  assign _zz_1342_ = _zz_1323_[18];
  assign _zz_1343_ = _zz_1323_[19];
  assign _zz_1344_ = _zz_1323_[20];
  assign _zz_1345_ = _zz_1323_[21];
  assign _zz_1346_ = _zz_1323_[22];
  assign _zz_1347_ = _zz_1323_[23];
  assign _zz_1348_ = _zz_1323_[24];
  assign _zz_1349_ = _zz_1323_[25];
  assign _zz_1350_ = _zz_1323_[26];
  assign _zz_1351_ = _zz_1323_[27];
  assign _zz_1352_ = _zz_1323_[28];
  assign _zz_1353_ = _zz_1323_[29];
  assign _zz_1354_ = _zz_1323_[30];
  assign _zz_1355_ = _zz_1323_[31];
  assign _zz_1356_ = _zz_1323_[32];
  assign _zz_1357_ = _zz_1323_[33];
  assign _zz_1358_ = _zz_1323_[34];
  assign _zz_1359_ = _zz_1323_[35];
  assign _zz_1360_ = _zz_1323_[36];
  assign _zz_1361_ = _zz_1323_[37];
  assign _zz_1362_ = _zz_1323_[38];
  assign _zz_1363_ = _zz_1323_[39];
  assign _zz_1364_ = _zz_1323_[40];
  assign _zz_1365_ = _zz_1323_[41];
  assign _zz_1366_ = _zz_1323_[42];
  assign _zz_1367_ = _zz_1323_[43];
  assign _zz_1368_ = _zz_1323_[44];
  assign _zz_1369_ = _zz_1323_[45];
  assign _zz_1370_ = _zz_1323_[46];
  assign _zz_1371_ = _zz_1323_[47];
  assign _zz_1372_ = _zz_1323_[48];
  assign _zz_1373_ = _zz_1323_[49];
  assign _zz_1374_ = (((32'h00000802 <= load_data_area_current_addr) && (load_data_area_current_addr < 32'h00000834)) ? axi4_w_payload_data_regNext : {_zz_2801_,_zz_2802_});
  assign _zz_1375_ = _zz_1374_[15 : 0];
  assign _zz_1376_ = _zz_1374_[31 : 16];
  assign _zz_1377_ = _zz_2882_[5:0];
  assign _zz_1378_ = ({63'd0,(1'b1)} <<< _zz_1377_);
  assign _zz_1379_ = _zz_1378_[0];
  assign _zz_1380_ = _zz_1378_[1];
  assign _zz_1381_ = _zz_1378_[2];
  assign _zz_1382_ = _zz_1378_[3];
  assign _zz_1383_ = _zz_1378_[4];
  assign _zz_1384_ = _zz_1378_[5];
  assign _zz_1385_ = _zz_1378_[6];
  assign _zz_1386_ = _zz_1378_[7];
  assign _zz_1387_ = _zz_1378_[8];
  assign _zz_1388_ = _zz_1378_[9];
  assign _zz_1389_ = _zz_1378_[10];
  assign _zz_1390_ = _zz_1378_[11];
  assign _zz_1391_ = _zz_1378_[12];
  assign _zz_1392_ = _zz_1378_[13];
  assign _zz_1393_ = _zz_1378_[14];
  assign _zz_1394_ = _zz_1378_[15];
  assign _zz_1395_ = _zz_1378_[16];
  assign _zz_1396_ = _zz_1378_[17];
  assign _zz_1397_ = _zz_1378_[18];
  assign _zz_1398_ = _zz_1378_[19];
  assign _zz_1399_ = _zz_1378_[20];
  assign _zz_1400_ = _zz_1378_[21];
  assign _zz_1401_ = _zz_1378_[22];
  assign _zz_1402_ = _zz_1378_[23];
  assign _zz_1403_ = _zz_1378_[24];
  assign _zz_1404_ = _zz_1378_[25];
  assign _zz_1405_ = _zz_1378_[26];
  assign _zz_1406_ = _zz_1378_[27];
  assign _zz_1407_ = _zz_1378_[28];
  assign _zz_1408_ = _zz_1378_[29];
  assign _zz_1409_ = _zz_1378_[30];
  assign _zz_1410_ = _zz_1378_[31];
  assign _zz_1411_ = _zz_1378_[32];
  assign _zz_1412_ = _zz_1378_[33];
  assign _zz_1413_ = _zz_1378_[34];
  assign _zz_1414_ = _zz_1378_[35];
  assign _zz_1415_ = _zz_1378_[36];
  assign _zz_1416_ = _zz_1378_[37];
  assign _zz_1417_ = _zz_1378_[38];
  assign _zz_1418_ = _zz_1378_[39];
  assign _zz_1419_ = _zz_1378_[40];
  assign _zz_1420_ = _zz_1378_[41];
  assign _zz_1421_ = _zz_1378_[42];
  assign _zz_1422_ = _zz_1378_[43];
  assign _zz_1423_ = _zz_1378_[44];
  assign _zz_1424_ = _zz_1378_[45];
  assign _zz_1425_ = _zz_1378_[46];
  assign _zz_1426_ = _zz_1378_[47];
  assign _zz_1427_ = _zz_1378_[48];
  assign _zz_1428_ = _zz_1378_[49];
  assign _zz_1429_ = (((32'h0000076c <= load_data_area_current_addr) && (load_data_area_current_addr < 32'h0000079e)) ? axi4_w_payload_data_regNext : {_zz_2803_,_zz_2804_});
  assign _zz_1430_ = _zz_1429_[15 : 0];
  assign _zz_1431_ = _zz_1429_[31 : 16];
  assign _zz_1432_ = _zz_2883_[5:0];
  assign _zz_1433_ = ({63'd0,(1'b1)} <<< _zz_1432_);
  assign _zz_1434_ = _zz_1433_[0];
  assign _zz_1435_ = _zz_1433_[1];
  assign _zz_1436_ = _zz_1433_[2];
  assign _zz_1437_ = _zz_1433_[3];
  assign _zz_1438_ = _zz_1433_[4];
  assign _zz_1439_ = _zz_1433_[5];
  assign _zz_1440_ = _zz_1433_[6];
  assign _zz_1441_ = _zz_1433_[7];
  assign _zz_1442_ = _zz_1433_[8];
  assign _zz_1443_ = _zz_1433_[9];
  assign _zz_1444_ = _zz_1433_[10];
  assign _zz_1445_ = _zz_1433_[11];
  assign _zz_1446_ = _zz_1433_[12];
  assign _zz_1447_ = _zz_1433_[13];
  assign _zz_1448_ = _zz_1433_[14];
  assign _zz_1449_ = _zz_1433_[15];
  assign _zz_1450_ = _zz_1433_[16];
  assign _zz_1451_ = _zz_1433_[17];
  assign _zz_1452_ = _zz_1433_[18];
  assign _zz_1453_ = _zz_1433_[19];
  assign _zz_1454_ = _zz_1433_[20];
  assign _zz_1455_ = _zz_1433_[21];
  assign _zz_1456_ = _zz_1433_[22];
  assign _zz_1457_ = _zz_1433_[23];
  assign _zz_1458_ = _zz_1433_[24];
  assign _zz_1459_ = _zz_1433_[25];
  assign _zz_1460_ = _zz_1433_[26];
  assign _zz_1461_ = _zz_1433_[27];
  assign _zz_1462_ = _zz_1433_[28];
  assign _zz_1463_ = _zz_1433_[29];
  assign _zz_1464_ = _zz_1433_[30];
  assign _zz_1465_ = _zz_1433_[31];
  assign _zz_1466_ = _zz_1433_[32];
  assign _zz_1467_ = _zz_1433_[33];
  assign _zz_1468_ = _zz_1433_[34];
  assign _zz_1469_ = _zz_1433_[35];
  assign _zz_1470_ = _zz_1433_[36];
  assign _zz_1471_ = _zz_1433_[37];
  assign _zz_1472_ = _zz_1433_[38];
  assign _zz_1473_ = _zz_1433_[39];
  assign _zz_1474_ = _zz_1433_[40];
  assign _zz_1475_ = _zz_1433_[41];
  assign _zz_1476_ = _zz_1433_[42];
  assign _zz_1477_ = _zz_1433_[43];
  assign _zz_1478_ = _zz_1433_[44];
  assign _zz_1479_ = _zz_1433_[45];
  assign _zz_1480_ = _zz_1433_[46];
  assign _zz_1481_ = _zz_1433_[47];
  assign _zz_1482_ = _zz_1433_[48];
  assign _zz_1483_ = _zz_1433_[49];
  assign _zz_1484_ = (((32'h00000096 <= load_data_area_current_addr) && (load_data_area_current_addr < 32'h000000c8)) ? axi4_w_payload_data_regNext : {_zz_2805_,_zz_2806_});
  assign _zz_1485_ = _zz_1484_[15 : 0];
  assign _zz_1486_ = _zz_1484_[31 : 16];
  assign _zz_1487_ = _zz_2884_[5:0];
  assign _zz_1488_ = ({63'd0,(1'b1)} <<< _zz_1487_);
  assign _zz_1489_ = _zz_1488_[0];
  assign _zz_1490_ = _zz_1488_[1];
  assign _zz_1491_ = _zz_1488_[2];
  assign _zz_1492_ = _zz_1488_[3];
  assign _zz_1493_ = _zz_1488_[4];
  assign _zz_1494_ = _zz_1488_[5];
  assign _zz_1495_ = _zz_1488_[6];
  assign _zz_1496_ = _zz_1488_[7];
  assign _zz_1497_ = _zz_1488_[8];
  assign _zz_1498_ = _zz_1488_[9];
  assign _zz_1499_ = _zz_1488_[10];
  assign _zz_1500_ = _zz_1488_[11];
  assign _zz_1501_ = _zz_1488_[12];
  assign _zz_1502_ = _zz_1488_[13];
  assign _zz_1503_ = _zz_1488_[14];
  assign _zz_1504_ = _zz_1488_[15];
  assign _zz_1505_ = _zz_1488_[16];
  assign _zz_1506_ = _zz_1488_[17];
  assign _zz_1507_ = _zz_1488_[18];
  assign _zz_1508_ = _zz_1488_[19];
  assign _zz_1509_ = _zz_1488_[20];
  assign _zz_1510_ = _zz_1488_[21];
  assign _zz_1511_ = _zz_1488_[22];
  assign _zz_1512_ = _zz_1488_[23];
  assign _zz_1513_ = _zz_1488_[24];
  assign _zz_1514_ = _zz_1488_[25];
  assign _zz_1515_ = _zz_1488_[26];
  assign _zz_1516_ = _zz_1488_[27];
  assign _zz_1517_ = _zz_1488_[28];
  assign _zz_1518_ = _zz_1488_[29];
  assign _zz_1519_ = _zz_1488_[30];
  assign _zz_1520_ = _zz_1488_[31];
  assign _zz_1521_ = _zz_1488_[32];
  assign _zz_1522_ = _zz_1488_[33];
  assign _zz_1523_ = _zz_1488_[34];
  assign _zz_1524_ = _zz_1488_[35];
  assign _zz_1525_ = _zz_1488_[36];
  assign _zz_1526_ = _zz_1488_[37];
  assign _zz_1527_ = _zz_1488_[38];
  assign _zz_1528_ = _zz_1488_[39];
  assign _zz_1529_ = _zz_1488_[40];
  assign _zz_1530_ = _zz_1488_[41];
  assign _zz_1531_ = _zz_1488_[42];
  assign _zz_1532_ = _zz_1488_[43];
  assign _zz_1533_ = _zz_1488_[44];
  assign _zz_1534_ = _zz_1488_[45];
  assign _zz_1535_ = _zz_1488_[46];
  assign _zz_1536_ = _zz_1488_[47];
  assign _zz_1537_ = _zz_1488_[48];
  assign _zz_1538_ = _zz_1488_[49];
  assign _zz_1539_ = (((32'h000006a4 <= load_data_area_current_addr) && (load_data_area_current_addr < 32'h000006d6)) ? axi4_w_payload_data_regNext : {_zz_2807_,_zz_2808_});
  assign _zz_1540_ = _zz_1539_[15 : 0];
  assign _zz_1541_ = _zz_1539_[31 : 16];
  assign _zz_1542_ = _zz_2885_[5:0];
  assign _zz_1543_ = ({63'd0,(1'b1)} <<< _zz_1542_);
  assign _zz_1544_ = _zz_1543_[0];
  assign _zz_1545_ = _zz_1543_[1];
  assign _zz_1546_ = _zz_1543_[2];
  assign _zz_1547_ = _zz_1543_[3];
  assign _zz_1548_ = _zz_1543_[4];
  assign _zz_1549_ = _zz_1543_[5];
  assign _zz_1550_ = _zz_1543_[6];
  assign _zz_1551_ = _zz_1543_[7];
  assign _zz_1552_ = _zz_1543_[8];
  assign _zz_1553_ = _zz_1543_[9];
  assign _zz_1554_ = _zz_1543_[10];
  assign _zz_1555_ = _zz_1543_[11];
  assign _zz_1556_ = _zz_1543_[12];
  assign _zz_1557_ = _zz_1543_[13];
  assign _zz_1558_ = _zz_1543_[14];
  assign _zz_1559_ = _zz_1543_[15];
  assign _zz_1560_ = _zz_1543_[16];
  assign _zz_1561_ = _zz_1543_[17];
  assign _zz_1562_ = _zz_1543_[18];
  assign _zz_1563_ = _zz_1543_[19];
  assign _zz_1564_ = _zz_1543_[20];
  assign _zz_1565_ = _zz_1543_[21];
  assign _zz_1566_ = _zz_1543_[22];
  assign _zz_1567_ = _zz_1543_[23];
  assign _zz_1568_ = _zz_1543_[24];
  assign _zz_1569_ = _zz_1543_[25];
  assign _zz_1570_ = _zz_1543_[26];
  assign _zz_1571_ = _zz_1543_[27];
  assign _zz_1572_ = _zz_1543_[28];
  assign _zz_1573_ = _zz_1543_[29];
  assign _zz_1574_ = _zz_1543_[30];
  assign _zz_1575_ = _zz_1543_[31];
  assign _zz_1576_ = _zz_1543_[32];
  assign _zz_1577_ = _zz_1543_[33];
  assign _zz_1578_ = _zz_1543_[34];
  assign _zz_1579_ = _zz_1543_[35];
  assign _zz_1580_ = _zz_1543_[36];
  assign _zz_1581_ = _zz_1543_[37];
  assign _zz_1582_ = _zz_1543_[38];
  assign _zz_1583_ = _zz_1543_[39];
  assign _zz_1584_ = _zz_1543_[40];
  assign _zz_1585_ = _zz_1543_[41];
  assign _zz_1586_ = _zz_1543_[42];
  assign _zz_1587_ = _zz_1543_[43];
  assign _zz_1588_ = _zz_1543_[44];
  assign _zz_1589_ = _zz_1543_[45];
  assign _zz_1590_ = _zz_1543_[46];
  assign _zz_1591_ = _zz_1543_[47];
  assign _zz_1592_ = _zz_1543_[48];
  assign _zz_1593_ = _zz_1543_[49];
  assign _zz_1594_ = (((32'h0000015e <= load_data_area_current_addr) && (load_data_area_current_addr < 32'h00000190)) ? axi4_w_payload_data_regNext : {_zz_2809_,_zz_2810_});
  assign _zz_1595_ = _zz_1594_[15 : 0];
  assign _zz_1596_ = _zz_1594_[31 : 16];
  assign _zz_1597_ = _zz_2886_[5:0];
  assign _zz_1598_ = ({63'd0,(1'b1)} <<< _zz_1597_);
  assign _zz_1599_ = _zz_1598_[0];
  assign _zz_1600_ = _zz_1598_[1];
  assign _zz_1601_ = _zz_1598_[2];
  assign _zz_1602_ = _zz_1598_[3];
  assign _zz_1603_ = _zz_1598_[4];
  assign _zz_1604_ = _zz_1598_[5];
  assign _zz_1605_ = _zz_1598_[6];
  assign _zz_1606_ = _zz_1598_[7];
  assign _zz_1607_ = _zz_1598_[8];
  assign _zz_1608_ = _zz_1598_[9];
  assign _zz_1609_ = _zz_1598_[10];
  assign _zz_1610_ = _zz_1598_[11];
  assign _zz_1611_ = _zz_1598_[12];
  assign _zz_1612_ = _zz_1598_[13];
  assign _zz_1613_ = _zz_1598_[14];
  assign _zz_1614_ = _zz_1598_[15];
  assign _zz_1615_ = _zz_1598_[16];
  assign _zz_1616_ = _zz_1598_[17];
  assign _zz_1617_ = _zz_1598_[18];
  assign _zz_1618_ = _zz_1598_[19];
  assign _zz_1619_ = _zz_1598_[20];
  assign _zz_1620_ = _zz_1598_[21];
  assign _zz_1621_ = _zz_1598_[22];
  assign _zz_1622_ = _zz_1598_[23];
  assign _zz_1623_ = _zz_1598_[24];
  assign _zz_1624_ = _zz_1598_[25];
  assign _zz_1625_ = _zz_1598_[26];
  assign _zz_1626_ = _zz_1598_[27];
  assign _zz_1627_ = _zz_1598_[28];
  assign _zz_1628_ = _zz_1598_[29];
  assign _zz_1629_ = _zz_1598_[30];
  assign _zz_1630_ = _zz_1598_[31];
  assign _zz_1631_ = _zz_1598_[32];
  assign _zz_1632_ = _zz_1598_[33];
  assign _zz_1633_ = _zz_1598_[34];
  assign _zz_1634_ = _zz_1598_[35];
  assign _zz_1635_ = _zz_1598_[36];
  assign _zz_1636_ = _zz_1598_[37];
  assign _zz_1637_ = _zz_1598_[38];
  assign _zz_1638_ = _zz_1598_[39];
  assign _zz_1639_ = _zz_1598_[40];
  assign _zz_1640_ = _zz_1598_[41];
  assign _zz_1641_ = _zz_1598_[42];
  assign _zz_1642_ = _zz_1598_[43];
  assign _zz_1643_ = _zz_1598_[44];
  assign _zz_1644_ = _zz_1598_[45];
  assign _zz_1645_ = _zz_1598_[46];
  assign _zz_1646_ = _zz_1598_[47];
  assign _zz_1647_ = _zz_1598_[48];
  assign _zz_1648_ = _zz_1598_[49];
  assign _zz_1649_ = (((32'h000001c2 <= load_data_area_current_addr) && (load_data_area_current_addr < 32'h000001f4)) ? axi4_w_payload_data_regNext : {_zz_2811_,_zz_2812_});
  assign _zz_1650_ = _zz_1649_[15 : 0];
  assign _zz_1651_ = _zz_1649_[31 : 16];
  assign _zz_1652_ = _zz_2887_[5:0];
  assign _zz_1653_ = ({63'd0,(1'b1)} <<< _zz_1652_);
  assign _zz_1654_ = _zz_1653_[0];
  assign _zz_1655_ = _zz_1653_[1];
  assign _zz_1656_ = _zz_1653_[2];
  assign _zz_1657_ = _zz_1653_[3];
  assign _zz_1658_ = _zz_1653_[4];
  assign _zz_1659_ = _zz_1653_[5];
  assign _zz_1660_ = _zz_1653_[6];
  assign _zz_1661_ = _zz_1653_[7];
  assign _zz_1662_ = _zz_1653_[8];
  assign _zz_1663_ = _zz_1653_[9];
  assign _zz_1664_ = _zz_1653_[10];
  assign _zz_1665_ = _zz_1653_[11];
  assign _zz_1666_ = _zz_1653_[12];
  assign _zz_1667_ = _zz_1653_[13];
  assign _zz_1668_ = _zz_1653_[14];
  assign _zz_1669_ = _zz_1653_[15];
  assign _zz_1670_ = _zz_1653_[16];
  assign _zz_1671_ = _zz_1653_[17];
  assign _zz_1672_ = _zz_1653_[18];
  assign _zz_1673_ = _zz_1653_[19];
  assign _zz_1674_ = _zz_1653_[20];
  assign _zz_1675_ = _zz_1653_[21];
  assign _zz_1676_ = _zz_1653_[22];
  assign _zz_1677_ = _zz_1653_[23];
  assign _zz_1678_ = _zz_1653_[24];
  assign _zz_1679_ = _zz_1653_[25];
  assign _zz_1680_ = _zz_1653_[26];
  assign _zz_1681_ = _zz_1653_[27];
  assign _zz_1682_ = _zz_1653_[28];
  assign _zz_1683_ = _zz_1653_[29];
  assign _zz_1684_ = _zz_1653_[30];
  assign _zz_1685_ = _zz_1653_[31];
  assign _zz_1686_ = _zz_1653_[32];
  assign _zz_1687_ = _zz_1653_[33];
  assign _zz_1688_ = _zz_1653_[34];
  assign _zz_1689_ = _zz_1653_[35];
  assign _zz_1690_ = _zz_1653_[36];
  assign _zz_1691_ = _zz_1653_[37];
  assign _zz_1692_ = _zz_1653_[38];
  assign _zz_1693_ = _zz_1653_[39];
  assign _zz_1694_ = _zz_1653_[40];
  assign _zz_1695_ = _zz_1653_[41];
  assign _zz_1696_ = _zz_1653_[42];
  assign _zz_1697_ = _zz_1653_[43];
  assign _zz_1698_ = _zz_1653_[44];
  assign _zz_1699_ = _zz_1653_[45];
  assign _zz_1700_ = _zz_1653_[46];
  assign _zz_1701_ = _zz_1653_[47];
  assign _zz_1702_ = _zz_1653_[48];
  assign _zz_1703_ = _zz_1653_[49];
  assign _zz_1704_ = (((32'h00000190 <= load_data_area_current_addr) && (load_data_area_current_addr < 32'h000001c2)) ? axi4_w_payload_data_regNext : {_zz_2813_,_zz_2814_});
  assign _zz_1705_ = _zz_1704_[15 : 0];
  assign _zz_1706_ = _zz_1704_[31 : 16];
  assign _zz_1707_ = _zz_2888_[5:0];
  assign _zz_1708_ = ({63'd0,(1'b1)} <<< _zz_1707_);
  assign _zz_1709_ = _zz_1708_[0];
  assign _zz_1710_ = _zz_1708_[1];
  assign _zz_1711_ = _zz_1708_[2];
  assign _zz_1712_ = _zz_1708_[3];
  assign _zz_1713_ = _zz_1708_[4];
  assign _zz_1714_ = _zz_1708_[5];
  assign _zz_1715_ = _zz_1708_[6];
  assign _zz_1716_ = _zz_1708_[7];
  assign _zz_1717_ = _zz_1708_[8];
  assign _zz_1718_ = _zz_1708_[9];
  assign _zz_1719_ = _zz_1708_[10];
  assign _zz_1720_ = _zz_1708_[11];
  assign _zz_1721_ = _zz_1708_[12];
  assign _zz_1722_ = _zz_1708_[13];
  assign _zz_1723_ = _zz_1708_[14];
  assign _zz_1724_ = _zz_1708_[15];
  assign _zz_1725_ = _zz_1708_[16];
  assign _zz_1726_ = _zz_1708_[17];
  assign _zz_1727_ = _zz_1708_[18];
  assign _zz_1728_ = _zz_1708_[19];
  assign _zz_1729_ = _zz_1708_[20];
  assign _zz_1730_ = _zz_1708_[21];
  assign _zz_1731_ = _zz_1708_[22];
  assign _zz_1732_ = _zz_1708_[23];
  assign _zz_1733_ = _zz_1708_[24];
  assign _zz_1734_ = _zz_1708_[25];
  assign _zz_1735_ = _zz_1708_[26];
  assign _zz_1736_ = _zz_1708_[27];
  assign _zz_1737_ = _zz_1708_[28];
  assign _zz_1738_ = _zz_1708_[29];
  assign _zz_1739_ = _zz_1708_[30];
  assign _zz_1740_ = _zz_1708_[31];
  assign _zz_1741_ = _zz_1708_[32];
  assign _zz_1742_ = _zz_1708_[33];
  assign _zz_1743_ = _zz_1708_[34];
  assign _zz_1744_ = _zz_1708_[35];
  assign _zz_1745_ = _zz_1708_[36];
  assign _zz_1746_ = _zz_1708_[37];
  assign _zz_1747_ = _zz_1708_[38];
  assign _zz_1748_ = _zz_1708_[39];
  assign _zz_1749_ = _zz_1708_[40];
  assign _zz_1750_ = _zz_1708_[41];
  assign _zz_1751_ = _zz_1708_[42];
  assign _zz_1752_ = _zz_1708_[43];
  assign _zz_1753_ = _zz_1708_[44];
  assign _zz_1754_ = _zz_1708_[45];
  assign _zz_1755_ = _zz_1708_[46];
  assign _zz_1756_ = _zz_1708_[47];
  assign _zz_1757_ = _zz_1708_[48];
  assign _zz_1758_ = _zz_1708_[49];
  assign _zz_1759_ = (((32'h00000384 <= load_data_area_current_addr) && (load_data_area_current_addr < 32'h000003b6)) ? axi4_w_payload_data_regNext : {_zz_2815_,_zz_2816_});
  assign _zz_1760_ = _zz_1759_[15 : 0];
  assign _zz_1761_ = _zz_1759_[31 : 16];
  assign _zz_1762_ = _zz_2889_[5:0];
  assign _zz_1763_ = ({63'd0,(1'b1)} <<< _zz_1762_);
  assign _zz_1764_ = _zz_1763_[0];
  assign _zz_1765_ = _zz_1763_[1];
  assign _zz_1766_ = _zz_1763_[2];
  assign _zz_1767_ = _zz_1763_[3];
  assign _zz_1768_ = _zz_1763_[4];
  assign _zz_1769_ = _zz_1763_[5];
  assign _zz_1770_ = _zz_1763_[6];
  assign _zz_1771_ = _zz_1763_[7];
  assign _zz_1772_ = _zz_1763_[8];
  assign _zz_1773_ = _zz_1763_[9];
  assign _zz_1774_ = _zz_1763_[10];
  assign _zz_1775_ = _zz_1763_[11];
  assign _zz_1776_ = _zz_1763_[12];
  assign _zz_1777_ = _zz_1763_[13];
  assign _zz_1778_ = _zz_1763_[14];
  assign _zz_1779_ = _zz_1763_[15];
  assign _zz_1780_ = _zz_1763_[16];
  assign _zz_1781_ = _zz_1763_[17];
  assign _zz_1782_ = _zz_1763_[18];
  assign _zz_1783_ = _zz_1763_[19];
  assign _zz_1784_ = _zz_1763_[20];
  assign _zz_1785_ = _zz_1763_[21];
  assign _zz_1786_ = _zz_1763_[22];
  assign _zz_1787_ = _zz_1763_[23];
  assign _zz_1788_ = _zz_1763_[24];
  assign _zz_1789_ = _zz_1763_[25];
  assign _zz_1790_ = _zz_1763_[26];
  assign _zz_1791_ = _zz_1763_[27];
  assign _zz_1792_ = _zz_1763_[28];
  assign _zz_1793_ = _zz_1763_[29];
  assign _zz_1794_ = _zz_1763_[30];
  assign _zz_1795_ = _zz_1763_[31];
  assign _zz_1796_ = _zz_1763_[32];
  assign _zz_1797_ = _zz_1763_[33];
  assign _zz_1798_ = _zz_1763_[34];
  assign _zz_1799_ = _zz_1763_[35];
  assign _zz_1800_ = _zz_1763_[36];
  assign _zz_1801_ = _zz_1763_[37];
  assign _zz_1802_ = _zz_1763_[38];
  assign _zz_1803_ = _zz_1763_[39];
  assign _zz_1804_ = _zz_1763_[40];
  assign _zz_1805_ = _zz_1763_[41];
  assign _zz_1806_ = _zz_1763_[42];
  assign _zz_1807_ = _zz_1763_[43];
  assign _zz_1808_ = _zz_1763_[44];
  assign _zz_1809_ = _zz_1763_[45];
  assign _zz_1810_ = _zz_1763_[46];
  assign _zz_1811_ = _zz_1763_[47];
  assign _zz_1812_ = _zz_1763_[48];
  assign _zz_1813_ = _zz_1763_[49];
  assign _zz_1814_ = (((32'h00000866 <= load_data_area_current_addr) && (load_data_area_current_addr < 32'h00000898)) ? axi4_w_payload_data_regNext : {_zz_2817_,_zz_2818_});
  assign _zz_1815_ = _zz_1814_[15 : 0];
  assign _zz_1816_ = _zz_1814_[31 : 16];
  assign _zz_1817_ = _zz_2890_[5:0];
  assign _zz_1818_ = ({63'd0,(1'b1)} <<< _zz_1817_);
  assign _zz_1819_ = _zz_1818_[0];
  assign _zz_1820_ = _zz_1818_[1];
  assign _zz_1821_ = _zz_1818_[2];
  assign _zz_1822_ = _zz_1818_[3];
  assign _zz_1823_ = _zz_1818_[4];
  assign _zz_1824_ = _zz_1818_[5];
  assign _zz_1825_ = _zz_1818_[6];
  assign _zz_1826_ = _zz_1818_[7];
  assign _zz_1827_ = _zz_1818_[8];
  assign _zz_1828_ = _zz_1818_[9];
  assign _zz_1829_ = _zz_1818_[10];
  assign _zz_1830_ = _zz_1818_[11];
  assign _zz_1831_ = _zz_1818_[12];
  assign _zz_1832_ = _zz_1818_[13];
  assign _zz_1833_ = _zz_1818_[14];
  assign _zz_1834_ = _zz_1818_[15];
  assign _zz_1835_ = _zz_1818_[16];
  assign _zz_1836_ = _zz_1818_[17];
  assign _zz_1837_ = _zz_1818_[18];
  assign _zz_1838_ = _zz_1818_[19];
  assign _zz_1839_ = _zz_1818_[20];
  assign _zz_1840_ = _zz_1818_[21];
  assign _zz_1841_ = _zz_1818_[22];
  assign _zz_1842_ = _zz_1818_[23];
  assign _zz_1843_ = _zz_1818_[24];
  assign _zz_1844_ = _zz_1818_[25];
  assign _zz_1845_ = _zz_1818_[26];
  assign _zz_1846_ = _zz_1818_[27];
  assign _zz_1847_ = _zz_1818_[28];
  assign _zz_1848_ = _zz_1818_[29];
  assign _zz_1849_ = _zz_1818_[30];
  assign _zz_1850_ = _zz_1818_[31];
  assign _zz_1851_ = _zz_1818_[32];
  assign _zz_1852_ = _zz_1818_[33];
  assign _zz_1853_ = _zz_1818_[34];
  assign _zz_1854_ = _zz_1818_[35];
  assign _zz_1855_ = _zz_1818_[36];
  assign _zz_1856_ = _zz_1818_[37];
  assign _zz_1857_ = _zz_1818_[38];
  assign _zz_1858_ = _zz_1818_[39];
  assign _zz_1859_ = _zz_1818_[40];
  assign _zz_1860_ = _zz_1818_[41];
  assign _zz_1861_ = _zz_1818_[42];
  assign _zz_1862_ = _zz_1818_[43];
  assign _zz_1863_ = _zz_1818_[44];
  assign _zz_1864_ = _zz_1818_[45];
  assign _zz_1865_ = _zz_1818_[46];
  assign _zz_1866_ = _zz_1818_[47];
  assign _zz_1867_ = _zz_1818_[48];
  assign _zz_1868_ = _zz_1818_[49];
  assign _zz_1869_ = (((32'h00000960 <= load_data_area_current_addr) && (load_data_area_current_addr < 32'h00000992)) ? axi4_w_payload_data_regNext : {_zz_2819_,_zz_2820_});
  assign _zz_1870_ = _zz_1869_[15 : 0];
  assign _zz_1871_ = _zz_1869_[31 : 16];
  assign _zz_1872_ = _zz_2891_[5:0];
  assign _zz_1873_ = ({63'd0,(1'b1)} <<< _zz_1872_);
  assign _zz_1874_ = _zz_1873_[0];
  assign _zz_1875_ = _zz_1873_[1];
  assign _zz_1876_ = _zz_1873_[2];
  assign _zz_1877_ = _zz_1873_[3];
  assign _zz_1878_ = _zz_1873_[4];
  assign _zz_1879_ = _zz_1873_[5];
  assign _zz_1880_ = _zz_1873_[6];
  assign _zz_1881_ = _zz_1873_[7];
  assign _zz_1882_ = _zz_1873_[8];
  assign _zz_1883_ = _zz_1873_[9];
  assign _zz_1884_ = _zz_1873_[10];
  assign _zz_1885_ = _zz_1873_[11];
  assign _zz_1886_ = _zz_1873_[12];
  assign _zz_1887_ = _zz_1873_[13];
  assign _zz_1888_ = _zz_1873_[14];
  assign _zz_1889_ = _zz_1873_[15];
  assign _zz_1890_ = _zz_1873_[16];
  assign _zz_1891_ = _zz_1873_[17];
  assign _zz_1892_ = _zz_1873_[18];
  assign _zz_1893_ = _zz_1873_[19];
  assign _zz_1894_ = _zz_1873_[20];
  assign _zz_1895_ = _zz_1873_[21];
  assign _zz_1896_ = _zz_1873_[22];
  assign _zz_1897_ = _zz_1873_[23];
  assign _zz_1898_ = _zz_1873_[24];
  assign _zz_1899_ = _zz_1873_[25];
  assign _zz_1900_ = _zz_1873_[26];
  assign _zz_1901_ = _zz_1873_[27];
  assign _zz_1902_ = _zz_1873_[28];
  assign _zz_1903_ = _zz_1873_[29];
  assign _zz_1904_ = _zz_1873_[30];
  assign _zz_1905_ = _zz_1873_[31];
  assign _zz_1906_ = _zz_1873_[32];
  assign _zz_1907_ = _zz_1873_[33];
  assign _zz_1908_ = _zz_1873_[34];
  assign _zz_1909_ = _zz_1873_[35];
  assign _zz_1910_ = _zz_1873_[36];
  assign _zz_1911_ = _zz_1873_[37];
  assign _zz_1912_ = _zz_1873_[38];
  assign _zz_1913_ = _zz_1873_[39];
  assign _zz_1914_ = _zz_1873_[40];
  assign _zz_1915_ = _zz_1873_[41];
  assign _zz_1916_ = _zz_1873_[42];
  assign _zz_1917_ = _zz_1873_[43];
  assign _zz_1918_ = _zz_1873_[44];
  assign _zz_1919_ = _zz_1873_[45];
  assign _zz_1920_ = _zz_1873_[46];
  assign _zz_1921_ = _zz_1873_[47];
  assign _zz_1922_ = _zz_1873_[48];
  assign _zz_1923_ = _zz_1873_[49];
  assign _zz_1924_ = (((32'h00000578 <= load_data_area_current_addr) && (load_data_area_current_addr < 32'h000005aa)) ? axi4_w_payload_data_regNext : {_zz_2821_,_zz_2822_});
  assign _zz_1925_ = _zz_1924_[15 : 0];
  assign _zz_1926_ = _zz_1924_[31 : 16];
  assign _zz_1927_ = _zz_2892_[5:0];
  assign _zz_1928_ = ({63'd0,(1'b1)} <<< _zz_1927_);
  assign _zz_1929_ = _zz_1928_[0];
  assign _zz_1930_ = _zz_1928_[1];
  assign _zz_1931_ = _zz_1928_[2];
  assign _zz_1932_ = _zz_1928_[3];
  assign _zz_1933_ = _zz_1928_[4];
  assign _zz_1934_ = _zz_1928_[5];
  assign _zz_1935_ = _zz_1928_[6];
  assign _zz_1936_ = _zz_1928_[7];
  assign _zz_1937_ = _zz_1928_[8];
  assign _zz_1938_ = _zz_1928_[9];
  assign _zz_1939_ = _zz_1928_[10];
  assign _zz_1940_ = _zz_1928_[11];
  assign _zz_1941_ = _zz_1928_[12];
  assign _zz_1942_ = _zz_1928_[13];
  assign _zz_1943_ = _zz_1928_[14];
  assign _zz_1944_ = _zz_1928_[15];
  assign _zz_1945_ = _zz_1928_[16];
  assign _zz_1946_ = _zz_1928_[17];
  assign _zz_1947_ = _zz_1928_[18];
  assign _zz_1948_ = _zz_1928_[19];
  assign _zz_1949_ = _zz_1928_[20];
  assign _zz_1950_ = _zz_1928_[21];
  assign _zz_1951_ = _zz_1928_[22];
  assign _zz_1952_ = _zz_1928_[23];
  assign _zz_1953_ = _zz_1928_[24];
  assign _zz_1954_ = _zz_1928_[25];
  assign _zz_1955_ = _zz_1928_[26];
  assign _zz_1956_ = _zz_1928_[27];
  assign _zz_1957_ = _zz_1928_[28];
  assign _zz_1958_ = _zz_1928_[29];
  assign _zz_1959_ = _zz_1928_[30];
  assign _zz_1960_ = _zz_1928_[31];
  assign _zz_1961_ = _zz_1928_[32];
  assign _zz_1962_ = _zz_1928_[33];
  assign _zz_1963_ = _zz_1928_[34];
  assign _zz_1964_ = _zz_1928_[35];
  assign _zz_1965_ = _zz_1928_[36];
  assign _zz_1966_ = _zz_1928_[37];
  assign _zz_1967_ = _zz_1928_[38];
  assign _zz_1968_ = _zz_1928_[39];
  assign _zz_1969_ = _zz_1928_[40];
  assign _zz_1970_ = _zz_1928_[41];
  assign _zz_1971_ = _zz_1928_[42];
  assign _zz_1972_ = _zz_1928_[43];
  assign _zz_1973_ = _zz_1928_[44];
  assign _zz_1974_ = _zz_1928_[45];
  assign _zz_1975_ = _zz_1928_[46];
  assign _zz_1976_ = _zz_1928_[47];
  assign _zz_1977_ = _zz_1928_[48];
  assign _zz_1978_ = _zz_1928_[49];
  assign _zz_1979_ = (((32'h000006d6 <= load_data_area_current_addr) && (load_data_area_current_addr < 32'h00000708)) ? axi4_w_payload_data_regNext : {_zz_2823_,_zz_2824_});
  assign _zz_1980_ = _zz_1979_[15 : 0];
  assign _zz_1981_ = _zz_1979_[31 : 16];
  assign _zz_1982_ = _zz_2893_[5:0];
  assign _zz_1983_ = ({63'd0,(1'b1)} <<< _zz_1982_);
  assign _zz_1984_ = _zz_1983_[0];
  assign _zz_1985_ = _zz_1983_[1];
  assign _zz_1986_ = _zz_1983_[2];
  assign _zz_1987_ = _zz_1983_[3];
  assign _zz_1988_ = _zz_1983_[4];
  assign _zz_1989_ = _zz_1983_[5];
  assign _zz_1990_ = _zz_1983_[6];
  assign _zz_1991_ = _zz_1983_[7];
  assign _zz_1992_ = _zz_1983_[8];
  assign _zz_1993_ = _zz_1983_[9];
  assign _zz_1994_ = _zz_1983_[10];
  assign _zz_1995_ = _zz_1983_[11];
  assign _zz_1996_ = _zz_1983_[12];
  assign _zz_1997_ = _zz_1983_[13];
  assign _zz_1998_ = _zz_1983_[14];
  assign _zz_1999_ = _zz_1983_[15];
  assign _zz_2000_ = _zz_1983_[16];
  assign _zz_2001_ = _zz_1983_[17];
  assign _zz_2002_ = _zz_1983_[18];
  assign _zz_2003_ = _zz_1983_[19];
  assign _zz_2004_ = _zz_1983_[20];
  assign _zz_2005_ = _zz_1983_[21];
  assign _zz_2006_ = _zz_1983_[22];
  assign _zz_2007_ = _zz_1983_[23];
  assign _zz_2008_ = _zz_1983_[24];
  assign _zz_2009_ = _zz_1983_[25];
  assign _zz_2010_ = _zz_1983_[26];
  assign _zz_2011_ = _zz_1983_[27];
  assign _zz_2012_ = _zz_1983_[28];
  assign _zz_2013_ = _zz_1983_[29];
  assign _zz_2014_ = _zz_1983_[30];
  assign _zz_2015_ = _zz_1983_[31];
  assign _zz_2016_ = _zz_1983_[32];
  assign _zz_2017_ = _zz_1983_[33];
  assign _zz_2018_ = _zz_1983_[34];
  assign _zz_2019_ = _zz_1983_[35];
  assign _zz_2020_ = _zz_1983_[36];
  assign _zz_2021_ = _zz_1983_[37];
  assign _zz_2022_ = _zz_1983_[38];
  assign _zz_2023_ = _zz_1983_[39];
  assign _zz_2024_ = _zz_1983_[40];
  assign _zz_2025_ = _zz_1983_[41];
  assign _zz_2026_ = _zz_1983_[42];
  assign _zz_2027_ = _zz_1983_[43];
  assign _zz_2028_ = _zz_1983_[44];
  assign _zz_2029_ = _zz_1983_[45];
  assign _zz_2030_ = _zz_1983_[46];
  assign _zz_2031_ = _zz_1983_[47];
  assign _zz_2032_ = _zz_1983_[48];
  assign _zz_2033_ = _zz_1983_[49];
  assign _zz_2034_ = (((32'h000000c8 <= load_data_area_current_addr) && (load_data_area_current_addr < 32'h000000fa)) ? axi4_w_payload_data_regNext : {_zz_2825_,_zz_2826_});
  assign _zz_2035_ = _zz_2034_[15 : 0];
  assign _zz_2036_ = _zz_2034_[31 : 16];
  assign _zz_2037_ = _zz_2894_[5:0];
  assign _zz_2038_ = ({63'd0,(1'b1)} <<< _zz_2037_);
  assign _zz_2039_ = _zz_2038_[0];
  assign _zz_2040_ = _zz_2038_[1];
  assign _zz_2041_ = _zz_2038_[2];
  assign _zz_2042_ = _zz_2038_[3];
  assign _zz_2043_ = _zz_2038_[4];
  assign _zz_2044_ = _zz_2038_[5];
  assign _zz_2045_ = _zz_2038_[6];
  assign _zz_2046_ = _zz_2038_[7];
  assign _zz_2047_ = _zz_2038_[8];
  assign _zz_2048_ = _zz_2038_[9];
  assign _zz_2049_ = _zz_2038_[10];
  assign _zz_2050_ = _zz_2038_[11];
  assign _zz_2051_ = _zz_2038_[12];
  assign _zz_2052_ = _zz_2038_[13];
  assign _zz_2053_ = _zz_2038_[14];
  assign _zz_2054_ = _zz_2038_[15];
  assign _zz_2055_ = _zz_2038_[16];
  assign _zz_2056_ = _zz_2038_[17];
  assign _zz_2057_ = _zz_2038_[18];
  assign _zz_2058_ = _zz_2038_[19];
  assign _zz_2059_ = _zz_2038_[20];
  assign _zz_2060_ = _zz_2038_[21];
  assign _zz_2061_ = _zz_2038_[22];
  assign _zz_2062_ = _zz_2038_[23];
  assign _zz_2063_ = _zz_2038_[24];
  assign _zz_2064_ = _zz_2038_[25];
  assign _zz_2065_ = _zz_2038_[26];
  assign _zz_2066_ = _zz_2038_[27];
  assign _zz_2067_ = _zz_2038_[28];
  assign _zz_2068_ = _zz_2038_[29];
  assign _zz_2069_ = _zz_2038_[30];
  assign _zz_2070_ = _zz_2038_[31];
  assign _zz_2071_ = _zz_2038_[32];
  assign _zz_2072_ = _zz_2038_[33];
  assign _zz_2073_ = _zz_2038_[34];
  assign _zz_2074_ = _zz_2038_[35];
  assign _zz_2075_ = _zz_2038_[36];
  assign _zz_2076_ = _zz_2038_[37];
  assign _zz_2077_ = _zz_2038_[38];
  assign _zz_2078_ = _zz_2038_[39];
  assign _zz_2079_ = _zz_2038_[40];
  assign _zz_2080_ = _zz_2038_[41];
  assign _zz_2081_ = _zz_2038_[42];
  assign _zz_2082_ = _zz_2038_[43];
  assign _zz_2083_ = _zz_2038_[44];
  assign _zz_2084_ = _zz_2038_[45];
  assign _zz_2085_ = _zz_2038_[46];
  assign _zz_2086_ = _zz_2038_[47];
  assign _zz_2087_ = _zz_2038_[48];
  assign _zz_2088_ = _zz_2038_[49];
  assign _zz_2089_ = (((32'h00000032 <= load_data_area_current_addr) && (load_data_area_current_addr < 32'h00000064)) ? axi4_w_payload_data_regNext : {_zz_2827_,_zz_2828_});
  assign _zz_2090_ = _zz_2089_[15 : 0];
  assign _zz_2091_ = _zz_2089_[31 : 16];
  assign _zz_2092_ = _zz_2895_[5:0];
  assign _zz_2093_ = ({63'd0,(1'b1)} <<< _zz_2092_);
  assign _zz_2094_ = _zz_2093_[0];
  assign _zz_2095_ = _zz_2093_[1];
  assign _zz_2096_ = _zz_2093_[2];
  assign _zz_2097_ = _zz_2093_[3];
  assign _zz_2098_ = _zz_2093_[4];
  assign _zz_2099_ = _zz_2093_[5];
  assign _zz_2100_ = _zz_2093_[6];
  assign _zz_2101_ = _zz_2093_[7];
  assign _zz_2102_ = _zz_2093_[8];
  assign _zz_2103_ = _zz_2093_[9];
  assign _zz_2104_ = _zz_2093_[10];
  assign _zz_2105_ = _zz_2093_[11];
  assign _zz_2106_ = _zz_2093_[12];
  assign _zz_2107_ = _zz_2093_[13];
  assign _zz_2108_ = _zz_2093_[14];
  assign _zz_2109_ = _zz_2093_[15];
  assign _zz_2110_ = _zz_2093_[16];
  assign _zz_2111_ = _zz_2093_[17];
  assign _zz_2112_ = _zz_2093_[18];
  assign _zz_2113_ = _zz_2093_[19];
  assign _zz_2114_ = _zz_2093_[20];
  assign _zz_2115_ = _zz_2093_[21];
  assign _zz_2116_ = _zz_2093_[22];
  assign _zz_2117_ = _zz_2093_[23];
  assign _zz_2118_ = _zz_2093_[24];
  assign _zz_2119_ = _zz_2093_[25];
  assign _zz_2120_ = _zz_2093_[26];
  assign _zz_2121_ = _zz_2093_[27];
  assign _zz_2122_ = _zz_2093_[28];
  assign _zz_2123_ = _zz_2093_[29];
  assign _zz_2124_ = _zz_2093_[30];
  assign _zz_2125_ = _zz_2093_[31];
  assign _zz_2126_ = _zz_2093_[32];
  assign _zz_2127_ = _zz_2093_[33];
  assign _zz_2128_ = _zz_2093_[34];
  assign _zz_2129_ = _zz_2093_[35];
  assign _zz_2130_ = _zz_2093_[36];
  assign _zz_2131_ = _zz_2093_[37];
  assign _zz_2132_ = _zz_2093_[38];
  assign _zz_2133_ = _zz_2093_[39];
  assign _zz_2134_ = _zz_2093_[40];
  assign _zz_2135_ = _zz_2093_[41];
  assign _zz_2136_ = _zz_2093_[42];
  assign _zz_2137_ = _zz_2093_[43];
  assign _zz_2138_ = _zz_2093_[44];
  assign _zz_2139_ = _zz_2093_[45];
  assign _zz_2140_ = _zz_2093_[46];
  assign _zz_2141_ = _zz_2093_[47];
  assign _zz_2142_ = _zz_2093_[48];
  assign _zz_2143_ = _zz_2093_[49];
  assign _zz_2144_ = (((32'h000002ee <= load_data_area_current_addr) && (load_data_area_current_addr < 32'h00000320)) ? axi4_w_payload_data_regNext : {_zz_2829_,_zz_2830_});
  assign _zz_2145_ = _zz_2144_[15 : 0];
  assign _zz_2146_ = _zz_2144_[31 : 16];
  assign _zz_2147_ = _zz_2896_[5:0];
  assign _zz_2148_ = ({63'd0,(1'b1)} <<< _zz_2147_);
  assign _zz_2149_ = _zz_2148_[0];
  assign _zz_2150_ = _zz_2148_[1];
  assign _zz_2151_ = _zz_2148_[2];
  assign _zz_2152_ = _zz_2148_[3];
  assign _zz_2153_ = _zz_2148_[4];
  assign _zz_2154_ = _zz_2148_[5];
  assign _zz_2155_ = _zz_2148_[6];
  assign _zz_2156_ = _zz_2148_[7];
  assign _zz_2157_ = _zz_2148_[8];
  assign _zz_2158_ = _zz_2148_[9];
  assign _zz_2159_ = _zz_2148_[10];
  assign _zz_2160_ = _zz_2148_[11];
  assign _zz_2161_ = _zz_2148_[12];
  assign _zz_2162_ = _zz_2148_[13];
  assign _zz_2163_ = _zz_2148_[14];
  assign _zz_2164_ = _zz_2148_[15];
  assign _zz_2165_ = _zz_2148_[16];
  assign _zz_2166_ = _zz_2148_[17];
  assign _zz_2167_ = _zz_2148_[18];
  assign _zz_2168_ = _zz_2148_[19];
  assign _zz_2169_ = _zz_2148_[20];
  assign _zz_2170_ = _zz_2148_[21];
  assign _zz_2171_ = _zz_2148_[22];
  assign _zz_2172_ = _zz_2148_[23];
  assign _zz_2173_ = _zz_2148_[24];
  assign _zz_2174_ = _zz_2148_[25];
  assign _zz_2175_ = _zz_2148_[26];
  assign _zz_2176_ = _zz_2148_[27];
  assign _zz_2177_ = _zz_2148_[28];
  assign _zz_2178_ = _zz_2148_[29];
  assign _zz_2179_ = _zz_2148_[30];
  assign _zz_2180_ = _zz_2148_[31];
  assign _zz_2181_ = _zz_2148_[32];
  assign _zz_2182_ = _zz_2148_[33];
  assign _zz_2183_ = _zz_2148_[34];
  assign _zz_2184_ = _zz_2148_[35];
  assign _zz_2185_ = _zz_2148_[36];
  assign _zz_2186_ = _zz_2148_[37];
  assign _zz_2187_ = _zz_2148_[38];
  assign _zz_2188_ = _zz_2148_[39];
  assign _zz_2189_ = _zz_2148_[40];
  assign _zz_2190_ = _zz_2148_[41];
  assign _zz_2191_ = _zz_2148_[42];
  assign _zz_2192_ = _zz_2148_[43];
  assign _zz_2193_ = _zz_2148_[44];
  assign _zz_2194_ = _zz_2148_[45];
  assign _zz_2195_ = _zz_2148_[46];
  assign _zz_2196_ = _zz_2148_[47];
  assign _zz_2197_ = _zz_2148_[48];
  assign _zz_2198_ = _zz_2148_[49];
  assign _zz_2199_ = (((32'h000008fc <= load_data_area_current_addr) && (load_data_area_current_addr < 32'h0000092e)) ? axi4_w_payload_data_regNext : {_zz_2831_,_zz_2832_});
  assign _zz_2200_ = _zz_2199_[15 : 0];
  assign _zz_2201_ = _zz_2199_[31 : 16];
  assign _zz_2202_ = _zz_2897_[5:0];
  assign _zz_2203_ = ({63'd0,(1'b1)} <<< _zz_2202_);
  assign _zz_2204_ = _zz_2203_[0];
  assign _zz_2205_ = _zz_2203_[1];
  assign _zz_2206_ = _zz_2203_[2];
  assign _zz_2207_ = _zz_2203_[3];
  assign _zz_2208_ = _zz_2203_[4];
  assign _zz_2209_ = _zz_2203_[5];
  assign _zz_2210_ = _zz_2203_[6];
  assign _zz_2211_ = _zz_2203_[7];
  assign _zz_2212_ = _zz_2203_[8];
  assign _zz_2213_ = _zz_2203_[9];
  assign _zz_2214_ = _zz_2203_[10];
  assign _zz_2215_ = _zz_2203_[11];
  assign _zz_2216_ = _zz_2203_[12];
  assign _zz_2217_ = _zz_2203_[13];
  assign _zz_2218_ = _zz_2203_[14];
  assign _zz_2219_ = _zz_2203_[15];
  assign _zz_2220_ = _zz_2203_[16];
  assign _zz_2221_ = _zz_2203_[17];
  assign _zz_2222_ = _zz_2203_[18];
  assign _zz_2223_ = _zz_2203_[19];
  assign _zz_2224_ = _zz_2203_[20];
  assign _zz_2225_ = _zz_2203_[21];
  assign _zz_2226_ = _zz_2203_[22];
  assign _zz_2227_ = _zz_2203_[23];
  assign _zz_2228_ = _zz_2203_[24];
  assign _zz_2229_ = _zz_2203_[25];
  assign _zz_2230_ = _zz_2203_[26];
  assign _zz_2231_ = _zz_2203_[27];
  assign _zz_2232_ = _zz_2203_[28];
  assign _zz_2233_ = _zz_2203_[29];
  assign _zz_2234_ = _zz_2203_[30];
  assign _zz_2235_ = _zz_2203_[31];
  assign _zz_2236_ = _zz_2203_[32];
  assign _zz_2237_ = _zz_2203_[33];
  assign _zz_2238_ = _zz_2203_[34];
  assign _zz_2239_ = _zz_2203_[35];
  assign _zz_2240_ = _zz_2203_[36];
  assign _zz_2241_ = _zz_2203_[37];
  assign _zz_2242_ = _zz_2203_[38];
  assign _zz_2243_ = _zz_2203_[39];
  assign _zz_2244_ = _zz_2203_[40];
  assign _zz_2245_ = _zz_2203_[41];
  assign _zz_2246_ = _zz_2203_[42];
  assign _zz_2247_ = _zz_2203_[43];
  assign _zz_2248_ = _zz_2203_[44];
  assign _zz_2249_ = _zz_2203_[45];
  assign _zz_2250_ = _zz_2203_[46];
  assign _zz_2251_ = _zz_2203_[47];
  assign _zz_2252_ = _zz_2203_[48];
  assign _zz_2253_ = _zz_2203_[49];
  assign _zz_2254_ = (((32'h0 <= load_data_area_current_addr) && (load_data_area_current_addr < 32'h00000032)) ? axi4_w_payload_data_regNext : {_zz_2833_,_zz_2834_});
  assign _zz_2255_ = _zz_2254_[15 : 0];
  assign _zz_2256_ = _zz_2254_[31 : 16];
  assign _zz_2257_ = _zz_2898_[5:0];
  assign _zz_2258_ = ({63'd0,(1'b1)} <<< _zz_2257_);
  assign _zz_2259_ = _zz_2258_[0];
  assign _zz_2260_ = _zz_2258_[1];
  assign _zz_2261_ = _zz_2258_[2];
  assign _zz_2262_ = _zz_2258_[3];
  assign _zz_2263_ = _zz_2258_[4];
  assign _zz_2264_ = _zz_2258_[5];
  assign _zz_2265_ = _zz_2258_[6];
  assign _zz_2266_ = _zz_2258_[7];
  assign _zz_2267_ = _zz_2258_[8];
  assign _zz_2268_ = _zz_2258_[9];
  assign _zz_2269_ = _zz_2258_[10];
  assign _zz_2270_ = _zz_2258_[11];
  assign _zz_2271_ = _zz_2258_[12];
  assign _zz_2272_ = _zz_2258_[13];
  assign _zz_2273_ = _zz_2258_[14];
  assign _zz_2274_ = _zz_2258_[15];
  assign _zz_2275_ = _zz_2258_[16];
  assign _zz_2276_ = _zz_2258_[17];
  assign _zz_2277_ = _zz_2258_[18];
  assign _zz_2278_ = _zz_2258_[19];
  assign _zz_2279_ = _zz_2258_[20];
  assign _zz_2280_ = _zz_2258_[21];
  assign _zz_2281_ = _zz_2258_[22];
  assign _zz_2282_ = _zz_2258_[23];
  assign _zz_2283_ = _zz_2258_[24];
  assign _zz_2284_ = _zz_2258_[25];
  assign _zz_2285_ = _zz_2258_[26];
  assign _zz_2286_ = _zz_2258_[27];
  assign _zz_2287_ = _zz_2258_[28];
  assign _zz_2288_ = _zz_2258_[29];
  assign _zz_2289_ = _zz_2258_[30];
  assign _zz_2290_ = _zz_2258_[31];
  assign _zz_2291_ = _zz_2258_[32];
  assign _zz_2292_ = _zz_2258_[33];
  assign _zz_2293_ = _zz_2258_[34];
  assign _zz_2294_ = _zz_2258_[35];
  assign _zz_2295_ = _zz_2258_[36];
  assign _zz_2296_ = _zz_2258_[37];
  assign _zz_2297_ = _zz_2258_[38];
  assign _zz_2298_ = _zz_2258_[39];
  assign _zz_2299_ = _zz_2258_[40];
  assign _zz_2300_ = _zz_2258_[41];
  assign _zz_2301_ = _zz_2258_[42];
  assign _zz_2302_ = _zz_2258_[43];
  assign _zz_2303_ = _zz_2258_[44];
  assign _zz_2304_ = _zz_2258_[45];
  assign _zz_2305_ = _zz_2258_[46];
  assign _zz_2306_ = _zz_2258_[47];
  assign _zz_2307_ = _zz_2258_[48];
  assign _zz_2308_ = _zz_2258_[49];
  assign _zz_2309_ = (((32'h0000044c <= load_data_area_current_addr) && (load_data_area_current_addr < 32'h0000047e)) ? axi4_w_payload_data_regNext : {_zz_2835_,_zz_2836_});
  assign _zz_2310_ = _zz_2309_[15 : 0];
  assign _zz_2311_ = _zz_2309_[31 : 16];
  assign _zz_2312_ = _zz_2899_[5:0];
  assign _zz_2313_ = ({63'd0,(1'b1)} <<< _zz_2312_);
  assign _zz_2314_ = _zz_2313_[0];
  assign _zz_2315_ = _zz_2313_[1];
  assign _zz_2316_ = _zz_2313_[2];
  assign _zz_2317_ = _zz_2313_[3];
  assign _zz_2318_ = _zz_2313_[4];
  assign _zz_2319_ = _zz_2313_[5];
  assign _zz_2320_ = _zz_2313_[6];
  assign _zz_2321_ = _zz_2313_[7];
  assign _zz_2322_ = _zz_2313_[8];
  assign _zz_2323_ = _zz_2313_[9];
  assign _zz_2324_ = _zz_2313_[10];
  assign _zz_2325_ = _zz_2313_[11];
  assign _zz_2326_ = _zz_2313_[12];
  assign _zz_2327_ = _zz_2313_[13];
  assign _zz_2328_ = _zz_2313_[14];
  assign _zz_2329_ = _zz_2313_[15];
  assign _zz_2330_ = _zz_2313_[16];
  assign _zz_2331_ = _zz_2313_[17];
  assign _zz_2332_ = _zz_2313_[18];
  assign _zz_2333_ = _zz_2313_[19];
  assign _zz_2334_ = _zz_2313_[20];
  assign _zz_2335_ = _zz_2313_[21];
  assign _zz_2336_ = _zz_2313_[22];
  assign _zz_2337_ = _zz_2313_[23];
  assign _zz_2338_ = _zz_2313_[24];
  assign _zz_2339_ = _zz_2313_[25];
  assign _zz_2340_ = _zz_2313_[26];
  assign _zz_2341_ = _zz_2313_[27];
  assign _zz_2342_ = _zz_2313_[28];
  assign _zz_2343_ = _zz_2313_[29];
  assign _zz_2344_ = _zz_2313_[30];
  assign _zz_2345_ = _zz_2313_[31];
  assign _zz_2346_ = _zz_2313_[32];
  assign _zz_2347_ = _zz_2313_[33];
  assign _zz_2348_ = _zz_2313_[34];
  assign _zz_2349_ = _zz_2313_[35];
  assign _zz_2350_ = _zz_2313_[36];
  assign _zz_2351_ = _zz_2313_[37];
  assign _zz_2352_ = _zz_2313_[38];
  assign _zz_2353_ = _zz_2313_[39];
  assign _zz_2354_ = _zz_2313_[40];
  assign _zz_2355_ = _zz_2313_[41];
  assign _zz_2356_ = _zz_2313_[42];
  assign _zz_2357_ = _zz_2313_[43];
  assign _zz_2358_ = _zz_2313_[44];
  assign _zz_2359_ = _zz_2313_[45];
  assign _zz_2360_ = _zz_2313_[46];
  assign _zz_2361_ = _zz_2313_[47];
  assign _zz_2362_ = _zz_2313_[48];
  assign _zz_2363_ = _zz_2313_[49];
  assign _zz_2364_ = (((32'h00000514 <= load_data_area_current_addr) && (load_data_area_current_addr < 32'h00000546)) ? axi4_w_payload_data_regNext : {_zz_2837_,_zz_2838_});
  assign _zz_2365_ = _zz_2364_[15 : 0];
  assign _zz_2366_ = _zz_2364_[31 : 16];
  assign _zz_2367_ = _zz_2900_[5:0];
  assign _zz_2368_ = ({63'd0,(1'b1)} <<< _zz_2367_);
  assign _zz_2369_ = _zz_2368_[0];
  assign _zz_2370_ = _zz_2368_[1];
  assign _zz_2371_ = _zz_2368_[2];
  assign _zz_2372_ = _zz_2368_[3];
  assign _zz_2373_ = _zz_2368_[4];
  assign _zz_2374_ = _zz_2368_[5];
  assign _zz_2375_ = _zz_2368_[6];
  assign _zz_2376_ = _zz_2368_[7];
  assign _zz_2377_ = _zz_2368_[8];
  assign _zz_2378_ = _zz_2368_[9];
  assign _zz_2379_ = _zz_2368_[10];
  assign _zz_2380_ = _zz_2368_[11];
  assign _zz_2381_ = _zz_2368_[12];
  assign _zz_2382_ = _zz_2368_[13];
  assign _zz_2383_ = _zz_2368_[14];
  assign _zz_2384_ = _zz_2368_[15];
  assign _zz_2385_ = _zz_2368_[16];
  assign _zz_2386_ = _zz_2368_[17];
  assign _zz_2387_ = _zz_2368_[18];
  assign _zz_2388_ = _zz_2368_[19];
  assign _zz_2389_ = _zz_2368_[20];
  assign _zz_2390_ = _zz_2368_[21];
  assign _zz_2391_ = _zz_2368_[22];
  assign _zz_2392_ = _zz_2368_[23];
  assign _zz_2393_ = _zz_2368_[24];
  assign _zz_2394_ = _zz_2368_[25];
  assign _zz_2395_ = _zz_2368_[26];
  assign _zz_2396_ = _zz_2368_[27];
  assign _zz_2397_ = _zz_2368_[28];
  assign _zz_2398_ = _zz_2368_[29];
  assign _zz_2399_ = _zz_2368_[30];
  assign _zz_2400_ = _zz_2368_[31];
  assign _zz_2401_ = _zz_2368_[32];
  assign _zz_2402_ = _zz_2368_[33];
  assign _zz_2403_ = _zz_2368_[34];
  assign _zz_2404_ = _zz_2368_[35];
  assign _zz_2405_ = _zz_2368_[36];
  assign _zz_2406_ = _zz_2368_[37];
  assign _zz_2407_ = _zz_2368_[38];
  assign _zz_2408_ = _zz_2368_[39];
  assign _zz_2409_ = _zz_2368_[40];
  assign _zz_2410_ = _zz_2368_[41];
  assign _zz_2411_ = _zz_2368_[42];
  assign _zz_2412_ = _zz_2368_[43];
  assign _zz_2413_ = _zz_2368_[44];
  assign _zz_2414_ = _zz_2368_[45];
  assign _zz_2415_ = _zz_2368_[46];
  assign _zz_2416_ = _zz_2368_[47];
  assign _zz_2417_ = _zz_2368_[48];
  assign _zz_2418_ = _zz_2368_[49];
  assign _zz_2419_ = (((32'h0000092e <= load_data_area_current_addr) && (load_data_area_current_addr < 32'h00000960)) ? axi4_w_payload_data_regNext : {_zz_2839_,_zz_2840_});
  assign _zz_2420_ = _zz_2419_[15 : 0];
  assign _zz_2421_ = _zz_2419_[31 : 16];
  assign _zz_2422_ = _zz_2901_[5:0];
  assign _zz_2423_ = ({63'd0,(1'b1)} <<< _zz_2422_);
  assign _zz_2424_ = _zz_2423_[0];
  assign _zz_2425_ = _zz_2423_[1];
  assign _zz_2426_ = _zz_2423_[2];
  assign _zz_2427_ = _zz_2423_[3];
  assign _zz_2428_ = _zz_2423_[4];
  assign _zz_2429_ = _zz_2423_[5];
  assign _zz_2430_ = _zz_2423_[6];
  assign _zz_2431_ = _zz_2423_[7];
  assign _zz_2432_ = _zz_2423_[8];
  assign _zz_2433_ = _zz_2423_[9];
  assign _zz_2434_ = _zz_2423_[10];
  assign _zz_2435_ = _zz_2423_[11];
  assign _zz_2436_ = _zz_2423_[12];
  assign _zz_2437_ = _zz_2423_[13];
  assign _zz_2438_ = _zz_2423_[14];
  assign _zz_2439_ = _zz_2423_[15];
  assign _zz_2440_ = _zz_2423_[16];
  assign _zz_2441_ = _zz_2423_[17];
  assign _zz_2442_ = _zz_2423_[18];
  assign _zz_2443_ = _zz_2423_[19];
  assign _zz_2444_ = _zz_2423_[20];
  assign _zz_2445_ = _zz_2423_[21];
  assign _zz_2446_ = _zz_2423_[22];
  assign _zz_2447_ = _zz_2423_[23];
  assign _zz_2448_ = _zz_2423_[24];
  assign _zz_2449_ = _zz_2423_[25];
  assign _zz_2450_ = _zz_2423_[26];
  assign _zz_2451_ = _zz_2423_[27];
  assign _zz_2452_ = _zz_2423_[28];
  assign _zz_2453_ = _zz_2423_[29];
  assign _zz_2454_ = _zz_2423_[30];
  assign _zz_2455_ = _zz_2423_[31];
  assign _zz_2456_ = _zz_2423_[32];
  assign _zz_2457_ = _zz_2423_[33];
  assign _zz_2458_ = _zz_2423_[34];
  assign _zz_2459_ = _zz_2423_[35];
  assign _zz_2460_ = _zz_2423_[36];
  assign _zz_2461_ = _zz_2423_[37];
  assign _zz_2462_ = _zz_2423_[38];
  assign _zz_2463_ = _zz_2423_[39];
  assign _zz_2464_ = _zz_2423_[40];
  assign _zz_2465_ = _zz_2423_[41];
  assign _zz_2466_ = _zz_2423_[42];
  assign _zz_2467_ = _zz_2423_[43];
  assign _zz_2468_ = _zz_2423_[44];
  assign _zz_2469_ = _zz_2423_[45];
  assign _zz_2470_ = _zz_2423_[46];
  assign _zz_2471_ = _zz_2423_[47];
  assign _zz_2472_ = _zz_2423_[48];
  assign _zz_2473_ = _zz_2423_[49];
  assign _zz_2474_ = (((32'h00000708 <= load_data_area_current_addr) && (load_data_area_current_addr < 32'h0000073a)) ? axi4_w_payload_data_regNext : {_zz_2841_,_zz_2842_});
  assign _zz_2475_ = _zz_2474_[15 : 0];
  assign _zz_2476_ = _zz_2474_[31 : 16];
  assign _zz_2477_ = _zz_2902_[5:0];
  assign _zz_2478_ = ({63'd0,(1'b1)} <<< _zz_2477_);
  assign _zz_2479_ = _zz_2478_[0];
  assign _zz_2480_ = _zz_2478_[1];
  assign _zz_2481_ = _zz_2478_[2];
  assign _zz_2482_ = _zz_2478_[3];
  assign _zz_2483_ = _zz_2478_[4];
  assign _zz_2484_ = _zz_2478_[5];
  assign _zz_2485_ = _zz_2478_[6];
  assign _zz_2486_ = _zz_2478_[7];
  assign _zz_2487_ = _zz_2478_[8];
  assign _zz_2488_ = _zz_2478_[9];
  assign _zz_2489_ = _zz_2478_[10];
  assign _zz_2490_ = _zz_2478_[11];
  assign _zz_2491_ = _zz_2478_[12];
  assign _zz_2492_ = _zz_2478_[13];
  assign _zz_2493_ = _zz_2478_[14];
  assign _zz_2494_ = _zz_2478_[15];
  assign _zz_2495_ = _zz_2478_[16];
  assign _zz_2496_ = _zz_2478_[17];
  assign _zz_2497_ = _zz_2478_[18];
  assign _zz_2498_ = _zz_2478_[19];
  assign _zz_2499_ = _zz_2478_[20];
  assign _zz_2500_ = _zz_2478_[21];
  assign _zz_2501_ = _zz_2478_[22];
  assign _zz_2502_ = _zz_2478_[23];
  assign _zz_2503_ = _zz_2478_[24];
  assign _zz_2504_ = _zz_2478_[25];
  assign _zz_2505_ = _zz_2478_[26];
  assign _zz_2506_ = _zz_2478_[27];
  assign _zz_2507_ = _zz_2478_[28];
  assign _zz_2508_ = _zz_2478_[29];
  assign _zz_2509_ = _zz_2478_[30];
  assign _zz_2510_ = _zz_2478_[31];
  assign _zz_2511_ = _zz_2478_[32];
  assign _zz_2512_ = _zz_2478_[33];
  assign _zz_2513_ = _zz_2478_[34];
  assign _zz_2514_ = _zz_2478_[35];
  assign _zz_2515_ = _zz_2478_[36];
  assign _zz_2516_ = _zz_2478_[37];
  assign _zz_2517_ = _zz_2478_[38];
  assign _zz_2518_ = _zz_2478_[39];
  assign _zz_2519_ = _zz_2478_[40];
  assign _zz_2520_ = _zz_2478_[41];
  assign _zz_2521_ = _zz_2478_[42];
  assign _zz_2522_ = _zz_2478_[43];
  assign _zz_2523_ = _zz_2478_[44];
  assign _zz_2524_ = _zz_2478_[45];
  assign _zz_2525_ = _zz_2478_[46];
  assign _zz_2526_ = _zz_2478_[47];
  assign _zz_2527_ = _zz_2478_[48];
  assign _zz_2528_ = _zz_2478_[49];
  assign _zz_2529_ = (((32'h0000060e <= load_data_area_current_addr) && (load_data_area_current_addr < 32'h00000640)) ? axi4_w_payload_data_regNext : {_zz_2843_,_zz_2844_});
  assign _zz_2530_ = _zz_2529_[15 : 0];
  assign _zz_2531_ = _zz_2529_[31 : 16];
  assign _zz_2532_ = _zz_2903_[5:0];
  assign _zz_2533_ = ({63'd0,(1'b1)} <<< _zz_2532_);
  assign _zz_2534_ = _zz_2533_[0];
  assign _zz_2535_ = _zz_2533_[1];
  assign _zz_2536_ = _zz_2533_[2];
  assign _zz_2537_ = _zz_2533_[3];
  assign _zz_2538_ = _zz_2533_[4];
  assign _zz_2539_ = _zz_2533_[5];
  assign _zz_2540_ = _zz_2533_[6];
  assign _zz_2541_ = _zz_2533_[7];
  assign _zz_2542_ = _zz_2533_[8];
  assign _zz_2543_ = _zz_2533_[9];
  assign _zz_2544_ = _zz_2533_[10];
  assign _zz_2545_ = _zz_2533_[11];
  assign _zz_2546_ = _zz_2533_[12];
  assign _zz_2547_ = _zz_2533_[13];
  assign _zz_2548_ = _zz_2533_[14];
  assign _zz_2549_ = _zz_2533_[15];
  assign _zz_2550_ = _zz_2533_[16];
  assign _zz_2551_ = _zz_2533_[17];
  assign _zz_2552_ = _zz_2533_[18];
  assign _zz_2553_ = _zz_2533_[19];
  assign _zz_2554_ = _zz_2533_[20];
  assign _zz_2555_ = _zz_2533_[21];
  assign _zz_2556_ = _zz_2533_[22];
  assign _zz_2557_ = _zz_2533_[23];
  assign _zz_2558_ = _zz_2533_[24];
  assign _zz_2559_ = _zz_2533_[25];
  assign _zz_2560_ = _zz_2533_[26];
  assign _zz_2561_ = _zz_2533_[27];
  assign _zz_2562_ = _zz_2533_[28];
  assign _zz_2563_ = _zz_2533_[29];
  assign _zz_2564_ = _zz_2533_[30];
  assign _zz_2565_ = _zz_2533_[31];
  assign _zz_2566_ = _zz_2533_[32];
  assign _zz_2567_ = _zz_2533_[33];
  assign _zz_2568_ = _zz_2533_[34];
  assign _zz_2569_ = _zz_2533_[35];
  assign _zz_2570_ = _zz_2533_[36];
  assign _zz_2571_ = _zz_2533_[37];
  assign _zz_2572_ = _zz_2533_[38];
  assign _zz_2573_ = _zz_2533_[39];
  assign _zz_2574_ = _zz_2533_[40];
  assign _zz_2575_ = _zz_2533_[41];
  assign _zz_2576_ = _zz_2533_[42];
  assign _zz_2577_ = _zz_2533_[43];
  assign _zz_2578_ = _zz_2533_[44];
  assign _zz_2579_ = _zz_2533_[45];
  assign _zz_2580_ = _zz_2533_[46];
  assign _zz_2581_ = _zz_2533_[47];
  assign _zz_2582_ = _zz_2533_[48];
  assign _zz_2583_ = _zz_2533_[49];
  assign _zz_2584_ = (((32'h000000fa <= load_data_area_current_addr) && (load_data_area_current_addr < 32'h0000012c)) ? axi4_w_payload_data_regNext : {_zz_2845_,_zz_2846_});
  assign _zz_2585_ = _zz_2584_[15 : 0];
  assign _zz_2586_ = _zz_2584_[31 : 16];
  assign _zz_2587_ = _zz_2904_[5:0];
  assign _zz_2588_ = ({63'd0,(1'b1)} <<< _zz_2587_);
  assign _zz_2589_ = _zz_2588_[0];
  assign _zz_2590_ = _zz_2588_[1];
  assign _zz_2591_ = _zz_2588_[2];
  assign _zz_2592_ = _zz_2588_[3];
  assign _zz_2593_ = _zz_2588_[4];
  assign _zz_2594_ = _zz_2588_[5];
  assign _zz_2595_ = _zz_2588_[6];
  assign _zz_2596_ = _zz_2588_[7];
  assign _zz_2597_ = _zz_2588_[8];
  assign _zz_2598_ = _zz_2588_[9];
  assign _zz_2599_ = _zz_2588_[10];
  assign _zz_2600_ = _zz_2588_[11];
  assign _zz_2601_ = _zz_2588_[12];
  assign _zz_2602_ = _zz_2588_[13];
  assign _zz_2603_ = _zz_2588_[14];
  assign _zz_2604_ = _zz_2588_[15];
  assign _zz_2605_ = _zz_2588_[16];
  assign _zz_2606_ = _zz_2588_[17];
  assign _zz_2607_ = _zz_2588_[18];
  assign _zz_2608_ = _zz_2588_[19];
  assign _zz_2609_ = _zz_2588_[20];
  assign _zz_2610_ = _zz_2588_[21];
  assign _zz_2611_ = _zz_2588_[22];
  assign _zz_2612_ = _zz_2588_[23];
  assign _zz_2613_ = _zz_2588_[24];
  assign _zz_2614_ = _zz_2588_[25];
  assign _zz_2615_ = _zz_2588_[26];
  assign _zz_2616_ = _zz_2588_[27];
  assign _zz_2617_ = _zz_2588_[28];
  assign _zz_2618_ = _zz_2588_[29];
  assign _zz_2619_ = _zz_2588_[30];
  assign _zz_2620_ = _zz_2588_[31];
  assign _zz_2621_ = _zz_2588_[32];
  assign _zz_2622_ = _zz_2588_[33];
  assign _zz_2623_ = _zz_2588_[34];
  assign _zz_2624_ = _zz_2588_[35];
  assign _zz_2625_ = _zz_2588_[36];
  assign _zz_2626_ = _zz_2588_[37];
  assign _zz_2627_ = _zz_2588_[38];
  assign _zz_2628_ = _zz_2588_[39];
  assign _zz_2629_ = _zz_2588_[40];
  assign _zz_2630_ = _zz_2588_[41];
  assign _zz_2631_ = _zz_2588_[42];
  assign _zz_2632_ = _zz_2588_[43];
  assign _zz_2633_ = _zz_2588_[44];
  assign _zz_2634_ = _zz_2588_[45];
  assign _zz_2635_ = _zz_2588_[46];
  assign _zz_2636_ = _zz_2588_[47];
  assign _zz_2637_ = _zz_2588_[48];
  assign _zz_2638_ = _zz_2588_[49];
  assign _zz_2639_ = (((32'h000007d0 <= load_data_area_current_addr) && (load_data_area_current_addr < 32'h00000802)) ? axi4_w_payload_data_regNext : {_zz_2847_,_zz_2848_});
  assign _zz_2640_ = _zz_2639_[15 : 0];
  assign _zz_2641_ = _zz_2639_[31 : 16];
  assign _zz_2642_ = _zz_2905_[5:0];
  assign _zz_2643_ = ({63'd0,(1'b1)} <<< _zz_2642_);
  assign _zz_2644_ = _zz_2643_[0];
  assign _zz_2645_ = _zz_2643_[1];
  assign _zz_2646_ = _zz_2643_[2];
  assign _zz_2647_ = _zz_2643_[3];
  assign _zz_2648_ = _zz_2643_[4];
  assign _zz_2649_ = _zz_2643_[5];
  assign _zz_2650_ = _zz_2643_[6];
  assign _zz_2651_ = _zz_2643_[7];
  assign _zz_2652_ = _zz_2643_[8];
  assign _zz_2653_ = _zz_2643_[9];
  assign _zz_2654_ = _zz_2643_[10];
  assign _zz_2655_ = _zz_2643_[11];
  assign _zz_2656_ = _zz_2643_[12];
  assign _zz_2657_ = _zz_2643_[13];
  assign _zz_2658_ = _zz_2643_[14];
  assign _zz_2659_ = _zz_2643_[15];
  assign _zz_2660_ = _zz_2643_[16];
  assign _zz_2661_ = _zz_2643_[17];
  assign _zz_2662_ = _zz_2643_[18];
  assign _zz_2663_ = _zz_2643_[19];
  assign _zz_2664_ = _zz_2643_[20];
  assign _zz_2665_ = _zz_2643_[21];
  assign _zz_2666_ = _zz_2643_[22];
  assign _zz_2667_ = _zz_2643_[23];
  assign _zz_2668_ = _zz_2643_[24];
  assign _zz_2669_ = _zz_2643_[25];
  assign _zz_2670_ = _zz_2643_[26];
  assign _zz_2671_ = _zz_2643_[27];
  assign _zz_2672_ = _zz_2643_[28];
  assign _zz_2673_ = _zz_2643_[29];
  assign _zz_2674_ = _zz_2643_[30];
  assign _zz_2675_ = _zz_2643_[31];
  assign _zz_2676_ = _zz_2643_[32];
  assign _zz_2677_ = _zz_2643_[33];
  assign _zz_2678_ = _zz_2643_[34];
  assign _zz_2679_ = _zz_2643_[35];
  assign _zz_2680_ = _zz_2643_[36];
  assign _zz_2681_ = _zz_2643_[37];
  assign _zz_2682_ = _zz_2643_[38];
  assign _zz_2683_ = _zz_2643_[39];
  assign _zz_2684_ = _zz_2643_[40];
  assign _zz_2685_ = _zz_2643_[41];
  assign _zz_2686_ = _zz_2643_[42];
  assign _zz_2687_ = _zz_2643_[43];
  assign _zz_2688_ = _zz_2643_[44];
  assign _zz_2689_ = _zz_2643_[45];
  assign _zz_2690_ = _zz_2643_[46];
  assign _zz_2691_ = _zz_2643_[47];
  assign _zz_2692_ = _zz_2643_[48];
  assign _zz_2693_ = _zz_2643_[49];
  assign _zz_2694_ = (((32'h0000079e <= load_data_area_current_addr) && (load_data_area_current_addr < 32'h000007d0)) ? axi4_w_payload_data_regNext : {_zz_2849_,_zz_2850_});
  assign _zz_2695_ = _zz_2694_[15 : 0];
  assign _zz_2696_ = _zz_2694_[31 : 16];
  assign _zz_2697_ = _zz_2906_[5:0];
  assign _zz_2698_ = ({63'd0,(1'b1)} <<< _zz_2697_);
  assign _zz_2699_ = _zz_2698_[0];
  assign _zz_2700_ = _zz_2698_[1];
  assign _zz_2701_ = _zz_2698_[2];
  assign _zz_2702_ = _zz_2698_[3];
  assign _zz_2703_ = _zz_2698_[4];
  assign _zz_2704_ = _zz_2698_[5];
  assign _zz_2705_ = _zz_2698_[6];
  assign _zz_2706_ = _zz_2698_[7];
  assign _zz_2707_ = _zz_2698_[8];
  assign _zz_2708_ = _zz_2698_[9];
  assign _zz_2709_ = _zz_2698_[10];
  assign _zz_2710_ = _zz_2698_[11];
  assign _zz_2711_ = _zz_2698_[12];
  assign _zz_2712_ = _zz_2698_[13];
  assign _zz_2713_ = _zz_2698_[14];
  assign _zz_2714_ = _zz_2698_[15];
  assign _zz_2715_ = _zz_2698_[16];
  assign _zz_2716_ = _zz_2698_[17];
  assign _zz_2717_ = _zz_2698_[18];
  assign _zz_2718_ = _zz_2698_[19];
  assign _zz_2719_ = _zz_2698_[20];
  assign _zz_2720_ = _zz_2698_[21];
  assign _zz_2721_ = _zz_2698_[22];
  assign _zz_2722_ = _zz_2698_[23];
  assign _zz_2723_ = _zz_2698_[24];
  assign _zz_2724_ = _zz_2698_[25];
  assign _zz_2725_ = _zz_2698_[26];
  assign _zz_2726_ = _zz_2698_[27];
  assign _zz_2727_ = _zz_2698_[28];
  assign _zz_2728_ = _zz_2698_[29];
  assign _zz_2729_ = _zz_2698_[30];
  assign _zz_2730_ = _zz_2698_[31];
  assign _zz_2731_ = _zz_2698_[32];
  assign _zz_2732_ = _zz_2698_[33];
  assign _zz_2733_ = _zz_2698_[34];
  assign _zz_2734_ = _zz_2698_[35];
  assign _zz_2735_ = _zz_2698_[36];
  assign _zz_2736_ = _zz_2698_[37];
  assign _zz_2737_ = _zz_2698_[38];
  assign _zz_2738_ = _zz_2698_[39];
  assign _zz_2739_ = _zz_2698_[40];
  assign _zz_2740_ = _zz_2698_[41];
  assign _zz_2741_ = _zz_2698_[42];
  assign _zz_2742_ = _zz_2698_[43];
  assign _zz_2743_ = _zz_2698_[44];
  assign _zz_2744_ = _zz_2698_[45];
  assign _zz_2745_ = _zz_2698_[46];
  assign _zz_2746_ = _zz_2698_[47];
  assign _zz_2747_ = _zz_2698_[48];
  assign _zz_2748_ = _zz_2698_[49];
  assign _zz_2749_ = (((32'h0000012c <= load_data_area_current_addr) && (load_data_area_current_addr < 32'h0000015e)) ? axi4_w_payload_data_regNext : {_zz_2851_,_zz_2852_});
  assign _zz_2750_ = _zz_2749_[15 : 0];
  assign _zz_2751_ = _zz_2749_[31 : 16];
  assign io_coef_out_valid = transfer_done;
  assign io_coef_out_payload_0_0_0_real = int_reg_array_0_0_real;
  assign io_coef_out_payload_0_0_0_imag = int_reg_array_0_0_imag;
  assign io_coef_out_payload_0_0_1_real = int_reg_array_0_1_real;
  assign io_coef_out_payload_0_0_1_imag = int_reg_array_0_1_imag;
  assign io_coef_out_payload_0_0_2_real = int_reg_array_0_2_real;
  assign io_coef_out_payload_0_0_2_imag = int_reg_array_0_2_imag;
  assign io_coef_out_payload_0_0_3_real = int_reg_array_0_3_real;
  assign io_coef_out_payload_0_0_3_imag = int_reg_array_0_3_imag;
  assign io_coef_out_payload_0_0_4_real = int_reg_array_0_4_real;
  assign io_coef_out_payload_0_0_4_imag = int_reg_array_0_4_imag;
  assign io_coef_out_payload_0_0_5_real = int_reg_array_0_5_real;
  assign io_coef_out_payload_0_0_5_imag = int_reg_array_0_5_imag;
  assign io_coef_out_payload_0_0_6_real = int_reg_array_0_6_real;
  assign io_coef_out_payload_0_0_6_imag = int_reg_array_0_6_imag;
  assign io_coef_out_payload_0_0_7_real = int_reg_array_0_7_real;
  assign io_coef_out_payload_0_0_7_imag = int_reg_array_0_7_imag;
  assign io_coef_out_payload_0_0_8_real = int_reg_array_0_8_real;
  assign io_coef_out_payload_0_0_8_imag = int_reg_array_0_8_imag;
  assign io_coef_out_payload_0_0_9_real = int_reg_array_0_9_real;
  assign io_coef_out_payload_0_0_9_imag = int_reg_array_0_9_imag;
  assign io_coef_out_payload_0_0_10_real = int_reg_array_0_10_real;
  assign io_coef_out_payload_0_0_10_imag = int_reg_array_0_10_imag;
  assign io_coef_out_payload_0_0_11_real = int_reg_array_0_11_real;
  assign io_coef_out_payload_0_0_11_imag = int_reg_array_0_11_imag;
  assign io_coef_out_payload_0_0_12_real = int_reg_array_0_12_real;
  assign io_coef_out_payload_0_0_12_imag = int_reg_array_0_12_imag;
  assign io_coef_out_payload_0_0_13_real = int_reg_array_0_13_real;
  assign io_coef_out_payload_0_0_13_imag = int_reg_array_0_13_imag;
  assign io_coef_out_payload_0_0_14_real = int_reg_array_0_14_real;
  assign io_coef_out_payload_0_0_14_imag = int_reg_array_0_14_imag;
  assign io_coef_out_payload_0_0_15_real = int_reg_array_0_15_real;
  assign io_coef_out_payload_0_0_15_imag = int_reg_array_0_15_imag;
  assign io_coef_out_payload_0_0_16_real = int_reg_array_0_16_real;
  assign io_coef_out_payload_0_0_16_imag = int_reg_array_0_16_imag;
  assign io_coef_out_payload_0_0_17_real = int_reg_array_0_17_real;
  assign io_coef_out_payload_0_0_17_imag = int_reg_array_0_17_imag;
  assign io_coef_out_payload_0_0_18_real = int_reg_array_0_18_real;
  assign io_coef_out_payload_0_0_18_imag = int_reg_array_0_18_imag;
  assign io_coef_out_payload_0_0_19_real = int_reg_array_0_19_real;
  assign io_coef_out_payload_0_0_19_imag = int_reg_array_0_19_imag;
  assign io_coef_out_payload_0_0_20_real = int_reg_array_0_20_real;
  assign io_coef_out_payload_0_0_20_imag = int_reg_array_0_20_imag;
  assign io_coef_out_payload_0_0_21_real = int_reg_array_0_21_real;
  assign io_coef_out_payload_0_0_21_imag = int_reg_array_0_21_imag;
  assign io_coef_out_payload_0_0_22_real = int_reg_array_0_22_real;
  assign io_coef_out_payload_0_0_22_imag = int_reg_array_0_22_imag;
  assign io_coef_out_payload_0_0_23_real = int_reg_array_0_23_real;
  assign io_coef_out_payload_0_0_23_imag = int_reg_array_0_23_imag;
  assign io_coef_out_payload_0_0_24_real = int_reg_array_0_24_real;
  assign io_coef_out_payload_0_0_24_imag = int_reg_array_0_24_imag;
  assign io_coef_out_payload_0_0_25_real = int_reg_array_0_25_real;
  assign io_coef_out_payload_0_0_25_imag = int_reg_array_0_25_imag;
  assign io_coef_out_payload_0_0_26_real = int_reg_array_0_26_real;
  assign io_coef_out_payload_0_0_26_imag = int_reg_array_0_26_imag;
  assign io_coef_out_payload_0_0_27_real = int_reg_array_0_27_real;
  assign io_coef_out_payload_0_0_27_imag = int_reg_array_0_27_imag;
  assign io_coef_out_payload_0_0_28_real = int_reg_array_0_28_real;
  assign io_coef_out_payload_0_0_28_imag = int_reg_array_0_28_imag;
  assign io_coef_out_payload_0_0_29_real = int_reg_array_0_29_real;
  assign io_coef_out_payload_0_0_29_imag = int_reg_array_0_29_imag;
  assign io_coef_out_payload_0_0_30_real = int_reg_array_0_30_real;
  assign io_coef_out_payload_0_0_30_imag = int_reg_array_0_30_imag;
  assign io_coef_out_payload_0_0_31_real = int_reg_array_0_31_real;
  assign io_coef_out_payload_0_0_31_imag = int_reg_array_0_31_imag;
  assign io_coef_out_payload_0_0_32_real = int_reg_array_0_32_real;
  assign io_coef_out_payload_0_0_32_imag = int_reg_array_0_32_imag;
  assign io_coef_out_payload_0_0_33_real = int_reg_array_0_33_real;
  assign io_coef_out_payload_0_0_33_imag = int_reg_array_0_33_imag;
  assign io_coef_out_payload_0_0_34_real = int_reg_array_0_34_real;
  assign io_coef_out_payload_0_0_34_imag = int_reg_array_0_34_imag;
  assign io_coef_out_payload_0_0_35_real = int_reg_array_0_35_real;
  assign io_coef_out_payload_0_0_35_imag = int_reg_array_0_35_imag;
  assign io_coef_out_payload_0_0_36_real = int_reg_array_0_36_real;
  assign io_coef_out_payload_0_0_36_imag = int_reg_array_0_36_imag;
  assign io_coef_out_payload_0_0_37_real = int_reg_array_0_37_real;
  assign io_coef_out_payload_0_0_37_imag = int_reg_array_0_37_imag;
  assign io_coef_out_payload_0_0_38_real = int_reg_array_0_38_real;
  assign io_coef_out_payload_0_0_38_imag = int_reg_array_0_38_imag;
  assign io_coef_out_payload_0_0_39_real = int_reg_array_0_39_real;
  assign io_coef_out_payload_0_0_39_imag = int_reg_array_0_39_imag;
  assign io_coef_out_payload_0_0_40_real = int_reg_array_0_40_real;
  assign io_coef_out_payload_0_0_40_imag = int_reg_array_0_40_imag;
  assign io_coef_out_payload_0_0_41_real = int_reg_array_0_41_real;
  assign io_coef_out_payload_0_0_41_imag = int_reg_array_0_41_imag;
  assign io_coef_out_payload_0_0_42_real = int_reg_array_0_42_real;
  assign io_coef_out_payload_0_0_42_imag = int_reg_array_0_42_imag;
  assign io_coef_out_payload_0_0_43_real = int_reg_array_0_43_real;
  assign io_coef_out_payload_0_0_43_imag = int_reg_array_0_43_imag;
  assign io_coef_out_payload_0_0_44_real = int_reg_array_0_44_real;
  assign io_coef_out_payload_0_0_44_imag = int_reg_array_0_44_imag;
  assign io_coef_out_payload_0_0_45_real = int_reg_array_0_45_real;
  assign io_coef_out_payload_0_0_45_imag = int_reg_array_0_45_imag;
  assign io_coef_out_payload_0_0_46_real = int_reg_array_0_46_real;
  assign io_coef_out_payload_0_0_46_imag = int_reg_array_0_46_imag;
  assign io_coef_out_payload_0_0_47_real = int_reg_array_0_47_real;
  assign io_coef_out_payload_0_0_47_imag = int_reg_array_0_47_imag;
  assign io_coef_out_payload_0_0_48_real = int_reg_array_0_48_real;
  assign io_coef_out_payload_0_0_48_imag = int_reg_array_0_48_imag;
  assign io_coef_out_payload_0_0_49_real = int_reg_array_0_49_real;
  assign io_coef_out_payload_0_0_49_imag = int_reg_array_0_49_imag;
  assign io_coef_out_payload_0_1_0_real = int_reg_array_1_0_real;
  assign io_coef_out_payload_0_1_0_imag = int_reg_array_1_0_imag;
  assign io_coef_out_payload_0_1_1_real = int_reg_array_1_1_real;
  assign io_coef_out_payload_0_1_1_imag = int_reg_array_1_1_imag;
  assign io_coef_out_payload_0_1_2_real = int_reg_array_1_2_real;
  assign io_coef_out_payload_0_1_2_imag = int_reg_array_1_2_imag;
  assign io_coef_out_payload_0_1_3_real = int_reg_array_1_3_real;
  assign io_coef_out_payload_0_1_3_imag = int_reg_array_1_3_imag;
  assign io_coef_out_payload_0_1_4_real = int_reg_array_1_4_real;
  assign io_coef_out_payload_0_1_4_imag = int_reg_array_1_4_imag;
  assign io_coef_out_payload_0_1_5_real = int_reg_array_1_5_real;
  assign io_coef_out_payload_0_1_5_imag = int_reg_array_1_5_imag;
  assign io_coef_out_payload_0_1_6_real = int_reg_array_1_6_real;
  assign io_coef_out_payload_0_1_6_imag = int_reg_array_1_6_imag;
  assign io_coef_out_payload_0_1_7_real = int_reg_array_1_7_real;
  assign io_coef_out_payload_0_1_7_imag = int_reg_array_1_7_imag;
  assign io_coef_out_payload_0_1_8_real = int_reg_array_1_8_real;
  assign io_coef_out_payload_0_1_8_imag = int_reg_array_1_8_imag;
  assign io_coef_out_payload_0_1_9_real = int_reg_array_1_9_real;
  assign io_coef_out_payload_0_1_9_imag = int_reg_array_1_9_imag;
  assign io_coef_out_payload_0_1_10_real = int_reg_array_1_10_real;
  assign io_coef_out_payload_0_1_10_imag = int_reg_array_1_10_imag;
  assign io_coef_out_payload_0_1_11_real = int_reg_array_1_11_real;
  assign io_coef_out_payload_0_1_11_imag = int_reg_array_1_11_imag;
  assign io_coef_out_payload_0_1_12_real = int_reg_array_1_12_real;
  assign io_coef_out_payload_0_1_12_imag = int_reg_array_1_12_imag;
  assign io_coef_out_payload_0_1_13_real = int_reg_array_1_13_real;
  assign io_coef_out_payload_0_1_13_imag = int_reg_array_1_13_imag;
  assign io_coef_out_payload_0_1_14_real = int_reg_array_1_14_real;
  assign io_coef_out_payload_0_1_14_imag = int_reg_array_1_14_imag;
  assign io_coef_out_payload_0_1_15_real = int_reg_array_1_15_real;
  assign io_coef_out_payload_0_1_15_imag = int_reg_array_1_15_imag;
  assign io_coef_out_payload_0_1_16_real = int_reg_array_1_16_real;
  assign io_coef_out_payload_0_1_16_imag = int_reg_array_1_16_imag;
  assign io_coef_out_payload_0_1_17_real = int_reg_array_1_17_real;
  assign io_coef_out_payload_0_1_17_imag = int_reg_array_1_17_imag;
  assign io_coef_out_payload_0_1_18_real = int_reg_array_1_18_real;
  assign io_coef_out_payload_0_1_18_imag = int_reg_array_1_18_imag;
  assign io_coef_out_payload_0_1_19_real = int_reg_array_1_19_real;
  assign io_coef_out_payload_0_1_19_imag = int_reg_array_1_19_imag;
  assign io_coef_out_payload_0_1_20_real = int_reg_array_1_20_real;
  assign io_coef_out_payload_0_1_20_imag = int_reg_array_1_20_imag;
  assign io_coef_out_payload_0_1_21_real = int_reg_array_1_21_real;
  assign io_coef_out_payload_0_1_21_imag = int_reg_array_1_21_imag;
  assign io_coef_out_payload_0_1_22_real = int_reg_array_1_22_real;
  assign io_coef_out_payload_0_1_22_imag = int_reg_array_1_22_imag;
  assign io_coef_out_payload_0_1_23_real = int_reg_array_1_23_real;
  assign io_coef_out_payload_0_1_23_imag = int_reg_array_1_23_imag;
  assign io_coef_out_payload_0_1_24_real = int_reg_array_1_24_real;
  assign io_coef_out_payload_0_1_24_imag = int_reg_array_1_24_imag;
  assign io_coef_out_payload_0_1_25_real = int_reg_array_1_25_real;
  assign io_coef_out_payload_0_1_25_imag = int_reg_array_1_25_imag;
  assign io_coef_out_payload_0_1_26_real = int_reg_array_1_26_real;
  assign io_coef_out_payload_0_1_26_imag = int_reg_array_1_26_imag;
  assign io_coef_out_payload_0_1_27_real = int_reg_array_1_27_real;
  assign io_coef_out_payload_0_1_27_imag = int_reg_array_1_27_imag;
  assign io_coef_out_payload_0_1_28_real = int_reg_array_1_28_real;
  assign io_coef_out_payload_0_1_28_imag = int_reg_array_1_28_imag;
  assign io_coef_out_payload_0_1_29_real = int_reg_array_1_29_real;
  assign io_coef_out_payload_0_1_29_imag = int_reg_array_1_29_imag;
  assign io_coef_out_payload_0_1_30_real = int_reg_array_1_30_real;
  assign io_coef_out_payload_0_1_30_imag = int_reg_array_1_30_imag;
  assign io_coef_out_payload_0_1_31_real = int_reg_array_1_31_real;
  assign io_coef_out_payload_0_1_31_imag = int_reg_array_1_31_imag;
  assign io_coef_out_payload_0_1_32_real = int_reg_array_1_32_real;
  assign io_coef_out_payload_0_1_32_imag = int_reg_array_1_32_imag;
  assign io_coef_out_payload_0_1_33_real = int_reg_array_1_33_real;
  assign io_coef_out_payload_0_1_33_imag = int_reg_array_1_33_imag;
  assign io_coef_out_payload_0_1_34_real = int_reg_array_1_34_real;
  assign io_coef_out_payload_0_1_34_imag = int_reg_array_1_34_imag;
  assign io_coef_out_payload_0_1_35_real = int_reg_array_1_35_real;
  assign io_coef_out_payload_0_1_35_imag = int_reg_array_1_35_imag;
  assign io_coef_out_payload_0_1_36_real = int_reg_array_1_36_real;
  assign io_coef_out_payload_0_1_36_imag = int_reg_array_1_36_imag;
  assign io_coef_out_payload_0_1_37_real = int_reg_array_1_37_real;
  assign io_coef_out_payload_0_1_37_imag = int_reg_array_1_37_imag;
  assign io_coef_out_payload_0_1_38_real = int_reg_array_1_38_real;
  assign io_coef_out_payload_0_1_38_imag = int_reg_array_1_38_imag;
  assign io_coef_out_payload_0_1_39_real = int_reg_array_1_39_real;
  assign io_coef_out_payload_0_1_39_imag = int_reg_array_1_39_imag;
  assign io_coef_out_payload_0_1_40_real = int_reg_array_1_40_real;
  assign io_coef_out_payload_0_1_40_imag = int_reg_array_1_40_imag;
  assign io_coef_out_payload_0_1_41_real = int_reg_array_1_41_real;
  assign io_coef_out_payload_0_1_41_imag = int_reg_array_1_41_imag;
  assign io_coef_out_payload_0_1_42_real = int_reg_array_1_42_real;
  assign io_coef_out_payload_0_1_42_imag = int_reg_array_1_42_imag;
  assign io_coef_out_payload_0_1_43_real = int_reg_array_1_43_real;
  assign io_coef_out_payload_0_1_43_imag = int_reg_array_1_43_imag;
  assign io_coef_out_payload_0_1_44_real = int_reg_array_1_44_real;
  assign io_coef_out_payload_0_1_44_imag = int_reg_array_1_44_imag;
  assign io_coef_out_payload_0_1_45_real = int_reg_array_1_45_real;
  assign io_coef_out_payload_0_1_45_imag = int_reg_array_1_45_imag;
  assign io_coef_out_payload_0_1_46_real = int_reg_array_1_46_real;
  assign io_coef_out_payload_0_1_46_imag = int_reg_array_1_46_imag;
  assign io_coef_out_payload_0_1_47_real = int_reg_array_1_47_real;
  assign io_coef_out_payload_0_1_47_imag = int_reg_array_1_47_imag;
  assign io_coef_out_payload_0_1_48_real = int_reg_array_1_48_real;
  assign io_coef_out_payload_0_1_48_imag = int_reg_array_1_48_imag;
  assign io_coef_out_payload_0_1_49_real = int_reg_array_1_49_real;
  assign io_coef_out_payload_0_1_49_imag = int_reg_array_1_49_imag;
  assign io_coef_out_payload_0_2_0_real = int_reg_array_2_0_real;
  assign io_coef_out_payload_0_2_0_imag = int_reg_array_2_0_imag;
  assign io_coef_out_payload_0_2_1_real = int_reg_array_2_1_real;
  assign io_coef_out_payload_0_2_1_imag = int_reg_array_2_1_imag;
  assign io_coef_out_payload_0_2_2_real = int_reg_array_2_2_real;
  assign io_coef_out_payload_0_2_2_imag = int_reg_array_2_2_imag;
  assign io_coef_out_payload_0_2_3_real = int_reg_array_2_3_real;
  assign io_coef_out_payload_0_2_3_imag = int_reg_array_2_3_imag;
  assign io_coef_out_payload_0_2_4_real = int_reg_array_2_4_real;
  assign io_coef_out_payload_0_2_4_imag = int_reg_array_2_4_imag;
  assign io_coef_out_payload_0_2_5_real = int_reg_array_2_5_real;
  assign io_coef_out_payload_0_2_5_imag = int_reg_array_2_5_imag;
  assign io_coef_out_payload_0_2_6_real = int_reg_array_2_6_real;
  assign io_coef_out_payload_0_2_6_imag = int_reg_array_2_6_imag;
  assign io_coef_out_payload_0_2_7_real = int_reg_array_2_7_real;
  assign io_coef_out_payload_0_2_7_imag = int_reg_array_2_7_imag;
  assign io_coef_out_payload_0_2_8_real = int_reg_array_2_8_real;
  assign io_coef_out_payload_0_2_8_imag = int_reg_array_2_8_imag;
  assign io_coef_out_payload_0_2_9_real = int_reg_array_2_9_real;
  assign io_coef_out_payload_0_2_9_imag = int_reg_array_2_9_imag;
  assign io_coef_out_payload_0_2_10_real = int_reg_array_2_10_real;
  assign io_coef_out_payload_0_2_10_imag = int_reg_array_2_10_imag;
  assign io_coef_out_payload_0_2_11_real = int_reg_array_2_11_real;
  assign io_coef_out_payload_0_2_11_imag = int_reg_array_2_11_imag;
  assign io_coef_out_payload_0_2_12_real = int_reg_array_2_12_real;
  assign io_coef_out_payload_0_2_12_imag = int_reg_array_2_12_imag;
  assign io_coef_out_payload_0_2_13_real = int_reg_array_2_13_real;
  assign io_coef_out_payload_0_2_13_imag = int_reg_array_2_13_imag;
  assign io_coef_out_payload_0_2_14_real = int_reg_array_2_14_real;
  assign io_coef_out_payload_0_2_14_imag = int_reg_array_2_14_imag;
  assign io_coef_out_payload_0_2_15_real = int_reg_array_2_15_real;
  assign io_coef_out_payload_0_2_15_imag = int_reg_array_2_15_imag;
  assign io_coef_out_payload_0_2_16_real = int_reg_array_2_16_real;
  assign io_coef_out_payload_0_2_16_imag = int_reg_array_2_16_imag;
  assign io_coef_out_payload_0_2_17_real = int_reg_array_2_17_real;
  assign io_coef_out_payload_0_2_17_imag = int_reg_array_2_17_imag;
  assign io_coef_out_payload_0_2_18_real = int_reg_array_2_18_real;
  assign io_coef_out_payload_0_2_18_imag = int_reg_array_2_18_imag;
  assign io_coef_out_payload_0_2_19_real = int_reg_array_2_19_real;
  assign io_coef_out_payload_0_2_19_imag = int_reg_array_2_19_imag;
  assign io_coef_out_payload_0_2_20_real = int_reg_array_2_20_real;
  assign io_coef_out_payload_0_2_20_imag = int_reg_array_2_20_imag;
  assign io_coef_out_payload_0_2_21_real = int_reg_array_2_21_real;
  assign io_coef_out_payload_0_2_21_imag = int_reg_array_2_21_imag;
  assign io_coef_out_payload_0_2_22_real = int_reg_array_2_22_real;
  assign io_coef_out_payload_0_2_22_imag = int_reg_array_2_22_imag;
  assign io_coef_out_payload_0_2_23_real = int_reg_array_2_23_real;
  assign io_coef_out_payload_0_2_23_imag = int_reg_array_2_23_imag;
  assign io_coef_out_payload_0_2_24_real = int_reg_array_2_24_real;
  assign io_coef_out_payload_0_2_24_imag = int_reg_array_2_24_imag;
  assign io_coef_out_payload_0_2_25_real = int_reg_array_2_25_real;
  assign io_coef_out_payload_0_2_25_imag = int_reg_array_2_25_imag;
  assign io_coef_out_payload_0_2_26_real = int_reg_array_2_26_real;
  assign io_coef_out_payload_0_2_26_imag = int_reg_array_2_26_imag;
  assign io_coef_out_payload_0_2_27_real = int_reg_array_2_27_real;
  assign io_coef_out_payload_0_2_27_imag = int_reg_array_2_27_imag;
  assign io_coef_out_payload_0_2_28_real = int_reg_array_2_28_real;
  assign io_coef_out_payload_0_2_28_imag = int_reg_array_2_28_imag;
  assign io_coef_out_payload_0_2_29_real = int_reg_array_2_29_real;
  assign io_coef_out_payload_0_2_29_imag = int_reg_array_2_29_imag;
  assign io_coef_out_payload_0_2_30_real = int_reg_array_2_30_real;
  assign io_coef_out_payload_0_2_30_imag = int_reg_array_2_30_imag;
  assign io_coef_out_payload_0_2_31_real = int_reg_array_2_31_real;
  assign io_coef_out_payload_0_2_31_imag = int_reg_array_2_31_imag;
  assign io_coef_out_payload_0_2_32_real = int_reg_array_2_32_real;
  assign io_coef_out_payload_0_2_32_imag = int_reg_array_2_32_imag;
  assign io_coef_out_payload_0_2_33_real = int_reg_array_2_33_real;
  assign io_coef_out_payload_0_2_33_imag = int_reg_array_2_33_imag;
  assign io_coef_out_payload_0_2_34_real = int_reg_array_2_34_real;
  assign io_coef_out_payload_0_2_34_imag = int_reg_array_2_34_imag;
  assign io_coef_out_payload_0_2_35_real = int_reg_array_2_35_real;
  assign io_coef_out_payload_0_2_35_imag = int_reg_array_2_35_imag;
  assign io_coef_out_payload_0_2_36_real = int_reg_array_2_36_real;
  assign io_coef_out_payload_0_2_36_imag = int_reg_array_2_36_imag;
  assign io_coef_out_payload_0_2_37_real = int_reg_array_2_37_real;
  assign io_coef_out_payload_0_2_37_imag = int_reg_array_2_37_imag;
  assign io_coef_out_payload_0_2_38_real = int_reg_array_2_38_real;
  assign io_coef_out_payload_0_2_38_imag = int_reg_array_2_38_imag;
  assign io_coef_out_payload_0_2_39_real = int_reg_array_2_39_real;
  assign io_coef_out_payload_0_2_39_imag = int_reg_array_2_39_imag;
  assign io_coef_out_payload_0_2_40_real = int_reg_array_2_40_real;
  assign io_coef_out_payload_0_2_40_imag = int_reg_array_2_40_imag;
  assign io_coef_out_payload_0_2_41_real = int_reg_array_2_41_real;
  assign io_coef_out_payload_0_2_41_imag = int_reg_array_2_41_imag;
  assign io_coef_out_payload_0_2_42_real = int_reg_array_2_42_real;
  assign io_coef_out_payload_0_2_42_imag = int_reg_array_2_42_imag;
  assign io_coef_out_payload_0_2_43_real = int_reg_array_2_43_real;
  assign io_coef_out_payload_0_2_43_imag = int_reg_array_2_43_imag;
  assign io_coef_out_payload_0_2_44_real = int_reg_array_2_44_real;
  assign io_coef_out_payload_0_2_44_imag = int_reg_array_2_44_imag;
  assign io_coef_out_payload_0_2_45_real = int_reg_array_2_45_real;
  assign io_coef_out_payload_0_2_45_imag = int_reg_array_2_45_imag;
  assign io_coef_out_payload_0_2_46_real = int_reg_array_2_46_real;
  assign io_coef_out_payload_0_2_46_imag = int_reg_array_2_46_imag;
  assign io_coef_out_payload_0_2_47_real = int_reg_array_2_47_real;
  assign io_coef_out_payload_0_2_47_imag = int_reg_array_2_47_imag;
  assign io_coef_out_payload_0_2_48_real = int_reg_array_2_48_real;
  assign io_coef_out_payload_0_2_48_imag = int_reg_array_2_48_imag;
  assign io_coef_out_payload_0_2_49_real = int_reg_array_2_49_real;
  assign io_coef_out_payload_0_2_49_imag = int_reg_array_2_49_imag;
  assign io_coef_out_payload_0_3_0_real = int_reg_array_3_0_real;
  assign io_coef_out_payload_0_3_0_imag = int_reg_array_3_0_imag;
  assign io_coef_out_payload_0_3_1_real = int_reg_array_3_1_real;
  assign io_coef_out_payload_0_3_1_imag = int_reg_array_3_1_imag;
  assign io_coef_out_payload_0_3_2_real = int_reg_array_3_2_real;
  assign io_coef_out_payload_0_3_2_imag = int_reg_array_3_2_imag;
  assign io_coef_out_payload_0_3_3_real = int_reg_array_3_3_real;
  assign io_coef_out_payload_0_3_3_imag = int_reg_array_3_3_imag;
  assign io_coef_out_payload_0_3_4_real = int_reg_array_3_4_real;
  assign io_coef_out_payload_0_3_4_imag = int_reg_array_3_4_imag;
  assign io_coef_out_payload_0_3_5_real = int_reg_array_3_5_real;
  assign io_coef_out_payload_0_3_5_imag = int_reg_array_3_5_imag;
  assign io_coef_out_payload_0_3_6_real = int_reg_array_3_6_real;
  assign io_coef_out_payload_0_3_6_imag = int_reg_array_3_6_imag;
  assign io_coef_out_payload_0_3_7_real = int_reg_array_3_7_real;
  assign io_coef_out_payload_0_3_7_imag = int_reg_array_3_7_imag;
  assign io_coef_out_payload_0_3_8_real = int_reg_array_3_8_real;
  assign io_coef_out_payload_0_3_8_imag = int_reg_array_3_8_imag;
  assign io_coef_out_payload_0_3_9_real = int_reg_array_3_9_real;
  assign io_coef_out_payload_0_3_9_imag = int_reg_array_3_9_imag;
  assign io_coef_out_payload_0_3_10_real = int_reg_array_3_10_real;
  assign io_coef_out_payload_0_3_10_imag = int_reg_array_3_10_imag;
  assign io_coef_out_payload_0_3_11_real = int_reg_array_3_11_real;
  assign io_coef_out_payload_0_3_11_imag = int_reg_array_3_11_imag;
  assign io_coef_out_payload_0_3_12_real = int_reg_array_3_12_real;
  assign io_coef_out_payload_0_3_12_imag = int_reg_array_3_12_imag;
  assign io_coef_out_payload_0_3_13_real = int_reg_array_3_13_real;
  assign io_coef_out_payload_0_3_13_imag = int_reg_array_3_13_imag;
  assign io_coef_out_payload_0_3_14_real = int_reg_array_3_14_real;
  assign io_coef_out_payload_0_3_14_imag = int_reg_array_3_14_imag;
  assign io_coef_out_payload_0_3_15_real = int_reg_array_3_15_real;
  assign io_coef_out_payload_0_3_15_imag = int_reg_array_3_15_imag;
  assign io_coef_out_payload_0_3_16_real = int_reg_array_3_16_real;
  assign io_coef_out_payload_0_3_16_imag = int_reg_array_3_16_imag;
  assign io_coef_out_payload_0_3_17_real = int_reg_array_3_17_real;
  assign io_coef_out_payload_0_3_17_imag = int_reg_array_3_17_imag;
  assign io_coef_out_payload_0_3_18_real = int_reg_array_3_18_real;
  assign io_coef_out_payload_0_3_18_imag = int_reg_array_3_18_imag;
  assign io_coef_out_payload_0_3_19_real = int_reg_array_3_19_real;
  assign io_coef_out_payload_0_3_19_imag = int_reg_array_3_19_imag;
  assign io_coef_out_payload_0_3_20_real = int_reg_array_3_20_real;
  assign io_coef_out_payload_0_3_20_imag = int_reg_array_3_20_imag;
  assign io_coef_out_payload_0_3_21_real = int_reg_array_3_21_real;
  assign io_coef_out_payload_0_3_21_imag = int_reg_array_3_21_imag;
  assign io_coef_out_payload_0_3_22_real = int_reg_array_3_22_real;
  assign io_coef_out_payload_0_3_22_imag = int_reg_array_3_22_imag;
  assign io_coef_out_payload_0_3_23_real = int_reg_array_3_23_real;
  assign io_coef_out_payload_0_3_23_imag = int_reg_array_3_23_imag;
  assign io_coef_out_payload_0_3_24_real = int_reg_array_3_24_real;
  assign io_coef_out_payload_0_3_24_imag = int_reg_array_3_24_imag;
  assign io_coef_out_payload_0_3_25_real = int_reg_array_3_25_real;
  assign io_coef_out_payload_0_3_25_imag = int_reg_array_3_25_imag;
  assign io_coef_out_payload_0_3_26_real = int_reg_array_3_26_real;
  assign io_coef_out_payload_0_3_26_imag = int_reg_array_3_26_imag;
  assign io_coef_out_payload_0_3_27_real = int_reg_array_3_27_real;
  assign io_coef_out_payload_0_3_27_imag = int_reg_array_3_27_imag;
  assign io_coef_out_payload_0_3_28_real = int_reg_array_3_28_real;
  assign io_coef_out_payload_0_3_28_imag = int_reg_array_3_28_imag;
  assign io_coef_out_payload_0_3_29_real = int_reg_array_3_29_real;
  assign io_coef_out_payload_0_3_29_imag = int_reg_array_3_29_imag;
  assign io_coef_out_payload_0_3_30_real = int_reg_array_3_30_real;
  assign io_coef_out_payload_0_3_30_imag = int_reg_array_3_30_imag;
  assign io_coef_out_payload_0_3_31_real = int_reg_array_3_31_real;
  assign io_coef_out_payload_0_3_31_imag = int_reg_array_3_31_imag;
  assign io_coef_out_payload_0_3_32_real = int_reg_array_3_32_real;
  assign io_coef_out_payload_0_3_32_imag = int_reg_array_3_32_imag;
  assign io_coef_out_payload_0_3_33_real = int_reg_array_3_33_real;
  assign io_coef_out_payload_0_3_33_imag = int_reg_array_3_33_imag;
  assign io_coef_out_payload_0_3_34_real = int_reg_array_3_34_real;
  assign io_coef_out_payload_0_3_34_imag = int_reg_array_3_34_imag;
  assign io_coef_out_payload_0_3_35_real = int_reg_array_3_35_real;
  assign io_coef_out_payload_0_3_35_imag = int_reg_array_3_35_imag;
  assign io_coef_out_payload_0_3_36_real = int_reg_array_3_36_real;
  assign io_coef_out_payload_0_3_36_imag = int_reg_array_3_36_imag;
  assign io_coef_out_payload_0_3_37_real = int_reg_array_3_37_real;
  assign io_coef_out_payload_0_3_37_imag = int_reg_array_3_37_imag;
  assign io_coef_out_payload_0_3_38_real = int_reg_array_3_38_real;
  assign io_coef_out_payload_0_3_38_imag = int_reg_array_3_38_imag;
  assign io_coef_out_payload_0_3_39_real = int_reg_array_3_39_real;
  assign io_coef_out_payload_0_3_39_imag = int_reg_array_3_39_imag;
  assign io_coef_out_payload_0_3_40_real = int_reg_array_3_40_real;
  assign io_coef_out_payload_0_3_40_imag = int_reg_array_3_40_imag;
  assign io_coef_out_payload_0_3_41_real = int_reg_array_3_41_real;
  assign io_coef_out_payload_0_3_41_imag = int_reg_array_3_41_imag;
  assign io_coef_out_payload_0_3_42_real = int_reg_array_3_42_real;
  assign io_coef_out_payload_0_3_42_imag = int_reg_array_3_42_imag;
  assign io_coef_out_payload_0_3_43_real = int_reg_array_3_43_real;
  assign io_coef_out_payload_0_3_43_imag = int_reg_array_3_43_imag;
  assign io_coef_out_payload_0_3_44_real = int_reg_array_3_44_real;
  assign io_coef_out_payload_0_3_44_imag = int_reg_array_3_44_imag;
  assign io_coef_out_payload_0_3_45_real = int_reg_array_3_45_real;
  assign io_coef_out_payload_0_3_45_imag = int_reg_array_3_45_imag;
  assign io_coef_out_payload_0_3_46_real = int_reg_array_3_46_real;
  assign io_coef_out_payload_0_3_46_imag = int_reg_array_3_46_imag;
  assign io_coef_out_payload_0_3_47_real = int_reg_array_3_47_real;
  assign io_coef_out_payload_0_3_47_imag = int_reg_array_3_47_imag;
  assign io_coef_out_payload_0_3_48_real = int_reg_array_3_48_real;
  assign io_coef_out_payload_0_3_48_imag = int_reg_array_3_48_imag;
  assign io_coef_out_payload_0_3_49_real = int_reg_array_3_49_real;
  assign io_coef_out_payload_0_3_49_imag = int_reg_array_3_49_imag;
  assign io_coef_out_payload_0_4_0_real = int_reg_array_4_0_real;
  assign io_coef_out_payload_0_4_0_imag = int_reg_array_4_0_imag;
  assign io_coef_out_payload_0_4_1_real = int_reg_array_4_1_real;
  assign io_coef_out_payload_0_4_1_imag = int_reg_array_4_1_imag;
  assign io_coef_out_payload_0_4_2_real = int_reg_array_4_2_real;
  assign io_coef_out_payload_0_4_2_imag = int_reg_array_4_2_imag;
  assign io_coef_out_payload_0_4_3_real = int_reg_array_4_3_real;
  assign io_coef_out_payload_0_4_3_imag = int_reg_array_4_3_imag;
  assign io_coef_out_payload_0_4_4_real = int_reg_array_4_4_real;
  assign io_coef_out_payload_0_4_4_imag = int_reg_array_4_4_imag;
  assign io_coef_out_payload_0_4_5_real = int_reg_array_4_5_real;
  assign io_coef_out_payload_0_4_5_imag = int_reg_array_4_5_imag;
  assign io_coef_out_payload_0_4_6_real = int_reg_array_4_6_real;
  assign io_coef_out_payload_0_4_6_imag = int_reg_array_4_6_imag;
  assign io_coef_out_payload_0_4_7_real = int_reg_array_4_7_real;
  assign io_coef_out_payload_0_4_7_imag = int_reg_array_4_7_imag;
  assign io_coef_out_payload_0_4_8_real = int_reg_array_4_8_real;
  assign io_coef_out_payload_0_4_8_imag = int_reg_array_4_8_imag;
  assign io_coef_out_payload_0_4_9_real = int_reg_array_4_9_real;
  assign io_coef_out_payload_0_4_9_imag = int_reg_array_4_9_imag;
  assign io_coef_out_payload_0_4_10_real = int_reg_array_4_10_real;
  assign io_coef_out_payload_0_4_10_imag = int_reg_array_4_10_imag;
  assign io_coef_out_payload_0_4_11_real = int_reg_array_4_11_real;
  assign io_coef_out_payload_0_4_11_imag = int_reg_array_4_11_imag;
  assign io_coef_out_payload_0_4_12_real = int_reg_array_4_12_real;
  assign io_coef_out_payload_0_4_12_imag = int_reg_array_4_12_imag;
  assign io_coef_out_payload_0_4_13_real = int_reg_array_4_13_real;
  assign io_coef_out_payload_0_4_13_imag = int_reg_array_4_13_imag;
  assign io_coef_out_payload_0_4_14_real = int_reg_array_4_14_real;
  assign io_coef_out_payload_0_4_14_imag = int_reg_array_4_14_imag;
  assign io_coef_out_payload_0_4_15_real = int_reg_array_4_15_real;
  assign io_coef_out_payload_0_4_15_imag = int_reg_array_4_15_imag;
  assign io_coef_out_payload_0_4_16_real = int_reg_array_4_16_real;
  assign io_coef_out_payload_0_4_16_imag = int_reg_array_4_16_imag;
  assign io_coef_out_payload_0_4_17_real = int_reg_array_4_17_real;
  assign io_coef_out_payload_0_4_17_imag = int_reg_array_4_17_imag;
  assign io_coef_out_payload_0_4_18_real = int_reg_array_4_18_real;
  assign io_coef_out_payload_0_4_18_imag = int_reg_array_4_18_imag;
  assign io_coef_out_payload_0_4_19_real = int_reg_array_4_19_real;
  assign io_coef_out_payload_0_4_19_imag = int_reg_array_4_19_imag;
  assign io_coef_out_payload_0_4_20_real = int_reg_array_4_20_real;
  assign io_coef_out_payload_0_4_20_imag = int_reg_array_4_20_imag;
  assign io_coef_out_payload_0_4_21_real = int_reg_array_4_21_real;
  assign io_coef_out_payload_0_4_21_imag = int_reg_array_4_21_imag;
  assign io_coef_out_payload_0_4_22_real = int_reg_array_4_22_real;
  assign io_coef_out_payload_0_4_22_imag = int_reg_array_4_22_imag;
  assign io_coef_out_payload_0_4_23_real = int_reg_array_4_23_real;
  assign io_coef_out_payload_0_4_23_imag = int_reg_array_4_23_imag;
  assign io_coef_out_payload_0_4_24_real = int_reg_array_4_24_real;
  assign io_coef_out_payload_0_4_24_imag = int_reg_array_4_24_imag;
  assign io_coef_out_payload_0_4_25_real = int_reg_array_4_25_real;
  assign io_coef_out_payload_0_4_25_imag = int_reg_array_4_25_imag;
  assign io_coef_out_payload_0_4_26_real = int_reg_array_4_26_real;
  assign io_coef_out_payload_0_4_26_imag = int_reg_array_4_26_imag;
  assign io_coef_out_payload_0_4_27_real = int_reg_array_4_27_real;
  assign io_coef_out_payload_0_4_27_imag = int_reg_array_4_27_imag;
  assign io_coef_out_payload_0_4_28_real = int_reg_array_4_28_real;
  assign io_coef_out_payload_0_4_28_imag = int_reg_array_4_28_imag;
  assign io_coef_out_payload_0_4_29_real = int_reg_array_4_29_real;
  assign io_coef_out_payload_0_4_29_imag = int_reg_array_4_29_imag;
  assign io_coef_out_payload_0_4_30_real = int_reg_array_4_30_real;
  assign io_coef_out_payload_0_4_30_imag = int_reg_array_4_30_imag;
  assign io_coef_out_payload_0_4_31_real = int_reg_array_4_31_real;
  assign io_coef_out_payload_0_4_31_imag = int_reg_array_4_31_imag;
  assign io_coef_out_payload_0_4_32_real = int_reg_array_4_32_real;
  assign io_coef_out_payload_0_4_32_imag = int_reg_array_4_32_imag;
  assign io_coef_out_payload_0_4_33_real = int_reg_array_4_33_real;
  assign io_coef_out_payload_0_4_33_imag = int_reg_array_4_33_imag;
  assign io_coef_out_payload_0_4_34_real = int_reg_array_4_34_real;
  assign io_coef_out_payload_0_4_34_imag = int_reg_array_4_34_imag;
  assign io_coef_out_payload_0_4_35_real = int_reg_array_4_35_real;
  assign io_coef_out_payload_0_4_35_imag = int_reg_array_4_35_imag;
  assign io_coef_out_payload_0_4_36_real = int_reg_array_4_36_real;
  assign io_coef_out_payload_0_4_36_imag = int_reg_array_4_36_imag;
  assign io_coef_out_payload_0_4_37_real = int_reg_array_4_37_real;
  assign io_coef_out_payload_0_4_37_imag = int_reg_array_4_37_imag;
  assign io_coef_out_payload_0_4_38_real = int_reg_array_4_38_real;
  assign io_coef_out_payload_0_4_38_imag = int_reg_array_4_38_imag;
  assign io_coef_out_payload_0_4_39_real = int_reg_array_4_39_real;
  assign io_coef_out_payload_0_4_39_imag = int_reg_array_4_39_imag;
  assign io_coef_out_payload_0_4_40_real = int_reg_array_4_40_real;
  assign io_coef_out_payload_0_4_40_imag = int_reg_array_4_40_imag;
  assign io_coef_out_payload_0_4_41_real = int_reg_array_4_41_real;
  assign io_coef_out_payload_0_4_41_imag = int_reg_array_4_41_imag;
  assign io_coef_out_payload_0_4_42_real = int_reg_array_4_42_real;
  assign io_coef_out_payload_0_4_42_imag = int_reg_array_4_42_imag;
  assign io_coef_out_payload_0_4_43_real = int_reg_array_4_43_real;
  assign io_coef_out_payload_0_4_43_imag = int_reg_array_4_43_imag;
  assign io_coef_out_payload_0_4_44_real = int_reg_array_4_44_real;
  assign io_coef_out_payload_0_4_44_imag = int_reg_array_4_44_imag;
  assign io_coef_out_payload_0_4_45_real = int_reg_array_4_45_real;
  assign io_coef_out_payload_0_4_45_imag = int_reg_array_4_45_imag;
  assign io_coef_out_payload_0_4_46_real = int_reg_array_4_46_real;
  assign io_coef_out_payload_0_4_46_imag = int_reg_array_4_46_imag;
  assign io_coef_out_payload_0_4_47_real = int_reg_array_4_47_real;
  assign io_coef_out_payload_0_4_47_imag = int_reg_array_4_47_imag;
  assign io_coef_out_payload_0_4_48_real = int_reg_array_4_48_real;
  assign io_coef_out_payload_0_4_48_imag = int_reg_array_4_48_imag;
  assign io_coef_out_payload_0_4_49_real = int_reg_array_4_49_real;
  assign io_coef_out_payload_0_4_49_imag = int_reg_array_4_49_imag;
  assign io_coef_out_payload_0_5_0_real = int_reg_array_5_0_real;
  assign io_coef_out_payload_0_5_0_imag = int_reg_array_5_0_imag;
  assign io_coef_out_payload_0_5_1_real = int_reg_array_5_1_real;
  assign io_coef_out_payload_0_5_1_imag = int_reg_array_5_1_imag;
  assign io_coef_out_payload_0_5_2_real = int_reg_array_5_2_real;
  assign io_coef_out_payload_0_5_2_imag = int_reg_array_5_2_imag;
  assign io_coef_out_payload_0_5_3_real = int_reg_array_5_3_real;
  assign io_coef_out_payload_0_5_3_imag = int_reg_array_5_3_imag;
  assign io_coef_out_payload_0_5_4_real = int_reg_array_5_4_real;
  assign io_coef_out_payload_0_5_4_imag = int_reg_array_5_4_imag;
  assign io_coef_out_payload_0_5_5_real = int_reg_array_5_5_real;
  assign io_coef_out_payload_0_5_5_imag = int_reg_array_5_5_imag;
  assign io_coef_out_payload_0_5_6_real = int_reg_array_5_6_real;
  assign io_coef_out_payload_0_5_6_imag = int_reg_array_5_6_imag;
  assign io_coef_out_payload_0_5_7_real = int_reg_array_5_7_real;
  assign io_coef_out_payload_0_5_7_imag = int_reg_array_5_7_imag;
  assign io_coef_out_payload_0_5_8_real = int_reg_array_5_8_real;
  assign io_coef_out_payload_0_5_8_imag = int_reg_array_5_8_imag;
  assign io_coef_out_payload_0_5_9_real = int_reg_array_5_9_real;
  assign io_coef_out_payload_0_5_9_imag = int_reg_array_5_9_imag;
  assign io_coef_out_payload_0_5_10_real = int_reg_array_5_10_real;
  assign io_coef_out_payload_0_5_10_imag = int_reg_array_5_10_imag;
  assign io_coef_out_payload_0_5_11_real = int_reg_array_5_11_real;
  assign io_coef_out_payload_0_5_11_imag = int_reg_array_5_11_imag;
  assign io_coef_out_payload_0_5_12_real = int_reg_array_5_12_real;
  assign io_coef_out_payload_0_5_12_imag = int_reg_array_5_12_imag;
  assign io_coef_out_payload_0_5_13_real = int_reg_array_5_13_real;
  assign io_coef_out_payload_0_5_13_imag = int_reg_array_5_13_imag;
  assign io_coef_out_payload_0_5_14_real = int_reg_array_5_14_real;
  assign io_coef_out_payload_0_5_14_imag = int_reg_array_5_14_imag;
  assign io_coef_out_payload_0_5_15_real = int_reg_array_5_15_real;
  assign io_coef_out_payload_0_5_15_imag = int_reg_array_5_15_imag;
  assign io_coef_out_payload_0_5_16_real = int_reg_array_5_16_real;
  assign io_coef_out_payload_0_5_16_imag = int_reg_array_5_16_imag;
  assign io_coef_out_payload_0_5_17_real = int_reg_array_5_17_real;
  assign io_coef_out_payload_0_5_17_imag = int_reg_array_5_17_imag;
  assign io_coef_out_payload_0_5_18_real = int_reg_array_5_18_real;
  assign io_coef_out_payload_0_5_18_imag = int_reg_array_5_18_imag;
  assign io_coef_out_payload_0_5_19_real = int_reg_array_5_19_real;
  assign io_coef_out_payload_0_5_19_imag = int_reg_array_5_19_imag;
  assign io_coef_out_payload_0_5_20_real = int_reg_array_5_20_real;
  assign io_coef_out_payload_0_5_20_imag = int_reg_array_5_20_imag;
  assign io_coef_out_payload_0_5_21_real = int_reg_array_5_21_real;
  assign io_coef_out_payload_0_5_21_imag = int_reg_array_5_21_imag;
  assign io_coef_out_payload_0_5_22_real = int_reg_array_5_22_real;
  assign io_coef_out_payload_0_5_22_imag = int_reg_array_5_22_imag;
  assign io_coef_out_payload_0_5_23_real = int_reg_array_5_23_real;
  assign io_coef_out_payload_0_5_23_imag = int_reg_array_5_23_imag;
  assign io_coef_out_payload_0_5_24_real = int_reg_array_5_24_real;
  assign io_coef_out_payload_0_5_24_imag = int_reg_array_5_24_imag;
  assign io_coef_out_payload_0_5_25_real = int_reg_array_5_25_real;
  assign io_coef_out_payload_0_5_25_imag = int_reg_array_5_25_imag;
  assign io_coef_out_payload_0_5_26_real = int_reg_array_5_26_real;
  assign io_coef_out_payload_0_5_26_imag = int_reg_array_5_26_imag;
  assign io_coef_out_payload_0_5_27_real = int_reg_array_5_27_real;
  assign io_coef_out_payload_0_5_27_imag = int_reg_array_5_27_imag;
  assign io_coef_out_payload_0_5_28_real = int_reg_array_5_28_real;
  assign io_coef_out_payload_0_5_28_imag = int_reg_array_5_28_imag;
  assign io_coef_out_payload_0_5_29_real = int_reg_array_5_29_real;
  assign io_coef_out_payload_0_5_29_imag = int_reg_array_5_29_imag;
  assign io_coef_out_payload_0_5_30_real = int_reg_array_5_30_real;
  assign io_coef_out_payload_0_5_30_imag = int_reg_array_5_30_imag;
  assign io_coef_out_payload_0_5_31_real = int_reg_array_5_31_real;
  assign io_coef_out_payload_0_5_31_imag = int_reg_array_5_31_imag;
  assign io_coef_out_payload_0_5_32_real = int_reg_array_5_32_real;
  assign io_coef_out_payload_0_5_32_imag = int_reg_array_5_32_imag;
  assign io_coef_out_payload_0_5_33_real = int_reg_array_5_33_real;
  assign io_coef_out_payload_0_5_33_imag = int_reg_array_5_33_imag;
  assign io_coef_out_payload_0_5_34_real = int_reg_array_5_34_real;
  assign io_coef_out_payload_0_5_34_imag = int_reg_array_5_34_imag;
  assign io_coef_out_payload_0_5_35_real = int_reg_array_5_35_real;
  assign io_coef_out_payload_0_5_35_imag = int_reg_array_5_35_imag;
  assign io_coef_out_payload_0_5_36_real = int_reg_array_5_36_real;
  assign io_coef_out_payload_0_5_36_imag = int_reg_array_5_36_imag;
  assign io_coef_out_payload_0_5_37_real = int_reg_array_5_37_real;
  assign io_coef_out_payload_0_5_37_imag = int_reg_array_5_37_imag;
  assign io_coef_out_payload_0_5_38_real = int_reg_array_5_38_real;
  assign io_coef_out_payload_0_5_38_imag = int_reg_array_5_38_imag;
  assign io_coef_out_payload_0_5_39_real = int_reg_array_5_39_real;
  assign io_coef_out_payload_0_5_39_imag = int_reg_array_5_39_imag;
  assign io_coef_out_payload_0_5_40_real = int_reg_array_5_40_real;
  assign io_coef_out_payload_0_5_40_imag = int_reg_array_5_40_imag;
  assign io_coef_out_payload_0_5_41_real = int_reg_array_5_41_real;
  assign io_coef_out_payload_0_5_41_imag = int_reg_array_5_41_imag;
  assign io_coef_out_payload_0_5_42_real = int_reg_array_5_42_real;
  assign io_coef_out_payload_0_5_42_imag = int_reg_array_5_42_imag;
  assign io_coef_out_payload_0_5_43_real = int_reg_array_5_43_real;
  assign io_coef_out_payload_0_5_43_imag = int_reg_array_5_43_imag;
  assign io_coef_out_payload_0_5_44_real = int_reg_array_5_44_real;
  assign io_coef_out_payload_0_5_44_imag = int_reg_array_5_44_imag;
  assign io_coef_out_payload_0_5_45_real = int_reg_array_5_45_real;
  assign io_coef_out_payload_0_5_45_imag = int_reg_array_5_45_imag;
  assign io_coef_out_payload_0_5_46_real = int_reg_array_5_46_real;
  assign io_coef_out_payload_0_5_46_imag = int_reg_array_5_46_imag;
  assign io_coef_out_payload_0_5_47_real = int_reg_array_5_47_real;
  assign io_coef_out_payload_0_5_47_imag = int_reg_array_5_47_imag;
  assign io_coef_out_payload_0_5_48_real = int_reg_array_5_48_real;
  assign io_coef_out_payload_0_5_48_imag = int_reg_array_5_48_imag;
  assign io_coef_out_payload_0_5_49_real = int_reg_array_5_49_real;
  assign io_coef_out_payload_0_5_49_imag = int_reg_array_5_49_imag;
  assign io_coef_out_payload_0_6_0_real = int_reg_array_6_0_real;
  assign io_coef_out_payload_0_6_0_imag = int_reg_array_6_0_imag;
  assign io_coef_out_payload_0_6_1_real = int_reg_array_6_1_real;
  assign io_coef_out_payload_0_6_1_imag = int_reg_array_6_1_imag;
  assign io_coef_out_payload_0_6_2_real = int_reg_array_6_2_real;
  assign io_coef_out_payload_0_6_2_imag = int_reg_array_6_2_imag;
  assign io_coef_out_payload_0_6_3_real = int_reg_array_6_3_real;
  assign io_coef_out_payload_0_6_3_imag = int_reg_array_6_3_imag;
  assign io_coef_out_payload_0_6_4_real = int_reg_array_6_4_real;
  assign io_coef_out_payload_0_6_4_imag = int_reg_array_6_4_imag;
  assign io_coef_out_payload_0_6_5_real = int_reg_array_6_5_real;
  assign io_coef_out_payload_0_6_5_imag = int_reg_array_6_5_imag;
  assign io_coef_out_payload_0_6_6_real = int_reg_array_6_6_real;
  assign io_coef_out_payload_0_6_6_imag = int_reg_array_6_6_imag;
  assign io_coef_out_payload_0_6_7_real = int_reg_array_6_7_real;
  assign io_coef_out_payload_0_6_7_imag = int_reg_array_6_7_imag;
  assign io_coef_out_payload_0_6_8_real = int_reg_array_6_8_real;
  assign io_coef_out_payload_0_6_8_imag = int_reg_array_6_8_imag;
  assign io_coef_out_payload_0_6_9_real = int_reg_array_6_9_real;
  assign io_coef_out_payload_0_6_9_imag = int_reg_array_6_9_imag;
  assign io_coef_out_payload_0_6_10_real = int_reg_array_6_10_real;
  assign io_coef_out_payload_0_6_10_imag = int_reg_array_6_10_imag;
  assign io_coef_out_payload_0_6_11_real = int_reg_array_6_11_real;
  assign io_coef_out_payload_0_6_11_imag = int_reg_array_6_11_imag;
  assign io_coef_out_payload_0_6_12_real = int_reg_array_6_12_real;
  assign io_coef_out_payload_0_6_12_imag = int_reg_array_6_12_imag;
  assign io_coef_out_payload_0_6_13_real = int_reg_array_6_13_real;
  assign io_coef_out_payload_0_6_13_imag = int_reg_array_6_13_imag;
  assign io_coef_out_payload_0_6_14_real = int_reg_array_6_14_real;
  assign io_coef_out_payload_0_6_14_imag = int_reg_array_6_14_imag;
  assign io_coef_out_payload_0_6_15_real = int_reg_array_6_15_real;
  assign io_coef_out_payload_0_6_15_imag = int_reg_array_6_15_imag;
  assign io_coef_out_payload_0_6_16_real = int_reg_array_6_16_real;
  assign io_coef_out_payload_0_6_16_imag = int_reg_array_6_16_imag;
  assign io_coef_out_payload_0_6_17_real = int_reg_array_6_17_real;
  assign io_coef_out_payload_0_6_17_imag = int_reg_array_6_17_imag;
  assign io_coef_out_payload_0_6_18_real = int_reg_array_6_18_real;
  assign io_coef_out_payload_0_6_18_imag = int_reg_array_6_18_imag;
  assign io_coef_out_payload_0_6_19_real = int_reg_array_6_19_real;
  assign io_coef_out_payload_0_6_19_imag = int_reg_array_6_19_imag;
  assign io_coef_out_payload_0_6_20_real = int_reg_array_6_20_real;
  assign io_coef_out_payload_0_6_20_imag = int_reg_array_6_20_imag;
  assign io_coef_out_payload_0_6_21_real = int_reg_array_6_21_real;
  assign io_coef_out_payload_0_6_21_imag = int_reg_array_6_21_imag;
  assign io_coef_out_payload_0_6_22_real = int_reg_array_6_22_real;
  assign io_coef_out_payload_0_6_22_imag = int_reg_array_6_22_imag;
  assign io_coef_out_payload_0_6_23_real = int_reg_array_6_23_real;
  assign io_coef_out_payload_0_6_23_imag = int_reg_array_6_23_imag;
  assign io_coef_out_payload_0_6_24_real = int_reg_array_6_24_real;
  assign io_coef_out_payload_0_6_24_imag = int_reg_array_6_24_imag;
  assign io_coef_out_payload_0_6_25_real = int_reg_array_6_25_real;
  assign io_coef_out_payload_0_6_25_imag = int_reg_array_6_25_imag;
  assign io_coef_out_payload_0_6_26_real = int_reg_array_6_26_real;
  assign io_coef_out_payload_0_6_26_imag = int_reg_array_6_26_imag;
  assign io_coef_out_payload_0_6_27_real = int_reg_array_6_27_real;
  assign io_coef_out_payload_0_6_27_imag = int_reg_array_6_27_imag;
  assign io_coef_out_payload_0_6_28_real = int_reg_array_6_28_real;
  assign io_coef_out_payload_0_6_28_imag = int_reg_array_6_28_imag;
  assign io_coef_out_payload_0_6_29_real = int_reg_array_6_29_real;
  assign io_coef_out_payload_0_6_29_imag = int_reg_array_6_29_imag;
  assign io_coef_out_payload_0_6_30_real = int_reg_array_6_30_real;
  assign io_coef_out_payload_0_6_30_imag = int_reg_array_6_30_imag;
  assign io_coef_out_payload_0_6_31_real = int_reg_array_6_31_real;
  assign io_coef_out_payload_0_6_31_imag = int_reg_array_6_31_imag;
  assign io_coef_out_payload_0_6_32_real = int_reg_array_6_32_real;
  assign io_coef_out_payload_0_6_32_imag = int_reg_array_6_32_imag;
  assign io_coef_out_payload_0_6_33_real = int_reg_array_6_33_real;
  assign io_coef_out_payload_0_6_33_imag = int_reg_array_6_33_imag;
  assign io_coef_out_payload_0_6_34_real = int_reg_array_6_34_real;
  assign io_coef_out_payload_0_6_34_imag = int_reg_array_6_34_imag;
  assign io_coef_out_payload_0_6_35_real = int_reg_array_6_35_real;
  assign io_coef_out_payload_0_6_35_imag = int_reg_array_6_35_imag;
  assign io_coef_out_payload_0_6_36_real = int_reg_array_6_36_real;
  assign io_coef_out_payload_0_6_36_imag = int_reg_array_6_36_imag;
  assign io_coef_out_payload_0_6_37_real = int_reg_array_6_37_real;
  assign io_coef_out_payload_0_6_37_imag = int_reg_array_6_37_imag;
  assign io_coef_out_payload_0_6_38_real = int_reg_array_6_38_real;
  assign io_coef_out_payload_0_6_38_imag = int_reg_array_6_38_imag;
  assign io_coef_out_payload_0_6_39_real = int_reg_array_6_39_real;
  assign io_coef_out_payload_0_6_39_imag = int_reg_array_6_39_imag;
  assign io_coef_out_payload_0_6_40_real = int_reg_array_6_40_real;
  assign io_coef_out_payload_0_6_40_imag = int_reg_array_6_40_imag;
  assign io_coef_out_payload_0_6_41_real = int_reg_array_6_41_real;
  assign io_coef_out_payload_0_6_41_imag = int_reg_array_6_41_imag;
  assign io_coef_out_payload_0_6_42_real = int_reg_array_6_42_real;
  assign io_coef_out_payload_0_6_42_imag = int_reg_array_6_42_imag;
  assign io_coef_out_payload_0_6_43_real = int_reg_array_6_43_real;
  assign io_coef_out_payload_0_6_43_imag = int_reg_array_6_43_imag;
  assign io_coef_out_payload_0_6_44_real = int_reg_array_6_44_real;
  assign io_coef_out_payload_0_6_44_imag = int_reg_array_6_44_imag;
  assign io_coef_out_payload_0_6_45_real = int_reg_array_6_45_real;
  assign io_coef_out_payload_0_6_45_imag = int_reg_array_6_45_imag;
  assign io_coef_out_payload_0_6_46_real = int_reg_array_6_46_real;
  assign io_coef_out_payload_0_6_46_imag = int_reg_array_6_46_imag;
  assign io_coef_out_payload_0_6_47_real = int_reg_array_6_47_real;
  assign io_coef_out_payload_0_6_47_imag = int_reg_array_6_47_imag;
  assign io_coef_out_payload_0_6_48_real = int_reg_array_6_48_real;
  assign io_coef_out_payload_0_6_48_imag = int_reg_array_6_48_imag;
  assign io_coef_out_payload_0_6_49_real = int_reg_array_6_49_real;
  assign io_coef_out_payload_0_6_49_imag = int_reg_array_6_49_imag;
  assign io_coef_out_payload_0_7_0_real = int_reg_array_7_0_real;
  assign io_coef_out_payload_0_7_0_imag = int_reg_array_7_0_imag;
  assign io_coef_out_payload_0_7_1_real = int_reg_array_7_1_real;
  assign io_coef_out_payload_0_7_1_imag = int_reg_array_7_1_imag;
  assign io_coef_out_payload_0_7_2_real = int_reg_array_7_2_real;
  assign io_coef_out_payload_0_7_2_imag = int_reg_array_7_2_imag;
  assign io_coef_out_payload_0_7_3_real = int_reg_array_7_3_real;
  assign io_coef_out_payload_0_7_3_imag = int_reg_array_7_3_imag;
  assign io_coef_out_payload_0_7_4_real = int_reg_array_7_4_real;
  assign io_coef_out_payload_0_7_4_imag = int_reg_array_7_4_imag;
  assign io_coef_out_payload_0_7_5_real = int_reg_array_7_5_real;
  assign io_coef_out_payload_0_7_5_imag = int_reg_array_7_5_imag;
  assign io_coef_out_payload_0_7_6_real = int_reg_array_7_6_real;
  assign io_coef_out_payload_0_7_6_imag = int_reg_array_7_6_imag;
  assign io_coef_out_payload_0_7_7_real = int_reg_array_7_7_real;
  assign io_coef_out_payload_0_7_7_imag = int_reg_array_7_7_imag;
  assign io_coef_out_payload_0_7_8_real = int_reg_array_7_8_real;
  assign io_coef_out_payload_0_7_8_imag = int_reg_array_7_8_imag;
  assign io_coef_out_payload_0_7_9_real = int_reg_array_7_9_real;
  assign io_coef_out_payload_0_7_9_imag = int_reg_array_7_9_imag;
  assign io_coef_out_payload_0_7_10_real = int_reg_array_7_10_real;
  assign io_coef_out_payload_0_7_10_imag = int_reg_array_7_10_imag;
  assign io_coef_out_payload_0_7_11_real = int_reg_array_7_11_real;
  assign io_coef_out_payload_0_7_11_imag = int_reg_array_7_11_imag;
  assign io_coef_out_payload_0_7_12_real = int_reg_array_7_12_real;
  assign io_coef_out_payload_0_7_12_imag = int_reg_array_7_12_imag;
  assign io_coef_out_payload_0_7_13_real = int_reg_array_7_13_real;
  assign io_coef_out_payload_0_7_13_imag = int_reg_array_7_13_imag;
  assign io_coef_out_payload_0_7_14_real = int_reg_array_7_14_real;
  assign io_coef_out_payload_0_7_14_imag = int_reg_array_7_14_imag;
  assign io_coef_out_payload_0_7_15_real = int_reg_array_7_15_real;
  assign io_coef_out_payload_0_7_15_imag = int_reg_array_7_15_imag;
  assign io_coef_out_payload_0_7_16_real = int_reg_array_7_16_real;
  assign io_coef_out_payload_0_7_16_imag = int_reg_array_7_16_imag;
  assign io_coef_out_payload_0_7_17_real = int_reg_array_7_17_real;
  assign io_coef_out_payload_0_7_17_imag = int_reg_array_7_17_imag;
  assign io_coef_out_payload_0_7_18_real = int_reg_array_7_18_real;
  assign io_coef_out_payload_0_7_18_imag = int_reg_array_7_18_imag;
  assign io_coef_out_payload_0_7_19_real = int_reg_array_7_19_real;
  assign io_coef_out_payload_0_7_19_imag = int_reg_array_7_19_imag;
  assign io_coef_out_payload_0_7_20_real = int_reg_array_7_20_real;
  assign io_coef_out_payload_0_7_20_imag = int_reg_array_7_20_imag;
  assign io_coef_out_payload_0_7_21_real = int_reg_array_7_21_real;
  assign io_coef_out_payload_0_7_21_imag = int_reg_array_7_21_imag;
  assign io_coef_out_payload_0_7_22_real = int_reg_array_7_22_real;
  assign io_coef_out_payload_0_7_22_imag = int_reg_array_7_22_imag;
  assign io_coef_out_payload_0_7_23_real = int_reg_array_7_23_real;
  assign io_coef_out_payload_0_7_23_imag = int_reg_array_7_23_imag;
  assign io_coef_out_payload_0_7_24_real = int_reg_array_7_24_real;
  assign io_coef_out_payload_0_7_24_imag = int_reg_array_7_24_imag;
  assign io_coef_out_payload_0_7_25_real = int_reg_array_7_25_real;
  assign io_coef_out_payload_0_7_25_imag = int_reg_array_7_25_imag;
  assign io_coef_out_payload_0_7_26_real = int_reg_array_7_26_real;
  assign io_coef_out_payload_0_7_26_imag = int_reg_array_7_26_imag;
  assign io_coef_out_payload_0_7_27_real = int_reg_array_7_27_real;
  assign io_coef_out_payload_0_7_27_imag = int_reg_array_7_27_imag;
  assign io_coef_out_payload_0_7_28_real = int_reg_array_7_28_real;
  assign io_coef_out_payload_0_7_28_imag = int_reg_array_7_28_imag;
  assign io_coef_out_payload_0_7_29_real = int_reg_array_7_29_real;
  assign io_coef_out_payload_0_7_29_imag = int_reg_array_7_29_imag;
  assign io_coef_out_payload_0_7_30_real = int_reg_array_7_30_real;
  assign io_coef_out_payload_0_7_30_imag = int_reg_array_7_30_imag;
  assign io_coef_out_payload_0_7_31_real = int_reg_array_7_31_real;
  assign io_coef_out_payload_0_7_31_imag = int_reg_array_7_31_imag;
  assign io_coef_out_payload_0_7_32_real = int_reg_array_7_32_real;
  assign io_coef_out_payload_0_7_32_imag = int_reg_array_7_32_imag;
  assign io_coef_out_payload_0_7_33_real = int_reg_array_7_33_real;
  assign io_coef_out_payload_0_7_33_imag = int_reg_array_7_33_imag;
  assign io_coef_out_payload_0_7_34_real = int_reg_array_7_34_real;
  assign io_coef_out_payload_0_7_34_imag = int_reg_array_7_34_imag;
  assign io_coef_out_payload_0_7_35_real = int_reg_array_7_35_real;
  assign io_coef_out_payload_0_7_35_imag = int_reg_array_7_35_imag;
  assign io_coef_out_payload_0_7_36_real = int_reg_array_7_36_real;
  assign io_coef_out_payload_0_7_36_imag = int_reg_array_7_36_imag;
  assign io_coef_out_payload_0_7_37_real = int_reg_array_7_37_real;
  assign io_coef_out_payload_0_7_37_imag = int_reg_array_7_37_imag;
  assign io_coef_out_payload_0_7_38_real = int_reg_array_7_38_real;
  assign io_coef_out_payload_0_7_38_imag = int_reg_array_7_38_imag;
  assign io_coef_out_payload_0_7_39_real = int_reg_array_7_39_real;
  assign io_coef_out_payload_0_7_39_imag = int_reg_array_7_39_imag;
  assign io_coef_out_payload_0_7_40_real = int_reg_array_7_40_real;
  assign io_coef_out_payload_0_7_40_imag = int_reg_array_7_40_imag;
  assign io_coef_out_payload_0_7_41_real = int_reg_array_7_41_real;
  assign io_coef_out_payload_0_7_41_imag = int_reg_array_7_41_imag;
  assign io_coef_out_payload_0_7_42_real = int_reg_array_7_42_real;
  assign io_coef_out_payload_0_7_42_imag = int_reg_array_7_42_imag;
  assign io_coef_out_payload_0_7_43_real = int_reg_array_7_43_real;
  assign io_coef_out_payload_0_7_43_imag = int_reg_array_7_43_imag;
  assign io_coef_out_payload_0_7_44_real = int_reg_array_7_44_real;
  assign io_coef_out_payload_0_7_44_imag = int_reg_array_7_44_imag;
  assign io_coef_out_payload_0_7_45_real = int_reg_array_7_45_real;
  assign io_coef_out_payload_0_7_45_imag = int_reg_array_7_45_imag;
  assign io_coef_out_payload_0_7_46_real = int_reg_array_7_46_real;
  assign io_coef_out_payload_0_7_46_imag = int_reg_array_7_46_imag;
  assign io_coef_out_payload_0_7_47_real = int_reg_array_7_47_real;
  assign io_coef_out_payload_0_7_47_imag = int_reg_array_7_47_imag;
  assign io_coef_out_payload_0_7_48_real = int_reg_array_7_48_real;
  assign io_coef_out_payload_0_7_48_imag = int_reg_array_7_48_imag;
  assign io_coef_out_payload_0_7_49_real = int_reg_array_7_49_real;
  assign io_coef_out_payload_0_7_49_imag = int_reg_array_7_49_imag;
  assign io_coef_out_payload_0_8_0_real = int_reg_array_8_0_real;
  assign io_coef_out_payload_0_8_0_imag = int_reg_array_8_0_imag;
  assign io_coef_out_payload_0_8_1_real = int_reg_array_8_1_real;
  assign io_coef_out_payload_0_8_1_imag = int_reg_array_8_1_imag;
  assign io_coef_out_payload_0_8_2_real = int_reg_array_8_2_real;
  assign io_coef_out_payload_0_8_2_imag = int_reg_array_8_2_imag;
  assign io_coef_out_payload_0_8_3_real = int_reg_array_8_3_real;
  assign io_coef_out_payload_0_8_3_imag = int_reg_array_8_3_imag;
  assign io_coef_out_payload_0_8_4_real = int_reg_array_8_4_real;
  assign io_coef_out_payload_0_8_4_imag = int_reg_array_8_4_imag;
  assign io_coef_out_payload_0_8_5_real = int_reg_array_8_5_real;
  assign io_coef_out_payload_0_8_5_imag = int_reg_array_8_5_imag;
  assign io_coef_out_payload_0_8_6_real = int_reg_array_8_6_real;
  assign io_coef_out_payload_0_8_6_imag = int_reg_array_8_6_imag;
  assign io_coef_out_payload_0_8_7_real = int_reg_array_8_7_real;
  assign io_coef_out_payload_0_8_7_imag = int_reg_array_8_7_imag;
  assign io_coef_out_payload_0_8_8_real = int_reg_array_8_8_real;
  assign io_coef_out_payload_0_8_8_imag = int_reg_array_8_8_imag;
  assign io_coef_out_payload_0_8_9_real = int_reg_array_8_9_real;
  assign io_coef_out_payload_0_8_9_imag = int_reg_array_8_9_imag;
  assign io_coef_out_payload_0_8_10_real = int_reg_array_8_10_real;
  assign io_coef_out_payload_0_8_10_imag = int_reg_array_8_10_imag;
  assign io_coef_out_payload_0_8_11_real = int_reg_array_8_11_real;
  assign io_coef_out_payload_0_8_11_imag = int_reg_array_8_11_imag;
  assign io_coef_out_payload_0_8_12_real = int_reg_array_8_12_real;
  assign io_coef_out_payload_0_8_12_imag = int_reg_array_8_12_imag;
  assign io_coef_out_payload_0_8_13_real = int_reg_array_8_13_real;
  assign io_coef_out_payload_0_8_13_imag = int_reg_array_8_13_imag;
  assign io_coef_out_payload_0_8_14_real = int_reg_array_8_14_real;
  assign io_coef_out_payload_0_8_14_imag = int_reg_array_8_14_imag;
  assign io_coef_out_payload_0_8_15_real = int_reg_array_8_15_real;
  assign io_coef_out_payload_0_8_15_imag = int_reg_array_8_15_imag;
  assign io_coef_out_payload_0_8_16_real = int_reg_array_8_16_real;
  assign io_coef_out_payload_0_8_16_imag = int_reg_array_8_16_imag;
  assign io_coef_out_payload_0_8_17_real = int_reg_array_8_17_real;
  assign io_coef_out_payload_0_8_17_imag = int_reg_array_8_17_imag;
  assign io_coef_out_payload_0_8_18_real = int_reg_array_8_18_real;
  assign io_coef_out_payload_0_8_18_imag = int_reg_array_8_18_imag;
  assign io_coef_out_payload_0_8_19_real = int_reg_array_8_19_real;
  assign io_coef_out_payload_0_8_19_imag = int_reg_array_8_19_imag;
  assign io_coef_out_payload_0_8_20_real = int_reg_array_8_20_real;
  assign io_coef_out_payload_0_8_20_imag = int_reg_array_8_20_imag;
  assign io_coef_out_payload_0_8_21_real = int_reg_array_8_21_real;
  assign io_coef_out_payload_0_8_21_imag = int_reg_array_8_21_imag;
  assign io_coef_out_payload_0_8_22_real = int_reg_array_8_22_real;
  assign io_coef_out_payload_0_8_22_imag = int_reg_array_8_22_imag;
  assign io_coef_out_payload_0_8_23_real = int_reg_array_8_23_real;
  assign io_coef_out_payload_0_8_23_imag = int_reg_array_8_23_imag;
  assign io_coef_out_payload_0_8_24_real = int_reg_array_8_24_real;
  assign io_coef_out_payload_0_8_24_imag = int_reg_array_8_24_imag;
  assign io_coef_out_payload_0_8_25_real = int_reg_array_8_25_real;
  assign io_coef_out_payload_0_8_25_imag = int_reg_array_8_25_imag;
  assign io_coef_out_payload_0_8_26_real = int_reg_array_8_26_real;
  assign io_coef_out_payload_0_8_26_imag = int_reg_array_8_26_imag;
  assign io_coef_out_payload_0_8_27_real = int_reg_array_8_27_real;
  assign io_coef_out_payload_0_8_27_imag = int_reg_array_8_27_imag;
  assign io_coef_out_payload_0_8_28_real = int_reg_array_8_28_real;
  assign io_coef_out_payload_0_8_28_imag = int_reg_array_8_28_imag;
  assign io_coef_out_payload_0_8_29_real = int_reg_array_8_29_real;
  assign io_coef_out_payload_0_8_29_imag = int_reg_array_8_29_imag;
  assign io_coef_out_payload_0_8_30_real = int_reg_array_8_30_real;
  assign io_coef_out_payload_0_8_30_imag = int_reg_array_8_30_imag;
  assign io_coef_out_payload_0_8_31_real = int_reg_array_8_31_real;
  assign io_coef_out_payload_0_8_31_imag = int_reg_array_8_31_imag;
  assign io_coef_out_payload_0_8_32_real = int_reg_array_8_32_real;
  assign io_coef_out_payload_0_8_32_imag = int_reg_array_8_32_imag;
  assign io_coef_out_payload_0_8_33_real = int_reg_array_8_33_real;
  assign io_coef_out_payload_0_8_33_imag = int_reg_array_8_33_imag;
  assign io_coef_out_payload_0_8_34_real = int_reg_array_8_34_real;
  assign io_coef_out_payload_0_8_34_imag = int_reg_array_8_34_imag;
  assign io_coef_out_payload_0_8_35_real = int_reg_array_8_35_real;
  assign io_coef_out_payload_0_8_35_imag = int_reg_array_8_35_imag;
  assign io_coef_out_payload_0_8_36_real = int_reg_array_8_36_real;
  assign io_coef_out_payload_0_8_36_imag = int_reg_array_8_36_imag;
  assign io_coef_out_payload_0_8_37_real = int_reg_array_8_37_real;
  assign io_coef_out_payload_0_8_37_imag = int_reg_array_8_37_imag;
  assign io_coef_out_payload_0_8_38_real = int_reg_array_8_38_real;
  assign io_coef_out_payload_0_8_38_imag = int_reg_array_8_38_imag;
  assign io_coef_out_payload_0_8_39_real = int_reg_array_8_39_real;
  assign io_coef_out_payload_0_8_39_imag = int_reg_array_8_39_imag;
  assign io_coef_out_payload_0_8_40_real = int_reg_array_8_40_real;
  assign io_coef_out_payload_0_8_40_imag = int_reg_array_8_40_imag;
  assign io_coef_out_payload_0_8_41_real = int_reg_array_8_41_real;
  assign io_coef_out_payload_0_8_41_imag = int_reg_array_8_41_imag;
  assign io_coef_out_payload_0_8_42_real = int_reg_array_8_42_real;
  assign io_coef_out_payload_0_8_42_imag = int_reg_array_8_42_imag;
  assign io_coef_out_payload_0_8_43_real = int_reg_array_8_43_real;
  assign io_coef_out_payload_0_8_43_imag = int_reg_array_8_43_imag;
  assign io_coef_out_payload_0_8_44_real = int_reg_array_8_44_real;
  assign io_coef_out_payload_0_8_44_imag = int_reg_array_8_44_imag;
  assign io_coef_out_payload_0_8_45_real = int_reg_array_8_45_real;
  assign io_coef_out_payload_0_8_45_imag = int_reg_array_8_45_imag;
  assign io_coef_out_payload_0_8_46_real = int_reg_array_8_46_real;
  assign io_coef_out_payload_0_8_46_imag = int_reg_array_8_46_imag;
  assign io_coef_out_payload_0_8_47_real = int_reg_array_8_47_real;
  assign io_coef_out_payload_0_8_47_imag = int_reg_array_8_47_imag;
  assign io_coef_out_payload_0_8_48_real = int_reg_array_8_48_real;
  assign io_coef_out_payload_0_8_48_imag = int_reg_array_8_48_imag;
  assign io_coef_out_payload_0_8_49_real = int_reg_array_8_49_real;
  assign io_coef_out_payload_0_8_49_imag = int_reg_array_8_49_imag;
  assign io_coef_out_payload_0_9_0_real = int_reg_array_9_0_real;
  assign io_coef_out_payload_0_9_0_imag = int_reg_array_9_0_imag;
  assign io_coef_out_payload_0_9_1_real = int_reg_array_9_1_real;
  assign io_coef_out_payload_0_9_1_imag = int_reg_array_9_1_imag;
  assign io_coef_out_payload_0_9_2_real = int_reg_array_9_2_real;
  assign io_coef_out_payload_0_9_2_imag = int_reg_array_9_2_imag;
  assign io_coef_out_payload_0_9_3_real = int_reg_array_9_3_real;
  assign io_coef_out_payload_0_9_3_imag = int_reg_array_9_3_imag;
  assign io_coef_out_payload_0_9_4_real = int_reg_array_9_4_real;
  assign io_coef_out_payload_0_9_4_imag = int_reg_array_9_4_imag;
  assign io_coef_out_payload_0_9_5_real = int_reg_array_9_5_real;
  assign io_coef_out_payload_0_9_5_imag = int_reg_array_9_5_imag;
  assign io_coef_out_payload_0_9_6_real = int_reg_array_9_6_real;
  assign io_coef_out_payload_0_9_6_imag = int_reg_array_9_6_imag;
  assign io_coef_out_payload_0_9_7_real = int_reg_array_9_7_real;
  assign io_coef_out_payload_0_9_7_imag = int_reg_array_9_7_imag;
  assign io_coef_out_payload_0_9_8_real = int_reg_array_9_8_real;
  assign io_coef_out_payload_0_9_8_imag = int_reg_array_9_8_imag;
  assign io_coef_out_payload_0_9_9_real = int_reg_array_9_9_real;
  assign io_coef_out_payload_0_9_9_imag = int_reg_array_9_9_imag;
  assign io_coef_out_payload_0_9_10_real = int_reg_array_9_10_real;
  assign io_coef_out_payload_0_9_10_imag = int_reg_array_9_10_imag;
  assign io_coef_out_payload_0_9_11_real = int_reg_array_9_11_real;
  assign io_coef_out_payload_0_9_11_imag = int_reg_array_9_11_imag;
  assign io_coef_out_payload_0_9_12_real = int_reg_array_9_12_real;
  assign io_coef_out_payload_0_9_12_imag = int_reg_array_9_12_imag;
  assign io_coef_out_payload_0_9_13_real = int_reg_array_9_13_real;
  assign io_coef_out_payload_0_9_13_imag = int_reg_array_9_13_imag;
  assign io_coef_out_payload_0_9_14_real = int_reg_array_9_14_real;
  assign io_coef_out_payload_0_9_14_imag = int_reg_array_9_14_imag;
  assign io_coef_out_payload_0_9_15_real = int_reg_array_9_15_real;
  assign io_coef_out_payload_0_9_15_imag = int_reg_array_9_15_imag;
  assign io_coef_out_payload_0_9_16_real = int_reg_array_9_16_real;
  assign io_coef_out_payload_0_9_16_imag = int_reg_array_9_16_imag;
  assign io_coef_out_payload_0_9_17_real = int_reg_array_9_17_real;
  assign io_coef_out_payload_0_9_17_imag = int_reg_array_9_17_imag;
  assign io_coef_out_payload_0_9_18_real = int_reg_array_9_18_real;
  assign io_coef_out_payload_0_9_18_imag = int_reg_array_9_18_imag;
  assign io_coef_out_payload_0_9_19_real = int_reg_array_9_19_real;
  assign io_coef_out_payload_0_9_19_imag = int_reg_array_9_19_imag;
  assign io_coef_out_payload_0_9_20_real = int_reg_array_9_20_real;
  assign io_coef_out_payload_0_9_20_imag = int_reg_array_9_20_imag;
  assign io_coef_out_payload_0_9_21_real = int_reg_array_9_21_real;
  assign io_coef_out_payload_0_9_21_imag = int_reg_array_9_21_imag;
  assign io_coef_out_payload_0_9_22_real = int_reg_array_9_22_real;
  assign io_coef_out_payload_0_9_22_imag = int_reg_array_9_22_imag;
  assign io_coef_out_payload_0_9_23_real = int_reg_array_9_23_real;
  assign io_coef_out_payload_0_9_23_imag = int_reg_array_9_23_imag;
  assign io_coef_out_payload_0_9_24_real = int_reg_array_9_24_real;
  assign io_coef_out_payload_0_9_24_imag = int_reg_array_9_24_imag;
  assign io_coef_out_payload_0_9_25_real = int_reg_array_9_25_real;
  assign io_coef_out_payload_0_9_25_imag = int_reg_array_9_25_imag;
  assign io_coef_out_payload_0_9_26_real = int_reg_array_9_26_real;
  assign io_coef_out_payload_0_9_26_imag = int_reg_array_9_26_imag;
  assign io_coef_out_payload_0_9_27_real = int_reg_array_9_27_real;
  assign io_coef_out_payload_0_9_27_imag = int_reg_array_9_27_imag;
  assign io_coef_out_payload_0_9_28_real = int_reg_array_9_28_real;
  assign io_coef_out_payload_0_9_28_imag = int_reg_array_9_28_imag;
  assign io_coef_out_payload_0_9_29_real = int_reg_array_9_29_real;
  assign io_coef_out_payload_0_9_29_imag = int_reg_array_9_29_imag;
  assign io_coef_out_payload_0_9_30_real = int_reg_array_9_30_real;
  assign io_coef_out_payload_0_9_30_imag = int_reg_array_9_30_imag;
  assign io_coef_out_payload_0_9_31_real = int_reg_array_9_31_real;
  assign io_coef_out_payload_0_9_31_imag = int_reg_array_9_31_imag;
  assign io_coef_out_payload_0_9_32_real = int_reg_array_9_32_real;
  assign io_coef_out_payload_0_9_32_imag = int_reg_array_9_32_imag;
  assign io_coef_out_payload_0_9_33_real = int_reg_array_9_33_real;
  assign io_coef_out_payload_0_9_33_imag = int_reg_array_9_33_imag;
  assign io_coef_out_payload_0_9_34_real = int_reg_array_9_34_real;
  assign io_coef_out_payload_0_9_34_imag = int_reg_array_9_34_imag;
  assign io_coef_out_payload_0_9_35_real = int_reg_array_9_35_real;
  assign io_coef_out_payload_0_9_35_imag = int_reg_array_9_35_imag;
  assign io_coef_out_payload_0_9_36_real = int_reg_array_9_36_real;
  assign io_coef_out_payload_0_9_36_imag = int_reg_array_9_36_imag;
  assign io_coef_out_payload_0_9_37_real = int_reg_array_9_37_real;
  assign io_coef_out_payload_0_9_37_imag = int_reg_array_9_37_imag;
  assign io_coef_out_payload_0_9_38_real = int_reg_array_9_38_real;
  assign io_coef_out_payload_0_9_38_imag = int_reg_array_9_38_imag;
  assign io_coef_out_payload_0_9_39_real = int_reg_array_9_39_real;
  assign io_coef_out_payload_0_9_39_imag = int_reg_array_9_39_imag;
  assign io_coef_out_payload_0_9_40_real = int_reg_array_9_40_real;
  assign io_coef_out_payload_0_9_40_imag = int_reg_array_9_40_imag;
  assign io_coef_out_payload_0_9_41_real = int_reg_array_9_41_real;
  assign io_coef_out_payload_0_9_41_imag = int_reg_array_9_41_imag;
  assign io_coef_out_payload_0_9_42_real = int_reg_array_9_42_real;
  assign io_coef_out_payload_0_9_42_imag = int_reg_array_9_42_imag;
  assign io_coef_out_payload_0_9_43_real = int_reg_array_9_43_real;
  assign io_coef_out_payload_0_9_43_imag = int_reg_array_9_43_imag;
  assign io_coef_out_payload_0_9_44_real = int_reg_array_9_44_real;
  assign io_coef_out_payload_0_9_44_imag = int_reg_array_9_44_imag;
  assign io_coef_out_payload_0_9_45_real = int_reg_array_9_45_real;
  assign io_coef_out_payload_0_9_45_imag = int_reg_array_9_45_imag;
  assign io_coef_out_payload_0_9_46_real = int_reg_array_9_46_real;
  assign io_coef_out_payload_0_9_46_imag = int_reg_array_9_46_imag;
  assign io_coef_out_payload_0_9_47_real = int_reg_array_9_47_real;
  assign io_coef_out_payload_0_9_47_imag = int_reg_array_9_47_imag;
  assign io_coef_out_payload_0_9_48_real = int_reg_array_9_48_real;
  assign io_coef_out_payload_0_9_48_imag = int_reg_array_9_48_imag;
  assign io_coef_out_payload_0_9_49_real = int_reg_array_9_49_real;
  assign io_coef_out_payload_0_9_49_imag = int_reg_array_9_49_imag;
  assign io_coef_out_payload_0_10_0_real = int_reg_array_10_0_real;
  assign io_coef_out_payload_0_10_0_imag = int_reg_array_10_0_imag;
  assign io_coef_out_payload_0_10_1_real = int_reg_array_10_1_real;
  assign io_coef_out_payload_0_10_1_imag = int_reg_array_10_1_imag;
  assign io_coef_out_payload_0_10_2_real = int_reg_array_10_2_real;
  assign io_coef_out_payload_0_10_2_imag = int_reg_array_10_2_imag;
  assign io_coef_out_payload_0_10_3_real = int_reg_array_10_3_real;
  assign io_coef_out_payload_0_10_3_imag = int_reg_array_10_3_imag;
  assign io_coef_out_payload_0_10_4_real = int_reg_array_10_4_real;
  assign io_coef_out_payload_0_10_4_imag = int_reg_array_10_4_imag;
  assign io_coef_out_payload_0_10_5_real = int_reg_array_10_5_real;
  assign io_coef_out_payload_0_10_5_imag = int_reg_array_10_5_imag;
  assign io_coef_out_payload_0_10_6_real = int_reg_array_10_6_real;
  assign io_coef_out_payload_0_10_6_imag = int_reg_array_10_6_imag;
  assign io_coef_out_payload_0_10_7_real = int_reg_array_10_7_real;
  assign io_coef_out_payload_0_10_7_imag = int_reg_array_10_7_imag;
  assign io_coef_out_payload_0_10_8_real = int_reg_array_10_8_real;
  assign io_coef_out_payload_0_10_8_imag = int_reg_array_10_8_imag;
  assign io_coef_out_payload_0_10_9_real = int_reg_array_10_9_real;
  assign io_coef_out_payload_0_10_9_imag = int_reg_array_10_9_imag;
  assign io_coef_out_payload_0_10_10_real = int_reg_array_10_10_real;
  assign io_coef_out_payload_0_10_10_imag = int_reg_array_10_10_imag;
  assign io_coef_out_payload_0_10_11_real = int_reg_array_10_11_real;
  assign io_coef_out_payload_0_10_11_imag = int_reg_array_10_11_imag;
  assign io_coef_out_payload_0_10_12_real = int_reg_array_10_12_real;
  assign io_coef_out_payload_0_10_12_imag = int_reg_array_10_12_imag;
  assign io_coef_out_payload_0_10_13_real = int_reg_array_10_13_real;
  assign io_coef_out_payload_0_10_13_imag = int_reg_array_10_13_imag;
  assign io_coef_out_payload_0_10_14_real = int_reg_array_10_14_real;
  assign io_coef_out_payload_0_10_14_imag = int_reg_array_10_14_imag;
  assign io_coef_out_payload_0_10_15_real = int_reg_array_10_15_real;
  assign io_coef_out_payload_0_10_15_imag = int_reg_array_10_15_imag;
  assign io_coef_out_payload_0_10_16_real = int_reg_array_10_16_real;
  assign io_coef_out_payload_0_10_16_imag = int_reg_array_10_16_imag;
  assign io_coef_out_payload_0_10_17_real = int_reg_array_10_17_real;
  assign io_coef_out_payload_0_10_17_imag = int_reg_array_10_17_imag;
  assign io_coef_out_payload_0_10_18_real = int_reg_array_10_18_real;
  assign io_coef_out_payload_0_10_18_imag = int_reg_array_10_18_imag;
  assign io_coef_out_payload_0_10_19_real = int_reg_array_10_19_real;
  assign io_coef_out_payload_0_10_19_imag = int_reg_array_10_19_imag;
  assign io_coef_out_payload_0_10_20_real = int_reg_array_10_20_real;
  assign io_coef_out_payload_0_10_20_imag = int_reg_array_10_20_imag;
  assign io_coef_out_payload_0_10_21_real = int_reg_array_10_21_real;
  assign io_coef_out_payload_0_10_21_imag = int_reg_array_10_21_imag;
  assign io_coef_out_payload_0_10_22_real = int_reg_array_10_22_real;
  assign io_coef_out_payload_0_10_22_imag = int_reg_array_10_22_imag;
  assign io_coef_out_payload_0_10_23_real = int_reg_array_10_23_real;
  assign io_coef_out_payload_0_10_23_imag = int_reg_array_10_23_imag;
  assign io_coef_out_payload_0_10_24_real = int_reg_array_10_24_real;
  assign io_coef_out_payload_0_10_24_imag = int_reg_array_10_24_imag;
  assign io_coef_out_payload_0_10_25_real = int_reg_array_10_25_real;
  assign io_coef_out_payload_0_10_25_imag = int_reg_array_10_25_imag;
  assign io_coef_out_payload_0_10_26_real = int_reg_array_10_26_real;
  assign io_coef_out_payload_0_10_26_imag = int_reg_array_10_26_imag;
  assign io_coef_out_payload_0_10_27_real = int_reg_array_10_27_real;
  assign io_coef_out_payload_0_10_27_imag = int_reg_array_10_27_imag;
  assign io_coef_out_payload_0_10_28_real = int_reg_array_10_28_real;
  assign io_coef_out_payload_0_10_28_imag = int_reg_array_10_28_imag;
  assign io_coef_out_payload_0_10_29_real = int_reg_array_10_29_real;
  assign io_coef_out_payload_0_10_29_imag = int_reg_array_10_29_imag;
  assign io_coef_out_payload_0_10_30_real = int_reg_array_10_30_real;
  assign io_coef_out_payload_0_10_30_imag = int_reg_array_10_30_imag;
  assign io_coef_out_payload_0_10_31_real = int_reg_array_10_31_real;
  assign io_coef_out_payload_0_10_31_imag = int_reg_array_10_31_imag;
  assign io_coef_out_payload_0_10_32_real = int_reg_array_10_32_real;
  assign io_coef_out_payload_0_10_32_imag = int_reg_array_10_32_imag;
  assign io_coef_out_payload_0_10_33_real = int_reg_array_10_33_real;
  assign io_coef_out_payload_0_10_33_imag = int_reg_array_10_33_imag;
  assign io_coef_out_payload_0_10_34_real = int_reg_array_10_34_real;
  assign io_coef_out_payload_0_10_34_imag = int_reg_array_10_34_imag;
  assign io_coef_out_payload_0_10_35_real = int_reg_array_10_35_real;
  assign io_coef_out_payload_0_10_35_imag = int_reg_array_10_35_imag;
  assign io_coef_out_payload_0_10_36_real = int_reg_array_10_36_real;
  assign io_coef_out_payload_0_10_36_imag = int_reg_array_10_36_imag;
  assign io_coef_out_payload_0_10_37_real = int_reg_array_10_37_real;
  assign io_coef_out_payload_0_10_37_imag = int_reg_array_10_37_imag;
  assign io_coef_out_payload_0_10_38_real = int_reg_array_10_38_real;
  assign io_coef_out_payload_0_10_38_imag = int_reg_array_10_38_imag;
  assign io_coef_out_payload_0_10_39_real = int_reg_array_10_39_real;
  assign io_coef_out_payload_0_10_39_imag = int_reg_array_10_39_imag;
  assign io_coef_out_payload_0_10_40_real = int_reg_array_10_40_real;
  assign io_coef_out_payload_0_10_40_imag = int_reg_array_10_40_imag;
  assign io_coef_out_payload_0_10_41_real = int_reg_array_10_41_real;
  assign io_coef_out_payload_0_10_41_imag = int_reg_array_10_41_imag;
  assign io_coef_out_payload_0_10_42_real = int_reg_array_10_42_real;
  assign io_coef_out_payload_0_10_42_imag = int_reg_array_10_42_imag;
  assign io_coef_out_payload_0_10_43_real = int_reg_array_10_43_real;
  assign io_coef_out_payload_0_10_43_imag = int_reg_array_10_43_imag;
  assign io_coef_out_payload_0_10_44_real = int_reg_array_10_44_real;
  assign io_coef_out_payload_0_10_44_imag = int_reg_array_10_44_imag;
  assign io_coef_out_payload_0_10_45_real = int_reg_array_10_45_real;
  assign io_coef_out_payload_0_10_45_imag = int_reg_array_10_45_imag;
  assign io_coef_out_payload_0_10_46_real = int_reg_array_10_46_real;
  assign io_coef_out_payload_0_10_46_imag = int_reg_array_10_46_imag;
  assign io_coef_out_payload_0_10_47_real = int_reg_array_10_47_real;
  assign io_coef_out_payload_0_10_47_imag = int_reg_array_10_47_imag;
  assign io_coef_out_payload_0_10_48_real = int_reg_array_10_48_real;
  assign io_coef_out_payload_0_10_48_imag = int_reg_array_10_48_imag;
  assign io_coef_out_payload_0_10_49_real = int_reg_array_10_49_real;
  assign io_coef_out_payload_0_10_49_imag = int_reg_array_10_49_imag;
  assign io_coef_out_payload_0_11_0_real = int_reg_array_11_0_real;
  assign io_coef_out_payload_0_11_0_imag = int_reg_array_11_0_imag;
  assign io_coef_out_payload_0_11_1_real = int_reg_array_11_1_real;
  assign io_coef_out_payload_0_11_1_imag = int_reg_array_11_1_imag;
  assign io_coef_out_payload_0_11_2_real = int_reg_array_11_2_real;
  assign io_coef_out_payload_0_11_2_imag = int_reg_array_11_2_imag;
  assign io_coef_out_payload_0_11_3_real = int_reg_array_11_3_real;
  assign io_coef_out_payload_0_11_3_imag = int_reg_array_11_3_imag;
  assign io_coef_out_payload_0_11_4_real = int_reg_array_11_4_real;
  assign io_coef_out_payload_0_11_4_imag = int_reg_array_11_4_imag;
  assign io_coef_out_payload_0_11_5_real = int_reg_array_11_5_real;
  assign io_coef_out_payload_0_11_5_imag = int_reg_array_11_5_imag;
  assign io_coef_out_payload_0_11_6_real = int_reg_array_11_6_real;
  assign io_coef_out_payload_0_11_6_imag = int_reg_array_11_6_imag;
  assign io_coef_out_payload_0_11_7_real = int_reg_array_11_7_real;
  assign io_coef_out_payload_0_11_7_imag = int_reg_array_11_7_imag;
  assign io_coef_out_payload_0_11_8_real = int_reg_array_11_8_real;
  assign io_coef_out_payload_0_11_8_imag = int_reg_array_11_8_imag;
  assign io_coef_out_payload_0_11_9_real = int_reg_array_11_9_real;
  assign io_coef_out_payload_0_11_9_imag = int_reg_array_11_9_imag;
  assign io_coef_out_payload_0_11_10_real = int_reg_array_11_10_real;
  assign io_coef_out_payload_0_11_10_imag = int_reg_array_11_10_imag;
  assign io_coef_out_payload_0_11_11_real = int_reg_array_11_11_real;
  assign io_coef_out_payload_0_11_11_imag = int_reg_array_11_11_imag;
  assign io_coef_out_payload_0_11_12_real = int_reg_array_11_12_real;
  assign io_coef_out_payload_0_11_12_imag = int_reg_array_11_12_imag;
  assign io_coef_out_payload_0_11_13_real = int_reg_array_11_13_real;
  assign io_coef_out_payload_0_11_13_imag = int_reg_array_11_13_imag;
  assign io_coef_out_payload_0_11_14_real = int_reg_array_11_14_real;
  assign io_coef_out_payload_0_11_14_imag = int_reg_array_11_14_imag;
  assign io_coef_out_payload_0_11_15_real = int_reg_array_11_15_real;
  assign io_coef_out_payload_0_11_15_imag = int_reg_array_11_15_imag;
  assign io_coef_out_payload_0_11_16_real = int_reg_array_11_16_real;
  assign io_coef_out_payload_0_11_16_imag = int_reg_array_11_16_imag;
  assign io_coef_out_payload_0_11_17_real = int_reg_array_11_17_real;
  assign io_coef_out_payload_0_11_17_imag = int_reg_array_11_17_imag;
  assign io_coef_out_payload_0_11_18_real = int_reg_array_11_18_real;
  assign io_coef_out_payload_0_11_18_imag = int_reg_array_11_18_imag;
  assign io_coef_out_payload_0_11_19_real = int_reg_array_11_19_real;
  assign io_coef_out_payload_0_11_19_imag = int_reg_array_11_19_imag;
  assign io_coef_out_payload_0_11_20_real = int_reg_array_11_20_real;
  assign io_coef_out_payload_0_11_20_imag = int_reg_array_11_20_imag;
  assign io_coef_out_payload_0_11_21_real = int_reg_array_11_21_real;
  assign io_coef_out_payload_0_11_21_imag = int_reg_array_11_21_imag;
  assign io_coef_out_payload_0_11_22_real = int_reg_array_11_22_real;
  assign io_coef_out_payload_0_11_22_imag = int_reg_array_11_22_imag;
  assign io_coef_out_payload_0_11_23_real = int_reg_array_11_23_real;
  assign io_coef_out_payload_0_11_23_imag = int_reg_array_11_23_imag;
  assign io_coef_out_payload_0_11_24_real = int_reg_array_11_24_real;
  assign io_coef_out_payload_0_11_24_imag = int_reg_array_11_24_imag;
  assign io_coef_out_payload_0_11_25_real = int_reg_array_11_25_real;
  assign io_coef_out_payload_0_11_25_imag = int_reg_array_11_25_imag;
  assign io_coef_out_payload_0_11_26_real = int_reg_array_11_26_real;
  assign io_coef_out_payload_0_11_26_imag = int_reg_array_11_26_imag;
  assign io_coef_out_payload_0_11_27_real = int_reg_array_11_27_real;
  assign io_coef_out_payload_0_11_27_imag = int_reg_array_11_27_imag;
  assign io_coef_out_payload_0_11_28_real = int_reg_array_11_28_real;
  assign io_coef_out_payload_0_11_28_imag = int_reg_array_11_28_imag;
  assign io_coef_out_payload_0_11_29_real = int_reg_array_11_29_real;
  assign io_coef_out_payload_0_11_29_imag = int_reg_array_11_29_imag;
  assign io_coef_out_payload_0_11_30_real = int_reg_array_11_30_real;
  assign io_coef_out_payload_0_11_30_imag = int_reg_array_11_30_imag;
  assign io_coef_out_payload_0_11_31_real = int_reg_array_11_31_real;
  assign io_coef_out_payload_0_11_31_imag = int_reg_array_11_31_imag;
  assign io_coef_out_payload_0_11_32_real = int_reg_array_11_32_real;
  assign io_coef_out_payload_0_11_32_imag = int_reg_array_11_32_imag;
  assign io_coef_out_payload_0_11_33_real = int_reg_array_11_33_real;
  assign io_coef_out_payload_0_11_33_imag = int_reg_array_11_33_imag;
  assign io_coef_out_payload_0_11_34_real = int_reg_array_11_34_real;
  assign io_coef_out_payload_0_11_34_imag = int_reg_array_11_34_imag;
  assign io_coef_out_payload_0_11_35_real = int_reg_array_11_35_real;
  assign io_coef_out_payload_0_11_35_imag = int_reg_array_11_35_imag;
  assign io_coef_out_payload_0_11_36_real = int_reg_array_11_36_real;
  assign io_coef_out_payload_0_11_36_imag = int_reg_array_11_36_imag;
  assign io_coef_out_payload_0_11_37_real = int_reg_array_11_37_real;
  assign io_coef_out_payload_0_11_37_imag = int_reg_array_11_37_imag;
  assign io_coef_out_payload_0_11_38_real = int_reg_array_11_38_real;
  assign io_coef_out_payload_0_11_38_imag = int_reg_array_11_38_imag;
  assign io_coef_out_payload_0_11_39_real = int_reg_array_11_39_real;
  assign io_coef_out_payload_0_11_39_imag = int_reg_array_11_39_imag;
  assign io_coef_out_payload_0_11_40_real = int_reg_array_11_40_real;
  assign io_coef_out_payload_0_11_40_imag = int_reg_array_11_40_imag;
  assign io_coef_out_payload_0_11_41_real = int_reg_array_11_41_real;
  assign io_coef_out_payload_0_11_41_imag = int_reg_array_11_41_imag;
  assign io_coef_out_payload_0_11_42_real = int_reg_array_11_42_real;
  assign io_coef_out_payload_0_11_42_imag = int_reg_array_11_42_imag;
  assign io_coef_out_payload_0_11_43_real = int_reg_array_11_43_real;
  assign io_coef_out_payload_0_11_43_imag = int_reg_array_11_43_imag;
  assign io_coef_out_payload_0_11_44_real = int_reg_array_11_44_real;
  assign io_coef_out_payload_0_11_44_imag = int_reg_array_11_44_imag;
  assign io_coef_out_payload_0_11_45_real = int_reg_array_11_45_real;
  assign io_coef_out_payload_0_11_45_imag = int_reg_array_11_45_imag;
  assign io_coef_out_payload_0_11_46_real = int_reg_array_11_46_real;
  assign io_coef_out_payload_0_11_46_imag = int_reg_array_11_46_imag;
  assign io_coef_out_payload_0_11_47_real = int_reg_array_11_47_real;
  assign io_coef_out_payload_0_11_47_imag = int_reg_array_11_47_imag;
  assign io_coef_out_payload_0_11_48_real = int_reg_array_11_48_real;
  assign io_coef_out_payload_0_11_48_imag = int_reg_array_11_48_imag;
  assign io_coef_out_payload_0_11_49_real = int_reg_array_11_49_real;
  assign io_coef_out_payload_0_11_49_imag = int_reg_array_11_49_imag;
  assign io_coef_out_payload_0_12_0_real = int_reg_array_12_0_real;
  assign io_coef_out_payload_0_12_0_imag = int_reg_array_12_0_imag;
  assign io_coef_out_payload_0_12_1_real = int_reg_array_12_1_real;
  assign io_coef_out_payload_0_12_1_imag = int_reg_array_12_1_imag;
  assign io_coef_out_payload_0_12_2_real = int_reg_array_12_2_real;
  assign io_coef_out_payload_0_12_2_imag = int_reg_array_12_2_imag;
  assign io_coef_out_payload_0_12_3_real = int_reg_array_12_3_real;
  assign io_coef_out_payload_0_12_3_imag = int_reg_array_12_3_imag;
  assign io_coef_out_payload_0_12_4_real = int_reg_array_12_4_real;
  assign io_coef_out_payload_0_12_4_imag = int_reg_array_12_4_imag;
  assign io_coef_out_payload_0_12_5_real = int_reg_array_12_5_real;
  assign io_coef_out_payload_0_12_5_imag = int_reg_array_12_5_imag;
  assign io_coef_out_payload_0_12_6_real = int_reg_array_12_6_real;
  assign io_coef_out_payload_0_12_6_imag = int_reg_array_12_6_imag;
  assign io_coef_out_payload_0_12_7_real = int_reg_array_12_7_real;
  assign io_coef_out_payload_0_12_7_imag = int_reg_array_12_7_imag;
  assign io_coef_out_payload_0_12_8_real = int_reg_array_12_8_real;
  assign io_coef_out_payload_0_12_8_imag = int_reg_array_12_8_imag;
  assign io_coef_out_payload_0_12_9_real = int_reg_array_12_9_real;
  assign io_coef_out_payload_0_12_9_imag = int_reg_array_12_9_imag;
  assign io_coef_out_payload_0_12_10_real = int_reg_array_12_10_real;
  assign io_coef_out_payload_0_12_10_imag = int_reg_array_12_10_imag;
  assign io_coef_out_payload_0_12_11_real = int_reg_array_12_11_real;
  assign io_coef_out_payload_0_12_11_imag = int_reg_array_12_11_imag;
  assign io_coef_out_payload_0_12_12_real = int_reg_array_12_12_real;
  assign io_coef_out_payload_0_12_12_imag = int_reg_array_12_12_imag;
  assign io_coef_out_payload_0_12_13_real = int_reg_array_12_13_real;
  assign io_coef_out_payload_0_12_13_imag = int_reg_array_12_13_imag;
  assign io_coef_out_payload_0_12_14_real = int_reg_array_12_14_real;
  assign io_coef_out_payload_0_12_14_imag = int_reg_array_12_14_imag;
  assign io_coef_out_payload_0_12_15_real = int_reg_array_12_15_real;
  assign io_coef_out_payload_0_12_15_imag = int_reg_array_12_15_imag;
  assign io_coef_out_payload_0_12_16_real = int_reg_array_12_16_real;
  assign io_coef_out_payload_0_12_16_imag = int_reg_array_12_16_imag;
  assign io_coef_out_payload_0_12_17_real = int_reg_array_12_17_real;
  assign io_coef_out_payload_0_12_17_imag = int_reg_array_12_17_imag;
  assign io_coef_out_payload_0_12_18_real = int_reg_array_12_18_real;
  assign io_coef_out_payload_0_12_18_imag = int_reg_array_12_18_imag;
  assign io_coef_out_payload_0_12_19_real = int_reg_array_12_19_real;
  assign io_coef_out_payload_0_12_19_imag = int_reg_array_12_19_imag;
  assign io_coef_out_payload_0_12_20_real = int_reg_array_12_20_real;
  assign io_coef_out_payload_0_12_20_imag = int_reg_array_12_20_imag;
  assign io_coef_out_payload_0_12_21_real = int_reg_array_12_21_real;
  assign io_coef_out_payload_0_12_21_imag = int_reg_array_12_21_imag;
  assign io_coef_out_payload_0_12_22_real = int_reg_array_12_22_real;
  assign io_coef_out_payload_0_12_22_imag = int_reg_array_12_22_imag;
  assign io_coef_out_payload_0_12_23_real = int_reg_array_12_23_real;
  assign io_coef_out_payload_0_12_23_imag = int_reg_array_12_23_imag;
  assign io_coef_out_payload_0_12_24_real = int_reg_array_12_24_real;
  assign io_coef_out_payload_0_12_24_imag = int_reg_array_12_24_imag;
  assign io_coef_out_payload_0_12_25_real = int_reg_array_12_25_real;
  assign io_coef_out_payload_0_12_25_imag = int_reg_array_12_25_imag;
  assign io_coef_out_payload_0_12_26_real = int_reg_array_12_26_real;
  assign io_coef_out_payload_0_12_26_imag = int_reg_array_12_26_imag;
  assign io_coef_out_payload_0_12_27_real = int_reg_array_12_27_real;
  assign io_coef_out_payload_0_12_27_imag = int_reg_array_12_27_imag;
  assign io_coef_out_payload_0_12_28_real = int_reg_array_12_28_real;
  assign io_coef_out_payload_0_12_28_imag = int_reg_array_12_28_imag;
  assign io_coef_out_payload_0_12_29_real = int_reg_array_12_29_real;
  assign io_coef_out_payload_0_12_29_imag = int_reg_array_12_29_imag;
  assign io_coef_out_payload_0_12_30_real = int_reg_array_12_30_real;
  assign io_coef_out_payload_0_12_30_imag = int_reg_array_12_30_imag;
  assign io_coef_out_payload_0_12_31_real = int_reg_array_12_31_real;
  assign io_coef_out_payload_0_12_31_imag = int_reg_array_12_31_imag;
  assign io_coef_out_payload_0_12_32_real = int_reg_array_12_32_real;
  assign io_coef_out_payload_0_12_32_imag = int_reg_array_12_32_imag;
  assign io_coef_out_payload_0_12_33_real = int_reg_array_12_33_real;
  assign io_coef_out_payload_0_12_33_imag = int_reg_array_12_33_imag;
  assign io_coef_out_payload_0_12_34_real = int_reg_array_12_34_real;
  assign io_coef_out_payload_0_12_34_imag = int_reg_array_12_34_imag;
  assign io_coef_out_payload_0_12_35_real = int_reg_array_12_35_real;
  assign io_coef_out_payload_0_12_35_imag = int_reg_array_12_35_imag;
  assign io_coef_out_payload_0_12_36_real = int_reg_array_12_36_real;
  assign io_coef_out_payload_0_12_36_imag = int_reg_array_12_36_imag;
  assign io_coef_out_payload_0_12_37_real = int_reg_array_12_37_real;
  assign io_coef_out_payload_0_12_37_imag = int_reg_array_12_37_imag;
  assign io_coef_out_payload_0_12_38_real = int_reg_array_12_38_real;
  assign io_coef_out_payload_0_12_38_imag = int_reg_array_12_38_imag;
  assign io_coef_out_payload_0_12_39_real = int_reg_array_12_39_real;
  assign io_coef_out_payload_0_12_39_imag = int_reg_array_12_39_imag;
  assign io_coef_out_payload_0_12_40_real = int_reg_array_12_40_real;
  assign io_coef_out_payload_0_12_40_imag = int_reg_array_12_40_imag;
  assign io_coef_out_payload_0_12_41_real = int_reg_array_12_41_real;
  assign io_coef_out_payload_0_12_41_imag = int_reg_array_12_41_imag;
  assign io_coef_out_payload_0_12_42_real = int_reg_array_12_42_real;
  assign io_coef_out_payload_0_12_42_imag = int_reg_array_12_42_imag;
  assign io_coef_out_payload_0_12_43_real = int_reg_array_12_43_real;
  assign io_coef_out_payload_0_12_43_imag = int_reg_array_12_43_imag;
  assign io_coef_out_payload_0_12_44_real = int_reg_array_12_44_real;
  assign io_coef_out_payload_0_12_44_imag = int_reg_array_12_44_imag;
  assign io_coef_out_payload_0_12_45_real = int_reg_array_12_45_real;
  assign io_coef_out_payload_0_12_45_imag = int_reg_array_12_45_imag;
  assign io_coef_out_payload_0_12_46_real = int_reg_array_12_46_real;
  assign io_coef_out_payload_0_12_46_imag = int_reg_array_12_46_imag;
  assign io_coef_out_payload_0_12_47_real = int_reg_array_12_47_real;
  assign io_coef_out_payload_0_12_47_imag = int_reg_array_12_47_imag;
  assign io_coef_out_payload_0_12_48_real = int_reg_array_12_48_real;
  assign io_coef_out_payload_0_12_48_imag = int_reg_array_12_48_imag;
  assign io_coef_out_payload_0_12_49_real = int_reg_array_12_49_real;
  assign io_coef_out_payload_0_12_49_imag = int_reg_array_12_49_imag;
  assign io_coef_out_payload_0_13_0_real = int_reg_array_13_0_real;
  assign io_coef_out_payload_0_13_0_imag = int_reg_array_13_0_imag;
  assign io_coef_out_payload_0_13_1_real = int_reg_array_13_1_real;
  assign io_coef_out_payload_0_13_1_imag = int_reg_array_13_1_imag;
  assign io_coef_out_payload_0_13_2_real = int_reg_array_13_2_real;
  assign io_coef_out_payload_0_13_2_imag = int_reg_array_13_2_imag;
  assign io_coef_out_payload_0_13_3_real = int_reg_array_13_3_real;
  assign io_coef_out_payload_0_13_3_imag = int_reg_array_13_3_imag;
  assign io_coef_out_payload_0_13_4_real = int_reg_array_13_4_real;
  assign io_coef_out_payload_0_13_4_imag = int_reg_array_13_4_imag;
  assign io_coef_out_payload_0_13_5_real = int_reg_array_13_5_real;
  assign io_coef_out_payload_0_13_5_imag = int_reg_array_13_5_imag;
  assign io_coef_out_payload_0_13_6_real = int_reg_array_13_6_real;
  assign io_coef_out_payload_0_13_6_imag = int_reg_array_13_6_imag;
  assign io_coef_out_payload_0_13_7_real = int_reg_array_13_7_real;
  assign io_coef_out_payload_0_13_7_imag = int_reg_array_13_7_imag;
  assign io_coef_out_payload_0_13_8_real = int_reg_array_13_8_real;
  assign io_coef_out_payload_0_13_8_imag = int_reg_array_13_8_imag;
  assign io_coef_out_payload_0_13_9_real = int_reg_array_13_9_real;
  assign io_coef_out_payload_0_13_9_imag = int_reg_array_13_9_imag;
  assign io_coef_out_payload_0_13_10_real = int_reg_array_13_10_real;
  assign io_coef_out_payload_0_13_10_imag = int_reg_array_13_10_imag;
  assign io_coef_out_payload_0_13_11_real = int_reg_array_13_11_real;
  assign io_coef_out_payload_0_13_11_imag = int_reg_array_13_11_imag;
  assign io_coef_out_payload_0_13_12_real = int_reg_array_13_12_real;
  assign io_coef_out_payload_0_13_12_imag = int_reg_array_13_12_imag;
  assign io_coef_out_payload_0_13_13_real = int_reg_array_13_13_real;
  assign io_coef_out_payload_0_13_13_imag = int_reg_array_13_13_imag;
  assign io_coef_out_payload_0_13_14_real = int_reg_array_13_14_real;
  assign io_coef_out_payload_0_13_14_imag = int_reg_array_13_14_imag;
  assign io_coef_out_payload_0_13_15_real = int_reg_array_13_15_real;
  assign io_coef_out_payload_0_13_15_imag = int_reg_array_13_15_imag;
  assign io_coef_out_payload_0_13_16_real = int_reg_array_13_16_real;
  assign io_coef_out_payload_0_13_16_imag = int_reg_array_13_16_imag;
  assign io_coef_out_payload_0_13_17_real = int_reg_array_13_17_real;
  assign io_coef_out_payload_0_13_17_imag = int_reg_array_13_17_imag;
  assign io_coef_out_payload_0_13_18_real = int_reg_array_13_18_real;
  assign io_coef_out_payload_0_13_18_imag = int_reg_array_13_18_imag;
  assign io_coef_out_payload_0_13_19_real = int_reg_array_13_19_real;
  assign io_coef_out_payload_0_13_19_imag = int_reg_array_13_19_imag;
  assign io_coef_out_payload_0_13_20_real = int_reg_array_13_20_real;
  assign io_coef_out_payload_0_13_20_imag = int_reg_array_13_20_imag;
  assign io_coef_out_payload_0_13_21_real = int_reg_array_13_21_real;
  assign io_coef_out_payload_0_13_21_imag = int_reg_array_13_21_imag;
  assign io_coef_out_payload_0_13_22_real = int_reg_array_13_22_real;
  assign io_coef_out_payload_0_13_22_imag = int_reg_array_13_22_imag;
  assign io_coef_out_payload_0_13_23_real = int_reg_array_13_23_real;
  assign io_coef_out_payload_0_13_23_imag = int_reg_array_13_23_imag;
  assign io_coef_out_payload_0_13_24_real = int_reg_array_13_24_real;
  assign io_coef_out_payload_0_13_24_imag = int_reg_array_13_24_imag;
  assign io_coef_out_payload_0_13_25_real = int_reg_array_13_25_real;
  assign io_coef_out_payload_0_13_25_imag = int_reg_array_13_25_imag;
  assign io_coef_out_payload_0_13_26_real = int_reg_array_13_26_real;
  assign io_coef_out_payload_0_13_26_imag = int_reg_array_13_26_imag;
  assign io_coef_out_payload_0_13_27_real = int_reg_array_13_27_real;
  assign io_coef_out_payload_0_13_27_imag = int_reg_array_13_27_imag;
  assign io_coef_out_payload_0_13_28_real = int_reg_array_13_28_real;
  assign io_coef_out_payload_0_13_28_imag = int_reg_array_13_28_imag;
  assign io_coef_out_payload_0_13_29_real = int_reg_array_13_29_real;
  assign io_coef_out_payload_0_13_29_imag = int_reg_array_13_29_imag;
  assign io_coef_out_payload_0_13_30_real = int_reg_array_13_30_real;
  assign io_coef_out_payload_0_13_30_imag = int_reg_array_13_30_imag;
  assign io_coef_out_payload_0_13_31_real = int_reg_array_13_31_real;
  assign io_coef_out_payload_0_13_31_imag = int_reg_array_13_31_imag;
  assign io_coef_out_payload_0_13_32_real = int_reg_array_13_32_real;
  assign io_coef_out_payload_0_13_32_imag = int_reg_array_13_32_imag;
  assign io_coef_out_payload_0_13_33_real = int_reg_array_13_33_real;
  assign io_coef_out_payload_0_13_33_imag = int_reg_array_13_33_imag;
  assign io_coef_out_payload_0_13_34_real = int_reg_array_13_34_real;
  assign io_coef_out_payload_0_13_34_imag = int_reg_array_13_34_imag;
  assign io_coef_out_payload_0_13_35_real = int_reg_array_13_35_real;
  assign io_coef_out_payload_0_13_35_imag = int_reg_array_13_35_imag;
  assign io_coef_out_payload_0_13_36_real = int_reg_array_13_36_real;
  assign io_coef_out_payload_0_13_36_imag = int_reg_array_13_36_imag;
  assign io_coef_out_payload_0_13_37_real = int_reg_array_13_37_real;
  assign io_coef_out_payload_0_13_37_imag = int_reg_array_13_37_imag;
  assign io_coef_out_payload_0_13_38_real = int_reg_array_13_38_real;
  assign io_coef_out_payload_0_13_38_imag = int_reg_array_13_38_imag;
  assign io_coef_out_payload_0_13_39_real = int_reg_array_13_39_real;
  assign io_coef_out_payload_0_13_39_imag = int_reg_array_13_39_imag;
  assign io_coef_out_payload_0_13_40_real = int_reg_array_13_40_real;
  assign io_coef_out_payload_0_13_40_imag = int_reg_array_13_40_imag;
  assign io_coef_out_payload_0_13_41_real = int_reg_array_13_41_real;
  assign io_coef_out_payload_0_13_41_imag = int_reg_array_13_41_imag;
  assign io_coef_out_payload_0_13_42_real = int_reg_array_13_42_real;
  assign io_coef_out_payload_0_13_42_imag = int_reg_array_13_42_imag;
  assign io_coef_out_payload_0_13_43_real = int_reg_array_13_43_real;
  assign io_coef_out_payload_0_13_43_imag = int_reg_array_13_43_imag;
  assign io_coef_out_payload_0_13_44_real = int_reg_array_13_44_real;
  assign io_coef_out_payload_0_13_44_imag = int_reg_array_13_44_imag;
  assign io_coef_out_payload_0_13_45_real = int_reg_array_13_45_real;
  assign io_coef_out_payload_0_13_45_imag = int_reg_array_13_45_imag;
  assign io_coef_out_payload_0_13_46_real = int_reg_array_13_46_real;
  assign io_coef_out_payload_0_13_46_imag = int_reg_array_13_46_imag;
  assign io_coef_out_payload_0_13_47_real = int_reg_array_13_47_real;
  assign io_coef_out_payload_0_13_47_imag = int_reg_array_13_47_imag;
  assign io_coef_out_payload_0_13_48_real = int_reg_array_13_48_real;
  assign io_coef_out_payload_0_13_48_imag = int_reg_array_13_48_imag;
  assign io_coef_out_payload_0_13_49_real = int_reg_array_13_49_real;
  assign io_coef_out_payload_0_13_49_imag = int_reg_array_13_49_imag;
  assign io_coef_out_payload_0_14_0_real = int_reg_array_14_0_real;
  assign io_coef_out_payload_0_14_0_imag = int_reg_array_14_0_imag;
  assign io_coef_out_payload_0_14_1_real = int_reg_array_14_1_real;
  assign io_coef_out_payload_0_14_1_imag = int_reg_array_14_1_imag;
  assign io_coef_out_payload_0_14_2_real = int_reg_array_14_2_real;
  assign io_coef_out_payload_0_14_2_imag = int_reg_array_14_2_imag;
  assign io_coef_out_payload_0_14_3_real = int_reg_array_14_3_real;
  assign io_coef_out_payload_0_14_3_imag = int_reg_array_14_3_imag;
  assign io_coef_out_payload_0_14_4_real = int_reg_array_14_4_real;
  assign io_coef_out_payload_0_14_4_imag = int_reg_array_14_4_imag;
  assign io_coef_out_payload_0_14_5_real = int_reg_array_14_5_real;
  assign io_coef_out_payload_0_14_5_imag = int_reg_array_14_5_imag;
  assign io_coef_out_payload_0_14_6_real = int_reg_array_14_6_real;
  assign io_coef_out_payload_0_14_6_imag = int_reg_array_14_6_imag;
  assign io_coef_out_payload_0_14_7_real = int_reg_array_14_7_real;
  assign io_coef_out_payload_0_14_7_imag = int_reg_array_14_7_imag;
  assign io_coef_out_payload_0_14_8_real = int_reg_array_14_8_real;
  assign io_coef_out_payload_0_14_8_imag = int_reg_array_14_8_imag;
  assign io_coef_out_payload_0_14_9_real = int_reg_array_14_9_real;
  assign io_coef_out_payload_0_14_9_imag = int_reg_array_14_9_imag;
  assign io_coef_out_payload_0_14_10_real = int_reg_array_14_10_real;
  assign io_coef_out_payload_0_14_10_imag = int_reg_array_14_10_imag;
  assign io_coef_out_payload_0_14_11_real = int_reg_array_14_11_real;
  assign io_coef_out_payload_0_14_11_imag = int_reg_array_14_11_imag;
  assign io_coef_out_payload_0_14_12_real = int_reg_array_14_12_real;
  assign io_coef_out_payload_0_14_12_imag = int_reg_array_14_12_imag;
  assign io_coef_out_payload_0_14_13_real = int_reg_array_14_13_real;
  assign io_coef_out_payload_0_14_13_imag = int_reg_array_14_13_imag;
  assign io_coef_out_payload_0_14_14_real = int_reg_array_14_14_real;
  assign io_coef_out_payload_0_14_14_imag = int_reg_array_14_14_imag;
  assign io_coef_out_payload_0_14_15_real = int_reg_array_14_15_real;
  assign io_coef_out_payload_0_14_15_imag = int_reg_array_14_15_imag;
  assign io_coef_out_payload_0_14_16_real = int_reg_array_14_16_real;
  assign io_coef_out_payload_0_14_16_imag = int_reg_array_14_16_imag;
  assign io_coef_out_payload_0_14_17_real = int_reg_array_14_17_real;
  assign io_coef_out_payload_0_14_17_imag = int_reg_array_14_17_imag;
  assign io_coef_out_payload_0_14_18_real = int_reg_array_14_18_real;
  assign io_coef_out_payload_0_14_18_imag = int_reg_array_14_18_imag;
  assign io_coef_out_payload_0_14_19_real = int_reg_array_14_19_real;
  assign io_coef_out_payload_0_14_19_imag = int_reg_array_14_19_imag;
  assign io_coef_out_payload_0_14_20_real = int_reg_array_14_20_real;
  assign io_coef_out_payload_0_14_20_imag = int_reg_array_14_20_imag;
  assign io_coef_out_payload_0_14_21_real = int_reg_array_14_21_real;
  assign io_coef_out_payload_0_14_21_imag = int_reg_array_14_21_imag;
  assign io_coef_out_payload_0_14_22_real = int_reg_array_14_22_real;
  assign io_coef_out_payload_0_14_22_imag = int_reg_array_14_22_imag;
  assign io_coef_out_payload_0_14_23_real = int_reg_array_14_23_real;
  assign io_coef_out_payload_0_14_23_imag = int_reg_array_14_23_imag;
  assign io_coef_out_payload_0_14_24_real = int_reg_array_14_24_real;
  assign io_coef_out_payload_0_14_24_imag = int_reg_array_14_24_imag;
  assign io_coef_out_payload_0_14_25_real = int_reg_array_14_25_real;
  assign io_coef_out_payload_0_14_25_imag = int_reg_array_14_25_imag;
  assign io_coef_out_payload_0_14_26_real = int_reg_array_14_26_real;
  assign io_coef_out_payload_0_14_26_imag = int_reg_array_14_26_imag;
  assign io_coef_out_payload_0_14_27_real = int_reg_array_14_27_real;
  assign io_coef_out_payload_0_14_27_imag = int_reg_array_14_27_imag;
  assign io_coef_out_payload_0_14_28_real = int_reg_array_14_28_real;
  assign io_coef_out_payload_0_14_28_imag = int_reg_array_14_28_imag;
  assign io_coef_out_payload_0_14_29_real = int_reg_array_14_29_real;
  assign io_coef_out_payload_0_14_29_imag = int_reg_array_14_29_imag;
  assign io_coef_out_payload_0_14_30_real = int_reg_array_14_30_real;
  assign io_coef_out_payload_0_14_30_imag = int_reg_array_14_30_imag;
  assign io_coef_out_payload_0_14_31_real = int_reg_array_14_31_real;
  assign io_coef_out_payload_0_14_31_imag = int_reg_array_14_31_imag;
  assign io_coef_out_payload_0_14_32_real = int_reg_array_14_32_real;
  assign io_coef_out_payload_0_14_32_imag = int_reg_array_14_32_imag;
  assign io_coef_out_payload_0_14_33_real = int_reg_array_14_33_real;
  assign io_coef_out_payload_0_14_33_imag = int_reg_array_14_33_imag;
  assign io_coef_out_payload_0_14_34_real = int_reg_array_14_34_real;
  assign io_coef_out_payload_0_14_34_imag = int_reg_array_14_34_imag;
  assign io_coef_out_payload_0_14_35_real = int_reg_array_14_35_real;
  assign io_coef_out_payload_0_14_35_imag = int_reg_array_14_35_imag;
  assign io_coef_out_payload_0_14_36_real = int_reg_array_14_36_real;
  assign io_coef_out_payload_0_14_36_imag = int_reg_array_14_36_imag;
  assign io_coef_out_payload_0_14_37_real = int_reg_array_14_37_real;
  assign io_coef_out_payload_0_14_37_imag = int_reg_array_14_37_imag;
  assign io_coef_out_payload_0_14_38_real = int_reg_array_14_38_real;
  assign io_coef_out_payload_0_14_38_imag = int_reg_array_14_38_imag;
  assign io_coef_out_payload_0_14_39_real = int_reg_array_14_39_real;
  assign io_coef_out_payload_0_14_39_imag = int_reg_array_14_39_imag;
  assign io_coef_out_payload_0_14_40_real = int_reg_array_14_40_real;
  assign io_coef_out_payload_0_14_40_imag = int_reg_array_14_40_imag;
  assign io_coef_out_payload_0_14_41_real = int_reg_array_14_41_real;
  assign io_coef_out_payload_0_14_41_imag = int_reg_array_14_41_imag;
  assign io_coef_out_payload_0_14_42_real = int_reg_array_14_42_real;
  assign io_coef_out_payload_0_14_42_imag = int_reg_array_14_42_imag;
  assign io_coef_out_payload_0_14_43_real = int_reg_array_14_43_real;
  assign io_coef_out_payload_0_14_43_imag = int_reg_array_14_43_imag;
  assign io_coef_out_payload_0_14_44_real = int_reg_array_14_44_real;
  assign io_coef_out_payload_0_14_44_imag = int_reg_array_14_44_imag;
  assign io_coef_out_payload_0_14_45_real = int_reg_array_14_45_real;
  assign io_coef_out_payload_0_14_45_imag = int_reg_array_14_45_imag;
  assign io_coef_out_payload_0_14_46_real = int_reg_array_14_46_real;
  assign io_coef_out_payload_0_14_46_imag = int_reg_array_14_46_imag;
  assign io_coef_out_payload_0_14_47_real = int_reg_array_14_47_real;
  assign io_coef_out_payload_0_14_47_imag = int_reg_array_14_47_imag;
  assign io_coef_out_payload_0_14_48_real = int_reg_array_14_48_real;
  assign io_coef_out_payload_0_14_48_imag = int_reg_array_14_48_imag;
  assign io_coef_out_payload_0_14_49_real = int_reg_array_14_49_real;
  assign io_coef_out_payload_0_14_49_imag = int_reg_array_14_49_imag;
  assign io_coef_out_payload_0_15_0_real = int_reg_array_15_0_real;
  assign io_coef_out_payload_0_15_0_imag = int_reg_array_15_0_imag;
  assign io_coef_out_payload_0_15_1_real = int_reg_array_15_1_real;
  assign io_coef_out_payload_0_15_1_imag = int_reg_array_15_1_imag;
  assign io_coef_out_payload_0_15_2_real = int_reg_array_15_2_real;
  assign io_coef_out_payload_0_15_2_imag = int_reg_array_15_2_imag;
  assign io_coef_out_payload_0_15_3_real = int_reg_array_15_3_real;
  assign io_coef_out_payload_0_15_3_imag = int_reg_array_15_3_imag;
  assign io_coef_out_payload_0_15_4_real = int_reg_array_15_4_real;
  assign io_coef_out_payload_0_15_4_imag = int_reg_array_15_4_imag;
  assign io_coef_out_payload_0_15_5_real = int_reg_array_15_5_real;
  assign io_coef_out_payload_0_15_5_imag = int_reg_array_15_5_imag;
  assign io_coef_out_payload_0_15_6_real = int_reg_array_15_6_real;
  assign io_coef_out_payload_0_15_6_imag = int_reg_array_15_6_imag;
  assign io_coef_out_payload_0_15_7_real = int_reg_array_15_7_real;
  assign io_coef_out_payload_0_15_7_imag = int_reg_array_15_7_imag;
  assign io_coef_out_payload_0_15_8_real = int_reg_array_15_8_real;
  assign io_coef_out_payload_0_15_8_imag = int_reg_array_15_8_imag;
  assign io_coef_out_payload_0_15_9_real = int_reg_array_15_9_real;
  assign io_coef_out_payload_0_15_9_imag = int_reg_array_15_9_imag;
  assign io_coef_out_payload_0_15_10_real = int_reg_array_15_10_real;
  assign io_coef_out_payload_0_15_10_imag = int_reg_array_15_10_imag;
  assign io_coef_out_payload_0_15_11_real = int_reg_array_15_11_real;
  assign io_coef_out_payload_0_15_11_imag = int_reg_array_15_11_imag;
  assign io_coef_out_payload_0_15_12_real = int_reg_array_15_12_real;
  assign io_coef_out_payload_0_15_12_imag = int_reg_array_15_12_imag;
  assign io_coef_out_payload_0_15_13_real = int_reg_array_15_13_real;
  assign io_coef_out_payload_0_15_13_imag = int_reg_array_15_13_imag;
  assign io_coef_out_payload_0_15_14_real = int_reg_array_15_14_real;
  assign io_coef_out_payload_0_15_14_imag = int_reg_array_15_14_imag;
  assign io_coef_out_payload_0_15_15_real = int_reg_array_15_15_real;
  assign io_coef_out_payload_0_15_15_imag = int_reg_array_15_15_imag;
  assign io_coef_out_payload_0_15_16_real = int_reg_array_15_16_real;
  assign io_coef_out_payload_0_15_16_imag = int_reg_array_15_16_imag;
  assign io_coef_out_payload_0_15_17_real = int_reg_array_15_17_real;
  assign io_coef_out_payload_0_15_17_imag = int_reg_array_15_17_imag;
  assign io_coef_out_payload_0_15_18_real = int_reg_array_15_18_real;
  assign io_coef_out_payload_0_15_18_imag = int_reg_array_15_18_imag;
  assign io_coef_out_payload_0_15_19_real = int_reg_array_15_19_real;
  assign io_coef_out_payload_0_15_19_imag = int_reg_array_15_19_imag;
  assign io_coef_out_payload_0_15_20_real = int_reg_array_15_20_real;
  assign io_coef_out_payload_0_15_20_imag = int_reg_array_15_20_imag;
  assign io_coef_out_payload_0_15_21_real = int_reg_array_15_21_real;
  assign io_coef_out_payload_0_15_21_imag = int_reg_array_15_21_imag;
  assign io_coef_out_payload_0_15_22_real = int_reg_array_15_22_real;
  assign io_coef_out_payload_0_15_22_imag = int_reg_array_15_22_imag;
  assign io_coef_out_payload_0_15_23_real = int_reg_array_15_23_real;
  assign io_coef_out_payload_0_15_23_imag = int_reg_array_15_23_imag;
  assign io_coef_out_payload_0_15_24_real = int_reg_array_15_24_real;
  assign io_coef_out_payload_0_15_24_imag = int_reg_array_15_24_imag;
  assign io_coef_out_payload_0_15_25_real = int_reg_array_15_25_real;
  assign io_coef_out_payload_0_15_25_imag = int_reg_array_15_25_imag;
  assign io_coef_out_payload_0_15_26_real = int_reg_array_15_26_real;
  assign io_coef_out_payload_0_15_26_imag = int_reg_array_15_26_imag;
  assign io_coef_out_payload_0_15_27_real = int_reg_array_15_27_real;
  assign io_coef_out_payload_0_15_27_imag = int_reg_array_15_27_imag;
  assign io_coef_out_payload_0_15_28_real = int_reg_array_15_28_real;
  assign io_coef_out_payload_0_15_28_imag = int_reg_array_15_28_imag;
  assign io_coef_out_payload_0_15_29_real = int_reg_array_15_29_real;
  assign io_coef_out_payload_0_15_29_imag = int_reg_array_15_29_imag;
  assign io_coef_out_payload_0_15_30_real = int_reg_array_15_30_real;
  assign io_coef_out_payload_0_15_30_imag = int_reg_array_15_30_imag;
  assign io_coef_out_payload_0_15_31_real = int_reg_array_15_31_real;
  assign io_coef_out_payload_0_15_31_imag = int_reg_array_15_31_imag;
  assign io_coef_out_payload_0_15_32_real = int_reg_array_15_32_real;
  assign io_coef_out_payload_0_15_32_imag = int_reg_array_15_32_imag;
  assign io_coef_out_payload_0_15_33_real = int_reg_array_15_33_real;
  assign io_coef_out_payload_0_15_33_imag = int_reg_array_15_33_imag;
  assign io_coef_out_payload_0_15_34_real = int_reg_array_15_34_real;
  assign io_coef_out_payload_0_15_34_imag = int_reg_array_15_34_imag;
  assign io_coef_out_payload_0_15_35_real = int_reg_array_15_35_real;
  assign io_coef_out_payload_0_15_35_imag = int_reg_array_15_35_imag;
  assign io_coef_out_payload_0_15_36_real = int_reg_array_15_36_real;
  assign io_coef_out_payload_0_15_36_imag = int_reg_array_15_36_imag;
  assign io_coef_out_payload_0_15_37_real = int_reg_array_15_37_real;
  assign io_coef_out_payload_0_15_37_imag = int_reg_array_15_37_imag;
  assign io_coef_out_payload_0_15_38_real = int_reg_array_15_38_real;
  assign io_coef_out_payload_0_15_38_imag = int_reg_array_15_38_imag;
  assign io_coef_out_payload_0_15_39_real = int_reg_array_15_39_real;
  assign io_coef_out_payload_0_15_39_imag = int_reg_array_15_39_imag;
  assign io_coef_out_payload_0_15_40_real = int_reg_array_15_40_real;
  assign io_coef_out_payload_0_15_40_imag = int_reg_array_15_40_imag;
  assign io_coef_out_payload_0_15_41_real = int_reg_array_15_41_real;
  assign io_coef_out_payload_0_15_41_imag = int_reg_array_15_41_imag;
  assign io_coef_out_payload_0_15_42_real = int_reg_array_15_42_real;
  assign io_coef_out_payload_0_15_42_imag = int_reg_array_15_42_imag;
  assign io_coef_out_payload_0_15_43_real = int_reg_array_15_43_real;
  assign io_coef_out_payload_0_15_43_imag = int_reg_array_15_43_imag;
  assign io_coef_out_payload_0_15_44_real = int_reg_array_15_44_real;
  assign io_coef_out_payload_0_15_44_imag = int_reg_array_15_44_imag;
  assign io_coef_out_payload_0_15_45_real = int_reg_array_15_45_real;
  assign io_coef_out_payload_0_15_45_imag = int_reg_array_15_45_imag;
  assign io_coef_out_payload_0_15_46_real = int_reg_array_15_46_real;
  assign io_coef_out_payload_0_15_46_imag = int_reg_array_15_46_imag;
  assign io_coef_out_payload_0_15_47_real = int_reg_array_15_47_real;
  assign io_coef_out_payload_0_15_47_imag = int_reg_array_15_47_imag;
  assign io_coef_out_payload_0_15_48_real = int_reg_array_15_48_real;
  assign io_coef_out_payload_0_15_48_imag = int_reg_array_15_48_imag;
  assign io_coef_out_payload_0_15_49_real = int_reg_array_15_49_real;
  assign io_coef_out_payload_0_15_49_imag = int_reg_array_15_49_imag;
  assign io_coef_out_payload_0_16_0_real = int_reg_array_16_0_real;
  assign io_coef_out_payload_0_16_0_imag = int_reg_array_16_0_imag;
  assign io_coef_out_payload_0_16_1_real = int_reg_array_16_1_real;
  assign io_coef_out_payload_0_16_1_imag = int_reg_array_16_1_imag;
  assign io_coef_out_payload_0_16_2_real = int_reg_array_16_2_real;
  assign io_coef_out_payload_0_16_2_imag = int_reg_array_16_2_imag;
  assign io_coef_out_payload_0_16_3_real = int_reg_array_16_3_real;
  assign io_coef_out_payload_0_16_3_imag = int_reg_array_16_3_imag;
  assign io_coef_out_payload_0_16_4_real = int_reg_array_16_4_real;
  assign io_coef_out_payload_0_16_4_imag = int_reg_array_16_4_imag;
  assign io_coef_out_payload_0_16_5_real = int_reg_array_16_5_real;
  assign io_coef_out_payload_0_16_5_imag = int_reg_array_16_5_imag;
  assign io_coef_out_payload_0_16_6_real = int_reg_array_16_6_real;
  assign io_coef_out_payload_0_16_6_imag = int_reg_array_16_6_imag;
  assign io_coef_out_payload_0_16_7_real = int_reg_array_16_7_real;
  assign io_coef_out_payload_0_16_7_imag = int_reg_array_16_7_imag;
  assign io_coef_out_payload_0_16_8_real = int_reg_array_16_8_real;
  assign io_coef_out_payload_0_16_8_imag = int_reg_array_16_8_imag;
  assign io_coef_out_payload_0_16_9_real = int_reg_array_16_9_real;
  assign io_coef_out_payload_0_16_9_imag = int_reg_array_16_9_imag;
  assign io_coef_out_payload_0_16_10_real = int_reg_array_16_10_real;
  assign io_coef_out_payload_0_16_10_imag = int_reg_array_16_10_imag;
  assign io_coef_out_payload_0_16_11_real = int_reg_array_16_11_real;
  assign io_coef_out_payload_0_16_11_imag = int_reg_array_16_11_imag;
  assign io_coef_out_payload_0_16_12_real = int_reg_array_16_12_real;
  assign io_coef_out_payload_0_16_12_imag = int_reg_array_16_12_imag;
  assign io_coef_out_payload_0_16_13_real = int_reg_array_16_13_real;
  assign io_coef_out_payload_0_16_13_imag = int_reg_array_16_13_imag;
  assign io_coef_out_payload_0_16_14_real = int_reg_array_16_14_real;
  assign io_coef_out_payload_0_16_14_imag = int_reg_array_16_14_imag;
  assign io_coef_out_payload_0_16_15_real = int_reg_array_16_15_real;
  assign io_coef_out_payload_0_16_15_imag = int_reg_array_16_15_imag;
  assign io_coef_out_payload_0_16_16_real = int_reg_array_16_16_real;
  assign io_coef_out_payload_0_16_16_imag = int_reg_array_16_16_imag;
  assign io_coef_out_payload_0_16_17_real = int_reg_array_16_17_real;
  assign io_coef_out_payload_0_16_17_imag = int_reg_array_16_17_imag;
  assign io_coef_out_payload_0_16_18_real = int_reg_array_16_18_real;
  assign io_coef_out_payload_0_16_18_imag = int_reg_array_16_18_imag;
  assign io_coef_out_payload_0_16_19_real = int_reg_array_16_19_real;
  assign io_coef_out_payload_0_16_19_imag = int_reg_array_16_19_imag;
  assign io_coef_out_payload_0_16_20_real = int_reg_array_16_20_real;
  assign io_coef_out_payload_0_16_20_imag = int_reg_array_16_20_imag;
  assign io_coef_out_payload_0_16_21_real = int_reg_array_16_21_real;
  assign io_coef_out_payload_0_16_21_imag = int_reg_array_16_21_imag;
  assign io_coef_out_payload_0_16_22_real = int_reg_array_16_22_real;
  assign io_coef_out_payload_0_16_22_imag = int_reg_array_16_22_imag;
  assign io_coef_out_payload_0_16_23_real = int_reg_array_16_23_real;
  assign io_coef_out_payload_0_16_23_imag = int_reg_array_16_23_imag;
  assign io_coef_out_payload_0_16_24_real = int_reg_array_16_24_real;
  assign io_coef_out_payload_0_16_24_imag = int_reg_array_16_24_imag;
  assign io_coef_out_payload_0_16_25_real = int_reg_array_16_25_real;
  assign io_coef_out_payload_0_16_25_imag = int_reg_array_16_25_imag;
  assign io_coef_out_payload_0_16_26_real = int_reg_array_16_26_real;
  assign io_coef_out_payload_0_16_26_imag = int_reg_array_16_26_imag;
  assign io_coef_out_payload_0_16_27_real = int_reg_array_16_27_real;
  assign io_coef_out_payload_0_16_27_imag = int_reg_array_16_27_imag;
  assign io_coef_out_payload_0_16_28_real = int_reg_array_16_28_real;
  assign io_coef_out_payload_0_16_28_imag = int_reg_array_16_28_imag;
  assign io_coef_out_payload_0_16_29_real = int_reg_array_16_29_real;
  assign io_coef_out_payload_0_16_29_imag = int_reg_array_16_29_imag;
  assign io_coef_out_payload_0_16_30_real = int_reg_array_16_30_real;
  assign io_coef_out_payload_0_16_30_imag = int_reg_array_16_30_imag;
  assign io_coef_out_payload_0_16_31_real = int_reg_array_16_31_real;
  assign io_coef_out_payload_0_16_31_imag = int_reg_array_16_31_imag;
  assign io_coef_out_payload_0_16_32_real = int_reg_array_16_32_real;
  assign io_coef_out_payload_0_16_32_imag = int_reg_array_16_32_imag;
  assign io_coef_out_payload_0_16_33_real = int_reg_array_16_33_real;
  assign io_coef_out_payload_0_16_33_imag = int_reg_array_16_33_imag;
  assign io_coef_out_payload_0_16_34_real = int_reg_array_16_34_real;
  assign io_coef_out_payload_0_16_34_imag = int_reg_array_16_34_imag;
  assign io_coef_out_payload_0_16_35_real = int_reg_array_16_35_real;
  assign io_coef_out_payload_0_16_35_imag = int_reg_array_16_35_imag;
  assign io_coef_out_payload_0_16_36_real = int_reg_array_16_36_real;
  assign io_coef_out_payload_0_16_36_imag = int_reg_array_16_36_imag;
  assign io_coef_out_payload_0_16_37_real = int_reg_array_16_37_real;
  assign io_coef_out_payload_0_16_37_imag = int_reg_array_16_37_imag;
  assign io_coef_out_payload_0_16_38_real = int_reg_array_16_38_real;
  assign io_coef_out_payload_0_16_38_imag = int_reg_array_16_38_imag;
  assign io_coef_out_payload_0_16_39_real = int_reg_array_16_39_real;
  assign io_coef_out_payload_0_16_39_imag = int_reg_array_16_39_imag;
  assign io_coef_out_payload_0_16_40_real = int_reg_array_16_40_real;
  assign io_coef_out_payload_0_16_40_imag = int_reg_array_16_40_imag;
  assign io_coef_out_payload_0_16_41_real = int_reg_array_16_41_real;
  assign io_coef_out_payload_0_16_41_imag = int_reg_array_16_41_imag;
  assign io_coef_out_payload_0_16_42_real = int_reg_array_16_42_real;
  assign io_coef_out_payload_0_16_42_imag = int_reg_array_16_42_imag;
  assign io_coef_out_payload_0_16_43_real = int_reg_array_16_43_real;
  assign io_coef_out_payload_0_16_43_imag = int_reg_array_16_43_imag;
  assign io_coef_out_payload_0_16_44_real = int_reg_array_16_44_real;
  assign io_coef_out_payload_0_16_44_imag = int_reg_array_16_44_imag;
  assign io_coef_out_payload_0_16_45_real = int_reg_array_16_45_real;
  assign io_coef_out_payload_0_16_45_imag = int_reg_array_16_45_imag;
  assign io_coef_out_payload_0_16_46_real = int_reg_array_16_46_real;
  assign io_coef_out_payload_0_16_46_imag = int_reg_array_16_46_imag;
  assign io_coef_out_payload_0_16_47_real = int_reg_array_16_47_real;
  assign io_coef_out_payload_0_16_47_imag = int_reg_array_16_47_imag;
  assign io_coef_out_payload_0_16_48_real = int_reg_array_16_48_real;
  assign io_coef_out_payload_0_16_48_imag = int_reg_array_16_48_imag;
  assign io_coef_out_payload_0_16_49_real = int_reg_array_16_49_real;
  assign io_coef_out_payload_0_16_49_imag = int_reg_array_16_49_imag;
  assign io_coef_out_payload_0_17_0_real = int_reg_array_17_0_real;
  assign io_coef_out_payload_0_17_0_imag = int_reg_array_17_0_imag;
  assign io_coef_out_payload_0_17_1_real = int_reg_array_17_1_real;
  assign io_coef_out_payload_0_17_1_imag = int_reg_array_17_1_imag;
  assign io_coef_out_payload_0_17_2_real = int_reg_array_17_2_real;
  assign io_coef_out_payload_0_17_2_imag = int_reg_array_17_2_imag;
  assign io_coef_out_payload_0_17_3_real = int_reg_array_17_3_real;
  assign io_coef_out_payload_0_17_3_imag = int_reg_array_17_3_imag;
  assign io_coef_out_payload_0_17_4_real = int_reg_array_17_4_real;
  assign io_coef_out_payload_0_17_4_imag = int_reg_array_17_4_imag;
  assign io_coef_out_payload_0_17_5_real = int_reg_array_17_5_real;
  assign io_coef_out_payload_0_17_5_imag = int_reg_array_17_5_imag;
  assign io_coef_out_payload_0_17_6_real = int_reg_array_17_6_real;
  assign io_coef_out_payload_0_17_6_imag = int_reg_array_17_6_imag;
  assign io_coef_out_payload_0_17_7_real = int_reg_array_17_7_real;
  assign io_coef_out_payload_0_17_7_imag = int_reg_array_17_7_imag;
  assign io_coef_out_payload_0_17_8_real = int_reg_array_17_8_real;
  assign io_coef_out_payload_0_17_8_imag = int_reg_array_17_8_imag;
  assign io_coef_out_payload_0_17_9_real = int_reg_array_17_9_real;
  assign io_coef_out_payload_0_17_9_imag = int_reg_array_17_9_imag;
  assign io_coef_out_payload_0_17_10_real = int_reg_array_17_10_real;
  assign io_coef_out_payload_0_17_10_imag = int_reg_array_17_10_imag;
  assign io_coef_out_payload_0_17_11_real = int_reg_array_17_11_real;
  assign io_coef_out_payload_0_17_11_imag = int_reg_array_17_11_imag;
  assign io_coef_out_payload_0_17_12_real = int_reg_array_17_12_real;
  assign io_coef_out_payload_0_17_12_imag = int_reg_array_17_12_imag;
  assign io_coef_out_payload_0_17_13_real = int_reg_array_17_13_real;
  assign io_coef_out_payload_0_17_13_imag = int_reg_array_17_13_imag;
  assign io_coef_out_payload_0_17_14_real = int_reg_array_17_14_real;
  assign io_coef_out_payload_0_17_14_imag = int_reg_array_17_14_imag;
  assign io_coef_out_payload_0_17_15_real = int_reg_array_17_15_real;
  assign io_coef_out_payload_0_17_15_imag = int_reg_array_17_15_imag;
  assign io_coef_out_payload_0_17_16_real = int_reg_array_17_16_real;
  assign io_coef_out_payload_0_17_16_imag = int_reg_array_17_16_imag;
  assign io_coef_out_payload_0_17_17_real = int_reg_array_17_17_real;
  assign io_coef_out_payload_0_17_17_imag = int_reg_array_17_17_imag;
  assign io_coef_out_payload_0_17_18_real = int_reg_array_17_18_real;
  assign io_coef_out_payload_0_17_18_imag = int_reg_array_17_18_imag;
  assign io_coef_out_payload_0_17_19_real = int_reg_array_17_19_real;
  assign io_coef_out_payload_0_17_19_imag = int_reg_array_17_19_imag;
  assign io_coef_out_payload_0_17_20_real = int_reg_array_17_20_real;
  assign io_coef_out_payload_0_17_20_imag = int_reg_array_17_20_imag;
  assign io_coef_out_payload_0_17_21_real = int_reg_array_17_21_real;
  assign io_coef_out_payload_0_17_21_imag = int_reg_array_17_21_imag;
  assign io_coef_out_payload_0_17_22_real = int_reg_array_17_22_real;
  assign io_coef_out_payload_0_17_22_imag = int_reg_array_17_22_imag;
  assign io_coef_out_payload_0_17_23_real = int_reg_array_17_23_real;
  assign io_coef_out_payload_0_17_23_imag = int_reg_array_17_23_imag;
  assign io_coef_out_payload_0_17_24_real = int_reg_array_17_24_real;
  assign io_coef_out_payload_0_17_24_imag = int_reg_array_17_24_imag;
  assign io_coef_out_payload_0_17_25_real = int_reg_array_17_25_real;
  assign io_coef_out_payload_0_17_25_imag = int_reg_array_17_25_imag;
  assign io_coef_out_payload_0_17_26_real = int_reg_array_17_26_real;
  assign io_coef_out_payload_0_17_26_imag = int_reg_array_17_26_imag;
  assign io_coef_out_payload_0_17_27_real = int_reg_array_17_27_real;
  assign io_coef_out_payload_0_17_27_imag = int_reg_array_17_27_imag;
  assign io_coef_out_payload_0_17_28_real = int_reg_array_17_28_real;
  assign io_coef_out_payload_0_17_28_imag = int_reg_array_17_28_imag;
  assign io_coef_out_payload_0_17_29_real = int_reg_array_17_29_real;
  assign io_coef_out_payload_0_17_29_imag = int_reg_array_17_29_imag;
  assign io_coef_out_payload_0_17_30_real = int_reg_array_17_30_real;
  assign io_coef_out_payload_0_17_30_imag = int_reg_array_17_30_imag;
  assign io_coef_out_payload_0_17_31_real = int_reg_array_17_31_real;
  assign io_coef_out_payload_0_17_31_imag = int_reg_array_17_31_imag;
  assign io_coef_out_payload_0_17_32_real = int_reg_array_17_32_real;
  assign io_coef_out_payload_0_17_32_imag = int_reg_array_17_32_imag;
  assign io_coef_out_payload_0_17_33_real = int_reg_array_17_33_real;
  assign io_coef_out_payload_0_17_33_imag = int_reg_array_17_33_imag;
  assign io_coef_out_payload_0_17_34_real = int_reg_array_17_34_real;
  assign io_coef_out_payload_0_17_34_imag = int_reg_array_17_34_imag;
  assign io_coef_out_payload_0_17_35_real = int_reg_array_17_35_real;
  assign io_coef_out_payload_0_17_35_imag = int_reg_array_17_35_imag;
  assign io_coef_out_payload_0_17_36_real = int_reg_array_17_36_real;
  assign io_coef_out_payload_0_17_36_imag = int_reg_array_17_36_imag;
  assign io_coef_out_payload_0_17_37_real = int_reg_array_17_37_real;
  assign io_coef_out_payload_0_17_37_imag = int_reg_array_17_37_imag;
  assign io_coef_out_payload_0_17_38_real = int_reg_array_17_38_real;
  assign io_coef_out_payload_0_17_38_imag = int_reg_array_17_38_imag;
  assign io_coef_out_payload_0_17_39_real = int_reg_array_17_39_real;
  assign io_coef_out_payload_0_17_39_imag = int_reg_array_17_39_imag;
  assign io_coef_out_payload_0_17_40_real = int_reg_array_17_40_real;
  assign io_coef_out_payload_0_17_40_imag = int_reg_array_17_40_imag;
  assign io_coef_out_payload_0_17_41_real = int_reg_array_17_41_real;
  assign io_coef_out_payload_0_17_41_imag = int_reg_array_17_41_imag;
  assign io_coef_out_payload_0_17_42_real = int_reg_array_17_42_real;
  assign io_coef_out_payload_0_17_42_imag = int_reg_array_17_42_imag;
  assign io_coef_out_payload_0_17_43_real = int_reg_array_17_43_real;
  assign io_coef_out_payload_0_17_43_imag = int_reg_array_17_43_imag;
  assign io_coef_out_payload_0_17_44_real = int_reg_array_17_44_real;
  assign io_coef_out_payload_0_17_44_imag = int_reg_array_17_44_imag;
  assign io_coef_out_payload_0_17_45_real = int_reg_array_17_45_real;
  assign io_coef_out_payload_0_17_45_imag = int_reg_array_17_45_imag;
  assign io_coef_out_payload_0_17_46_real = int_reg_array_17_46_real;
  assign io_coef_out_payload_0_17_46_imag = int_reg_array_17_46_imag;
  assign io_coef_out_payload_0_17_47_real = int_reg_array_17_47_real;
  assign io_coef_out_payload_0_17_47_imag = int_reg_array_17_47_imag;
  assign io_coef_out_payload_0_17_48_real = int_reg_array_17_48_real;
  assign io_coef_out_payload_0_17_48_imag = int_reg_array_17_48_imag;
  assign io_coef_out_payload_0_17_49_real = int_reg_array_17_49_real;
  assign io_coef_out_payload_0_17_49_imag = int_reg_array_17_49_imag;
  assign io_coef_out_payload_0_18_0_real = int_reg_array_18_0_real;
  assign io_coef_out_payload_0_18_0_imag = int_reg_array_18_0_imag;
  assign io_coef_out_payload_0_18_1_real = int_reg_array_18_1_real;
  assign io_coef_out_payload_0_18_1_imag = int_reg_array_18_1_imag;
  assign io_coef_out_payload_0_18_2_real = int_reg_array_18_2_real;
  assign io_coef_out_payload_0_18_2_imag = int_reg_array_18_2_imag;
  assign io_coef_out_payload_0_18_3_real = int_reg_array_18_3_real;
  assign io_coef_out_payload_0_18_3_imag = int_reg_array_18_3_imag;
  assign io_coef_out_payload_0_18_4_real = int_reg_array_18_4_real;
  assign io_coef_out_payload_0_18_4_imag = int_reg_array_18_4_imag;
  assign io_coef_out_payload_0_18_5_real = int_reg_array_18_5_real;
  assign io_coef_out_payload_0_18_5_imag = int_reg_array_18_5_imag;
  assign io_coef_out_payload_0_18_6_real = int_reg_array_18_6_real;
  assign io_coef_out_payload_0_18_6_imag = int_reg_array_18_6_imag;
  assign io_coef_out_payload_0_18_7_real = int_reg_array_18_7_real;
  assign io_coef_out_payload_0_18_7_imag = int_reg_array_18_7_imag;
  assign io_coef_out_payload_0_18_8_real = int_reg_array_18_8_real;
  assign io_coef_out_payload_0_18_8_imag = int_reg_array_18_8_imag;
  assign io_coef_out_payload_0_18_9_real = int_reg_array_18_9_real;
  assign io_coef_out_payload_0_18_9_imag = int_reg_array_18_9_imag;
  assign io_coef_out_payload_0_18_10_real = int_reg_array_18_10_real;
  assign io_coef_out_payload_0_18_10_imag = int_reg_array_18_10_imag;
  assign io_coef_out_payload_0_18_11_real = int_reg_array_18_11_real;
  assign io_coef_out_payload_0_18_11_imag = int_reg_array_18_11_imag;
  assign io_coef_out_payload_0_18_12_real = int_reg_array_18_12_real;
  assign io_coef_out_payload_0_18_12_imag = int_reg_array_18_12_imag;
  assign io_coef_out_payload_0_18_13_real = int_reg_array_18_13_real;
  assign io_coef_out_payload_0_18_13_imag = int_reg_array_18_13_imag;
  assign io_coef_out_payload_0_18_14_real = int_reg_array_18_14_real;
  assign io_coef_out_payload_0_18_14_imag = int_reg_array_18_14_imag;
  assign io_coef_out_payload_0_18_15_real = int_reg_array_18_15_real;
  assign io_coef_out_payload_0_18_15_imag = int_reg_array_18_15_imag;
  assign io_coef_out_payload_0_18_16_real = int_reg_array_18_16_real;
  assign io_coef_out_payload_0_18_16_imag = int_reg_array_18_16_imag;
  assign io_coef_out_payload_0_18_17_real = int_reg_array_18_17_real;
  assign io_coef_out_payload_0_18_17_imag = int_reg_array_18_17_imag;
  assign io_coef_out_payload_0_18_18_real = int_reg_array_18_18_real;
  assign io_coef_out_payload_0_18_18_imag = int_reg_array_18_18_imag;
  assign io_coef_out_payload_0_18_19_real = int_reg_array_18_19_real;
  assign io_coef_out_payload_0_18_19_imag = int_reg_array_18_19_imag;
  assign io_coef_out_payload_0_18_20_real = int_reg_array_18_20_real;
  assign io_coef_out_payload_0_18_20_imag = int_reg_array_18_20_imag;
  assign io_coef_out_payload_0_18_21_real = int_reg_array_18_21_real;
  assign io_coef_out_payload_0_18_21_imag = int_reg_array_18_21_imag;
  assign io_coef_out_payload_0_18_22_real = int_reg_array_18_22_real;
  assign io_coef_out_payload_0_18_22_imag = int_reg_array_18_22_imag;
  assign io_coef_out_payload_0_18_23_real = int_reg_array_18_23_real;
  assign io_coef_out_payload_0_18_23_imag = int_reg_array_18_23_imag;
  assign io_coef_out_payload_0_18_24_real = int_reg_array_18_24_real;
  assign io_coef_out_payload_0_18_24_imag = int_reg_array_18_24_imag;
  assign io_coef_out_payload_0_18_25_real = int_reg_array_18_25_real;
  assign io_coef_out_payload_0_18_25_imag = int_reg_array_18_25_imag;
  assign io_coef_out_payload_0_18_26_real = int_reg_array_18_26_real;
  assign io_coef_out_payload_0_18_26_imag = int_reg_array_18_26_imag;
  assign io_coef_out_payload_0_18_27_real = int_reg_array_18_27_real;
  assign io_coef_out_payload_0_18_27_imag = int_reg_array_18_27_imag;
  assign io_coef_out_payload_0_18_28_real = int_reg_array_18_28_real;
  assign io_coef_out_payload_0_18_28_imag = int_reg_array_18_28_imag;
  assign io_coef_out_payload_0_18_29_real = int_reg_array_18_29_real;
  assign io_coef_out_payload_0_18_29_imag = int_reg_array_18_29_imag;
  assign io_coef_out_payload_0_18_30_real = int_reg_array_18_30_real;
  assign io_coef_out_payload_0_18_30_imag = int_reg_array_18_30_imag;
  assign io_coef_out_payload_0_18_31_real = int_reg_array_18_31_real;
  assign io_coef_out_payload_0_18_31_imag = int_reg_array_18_31_imag;
  assign io_coef_out_payload_0_18_32_real = int_reg_array_18_32_real;
  assign io_coef_out_payload_0_18_32_imag = int_reg_array_18_32_imag;
  assign io_coef_out_payload_0_18_33_real = int_reg_array_18_33_real;
  assign io_coef_out_payload_0_18_33_imag = int_reg_array_18_33_imag;
  assign io_coef_out_payload_0_18_34_real = int_reg_array_18_34_real;
  assign io_coef_out_payload_0_18_34_imag = int_reg_array_18_34_imag;
  assign io_coef_out_payload_0_18_35_real = int_reg_array_18_35_real;
  assign io_coef_out_payload_0_18_35_imag = int_reg_array_18_35_imag;
  assign io_coef_out_payload_0_18_36_real = int_reg_array_18_36_real;
  assign io_coef_out_payload_0_18_36_imag = int_reg_array_18_36_imag;
  assign io_coef_out_payload_0_18_37_real = int_reg_array_18_37_real;
  assign io_coef_out_payload_0_18_37_imag = int_reg_array_18_37_imag;
  assign io_coef_out_payload_0_18_38_real = int_reg_array_18_38_real;
  assign io_coef_out_payload_0_18_38_imag = int_reg_array_18_38_imag;
  assign io_coef_out_payload_0_18_39_real = int_reg_array_18_39_real;
  assign io_coef_out_payload_0_18_39_imag = int_reg_array_18_39_imag;
  assign io_coef_out_payload_0_18_40_real = int_reg_array_18_40_real;
  assign io_coef_out_payload_0_18_40_imag = int_reg_array_18_40_imag;
  assign io_coef_out_payload_0_18_41_real = int_reg_array_18_41_real;
  assign io_coef_out_payload_0_18_41_imag = int_reg_array_18_41_imag;
  assign io_coef_out_payload_0_18_42_real = int_reg_array_18_42_real;
  assign io_coef_out_payload_0_18_42_imag = int_reg_array_18_42_imag;
  assign io_coef_out_payload_0_18_43_real = int_reg_array_18_43_real;
  assign io_coef_out_payload_0_18_43_imag = int_reg_array_18_43_imag;
  assign io_coef_out_payload_0_18_44_real = int_reg_array_18_44_real;
  assign io_coef_out_payload_0_18_44_imag = int_reg_array_18_44_imag;
  assign io_coef_out_payload_0_18_45_real = int_reg_array_18_45_real;
  assign io_coef_out_payload_0_18_45_imag = int_reg_array_18_45_imag;
  assign io_coef_out_payload_0_18_46_real = int_reg_array_18_46_real;
  assign io_coef_out_payload_0_18_46_imag = int_reg_array_18_46_imag;
  assign io_coef_out_payload_0_18_47_real = int_reg_array_18_47_real;
  assign io_coef_out_payload_0_18_47_imag = int_reg_array_18_47_imag;
  assign io_coef_out_payload_0_18_48_real = int_reg_array_18_48_real;
  assign io_coef_out_payload_0_18_48_imag = int_reg_array_18_48_imag;
  assign io_coef_out_payload_0_18_49_real = int_reg_array_18_49_real;
  assign io_coef_out_payload_0_18_49_imag = int_reg_array_18_49_imag;
  assign io_coef_out_payload_0_19_0_real = int_reg_array_19_0_real;
  assign io_coef_out_payload_0_19_0_imag = int_reg_array_19_0_imag;
  assign io_coef_out_payload_0_19_1_real = int_reg_array_19_1_real;
  assign io_coef_out_payload_0_19_1_imag = int_reg_array_19_1_imag;
  assign io_coef_out_payload_0_19_2_real = int_reg_array_19_2_real;
  assign io_coef_out_payload_0_19_2_imag = int_reg_array_19_2_imag;
  assign io_coef_out_payload_0_19_3_real = int_reg_array_19_3_real;
  assign io_coef_out_payload_0_19_3_imag = int_reg_array_19_3_imag;
  assign io_coef_out_payload_0_19_4_real = int_reg_array_19_4_real;
  assign io_coef_out_payload_0_19_4_imag = int_reg_array_19_4_imag;
  assign io_coef_out_payload_0_19_5_real = int_reg_array_19_5_real;
  assign io_coef_out_payload_0_19_5_imag = int_reg_array_19_5_imag;
  assign io_coef_out_payload_0_19_6_real = int_reg_array_19_6_real;
  assign io_coef_out_payload_0_19_6_imag = int_reg_array_19_6_imag;
  assign io_coef_out_payload_0_19_7_real = int_reg_array_19_7_real;
  assign io_coef_out_payload_0_19_7_imag = int_reg_array_19_7_imag;
  assign io_coef_out_payload_0_19_8_real = int_reg_array_19_8_real;
  assign io_coef_out_payload_0_19_8_imag = int_reg_array_19_8_imag;
  assign io_coef_out_payload_0_19_9_real = int_reg_array_19_9_real;
  assign io_coef_out_payload_0_19_9_imag = int_reg_array_19_9_imag;
  assign io_coef_out_payload_0_19_10_real = int_reg_array_19_10_real;
  assign io_coef_out_payload_0_19_10_imag = int_reg_array_19_10_imag;
  assign io_coef_out_payload_0_19_11_real = int_reg_array_19_11_real;
  assign io_coef_out_payload_0_19_11_imag = int_reg_array_19_11_imag;
  assign io_coef_out_payload_0_19_12_real = int_reg_array_19_12_real;
  assign io_coef_out_payload_0_19_12_imag = int_reg_array_19_12_imag;
  assign io_coef_out_payload_0_19_13_real = int_reg_array_19_13_real;
  assign io_coef_out_payload_0_19_13_imag = int_reg_array_19_13_imag;
  assign io_coef_out_payload_0_19_14_real = int_reg_array_19_14_real;
  assign io_coef_out_payload_0_19_14_imag = int_reg_array_19_14_imag;
  assign io_coef_out_payload_0_19_15_real = int_reg_array_19_15_real;
  assign io_coef_out_payload_0_19_15_imag = int_reg_array_19_15_imag;
  assign io_coef_out_payload_0_19_16_real = int_reg_array_19_16_real;
  assign io_coef_out_payload_0_19_16_imag = int_reg_array_19_16_imag;
  assign io_coef_out_payload_0_19_17_real = int_reg_array_19_17_real;
  assign io_coef_out_payload_0_19_17_imag = int_reg_array_19_17_imag;
  assign io_coef_out_payload_0_19_18_real = int_reg_array_19_18_real;
  assign io_coef_out_payload_0_19_18_imag = int_reg_array_19_18_imag;
  assign io_coef_out_payload_0_19_19_real = int_reg_array_19_19_real;
  assign io_coef_out_payload_0_19_19_imag = int_reg_array_19_19_imag;
  assign io_coef_out_payload_0_19_20_real = int_reg_array_19_20_real;
  assign io_coef_out_payload_0_19_20_imag = int_reg_array_19_20_imag;
  assign io_coef_out_payload_0_19_21_real = int_reg_array_19_21_real;
  assign io_coef_out_payload_0_19_21_imag = int_reg_array_19_21_imag;
  assign io_coef_out_payload_0_19_22_real = int_reg_array_19_22_real;
  assign io_coef_out_payload_0_19_22_imag = int_reg_array_19_22_imag;
  assign io_coef_out_payload_0_19_23_real = int_reg_array_19_23_real;
  assign io_coef_out_payload_0_19_23_imag = int_reg_array_19_23_imag;
  assign io_coef_out_payload_0_19_24_real = int_reg_array_19_24_real;
  assign io_coef_out_payload_0_19_24_imag = int_reg_array_19_24_imag;
  assign io_coef_out_payload_0_19_25_real = int_reg_array_19_25_real;
  assign io_coef_out_payload_0_19_25_imag = int_reg_array_19_25_imag;
  assign io_coef_out_payload_0_19_26_real = int_reg_array_19_26_real;
  assign io_coef_out_payload_0_19_26_imag = int_reg_array_19_26_imag;
  assign io_coef_out_payload_0_19_27_real = int_reg_array_19_27_real;
  assign io_coef_out_payload_0_19_27_imag = int_reg_array_19_27_imag;
  assign io_coef_out_payload_0_19_28_real = int_reg_array_19_28_real;
  assign io_coef_out_payload_0_19_28_imag = int_reg_array_19_28_imag;
  assign io_coef_out_payload_0_19_29_real = int_reg_array_19_29_real;
  assign io_coef_out_payload_0_19_29_imag = int_reg_array_19_29_imag;
  assign io_coef_out_payload_0_19_30_real = int_reg_array_19_30_real;
  assign io_coef_out_payload_0_19_30_imag = int_reg_array_19_30_imag;
  assign io_coef_out_payload_0_19_31_real = int_reg_array_19_31_real;
  assign io_coef_out_payload_0_19_31_imag = int_reg_array_19_31_imag;
  assign io_coef_out_payload_0_19_32_real = int_reg_array_19_32_real;
  assign io_coef_out_payload_0_19_32_imag = int_reg_array_19_32_imag;
  assign io_coef_out_payload_0_19_33_real = int_reg_array_19_33_real;
  assign io_coef_out_payload_0_19_33_imag = int_reg_array_19_33_imag;
  assign io_coef_out_payload_0_19_34_real = int_reg_array_19_34_real;
  assign io_coef_out_payload_0_19_34_imag = int_reg_array_19_34_imag;
  assign io_coef_out_payload_0_19_35_real = int_reg_array_19_35_real;
  assign io_coef_out_payload_0_19_35_imag = int_reg_array_19_35_imag;
  assign io_coef_out_payload_0_19_36_real = int_reg_array_19_36_real;
  assign io_coef_out_payload_0_19_36_imag = int_reg_array_19_36_imag;
  assign io_coef_out_payload_0_19_37_real = int_reg_array_19_37_real;
  assign io_coef_out_payload_0_19_37_imag = int_reg_array_19_37_imag;
  assign io_coef_out_payload_0_19_38_real = int_reg_array_19_38_real;
  assign io_coef_out_payload_0_19_38_imag = int_reg_array_19_38_imag;
  assign io_coef_out_payload_0_19_39_real = int_reg_array_19_39_real;
  assign io_coef_out_payload_0_19_39_imag = int_reg_array_19_39_imag;
  assign io_coef_out_payload_0_19_40_real = int_reg_array_19_40_real;
  assign io_coef_out_payload_0_19_40_imag = int_reg_array_19_40_imag;
  assign io_coef_out_payload_0_19_41_real = int_reg_array_19_41_real;
  assign io_coef_out_payload_0_19_41_imag = int_reg_array_19_41_imag;
  assign io_coef_out_payload_0_19_42_real = int_reg_array_19_42_real;
  assign io_coef_out_payload_0_19_42_imag = int_reg_array_19_42_imag;
  assign io_coef_out_payload_0_19_43_real = int_reg_array_19_43_real;
  assign io_coef_out_payload_0_19_43_imag = int_reg_array_19_43_imag;
  assign io_coef_out_payload_0_19_44_real = int_reg_array_19_44_real;
  assign io_coef_out_payload_0_19_44_imag = int_reg_array_19_44_imag;
  assign io_coef_out_payload_0_19_45_real = int_reg_array_19_45_real;
  assign io_coef_out_payload_0_19_45_imag = int_reg_array_19_45_imag;
  assign io_coef_out_payload_0_19_46_real = int_reg_array_19_46_real;
  assign io_coef_out_payload_0_19_46_imag = int_reg_array_19_46_imag;
  assign io_coef_out_payload_0_19_47_real = int_reg_array_19_47_real;
  assign io_coef_out_payload_0_19_47_imag = int_reg_array_19_47_imag;
  assign io_coef_out_payload_0_19_48_real = int_reg_array_19_48_real;
  assign io_coef_out_payload_0_19_48_imag = int_reg_array_19_48_imag;
  assign io_coef_out_payload_0_19_49_real = int_reg_array_19_49_real;
  assign io_coef_out_payload_0_19_49_imag = int_reg_array_19_49_imag;
  assign io_coef_out_payload_0_20_0_real = int_reg_array_20_0_real;
  assign io_coef_out_payload_0_20_0_imag = int_reg_array_20_0_imag;
  assign io_coef_out_payload_0_20_1_real = int_reg_array_20_1_real;
  assign io_coef_out_payload_0_20_1_imag = int_reg_array_20_1_imag;
  assign io_coef_out_payload_0_20_2_real = int_reg_array_20_2_real;
  assign io_coef_out_payload_0_20_2_imag = int_reg_array_20_2_imag;
  assign io_coef_out_payload_0_20_3_real = int_reg_array_20_3_real;
  assign io_coef_out_payload_0_20_3_imag = int_reg_array_20_3_imag;
  assign io_coef_out_payload_0_20_4_real = int_reg_array_20_4_real;
  assign io_coef_out_payload_0_20_4_imag = int_reg_array_20_4_imag;
  assign io_coef_out_payload_0_20_5_real = int_reg_array_20_5_real;
  assign io_coef_out_payload_0_20_5_imag = int_reg_array_20_5_imag;
  assign io_coef_out_payload_0_20_6_real = int_reg_array_20_6_real;
  assign io_coef_out_payload_0_20_6_imag = int_reg_array_20_6_imag;
  assign io_coef_out_payload_0_20_7_real = int_reg_array_20_7_real;
  assign io_coef_out_payload_0_20_7_imag = int_reg_array_20_7_imag;
  assign io_coef_out_payload_0_20_8_real = int_reg_array_20_8_real;
  assign io_coef_out_payload_0_20_8_imag = int_reg_array_20_8_imag;
  assign io_coef_out_payload_0_20_9_real = int_reg_array_20_9_real;
  assign io_coef_out_payload_0_20_9_imag = int_reg_array_20_9_imag;
  assign io_coef_out_payload_0_20_10_real = int_reg_array_20_10_real;
  assign io_coef_out_payload_0_20_10_imag = int_reg_array_20_10_imag;
  assign io_coef_out_payload_0_20_11_real = int_reg_array_20_11_real;
  assign io_coef_out_payload_0_20_11_imag = int_reg_array_20_11_imag;
  assign io_coef_out_payload_0_20_12_real = int_reg_array_20_12_real;
  assign io_coef_out_payload_0_20_12_imag = int_reg_array_20_12_imag;
  assign io_coef_out_payload_0_20_13_real = int_reg_array_20_13_real;
  assign io_coef_out_payload_0_20_13_imag = int_reg_array_20_13_imag;
  assign io_coef_out_payload_0_20_14_real = int_reg_array_20_14_real;
  assign io_coef_out_payload_0_20_14_imag = int_reg_array_20_14_imag;
  assign io_coef_out_payload_0_20_15_real = int_reg_array_20_15_real;
  assign io_coef_out_payload_0_20_15_imag = int_reg_array_20_15_imag;
  assign io_coef_out_payload_0_20_16_real = int_reg_array_20_16_real;
  assign io_coef_out_payload_0_20_16_imag = int_reg_array_20_16_imag;
  assign io_coef_out_payload_0_20_17_real = int_reg_array_20_17_real;
  assign io_coef_out_payload_0_20_17_imag = int_reg_array_20_17_imag;
  assign io_coef_out_payload_0_20_18_real = int_reg_array_20_18_real;
  assign io_coef_out_payload_0_20_18_imag = int_reg_array_20_18_imag;
  assign io_coef_out_payload_0_20_19_real = int_reg_array_20_19_real;
  assign io_coef_out_payload_0_20_19_imag = int_reg_array_20_19_imag;
  assign io_coef_out_payload_0_20_20_real = int_reg_array_20_20_real;
  assign io_coef_out_payload_0_20_20_imag = int_reg_array_20_20_imag;
  assign io_coef_out_payload_0_20_21_real = int_reg_array_20_21_real;
  assign io_coef_out_payload_0_20_21_imag = int_reg_array_20_21_imag;
  assign io_coef_out_payload_0_20_22_real = int_reg_array_20_22_real;
  assign io_coef_out_payload_0_20_22_imag = int_reg_array_20_22_imag;
  assign io_coef_out_payload_0_20_23_real = int_reg_array_20_23_real;
  assign io_coef_out_payload_0_20_23_imag = int_reg_array_20_23_imag;
  assign io_coef_out_payload_0_20_24_real = int_reg_array_20_24_real;
  assign io_coef_out_payload_0_20_24_imag = int_reg_array_20_24_imag;
  assign io_coef_out_payload_0_20_25_real = int_reg_array_20_25_real;
  assign io_coef_out_payload_0_20_25_imag = int_reg_array_20_25_imag;
  assign io_coef_out_payload_0_20_26_real = int_reg_array_20_26_real;
  assign io_coef_out_payload_0_20_26_imag = int_reg_array_20_26_imag;
  assign io_coef_out_payload_0_20_27_real = int_reg_array_20_27_real;
  assign io_coef_out_payload_0_20_27_imag = int_reg_array_20_27_imag;
  assign io_coef_out_payload_0_20_28_real = int_reg_array_20_28_real;
  assign io_coef_out_payload_0_20_28_imag = int_reg_array_20_28_imag;
  assign io_coef_out_payload_0_20_29_real = int_reg_array_20_29_real;
  assign io_coef_out_payload_0_20_29_imag = int_reg_array_20_29_imag;
  assign io_coef_out_payload_0_20_30_real = int_reg_array_20_30_real;
  assign io_coef_out_payload_0_20_30_imag = int_reg_array_20_30_imag;
  assign io_coef_out_payload_0_20_31_real = int_reg_array_20_31_real;
  assign io_coef_out_payload_0_20_31_imag = int_reg_array_20_31_imag;
  assign io_coef_out_payload_0_20_32_real = int_reg_array_20_32_real;
  assign io_coef_out_payload_0_20_32_imag = int_reg_array_20_32_imag;
  assign io_coef_out_payload_0_20_33_real = int_reg_array_20_33_real;
  assign io_coef_out_payload_0_20_33_imag = int_reg_array_20_33_imag;
  assign io_coef_out_payload_0_20_34_real = int_reg_array_20_34_real;
  assign io_coef_out_payload_0_20_34_imag = int_reg_array_20_34_imag;
  assign io_coef_out_payload_0_20_35_real = int_reg_array_20_35_real;
  assign io_coef_out_payload_0_20_35_imag = int_reg_array_20_35_imag;
  assign io_coef_out_payload_0_20_36_real = int_reg_array_20_36_real;
  assign io_coef_out_payload_0_20_36_imag = int_reg_array_20_36_imag;
  assign io_coef_out_payload_0_20_37_real = int_reg_array_20_37_real;
  assign io_coef_out_payload_0_20_37_imag = int_reg_array_20_37_imag;
  assign io_coef_out_payload_0_20_38_real = int_reg_array_20_38_real;
  assign io_coef_out_payload_0_20_38_imag = int_reg_array_20_38_imag;
  assign io_coef_out_payload_0_20_39_real = int_reg_array_20_39_real;
  assign io_coef_out_payload_0_20_39_imag = int_reg_array_20_39_imag;
  assign io_coef_out_payload_0_20_40_real = int_reg_array_20_40_real;
  assign io_coef_out_payload_0_20_40_imag = int_reg_array_20_40_imag;
  assign io_coef_out_payload_0_20_41_real = int_reg_array_20_41_real;
  assign io_coef_out_payload_0_20_41_imag = int_reg_array_20_41_imag;
  assign io_coef_out_payload_0_20_42_real = int_reg_array_20_42_real;
  assign io_coef_out_payload_0_20_42_imag = int_reg_array_20_42_imag;
  assign io_coef_out_payload_0_20_43_real = int_reg_array_20_43_real;
  assign io_coef_out_payload_0_20_43_imag = int_reg_array_20_43_imag;
  assign io_coef_out_payload_0_20_44_real = int_reg_array_20_44_real;
  assign io_coef_out_payload_0_20_44_imag = int_reg_array_20_44_imag;
  assign io_coef_out_payload_0_20_45_real = int_reg_array_20_45_real;
  assign io_coef_out_payload_0_20_45_imag = int_reg_array_20_45_imag;
  assign io_coef_out_payload_0_20_46_real = int_reg_array_20_46_real;
  assign io_coef_out_payload_0_20_46_imag = int_reg_array_20_46_imag;
  assign io_coef_out_payload_0_20_47_real = int_reg_array_20_47_real;
  assign io_coef_out_payload_0_20_47_imag = int_reg_array_20_47_imag;
  assign io_coef_out_payload_0_20_48_real = int_reg_array_20_48_real;
  assign io_coef_out_payload_0_20_48_imag = int_reg_array_20_48_imag;
  assign io_coef_out_payload_0_20_49_real = int_reg_array_20_49_real;
  assign io_coef_out_payload_0_20_49_imag = int_reg_array_20_49_imag;
  assign io_coef_out_payload_0_21_0_real = int_reg_array_21_0_real;
  assign io_coef_out_payload_0_21_0_imag = int_reg_array_21_0_imag;
  assign io_coef_out_payload_0_21_1_real = int_reg_array_21_1_real;
  assign io_coef_out_payload_0_21_1_imag = int_reg_array_21_1_imag;
  assign io_coef_out_payload_0_21_2_real = int_reg_array_21_2_real;
  assign io_coef_out_payload_0_21_2_imag = int_reg_array_21_2_imag;
  assign io_coef_out_payload_0_21_3_real = int_reg_array_21_3_real;
  assign io_coef_out_payload_0_21_3_imag = int_reg_array_21_3_imag;
  assign io_coef_out_payload_0_21_4_real = int_reg_array_21_4_real;
  assign io_coef_out_payload_0_21_4_imag = int_reg_array_21_4_imag;
  assign io_coef_out_payload_0_21_5_real = int_reg_array_21_5_real;
  assign io_coef_out_payload_0_21_5_imag = int_reg_array_21_5_imag;
  assign io_coef_out_payload_0_21_6_real = int_reg_array_21_6_real;
  assign io_coef_out_payload_0_21_6_imag = int_reg_array_21_6_imag;
  assign io_coef_out_payload_0_21_7_real = int_reg_array_21_7_real;
  assign io_coef_out_payload_0_21_7_imag = int_reg_array_21_7_imag;
  assign io_coef_out_payload_0_21_8_real = int_reg_array_21_8_real;
  assign io_coef_out_payload_0_21_8_imag = int_reg_array_21_8_imag;
  assign io_coef_out_payload_0_21_9_real = int_reg_array_21_9_real;
  assign io_coef_out_payload_0_21_9_imag = int_reg_array_21_9_imag;
  assign io_coef_out_payload_0_21_10_real = int_reg_array_21_10_real;
  assign io_coef_out_payload_0_21_10_imag = int_reg_array_21_10_imag;
  assign io_coef_out_payload_0_21_11_real = int_reg_array_21_11_real;
  assign io_coef_out_payload_0_21_11_imag = int_reg_array_21_11_imag;
  assign io_coef_out_payload_0_21_12_real = int_reg_array_21_12_real;
  assign io_coef_out_payload_0_21_12_imag = int_reg_array_21_12_imag;
  assign io_coef_out_payload_0_21_13_real = int_reg_array_21_13_real;
  assign io_coef_out_payload_0_21_13_imag = int_reg_array_21_13_imag;
  assign io_coef_out_payload_0_21_14_real = int_reg_array_21_14_real;
  assign io_coef_out_payload_0_21_14_imag = int_reg_array_21_14_imag;
  assign io_coef_out_payload_0_21_15_real = int_reg_array_21_15_real;
  assign io_coef_out_payload_0_21_15_imag = int_reg_array_21_15_imag;
  assign io_coef_out_payload_0_21_16_real = int_reg_array_21_16_real;
  assign io_coef_out_payload_0_21_16_imag = int_reg_array_21_16_imag;
  assign io_coef_out_payload_0_21_17_real = int_reg_array_21_17_real;
  assign io_coef_out_payload_0_21_17_imag = int_reg_array_21_17_imag;
  assign io_coef_out_payload_0_21_18_real = int_reg_array_21_18_real;
  assign io_coef_out_payload_0_21_18_imag = int_reg_array_21_18_imag;
  assign io_coef_out_payload_0_21_19_real = int_reg_array_21_19_real;
  assign io_coef_out_payload_0_21_19_imag = int_reg_array_21_19_imag;
  assign io_coef_out_payload_0_21_20_real = int_reg_array_21_20_real;
  assign io_coef_out_payload_0_21_20_imag = int_reg_array_21_20_imag;
  assign io_coef_out_payload_0_21_21_real = int_reg_array_21_21_real;
  assign io_coef_out_payload_0_21_21_imag = int_reg_array_21_21_imag;
  assign io_coef_out_payload_0_21_22_real = int_reg_array_21_22_real;
  assign io_coef_out_payload_0_21_22_imag = int_reg_array_21_22_imag;
  assign io_coef_out_payload_0_21_23_real = int_reg_array_21_23_real;
  assign io_coef_out_payload_0_21_23_imag = int_reg_array_21_23_imag;
  assign io_coef_out_payload_0_21_24_real = int_reg_array_21_24_real;
  assign io_coef_out_payload_0_21_24_imag = int_reg_array_21_24_imag;
  assign io_coef_out_payload_0_21_25_real = int_reg_array_21_25_real;
  assign io_coef_out_payload_0_21_25_imag = int_reg_array_21_25_imag;
  assign io_coef_out_payload_0_21_26_real = int_reg_array_21_26_real;
  assign io_coef_out_payload_0_21_26_imag = int_reg_array_21_26_imag;
  assign io_coef_out_payload_0_21_27_real = int_reg_array_21_27_real;
  assign io_coef_out_payload_0_21_27_imag = int_reg_array_21_27_imag;
  assign io_coef_out_payload_0_21_28_real = int_reg_array_21_28_real;
  assign io_coef_out_payload_0_21_28_imag = int_reg_array_21_28_imag;
  assign io_coef_out_payload_0_21_29_real = int_reg_array_21_29_real;
  assign io_coef_out_payload_0_21_29_imag = int_reg_array_21_29_imag;
  assign io_coef_out_payload_0_21_30_real = int_reg_array_21_30_real;
  assign io_coef_out_payload_0_21_30_imag = int_reg_array_21_30_imag;
  assign io_coef_out_payload_0_21_31_real = int_reg_array_21_31_real;
  assign io_coef_out_payload_0_21_31_imag = int_reg_array_21_31_imag;
  assign io_coef_out_payload_0_21_32_real = int_reg_array_21_32_real;
  assign io_coef_out_payload_0_21_32_imag = int_reg_array_21_32_imag;
  assign io_coef_out_payload_0_21_33_real = int_reg_array_21_33_real;
  assign io_coef_out_payload_0_21_33_imag = int_reg_array_21_33_imag;
  assign io_coef_out_payload_0_21_34_real = int_reg_array_21_34_real;
  assign io_coef_out_payload_0_21_34_imag = int_reg_array_21_34_imag;
  assign io_coef_out_payload_0_21_35_real = int_reg_array_21_35_real;
  assign io_coef_out_payload_0_21_35_imag = int_reg_array_21_35_imag;
  assign io_coef_out_payload_0_21_36_real = int_reg_array_21_36_real;
  assign io_coef_out_payload_0_21_36_imag = int_reg_array_21_36_imag;
  assign io_coef_out_payload_0_21_37_real = int_reg_array_21_37_real;
  assign io_coef_out_payload_0_21_37_imag = int_reg_array_21_37_imag;
  assign io_coef_out_payload_0_21_38_real = int_reg_array_21_38_real;
  assign io_coef_out_payload_0_21_38_imag = int_reg_array_21_38_imag;
  assign io_coef_out_payload_0_21_39_real = int_reg_array_21_39_real;
  assign io_coef_out_payload_0_21_39_imag = int_reg_array_21_39_imag;
  assign io_coef_out_payload_0_21_40_real = int_reg_array_21_40_real;
  assign io_coef_out_payload_0_21_40_imag = int_reg_array_21_40_imag;
  assign io_coef_out_payload_0_21_41_real = int_reg_array_21_41_real;
  assign io_coef_out_payload_0_21_41_imag = int_reg_array_21_41_imag;
  assign io_coef_out_payload_0_21_42_real = int_reg_array_21_42_real;
  assign io_coef_out_payload_0_21_42_imag = int_reg_array_21_42_imag;
  assign io_coef_out_payload_0_21_43_real = int_reg_array_21_43_real;
  assign io_coef_out_payload_0_21_43_imag = int_reg_array_21_43_imag;
  assign io_coef_out_payload_0_21_44_real = int_reg_array_21_44_real;
  assign io_coef_out_payload_0_21_44_imag = int_reg_array_21_44_imag;
  assign io_coef_out_payload_0_21_45_real = int_reg_array_21_45_real;
  assign io_coef_out_payload_0_21_45_imag = int_reg_array_21_45_imag;
  assign io_coef_out_payload_0_21_46_real = int_reg_array_21_46_real;
  assign io_coef_out_payload_0_21_46_imag = int_reg_array_21_46_imag;
  assign io_coef_out_payload_0_21_47_real = int_reg_array_21_47_real;
  assign io_coef_out_payload_0_21_47_imag = int_reg_array_21_47_imag;
  assign io_coef_out_payload_0_21_48_real = int_reg_array_21_48_real;
  assign io_coef_out_payload_0_21_48_imag = int_reg_array_21_48_imag;
  assign io_coef_out_payload_0_21_49_real = int_reg_array_21_49_real;
  assign io_coef_out_payload_0_21_49_imag = int_reg_array_21_49_imag;
  assign io_coef_out_payload_0_22_0_real = int_reg_array_22_0_real;
  assign io_coef_out_payload_0_22_0_imag = int_reg_array_22_0_imag;
  assign io_coef_out_payload_0_22_1_real = int_reg_array_22_1_real;
  assign io_coef_out_payload_0_22_1_imag = int_reg_array_22_1_imag;
  assign io_coef_out_payload_0_22_2_real = int_reg_array_22_2_real;
  assign io_coef_out_payload_0_22_2_imag = int_reg_array_22_2_imag;
  assign io_coef_out_payload_0_22_3_real = int_reg_array_22_3_real;
  assign io_coef_out_payload_0_22_3_imag = int_reg_array_22_3_imag;
  assign io_coef_out_payload_0_22_4_real = int_reg_array_22_4_real;
  assign io_coef_out_payload_0_22_4_imag = int_reg_array_22_4_imag;
  assign io_coef_out_payload_0_22_5_real = int_reg_array_22_5_real;
  assign io_coef_out_payload_0_22_5_imag = int_reg_array_22_5_imag;
  assign io_coef_out_payload_0_22_6_real = int_reg_array_22_6_real;
  assign io_coef_out_payload_0_22_6_imag = int_reg_array_22_6_imag;
  assign io_coef_out_payload_0_22_7_real = int_reg_array_22_7_real;
  assign io_coef_out_payload_0_22_7_imag = int_reg_array_22_7_imag;
  assign io_coef_out_payload_0_22_8_real = int_reg_array_22_8_real;
  assign io_coef_out_payload_0_22_8_imag = int_reg_array_22_8_imag;
  assign io_coef_out_payload_0_22_9_real = int_reg_array_22_9_real;
  assign io_coef_out_payload_0_22_9_imag = int_reg_array_22_9_imag;
  assign io_coef_out_payload_0_22_10_real = int_reg_array_22_10_real;
  assign io_coef_out_payload_0_22_10_imag = int_reg_array_22_10_imag;
  assign io_coef_out_payload_0_22_11_real = int_reg_array_22_11_real;
  assign io_coef_out_payload_0_22_11_imag = int_reg_array_22_11_imag;
  assign io_coef_out_payload_0_22_12_real = int_reg_array_22_12_real;
  assign io_coef_out_payload_0_22_12_imag = int_reg_array_22_12_imag;
  assign io_coef_out_payload_0_22_13_real = int_reg_array_22_13_real;
  assign io_coef_out_payload_0_22_13_imag = int_reg_array_22_13_imag;
  assign io_coef_out_payload_0_22_14_real = int_reg_array_22_14_real;
  assign io_coef_out_payload_0_22_14_imag = int_reg_array_22_14_imag;
  assign io_coef_out_payload_0_22_15_real = int_reg_array_22_15_real;
  assign io_coef_out_payload_0_22_15_imag = int_reg_array_22_15_imag;
  assign io_coef_out_payload_0_22_16_real = int_reg_array_22_16_real;
  assign io_coef_out_payload_0_22_16_imag = int_reg_array_22_16_imag;
  assign io_coef_out_payload_0_22_17_real = int_reg_array_22_17_real;
  assign io_coef_out_payload_0_22_17_imag = int_reg_array_22_17_imag;
  assign io_coef_out_payload_0_22_18_real = int_reg_array_22_18_real;
  assign io_coef_out_payload_0_22_18_imag = int_reg_array_22_18_imag;
  assign io_coef_out_payload_0_22_19_real = int_reg_array_22_19_real;
  assign io_coef_out_payload_0_22_19_imag = int_reg_array_22_19_imag;
  assign io_coef_out_payload_0_22_20_real = int_reg_array_22_20_real;
  assign io_coef_out_payload_0_22_20_imag = int_reg_array_22_20_imag;
  assign io_coef_out_payload_0_22_21_real = int_reg_array_22_21_real;
  assign io_coef_out_payload_0_22_21_imag = int_reg_array_22_21_imag;
  assign io_coef_out_payload_0_22_22_real = int_reg_array_22_22_real;
  assign io_coef_out_payload_0_22_22_imag = int_reg_array_22_22_imag;
  assign io_coef_out_payload_0_22_23_real = int_reg_array_22_23_real;
  assign io_coef_out_payload_0_22_23_imag = int_reg_array_22_23_imag;
  assign io_coef_out_payload_0_22_24_real = int_reg_array_22_24_real;
  assign io_coef_out_payload_0_22_24_imag = int_reg_array_22_24_imag;
  assign io_coef_out_payload_0_22_25_real = int_reg_array_22_25_real;
  assign io_coef_out_payload_0_22_25_imag = int_reg_array_22_25_imag;
  assign io_coef_out_payload_0_22_26_real = int_reg_array_22_26_real;
  assign io_coef_out_payload_0_22_26_imag = int_reg_array_22_26_imag;
  assign io_coef_out_payload_0_22_27_real = int_reg_array_22_27_real;
  assign io_coef_out_payload_0_22_27_imag = int_reg_array_22_27_imag;
  assign io_coef_out_payload_0_22_28_real = int_reg_array_22_28_real;
  assign io_coef_out_payload_0_22_28_imag = int_reg_array_22_28_imag;
  assign io_coef_out_payload_0_22_29_real = int_reg_array_22_29_real;
  assign io_coef_out_payload_0_22_29_imag = int_reg_array_22_29_imag;
  assign io_coef_out_payload_0_22_30_real = int_reg_array_22_30_real;
  assign io_coef_out_payload_0_22_30_imag = int_reg_array_22_30_imag;
  assign io_coef_out_payload_0_22_31_real = int_reg_array_22_31_real;
  assign io_coef_out_payload_0_22_31_imag = int_reg_array_22_31_imag;
  assign io_coef_out_payload_0_22_32_real = int_reg_array_22_32_real;
  assign io_coef_out_payload_0_22_32_imag = int_reg_array_22_32_imag;
  assign io_coef_out_payload_0_22_33_real = int_reg_array_22_33_real;
  assign io_coef_out_payload_0_22_33_imag = int_reg_array_22_33_imag;
  assign io_coef_out_payload_0_22_34_real = int_reg_array_22_34_real;
  assign io_coef_out_payload_0_22_34_imag = int_reg_array_22_34_imag;
  assign io_coef_out_payload_0_22_35_real = int_reg_array_22_35_real;
  assign io_coef_out_payload_0_22_35_imag = int_reg_array_22_35_imag;
  assign io_coef_out_payload_0_22_36_real = int_reg_array_22_36_real;
  assign io_coef_out_payload_0_22_36_imag = int_reg_array_22_36_imag;
  assign io_coef_out_payload_0_22_37_real = int_reg_array_22_37_real;
  assign io_coef_out_payload_0_22_37_imag = int_reg_array_22_37_imag;
  assign io_coef_out_payload_0_22_38_real = int_reg_array_22_38_real;
  assign io_coef_out_payload_0_22_38_imag = int_reg_array_22_38_imag;
  assign io_coef_out_payload_0_22_39_real = int_reg_array_22_39_real;
  assign io_coef_out_payload_0_22_39_imag = int_reg_array_22_39_imag;
  assign io_coef_out_payload_0_22_40_real = int_reg_array_22_40_real;
  assign io_coef_out_payload_0_22_40_imag = int_reg_array_22_40_imag;
  assign io_coef_out_payload_0_22_41_real = int_reg_array_22_41_real;
  assign io_coef_out_payload_0_22_41_imag = int_reg_array_22_41_imag;
  assign io_coef_out_payload_0_22_42_real = int_reg_array_22_42_real;
  assign io_coef_out_payload_0_22_42_imag = int_reg_array_22_42_imag;
  assign io_coef_out_payload_0_22_43_real = int_reg_array_22_43_real;
  assign io_coef_out_payload_0_22_43_imag = int_reg_array_22_43_imag;
  assign io_coef_out_payload_0_22_44_real = int_reg_array_22_44_real;
  assign io_coef_out_payload_0_22_44_imag = int_reg_array_22_44_imag;
  assign io_coef_out_payload_0_22_45_real = int_reg_array_22_45_real;
  assign io_coef_out_payload_0_22_45_imag = int_reg_array_22_45_imag;
  assign io_coef_out_payload_0_22_46_real = int_reg_array_22_46_real;
  assign io_coef_out_payload_0_22_46_imag = int_reg_array_22_46_imag;
  assign io_coef_out_payload_0_22_47_real = int_reg_array_22_47_real;
  assign io_coef_out_payload_0_22_47_imag = int_reg_array_22_47_imag;
  assign io_coef_out_payload_0_22_48_real = int_reg_array_22_48_real;
  assign io_coef_out_payload_0_22_48_imag = int_reg_array_22_48_imag;
  assign io_coef_out_payload_0_22_49_real = int_reg_array_22_49_real;
  assign io_coef_out_payload_0_22_49_imag = int_reg_array_22_49_imag;
  assign io_coef_out_payload_0_23_0_real = int_reg_array_23_0_real;
  assign io_coef_out_payload_0_23_0_imag = int_reg_array_23_0_imag;
  assign io_coef_out_payload_0_23_1_real = int_reg_array_23_1_real;
  assign io_coef_out_payload_0_23_1_imag = int_reg_array_23_1_imag;
  assign io_coef_out_payload_0_23_2_real = int_reg_array_23_2_real;
  assign io_coef_out_payload_0_23_2_imag = int_reg_array_23_2_imag;
  assign io_coef_out_payload_0_23_3_real = int_reg_array_23_3_real;
  assign io_coef_out_payload_0_23_3_imag = int_reg_array_23_3_imag;
  assign io_coef_out_payload_0_23_4_real = int_reg_array_23_4_real;
  assign io_coef_out_payload_0_23_4_imag = int_reg_array_23_4_imag;
  assign io_coef_out_payload_0_23_5_real = int_reg_array_23_5_real;
  assign io_coef_out_payload_0_23_5_imag = int_reg_array_23_5_imag;
  assign io_coef_out_payload_0_23_6_real = int_reg_array_23_6_real;
  assign io_coef_out_payload_0_23_6_imag = int_reg_array_23_6_imag;
  assign io_coef_out_payload_0_23_7_real = int_reg_array_23_7_real;
  assign io_coef_out_payload_0_23_7_imag = int_reg_array_23_7_imag;
  assign io_coef_out_payload_0_23_8_real = int_reg_array_23_8_real;
  assign io_coef_out_payload_0_23_8_imag = int_reg_array_23_8_imag;
  assign io_coef_out_payload_0_23_9_real = int_reg_array_23_9_real;
  assign io_coef_out_payload_0_23_9_imag = int_reg_array_23_9_imag;
  assign io_coef_out_payload_0_23_10_real = int_reg_array_23_10_real;
  assign io_coef_out_payload_0_23_10_imag = int_reg_array_23_10_imag;
  assign io_coef_out_payload_0_23_11_real = int_reg_array_23_11_real;
  assign io_coef_out_payload_0_23_11_imag = int_reg_array_23_11_imag;
  assign io_coef_out_payload_0_23_12_real = int_reg_array_23_12_real;
  assign io_coef_out_payload_0_23_12_imag = int_reg_array_23_12_imag;
  assign io_coef_out_payload_0_23_13_real = int_reg_array_23_13_real;
  assign io_coef_out_payload_0_23_13_imag = int_reg_array_23_13_imag;
  assign io_coef_out_payload_0_23_14_real = int_reg_array_23_14_real;
  assign io_coef_out_payload_0_23_14_imag = int_reg_array_23_14_imag;
  assign io_coef_out_payload_0_23_15_real = int_reg_array_23_15_real;
  assign io_coef_out_payload_0_23_15_imag = int_reg_array_23_15_imag;
  assign io_coef_out_payload_0_23_16_real = int_reg_array_23_16_real;
  assign io_coef_out_payload_0_23_16_imag = int_reg_array_23_16_imag;
  assign io_coef_out_payload_0_23_17_real = int_reg_array_23_17_real;
  assign io_coef_out_payload_0_23_17_imag = int_reg_array_23_17_imag;
  assign io_coef_out_payload_0_23_18_real = int_reg_array_23_18_real;
  assign io_coef_out_payload_0_23_18_imag = int_reg_array_23_18_imag;
  assign io_coef_out_payload_0_23_19_real = int_reg_array_23_19_real;
  assign io_coef_out_payload_0_23_19_imag = int_reg_array_23_19_imag;
  assign io_coef_out_payload_0_23_20_real = int_reg_array_23_20_real;
  assign io_coef_out_payload_0_23_20_imag = int_reg_array_23_20_imag;
  assign io_coef_out_payload_0_23_21_real = int_reg_array_23_21_real;
  assign io_coef_out_payload_0_23_21_imag = int_reg_array_23_21_imag;
  assign io_coef_out_payload_0_23_22_real = int_reg_array_23_22_real;
  assign io_coef_out_payload_0_23_22_imag = int_reg_array_23_22_imag;
  assign io_coef_out_payload_0_23_23_real = int_reg_array_23_23_real;
  assign io_coef_out_payload_0_23_23_imag = int_reg_array_23_23_imag;
  assign io_coef_out_payload_0_23_24_real = int_reg_array_23_24_real;
  assign io_coef_out_payload_0_23_24_imag = int_reg_array_23_24_imag;
  assign io_coef_out_payload_0_23_25_real = int_reg_array_23_25_real;
  assign io_coef_out_payload_0_23_25_imag = int_reg_array_23_25_imag;
  assign io_coef_out_payload_0_23_26_real = int_reg_array_23_26_real;
  assign io_coef_out_payload_0_23_26_imag = int_reg_array_23_26_imag;
  assign io_coef_out_payload_0_23_27_real = int_reg_array_23_27_real;
  assign io_coef_out_payload_0_23_27_imag = int_reg_array_23_27_imag;
  assign io_coef_out_payload_0_23_28_real = int_reg_array_23_28_real;
  assign io_coef_out_payload_0_23_28_imag = int_reg_array_23_28_imag;
  assign io_coef_out_payload_0_23_29_real = int_reg_array_23_29_real;
  assign io_coef_out_payload_0_23_29_imag = int_reg_array_23_29_imag;
  assign io_coef_out_payload_0_23_30_real = int_reg_array_23_30_real;
  assign io_coef_out_payload_0_23_30_imag = int_reg_array_23_30_imag;
  assign io_coef_out_payload_0_23_31_real = int_reg_array_23_31_real;
  assign io_coef_out_payload_0_23_31_imag = int_reg_array_23_31_imag;
  assign io_coef_out_payload_0_23_32_real = int_reg_array_23_32_real;
  assign io_coef_out_payload_0_23_32_imag = int_reg_array_23_32_imag;
  assign io_coef_out_payload_0_23_33_real = int_reg_array_23_33_real;
  assign io_coef_out_payload_0_23_33_imag = int_reg_array_23_33_imag;
  assign io_coef_out_payload_0_23_34_real = int_reg_array_23_34_real;
  assign io_coef_out_payload_0_23_34_imag = int_reg_array_23_34_imag;
  assign io_coef_out_payload_0_23_35_real = int_reg_array_23_35_real;
  assign io_coef_out_payload_0_23_35_imag = int_reg_array_23_35_imag;
  assign io_coef_out_payload_0_23_36_real = int_reg_array_23_36_real;
  assign io_coef_out_payload_0_23_36_imag = int_reg_array_23_36_imag;
  assign io_coef_out_payload_0_23_37_real = int_reg_array_23_37_real;
  assign io_coef_out_payload_0_23_37_imag = int_reg_array_23_37_imag;
  assign io_coef_out_payload_0_23_38_real = int_reg_array_23_38_real;
  assign io_coef_out_payload_0_23_38_imag = int_reg_array_23_38_imag;
  assign io_coef_out_payload_0_23_39_real = int_reg_array_23_39_real;
  assign io_coef_out_payload_0_23_39_imag = int_reg_array_23_39_imag;
  assign io_coef_out_payload_0_23_40_real = int_reg_array_23_40_real;
  assign io_coef_out_payload_0_23_40_imag = int_reg_array_23_40_imag;
  assign io_coef_out_payload_0_23_41_real = int_reg_array_23_41_real;
  assign io_coef_out_payload_0_23_41_imag = int_reg_array_23_41_imag;
  assign io_coef_out_payload_0_23_42_real = int_reg_array_23_42_real;
  assign io_coef_out_payload_0_23_42_imag = int_reg_array_23_42_imag;
  assign io_coef_out_payload_0_23_43_real = int_reg_array_23_43_real;
  assign io_coef_out_payload_0_23_43_imag = int_reg_array_23_43_imag;
  assign io_coef_out_payload_0_23_44_real = int_reg_array_23_44_real;
  assign io_coef_out_payload_0_23_44_imag = int_reg_array_23_44_imag;
  assign io_coef_out_payload_0_23_45_real = int_reg_array_23_45_real;
  assign io_coef_out_payload_0_23_45_imag = int_reg_array_23_45_imag;
  assign io_coef_out_payload_0_23_46_real = int_reg_array_23_46_real;
  assign io_coef_out_payload_0_23_46_imag = int_reg_array_23_46_imag;
  assign io_coef_out_payload_0_23_47_real = int_reg_array_23_47_real;
  assign io_coef_out_payload_0_23_47_imag = int_reg_array_23_47_imag;
  assign io_coef_out_payload_0_23_48_real = int_reg_array_23_48_real;
  assign io_coef_out_payload_0_23_48_imag = int_reg_array_23_48_imag;
  assign io_coef_out_payload_0_23_49_real = int_reg_array_23_49_real;
  assign io_coef_out_payload_0_23_49_imag = int_reg_array_23_49_imag;
  assign io_coef_out_payload_0_24_0_real = int_reg_array_24_0_real;
  assign io_coef_out_payload_0_24_0_imag = int_reg_array_24_0_imag;
  assign io_coef_out_payload_0_24_1_real = int_reg_array_24_1_real;
  assign io_coef_out_payload_0_24_1_imag = int_reg_array_24_1_imag;
  assign io_coef_out_payload_0_24_2_real = int_reg_array_24_2_real;
  assign io_coef_out_payload_0_24_2_imag = int_reg_array_24_2_imag;
  assign io_coef_out_payload_0_24_3_real = int_reg_array_24_3_real;
  assign io_coef_out_payload_0_24_3_imag = int_reg_array_24_3_imag;
  assign io_coef_out_payload_0_24_4_real = int_reg_array_24_4_real;
  assign io_coef_out_payload_0_24_4_imag = int_reg_array_24_4_imag;
  assign io_coef_out_payload_0_24_5_real = int_reg_array_24_5_real;
  assign io_coef_out_payload_0_24_5_imag = int_reg_array_24_5_imag;
  assign io_coef_out_payload_0_24_6_real = int_reg_array_24_6_real;
  assign io_coef_out_payload_0_24_6_imag = int_reg_array_24_6_imag;
  assign io_coef_out_payload_0_24_7_real = int_reg_array_24_7_real;
  assign io_coef_out_payload_0_24_7_imag = int_reg_array_24_7_imag;
  assign io_coef_out_payload_0_24_8_real = int_reg_array_24_8_real;
  assign io_coef_out_payload_0_24_8_imag = int_reg_array_24_8_imag;
  assign io_coef_out_payload_0_24_9_real = int_reg_array_24_9_real;
  assign io_coef_out_payload_0_24_9_imag = int_reg_array_24_9_imag;
  assign io_coef_out_payload_0_24_10_real = int_reg_array_24_10_real;
  assign io_coef_out_payload_0_24_10_imag = int_reg_array_24_10_imag;
  assign io_coef_out_payload_0_24_11_real = int_reg_array_24_11_real;
  assign io_coef_out_payload_0_24_11_imag = int_reg_array_24_11_imag;
  assign io_coef_out_payload_0_24_12_real = int_reg_array_24_12_real;
  assign io_coef_out_payload_0_24_12_imag = int_reg_array_24_12_imag;
  assign io_coef_out_payload_0_24_13_real = int_reg_array_24_13_real;
  assign io_coef_out_payload_0_24_13_imag = int_reg_array_24_13_imag;
  assign io_coef_out_payload_0_24_14_real = int_reg_array_24_14_real;
  assign io_coef_out_payload_0_24_14_imag = int_reg_array_24_14_imag;
  assign io_coef_out_payload_0_24_15_real = int_reg_array_24_15_real;
  assign io_coef_out_payload_0_24_15_imag = int_reg_array_24_15_imag;
  assign io_coef_out_payload_0_24_16_real = int_reg_array_24_16_real;
  assign io_coef_out_payload_0_24_16_imag = int_reg_array_24_16_imag;
  assign io_coef_out_payload_0_24_17_real = int_reg_array_24_17_real;
  assign io_coef_out_payload_0_24_17_imag = int_reg_array_24_17_imag;
  assign io_coef_out_payload_0_24_18_real = int_reg_array_24_18_real;
  assign io_coef_out_payload_0_24_18_imag = int_reg_array_24_18_imag;
  assign io_coef_out_payload_0_24_19_real = int_reg_array_24_19_real;
  assign io_coef_out_payload_0_24_19_imag = int_reg_array_24_19_imag;
  assign io_coef_out_payload_0_24_20_real = int_reg_array_24_20_real;
  assign io_coef_out_payload_0_24_20_imag = int_reg_array_24_20_imag;
  assign io_coef_out_payload_0_24_21_real = int_reg_array_24_21_real;
  assign io_coef_out_payload_0_24_21_imag = int_reg_array_24_21_imag;
  assign io_coef_out_payload_0_24_22_real = int_reg_array_24_22_real;
  assign io_coef_out_payload_0_24_22_imag = int_reg_array_24_22_imag;
  assign io_coef_out_payload_0_24_23_real = int_reg_array_24_23_real;
  assign io_coef_out_payload_0_24_23_imag = int_reg_array_24_23_imag;
  assign io_coef_out_payload_0_24_24_real = int_reg_array_24_24_real;
  assign io_coef_out_payload_0_24_24_imag = int_reg_array_24_24_imag;
  assign io_coef_out_payload_0_24_25_real = int_reg_array_24_25_real;
  assign io_coef_out_payload_0_24_25_imag = int_reg_array_24_25_imag;
  assign io_coef_out_payload_0_24_26_real = int_reg_array_24_26_real;
  assign io_coef_out_payload_0_24_26_imag = int_reg_array_24_26_imag;
  assign io_coef_out_payload_0_24_27_real = int_reg_array_24_27_real;
  assign io_coef_out_payload_0_24_27_imag = int_reg_array_24_27_imag;
  assign io_coef_out_payload_0_24_28_real = int_reg_array_24_28_real;
  assign io_coef_out_payload_0_24_28_imag = int_reg_array_24_28_imag;
  assign io_coef_out_payload_0_24_29_real = int_reg_array_24_29_real;
  assign io_coef_out_payload_0_24_29_imag = int_reg_array_24_29_imag;
  assign io_coef_out_payload_0_24_30_real = int_reg_array_24_30_real;
  assign io_coef_out_payload_0_24_30_imag = int_reg_array_24_30_imag;
  assign io_coef_out_payload_0_24_31_real = int_reg_array_24_31_real;
  assign io_coef_out_payload_0_24_31_imag = int_reg_array_24_31_imag;
  assign io_coef_out_payload_0_24_32_real = int_reg_array_24_32_real;
  assign io_coef_out_payload_0_24_32_imag = int_reg_array_24_32_imag;
  assign io_coef_out_payload_0_24_33_real = int_reg_array_24_33_real;
  assign io_coef_out_payload_0_24_33_imag = int_reg_array_24_33_imag;
  assign io_coef_out_payload_0_24_34_real = int_reg_array_24_34_real;
  assign io_coef_out_payload_0_24_34_imag = int_reg_array_24_34_imag;
  assign io_coef_out_payload_0_24_35_real = int_reg_array_24_35_real;
  assign io_coef_out_payload_0_24_35_imag = int_reg_array_24_35_imag;
  assign io_coef_out_payload_0_24_36_real = int_reg_array_24_36_real;
  assign io_coef_out_payload_0_24_36_imag = int_reg_array_24_36_imag;
  assign io_coef_out_payload_0_24_37_real = int_reg_array_24_37_real;
  assign io_coef_out_payload_0_24_37_imag = int_reg_array_24_37_imag;
  assign io_coef_out_payload_0_24_38_real = int_reg_array_24_38_real;
  assign io_coef_out_payload_0_24_38_imag = int_reg_array_24_38_imag;
  assign io_coef_out_payload_0_24_39_real = int_reg_array_24_39_real;
  assign io_coef_out_payload_0_24_39_imag = int_reg_array_24_39_imag;
  assign io_coef_out_payload_0_24_40_real = int_reg_array_24_40_real;
  assign io_coef_out_payload_0_24_40_imag = int_reg_array_24_40_imag;
  assign io_coef_out_payload_0_24_41_real = int_reg_array_24_41_real;
  assign io_coef_out_payload_0_24_41_imag = int_reg_array_24_41_imag;
  assign io_coef_out_payload_0_24_42_real = int_reg_array_24_42_real;
  assign io_coef_out_payload_0_24_42_imag = int_reg_array_24_42_imag;
  assign io_coef_out_payload_0_24_43_real = int_reg_array_24_43_real;
  assign io_coef_out_payload_0_24_43_imag = int_reg_array_24_43_imag;
  assign io_coef_out_payload_0_24_44_real = int_reg_array_24_44_real;
  assign io_coef_out_payload_0_24_44_imag = int_reg_array_24_44_imag;
  assign io_coef_out_payload_0_24_45_real = int_reg_array_24_45_real;
  assign io_coef_out_payload_0_24_45_imag = int_reg_array_24_45_imag;
  assign io_coef_out_payload_0_24_46_real = int_reg_array_24_46_real;
  assign io_coef_out_payload_0_24_46_imag = int_reg_array_24_46_imag;
  assign io_coef_out_payload_0_24_47_real = int_reg_array_24_47_real;
  assign io_coef_out_payload_0_24_47_imag = int_reg_array_24_47_imag;
  assign io_coef_out_payload_0_24_48_real = int_reg_array_24_48_real;
  assign io_coef_out_payload_0_24_48_imag = int_reg_array_24_48_imag;
  assign io_coef_out_payload_0_24_49_real = int_reg_array_24_49_real;
  assign io_coef_out_payload_0_24_49_imag = int_reg_array_24_49_imag;
  assign io_coef_out_payload_0_25_0_real = int_reg_array_25_0_real;
  assign io_coef_out_payload_0_25_0_imag = int_reg_array_25_0_imag;
  assign io_coef_out_payload_0_25_1_real = int_reg_array_25_1_real;
  assign io_coef_out_payload_0_25_1_imag = int_reg_array_25_1_imag;
  assign io_coef_out_payload_0_25_2_real = int_reg_array_25_2_real;
  assign io_coef_out_payload_0_25_2_imag = int_reg_array_25_2_imag;
  assign io_coef_out_payload_0_25_3_real = int_reg_array_25_3_real;
  assign io_coef_out_payload_0_25_3_imag = int_reg_array_25_3_imag;
  assign io_coef_out_payload_0_25_4_real = int_reg_array_25_4_real;
  assign io_coef_out_payload_0_25_4_imag = int_reg_array_25_4_imag;
  assign io_coef_out_payload_0_25_5_real = int_reg_array_25_5_real;
  assign io_coef_out_payload_0_25_5_imag = int_reg_array_25_5_imag;
  assign io_coef_out_payload_0_25_6_real = int_reg_array_25_6_real;
  assign io_coef_out_payload_0_25_6_imag = int_reg_array_25_6_imag;
  assign io_coef_out_payload_0_25_7_real = int_reg_array_25_7_real;
  assign io_coef_out_payload_0_25_7_imag = int_reg_array_25_7_imag;
  assign io_coef_out_payload_0_25_8_real = int_reg_array_25_8_real;
  assign io_coef_out_payload_0_25_8_imag = int_reg_array_25_8_imag;
  assign io_coef_out_payload_0_25_9_real = int_reg_array_25_9_real;
  assign io_coef_out_payload_0_25_9_imag = int_reg_array_25_9_imag;
  assign io_coef_out_payload_0_25_10_real = int_reg_array_25_10_real;
  assign io_coef_out_payload_0_25_10_imag = int_reg_array_25_10_imag;
  assign io_coef_out_payload_0_25_11_real = int_reg_array_25_11_real;
  assign io_coef_out_payload_0_25_11_imag = int_reg_array_25_11_imag;
  assign io_coef_out_payload_0_25_12_real = int_reg_array_25_12_real;
  assign io_coef_out_payload_0_25_12_imag = int_reg_array_25_12_imag;
  assign io_coef_out_payload_0_25_13_real = int_reg_array_25_13_real;
  assign io_coef_out_payload_0_25_13_imag = int_reg_array_25_13_imag;
  assign io_coef_out_payload_0_25_14_real = int_reg_array_25_14_real;
  assign io_coef_out_payload_0_25_14_imag = int_reg_array_25_14_imag;
  assign io_coef_out_payload_0_25_15_real = int_reg_array_25_15_real;
  assign io_coef_out_payload_0_25_15_imag = int_reg_array_25_15_imag;
  assign io_coef_out_payload_0_25_16_real = int_reg_array_25_16_real;
  assign io_coef_out_payload_0_25_16_imag = int_reg_array_25_16_imag;
  assign io_coef_out_payload_0_25_17_real = int_reg_array_25_17_real;
  assign io_coef_out_payload_0_25_17_imag = int_reg_array_25_17_imag;
  assign io_coef_out_payload_0_25_18_real = int_reg_array_25_18_real;
  assign io_coef_out_payload_0_25_18_imag = int_reg_array_25_18_imag;
  assign io_coef_out_payload_0_25_19_real = int_reg_array_25_19_real;
  assign io_coef_out_payload_0_25_19_imag = int_reg_array_25_19_imag;
  assign io_coef_out_payload_0_25_20_real = int_reg_array_25_20_real;
  assign io_coef_out_payload_0_25_20_imag = int_reg_array_25_20_imag;
  assign io_coef_out_payload_0_25_21_real = int_reg_array_25_21_real;
  assign io_coef_out_payload_0_25_21_imag = int_reg_array_25_21_imag;
  assign io_coef_out_payload_0_25_22_real = int_reg_array_25_22_real;
  assign io_coef_out_payload_0_25_22_imag = int_reg_array_25_22_imag;
  assign io_coef_out_payload_0_25_23_real = int_reg_array_25_23_real;
  assign io_coef_out_payload_0_25_23_imag = int_reg_array_25_23_imag;
  assign io_coef_out_payload_0_25_24_real = int_reg_array_25_24_real;
  assign io_coef_out_payload_0_25_24_imag = int_reg_array_25_24_imag;
  assign io_coef_out_payload_0_25_25_real = int_reg_array_25_25_real;
  assign io_coef_out_payload_0_25_25_imag = int_reg_array_25_25_imag;
  assign io_coef_out_payload_0_25_26_real = int_reg_array_25_26_real;
  assign io_coef_out_payload_0_25_26_imag = int_reg_array_25_26_imag;
  assign io_coef_out_payload_0_25_27_real = int_reg_array_25_27_real;
  assign io_coef_out_payload_0_25_27_imag = int_reg_array_25_27_imag;
  assign io_coef_out_payload_0_25_28_real = int_reg_array_25_28_real;
  assign io_coef_out_payload_0_25_28_imag = int_reg_array_25_28_imag;
  assign io_coef_out_payload_0_25_29_real = int_reg_array_25_29_real;
  assign io_coef_out_payload_0_25_29_imag = int_reg_array_25_29_imag;
  assign io_coef_out_payload_0_25_30_real = int_reg_array_25_30_real;
  assign io_coef_out_payload_0_25_30_imag = int_reg_array_25_30_imag;
  assign io_coef_out_payload_0_25_31_real = int_reg_array_25_31_real;
  assign io_coef_out_payload_0_25_31_imag = int_reg_array_25_31_imag;
  assign io_coef_out_payload_0_25_32_real = int_reg_array_25_32_real;
  assign io_coef_out_payload_0_25_32_imag = int_reg_array_25_32_imag;
  assign io_coef_out_payload_0_25_33_real = int_reg_array_25_33_real;
  assign io_coef_out_payload_0_25_33_imag = int_reg_array_25_33_imag;
  assign io_coef_out_payload_0_25_34_real = int_reg_array_25_34_real;
  assign io_coef_out_payload_0_25_34_imag = int_reg_array_25_34_imag;
  assign io_coef_out_payload_0_25_35_real = int_reg_array_25_35_real;
  assign io_coef_out_payload_0_25_35_imag = int_reg_array_25_35_imag;
  assign io_coef_out_payload_0_25_36_real = int_reg_array_25_36_real;
  assign io_coef_out_payload_0_25_36_imag = int_reg_array_25_36_imag;
  assign io_coef_out_payload_0_25_37_real = int_reg_array_25_37_real;
  assign io_coef_out_payload_0_25_37_imag = int_reg_array_25_37_imag;
  assign io_coef_out_payload_0_25_38_real = int_reg_array_25_38_real;
  assign io_coef_out_payload_0_25_38_imag = int_reg_array_25_38_imag;
  assign io_coef_out_payload_0_25_39_real = int_reg_array_25_39_real;
  assign io_coef_out_payload_0_25_39_imag = int_reg_array_25_39_imag;
  assign io_coef_out_payload_0_25_40_real = int_reg_array_25_40_real;
  assign io_coef_out_payload_0_25_40_imag = int_reg_array_25_40_imag;
  assign io_coef_out_payload_0_25_41_real = int_reg_array_25_41_real;
  assign io_coef_out_payload_0_25_41_imag = int_reg_array_25_41_imag;
  assign io_coef_out_payload_0_25_42_real = int_reg_array_25_42_real;
  assign io_coef_out_payload_0_25_42_imag = int_reg_array_25_42_imag;
  assign io_coef_out_payload_0_25_43_real = int_reg_array_25_43_real;
  assign io_coef_out_payload_0_25_43_imag = int_reg_array_25_43_imag;
  assign io_coef_out_payload_0_25_44_real = int_reg_array_25_44_real;
  assign io_coef_out_payload_0_25_44_imag = int_reg_array_25_44_imag;
  assign io_coef_out_payload_0_25_45_real = int_reg_array_25_45_real;
  assign io_coef_out_payload_0_25_45_imag = int_reg_array_25_45_imag;
  assign io_coef_out_payload_0_25_46_real = int_reg_array_25_46_real;
  assign io_coef_out_payload_0_25_46_imag = int_reg_array_25_46_imag;
  assign io_coef_out_payload_0_25_47_real = int_reg_array_25_47_real;
  assign io_coef_out_payload_0_25_47_imag = int_reg_array_25_47_imag;
  assign io_coef_out_payload_0_25_48_real = int_reg_array_25_48_real;
  assign io_coef_out_payload_0_25_48_imag = int_reg_array_25_48_imag;
  assign io_coef_out_payload_0_25_49_real = int_reg_array_25_49_real;
  assign io_coef_out_payload_0_25_49_imag = int_reg_array_25_49_imag;
  assign io_coef_out_payload_0_26_0_real = int_reg_array_26_0_real;
  assign io_coef_out_payload_0_26_0_imag = int_reg_array_26_0_imag;
  assign io_coef_out_payload_0_26_1_real = int_reg_array_26_1_real;
  assign io_coef_out_payload_0_26_1_imag = int_reg_array_26_1_imag;
  assign io_coef_out_payload_0_26_2_real = int_reg_array_26_2_real;
  assign io_coef_out_payload_0_26_2_imag = int_reg_array_26_2_imag;
  assign io_coef_out_payload_0_26_3_real = int_reg_array_26_3_real;
  assign io_coef_out_payload_0_26_3_imag = int_reg_array_26_3_imag;
  assign io_coef_out_payload_0_26_4_real = int_reg_array_26_4_real;
  assign io_coef_out_payload_0_26_4_imag = int_reg_array_26_4_imag;
  assign io_coef_out_payload_0_26_5_real = int_reg_array_26_5_real;
  assign io_coef_out_payload_0_26_5_imag = int_reg_array_26_5_imag;
  assign io_coef_out_payload_0_26_6_real = int_reg_array_26_6_real;
  assign io_coef_out_payload_0_26_6_imag = int_reg_array_26_6_imag;
  assign io_coef_out_payload_0_26_7_real = int_reg_array_26_7_real;
  assign io_coef_out_payload_0_26_7_imag = int_reg_array_26_7_imag;
  assign io_coef_out_payload_0_26_8_real = int_reg_array_26_8_real;
  assign io_coef_out_payload_0_26_8_imag = int_reg_array_26_8_imag;
  assign io_coef_out_payload_0_26_9_real = int_reg_array_26_9_real;
  assign io_coef_out_payload_0_26_9_imag = int_reg_array_26_9_imag;
  assign io_coef_out_payload_0_26_10_real = int_reg_array_26_10_real;
  assign io_coef_out_payload_0_26_10_imag = int_reg_array_26_10_imag;
  assign io_coef_out_payload_0_26_11_real = int_reg_array_26_11_real;
  assign io_coef_out_payload_0_26_11_imag = int_reg_array_26_11_imag;
  assign io_coef_out_payload_0_26_12_real = int_reg_array_26_12_real;
  assign io_coef_out_payload_0_26_12_imag = int_reg_array_26_12_imag;
  assign io_coef_out_payload_0_26_13_real = int_reg_array_26_13_real;
  assign io_coef_out_payload_0_26_13_imag = int_reg_array_26_13_imag;
  assign io_coef_out_payload_0_26_14_real = int_reg_array_26_14_real;
  assign io_coef_out_payload_0_26_14_imag = int_reg_array_26_14_imag;
  assign io_coef_out_payload_0_26_15_real = int_reg_array_26_15_real;
  assign io_coef_out_payload_0_26_15_imag = int_reg_array_26_15_imag;
  assign io_coef_out_payload_0_26_16_real = int_reg_array_26_16_real;
  assign io_coef_out_payload_0_26_16_imag = int_reg_array_26_16_imag;
  assign io_coef_out_payload_0_26_17_real = int_reg_array_26_17_real;
  assign io_coef_out_payload_0_26_17_imag = int_reg_array_26_17_imag;
  assign io_coef_out_payload_0_26_18_real = int_reg_array_26_18_real;
  assign io_coef_out_payload_0_26_18_imag = int_reg_array_26_18_imag;
  assign io_coef_out_payload_0_26_19_real = int_reg_array_26_19_real;
  assign io_coef_out_payload_0_26_19_imag = int_reg_array_26_19_imag;
  assign io_coef_out_payload_0_26_20_real = int_reg_array_26_20_real;
  assign io_coef_out_payload_0_26_20_imag = int_reg_array_26_20_imag;
  assign io_coef_out_payload_0_26_21_real = int_reg_array_26_21_real;
  assign io_coef_out_payload_0_26_21_imag = int_reg_array_26_21_imag;
  assign io_coef_out_payload_0_26_22_real = int_reg_array_26_22_real;
  assign io_coef_out_payload_0_26_22_imag = int_reg_array_26_22_imag;
  assign io_coef_out_payload_0_26_23_real = int_reg_array_26_23_real;
  assign io_coef_out_payload_0_26_23_imag = int_reg_array_26_23_imag;
  assign io_coef_out_payload_0_26_24_real = int_reg_array_26_24_real;
  assign io_coef_out_payload_0_26_24_imag = int_reg_array_26_24_imag;
  assign io_coef_out_payload_0_26_25_real = int_reg_array_26_25_real;
  assign io_coef_out_payload_0_26_25_imag = int_reg_array_26_25_imag;
  assign io_coef_out_payload_0_26_26_real = int_reg_array_26_26_real;
  assign io_coef_out_payload_0_26_26_imag = int_reg_array_26_26_imag;
  assign io_coef_out_payload_0_26_27_real = int_reg_array_26_27_real;
  assign io_coef_out_payload_0_26_27_imag = int_reg_array_26_27_imag;
  assign io_coef_out_payload_0_26_28_real = int_reg_array_26_28_real;
  assign io_coef_out_payload_0_26_28_imag = int_reg_array_26_28_imag;
  assign io_coef_out_payload_0_26_29_real = int_reg_array_26_29_real;
  assign io_coef_out_payload_0_26_29_imag = int_reg_array_26_29_imag;
  assign io_coef_out_payload_0_26_30_real = int_reg_array_26_30_real;
  assign io_coef_out_payload_0_26_30_imag = int_reg_array_26_30_imag;
  assign io_coef_out_payload_0_26_31_real = int_reg_array_26_31_real;
  assign io_coef_out_payload_0_26_31_imag = int_reg_array_26_31_imag;
  assign io_coef_out_payload_0_26_32_real = int_reg_array_26_32_real;
  assign io_coef_out_payload_0_26_32_imag = int_reg_array_26_32_imag;
  assign io_coef_out_payload_0_26_33_real = int_reg_array_26_33_real;
  assign io_coef_out_payload_0_26_33_imag = int_reg_array_26_33_imag;
  assign io_coef_out_payload_0_26_34_real = int_reg_array_26_34_real;
  assign io_coef_out_payload_0_26_34_imag = int_reg_array_26_34_imag;
  assign io_coef_out_payload_0_26_35_real = int_reg_array_26_35_real;
  assign io_coef_out_payload_0_26_35_imag = int_reg_array_26_35_imag;
  assign io_coef_out_payload_0_26_36_real = int_reg_array_26_36_real;
  assign io_coef_out_payload_0_26_36_imag = int_reg_array_26_36_imag;
  assign io_coef_out_payload_0_26_37_real = int_reg_array_26_37_real;
  assign io_coef_out_payload_0_26_37_imag = int_reg_array_26_37_imag;
  assign io_coef_out_payload_0_26_38_real = int_reg_array_26_38_real;
  assign io_coef_out_payload_0_26_38_imag = int_reg_array_26_38_imag;
  assign io_coef_out_payload_0_26_39_real = int_reg_array_26_39_real;
  assign io_coef_out_payload_0_26_39_imag = int_reg_array_26_39_imag;
  assign io_coef_out_payload_0_26_40_real = int_reg_array_26_40_real;
  assign io_coef_out_payload_0_26_40_imag = int_reg_array_26_40_imag;
  assign io_coef_out_payload_0_26_41_real = int_reg_array_26_41_real;
  assign io_coef_out_payload_0_26_41_imag = int_reg_array_26_41_imag;
  assign io_coef_out_payload_0_26_42_real = int_reg_array_26_42_real;
  assign io_coef_out_payload_0_26_42_imag = int_reg_array_26_42_imag;
  assign io_coef_out_payload_0_26_43_real = int_reg_array_26_43_real;
  assign io_coef_out_payload_0_26_43_imag = int_reg_array_26_43_imag;
  assign io_coef_out_payload_0_26_44_real = int_reg_array_26_44_real;
  assign io_coef_out_payload_0_26_44_imag = int_reg_array_26_44_imag;
  assign io_coef_out_payload_0_26_45_real = int_reg_array_26_45_real;
  assign io_coef_out_payload_0_26_45_imag = int_reg_array_26_45_imag;
  assign io_coef_out_payload_0_26_46_real = int_reg_array_26_46_real;
  assign io_coef_out_payload_0_26_46_imag = int_reg_array_26_46_imag;
  assign io_coef_out_payload_0_26_47_real = int_reg_array_26_47_real;
  assign io_coef_out_payload_0_26_47_imag = int_reg_array_26_47_imag;
  assign io_coef_out_payload_0_26_48_real = int_reg_array_26_48_real;
  assign io_coef_out_payload_0_26_48_imag = int_reg_array_26_48_imag;
  assign io_coef_out_payload_0_26_49_real = int_reg_array_26_49_real;
  assign io_coef_out_payload_0_26_49_imag = int_reg_array_26_49_imag;
  assign io_coef_out_payload_0_27_0_real = int_reg_array_27_0_real;
  assign io_coef_out_payload_0_27_0_imag = int_reg_array_27_0_imag;
  assign io_coef_out_payload_0_27_1_real = int_reg_array_27_1_real;
  assign io_coef_out_payload_0_27_1_imag = int_reg_array_27_1_imag;
  assign io_coef_out_payload_0_27_2_real = int_reg_array_27_2_real;
  assign io_coef_out_payload_0_27_2_imag = int_reg_array_27_2_imag;
  assign io_coef_out_payload_0_27_3_real = int_reg_array_27_3_real;
  assign io_coef_out_payload_0_27_3_imag = int_reg_array_27_3_imag;
  assign io_coef_out_payload_0_27_4_real = int_reg_array_27_4_real;
  assign io_coef_out_payload_0_27_4_imag = int_reg_array_27_4_imag;
  assign io_coef_out_payload_0_27_5_real = int_reg_array_27_5_real;
  assign io_coef_out_payload_0_27_5_imag = int_reg_array_27_5_imag;
  assign io_coef_out_payload_0_27_6_real = int_reg_array_27_6_real;
  assign io_coef_out_payload_0_27_6_imag = int_reg_array_27_6_imag;
  assign io_coef_out_payload_0_27_7_real = int_reg_array_27_7_real;
  assign io_coef_out_payload_0_27_7_imag = int_reg_array_27_7_imag;
  assign io_coef_out_payload_0_27_8_real = int_reg_array_27_8_real;
  assign io_coef_out_payload_0_27_8_imag = int_reg_array_27_8_imag;
  assign io_coef_out_payload_0_27_9_real = int_reg_array_27_9_real;
  assign io_coef_out_payload_0_27_9_imag = int_reg_array_27_9_imag;
  assign io_coef_out_payload_0_27_10_real = int_reg_array_27_10_real;
  assign io_coef_out_payload_0_27_10_imag = int_reg_array_27_10_imag;
  assign io_coef_out_payload_0_27_11_real = int_reg_array_27_11_real;
  assign io_coef_out_payload_0_27_11_imag = int_reg_array_27_11_imag;
  assign io_coef_out_payload_0_27_12_real = int_reg_array_27_12_real;
  assign io_coef_out_payload_0_27_12_imag = int_reg_array_27_12_imag;
  assign io_coef_out_payload_0_27_13_real = int_reg_array_27_13_real;
  assign io_coef_out_payload_0_27_13_imag = int_reg_array_27_13_imag;
  assign io_coef_out_payload_0_27_14_real = int_reg_array_27_14_real;
  assign io_coef_out_payload_0_27_14_imag = int_reg_array_27_14_imag;
  assign io_coef_out_payload_0_27_15_real = int_reg_array_27_15_real;
  assign io_coef_out_payload_0_27_15_imag = int_reg_array_27_15_imag;
  assign io_coef_out_payload_0_27_16_real = int_reg_array_27_16_real;
  assign io_coef_out_payload_0_27_16_imag = int_reg_array_27_16_imag;
  assign io_coef_out_payload_0_27_17_real = int_reg_array_27_17_real;
  assign io_coef_out_payload_0_27_17_imag = int_reg_array_27_17_imag;
  assign io_coef_out_payload_0_27_18_real = int_reg_array_27_18_real;
  assign io_coef_out_payload_0_27_18_imag = int_reg_array_27_18_imag;
  assign io_coef_out_payload_0_27_19_real = int_reg_array_27_19_real;
  assign io_coef_out_payload_0_27_19_imag = int_reg_array_27_19_imag;
  assign io_coef_out_payload_0_27_20_real = int_reg_array_27_20_real;
  assign io_coef_out_payload_0_27_20_imag = int_reg_array_27_20_imag;
  assign io_coef_out_payload_0_27_21_real = int_reg_array_27_21_real;
  assign io_coef_out_payload_0_27_21_imag = int_reg_array_27_21_imag;
  assign io_coef_out_payload_0_27_22_real = int_reg_array_27_22_real;
  assign io_coef_out_payload_0_27_22_imag = int_reg_array_27_22_imag;
  assign io_coef_out_payload_0_27_23_real = int_reg_array_27_23_real;
  assign io_coef_out_payload_0_27_23_imag = int_reg_array_27_23_imag;
  assign io_coef_out_payload_0_27_24_real = int_reg_array_27_24_real;
  assign io_coef_out_payload_0_27_24_imag = int_reg_array_27_24_imag;
  assign io_coef_out_payload_0_27_25_real = int_reg_array_27_25_real;
  assign io_coef_out_payload_0_27_25_imag = int_reg_array_27_25_imag;
  assign io_coef_out_payload_0_27_26_real = int_reg_array_27_26_real;
  assign io_coef_out_payload_0_27_26_imag = int_reg_array_27_26_imag;
  assign io_coef_out_payload_0_27_27_real = int_reg_array_27_27_real;
  assign io_coef_out_payload_0_27_27_imag = int_reg_array_27_27_imag;
  assign io_coef_out_payload_0_27_28_real = int_reg_array_27_28_real;
  assign io_coef_out_payload_0_27_28_imag = int_reg_array_27_28_imag;
  assign io_coef_out_payload_0_27_29_real = int_reg_array_27_29_real;
  assign io_coef_out_payload_0_27_29_imag = int_reg_array_27_29_imag;
  assign io_coef_out_payload_0_27_30_real = int_reg_array_27_30_real;
  assign io_coef_out_payload_0_27_30_imag = int_reg_array_27_30_imag;
  assign io_coef_out_payload_0_27_31_real = int_reg_array_27_31_real;
  assign io_coef_out_payload_0_27_31_imag = int_reg_array_27_31_imag;
  assign io_coef_out_payload_0_27_32_real = int_reg_array_27_32_real;
  assign io_coef_out_payload_0_27_32_imag = int_reg_array_27_32_imag;
  assign io_coef_out_payload_0_27_33_real = int_reg_array_27_33_real;
  assign io_coef_out_payload_0_27_33_imag = int_reg_array_27_33_imag;
  assign io_coef_out_payload_0_27_34_real = int_reg_array_27_34_real;
  assign io_coef_out_payload_0_27_34_imag = int_reg_array_27_34_imag;
  assign io_coef_out_payload_0_27_35_real = int_reg_array_27_35_real;
  assign io_coef_out_payload_0_27_35_imag = int_reg_array_27_35_imag;
  assign io_coef_out_payload_0_27_36_real = int_reg_array_27_36_real;
  assign io_coef_out_payload_0_27_36_imag = int_reg_array_27_36_imag;
  assign io_coef_out_payload_0_27_37_real = int_reg_array_27_37_real;
  assign io_coef_out_payload_0_27_37_imag = int_reg_array_27_37_imag;
  assign io_coef_out_payload_0_27_38_real = int_reg_array_27_38_real;
  assign io_coef_out_payload_0_27_38_imag = int_reg_array_27_38_imag;
  assign io_coef_out_payload_0_27_39_real = int_reg_array_27_39_real;
  assign io_coef_out_payload_0_27_39_imag = int_reg_array_27_39_imag;
  assign io_coef_out_payload_0_27_40_real = int_reg_array_27_40_real;
  assign io_coef_out_payload_0_27_40_imag = int_reg_array_27_40_imag;
  assign io_coef_out_payload_0_27_41_real = int_reg_array_27_41_real;
  assign io_coef_out_payload_0_27_41_imag = int_reg_array_27_41_imag;
  assign io_coef_out_payload_0_27_42_real = int_reg_array_27_42_real;
  assign io_coef_out_payload_0_27_42_imag = int_reg_array_27_42_imag;
  assign io_coef_out_payload_0_27_43_real = int_reg_array_27_43_real;
  assign io_coef_out_payload_0_27_43_imag = int_reg_array_27_43_imag;
  assign io_coef_out_payload_0_27_44_real = int_reg_array_27_44_real;
  assign io_coef_out_payload_0_27_44_imag = int_reg_array_27_44_imag;
  assign io_coef_out_payload_0_27_45_real = int_reg_array_27_45_real;
  assign io_coef_out_payload_0_27_45_imag = int_reg_array_27_45_imag;
  assign io_coef_out_payload_0_27_46_real = int_reg_array_27_46_real;
  assign io_coef_out_payload_0_27_46_imag = int_reg_array_27_46_imag;
  assign io_coef_out_payload_0_27_47_real = int_reg_array_27_47_real;
  assign io_coef_out_payload_0_27_47_imag = int_reg_array_27_47_imag;
  assign io_coef_out_payload_0_27_48_real = int_reg_array_27_48_real;
  assign io_coef_out_payload_0_27_48_imag = int_reg_array_27_48_imag;
  assign io_coef_out_payload_0_27_49_real = int_reg_array_27_49_real;
  assign io_coef_out_payload_0_27_49_imag = int_reg_array_27_49_imag;
  assign io_coef_out_payload_0_28_0_real = int_reg_array_28_0_real;
  assign io_coef_out_payload_0_28_0_imag = int_reg_array_28_0_imag;
  assign io_coef_out_payload_0_28_1_real = int_reg_array_28_1_real;
  assign io_coef_out_payload_0_28_1_imag = int_reg_array_28_1_imag;
  assign io_coef_out_payload_0_28_2_real = int_reg_array_28_2_real;
  assign io_coef_out_payload_0_28_2_imag = int_reg_array_28_2_imag;
  assign io_coef_out_payload_0_28_3_real = int_reg_array_28_3_real;
  assign io_coef_out_payload_0_28_3_imag = int_reg_array_28_3_imag;
  assign io_coef_out_payload_0_28_4_real = int_reg_array_28_4_real;
  assign io_coef_out_payload_0_28_4_imag = int_reg_array_28_4_imag;
  assign io_coef_out_payload_0_28_5_real = int_reg_array_28_5_real;
  assign io_coef_out_payload_0_28_5_imag = int_reg_array_28_5_imag;
  assign io_coef_out_payload_0_28_6_real = int_reg_array_28_6_real;
  assign io_coef_out_payload_0_28_6_imag = int_reg_array_28_6_imag;
  assign io_coef_out_payload_0_28_7_real = int_reg_array_28_7_real;
  assign io_coef_out_payload_0_28_7_imag = int_reg_array_28_7_imag;
  assign io_coef_out_payload_0_28_8_real = int_reg_array_28_8_real;
  assign io_coef_out_payload_0_28_8_imag = int_reg_array_28_8_imag;
  assign io_coef_out_payload_0_28_9_real = int_reg_array_28_9_real;
  assign io_coef_out_payload_0_28_9_imag = int_reg_array_28_9_imag;
  assign io_coef_out_payload_0_28_10_real = int_reg_array_28_10_real;
  assign io_coef_out_payload_0_28_10_imag = int_reg_array_28_10_imag;
  assign io_coef_out_payload_0_28_11_real = int_reg_array_28_11_real;
  assign io_coef_out_payload_0_28_11_imag = int_reg_array_28_11_imag;
  assign io_coef_out_payload_0_28_12_real = int_reg_array_28_12_real;
  assign io_coef_out_payload_0_28_12_imag = int_reg_array_28_12_imag;
  assign io_coef_out_payload_0_28_13_real = int_reg_array_28_13_real;
  assign io_coef_out_payload_0_28_13_imag = int_reg_array_28_13_imag;
  assign io_coef_out_payload_0_28_14_real = int_reg_array_28_14_real;
  assign io_coef_out_payload_0_28_14_imag = int_reg_array_28_14_imag;
  assign io_coef_out_payload_0_28_15_real = int_reg_array_28_15_real;
  assign io_coef_out_payload_0_28_15_imag = int_reg_array_28_15_imag;
  assign io_coef_out_payload_0_28_16_real = int_reg_array_28_16_real;
  assign io_coef_out_payload_0_28_16_imag = int_reg_array_28_16_imag;
  assign io_coef_out_payload_0_28_17_real = int_reg_array_28_17_real;
  assign io_coef_out_payload_0_28_17_imag = int_reg_array_28_17_imag;
  assign io_coef_out_payload_0_28_18_real = int_reg_array_28_18_real;
  assign io_coef_out_payload_0_28_18_imag = int_reg_array_28_18_imag;
  assign io_coef_out_payload_0_28_19_real = int_reg_array_28_19_real;
  assign io_coef_out_payload_0_28_19_imag = int_reg_array_28_19_imag;
  assign io_coef_out_payload_0_28_20_real = int_reg_array_28_20_real;
  assign io_coef_out_payload_0_28_20_imag = int_reg_array_28_20_imag;
  assign io_coef_out_payload_0_28_21_real = int_reg_array_28_21_real;
  assign io_coef_out_payload_0_28_21_imag = int_reg_array_28_21_imag;
  assign io_coef_out_payload_0_28_22_real = int_reg_array_28_22_real;
  assign io_coef_out_payload_0_28_22_imag = int_reg_array_28_22_imag;
  assign io_coef_out_payload_0_28_23_real = int_reg_array_28_23_real;
  assign io_coef_out_payload_0_28_23_imag = int_reg_array_28_23_imag;
  assign io_coef_out_payload_0_28_24_real = int_reg_array_28_24_real;
  assign io_coef_out_payload_0_28_24_imag = int_reg_array_28_24_imag;
  assign io_coef_out_payload_0_28_25_real = int_reg_array_28_25_real;
  assign io_coef_out_payload_0_28_25_imag = int_reg_array_28_25_imag;
  assign io_coef_out_payload_0_28_26_real = int_reg_array_28_26_real;
  assign io_coef_out_payload_0_28_26_imag = int_reg_array_28_26_imag;
  assign io_coef_out_payload_0_28_27_real = int_reg_array_28_27_real;
  assign io_coef_out_payload_0_28_27_imag = int_reg_array_28_27_imag;
  assign io_coef_out_payload_0_28_28_real = int_reg_array_28_28_real;
  assign io_coef_out_payload_0_28_28_imag = int_reg_array_28_28_imag;
  assign io_coef_out_payload_0_28_29_real = int_reg_array_28_29_real;
  assign io_coef_out_payload_0_28_29_imag = int_reg_array_28_29_imag;
  assign io_coef_out_payload_0_28_30_real = int_reg_array_28_30_real;
  assign io_coef_out_payload_0_28_30_imag = int_reg_array_28_30_imag;
  assign io_coef_out_payload_0_28_31_real = int_reg_array_28_31_real;
  assign io_coef_out_payload_0_28_31_imag = int_reg_array_28_31_imag;
  assign io_coef_out_payload_0_28_32_real = int_reg_array_28_32_real;
  assign io_coef_out_payload_0_28_32_imag = int_reg_array_28_32_imag;
  assign io_coef_out_payload_0_28_33_real = int_reg_array_28_33_real;
  assign io_coef_out_payload_0_28_33_imag = int_reg_array_28_33_imag;
  assign io_coef_out_payload_0_28_34_real = int_reg_array_28_34_real;
  assign io_coef_out_payload_0_28_34_imag = int_reg_array_28_34_imag;
  assign io_coef_out_payload_0_28_35_real = int_reg_array_28_35_real;
  assign io_coef_out_payload_0_28_35_imag = int_reg_array_28_35_imag;
  assign io_coef_out_payload_0_28_36_real = int_reg_array_28_36_real;
  assign io_coef_out_payload_0_28_36_imag = int_reg_array_28_36_imag;
  assign io_coef_out_payload_0_28_37_real = int_reg_array_28_37_real;
  assign io_coef_out_payload_0_28_37_imag = int_reg_array_28_37_imag;
  assign io_coef_out_payload_0_28_38_real = int_reg_array_28_38_real;
  assign io_coef_out_payload_0_28_38_imag = int_reg_array_28_38_imag;
  assign io_coef_out_payload_0_28_39_real = int_reg_array_28_39_real;
  assign io_coef_out_payload_0_28_39_imag = int_reg_array_28_39_imag;
  assign io_coef_out_payload_0_28_40_real = int_reg_array_28_40_real;
  assign io_coef_out_payload_0_28_40_imag = int_reg_array_28_40_imag;
  assign io_coef_out_payload_0_28_41_real = int_reg_array_28_41_real;
  assign io_coef_out_payload_0_28_41_imag = int_reg_array_28_41_imag;
  assign io_coef_out_payload_0_28_42_real = int_reg_array_28_42_real;
  assign io_coef_out_payload_0_28_42_imag = int_reg_array_28_42_imag;
  assign io_coef_out_payload_0_28_43_real = int_reg_array_28_43_real;
  assign io_coef_out_payload_0_28_43_imag = int_reg_array_28_43_imag;
  assign io_coef_out_payload_0_28_44_real = int_reg_array_28_44_real;
  assign io_coef_out_payload_0_28_44_imag = int_reg_array_28_44_imag;
  assign io_coef_out_payload_0_28_45_real = int_reg_array_28_45_real;
  assign io_coef_out_payload_0_28_45_imag = int_reg_array_28_45_imag;
  assign io_coef_out_payload_0_28_46_real = int_reg_array_28_46_real;
  assign io_coef_out_payload_0_28_46_imag = int_reg_array_28_46_imag;
  assign io_coef_out_payload_0_28_47_real = int_reg_array_28_47_real;
  assign io_coef_out_payload_0_28_47_imag = int_reg_array_28_47_imag;
  assign io_coef_out_payload_0_28_48_real = int_reg_array_28_48_real;
  assign io_coef_out_payload_0_28_48_imag = int_reg_array_28_48_imag;
  assign io_coef_out_payload_0_28_49_real = int_reg_array_28_49_real;
  assign io_coef_out_payload_0_28_49_imag = int_reg_array_28_49_imag;
  assign io_coef_out_payload_0_29_0_real = int_reg_array_29_0_real;
  assign io_coef_out_payload_0_29_0_imag = int_reg_array_29_0_imag;
  assign io_coef_out_payload_0_29_1_real = int_reg_array_29_1_real;
  assign io_coef_out_payload_0_29_1_imag = int_reg_array_29_1_imag;
  assign io_coef_out_payload_0_29_2_real = int_reg_array_29_2_real;
  assign io_coef_out_payload_0_29_2_imag = int_reg_array_29_2_imag;
  assign io_coef_out_payload_0_29_3_real = int_reg_array_29_3_real;
  assign io_coef_out_payload_0_29_3_imag = int_reg_array_29_3_imag;
  assign io_coef_out_payload_0_29_4_real = int_reg_array_29_4_real;
  assign io_coef_out_payload_0_29_4_imag = int_reg_array_29_4_imag;
  assign io_coef_out_payload_0_29_5_real = int_reg_array_29_5_real;
  assign io_coef_out_payload_0_29_5_imag = int_reg_array_29_5_imag;
  assign io_coef_out_payload_0_29_6_real = int_reg_array_29_6_real;
  assign io_coef_out_payload_0_29_6_imag = int_reg_array_29_6_imag;
  assign io_coef_out_payload_0_29_7_real = int_reg_array_29_7_real;
  assign io_coef_out_payload_0_29_7_imag = int_reg_array_29_7_imag;
  assign io_coef_out_payload_0_29_8_real = int_reg_array_29_8_real;
  assign io_coef_out_payload_0_29_8_imag = int_reg_array_29_8_imag;
  assign io_coef_out_payload_0_29_9_real = int_reg_array_29_9_real;
  assign io_coef_out_payload_0_29_9_imag = int_reg_array_29_9_imag;
  assign io_coef_out_payload_0_29_10_real = int_reg_array_29_10_real;
  assign io_coef_out_payload_0_29_10_imag = int_reg_array_29_10_imag;
  assign io_coef_out_payload_0_29_11_real = int_reg_array_29_11_real;
  assign io_coef_out_payload_0_29_11_imag = int_reg_array_29_11_imag;
  assign io_coef_out_payload_0_29_12_real = int_reg_array_29_12_real;
  assign io_coef_out_payload_0_29_12_imag = int_reg_array_29_12_imag;
  assign io_coef_out_payload_0_29_13_real = int_reg_array_29_13_real;
  assign io_coef_out_payload_0_29_13_imag = int_reg_array_29_13_imag;
  assign io_coef_out_payload_0_29_14_real = int_reg_array_29_14_real;
  assign io_coef_out_payload_0_29_14_imag = int_reg_array_29_14_imag;
  assign io_coef_out_payload_0_29_15_real = int_reg_array_29_15_real;
  assign io_coef_out_payload_0_29_15_imag = int_reg_array_29_15_imag;
  assign io_coef_out_payload_0_29_16_real = int_reg_array_29_16_real;
  assign io_coef_out_payload_0_29_16_imag = int_reg_array_29_16_imag;
  assign io_coef_out_payload_0_29_17_real = int_reg_array_29_17_real;
  assign io_coef_out_payload_0_29_17_imag = int_reg_array_29_17_imag;
  assign io_coef_out_payload_0_29_18_real = int_reg_array_29_18_real;
  assign io_coef_out_payload_0_29_18_imag = int_reg_array_29_18_imag;
  assign io_coef_out_payload_0_29_19_real = int_reg_array_29_19_real;
  assign io_coef_out_payload_0_29_19_imag = int_reg_array_29_19_imag;
  assign io_coef_out_payload_0_29_20_real = int_reg_array_29_20_real;
  assign io_coef_out_payload_0_29_20_imag = int_reg_array_29_20_imag;
  assign io_coef_out_payload_0_29_21_real = int_reg_array_29_21_real;
  assign io_coef_out_payload_0_29_21_imag = int_reg_array_29_21_imag;
  assign io_coef_out_payload_0_29_22_real = int_reg_array_29_22_real;
  assign io_coef_out_payload_0_29_22_imag = int_reg_array_29_22_imag;
  assign io_coef_out_payload_0_29_23_real = int_reg_array_29_23_real;
  assign io_coef_out_payload_0_29_23_imag = int_reg_array_29_23_imag;
  assign io_coef_out_payload_0_29_24_real = int_reg_array_29_24_real;
  assign io_coef_out_payload_0_29_24_imag = int_reg_array_29_24_imag;
  assign io_coef_out_payload_0_29_25_real = int_reg_array_29_25_real;
  assign io_coef_out_payload_0_29_25_imag = int_reg_array_29_25_imag;
  assign io_coef_out_payload_0_29_26_real = int_reg_array_29_26_real;
  assign io_coef_out_payload_0_29_26_imag = int_reg_array_29_26_imag;
  assign io_coef_out_payload_0_29_27_real = int_reg_array_29_27_real;
  assign io_coef_out_payload_0_29_27_imag = int_reg_array_29_27_imag;
  assign io_coef_out_payload_0_29_28_real = int_reg_array_29_28_real;
  assign io_coef_out_payload_0_29_28_imag = int_reg_array_29_28_imag;
  assign io_coef_out_payload_0_29_29_real = int_reg_array_29_29_real;
  assign io_coef_out_payload_0_29_29_imag = int_reg_array_29_29_imag;
  assign io_coef_out_payload_0_29_30_real = int_reg_array_29_30_real;
  assign io_coef_out_payload_0_29_30_imag = int_reg_array_29_30_imag;
  assign io_coef_out_payload_0_29_31_real = int_reg_array_29_31_real;
  assign io_coef_out_payload_0_29_31_imag = int_reg_array_29_31_imag;
  assign io_coef_out_payload_0_29_32_real = int_reg_array_29_32_real;
  assign io_coef_out_payload_0_29_32_imag = int_reg_array_29_32_imag;
  assign io_coef_out_payload_0_29_33_real = int_reg_array_29_33_real;
  assign io_coef_out_payload_0_29_33_imag = int_reg_array_29_33_imag;
  assign io_coef_out_payload_0_29_34_real = int_reg_array_29_34_real;
  assign io_coef_out_payload_0_29_34_imag = int_reg_array_29_34_imag;
  assign io_coef_out_payload_0_29_35_real = int_reg_array_29_35_real;
  assign io_coef_out_payload_0_29_35_imag = int_reg_array_29_35_imag;
  assign io_coef_out_payload_0_29_36_real = int_reg_array_29_36_real;
  assign io_coef_out_payload_0_29_36_imag = int_reg_array_29_36_imag;
  assign io_coef_out_payload_0_29_37_real = int_reg_array_29_37_real;
  assign io_coef_out_payload_0_29_37_imag = int_reg_array_29_37_imag;
  assign io_coef_out_payload_0_29_38_real = int_reg_array_29_38_real;
  assign io_coef_out_payload_0_29_38_imag = int_reg_array_29_38_imag;
  assign io_coef_out_payload_0_29_39_real = int_reg_array_29_39_real;
  assign io_coef_out_payload_0_29_39_imag = int_reg_array_29_39_imag;
  assign io_coef_out_payload_0_29_40_real = int_reg_array_29_40_real;
  assign io_coef_out_payload_0_29_40_imag = int_reg_array_29_40_imag;
  assign io_coef_out_payload_0_29_41_real = int_reg_array_29_41_real;
  assign io_coef_out_payload_0_29_41_imag = int_reg_array_29_41_imag;
  assign io_coef_out_payload_0_29_42_real = int_reg_array_29_42_real;
  assign io_coef_out_payload_0_29_42_imag = int_reg_array_29_42_imag;
  assign io_coef_out_payload_0_29_43_real = int_reg_array_29_43_real;
  assign io_coef_out_payload_0_29_43_imag = int_reg_array_29_43_imag;
  assign io_coef_out_payload_0_29_44_real = int_reg_array_29_44_real;
  assign io_coef_out_payload_0_29_44_imag = int_reg_array_29_44_imag;
  assign io_coef_out_payload_0_29_45_real = int_reg_array_29_45_real;
  assign io_coef_out_payload_0_29_45_imag = int_reg_array_29_45_imag;
  assign io_coef_out_payload_0_29_46_real = int_reg_array_29_46_real;
  assign io_coef_out_payload_0_29_46_imag = int_reg_array_29_46_imag;
  assign io_coef_out_payload_0_29_47_real = int_reg_array_29_47_real;
  assign io_coef_out_payload_0_29_47_imag = int_reg_array_29_47_imag;
  assign io_coef_out_payload_0_29_48_real = int_reg_array_29_48_real;
  assign io_coef_out_payload_0_29_48_imag = int_reg_array_29_48_imag;
  assign io_coef_out_payload_0_29_49_real = int_reg_array_29_49_real;
  assign io_coef_out_payload_0_29_49_imag = int_reg_array_29_49_imag;
  assign io_coef_out_payload_0_30_0_real = int_reg_array_30_0_real;
  assign io_coef_out_payload_0_30_0_imag = int_reg_array_30_0_imag;
  assign io_coef_out_payload_0_30_1_real = int_reg_array_30_1_real;
  assign io_coef_out_payload_0_30_1_imag = int_reg_array_30_1_imag;
  assign io_coef_out_payload_0_30_2_real = int_reg_array_30_2_real;
  assign io_coef_out_payload_0_30_2_imag = int_reg_array_30_2_imag;
  assign io_coef_out_payload_0_30_3_real = int_reg_array_30_3_real;
  assign io_coef_out_payload_0_30_3_imag = int_reg_array_30_3_imag;
  assign io_coef_out_payload_0_30_4_real = int_reg_array_30_4_real;
  assign io_coef_out_payload_0_30_4_imag = int_reg_array_30_4_imag;
  assign io_coef_out_payload_0_30_5_real = int_reg_array_30_5_real;
  assign io_coef_out_payload_0_30_5_imag = int_reg_array_30_5_imag;
  assign io_coef_out_payload_0_30_6_real = int_reg_array_30_6_real;
  assign io_coef_out_payload_0_30_6_imag = int_reg_array_30_6_imag;
  assign io_coef_out_payload_0_30_7_real = int_reg_array_30_7_real;
  assign io_coef_out_payload_0_30_7_imag = int_reg_array_30_7_imag;
  assign io_coef_out_payload_0_30_8_real = int_reg_array_30_8_real;
  assign io_coef_out_payload_0_30_8_imag = int_reg_array_30_8_imag;
  assign io_coef_out_payload_0_30_9_real = int_reg_array_30_9_real;
  assign io_coef_out_payload_0_30_9_imag = int_reg_array_30_9_imag;
  assign io_coef_out_payload_0_30_10_real = int_reg_array_30_10_real;
  assign io_coef_out_payload_0_30_10_imag = int_reg_array_30_10_imag;
  assign io_coef_out_payload_0_30_11_real = int_reg_array_30_11_real;
  assign io_coef_out_payload_0_30_11_imag = int_reg_array_30_11_imag;
  assign io_coef_out_payload_0_30_12_real = int_reg_array_30_12_real;
  assign io_coef_out_payload_0_30_12_imag = int_reg_array_30_12_imag;
  assign io_coef_out_payload_0_30_13_real = int_reg_array_30_13_real;
  assign io_coef_out_payload_0_30_13_imag = int_reg_array_30_13_imag;
  assign io_coef_out_payload_0_30_14_real = int_reg_array_30_14_real;
  assign io_coef_out_payload_0_30_14_imag = int_reg_array_30_14_imag;
  assign io_coef_out_payload_0_30_15_real = int_reg_array_30_15_real;
  assign io_coef_out_payload_0_30_15_imag = int_reg_array_30_15_imag;
  assign io_coef_out_payload_0_30_16_real = int_reg_array_30_16_real;
  assign io_coef_out_payload_0_30_16_imag = int_reg_array_30_16_imag;
  assign io_coef_out_payload_0_30_17_real = int_reg_array_30_17_real;
  assign io_coef_out_payload_0_30_17_imag = int_reg_array_30_17_imag;
  assign io_coef_out_payload_0_30_18_real = int_reg_array_30_18_real;
  assign io_coef_out_payload_0_30_18_imag = int_reg_array_30_18_imag;
  assign io_coef_out_payload_0_30_19_real = int_reg_array_30_19_real;
  assign io_coef_out_payload_0_30_19_imag = int_reg_array_30_19_imag;
  assign io_coef_out_payload_0_30_20_real = int_reg_array_30_20_real;
  assign io_coef_out_payload_0_30_20_imag = int_reg_array_30_20_imag;
  assign io_coef_out_payload_0_30_21_real = int_reg_array_30_21_real;
  assign io_coef_out_payload_0_30_21_imag = int_reg_array_30_21_imag;
  assign io_coef_out_payload_0_30_22_real = int_reg_array_30_22_real;
  assign io_coef_out_payload_0_30_22_imag = int_reg_array_30_22_imag;
  assign io_coef_out_payload_0_30_23_real = int_reg_array_30_23_real;
  assign io_coef_out_payload_0_30_23_imag = int_reg_array_30_23_imag;
  assign io_coef_out_payload_0_30_24_real = int_reg_array_30_24_real;
  assign io_coef_out_payload_0_30_24_imag = int_reg_array_30_24_imag;
  assign io_coef_out_payload_0_30_25_real = int_reg_array_30_25_real;
  assign io_coef_out_payload_0_30_25_imag = int_reg_array_30_25_imag;
  assign io_coef_out_payload_0_30_26_real = int_reg_array_30_26_real;
  assign io_coef_out_payload_0_30_26_imag = int_reg_array_30_26_imag;
  assign io_coef_out_payload_0_30_27_real = int_reg_array_30_27_real;
  assign io_coef_out_payload_0_30_27_imag = int_reg_array_30_27_imag;
  assign io_coef_out_payload_0_30_28_real = int_reg_array_30_28_real;
  assign io_coef_out_payload_0_30_28_imag = int_reg_array_30_28_imag;
  assign io_coef_out_payload_0_30_29_real = int_reg_array_30_29_real;
  assign io_coef_out_payload_0_30_29_imag = int_reg_array_30_29_imag;
  assign io_coef_out_payload_0_30_30_real = int_reg_array_30_30_real;
  assign io_coef_out_payload_0_30_30_imag = int_reg_array_30_30_imag;
  assign io_coef_out_payload_0_30_31_real = int_reg_array_30_31_real;
  assign io_coef_out_payload_0_30_31_imag = int_reg_array_30_31_imag;
  assign io_coef_out_payload_0_30_32_real = int_reg_array_30_32_real;
  assign io_coef_out_payload_0_30_32_imag = int_reg_array_30_32_imag;
  assign io_coef_out_payload_0_30_33_real = int_reg_array_30_33_real;
  assign io_coef_out_payload_0_30_33_imag = int_reg_array_30_33_imag;
  assign io_coef_out_payload_0_30_34_real = int_reg_array_30_34_real;
  assign io_coef_out_payload_0_30_34_imag = int_reg_array_30_34_imag;
  assign io_coef_out_payload_0_30_35_real = int_reg_array_30_35_real;
  assign io_coef_out_payload_0_30_35_imag = int_reg_array_30_35_imag;
  assign io_coef_out_payload_0_30_36_real = int_reg_array_30_36_real;
  assign io_coef_out_payload_0_30_36_imag = int_reg_array_30_36_imag;
  assign io_coef_out_payload_0_30_37_real = int_reg_array_30_37_real;
  assign io_coef_out_payload_0_30_37_imag = int_reg_array_30_37_imag;
  assign io_coef_out_payload_0_30_38_real = int_reg_array_30_38_real;
  assign io_coef_out_payload_0_30_38_imag = int_reg_array_30_38_imag;
  assign io_coef_out_payload_0_30_39_real = int_reg_array_30_39_real;
  assign io_coef_out_payload_0_30_39_imag = int_reg_array_30_39_imag;
  assign io_coef_out_payload_0_30_40_real = int_reg_array_30_40_real;
  assign io_coef_out_payload_0_30_40_imag = int_reg_array_30_40_imag;
  assign io_coef_out_payload_0_30_41_real = int_reg_array_30_41_real;
  assign io_coef_out_payload_0_30_41_imag = int_reg_array_30_41_imag;
  assign io_coef_out_payload_0_30_42_real = int_reg_array_30_42_real;
  assign io_coef_out_payload_0_30_42_imag = int_reg_array_30_42_imag;
  assign io_coef_out_payload_0_30_43_real = int_reg_array_30_43_real;
  assign io_coef_out_payload_0_30_43_imag = int_reg_array_30_43_imag;
  assign io_coef_out_payload_0_30_44_real = int_reg_array_30_44_real;
  assign io_coef_out_payload_0_30_44_imag = int_reg_array_30_44_imag;
  assign io_coef_out_payload_0_30_45_real = int_reg_array_30_45_real;
  assign io_coef_out_payload_0_30_45_imag = int_reg_array_30_45_imag;
  assign io_coef_out_payload_0_30_46_real = int_reg_array_30_46_real;
  assign io_coef_out_payload_0_30_46_imag = int_reg_array_30_46_imag;
  assign io_coef_out_payload_0_30_47_real = int_reg_array_30_47_real;
  assign io_coef_out_payload_0_30_47_imag = int_reg_array_30_47_imag;
  assign io_coef_out_payload_0_30_48_real = int_reg_array_30_48_real;
  assign io_coef_out_payload_0_30_48_imag = int_reg_array_30_48_imag;
  assign io_coef_out_payload_0_30_49_real = int_reg_array_30_49_real;
  assign io_coef_out_payload_0_30_49_imag = int_reg_array_30_49_imag;
  assign io_coef_out_payload_0_31_0_real = int_reg_array_31_0_real;
  assign io_coef_out_payload_0_31_0_imag = int_reg_array_31_0_imag;
  assign io_coef_out_payload_0_31_1_real = int_reg_array_31_1_real;
  assign io_coef_out_payload_0_31_1_imag = int_reg_array_31_1_imag;
  assign io_coef_out_payload_0_31_2_real = int_reg_array_31_2_real;
  assign io_coef_out_payload_0_31_2_imag = int_reg_array_31_2_imag;
  assign io_coef_out_payload_0_31_3_real = int_reg_array_31_3_real;
  assign io_coef_out_payload_0_31_3_imag = int_reg_array_31_3_imag;
  assign io_coef_out_payload_0_31_4_real = int_reg_array_31_4_real;
  assign io_coef_out_payload_0_31_4_imag = int_reg_array_31_4_imag;
  assign io_coef_out_payload_0_31_5_real = int_reg_array_31_5_real;
  assign io_coef_out_payload_0_31_5_imag = int_reg_array_31_5_imag;
  assign io_coef_out_payload_0_31_6_real = int_reg_array_31_6_real;
  assign io_coef_out_payload_0_31_6_imag = int_reg_array_31_6_imag;
  assign io_coef_out_payload_0_31_7_real = int_reg_array_31_7_real;
  assign io_coef_out_payload_0_31_7_imag = int_reg_array_31_7_imag;
  assign io_coef_out_payload_0_31_8_real = int_reg_array_31_8_real;
  assign io_coef_out_payload_0_31_8_imag = int_reg_array_31_8_imag;
  assign io_coef_out_payload_0_31_9_real = int_reg_array_31_9_real;
  assign io_coef_out_payload_0_31_9_imag = int_reg_array_31_9_imag;
  assign io_coef_out_payload_0_31_10_real = int_reg_array_31_10_real;
  assign io_coef_out_payload_0_31_10_imag = int_reg_array_31_10_imag;
  assign io_coef_out_payload_0_31_11_real = int_reg_array_31_11_real;
  assign io_coef_out_payload_0_31_11_imag = int_reg_array_31_11_imag;
  assign io_coef_out_payload_0_31_12_real = int_reg_array_31_12_real;
  assign io_coef_out_payload_0_31_12_imag = int_reg_array_31_12_imag;
  assign io_coef_out_payload_0_31_13_real = int_reg_array_31_13_real;
  assign io_coef_out_payload_0_31_13_imag = int_reg_array_31_13_imag;
  assign io_coef_out_payload_0_31_14_real = int_reg_array_31_14_real;
  assign io_coef_out_payload_0_31_14_imag = int_reg_array_31_14_imag;
  assign io_coef_out_payload_0_31_15_real = int_reg_array_31_15_real;
  assign io_coef_out_payload_0_31_15_imag = int_reg_array_31_15_imag;
  assign io_coef_out_payload_0_31_16_real = int_reg_array_31_16_real;
  assign io_coef_out_payload_0_31_16_imag = int_reg_array_31_16_imag;
  assign io_coef_out_payload_0_31_17_real = int_reg_array_31_17_real;
  assign io_coef_out_payload_0_31_17_imag = int_reg_array_31_17_imag;
  assign io_coef_out_payload_0_31_18_real = int_reg_array_31_18_real;
  assign io_coef_out_payload_0_31_18_imag = int_reg_array_31_18_imag;
  assign io_coef_out_payload_0_31_19_real = int_reg_array_31_19_real;
  assign io_coef_out_payload_0_31_19_imag = int_reg_array_31_19_imag;
  assign io_coef_out_payload_0_31_20_real = int_reg_array_31_20_real;
  assign io_coef_out_payload_0_31_20_imag = int_reg_array_31_20_imag;
  assign io_coef_out_payload_0_31_21_real = int_reg_array_31_21_real;
  assign io_coef_out_payload_0_31_21_imag = int_reg_array_31_21_imag;
  assign io_coef_out_payload_0_31_22_real = int_reg_array_31_22_real;
  assign io_coef_out_payload_0_31_22_imag = int_reg_array_31_22_imag;
  assign io_coef_out_payload_0_31_23_real = int_reg_array_31_23_real;
  assign io_coef_out_payload_0_31_23_imag = int_reg_array_31_23_imag;
  assign io_coef_out_payload_0_31_24_real = int_reg_array_31_24_real;
  assign io_coef_out_payload_0_31_24_imag = int_reg_array_31_24_imag;
  assign io_coef_out_payload_0_31_25_real = int_reg_array_31_25_real;
  assign io_coef_out_payload_0_31_25_imag = int_reg_array_31_25_imag;
  assign io_coef_out_payload_0_31_26_real = int_reg_array_31_26_real;
  assign io_coef_out_payload_0_31_26_imag = int_reg_array_31_26_imag;
  assign io_coef_out_payload_0_31_27_real = int_reg_array_31_27_real;
  assign io_coef_out_payload_0_31_27_imag = int_reg_array_31_27_imag;
  assign io_coef_out_payload_0_31_28_real = int_reg_array_31_28_real;
  assign io_coef_out_payload_0_31_28_imag = int_reg_array_31_28_imag;
  assign io_coef_out_payload_0_31_29_real = int_reg_array_31_29_real;
  assign io_coef_out_payload_0_31_29_imag = int_reg_array_31_29_imag;
  assign io_coef_out_payload_0_31_30_real = int_reg_array_31_30_real;
  assign io_coef_out_payload_0_31_30_imag = int_reg_array_31_30_imag;
  assign io_coef_out_payload_0_31_31_real = int_reg_array_31_31_real;
  assign io_coef_out_payload_0_31_31_imag = int_reg_array_31_31_imag;
  assign io_coef_out_payload_0_31_32_real = int_reg_array_31_32_real;
  assign io_coef_out_payload_0_31_32_imag = int_reg_array_31_32_imag;
  assign io_coef_out_payload_0_31_33_real = int_reg_array_31_33_real;
  assign io_coef_out_payload_0_31_33_imag = int_reg_array_31_33_imag;
  assign io_coef_out_payload_0_31_34_real = int_reg_array_31_34_real;
  assign io_coef_out_payload_0_31_34_imag = int_reg_array_31_34_imag;
  assign io_coef_out_payload_0_31_35_real = int_reg_array_31_35_real;
  assign io_coef_out_payload_0_31_35_imag = int_reg_array_31_35_imag;
  assign io_coef_out_payload_0_31_36_real = int_reg_array_31_36_real;
  assign io_coef_out_payload_0_31_36_imag = int_reg_array_31_36_imag;
  assign io_coef_out_payload_0_31_37_real = int_reg_array_31_37_real;
  assign io_coef_out_payload_0_31_37_imag = int_reg_array_31_37_imag;
  assign io_coef_out_payload_0_31_38_real = int_reg_array_31_38_real;
  assign io_coef_out_payload_0_31_38_imag = int_reg_array_31_38_imag;
  assign io_coef_out_payload_0_31_39_real = int_reg_array_31_39_real;
  assign io_coef_out_payload_0_31_39_imag = int_reg_array_31_39_imag;
  assign io_coef_out_payload_0_31_40_real = int_reg_array_31_40_real;
  assign io_coef_out_payload_0_31_40_imag = int_reg_array_31_40_imag;
  assign io_coef_out_payload_0_31_41_real = int_reg_array_31_41_real;
  assign io_coef_out_payload_0_31_41_imag = int_reg_array_31_41_imag;
  assign io_coef_out_payload_0_31_42_real = int_reg_array_31_42_real;
  assign io_coef_out_payload_0_31_42_imag = int_reg_array_31_42_imag;
  assign io_coef_out_payload_0_31_43_real = int_reg_array_31_43_real;
  assign io_coef_out_payload_0_31_43_imag = int_reg_array_31_43_imag;
  assign io_coef_out_payload_0_31_44_real = int_reg_array_31_44_real;
  assign io_coef_out_payload_0_31_44_imag = int_reg_array_31_44_imag;
  assign io_coef_out_payload_0_31_45_real = int_reg_array_31_45_real;
  assign io_coef_out_payload_0_31_45_imag = int_reg_array_31_45_imag;
  assign io_coef_out_payload_0_31_46_real = int_reg_array_31_46_real;
  assign io_coef_out_payload_0_31_46_imag = int_reg_array_31_46_imag;
  assign io_coef_out_payload_0_31_47_real = int_reg_array_31_47_real;
  assign io_coef_out_payload_0_31_47_imag = int_reg_array_31_47_imag;
  assign io_coef_out_payload_0_31_48_real = int_reg_array_31_48_real;
  assign io_coef_out_payload_0_31_48_imag = int_reg_array_31_48_imag;
  assign io_coef_out_payload_0_31_49_real = int_reg_array_31_49_real;
  assign io_coef_out_payload_0_31_49_imag = int_reg_array_31_49_imag;
  assign io_coef_out_payload_0_32_0_real = int_reg_array_32_0_real;
  assign io_coef_out_payload_0_32_0_imag = int_reg_array_32_0_imag;
  assign io_coef_out_payload_0_32_1_real = int_reg_array_32_1_real;
  assign io_coef_out_payload_0_32_1_imag = int_reg_array_32_1_imag;
  assign io_coef_out_payload_0_32_2_real = int_reg_array_32_2_real;
  assign io_coef_out_payload_0_32_2_imag = int_reg_array_32_2_imag;
  assign io_coef_out_payload_0_32_3_real = int_reg_array_32_3_real;
  assign io_coef_out_payload_0_32_3_imag = int_reg_array_32_3_imag;
  assign io_coef_out_payload_0_32_4_real = int_reg_array_32_4_real;
  assign io_coef_out_payload_0_32_4_imag = int_reg_array_32_4_imag;
  assign io_coef_out_payload_0_32_5_real = int_reg_array_32_5_real;
  assign io_coef_out_payload_0_32_5_imag = int_reg_array_32_5_imag;
  assign io_coef_out_payload_0_32_6_real = int_reg_array_32_6_real;
  assign io_coef_out_payload_0_32_6_imag = int_reg_array_32_6_imag;
  assign io_coef_out_payload_0_32_7_real = int_reg_array_32_7_real;
  assign io_coef_out_payload_0_32_7_imag = int_reg_array_32_7_imag;
  assign io_coef_out_payload_0_32_8_real = int_reg_array_32_8_real;
  assign io_coef_out_payload_0_32_8_imag = int_reg_array_32_8_imag;
  assign io_coef_out_payload_0_32_9_real = int_reg_array_32_9_real;
  assign io_coef_out_payload_0_32_9_imag = int_reg_array_32_9_imag;
  assign io_coef_out_payload_0_32_10_real = int_reg_array_32_10_real;
  assign io_coef_out_payload_0_32_10_imag = int_reg_array_32_10_imag;
  assign io_coef_out_payload_0_32_11_real = int_reg_array_32_11_real;
  assign io_coef_out_payload_0_32_11_imag = int_reg_array_32_11_imag;
  assign io_coef_out_payload_0_32_12_real = int_reg_array_32_12_real;
  assign io_coef_out_payload_0_32_12_imag = int_reg_array_32_12_imag;
  assign io_coef_out_payload_0_32_13_real = int_reg_array_32_13_real;
  assign io_coef_out_payload_0_32_13_imag = int_reg_array_32_13_imag;
  assign io_coef_out_payload_0_32_14_real = int_reg_array_32_14_real;
  assign io_coef_out_payload_0_32_14_imag = int_reg_array_32_14_imag;
  assign io_coef_out_payload_0_32_15_real = int_reg_array_32_15_real;
  assign io_coef_out_payload_0_32_15_imag = int_reg_array_32_15_imag;
  assign io_coef_out_payload_0_32_16_real = int_reg_array_32_16_real;
  assign io_coef_out_payload_0_32_16_imag = int_reg_array_32_16_imag;
  assign io_coef_out_payload_0_32_17_real = int_reg_array_32_17_real;
  assign io_coef_out_payload_0_32_17_imag = int_reg_array_32_17_imag;
  assign io_coef_out_payload_0_32_18_real = int_reg_array_32_18_real;
  assign io_coef_out_payload_0_32_18_imag = int_reg_array_32_18_imag;
  assign io_coef_out_payload_0_32_19_real = int_reg_array_32_19_real;
  assign io_coef_out_payload_0_32_19_imag = int_reg_array_32_19_imag;
  assign io_coef_out_payload_0_32_20_real = int_reg_array_32_20_real;
  assign io_coef_out_payload_0_32_20_imag = int_reg_array_32_20_imag;
  assign io_coef_out_payload_0_32_21_real = int_reg_array_32_21_real;
  assign io_coef_out_payload_0_32_21_imag = int_reg_array_32_21_imag;
  assign io_coef_out_payload_0_32_22_real = int_reg_array_32_22_real;
  assign io_coef_out_payload_0_32_22_imag = int_reg_array_32_22_imag;
  assign io_coef_out_payload_0_32_23_real = int_reg_array_32_23_real;
  assign io_coef_out_payload_0_32_23_imag = int_reg_array_32_23_imag;
  assign io_coef_out_payload_0_32_24_real = int_reg_array_32_24_real;
  assign io_coef_out_payload_0_32_24_imag = int_reg_array_32_24_imag;
  assign io_coef_out_payload_0_32_25_real = int_reg_array_32_25_real;
  assign io_coef_out_payload_0_32_25_imag = int_reg_array_32_25_imag;
  assign io_coef_out_payload_0_32_26_real = int_reg_array_32_26_real;
  assign io_coef_out_payload_0_32_26_imag = int_reg_array_32_26_imag;
  assign io_coef_out_payload_0_32_27_real = int_reg_array_32_27_real;
  assign io_coef_out_payload_0_32_27_imag = int_reg_array_32_27_imag;
  assign io_coef_out_payload_0_32_28_real = int_reg_array_32_28_real;
  assign io_coef_out_payload_0_32_28_imag = int_reg_array_32_28_imag;
  assign io_coef_out_payload_0_32_29_real = int_reg_array_32_29_real;
  assign io_coef_out_payload_0_32_29_imag = int_reg_array_32_29_imag;
  assign io_coef_out_payload_0_32_30_real = int_reg_array_32_30_real;
  assign io_coef_out_payload_0_32_30_imag = int_reg_array_32_30_imag;
  assign io_coef_out_payload_0_32_31_real = int_reg_array_32_31_real;
  assign io_coef_out_payload_0_32_31_imag = int_reg_array_32_31_imag;
  assign io_coef_out_payload_0_32_32_real = int_reg_array_32_32_real;
  assign io_coef_out_payload_0_32_32_imag = int_reg_array_32_32_imag;
  assign io_coef_out_payload_0_32_33_real = int_reg_array_32_33_real;
  assign io_coef_out_payload_0_32_33_imag = int_reg_array_32_33_imag;
  assign io_coef_out_payload_0_32_34_real = int_reg_array_32_34_real;
  assign io_coef_out_payload_0_32_34_imag = int_reg_array_32_34_imag;
  assign io_coef_out_payload_0_32_35_real = int_reg_array_32_35_real;
  assign io_coef_out_payload_0_32_35_imag = int_reg_array_32_35_imag;
  assign io_coef_out_payload_0_32_36_real = int_reg_array_32_36_real;
  assign io_coef_out_payload_0_32_36_imag = int_reg_array_32_36_imag;
  assign io_coef_out_payload_0_32_37_real = int_reg_array_32_37_real;
  assign io_coef_out_payload_0_32_37_imag = int_reg_array_32_37_imag;
  assign io_coef_out_payload_0_32_38_real = int_reg_array_32_38_real;
  assign io_coef_out_payload_0_32_38_imag = int_reg_array_32_38_imag;
  assign io_coef_out_payload_0_32_39_real = int_reg_array_32_39_real;
  assign io_coef_out_payload_0_32_39_imag = int_reg_array_32_39_imag;
  assign io_coef_out_payload_0_32_40_real = int_reg_array_32_40_real;
  assign io_coef_out_payload_0_32_40_imag = int_reg_array_32_40_imag;
  assign io_coef_out_payload_0_32_41_real = int_reg_array_32_41_real;
  assign io_coef_out_payload_0_32_41_imag = int_reg_array_32_41_imag;
  assign io_coef_out_payload_0_32_42_real = int_reg_array_32_42_real;
  assign io_coef_out_payload_0_32_42_imag = int_reg_array_32_42_imag;
  assign io_coef_out_payload_0_32_43_real = int_reg_array_32_43_real;
  assign io_coef_out_payload_0_32_43_imag = int_reg_array_32_43_imag;
  assign io_coef_out_payload_0_32_44_real = int_reg_array_32_44_real;
  assign io_coef_out_payload_0_32_44_imag = int_reg_array_32_44_imag;
  assign io_coef_out_payload_0_32_45_real = int_reg_array_32_45_real;
  assign io_coef_out_payload_0_32_45_imag = int_reg_array_32_45_imag;
  assign io_coef_out_payload_0_32_46_real = int_reg_array_32_46_real;
  assign io_coef_out_payload_0_32_46_imag = int_reg_array_32_46_imag;
  assign io_coef_out_payload_0_32_47_real = int_reg_array_32_47_real;
  assign io_coef_out_payload_0_32_47_imag = int_reg_array_32_47_imag;
  assign io_coef_out_payload_0_32_48_real = int_reg_array_32_48_real;
  assign io_coef_out_payload_0_32_48_imag = int_reg_array_32_48_imag;
  assign io_coef_out_payload_0_32_49_real = int_reg_array_32_49_real;
  assign io_coef_out_payload_0_32_49_imag = int_reg_array_32_49_imag;
  assign io_coef_out_payload_0_33_0_real = int_reg_array_33_0_real;
  assign io_coef_out_payload_0_33_0_imag = int_reg_array_33_0_imag;
  assign io_coef_out_payload_0_33_1_real = int_reg_array_33_1_real;
  assign io_coef_out_payload_0_33_1_imag = int_reg_array_33_1_imag;
  assign io_coef_out_payload_0_33_2_real = int_reg_array_33_2_real;
  assign io_coef_out_payload_0_33_2_imag = int_reg_array_33_2_imag;
  assign io_coef_out_payload_0_33_3_real = int_reg_array_33_3_real;
  assign io_coef_out_payload_0_33_3_imag = int_reg_array_33_3_imag;
  assign io_coef_out_payload_0_33_4_real = int_reg_array_33_4_real;
  assign io_coef_out_payload_0_33_4_imag = int_reg_array_33_4_imag;
  assign io_coef_out_payload_0_33_5_real = int_reg_array_33_5_real;
  assign io_coef_out_payload_0_33_5_imag = int_reg_array_33_5_imag;
  assign io_coef_out_payload_0_33_6_real = int_reg_array_33_6_real;
  assign io_coef_out_payload_0_33_6_imag = int_reg_array_33_6_imag;
  assign io_coef_out_payload_0_33_7_real = int_reg_array_33_7_real;
  assign io_coef_out_payload_0_33_7_imag = int_reg_array_33_7_imag;
  assign io_coef_out_payload_0_33_8_real = int_reg_array_33_8_real;
  assign io_coef_out_payload_0_33_8_imag = int_reg_array_33_8_imag;
  assign io_coef_out_payload_0_33_9_real = int_reg_array_33_9_real;
  assign io_coef_out_payload_0_33_9_imag = int_reg_array_33_9_imag;
  assign io_coef_out_payload_0_33_10_real = int_reg_array_33_10_real;
  assign io_coef_out_payload_0_33_10_imag = int_reg_array_33_10_imag;
  assign io_coef_out_payload_0_33_11_real = int_reg_array_33_11_real;
  assign io_coef_out_payload_0_33_11_imag = int_reg_array_33_11_imag;
  assign io_coef_out_payload_0_33_12_real = int_reg_array_33_12_real;
  assign io_coef_out_payload_0_33_12_imag = int_reg_array_33_12_imag;
  assign io_coef_out_payload_0_33_13_real = int_reg_array_33_13_real;
  assign io_coef_out_payload_0_33_13_imag = int_reg_array_33_13_imag;
  assign io_coef_out_payload_0_33_14_real = int_reg_array_33_14_real;
  assign io_coef_out_payload_0_33_14_imag = int_reg_array_33_14_imag;
  assign io_coef_out_payload_0_33_15_real = int_reg_array_33_15_real;
  assign io_coef_out_payload_0_33_15_imag = int_reg_array_33_15_imag;
  assign io_coef_out_payload_0_33_16_real = int_reg_array_33_16_real;
  assign io_coef_out_payload_0_33_16_imag = int_reg_array_33_16_imag;
  assign io_coef_out_payload_0_33_17_real = int_reg_array_33_17_real;
  assign io_coef_out_payload_0_33_17_imag = int_reg_array_33_17_imag;
  assign io_coef_out_payload_0_33_18_real = int_reg_array_33_18_real;
  assign io_coef_out_payload_0_33_18_imag = int_reg_array_33_18_imag;
  assign io_coef_out_payload_0_33_19_real = int_reg_array_33_19_real;
  assign io_coef_out_payload_0_33_19_imag = int_reg_array_33_19_imag;
  assign io_coef_out_payload_0_33_20_real = int_reg_array_33_20_real;
  assign io_coef_out_payload_0_33_20_imag = int_reg_array_33_20_imag;
  assign io_coef_out_payload_0_33_21_real = int_reg_array_33_21_real;
  assign io_coef_out_payload_0_33_21_imag = int_reg_array_33_21_imag;
  assign io_coef_out_payload_0_33_22_real = int_reg_array_33_22_real;
  assign io_coef_out_payload_0_33_22_imag = int_reg_array_33_22_imag;
  assign io_coef_out_payload_0_33_23_real = int_reg_array_33_23_real;
  assign io_coef_out_payload_0_33_23_imag = int_reg_array_33_23_imag;
  assign io_coef_out_payload_0_33_24_real = int_reg_array_33_24_real;
  assign io_coef_out_payload_0_33_24_imag = int_reg_array_33_24_imag;
  assign io_coef_out_payload_0_33_25_real = int_reg_array_33_25_real;
  assign io_coef_out_payload_0_33_25_imag = int_reg_array_33_25_imag;
  assign io_coef_out_payload_0_33_26_real = int_reg_array_33_26_real;
  assign io_coef_out_payload_0_33_26_imag = int_reg_array_33_26_imag;
  assign io_coef_out_payload_0_33_27_real = int_reg_array_33_27_real;
  assign io_coef_out_payload_0_33_27_imag = int_reg_array_33_27_imag;
  assign io_coef_out_payload_0_33_28_real = int_reg_array_33_28_real;
  assign io_coef_out_payload_0_33_28_imag = int_reg_array_33_28_imag;
  assign io_coef_out_payload_0_33_29_real = int_reg_array_33_29_real;
  assign io_coef_out_payload_0_33_29_imag = int_reg_array_33_29_imag;
  assign io_coef_out_payload_0_33_30_real = int_reg_array_33_30_real;
  assign io_coef_out_payload_0_33_30_imag = int_reg_array_33_30_imag;
  assign io_coef_out_payload_0_33_31_real = int_reg_array_33_31_real;
  assign io_coef_out_payload_0_33_31_imag = int_reg_array_33_31_imag;
  assign io_coef_out_payload_0_33_32_real = int_reg_array_33_32_real;
  assign io_coef_out_payload_0_33_32_imag = int_reg_array_33_32_imag;
  assign io_coef_out_payload_0_33_33_real = int_reg_array_33_33_real;
  assign io_coef_out_payload_0_33_33_imag = int_reg_array_33_33_imag;
  assign io_coef_out_payload_0_33_34_real = int_reg_array_33_34_real;
  assign io_coef_out_payload_0_33_34_imag = int_reg_array_33_34_imag;
  assign io_coef_out_payload_0_33_35_real = int_reg_array_33_35_real;
  assign io_coef_out_payload_0_33_35_imag = int_reg_array_33_35_imag;
  assign io_coef_out_payload_0_33_36_real = int_reg_array_33_36_real;
  assign io_coef_out_payload_0_33_36_imag = int_reg_array_33_36_imag;
  assign io_coef_out_payload_0_33_37_real = int_reg_array_33_37_real;
  assign io_coef_out_payload_0_33_37_imag = int_reg_array_33_37_imag;
  assign io_coef_out_payload_0_33_38_real = int_reg_array_33_38_real;
  assign io_coef_out_payload_0_33_38_imag = int_reg_array_33_38_imag;
  assign io_coef_out_payload_0_33_39_real = int_reg_array_33_39_real;
  assign io_coef_out_payload_0_33_39_imag = int_reg_array_33_39_imag;
  assign io_coef_out_payload_0_33_40_real = int_reg_array_33_40_real;
  assign io_coef_out_payload_0_33_40_imag = int_reg_array_33_40_imag;
  assign io_coef_out_payload_0_33_41_real = int_reg_array_33_41_real;
  assign io_coef_out_payload_0_33_41_imag = int_reg_array_33_41_imag;
  assign io_coef_out_payload_0_33_42_real = int_reg_array_33_42_real;
  assign io_coef_out_payload_0_33_42_imag = int_reg_array_33_42_imag;
  assign io_coef_out_payload_0_33_43_real = int_reg_array_33_43_real;
  assign io_coef_out_payload_0_33_43_imag = int_reg_array_33_43_imag;
  assign io_coef_out_payload_0_33_44_real = int_reg_array_33_44_real;
  assign io_coef_out_payload_0_33_44_imag = int_reg_array_33_44_imag;
  assign io_coef_out_payload_0_33_45_real = int_reg_array_33_45_real;
  assign io_coef_out_payload_0_33_45_imag = int_reg_array_33_45_imag;
  assign io_coef_out_payload_0_33_46_real = int_reg_array_33_46_real;
  assign io_coef_out_payload_0_33_46_imag = int_reg_array_33_46_imag;
  assign io_coef_out_payload_0_33_47_real = int_reg_array_33_47_real;
  assign io_coef_out_payload_0_33_47_imag = int_reg_array_33_47_imag;
  assign io_coef_out_payload_0_33_48_real = int_reg_array_33_48_real;
  assign io_coef_out_payload_0_33_48_imag = int_reg_array_33_48_imag;
  assign io_coef_out_payload_0_33_49_real = int_reg_array_33_49_real;
  assign io_coef_out_payload_0_33_49_imag = int_reg_array_33_49_imag;
  assign io_coef_out_payload_0_34_0_real = int_reg_array_34_0_real;
  assign io_coef_out_payload_0_34_0_imag = int_reg_array_34_0_imag;
  assign io_coef_out_payload_0_34_1_real = int_reg_array_34_1_real;
  assign io_coef_out_payload_0_34_1_imag = int_reg_array_34_1_imag;
  assign io_coef_out_payload_0_34_2_real = int_reg_array_34_2_real;
  assign io_coef_out_payload_0_34_2_imag = int_reg_array_34_2_imag;
  assign io_coef_out_payload_0_34_3_real = int_reg_array_34_3_real;
  assign io_coef_out_payload_0_34_3_imag = int_reg_array_34_3_imag;
  assign io_coef_out_payload_0_34_4_real = int_reg_array_34_4_real;
  assign io_coef_out_payload_0_34_4_imag = int_reg_array_34_4_imag;
  assign io_coef_out_payload_0_34_5_real = int_reg_array_34_5_real;
  assign io_coef_out_payload_0_34_5_imag = int_reg_array_34_5_imag;
  assign io_coef_out_payload_0_34_6_real = int_reg_array_34_6_real;
  assign io_coef_out_payload_0_34_6_imag = int_reg_array_34_6_imag;
  assign io_coef_out_payload_0_34_7_real = int_reg_array_34_7_real;
  assign io_coef_out_payload_0_34_7_imag = int_reg_array_34_7_imag;
  assign io_coef_out_payload_0_34_8_real = int_reg_array_34_8_real;
  assign io_coef_out_payload_0_34_8_imag = int_reg_array_34_8_imag;
  assign io_coef_out_payload_0_34_9_real = int_reg_array_34_9_real;
  assign io_coef_out_payload_0_34_9_imag = int_reg_array_34_9_imag;
  assign io_coef_out_payload_0_34_10_real = int_reg_array_34_10_real;
  assign io_coef_out_payload_0_34_10_imag = int_reg_array_34_10_imag;
  assign io_coef_out_payload_0_34_11_real = int_reg_array_34_11_real;
  assign io_coef_out_payload_0_34_11_imag = int_reg_array_34_11_imag;
  assign io_coef_out_payload_0_34_12_real = int_reg_array_34_12_real;
  assign io_coef_out_payload_0_34_12_imag = int_reg_array_34_12_imag;
  assign io_coef_out_payload_0_34_13_real = int_reg_array_34_13_real;
  assign io_coef_out_payload_0_34_13_imag = int_reg_array_34_13_imag;
  assign io_coef_out_payload_0_34_14_real = int_reg_array_34_14_real;
  assign io_coef_out_payload_0_34_14_imag = int_reg_array_34_14_imag;
  assign io_coef_out_payload_0_34_15_real = int_reg_array_34_15_real;
  assign io_coef_out_payload_0_34_15_imag = int_reg_array_34_15_imag;
  assign io_coef_out_payload_0_34_16_real = int_reg_array_34_16_real;
  assign io_coef_out_payload_0_34_16_imag = int_reg_array_34_16_imag;
  assign io_coef_out_payload_0_34_17_real = int_reg_array_34_17_real;
  assign io_coef_out_payload_0_34_17_imag = int_reg_array_34_17_imag;
  assign io_coef_out_payload_0_34_18_real = int_reg_array_34_18_real;
  assign io_coef_out_payload_0_34_18_imag = int_reg_array_34_18_imag;
  assign io_coef_out_payload_0_34_19_real = int_reg_array_34_19_real;
  assign io_coef_out_payload_0_34_19_imag = int_reg_array_34_19_imag;
  assign io_coef_out_payload_0_34_20_real = int_reg_array_34_20_real;
  assign io_coef_out_payload_0_34_20_imag = int_reg_array_34_20_imag;
  assign io_coef_out_payload_0_34_21_real = int_reg_array_34_21_real;
  assign io_coef_out_payload_0_34_21_imag = int_reg_array_34_21_imag;
  assign io_coef_out_payload_0_34_22_real = int_reg_array_34_22_real;
  assign io_coef_out_payload_0_34_22_imag = int_reg_array_34_22_imag;
  assign io_coef_out_payload_0_34_23_real = int_reg_array_34_23_real;
  assign io_coef_out_payload_0_34_23_imag = int_reg_array_34_23_imag;
  assign io_coef_out_payload_0_34_24_real = int_reg_array_34_24_real;
  assign io_coef_out_payload_0_34_24_imag = int_reg_array_34_24_imag;
  assign io_coef_out_payload_0_34_25_real = int_reg_array_34_25_real;
  assign io_coef_out_payload_0_34_25_imag = int_reg_array_34_25_imag;
  assign io_coef_out_payload_0_34_26_real = int_reg_array_34_26_real;
  assign io_coef_out_payload_0_34_26_imag = int_reg_array_34_26_imag;
  assign io_coef_out_payload_0_34_27_real = int_reg_array_34_27_real;
  assign io_coef_out_payload_0_34_27_imag = int_reg_array_34_27_imag;
  assign io_coef_out_payload_0_34_28_real = int_reg_array_34_28_real;
  assign io_coef_out_payload_0_34_28_imag = int_reg_array_34_28_imag;
  assign io_coef_out_payload_0_34_29_real = int_reg_array_34_29_real;
  assign io_coef_out_payload_0_34_29_imag = int_reg_array_34_29_imag;
  assign io_coef_out_payload_0_34_30_real = int_reg_array_34_30_real;
  assign io_coef_out_payload_0_34_30_imag = int_reg_array_34_30_imag;
  assign io_coef_out_payload_0_34_31_real = int_reg_array_34_31_real;
  assign io_coef_out_payload_0_34_31_imag = int_reg_array_34_31_imag;
  assign io_coef_out_payload_0_34_32_real = int_reg_array_34_32_real;
  assign io_coef_out_payload_0_34_32_imag = int_reg_array_34_32_imag;
  assign io_coef_out_payload_0_34_33_real = int_reg_array_34_33_real;
  assign io_coef_out_payload_0_34_33_imag = int_reg_array_34_33_imag;
  assign io_coef_out_payload_0_34_34_real = int_reg_array_34_34_real;
  assign io_coef_out_payload_0_34_34_imag = int_reg_array_34_34_imag;
  assign io_coef_out_payload_0_34_35_real = int_reg_array_34_35_real;
  assign io_coef_out_payload_0_34_35_imag = int_reg_array_34_35_imag;
  assign io_coef_out_payload_0_34_36_real = int_reg_array_34_36_real;
  assign io_coef_out_payload_0_34_36_imag = int_reg_array_34_36_imag;
  assign io_coef_out_payload_0_34_37_real = int_reg_array_34_37_real;
  assign io_coef_out_payload_0_34_37_imag = int_reg_array_34_37_imag;
  assign io_coef_out_payload_0_34_38_real = int_reg_array_34_38_real;
  assign io_coef_out_payload_0_34_38_imag = int_reg_array_34_38_imag;
  assign io_coef_out_payload_0_34_39_real = int_reg_array_34_39_real;
  assign io_coef_out_payload_0_34_39_imag = int_reg_array_34_39_imag;
  assign io_coef_out_payload_0_34_40_real = int_reg_array_34_40_real;
  assign io_coef_out_payload_0_34_40_imag = int_reg_array_34_40_imag;
  assign io_coef_out_payload_0_34_41_real = int_reg_array_34_41_real;
  assign io_coef_out_payload_0_34_41_imag = int_reg_array_34_41_imag;
  assign io_coef_out_payload_0_34_42_real = int_reg_array_34_42_real;
  assign io_coef_out_payload_0_34_42_imag = int_reg_array_34_42_imag;
  assign io_coef_out_payload_0_34_43_real = int_reg_array_34_43_real;
  assign io_coef_out_payload_0_34_43_imag = int_reg_array_34_43_imag;
  assign io_coef_out_payload_0_34_44_real = int_reg_array_34_44_real;
  assign io_coef_out_payload_0_34_44_imag = int_reg_array_34_44_imag;
  assign io_coef_out_payload_0_34_45_real = int_reg_array_34_45_real;
  assign io_coef_out_payload_0_34_45_imag = int_reg_array_34_45_imag;
  assign io_coef_out_payload_0_34_46_real = int_reg_array_34_46_real;
  assign io_coef_out_payload_0_34_46_imag = int_reg_array_34_46_imag;
  assign io_coef_out_payload_0_34_47_real = int_reg_array_34_47_real;
  assign io_coef_out_payload_0_34_47_imag = int_reg_array_34_47_imag;
  assign io_coef_out_payload_0_34_48_real = int_reg_array_34_48_real;
  assign io_coef_out_payload_0_34_48_imag = int_reg_array_34_48_imag;
  assign io_coef_out_payload_0_34_49_real = int_reg_array_34_49_real;
  assign io_coef_out_payload_0_34_49_imag = int_reg_array_34_49_imag;
  assign io_coef_out_payload_0_35_0_real = int_reg_array_35_0_real;
  assign io_coef_out_payload_0_35_0_imag = int_reg_array_35_0_imag;
  assign io_coef_out_payload_0_35_1_real = int_reg_array_35_1_real;
  assign io_coef_out_payload_0_35_1_imag = int_reg_array_35_1_imag;
  assign io_coef_out_payload_0_35_2_real = int_reg_array_35_2_real;
  assign io_coef_out_payload_0_35_2_imag = int_reg_array_35_2_imag;
  assign io_coef_out_payload_0_35_3_real = int_reg_array_35_3_real;
  assign io_coef_out_payload_0_35_3_imag = int_reg_array_35_3_imag;
  assign io_coef_out_payload_0_35_4_real = int_reg_array_35_4_real;
  assign io_coef_out_payload_0_35_4_imag = int_reg_array_35_4_imag;
  assign io_coef_out_payload_0_35_5_real = int_reg_array_35_5_real;
  assign io_coef_out_payload_0_35_5_imag = int_reg_array_35_5_imag;
  assign io_coef_out_payload_0_35_6_real = int_reg_array_35_6_real;
  assign io_coef_out_payload_0_35_6_imag = int_reg_array_35_6_imag;
  assign io_coef_out_payload_0_35_7_real = int_reg_array_35_7_real;
  assign io_coef_out_payload_0_35_7_imag = int_reg_array_35_7_imag;
  assign io_coef_out_payload_0_35_8_real = int_reg_array_35_8_real;
  assign io_coef_out_payload_0_35_8_imag = int_reg_array_35_8_imag;
  assign io_coef_out_payload_0_35_9_real = int_reg_array_35_9_real;
  assign io_coef_out_payload_0_35_9_imag = int_reg_array_35_9_imag;
  assign io_coef_out_payload_0_35_10_real = int_reg_array_35_10_real;
  assign io_coef_out_payload_0_35_10_imag = int_reg_array_35_10_imag;
  assign io_coef_out_payload_0_35_11_real = int_reg_array_35_11_real;
  assign io_coef_out_payload_0_35_11_imag = int_reg_array_35_11_imag;
  assign io_coef_out_payload_0_35_12_real = int_reg_array_35_12_real;
  assign io_coef_out_payload_0_35_12_imag = int_reg_array_35_12_imag;
  assign io_coef_out_payload_0_35_13_real = int_reg_array_35_13_real;
  assign io_coef_out_payload_0_35_13_imag = int_reg_array_35_13_imag;
  assign io_coef_out_payload_0_35_14_real = int_reg_array_35_14_real;
  assign io_coef_out_payload_0_35_14_imag = int_reg_array_35_14_imag;
  assign io_coef_out_payload_0_35_15_real = int_reg_array_35_15_real;
  assign io_coef_out_payload_0_35_15_imag = int_reg_array_35_15_imag;
  assign io_coef_out_payload_0_35_16_real = int_reg_array_35_16_real;
  assign io_coef_out_payload_0_35_16_imag = int_reg_array_35_16_imag;
  assign io_coef_out_payload_0_35_17_real = int_reg_array_35_17_real;
  assign io_coef_out_payload_0_35_17_imag = int_reg_array_35_17_imag;
  assign io_coef_out_payload_0_35_18_real = int_reg_array_35_18_real;
  assign io_coef_out_payload_0_35_18_imag = int_reg_array_35_18_imag;
  assign io_coef_out_payload_0_35_19_real = int_reg_array_35_19_real;
  assign io_coef_out_payload_0_35_19_imag = int_reg_array_35_19_imag;
  assign io_coef_out_payload_0_35_20_real = int_reg_array_35_20_real;
  assign io_coef_out_payload_0_35_20_imag = int_reg_array_35_20_imag;
  assign io_coef_out_payload_0_35_21_real = int_reg_array_35_21_real;
  assign io_coef_out_payload_0_35_21_imag = int_reg_array_35_21_imag;
  assign io_coef_out_payload_0_35_22_real = int_reg_array_35_22_real;
  assign io_coef_out_payload_0_35_22_imag = int_reg_array_35_22_imag;
  assign io_coef_out_payload_0_35_23_real = int_reg_array_35_23_real;
  assign io_coef_out_payload_0_35_23_imag = int_reg_array_35_23_imag;
  assign io_coef_out_payload_0_35_24_real = int_reg_array_35_24_real;
  assign io_coef_out_payload_0_35_24_imag = int_reg_array_35_24_imag;
  assign io_coef_out_payload_0_35_25_real = int_reg_array_35_25_real;
  assign io_coef_out_payload_0_35_25_imag = int_reg_array_35_25_imag;
  assign io_coef_out_payload_0_35_26_real = int_reg_array_35_26_real;
  assign io_coef_out_payload_0_35_26_imag = int_reg_array_35_26_imag;
  assign io_coef_out_payload_0_35_27_real = int_reg_array_35_27_real;
  assign io_coef_out_payload_0_35_27_imag = int_reg_array_35_27_imag;
  assign io_coef_out_payload_0_35_28_real = int_reg_array_35_28_real;
  assign io_coef_out_payload_0_35_28_imag = int_reg_array_35_28_imag;
  assign io_coef_out_payload_0_35_29_real = int_reg_array_35_29_real;
  assign io_coef_out_payload_0_35_29_imag = int_reg_array_35_29_imag;
  assign io_coef_out_payload_0_35_30_real = int_reg_array_35_30_real;
  assign io_coef_out_payload_0_35_30_imag = int_reg_array_35_30_imag;
  assign io_coef_out_payload_0_35_31_real = int_reg_array_35_31_real;
  assign io_coef_out_payload_0_35_31_imag = int_reg_array_35_31_imag;
  assign io_coef_out_payload_0_35_32_real = int_reg_array_35_32_real;
  assign io_coef_out_payload_0_35_32_imag = int_reg_array_35_32_imag;
  assign io_coef_out_payload_0_35_33_real = int_reg_array_35_33_real;
  assign io_coef_out_payload_0_35_33_imag = int_reg_array_35_33_imag;
  assign io_coef_out_payload_0_35_34_real = int_reg_array_35_34_real;
  assign io_coef_out_payload_0_35_34_imag = int_reg_array_35_34_imag;
  assign io_coef_out_payload_0_35_35_real = int_reg_array_35_35_real;
  assign io_coef_out_payload_0_35_35_imag = int_reg_array_35_35_imag;
  assign io_coef_out_payload_0_35_36_real = int_reg_array_35_36_real;
  assign io_coef_out_payload_0_35_36_imag = int_reg_array_35_36_imag;
  assign io_coef_out_payload_0_35_37_real = int_reg_array_35_37_real;
  assign io_coef_out_payload_0_35_37_imag = int_reg_array_35_37_imag;
  assign io_coef_out_payload_0_35_38_real = int_reg_array_35_38_real;
  assign io_coef_out_payload_0_35_38_imag = int_reg_array_35_38_imag;
  assign io_coef_out_payload_0_35_39_real = int_reg_array_35_39_real;
  assign io_coef_out_payload_0_35_39_imag = int_reg_array_35_39_imag;
  assign io_coef_out_payload_0_35_40_real = int_reg_array_35_40_real;
  assign io_coef_out_payload_0_35_40_imag = int_reg_array_35_40_imag;
  assign io_coef_out_payload_0_35_41_real = int_reg_array_35_41_real;
  assign io_coef_out_payload_0_35_41_imag = int_reg_array_35_41_imag;
  assign io_coef_out_payload_0_35_42_real = int_reg_array_35_42_real;
  assign io_coef_out_payload_0_35_42_imag = int_reg_array_35_42_imag;
  assign io_coef_out_payload_0_35_43_real = int_reg_array_35_43_real;
  assign io_coef_out_payload_0_35_43_imag = int_reg_array_35_43_imag;
  assign io_coef_out_payload_0_35_44_real = int_reg_array_35_44_real;
  assign io_coef_out_payload_0_35_44_imag = int_reg_array_35_44_imag;
  assign io_coef_out_payload_0_35_45_real = int_reg_array_35_45_real;
  assign io_coef_out_payload_0_35_45_imag = int_reg_array_35_45_imag;
  assign io_coef_out_payload_0_35_46_real = int_reg_array_35_46_real;
  assign io_coef_out_payload_0_35_46_imag = int_reg_array_35_46_imag;
  assign io_coef_out_payload_0_35_47_real = int_reg_array_35_47_real;
  assign io_coef_out_payload_0_35_47_imag = int_reg_array_35_47_imag;
  assign io_coef_out_payload_0_35_48_real = int_reg_array_35_48_real;
  assign io_coef_out_payload_0_35_48_imag = int_reg_array_35_48_imag;
  assign io_coef_out_payload_0_35_49_real = int_reg_array_35_49_real;
  assign io_coef_out_payload_0_35_49_imag = int_reg_array_35_49_imag;
  assign io_coef_out_payload_0_36_0_real = int_reg_array_36_0_real;
  assign io_coef_out_payload_0_36_0_imag = int_reg_array_36_0_imag;
  assign io_coef_out_payload_0_36_1_real = int_reg_array_36_1_real;
  assign io_coef_out_payload_0_36_1_imag = int_reg_array_36_1_imag;
  assign io_coef_out_payload_0_36_2_real = int_reg_array_36_2_real;
  assign io_coef_out_payload_0_36_2_imag = int_reg_array_36_2_imag;
  assign io_coef_out_payload_0_36_3_real = int_reg_array_36_3_real;
  assign io_coef_out_payload_0_36_3_imag = int_reg_array_36_3_imag;
  assign io_coef_out_payload_0_36_4_real = int_reg_array_36_4_real;
  assign io_coef_out_payload_0_36_4_imag = int_reg_array_36_4_imag;
  assign io_coef_out_payload_0_36_5_real = int_reg_array_36_5_real;
  assign io_coef_out_payload_0_36_5_imag = int_reg_array_36_5_imag;
  assign io_coef_out_payload_0_36_6_real = int_reg_array_36_6_real;
  assign io_coef_out_payload_0_36_6_imag = int_reg_array_36_6_imag;
  assign io_coef_out_payload_0_36_7_real = int_reg_array_36_7_real;
  assign io_coef_out_payload_0_36_7_imag = int_reg_array_36_7_imag;
  assign io_coef_out_payload_0_36_8_real = int_reg_array_36_8_real;
  assign io_coef_out_payload_0_36_8_imag = int_reg_array_36_8_imag;
  assign io_coef_out_payload_0_36_9_real = int_reg_array_36_9_real;
  assign io_coef_out_payload_0_36_9_imag = int_reg_array_36_9_imag;
  assign io_coef_out_payload_0_36_10_real = int_reg_array_36_10_real;
  assign io_coef_out_payload_0_36_10_imag = int_reg_array_36_10_imag;
  assign io_coef_out_payload_0_36_11_real = int_reg_array_36_11_real;
  assign io_coef_out_payload_0_36_11_imag = int_reg_array_36_11_imag;
  assign io_coef_out_payload_0_36_12_real = int_reg_array_36_12_real;
  assign io_coef_out_payload_0_36_12_imag = int_reg_array_36_12_imag;
  assign io_coef_out_payload_0_36_13_real = int_reg_array_36_13_real;
  assign io_coef_out_payload_0_36_13_imag = int_reg_array_36_13_imag;
  assign io_coef_out_payload_0_36_14_real = int_reg_array_36_14_real;
  assign io_coef_out_payload_0_36_14_imag = int_reg_array_36_14_imag;
  assign io_coef_out_payload_0_36_15_real = int_reg_array_36_15_real;
  assign io_coef_out_payload_0_36_15_imag = int_reg_array_36_15_imag;
  assign io_coef_out_payload_0_36_16_real = int_reg_array_36_16_real;
  assign io_coef_out_payload_0_36_16_imag = int_reg_array_36_16_imag;
  assign io_coef_out_payload_0_36_17_real = int_reg_array_36_17_real;
  assign io_coef_out_payload_0_36_17_imag = int_reg_array_36_17_imag;
  assign io_coef_out_payload_0_36_18_real = int_reg_array_36_18_real;
  assign io_coef_out_payload_0_36_18_imag = int_reg_array_36_18_imag;
  assign io_coef_out_payload_0_36_19_real = int_reg_array_36_19_real;
  assign io_coef_out_payload_0_36_19_imag = int_reg_array_36_19_imag;
  assign io_coef_out_payload_0_36_20_real = int_reg_array_36_20_real;
  assign io_coef_out_payload_0_36_20_imag = int_reg_array_36_20_imag;
  assign io_coef_out_payload_0_36_21_real = int_reg_array_36_21_real;
  assign io_coef_out_payload_0_36_21_imag = int_reg_array_36_21_imag;
  assign io_coef_out_payload_0_36_22_real = int_reg_array_36_22_real;
  assign io_coef_out_payload_0_36_22_imag = int_reg_array_36_22_imag;
  assign io_coef_out_payload_0_36_23_real = int_reg_array_36_23_real;
  assign io_coef_out_payload_0_36_23_imag = int_reg_array_36_23_imag;
  assign io_coef_out_payload_0_36_24_real = int_reg_array_36_24_real;
  assign io_coef_out_payload_0_36_24_imag = int_reg_array_36_24_imag;
  assign io_coef_out_payload_0_36_25_real = int_reg_array_36_25_real;
  assign io_coef_out_payload_0_36_25_imag = int_reg_array_36_25_imag;
  assign io_coef_out_payload_0_36_26_real = int_reg_array_36_26_real;
  assign io_coef_out_payload_0_36_26_imag = int_reg_array_36_26_imag;
  assign io_coef_out_payload_0_36_27_real = int_reg_array_36_27_real;
  assign io_coef_out_payload_0_36_27_imag = int_reg_array_36_27_imag;
  assign io_coef_out_payload_0_36_28_real = int_reg_array_36_28_real;
  assign io_coef_out_payload_0_36_28_imag = int_reg_array_36_28_imag;
  assign io_coef_out_payload_0_36_29_real = int_reg_array_36_29_real;
  assign io_coef_out_payload_0_36_29_imag = int_reg_array_36_29_imag;
  assign io_coef_out_payload_0_36_30_real = int_reg_array_36_30_real;
  assign io_coef_out_payload_0_36_30_imag = int_reg_array_36_30_imag;
  assign io_coef_out_payload_0_36_31_real = int_reg_array_36_31_real;
  assign io_coef_out_payload_0_36_31_imag = int_reg_array_36_31_imag;
  assign io_coef_out_payload_0_36_32_real = int_reg_array_36_32_real;
  assign io_coef_out_payload_0_36_32_imag = int_reg_array_36_32_imag;
  assign io_coef_out_payload_0_36_33_real = int_reg_array_36_33_real;
  assign io_coef_out_payload_0_36_33_imag = int_reg_array_36_33_imag;
  assign io_coef_out_payload_0_36_34_real = int_reg_array_36_34_real;
  assign io_coef_out_payload_0_36_34_imag = int_reg_array_36_34_imag;
  assign io_coef_out_payload_0_36_35_real = int_reg_array_36_35_real;
  assign io_coef_out_payload_0_36_35_imag = int_reg_array_36_35_imag;
  assign io_coef_out_payload_0_36_36_real = int_reg_array_36_36_real;
  assign io_coef_out_payload_0_36_36_imag = int_reg_array_36_36_imag;
  assign io_coef_out_payload_0_36_37_real = int_reg_array_36_37_real;
  assign io_coef_out_payload_0_36_37_imag = int_reg_array_36_37_imag;
  assign io_coef_out_payload_0_36_38_real = int_reg_array_36_38_real;
  assign io_coef_out_payload_0_36_38_imag = int_reg_array_36_38_imag;
  assign io_coef_out_payload_0_36_39_real = int_reg_array_36_39_real;
  assign io_coef_out_payload_0_36_39_imag = int_reg_array_36_39_imag;
  assign io_coef_out_payload_0_36_40_real = int_reg_array_36_40_real;
  assign io_coef_out_payload_0_36_40_imag = int_reg_array_36_40_imag;
  assign io_coef_out_payload_0_36_41_real = int_reg_array_36_41_real;
  assign io_coef_out_payload_0_36_41_imag = int_reg_array_36_41_imag;
  assign io_coef_out_payload_0_36_42_real = int_reg_array_36_42_real;
  assign io_coef_out_payload_0_36_42_imag = int_reg_array_36_42_imag;
  assign io_coef_out_payload_0_36_43_real = int_reg_array_36_43_real;
  assign io_coef_out_payload_0_36_43_imag = int_reg_array_36_43_imag;
  assign io_coef_out_payload_0_36_44_real = int_reg_array_36_44_real;
  assign io_coef_out_payload_0_36_44_imag = int_reg_array_36_44_imag;
  assign io_coef_out_payload_0_36_45_real = int_reg_array_36_45_real;
  assign io_coef_out_payload_0_36_45_imag = int_reg_array_36_45_imag;
  assign io_coef_out_payload_0_36_46_real = int_reg_array_36_46_real;
  assign io_coef_out_payload_0_36_46_imag = int_reg_array_36_46_imag;
  assign io_coef_out_payload_0_36_47_real = int_reg_array_36_47_real;
  assign io_coef_out_payload_0_36_47_imag = int_reg_array_36_47_imag;
  assign io_coef_out_payload_0_36_48_real = int_reg_array_36_48_real;
  assign io_coef_out_payload_0_36_48_imag = int_reg_array_36_48_imag;
  assign io_coef_out_payload_0_36_49_real = int_reg_array_36_49_real;
  assign io_coef_out_payload_0_36_49_imag = int_reg_array_36_49_imag;
  assign io_coef_out_payload_0_37_0_real = int_reg_array_37_0_real;
  assign io_coef_out_payload_0_37_0_imag = int_reg_array_37_0_imag;
  assign io_coef_out_payload_0_37_1_real = int_reg_array_37_1_real;
  assign io_coef_out_payload_0_37_1_imag = int_reg_array_37_1_imag;
  assign io_coef_out_payload_0_37_2_real = int_reg_array_37_2_real;
  assign io_coef_out_payload_0_37_2_imag = int_reg_array_37_2_imag;
  assign io_coef_out_payload_0_37_3_real = int_reg_array_37_3_real;
  assign io_coef_out_payload_0_37_3_imag = int_reg_array_37_3_imag;
  assign io_coef_out_payload_0_37_4_real = int_reg_array_37_4_real;
  assign io_coef_out_payload_0_37_4_imag = int_reg_array_37_4_imag;
  assign io_coef_out_payload_0_37_5_real = int_reg_array_37_5_real;
  assign io_coef_out_payload_0_37_5_imag = int_reg_array_37_5_imag;
  assign io_coef_out_payload_0_37_6_real = int_reg_array_37_6_real;
  assign io_coef_out_payload_0_37_6_imag = int_reg_array_37_6_imag;
  assign io_coef_out_payload_0_37_7_real = int_reg_array_37_7_real;
  assign io_coef_out_payload_0_37_7_imag = int_reg_array_37_7_imag;
  assign io_coef_out_payload_0_37_8_real = int_reg_array_37_8_real;
  assign io_coef_out_payload_0_37_8_imag = int_reg_array_37_8_imag;
  assign io_coef_out_payload_0_37_9_real = int_reg_array_37_9_real;
  assign io_coef_out_payload_0_37_9_imag = int_reg_array_37_9_imag;
  assign io_coef_out_payload_0_37_10_real = int_reg_array_37_10_real;
  assign io_coef_out_payload_0_37_10_imag = int_reg_array_37_10_imag;
  assign io_coef_out_payload_0_37_11_real = int_reg_array_37_11_real;
  assign io_coef_out_payload_0_37_11_imag = int_reg_array_37_11_imag;
  assign io_coef_out_payload_0_37_12_real = int_reg_array_37_12_real;
  assign io_coef_out_payload_0_37_12_imag = int_reg_array_37_12_imag;
  assign io_coef_out_payload_0_37_13_real = int_reg_array_37_13_real;
  assign io_coef_out_payload_0_37_13_imag = int_reg_array_37_13_imag;
  assign io_coef_out_payload_0_37_14_real = int_reg_array_37_14_real;
  assign io_coef_out_payload_0_37_14_imag = int_reg_array_37_14_imag;
  assign io_coef_out_payload_0_37_15_real = int_reg_array_37_15_real;
  assign io_coef_out_payload_0_37_15_imag = int_reg_array_37_15_imag;
  assign io_coef_out_payload_0_37_16_real = int_reg_array_37_16_real;
  assign io_coef_out_payload_0_37_16_imag = int_reg_array_37_16_imag;
  assign io_coef_out_payload_0_37_17_real = int_reg_array_37_17_real;
  assign io_coef_out_payload_0_37_17_imag = int_reg_array_37_17_imag;
  assign io_coef_out_payload_0_37_18_real = int_reg_array_37_18_real;
  assign io_coef_out_payload_0_37_18_imag = int_reg_array_37_18_imag;
  assign io_coef_out_payload_0_37_19_real = int_reg_array_37_19_real;
  assign io_coef_out_payload_0_37_19_imag = int_reg_array_37_19_imag;
  assign io_coef_out_payload_0_37_20_real = int_reg_array_37_20_real;
  assign io_coef_out_payload_0_37_20_imag = int_reg_array_37_20_imag;
  assign io_coef_out_payload_0_37_21_real = int_reg_array_37_21_real;
  assign io_coef_out_payload_0_37_21_imag = int_reg_array_37_21_imag;
  assign io_coef_out_payload_0_37_22_real = int_reg_array_37_22_real;
  assign io_coef_out_payload_0_37_22_imag = int_reg_array_37_22_imag;
  assign io_coef_out_payload_0_37_23_real = int_reg_array_37_23_real;
  assign io_coef_out_payload_0_37_23_imag = int_reg_array_37_23_imag;
  assign io_coef_out_payload_0_37_24_real = int_reg_array_37_24_real;
  assign io_coef_out_payload_0_37_24_imag = int_reg_array_37_24_imag;
  assign io_coef_out_payload_0_37_25_real = int_reg_array_37_25_real;
  assign io_coef_out_payload_0_37_25_imag = int_reg_array_37_25_imag;
  assign io_coef_out_payload_0_37_26_real = int_reg_array_37_26_real;
  assign io_coef_out_payload_0_37_26_imag = int_reg_array_37_26_imag;
  assign io_coef_out_payload_0_37_27_real = int_reg_array_37_27_real;
  assign io_coef_out_payload_0_37_27_imag = int_reg_array_37_27_imag;
  assign io_coef_out_payload_0_37_28_real = int_reg_array_37_28_real;
  assign io_coef_out_payload_0_37_28_imag = int_reg_array_37_28_imag;
  assign io_coef_out_payload_0_37_29_real = int_reg_array_37_29_real;
  assign io_coef_out_payload_0_37_29_imag = int_reg_array_37_29_imag;
  assign io_coef_out_payload_0_37_30_real = int_reg_array_37_30_real;
  assign io_coef_out_payload_0_37_30_imag = int_reg_array_37_30_imag;
  assign io_coef_out_payload_0_37_31_real = int_reg_array_37_31_real;
  assign io_coef_out_payload_0_37_31_imag = int_reg_array_37_31_imag;
  assign io_coef_out_payload_0_37_32_real = int_reg_array_37_32_real;
  assign io_coef_out_payload_0_37_32_imag = int_reg_array_37_32_imag;
  assign io_coef_out_payload_0_37_33_real = int_reg_array_37_33_real;
  assign io_coef_out_payload_0_37_33_imag = int_reg_array_37_33_imag;
  assign io_coef_out_payload_0_37_34_real = int_reg_array_37_34_real;
  assign io_coef_out_payload_0_37_34_imag = int_reg_array_37_34_imag;
  assign io_coef_out_payload_0_37_35_real = int_reg_array_37_35_real;
  assign io_coef_out_payload_0_37_35_imag = int_reg_array_37_35_imag;
  assign io_coef_out_payload_0_37_36_real = int_reg_array_37_36_real;
  assign io_coef_out_payload_0_37_36_imag = int_reg_array_37_36_imag;
  assign io_coef_out_payload_0_37_37_real = int_reg_array_37_37_real;
  assign io_coef_out_payload_0_37_37_imag = int_reg_array_37_37_imag;
  assign io_coef_out_payload_0_37_38_real = int_reg_array_37_38_real;
  assign io_coef_out_payload_0_37_38_imag = int_reg_array_37_38_imag;
  assign io_coef_out_payload_0_37_39_real = int_reg_array_37_39_real;
  assign io_coef_out_payload_0_37_39_imag = int_reg_array_37_39_imag;
  assign io_coef_out_payload_0_37_40_real = int_reg_array_37_40_real;
  assign io_coef_out_payload_0_37_40_imag = int_reg_array_37_40_imag;
  assign io_coef_out_payload_0_37_41_real = int_reg_array_37_41_real;
  assign io_coef_out_payload_0_37_41_imag = int_reg_array_37_41_imag;
  assign io_coef_out_payload_0_37_42_real = int_reg_array_37_42_real;
  assign io_coef_out_payload_0_37_42_imag = int_reg_array_37_42_imag;
  assign io_coef_out_payload_0_37_43_real = int_reg_array_37_43_real;
  assign io_coef_out_payload_0_37_43_imag = int_reg_array_37_43_imag;
  assign io_coef_out_payload_0_37_44_real = int_reg_array_37_44_real;
  assign io_coef_out_payload_0_37_44_imag = int_reg_array_37_44_imag;
  assign io_coef_out_payload_0_37_45_real = int_reg_array_37_45_real;
  assign io_coef_out_payload_0_37_45_imag = int_reg_array_37_45_imag;
  assign io_coef_out_payload_0_37_46_real = int_reg_array_37_46_real;
  assign io_coef_out_payload_0_37_46_imag = int_reg_array_37_46_imag;
  assign io_coef_out_payload_0_37_47_real = int_reg_array_37_47_real;
  assign io_coef_out_payload_0_37_47_imag = int_reg_array_37_47_imag;
  assign io_coef_out_payload_0_37_48_real = int_reg_array_37_48_real;
  assign io_coef_out_payload_0_37_48_imag = int_reg_array_37_48_imag;
  assign io_coef_out_payload_0_37_49_real = int_reg_array_37_49_real;
  assign io_coef_out_payload_0_37_49_imag = int_reg_array_37_49_imag;
  assign io_coef_out_payload_0_38_0_real = int_reg_array_38_0_real;
  assign io_coef_out_payload_0_38_0_imag = int_reg_array_38_0_imag;
  assign io_coef_out_payload_0_38_1_real = int_reg_array_38_1_real;
  assign io_coef_out_payload_0_38_1_imag = int_reg_array_38_1_imag;
  assign io_coef_out_payload_0_38_2_real = int_reg_array_38_2_real;
  assign io_coef_out_payload_0_38_2_imag = int_reg_array_38_2_imag;
  assign io_coef_out_payload_0_38_3_real = int_reg_array_38_3_real;
  assign io_coef_out_payload_0_38_3_imag = int_reg_array_38_3_imag;
  assign io_coef_out_payload_0_38_4_real = int_reg_array_38_4_real;
  assign io_coef_out_payload_0_38_4_imag = int_reg_array_38_4_imag;
  assign io_coef_out_payload_0_38_5_real = int_reg_array_38_5_real;
  assign io_coef_out_payload_0_38_5_imag = int_reg_array_38_5_imag;
  assign io_coef_out_payload_0_38_6_real = int_reg_array_38_6_real;
  assign io_coef_out_payload_0_38_6_imag = int_reg_array_38_6_imag;
  assign io_coef_out_payload_0_38_7_real = int_reg_array_38_7_real;
  assign io_coef_out_payload_0_38_7_imag = int_reg_array_38_7_imag;
  assign io_coef_out_payload_0_38_8_real = int_reg_array_38_8_real;
  assign io_coef_out_payload_0_38_8_imag = int_reg_array_38_8_imag;
  assign io_coef_out_payload_0_38_9_real = int_reg_array_38_9_real;
  assign io_coef_out_payload_0_38_9_imag = int_reg_array_38_9_imag;
  assign io_coef_out_payload_0_38_10_real = int_reg_array_38_10_real;
  assign io_coef_out_payload_0_38_10_imag = int_reg_array_38_10_imag;
  assign io_coef_out_payload_0_38_11_real = int_reg_array_38_11_real;
  assign io_coef_out_payload_0_38_11_imag = int_reg_array_38_11_imag;
  assign io_coef_out_payload_0_38_12_real = int_reg_array_38_12_real;
  assign io_coef_out_payload_0_38_12_imag = int_reg_array_38_12_imag;
  assign io_coef_out_payload_0_38_13_real = int_reg_array_38_13_real;
  assign io_coef_out_payload_0_38_13_imag = int_reg_array_38_13_imag;
  assign io_coef_out_payload_0_38_14_real = int_reg_array_38_14_real;
  assign io_coef_out_payload_0_38_14_imag = int_reg_array_38_14_imag;
  assign io_coef_out_payload_0_38_15_real = int_reg_array_38_15_real;
  assign io_coef_out_payload_0_38_15_imag = int_reg_array_38_15_imag;
  assign io_coef_out_payload_0_38_16_real = int_reg_array_38_16_real;
  assign io_coef_out_payload_0_38_16_imag = int_reg_array_38_16_imag;
  assign io_coef_out_payload_0_38_17_real = int_reg_array_38_17_real;
  assign io_coef_out_payload_0_38_17_imag = int_reg_array_38_17_imag;
  assign io_coef_out_payload_0_38_18_real = int_reg_array_38_18_real;
  assign io_coef_out_payload_0_38_18_imag = int_reg_array_38_18_imag;
  assign io_coef_out_payload_0_38_19_real = int_reg_array_38_19_real;
  assign io_coef_out_payload_0_38_19_imag = int_reg_array_38_19_imag;
  assign io_coef_out_payload_0_38_20_real = int_reg_array_38_20_real;
  assign io_coef_out_payload_0_38_20_imag = int_reg_array_38_20_imag;
  assign io_coef_out_payload_0_38_21_real = int_reg_array_38_21_real;
  assign io_coef_out_payload_0_38_21_imag = int_reg_array_38_21_imag;
  assign io_coef_out_payload_0_38_22_real = int_reg_array_38_22_real;
  assign io_coef_out_payload_0_38_22_imag = int_reg_array_38_22_imag;
  assign io_coef_out_payload_0_38_23_real = int_reg_array_38_23_real;
  assign io_coef_out_payload_0_38_23_imag = int_reg_array_38_23_imag;
  assign io_coef_out_payload_0_38_24_real = int_reg_array_38_24_real;
  assign io_coef_out_payload_0_38_24_imag = int_reg_array_38_24_imag;
  assign io_coef_out_payload_0_38_25_real = int_reg_array_38_25_real;
  assign io_coef_out_payload_0_38_25_imag = int_reg_array_38_25_imag;
  assign io_coef_out_payload_0_38_26_real = int_reg_array_38_26_real;
  assign io_coef_out_payload_0_38_26_imag = int_reg_array_38_26_imag;
  assign io_coef_out_payload_0_38_27_real = int_reg_array_38_27_real;
  assign io_coef_out_payload_0_38_27_imag = int_reg_array_38_27_imag;
  assign io_coef_out_payload_0_38_28_real = int_reg_array_38_28_real;
  assign io_coef_out_payload_0_38_28_imag = int_reg_array_38_28_imag;
  assign io_coef_out_payload_0_38_29_real = int_reg_array_38_29_real;
  assign io_coef_out_payload_0_38_29_imag = int_reg_array_38_29_imag;
  assign io_coef_out_payload_0_38_30_real = int_reg_array_38_30_real;
  assign io_coef_out_payload_0_38_30_imag = int_reg_array_38_30_imag;
  assign io_coef_out_payload_0_38_31_real = int_reg_array_38_31_real;
  assign io_coef_out_payload_0_38_31_imag = int_reg_array_38_31_imag;
  assign io_coef_out_payload_0_38_32_real = int_reg_array_38_32_real;
  assign io_coef_out_payload_0_38_32_imag = int_reg_array_38_32_imag;
  assign io_coef_out_payload_0_38_33_real = int_reg_array_38_33_real;
  assign io_coef_out_payload_0_38_33_imag = int_reg_array_38_33_imag;
  assign io_coef_out_payload_0_38_34_real = int_reg_array_38_34_real;
  assign io_coef_out_payload_0_38_34_imag = int_reg_array_38_34_imag;
  assign io_coef_out_payload_0_38_35_real = int_reg_array_38_35_real;
  assign io_coef_out_payload_0_38_35_imag = int_reg_array_38_35_imag;
  assign io_coef_out_payload_0_38_36_real = int_reg_array_38_36_real;
  assign io_coef_out_payload_0_38_36_imag = int_reg_array_38_36_imag;
  assign io_coef_out_payload_0_38_37_real = int_reg_array_38_37_real;
  assign io_coef_out_payload_0_38_37_imag = int_reg_array_38_37_imag;
  assign io_coef_out_payload_0_38_38_real = int_reg_array_38_38_real;
  assign io_coef_out_payload_0_38_38_imag = int_reg_array_38_38_imag;
  assign io_coef_out_payload_0_38_39_real = int_reg_array_38_39_real;
  assign io_coef_out_payload_0_38_39_imag = int_reg_array_38_39_imag;
  assign io_coef_out_payload_0_38_40_real = int_reg_array_38_40_real;
  assign io_coef_out_payload_0_38_40_imag = int_reg_array_38_40_imag;
  assign io_coef_out_payload_0_38_41_real = int_reg_array_38_41_real;
  assign io_coef_out_payload_0_38_41_imag = int_reg_array_38_41_imag;
  assign io_coef_out_payload_0_38_42_real = int_reg_array_38_42_real;
  assign io_coef_out_payload_0_38_42_imag = int_reg_array_38_42_imag;
  assign io_coef_out_payload_0_38_43_real = int_reg_array_38_43_real;
  assign io_coef_out_payload_0_38_43_imag = int_reg_array_38_43_imag;
  assign io_coef_out_payload_0_38_44_real = int_reg_array_38_44_real;
  assign io_coef_out_payload_0_38_44_imag = int_reg_array_38_44_imag;
  assign io_coef_out_payload_0_38_45_real = int_reg_array_38_45_real;
  assign io_coef_out_payload_0_38_45_imag = int_reg_array_38_45_imag;
  assign io_coef_out_payload_0_38_46_real = int_reg_array_38_46_real;
  assign io_coef_out_payload_0_38_46_imag = int_reg_array_38_46_imag;
  assign io_coef_out_payload_0_38_47_real = int_reg_array_38_47_real;
  assign io_coef_out_payload_0_38_47_imag = int_reg_array_38_47_imag;
  assign io_coef_out_payload_0_38_48_real = int_reg_array_38_48_real;
  assign io_coef_out_payload_0_38_48_imag = int_reg_array_38_48_imag;
  assign io_coef_out_payload_0_38_49_real = int_reg_array_38_49_real;
  assign io_coef_out_payload_0_38_49_imag = int_reg_array_38_49_imag;
  assign io_coef_out_payload_0_39_0_real = int_reg_array_39_0_real;
  assign io_coef_out_payload_0_39_0_imag = int_reg_array_39_0_imag;
  assign io_coef_out_payload_0_39_1_real = int_reg_array_39_1_real;
  assign io_coef_out_payload_0_39_1_imag = int_reg_array_39_1_imag;
  assign io_coef_out_payload_0_39_2_real = int_reg_array_39_2_real;
  assign io_coef_out_payload_0_39_2_imag = int_reg_array_39_2_imag;
  assign io_coef_out_payload_0_39_3_real = int_reg_array_39_3_real;
  assign io_coef_out_payload_0_39_3_imag = int_reg_array_39_3_imag;
  assign io_coef_out_payload_0_39_4_real = int_reg_array_39_4_real;
  assign io_coef_out_payload_0_39_4_imag = int_reg_array_39_4_imag;
  assign io_coef_out_payload_0_39_5_real = int_reg_array_39_5_real;
  assign io_coef_out_payload_0_39_5_imag = int_reg_array_39_5_imag;
  assign io_coef_out_payload_0_39_6_real = int_reg_array_39_6_real;
  assign io_coef_out_payload_0_39_6_imag = int_reg_array_39_6_imag;
  assign io_coef_out_payload_0_39_7_real = int_reg_array_39_7_real;
  assign io_coef_out_payload_0_39_7_imag = int_reg_array_39_7_imag;
  assign io_coef_out_payload_0_39_8_real = int_reg_array_39_8_real;
  assign io_coef_out_payload_0_39_8_imag = int_reg_array_39_8_imag;
  assign io_coef_out_payload_0_39_9_real = int_reg_array_39_9_real;
  assign io_coef_out_payload_0_39_9_imag = int_reg_array_39_9_imag;
  assign io_coef_out_payload_0_39_10_real = int_reg_array_39_10_real;
  assign io_coef_out_payload_0_39_10_imag = int_reg_array_39_10_imag;
  assign io_coef_out_payload_0_39_11_real = int_reg_array_39_11_real;
  assign io_coef_out_payload_0_39_11_imag = int_reg_array_39_11_imag;
  assign io_coef_out_payload_0_39_12_real = int_reg_array_39_12_real;
  assign io_coef_out_payload_0_39_12_imag = int_reg_array_39_12_imag;
  assign io_coef_out_payload_0_39_13_real = int_reg_array_39_13_real;
  assign io_coef_out_payload_0_39_13_imag = int_reg_array_39_13_imag;
  assign io_coef_out_payload_0_39_14_real = int_reg_array_39_14_real;
  assign io_coef_out_payload_0_39_14_imag = int_reg_array_39_14_imag;
  assign io_coef_out_payload_0_39_15_real = int_reg_array_39_15_real;
  assign io_coef_out_payload_0_39_15_imag = int_reg_array_39_15_imag;
  assign io_coef_out_payload_0_39_16_real = int_reg_array_39_16_real;
  assign io_coef_out_payload_0_39_16_imag = int_reg_array_39_16_imag;
  assign io_coef_out_payload_0_39_17_real = int_reg_array_39_17_real;
  assign io_coef_out_payload_0_39_17_imag = int_reg_array_39_17_imag;
  assign io_coef_out_payload_0_39_18_real = int_reg_array_39_18_real;
  assign io_coef_out_payload_0_39_18_imag = int_reg_array_39_18_imag;
  assign io_coef_out_payload_0_39_19_real = int_reg_array_39_19_real;
  assign io_coef_out_payload_0_39_19_imag = int_reg_array_39_19_imag;
  assign io_coef_out_payload_0_39_20_real = int_reg_array_39_20_real;
  assign io_coef_out_payload_0_39_20_imag = int_reg_array_39_20_imag;
  assign io_coef_out_payload_0_39_21_real = int_reg_array_39_21_real;
  assign io_coef_out_payload_0_39_21_imag = int_reg_array_39_21_imag;
  assign io_coef_out_payload_0_39_22_real = int_reg_array_39_22_real;
  assign io_coef_out_payload_0_39_22_imag = int_reg_array_39_22_imag;
  assign io_coef_out_payload_0_39_23_real = int_reg_array_39_23_real;
  assign io_coef_out_payload_0_39_23_imag = int_reg_array_39_23_imag;
  assign io_coef_out_payload_0_39_24_real = int_reg_array_39_24_real;
  assign io_coef_out_payload_0_39_24_imag = int_reg_array_39_24_imag;
  assign io_coef_out_payload_0_39_25_real = int_reg_array_39_25_real;
  assign io_coef_out_payload_0_39_25_imag = int_reg_array_39_25_imag;
  assign io_coef_out_payload_0_39_26_real = int_reg_array_39_26_real;
  assign io_coef_out_payload_0_39_26_imag = int_reg_array_39_26_imag;
  assign io_coef_out_payload_0_39_27_real = int_reg_array_39_27_real;
  assign io_coef_out_payload_0_39_27_imag = int_reg_array_39_27_imag;
  assign io_coef_out_payload_0_39_28_real = int_reg_array_39_28_real;
  assign io_coef_out_payload_0_39_28_imag = int_reg_array_39_28_imag;
  assign io_coef_out_payload_0_39_29_real = int_reg_array_39_29_real;
  assign io_coef_out_payload_0_39_29_imag = int_reg_array_39_29_imag;
  assign io_coef_out_payload_0_39_30_real = int_reg_array_39_30_real;
  assign io_coef_out_payload_0_39_30_imag = int_reg_array_39_30_imag;
  assign io_coef_out_payload_0_39_31_real = int_reg_array_39_31_real;
  assign io_coef_out_payload_0_39_31_imag = int_reg_array_39_31_imag;
  assign io_coef_out_payload_0_39_32_real = int_reg_array_39_32_real;
  assign io_coef_out_payload_0_39_32_imag = int_reg_array_39_32_imag;
  assign io_coef_out_payload_0_39_33_real = int_reg_array_39_33_real;
  assign io_coef_out_payload_0_39_33_imag = int_reg_array_39_33_imag;
  assign io_coef_out_payload_0_39_34_real = int_reg_array_39_34_real;
  assign io_coef_out_payload_0_39_34_imag = int_reg_array_39_34_imag;
  assign io_coef_out_payload_0_39_35_real = int_reg_array_39_35_real;
  assign io_coef_out_payload_0_39_35_imag = int_reg_array_39_35_imag;
  assign io_coef_out_payload_0_39_36_real = int_reg_array_39_36_real;
  assign io_coef_out_payload_0_39_36_imag = int_reg_array_39_36_imag;
  assign io_coef_out_payload_0_39_37_real = int_reg_array_39_37_real;
  assign io_coef_out_payload_0_39_37_imag = int_reg_array_39_37_imag;
  assign io_coef_out_payload_0_39_38_real = int_reg_array_39_38_real;
  assign io_coef_out_payload_0_39_38_imag = int_reg_array_39_38_imag;
  assign io_coef_out_payload_0_39_39_real = int_reg_array_39_39_real;
  assign io_coef_out_payload_0_39_39_imag = int_reg_array_39_39_imag;
  assign io_coef_out_payload_0_39_40_real = int_reg_array_39_40_real;
  assign io_coef_out_payload_0_39_40_imag = int_reg_array_39_40_imag;
  assign io_coef_out_payload_0_39_41_real = int_reg_array_39_41_real;
  assign io_coef_out_payload_0_39_41_imag = int_reg_array_39_41_imag;
  assign io_coef_out_payload_0_39_42_real = int_reg_array_39_42_real;
  assign io_coef_out_payload_0_39_42_imag = int_reg_array_39_42_imag;
  assign io_coef_out_payload_0_39_43_real = int_reg_array_39_43_real;
  assign io_coef_out_payload_0_39_43_imag = int_reg_array_39_43_imag;
  assign io_coef_out_payload_0_39_44_real = int_reg_array_39_44_real;
  assign io_coef_out_payload_0_39_44_imag = int_reg_array_39_44_imag;
  assign io_coef_out_payload_0_39_45_real = int_reg_array_39_45_real;
  assign io_coef_out_payload_0_39_45_imag = int_reg_array_39_45_imag;
  assign io_coef_out_payload_0_39_46_real = int_reg_array_39_46_real;
  assign io_coef_out_payload_0_39_46_imag = int_reg_array_39_46_imag;
  assign io_coef_out_payload_0_39_47_real = int_reg_array_39_47_real;
  assign io_coef_out_payload_0_39_47_imag = int_reg_array_39_47_imag;
  assign io_coef_out_payload_0_39_48_real = int_reg_array_39_48_real;
  assign io_coef_out_payload_0_39_48_imag = int_reg_array_39_48_imag;
  assign io_coef_out_payload_0_39_49_real = int_reg_array_39_49_real;
  assign io_coef_out_payload_0_39_49_imag = int_reg_array_39_49_imag;
  assign io_coef_out_payload_0_40_0_real = int_reg_array_40_0_real;
  assign io_coef_out_payload_0_40_0_imag = int_reg_array_40_0_imag;
  assign io_coef_out_payload_0_40_1_real = int_reg_array_40_1_real;
  assign io_coef_out_payload_0_40_1_imag = int_reg_array_40_1_imag;
  assign io_coef_out_payload_0_40_2_real = int_reg_array_40_2_real;
  assign io_coef_out_payload_0_40_2_imag = int_reg_array_40_2_imag;
  assign io_coef_out_payload_0_40_3_real = int_reg_array_40_3_real;
  assign io_coef_out_payload_0_40_3_imag = int_reg_array_40_3_imag;
  assign io_coef_out_payload_0_40_4_real = int_reg_array_40_4_real;
  assign io_coef_out_payload_0_40_4_imag = int_reg_array_40_4_imag;
  assign io_coef_out_payload_0_40_5_real = int_reg_array_40_5_real;
  assign io_coef_out_payload_0_40_5_imag = int_reg_array_40_5_imag;
  assign io_coef_out_payload_0_40_6_real = int_reg_array_40_6_real;
  assign io_coef_out_payload_0_40_6_imag = int_reg_array_40_6_imag;
  assign io_coef_out_payload_0_40_7_real = int_reg_array_40_7_real;
  assign io_coef_out_payload_0_40_7_imag = int_reg_array_40_7_imag;
  assign io_coef_out_payload_0_40_8_real = int_reg_array_40_8_real;
  assign io_coef_out_payload_0_40_8_imag = int_reg_array_40_8_imag;
  assign io_coef_out_payload_0_40_9_real = int_reg_array_40_9_real;
  assign io_coef_out_payload_0_40_9_imag = int_reg_array_40_9_imag;
  assign io_coef_out_payload_0_40_10_real = int_reg_array_40_10_real;
  assign io_coef_out_payload_0_40_10_imag = int_reg_array_40_10_imag;
  assign io_coef_out_payload_0_40_11_real = int_reg_array_40_11_real;
  assign io_coef_out_payload_0_40_11_imag = int_reg_array_40_11_imag;
  assign io_coef_out_payload_0_40_12_real = int_reg_array_40_12_real;
  assign io_coef_out_payload_0_40_12_imag = int_reg_array_40_12_imag;
  assign io_coef_out_payload_0_40_13_real = int_reg_array_40_13_real;
  assign io_coef_out_payload_0_40_13_imag = int_reg_array_40_13_imag;
  assign io_coef_out_payload_0_40_14_real = int_reg_array_40_14_real;
  assign io_coef_out_payload_0_40_14_imag = int_reg_array_40_14_imag;
  assign io_coef_out_payload_0_40_15_real = int_reg_array_40_15_real;
  assign io_coef_out_payload_0_40_15_imag = int_reg_array_40_15_imag;
  assign io_coef_out_payload_0_40_16_real = int_reg_array_40_16_real;
  assign io_coef_out_payload_0_40_16_imag = int_reg_array_40_16_imag;
  assign io_coef_out_payload_0_40_17_real = int_reg_array_40_17_real;
  assign io_coef_out_payload_0_40_17_imag = int_reg_array_40_17_imag;
  assign io_coef_out_payload_0_40_18_real = int_reg_array_40_18_real;
  assign io_coef_out_payload_0_40_18_imag = int_reg_array_40_18_imag;
  assign io_coef_out_payload_0_40_19_real = int_reg_array_40_19_real;
  assign io_coef_out_payload_0_40_19_imag = int_reg_array_40_19_imag;
  assign io_coef_out_payload_0_40_20_real = int_reg_array_40_20_real;
  assign io_coef_out_payload_0_40_20_imag = int_reg_array_40_20_imag;
  assign io_coef_out_payload_0_40_21_real = int_reg_array_40_21_real;
  assign io_coef_out_payload_0_40_21_imag = int_reg_array_40_21_imag;
  assign io_coef_out_payload_0_40_22_real = int_reg_array_40_22_real;
  assign io_coef_out_payload_0_40_22_imag = int_reg_array_40_22_imag;
  assign io_coef_out_payload_0_40_23_real = int_reg_array_40_23_real;
  assign io_coef_out_payload_0_40_23_imag = int_reg_array_40_23_imag;
  assign io_coef_out_payload_0_40_24_real = int_reg_array_40_24_real;
  assign io_coef_out_payload_0_40_24_imag = int_reg_array_40_24_imag;
  assign io_coef_out_payload_0_40_25_real = int_reg_array_40_25_real;
  assign io_coef_out_payload_0_40_25_imag = int_reg_array_40_25_imag;
  assign io_coef_out_payload_0_40_26_real = int_reg_array_40_26_real;
  assign io_coef_out_payload_0_40_26_imag = int_reg_array_40_26_imag;
  assign io_coef_out_payload_0_40_27_real = int_reg_array_40_27_real;
  assign io_coef_out_payload_0_40_27_imag = int_reg_array_40_27_imag;
  assign io_coef_out_payload_0_40_28_real = int_reg_array_40_28_real;
  assign io_coef_out_payload_0_40_28_imag = int_reg_array_40_28_imag;
  assign io_coef_out_payload_0_40_29_real = int_reg_array_40_29_real;
  assign io_coef_out_payload_0_40_29_imag = int_reg_array_40_29_imag;
  assign io_coef_out_payload_0_40_30_real = int_reg_array_40_30_real;
  assign io_coef_out_payload_0_40_30_imag = int_reg_array_40_30_imag;
  assign io_coef_out_payload_0_40_31_real = int_reg_array_40_31_real;
  assign io_coef_out_payload_0_40_31_imag = int_reg_array_40_31_imag;
  assign io_coef_out_payload_0_40_32_real = int_reg_array_40_32_real;
  assign io_coef_out_payload_0_40_32_imag = int_reg_array_40_32_imag;
  assign io_coef_out_payload_0_40_33_real = int_reg_array_40_33_real;
  assign io_coef_out_payload_0_40_33_imag = int_reg_array_40_33_imag;
  assign io_coef_out_payload_0_40_34_real = int_reg_array_40_34_real;
  assign io_coef_out_payload_0_40_34_imag = int_reg_array_40_34_imag;
  assign io_coef_out_payload_0_40_35_real = int_reg_array_40_35_real;
  assign io_coef_out_payload_0_40_35_imag = int_reg_array_40_35_imag;
  assign io_coef_out_payload_0_40_36_real = int_reg_array_40_36_real;
  assign io_coef_out_payload_0_40_36_imag = int_reg_array_40_36_imag;
  assign io_coef_out_payload_0_40_37_real = int_reg_array_40_37_real;
  assign io_coef_out_payload_0_40_37_imag = int_reg_array_40_37_imag;
  assign io_coef_out_payload_0_40_38_real = int_reg_array_40_38_real;
  assign io_coef_out_payload_0_40_38_imag = int_reg_array_40_38_imag;
  assign io_coef_out_payload_0_40_39_real = int_reg_array_40_39_real;
  assign io_coef_out_payload_0_40_39_imag = int_reg_array_40_39_imag;
  assign io_coef_out_payload_0_40_40_real = int_reg_array_40_40_real;
  assign io_coef_out_payload_0_40_40_imag = int_reg_array_40_40_imag;
  assign io_coef_out_payload_0_40_41_real = int_reg_array_40_41_real;
  assign io_coef_out_payload_0_40_41_imag = int_reg_array_40_41_imag;
  assign io_coef_out_payload_0_40_42_real = int_reg_array_40_42_real;
  assign io_coef_out_payload_0_40_42_imag = int_reg_array_40_42_imag;
  assign io_coef_out_payload_0_40_43_real = int_reg_array_40_43_real;
  assign io_coef_out_payload_0_40_43_imag = int_reg_array_40_43_imag;
  assign io_coef_out_payload_0_40_44_real = int_reg_array_40_44_real;
  assign io_coef_out_payload_0_40_44_imag = int_reg_array_40_44_imag;
  assign io_coef_out_payload_0_40_45_real = int_reg_array_40_45_real;
  assign io_coef_out_payload_0_40_45_imag = int_reg_array_40_45_imag;
  assign io_coef_out_payload_0_40_46_real = int_reg_array_40_46_real;
  assign io_coef_out_payload_0_40_46_imag = int_reg_array_40_46_imag;
  assign io_coef_out_payload_0_40_47_real = int_reg_array_40_47_real;
  assign io_coef_out_payload_0_40_47_imag = int_reg_array_40_47_imag;
  assign io_coef_out_payload_0_40_48_real = int_reg_array_40_48_real;
  assign io_coef_out_payload_0_40_48_imag = int_reg_array_40_48_imag;
  assign io_coef_out_payload_0_40_49_real = int_reg_array_40_49_real;
  assign io_coef_out_payload_0_40_49_imag = int_reg_array_40_49_imag;
  assign io_coef_out_payload_0_41_0_real = int_reg_array_41_0_real;
  assign io_coef_out_payload_0_41_0_imag = int_reg_array_41_0_imag;
  assign io_coef_out_payload_0_41_1_real = int_reg_array_41_1_real;
  assign io_coef_out_payload_0_41_1_imag = int_reg_array_41_1_imag;
  assign io_coef_out_payload_0_41_2_real = int_reg_array_41_2_real;
  assign io_coef_out_payload_0_41_2_imag = int_reg_array_41_2_imag;
  assign io_coef_out_payload_0_41_3_real = int_reg_array_41_3_real;
  assign io_coef_out_payload_0_41_3_imag = int_reg_array_41_3_imag;
  assign io_coef_out_payload_0_41_4_real = int_reg_array_41_4_real;
  assign io_coef_out_payload_0_41_4_imag = int_reg_array_41_4_imag;
  assign io_coef_out_payload_0_41_5_real = int_reg_array_41_5_real;
  assign io_coef_out_payload_0_41_5_imag = int_reg_array_41_5_imag;
  assign io_coef_out_payload_0_41_6_real = int_reg_array_41_6_real;
  assign io_coef_out_payload_0_41_6_imag = int_reg_array_41_6_imag;
  assign io_coef_out_payload_0_41_7_real = int_reg_array_41_7_real;
  assign io_coef_out_payload_0_41_7_imag = int_reg_array_41_7_imag;
  assign io_coef_out_payload_0_41_8_real = int_reg_array_41_8_real;
  assign io_coef_out_payload_0_41_8_imag = int_reg_array_41_8_imag;
  assign io_coef_out_payload_0_41_9_real = int_reg_array_41_9_real;
  assign io_coef_out_payload_0_41_9_imag = int_reg_array_41_9_imag;
  assign io_coef_out_payload_0_41_10_real = int_reg_array_41_10_real;
  assign io_coef_out_payload_0_41_10_imag = int_reg_array_41_10_imag;
  assign io_coef_out_payload_0_41_11_real = int_reg_array_41_11_real;
  assign io_coef_out_payload_0_41_11_imag = int_reg_array_41_11_imag;
  assign io_coef_out_payload_0_41_12_real = int_reg_array_41_12_real;
  assign io_coef_out_payload_0_41_12_imag = int_reg_array_41_12_imag;
  assign io_coef_out_payload_0_41_13_real = int_reg_array_41_13_real;
  assign io_coef_out_payload_0_41_13_imag = int_reg_array_41_13_imag;
  assign io_coef_out_payload_0_41_14_real = int_reg_array_41_14_real;
  assign io_coef_out_payload_0_41_14_imag = int_reg_array_41_14_imag;
  assign io_coef_out_payload_0_41_15_real = int_reg_array_41_15_real;
  assign io_coef_out_payload_0_41_15_imag = int_reg_array_41_15_imag;
  assign io_coef_out_payload_0_41_16_real = int_reg_array_41_16_real;
  assign io_coef_out_payload_0_41_16_imag = int_reg_array_41_16_imag;
  assign io_coef_out_payload_0_41_17_real = int_reg_array_41_17_real;
  assign io_coef_out_payload_0_41_17_imag = int_reg_array_41_17_imag;
  assign io_coef_out_payload_0_41_18_real = int_reg_array_41_18_real;
  assign io_coef_out_payload_0_41_18_imag = int_reg_array_41_18_imag;
  assign io_coef_out_payload_0_41_19_real = int_reg_array_41_19_real;
  assign io_coef_out_payload_0_41_19_imag = int_reg_array_41_19_imag;
  assign io_coef_out_payload_0_41_20_real = int_reg_array_41_20_real;
  assign io_coef_out_payload_0_41_20_imag = int_reg_array_41_20_imag;
  assign io_coef_out_payload_0_41_21_real = int_reg_array_41_21_real;
  assign io_coef_out_payload_0_41_21_imag = int_reg_array_41_21_imag;
  assign io_coef_out_payload_0_41_22_real = int_reg_array_41_22_real;
  assign io_coef_out_payload_0_41_22_imag = int_reg_array_41_22_imag;
  assign io_coef_out_payload_0_41_23_real = int_reg_array_41_23_real;
  assign io_coef_out_payload_0_41_23_imag = int_reg_array_41_23_imag;
  assign io_coef_out_payload_0_41_24_real = int_reg_array_41_24_real;
  assign io_coef_out_payload_0_41_24_imag = int_reg_array_41_24_imag;
  assign io_coef_out_payload_0_41_25_real = int_reg_array_41_25_real;
  assign io_coef_out_payload_0_41_25_imag = int_reg_array_41_25_imag;
  assign io_coef_out_payload_0_41_26_real = int_reg_array_41_26_real;
  assign io_coef_out_payload_0_41_26_imag = int_reg_array_41_26_imag;
  assign io_coef_out_payload_0_41_27_real = int_reg_array_41_27_real;
  assign io_coef_out_payload_0_41_27_imag = int_reg_array_41_27_imag;
  assign io_coef_out_payload_0_41_28_real = int_reg_array_41_28_real;
  assign io_coef_out_payload_0_41_28_imag = int_reg_array_41_28_imag;
  assign io_coef_out_payload_0_41_29_real = int_reg_array_41_29_real;
  assign io_coef_out_payload_0_41_29_imag = int_reg_array_41_29_imag;
  assign io_coef_out_payload_0_41_30_real = int_reg_array_41_30_real;
  assign io_coef_out_payload_0_41_30_imag = int_reg_array_41_30_imag;
  assign io_coef_out_payload_0_41_31_real = int_reg_array_41_31_real;
  assign io_coef_out_payload_0_41_31_imag = int_reg_array_41_31_imag;
  assign io_coef_out_payload_0_41_32_real = int_reg_array_41_32_real;
  assign io_coef_out_payload_0_41_32_imag = int_reg_array_41_32_imag;
  assign io_coef_out_payload_0_41_33_real = int_reg_array_41_33_real;
  assign io_coef_out_payload_0_41_33_imag = int_reg_array_41_33_imag;
  assign io_coef_out_payload_0_41_34_real = int_reg_array_41_34_real;
  assign io_coef_out_payload_0_41_34_imag = int_reg_array_41_34_imag;
  assign io_coef_out_payload_0_41_35_real = int_reg_array_41_35_real;
  assign io_coef_out_payload_0_41_35_imag = int_reg_array_41_35_imag;
  assign io_coef_out_payload_0_41_36_real = int_reg_array_41_36_real;
  assign io_coef_out_payload_0_41_36_imag = int_reg_array_41_36_imag;
  assign io_coef_out_payload_0_41_37_real = int_reg_array_41_37_real;
  assign io_coef_out_payload_0_41_37_imag = int_reg_array_41_37_imag;
  assign io_coef_out_payload_0_41_38_real = int_reg_array_41_38_real;
  assign io_coef_out_payload_0_41_38_imag = int_reg_array_41_38_imag;
  assign io_coef_out_payload_0_41_39_real = int_reg_array_41_39_real;
  assign io_coef_out_payload_0_41_39_imag = int_reg_array_41_39_imag;
  assign io_coef_out_payload_0_41_40_real = int_reg_array_41_40_real;
  assign io_coef_out_payload_0_41_40_imag = int_reg_array_41_40_imag;
  assign io_coef_out_payload_0_41_41_real = int_reg_array_41_41_real;
  assign io_coef_out_payload_0_41_41_imag = int_reg_array_41_41_imag;
  assign io_coef_out_payload_0_41_42_real = int_reg_array_41_42_real;
  assign io_coef_out_payload_0_41_42_imag = int_reg_array_41_42_imag;
  assign io_coef_out_payload_0_41_43_real = int_reg_array_41_43_real;
  assign io_coef_out_payload_0_41_43_imag = int_reg_array_41_43_imag;
  assign io_coef_out_payload_0_41_44_real = int_reg_array_41_44_real;
  assign io_coef_out_payload_0_41_44_imag = int_reg_array_41_44_imag;
  assign io_coef_out_payload_0_41_45_real = int_reg_array_41_45_real;
  assign io_coef_out_payload_0_41_45_imag = int_reg_array_41_45_imag;
  assign io_coef_out_payload_0_41_46_real = int_reg_array_41_46_real;
  assign io_coef_out_payload_0_41_46_imag = int_reg_array_41_46_imag;
  assign io_coef_out_payload_0_41_47_real = int_reg_array_41_47_real;
  assign io_coef_out_payload_0_41_47_imag = int_reg_array_41_47_imag;
  assign io_coef_out_payload_0_41_48_real = int_reg_array_41_48_real;
  assign io_coef_out_payload_0_41_48_imag = int_reg_array_41_48_imag;
  assign io_coef_out_payload_0_41_49_real = int_reg_array_41_49_real;
  assign io_coef_out_payload_0_41_49_imag = int_reg_array_41_49_imag;
  assign io_coef_out_payload_0_42_0_real = int_reg_array_42_0_real;
  assign io_coef_out_payload_0_42_0_imag = int_reg_array_42_0_imag;
  assign io_coef_out_payload_0_42_1_real = int_reg_array_42_1_real;
  assign io_coef_out_payload_0_42_1_imag = int_reg_array_42_1_imag;
  assign io_coef_out_payload_0_42_2_real = int_reg_array_42_2_real;
  assign io_coef_out_payload_0_42_2_imag = int_reg_array_42_2_imag;
  assign io_coef_out_payload_0_42_3_real = int_reg_array_42_3_real;
  assign io_coef_out_payload_0_42_3_imag = int_reg_array_42_3_imag;
  assign io_coef_out_payload_0_42_4_real = int_reg_array_42_4_real;
  assign io_coef_out_payload_0_42_4_imag = int_reg_array_42_4_imag;
  assign io_coef_out_payload_0_42_5_real = int_reg_array_42_5_real;
  assign io_coef_out_payload_0_42_5_imag = int_reg_array_42_5_imag;
  assign io_coef_out_payload_0_42_6_real = int_reg_array_42_6_real;
  assign io_coef_out_payload_0_42_6_imag = int_reg_array_42_6_imag;
  assign io_coef_out_payload_0_42_7_real = int_reg_array_42_7_real;
  assign io_coef_out_payload_0_42_7_imag = int_reg_array_42_7_imag;
  assign io_coef_out_payload_0_42_8_real = int_reg_array_42_8_real;
  assign io_coef_out_payload_0_42_8_imag = int_reg_array_42_8_imag;
  assign io_coef_out_payload_0_42_9_real = int_reg_array_42_9_real;
  assign io_coef_out_payload_0_42_9_imag = int_reg_array_42_9_imag;
  assign io_coef_out_payload_0_42_10_real = int_reg_array_42_10_real;
  assign io_coef_out_payload_0_42_10_imag = int_reg_array_42_10_imag;
  assign io_coef_out_payload_0_42_11_real = int_reg_array_42_11_real;
  assign io_coef_out_payload_0_42_11_imag = int_reg_array_42_11_imag;
  assign io_coef_out_payload_0_42_12_real = int_reg_array_42_12_real;
  assign io_coef_out_payload_0_42_12_imag = int_reg_array_42_12_imag;
  assign io_coef_out_payload_0_42_13_real = int_reg_array_42_13_real;
  assign io_coef_out_payload_0_42_13_imag = int_reg_array_42_13_imag;
  assign io_coef_out_payload_0_42_14_real = int_reg_array_42_14_real;
  assign io_coef_out_payload_0_42_14_imag = int_reg_array_42_14_imag;
  assign io_coef_out_payload_0_42_15_real = int_reg_array_42_15_real;
  assign io_coef_out_payload_0_42_15_imag = int_reg_array_42_15_imag;
  assign io_coef_out_payload_0_42_16_real = int_reg_array_42_16_real;
  assign io_coef_out_payload_0_42_16_imag = int_reg_array_42_16_imag;
  assign io_coef_out_payload_0_42_17_real = int_reg_array_42_17_real;
  assign io_coef_out_payload_0_42_17_imag = int_reg_array_42_17_imag;
  assign io_coef_out_payload_0_42_18_real = int_reg_array_42_18_real;
  assign io_coef_out_payload_0_42_18_imag = int_reg_array_42_18_imag;
  assign io_coef_out_payload_0_42_19_real = int_reg_array_42_19_real;
  assign io_coef_out_payload_0_42_19_imag = int_reg_array_42_19_imag;
  assign io_coef_out_payload_0_42_20_real = int_reg_array_42_20_real;
  assign io_coef_out_payload_0_42_20_imag = int_reg_array_42_20_imag;
  assign io_coef_out_payload_0_42_21_real = int_reg_array_42_21_real;
  assign io_coef_out_payload_0_42_21_imag = int_reg_array_42_21_imag;
  assign io_coef_out_payload_0_42_22_real = int_reg_array_42_22_real;
  assign io_coef_out_payload_0_42_22_imag = int_reg_array_42_22_imag;
  assign io_coef_out_payload_0_42_23_real = int_reg_array_42_23_real;
  assign io_coef_out_payload_0_42_23_imag = int_reg_array_42_23_imag;
  assign io_coef_out_payload_0_42_24_real = int_reg_array_42_24_real;
  assign io_coef_out_payload_0_42_24_imag = int_reg_array_42_24_imag;
  assign io_coef_out_payload_0_42_25_real = int_reg_array_42_25_real;
  assign io_coef_out_payload_0_42_25_imag = int_reg_array_42_25_imag;
  assign io_coef_out_payload_0_42_26_real = int_reg_array_42_26_real;
  assign io_coef_out_payload_0_42_26_imag = int_reg_array_42_26_imag;
  assign io_coef_out_payload_0_42_27_real = int_reg_array_42_27_real;
  assign io_coef_out_payload_0_42_27_imag = int_reg_array_42_27_imag;
  assign io_coef_out_payload_0_42_28_real = int_reg_array_42_28_real;
  assign io_coef_out_payload_0_42_28_imag = int_reg_array_42_28_imag;
  assign io_coef_out_payload_0_42_29_real = int_reg_array_42_29_real;
  assign io_coef_out_payload_0_42_29_imag = int_reg_array_42_29_imag;
  assign io_coef_out_payload_0_42_30_real = int_reg_array_42_30_real;
  assign io_coef_out_payload_0_42_30_imag = int_reg_array_42_30_imag;
  assign io_coef_out_payload_0_42_31_real = int_reg_array_42_31_real;
  assign io_coef_out_payload_0_42_31_imag = int_reg_array_42_31_imag;
  assign io_coef_out_payload_0_42_32_real = int_reg_array_42_32_real;
  assign io_coef_out_payload_0_42_32_imag = int_reg_array_42_32_imag;
  assign io_coef_out_payload_0_42_33_real = int_reg_array_42_33_real;
  assign io_coef_out_payload_0_42_33_imag = int_reg_array_42_33_imag;
  assign io_coef_out_payload_0_42_34_real = int_reg_array_42_34_real;
  assign io_coef_out_payload_0_42_34_imag = int_reg_array_42_34_imag;
  assign io_coef_out_payload_0_42_35_real = int_reg_array_42_35_real;
  assign io_coef_out_payload_0_42_35_imag = int_reg_array_42_35_imag;
  assign io_coef_out_payload_0_42_36_real = int_reg_array_42_36_real;
  assign io_coef_out_payload_0_42_36_imag = int_reg_array_42_36_imag;
  assign io_coef_out_payload_0_42_37_real = int_reg_array_42_37_real;
  assign io_coef_out_payload_0_42_37_imag = int_reg_array_42_37_imag;
  assign io_coef_out_payload_0_42_38_real = int_reg_array_42_38_real;
  assign io_coef_out_payload_0_42_38_imag = int_reg_array_42_38_imag;
  assign io_coef_out_payload_0_42_39_real = int_reg_array_42_39_real;
  assign io_coef_out_payload_0_42_39_imag = int_reg_array_42_39_imag;
  assign io_coef_out_payload_0_42_40_real = int_reg_array_42_40_real;
  assign io_coef_out_payload_0_42_40_imag = int_reg_array_42_40_imag;
  assign io_coef_out_payload_0_42_41_real = int_reg_array_42_41_real;
  assign io_coef_out_payload_0_42_41_imag = int_reg_array_42_41_imag;
  assign io_coef_out_payload_0_42_42_real = int_reg_array_42_42_real;
  assign io_coef_out_payload_0_42_42_imag = int_reg_array_42_42_imag;
  assign io_coef_out_payload_0_42_43_real = int_reg_array_42_43_real;
  assign io_coef_out_payload_0_42_43_imag = int_reg_array_42_43_imag;
  assign io_coef_out_payload_0_42_44_real = int_reg_array_42_44_real;
  assign io_coef_out_payload_0_42_44_imag = int_reg_array_42_44_imag;
  assign io_coef_out_payload_0_42_45_real = int_reg_array_42_45_real;
  assign io_coef_out_payload_0_42_45_imag = int_reg_array_42_45_imag;
  assign io_coef_out_payload_0_42_46_real = int_reg_array_42_46_real;
  assign io_coef_out_payload_0_42_46_imag = int_reg_array_42_46_imag;
  assign io_coef_out_payload_0_42_47_real = int_reg_array_42_47_real;
  assign io_coef_out_payload_0_42_47_imag = int_reg_array_42_47_imag;
  assign io_coef_out_payload_0_42_48_real = int_reg_array_42_48_real;
  assign io_coef_out_payload_0_42_48_imag = int_reg_array_42_48_imag;
  assign io_coef_out_payload_0_42_49_real = int_reg_array_42_49_real;
  assign io_coef_out_payload_0_42_49_imag = int_reg_array_42_49_imag;
  assign io_coef_out_payload_0_43_0_real = int_reg_array_43_0_real;
  assign io_coef_out_payload_0_43_0_imag = int_reg_array_43_0_imag;
  assign io_coef_out_payload_0_43_1_real = int_reg_array_43_1_real;
  assign io_coef_out_payload_0_43_1_imag = int_reg_array_43_1_imag;
  assign io_coef_out_payload_0_43_2_real = int_reg_array_43_2_real;
  assign io_coef_out_payload_0_43_2_imag = int_reg_array_43_2_imag;
  assign io_coef_out_payload_0_43_3_real = int_reg_array_43_3_real;
  assign io_coef_out_payload_0_43_3_imag = int_reg_array_43_3_imag;
  assign io_coef_out_payload_0_43_4_real = int_reg_array_43_4_real;
  assign io_coef_out_payload_0_43_4_imag = int_reg_array_43_4_imag;
  assign io_coef_out_payload_0_43_5_real = int_reg_array_43_5_real;
  assign io_coef_out_payload_0_43_5_imag = int_reg_array_43_5_imag;
  assign io_coef_out_payload_0_43_6_real = int_reg_array_43_6_real;
  assign io_coef_out_payload_0_43_6_imag = int_reg_array_43_6_imag;
  assign io_coef_out_payload_0_43_7_real = int_reg_array_43_7_real;
  assign io_coef_out_payload_0_43_7_imag = int_reg_array_43_7_imag;
  assign io_coef_out_payload_0_43_8_real = int_reg_array_43_8_real;
  assign io_coef_out_payload_0_43_8_imag = int_reg_array_43_8_imag;
  assign io_coef_out_payload_0_43_9_real = int_reg_array_43_9_real;
  assign io_coef_out_payload_0_43_9_imag = int_reg_array_43_9_imag;
  assign io_coef_out_payload_0_43_10_real = int_reg_array_43_10_real;
  assign io_coef_out_payload_0_43_10_imag = int_reg_array_43_10_imag;
  assign io_coef_out_payload_0_43_11_real = int_reg_array_43_11_real;
  assign io_coef_out_payload_0_43_11_imag = int_reg_array_43_11_imag;
  assign io_coef_out_payload_0_43_12_real = int_reg_array_43_12_real;
  assign io_coef_out_payload_0_43_12_imag = int_reg_array_43_12_imag;
  assign io_coef_out_payload_0_43_13_real = int_reg_array_43_13_real;
  assign io_coef_out_payload_0_43_13_imag = int_reg_array_43_13_imag;
  assign io_coef_out_payload_0_43_14_real = int_reg_array_43_14_real;
  assign io_coef_out_payload_0_43_14_imag = int_reg_array_43_14_imag;
  assign io_coef_out_payload_0_43_15_real = int_reg_array_43_15_real;
  assign io_coef_out_payload_0_43_15_imag = int_reg_array_43_15_imag;
  assign io_coef_out_payload_0_43_16_real = int_reg_array_43_16_real;
  assign io_coef_out_payload_0_43_16_imag = int_reg_array_43_16_imag;
  assign io_coef_out_payload_0_43_17_real = int_reg_array_43_17_real;
  assign io_coef_out_payload_0_43_17_imag = int_reg_array_43_17_imag;
  assign io_coef_out_payload_0_43_18_real = int_reg_array_43_18_real;
  assign io_coef_out_payload_0_43_18_imag = int_reg_array_43_18_imag;
  assign io_coef_out_payload_0_43_19_real = int_reg_array_43_19_real;
  assign io_coef_out_payload_0_43_19_imag = int_reg_array_43_19_imag;
  assign io_coef_out_payload_0_43_20_real = int_reg_array_43_20_real;
  assign io_coef_out_payload_0_43_20_imag = int_reg_array_43_20_imag;
  assign io_coef_out_payload_0_43_21_real = int_reg_array_43_21_real;
  assign io_coef_out_payload_0_43_21_imag = int_reg_array_43_21_imag;
  assign io_coef_out_payload_0_43_22_real = int_reg_array_43_22_real;
  assign io_coef_out_payload_0_43_22_imag = int_reg_array_43_22_imag;
  assign io_coef_out_payload_0_43_23_real = int_reg_array_43_23_real;
  assign io_coef_out_payload_0_43_23_imag = int_reg_array_43_23_imag;
  assign io_coef_out_payload_0_43_24_real = int_reg_array_43_24_real;
  assign io_coef_out_payload_0_43_24_imag = int_reg_array_43_24_imag;
  assign io_coef_out_payload_0_43_25_real = int_reg_array_43_25_real;
  assign io_coef_out_payload_0_43_25_imag = int_reg_array_43_25_imag;
  assign io_coef_out_payload_0_43_26_real = int_reg_array_43_26_real;
  assign io_coef_out_payload_0_43_26_imag = int_reg_array_43_26_imag;
  assign io_coef_out_payload_0_43_27_real = int_reg_array_43_27_real;
  assign io_coef_out_payload_0_43_27_imag = int_reg_array_43_27_imag;
  assign io_coef_out_payload_0_43_28_real = int_reg_array_43_28_real;
  assign io_coef_out_payload_0_43_28_imag = int_reg_array_43_28_imag;
  assign io_coef_out_payload_0_43_29_real = int_reg_array_43_29_real;
  assign io_coef_out_payload_0_43_29_imag = int_reg_array_43_29_imag;
  assign io_coef_out_payload_0_43_30_real = int_reg_array_43_30_real;
  assign io_coef_out_payload_0_43_30_imag = int_reg_array_43_30_imag;
  assign io_coef_out_payload_0_43_31_real = int_reg_array_43_31_real;
  assign io_coef_out_payload_0_43_31_imag = int_reg_array_43_31_imag;
  assign io_coef_out_payload_0_43_32_real = int_reg_array_43_32_real;
  assign io_coef_out_payload_0_43_32_imag = int_reg_array_43_32_imag;
  assign io_coef_out_payload_0_43_33_real = int_reg_array_43_33_real;
  assign io_coef_out_payload_0_43_33_imag = int_reg_array_43_33_imag;
  assign io_coef_out_payload_0_43_34_real = int_reg_array_43_34_real;
  assign io_coef_out_payload_0_43_34_imag = int_reg_array_43_34_imag;
  assign io_coef_out_payload_0_43_35_real = int_reg_array_43_35_real;
  assign io_coef_out_payload_0_43_35_imag = int_reg_array_43_35_imag;
  assign io_coef_out_payload_0_43_36_real = int_reg_array_43_36_real;
  assign io_coef_out_payload_0_43_36_imag = int_reg_array_43_36_imag;
  assign io_coef_out_payload_0_43_37_real = int_reg_array_43_37_real;
  assign io_coef_out_payload_0_43_37_imag = int_reg_array_43_37_imag;
  assign io_coef_out_payload_0_43_38_real = int_reg_array_43_38_real;
  assign io_coef_out_payload_0_43_38_imag = int_reg_array_43_38_imag;
  assign io_coef_out_payload_0_43_39_real = int_reg_array_43_39_real;
  assign io_coef_out_payload_0_43_39_imag = int_reg_array_43_39_imag;
  assign io_coef_out_payload_0_43_40_real = int_reg_array_43_40_real;
  assign io_coef_out_payload_0_43_40_imag = int_reg_array_43_40_imag;
  assign io_coef_out_payload_0_43_41_real = int_reg_array_43_41_real;
  assign io_coef_out_payload_0_43_41_imag = int_reg_array_43_41_imag;
  assign io_coef_out_payload_0_43_42_real = int_reg_array_43_42_real;
  assign io_coef_out_payload_0_43_42_imag = int_reg_array_43_42_imag;
  assign io_coef_out_payload_0_43_43_real = int_reg_array_43_43_real;
  assign io_coef_out_payload_0_43_43_imag = int_reg_array_43_43_imag;
  assign io_coef_out_payload_0_43_44_real = int_reg_array_43_44_real;
  assign io_coef_out_payload_0_43_44_imag = int_reg_array_43_44_imag;
  assign io_coef_out_payload_0_43_45_real = int_reg_array_43_45_real;
  assign io_coef_out_payload_0_43_45_imag = int_reg_array_43_45_imag;
  assign io_coef_out_payload_0_43_46_real = int_reg_array_43_46_real;
  assign io_coef_out_payload_0_43_46_imag = int_reg_array_43_46_imag;
  assign io_coef_out_payload_0_43_47_real = int_reg_array_43_47_real;
  assign io_coef_out_payload_0_43_47_imag = int_reg_array_43_47_imag;
  assign io_coef_out_payload_0_43_48_real = int_reg_array_43_48_real;
  assign io_coef_out_payload_0_43_48_imag = int_reg_array_43_48_imag;
  assign io_coef_out_payload_0_43_49_real = int_reg_array_43_49_real;
  assign io_coef_out_payload_0_43_49_imag = int_reg_array_43_49_imag;
  assign io_coef_out_payload_0_44_0_real = int_reg_array_44_0_real;
  assign io_coef_out_payload_0_44_0_imag = int_reg_array_44_0_imag;
  assign io_coef_out_payload_0_44_1_real = int_reg_array_44_1_real;
  assign io_coef_out_payload_0_44_1_imag = int_reg_array_44_1_imag;
  assign io_coef_out_payload_0_44_2_real = int_reg_array_44_2_real;
  assign io_coef_out_payload_0_44_2_imag = int_reg_array_44_2_imag;
  assign io_coef_out_payload_0_44_3_real = int_reg_array_44_3_real;
  assign io_coef_out_payload_0_44_3_imag = int_reg_array_44_3_imag;
  assign io_coef_out_payload_0_44_4_real = int_reg_array_44_4_real;
  assign io_coef_out_payload_0_44_4_imag = int_reg_array_44_4_imag;
  assign io_coef_out_payload_0_44_5_real = int_reg_array_44_5_real;
  assign io_coef_out_payload_0_44_5_imag = int_reg_array_44_5_imag;
  assign io_coef_out_payload_0_44_6_real = int_reg_array_44_6_real;
  assign io_coef_out_payload_0_44_6_imag = int_reg_array_44_6_imag;
  assign io_coef_out_payload_0_44_7_real = int_reg_array_44_7_real;
  assign io_coef_out_payload_0_44_7_imag = int_reg_array_44_7_imag;
  assign io_coef_out_payload_0_44_8_real = int_reg_array_44_8_real;
  assign io_coef_out_payload_0_44_8_imag = int_reg_array_44_8_imag;
  assign io_coef_out_payload_0_44_9_real = int_reg_array_44_9_real;
  assign io_coef_out_payload_0_44_9_imag = int_reg_array_44_9_imag;
  assign io_coef_out_payload_0_44_10_real = int_reg_array_44_10_real;
  assign io_coef_out_payload_0_44_10_imag = int_reg_array_44_10_imag;
  assign io_coef_out_payload_0_44_11_real = int_reg_array_44_11_real;
  assign io_coef_out_payload_0_44_11_imag = int_reg_array_44_11_imag;
  assign io_coef_out_payload_0_44_12_real = int_reg_array_44_12_real;
  assign io_coef_out_payload_0_44_12_imag = int_reg_array_44_12_imag;
  assign io_coef_out_payload_0_44_13_real = int_reg_array_44_13_real;
  assign io_coef_out_payload_0_44_13_imag = int_reg_array_44_13_imag;
  assign io_coef_out_payload_0_44_14_real = int_reg_array_44_14_real;
  assign io_coef_out_payload_0_44_14_imag = int_reg_array_44_14_imag;
  assign io_coef_out_payload_0_44_15_real = int_reg_array_44_15_real;
  assign io_coef_out_payload_0_44_15_imag = int_reg_array_44_15_imag;
  assign io_coef_out_payload_0_44_16_real = int_reg_array_44_16_real;
  assign io_coef_out_payload_0_44_16_imag = int_reg_array_44_16_imag;
  assign io_coef_out_payload_0_44_17_real = int_reg_array_44_17_real;
  assign io_coef_out_payload_0_44_17_imag = int_reg_array_44_17_imag;
  assign io_coef_out_payload_0_44_18_real = int_reg_array_44_18_real;
  assign io_coef_out_payload_0_44_18_imag = int_reg_array_44_18_imag;
  assign io_coef_out_payload_0_44_19_real = int_reg_array_44_19_real;
  assign io_coef_out_payload_0_44_19_imag = int_reg_array_44_19_imag;
  assign io_coef_out_payload_0_44_20_real = int_reg_array_44_20_real;
  assign io_coef_out_payload_0_44_20_imag = int_reg_array_44_20_imag;
  assign io_coef_out_payload_0_44_21_real = int_reg_array_44_21_real;
  assign io_coef_out_payload_0_44_21_imag = int_reg_array_44_21_imag;
  assign io_coef_out_payload_0_44_22_real = int_reg_array_44_22_real;
  assign io_coef_out_payload_0_44_22_imag = int_reg_array_44_22_imag;
  assign io_coef_out_payload_0_44_23_real = int_reg_array_44_23_real;
  assign io_coef_out_payload_0_44_23_imag = int_reg_array_44_23_imag;
  assign io_coef_out_payload_0_44_24_real = int_reg_array_44_24_real;
  assign io_coef_out_payload_0_44_24_imag = int_reg_array_44_24_imag;
  assign io_coef_out_payload_0_44_25_real = int_reg_array_44_25_real;
  assign io_coef_out_payload_0_44_25_imag = int_reg_array_44_25_imag;
  assign io_coef_out_payload_0_44_26_real = int_reg_array_44_26_real;
  assign io_coef_out_payload_0_44_26_imag = int_reg_array_44_26_imag;
  assign io_coef_out_payload_0_44_27_real = int_reg_array_44_27_real;
  assign io_coef_out_payload_0_44_27_imag = int_reg_array_44_27_imag;
  assign io_coef_out_payload_0_44_28_real = int_reg_array_44_28_real;
  assign io_coef_out_payload_0_44_28_imag = int_reg_array_44_28_imag;
  assign io_coef_out_payload_0_44_29_real = int_reg_array_44_29_real;
  assign io_coef_out_payload_0_44_29_imag = int_reg_array_44_29_imag;
  assign io_coef_out_payload_0_44_30_real = int_reg_array_44_30_real;
  assign io_coef_out_payload_0_44_30_imag = int_reg_array_44_30_imag;
  assign io_coef_out_payload_0_44_31_real = int_reg_array_44_31_real;
  assign io_coef_out_payload_0_44_31_imag = int_reg_array_44_31_imag;
  assign io_coef_out_payload_0_44_32_real = int_reg_array_44_32_real;
  assign io_coef_out_payload_0_44_32_imag = int_reg_array_44_32_imag;
  assign io_coef_out_payload_0_44_33_real = int_reg_array_44_33_real;
  assign io_coef_out_payload_0_44_33_imag = int_reg_array_44_33_imag;
  assign io_coef_out_payload_0_44_34_real = int_reg_array_44_34_real;
  assign io_coef_out_payload_0_44_34_imag = int_reg_array_44_34_imag;
  assign io_coef_out_payload_0_44_35_real = int_reg_array_44_35_real;
  assign io_coef_out_payload_0_44_35_imag = int_reg_array_44_35_imag;
  assign io_coef_out_payload_0_44_36_real = int_reg_array_44_36_real;
  assign io_coef_out_payload_0_44_36_imag = int_reg_array_44_36_imag;
  assign io_coef_out_payload_0_44_37_real = int_reg_array_44_37_real;
  assign io_coef_out_payload_0_44_37_imag = int_reg_array_44_37_imag;
  assign io_coef_out_payload_0_44_38_real = int_reg_array_44_38_real;
  assign io_coef_out_payload_0_44_38_imag = int_reg_array_44_38_imag;
  assign io_coef_out_payload_0_44_39_real = int_reg_array_44_39_real;
  assign io_coef_out_payload_0_44_39_imag = int_reg_array_44_39_imag;
  assign io_coef_out_payload_0_44_40_real = int_reg_array_44_40_real;
  assign io_coef_out_payload_0_44_40_imag = int_reg_array_44_40_imag;
  assign io_coef_out_payload_0_44_41_real = int_reg_array_44_41_real;
  assign io_coef_out_payload_0_44_41_imag = int_reg_array_44_41_imag;
  assign io_coef_out_payload_0_44_42_real = int_reg_array_44_42_real;
  assign io_coef_out_payload_0_44_42_imag = int_reg_array_44_42_imag;
  assign io_coef_out_payload_0_44_43_real = int_reg_array_44_43_real;
  assign io_coef_out_payload_0_44_43_imag = int_reg_array_44_43_imag;
  assign io_coef_out_payload_0_44_44_real = int_reg_array_44_44_real;
  assign io_coef_out_payload_0_44_44_imag = int_reg_array_44_44_imag;
  assign io_coef_out_payload_0_44_45_real = int_reg_array_44_45_real;
  assign io_coef_out_payload_0_44_45_imag = int_reg_array_44_45_imag;
  assign io_coef_out_payload_0_44_46_real = int_reg_array_44_46_real;
  assign io_coef_out_payload_0_44_46_imag = int_reg_array_44_46_imag;
  assign io_coef_out_payload_0_44_47_real = int_reg_array_44_47_real;
  assign io_coef_out_payload_0_44_47_imag = int_reg_array_44_47_imag;
  assign io_coef_out_payload_0_44_48_real = int_reg_array_44_48_real;
  assign io_coef_out_payload_0_44_48_imag = int_reg_array_44_48_imag;
  assign io_coef_out_payload_0_44_49_real = int_reg_array_44_49_real;
  assign io_coef_out_payload_0_44_49_imag = int_reg_array_44_49_imag;
  assign io_coef_out_payload_0_45_0_real = int_reg_array_45_0_real;
  assign io_coef_out_payload_0_45_0_imag = int_reg_array_45_0_imag;
  assign io_coef_out_payload_0_45_1_real = int_reg_array_45_1_real;
  assign io_coef_out_payload_0_45_1_imag = int_reg_array_45_1_imag;
  assign io_coef_out_payload_0_45_2_real = int_reg_array_45_2_real;
  assign io_coef_out_payload_0_45_2_imag = int_reg_array_45_2_imag;
  assign io_coef_out_payload_0_45_3_real = int_reg_array_45_3_real;
  assign io_coef_out_payload_0_45_3_imag = int_reg_array_45_3_imag;
  assign io_coef_out_payload_0_45_4_real = int_reg_array_45_4_real;
  assign io_coef_out_payload_0_45_4_imag = int_reg_array_45_4_imag;
  assign io_coef_out_payload_0_45_5_real = int_reg_array_45_5_real;
  assign io_coef_out_payload_0_45_5_imag = int_reg_array_45_5_imag;
  assign io_coef_out_payload_0_45_6_real = int_reg_array_45_6_real;
  assign io_coef_out_payload_0_45_6_imag = int_reg_array_45_6_imag;
  assign io_coef_out_payload_0_45_7_real = int_reg_array_45_7_real;
  assign io_coef_out_payload_0_45_7_imag = int_reg_array_45_7_imag;
  assign io_coef_out_payload_0_45_8_real = int_reg_array_45_8_real;
  assign io_coef_out_payload_0_45_8_imag = int_reg_array_45_8_imag;
  assign io_coef_out_payload_0_45_9_real = int_reg_array_45_9_real;
  assign io_coef_out_payload_0_45_9_imag = int_reg_array_45_9_imag;
  assign io_coef_out_payload_0_45_10_real = int_reg_array_45_10_real;
  assign io_coef_out_payload_0_45_10_imag = int_reg_array_45_10_imag;
  assign io_coef_out_payload_0_45_11_real = int_reg_array_45_11_real;
  assign io_coef_out_payload_0_45_11_imag = int_reg_array_45_11_imag;
  assign io_coef_out_payload_0_45_12_real = int_reg_array_45_12_real;
  assign io_coef_out_payload_0_45_12_imag = int_reg_array_45_12_imag;
  assign io_coef_out_payload_0_45_13_real = int_reg_array_45_13_real;
  assign io_coef_out_payload_0_45_13_imag = int_reg_array_45_13_imag;
  assign io_coef_out_payload_0_45_14_real = int_reg_array_45_14_real;
  assign io_coef_out_payload_0_45_14_imag = int_reg_array_45_14_imag;
  assign io_coef_out_payload_0_45_15_real = int_reg_array_45_15_real;
  assign io_coef_out_payload_0_45_15_imag = int_reg_array_45_15_imag;
  assign io_coef_out_payload_0_45_16_real = int_reg_array_45_16_real;
  assign io_coef_out_payload_0_45_16_imag = int_reg_array_45_16_imag;
  assign io_coef_out_payload_0_45_17_real = int_reg_array_45_17_real;
  assign io_coef_out_payload_0_45_17_imag = int_reg_array_45_17_imag;
  assign io_coef_out_payload_0_45_18_real = int_reg_array_45_18_real;
  assign io_coef_out_payload_0_45_18_imag = int_reg_array_45_18_imag;
  assign io_coef_out_payload_0_45_19_real = int_reg_array_45_19_real;
  assign io_coef_out_payload_0_45_19_imag = int_reg_array_45_19_imag;
  assign io_coef_out_payload_0_45_20_real = int_reg_array_45_20_real;
  assign io_coef_out_payload_0_45_20_imag = int_reg_array_45_20_imag;
  assign io_coef_out_payload_0_45_21_real = int_reg_array_45_21_real;
  assign io_coef_out_payload_0_45_21_imag = int_reg_array_45_21_imag;
  assign io_coef_out_payload_0_45_22_real = int_reg_array_45_22_real;
  assign io_coef_out_payload_0_45_22_imag = int_reg_array_45_22_imag;
  assign io_coef_out_payload_0_45_23_real = int_reg_array_45_23_real;
  assign io_coef_out_payload_0_45_23_imag = int_reg_array_45_23_imag;
  assign io_coef_out_payload_0_45_24_real = int_reg_array_45_24_real;
  assign io_coef_out_payload_0_45_24_imag = int_reg_array_45_24_imag;
  assign io_coef_out_payload_0_45_25_real = int_reg_array_45_25_real;
  assign io_coef_out_payload_0_45_25_imag = int_reg_array_45_25_imag;
  assign io_coef_out_payload_0_45_26_real = int_reg_array_45_26_real;
  assign io_coef_out_payload_0_45_26_imag = int_reg_array_45_26_imag;
  assign io_coef_out_payload_0_45_27_real = int_reg_array_45_27_real;
  assign io_coef_out_payload_0_45_27_imag = int_reg_array_45_27_imag;
  assign io_coef_out_payload_0_45_28_real = int_reg_array_45_28_real;
  assign io_coef_out_payload_0_45_28_imag = int_reg_array_45_28_imag;
  assign io_coef_out_payload_0_45_29_real = int_reg_array_45_29_real;
  assign io_coef_out_payload_0_45_29_imag = int_reg_array_45_29_imag;
  assign io_coef_out_payload_0_45_30_real = int_reg_array_45_30_real;
  assign io_coef_out_payload_0_45_30_imag = int_reg_array_45_30_imag;
  assign io_coef_out_payload_0_45_31_real = int_reg_array_45_31_real;
  assign io_coef_out_payload_0_45_31_imag = int_reg_array_45_31_imag;
  assign io_coef_out_payload_0_45_32_real = int_reg_array_45_32_real;
  assign io_coef_out_payload_0_45_32_imag = int_reg_array_45_32_imag;
  assign io_coef_out_payload_0_45_33_real = int_reg_array_45_33_real;
  assign io_coef_out_payload_0_45_33_imag = int_reg_array_45_33_imag;
  assign io_coef_out_payload_0_45_34_real = int_reg_array_45_34_real;
  assign io_coef_out_payload_0_45_34_imag = int_reg_array_45_34_imag;
  assign io_coef_out_payload_0_45_35_real = int_reg_array_45_35_real;
  assign io_coef_out_payload_0_45_35_imag = int_reg_array_45_35_imag;
  assign io_coef_out_payload_0_45_36_real = int_reg_array_45_36_real;
  assign io_coef_out_payload_0_45_36_imag = int_reg_array_45_36_imag;
  assign io_coef_out_payload_0_45_37_real = int_reg_array_45_37_real;
  assign io_coef_out_payload_0_45_37_imag = int_reg_array_45_37_imag;
  assign io_coef_out_payload_0_45_38_real = int_reg_array_45_38_real;
  assign io_coef_out_payload_0_45_38_imag = int_reg_array_45_38_imag;
  assign io_coef_out_payload_0_45_39_real = int_reg_array_45_39_real;
  assign io_coef_out_payload_0_45_39_imag = int_reg_array_45_39_imag;
  assign io_coef_out_payload_0_45_40_real = int_reg_array_45_40_real;
  assign io_coef_out_payload_0_45_40_imag = int_reg_array_45_40_imag;
  assign io_coef_out_payload_0_45_41_real = int_reg_array_45_41_real;
  assign io_coef_out_payload_0_45_41_imag = int_reg_array_45_41_imag;
  assign io_coef_out_payload_0_45_42_real = int_reg_array_45_42_real;
  assign io_coef_out_payload_0_45_42_imag = int_reg_array_45_42_imag;
  assign io_coef_out_payload_0_45_43_real = int_reg_array_45_43_real;
  assign io_coef_out_payload_0_45_43_imag = int_reg_array_45_43_imag;
  assign io_coef_out_payload_0_45_44_real = int_reg_array_45_44_real;
  assign io_coef_out_payload_0_45_44_imag = int_reg_array_45_44_imag;
  assign io_coef_out_payload_0_45_45_real = int_reg_array_45_45_real;
  assign io_coef_out_payload_0_45_45_imag = int_reg_array_45_45_imag;
  assign io_coef_out_payload_0_45_46_real = int_reg_array_45_46_real;
  assign io_coef_out_payload_0_45_46_imag = int_reg_array_45_46_imag;
  assign io_coef_out_payload_0_45_47_real = int_reg_array_45_47_real;
  assign io_coef_out_payload_0_45_47_imag = int_reg_array_45_47_imag;
  assign io_coef_out_payload_0_45_48_real = int_reg_array_45_48_real;
  assign io_coef_out_payload_0_45_48_imag = int_reg_array_45_48_imag;
  assign io_coef_out_payload_0_45_49_real = int_reg_array_45_49_real;
  assign io_coef_out_payload_0_45_49_imag = int_reg_array_45_49_imag;
  assign io_coef_out_payload_0_46_0_real = int_reg_array_46_0_real;
  assign io_coef_out_payload_0_46_0_imag = int_reg_array_46_0_imag;
  assign io_coef_out_payload_0_46_1_real = int_reg_array_46_1_real;
  assign io_coef_out_payload_0_46_1_imag = int_reg_array_46_1_imag;
  assign io_coef_out_payload_0_46_2_real = int_reg_array_46_2_real;
  assign io_coef_out_payload_0_46_2_imag = int_reg_array_46_2_imag;
  assign io_coef_out_payload_0_46_3_real = int_reg_array_46_3_real;
  assign io_coef_out_payload_0_46_3_imag = int_reg_array_46_3_imag;
  assign io_coef_out_payload_0_46_4_real = int_reg_array_46_4_real;
  assign io_coef_out_payload_0_46_4_imag = int_reg_array_46_4_imag;
  assign io_coef_out_payload_0_46_5_real = int_reg_array_46_5_real;
  assign io_coef_out_payload_0_46_5_imag = int_reg_array_46_5_imag;
  assign io_coef_out_payload_0_46_6_real = int_reg_array_46_6_real;
  assign io_coef_out_payload_0_46_6_imag = int_reg_array_46_6_imag;
  assign io_coef_out_payload_0_46_7_real = int_reg_array_46_7_real;
  assign io_coef_out_payload_0_46_7_imag = int_reg_array_46_7_imag;
  assign io_coef_out_payload_0_46_8_real = int_reg_array_46_8_real;
  assign io_coef_out_payload_0_46_8_imag = int_reg_array_46_8_imag;
  assign io_coef_out_payload_0_46_9_real = int_reg_array_46_9_real;
  assign io_coef_out_payload_0_46_9_imag = int_reg_array_46_9_imag;
  assign io_coef_out_payload_0_46_10_real = int_reg_array_46_10_real;
  assign io_coef_out_payload_0_46_10_imag = int_reg_array_46_10_imag;
  assign io_coef_out_payload_0_46_11_real = int_reg_array_46_11_real;
  assign io_coef_out_payload_0_46_11_imag = int_reg_array_46_11_imag;
  assign io_coef_out_payload_0_46_12_real = int_reg_array_46_12_real;
  assign io_coef_out_payload_0_46_12_imag = int_reg_array_46_12_imag;
  assign io_coef_out_payload_0_46_13_real = int_reg_array_46_13_real;
  assign io_coef_out_payload_0_46_13_imag = int_reg_array_46_13_imag;
  assign io_coef_out_payload_0_46_14_real = int_reg_array_46_14_real;
  assign io_coef_out_payload_0_46_14_imag = int_reg_array_46_14_imag;
  assign io_coef_out_payload_0_46_15_real = int_reg_array_46_15_real;
  assign io_coef_out_payload_0_46_15_imag = int_reg_array_46_15_imag;
  assign io_coef_out_payload_0_46_16_real = int_reg_array_46_16_real;
  assign io_coef_out_payload_0_46_16_imag = int_reg_array_46_16_imag;
  assign io_coef_out_payload_0_46_17_real = int_reg_array_46_17_real;
  assign io_coef_out_payload_0_46_17_imag = int_reg_array_46_17_imag;
  assign io_coef_out_payload_0_46_18_real = int_reg_array_46_18_real;
  assign io_coef_out_payload_0_46_18_imag = int_reg_array_46_18_imag;
  assign io_coef_out_payload_0_46_19_real = int_reg_array_46_19_real;
  assign io_coef_out_payload_0_46_19_imag = int_reg_array_46_19_imag;
  assign io_coef_out_payload_0_46_20_real = int_reg_array_46_20_real;
  assign io_coef_out_payload_0_46_20_imag = int_reg_array_46_20_imag;
  assign io_coef_out_payload_0_46_21_real = int_reg_array_46_21_real;
  assign io_coef_out_payload_0_46_21_imag = int_reg_array_46_21_imag;
  assign io_coef_out_payload_0_46_22_real = int_reg_array_46_22_real;
  assign io_coef_out_payload_0_46_22_imag = int_reg_array_46_22_imag;
  assign io_coef_out_payload_0_46_23_real = int_reg_array_46_23_real;
  assign io_coef_out_payload_0_46_23_imag = int_reg_array_46_23_imag;
  assign io_coef_out_payload_0_46_24_real = int_reg_array_46_24_real;
  assign io_coef_out_payload_0_46_24_imag = int_reg_array_46_24_imag;
  assign io_coef_out_payload_0_46_25_real = int_reg_array_46_25_real;
  assign io_coef_out_payload_0_46_25_imag = int_reg_array_46_25_imag;
  assign io_coef_out_payload_0_46_26_real = int_reg_array_46_26_real;
  assign io_coef_out_payload_0_46_26_imag = int_reg_array_46_26_imag;
  assign io_coef_out_payload_0_46_27_real = int_reg_array_46_27_real;
  assign io_coef_out_payload_0_46_27_imag = int_reg_array_46_27_imag;
  assign io_coef_out_payload_0_46_28_real = int_reg_array_46_28_real;
  assign io_coef_out_payload_0_46_28_imag = int_reg_array_46_28_imag;
  assign io_coef_out_payload_0_46_29_real = int_reg_array_46_29_real;
  assign io_coef_out_payload_0_46_29_imag = int_reg_array_46_29_imag;
  assign io_coef_out_payload_0_46_30_real = int_reg_array_46_30_real;
  assign io_coef_out_payload_0_46_30_imag = int_reg_array_46_30_imag;
  assign io_coef_out_payload_0_46_31_real = int_reg_array_46_31_real;
  assign io_coef_out_payload_0_46_31_imag = int_reg_array_46_31_imag;
  assign io_coef_out_payload_0_46_32_real = int_reg_array_46_32_real;
  assign io_coef_out_payload_0_46_32_imag = int_reg_array_46_32_imag;
  assign io_coef_out_payload_0_46_33_real = int_reg_array_46_33_real;
  assign io_coef_out_payload_0_46_33_imag = int_reg_array_46_33_imag;
  assign io_coef_out_payload_0_46_34_real = int_reg_array_46_34_real;
  assign io_coef_out_payload_0_46_34_imag = int_reg_array_46_34_imag;
  assign io_coef_out_payload_0_46_35_real = int_reg_array_46_35_real;
  assign io_coef_out_payload_0_46_35_imag = int_reg_array_46_35_imag;
  assign io_coef_out_payload_0_46_36_real = int_reg_array_46_36_real;
  assign io_coef_out_payload_0_46_36_imag = int_reg_array_46_36_imag;
  assign io_coef_out_payload_0_46_37_real = int_reg_array_46_37_real;
  assign io_coef_out_payload_0_46_37_imag = int_reg_array_46_37_imag;
  assign io_coef_out_payload_0_46_38_real = int_reg_array_46_38_real;
  assign io_coef_out_payload_0_46_38_imag = int_reg_array_46_38_imag;
  assign io_coef_out_payload_0_46_39_real = int_reg_array_46_39_real;
  assign io_coef_out_payload_0_46_39_imag = int_reg_array_46_39_imag;
  assign io_coef_out_payload_0_46_40_real = int_reg_array_46_40_real;
  assign io_coef_out_payload_0_46_40_imag = int_reg_array_46_40_imag;
  assign io_coef_out_payload_0_46_41_real = int_reg_array_46_41_real;
  assign io_coef_out_payload_0_46_41_imag = int_reg_array_46_41_imag;
  assign io_coef_out_payload_0_46_42_real = int_reg_array_46_42_real;
  assign io_coef_out_payload_0_46_42_imag = int_reg_array_46_42_imag;
  assign io_coef_out_payload_0_46_43_real = int_reg_array_46_43_real;
  assign io_coef_out_payload_0_46_43_imag = int_reg_array_46_43_imag;
  assign io_coef_out_payload_0_46_44_real = int_reg_array_46_44_real;
  assign io_coef_out_payload_0_46_44_imag = int_reg_array_46_44_imag;
  assign io_coef_out_payload_0_46_45_real = int_reg_array_46_45_real;
  assign io_coef_out_payload_0_46_45_imag = int_reg_array_46_45_imag;
  assign io_coef_out_payload_0_46_46_real = int_reg_array_46_46_real;
  assign io_coef_out_payload_0_46_46_imag = int_reg_array_46_46_imag;
  assign io_coef_out_payload_0_46_47_real = int_reg_array_46_47_real;
  assign io_coef_out_payload_0_46_47_imag = int_reg_array_46_47_imag;
  assign io_coef_out_payload_0_46_48_real = int_reg_array_46_48_real;
  assign io_coef_out_payload_0_46_48_imag = int_reg_array_46_48_imag;
  assign io_coef_out_payload_0_46_49_real = int_reg_array_46_49_real;
  assign io_coef_out_payload_0_46_49_imag = int_reg_array_46_49_imag;
  assign io_coef_out_payload_0_47_0_real = int_reg_array_47_0_real;
  assign io_coef_out_payload_0_47_0_imag = int_reg_array_47_0_imag;
  assign io_coef_out_payload_0_47_1_real = int_reg_array_47_1_real;
  assign io_coef_out_payload_0_47_1_imag = int_reg_array_47_1_imag;
  assign io_coef_out_payload_0_47_2_real = int_reg_array_47_2_real;
  assign io_coef_out_payload_0_47_2_imag = int_reg_array_47_2_imag;
  assign io_coef_out_payload_0_47_3_real = int_reg_array_47_3_real;
  assign io_coef_out_payload_0_47_3_imag = int_reg_array_47_3_imag;
  assign io_coef_out_payload_0_47_4_real = int_reg_array_47_4_real;
  assign io_coef_out_payload_0_47_4_imag = int_reg_array_47_4_imag;
  assign io_coef_out_payload_0_47_5_real = int_reg_array_47_5_real;
  assign io_coef_out_payload_0_47_5_imag = int_reg_array_47_5_imag;
  assign io_coef_out_payload_0_47_6_real = int_reg_array_47_6_real;
  assign io_coef_out_payload_0_47_6_imag = int_reg_array_47_6_imag;
  assign io_coef_out_payload_0_47_7_real = int_reg_array_47_7_real;
  assign io_coef_out_payload_0_47_7_imag = int_reg_array_47_7_imag;
  assign io_coef_out_payload_0_47_8_real = int_reg_array_47_8_real;
  assign io_coef_out_payload_0_47_8_imag = int_reg_array_47_8_imag;
  assign io_coef_out_payload_0_47_9_real = int_reg_array_47_9_real;
  assign io_coef_out_payload_0_47_9_imag = int_reg_array_47_9_imag;
  assign io_coef_out_payload_0_47_10_real = int_reg_array_47_10_real;
  assign io_coef_out_payload_0_47_10_imag = int_reg_array_47_10_imag;
  assign io_coef_out_payload_0_47_11_real = int_reg_array_47_11_real;
  assign io_coef_out_payload_0_47_11_imag = int_reg_array_47_11_imag;
  assign io_coef_out_payload_0_47_12_real = int_reg_array_47_12_real;
  assign io_coef_out_payload_0_47_12_imag = int_reg_array_47_12_imag;
  assign io_coef_out_payload_0_47_13_real = int_reg_array_47_13_real;
  assign io_coef_out_payload_0_47_13_imag = int_reg_array_47_13_imag;
  assign io_coef_out_payload_0_47_14_real = int_reg_array_47_14_real;
  assign io_coef_out_payload_0_47_14_imag = int_reg_array_47_14_imag;
  assign io_coef_out_payload_0_47_15_real = int_reg_array_47_15_real;
  assign io_coef_out_payload_0_47_15_imag = int_reg_array_47_15_imag;
  assign io_coef_out_payload_0_47_16_real = int_reg_array_47_16_real;
  assign io_coef_out_payload_0_47_16_imag = int_reg_array_47_16_imag;
  assign io_coef_out_payload_0_47_17_real = int_reg_array_47_17_real;
  assign io_coef_out_payload_0_47_17_imag = int_reg_array_47_17_imag;
  assign io_coef_out_payload_0_47_18_real = int_reg_array_47_18_real;
  assign io_coef_out_payload_0_47_18_imag = int_reg_array_47_18_imag;
  assign io_coef_out_payload_0_47_19_real = int_reg_array_47_19_real;
  assign io_coef_out_payload_0_47_19_imag = int_reg_array_47_19_imag;
  assign io_coef_out_payload_0_47_20_real = int_reg_array_47_20_real;
  assign io_coef_out_payload_0_47_20_imag = int_reg_array_47_20_imag;
  assign io_coef_out_payload_0_47_21_real = int_reg_array_47_21_real;
  assign io_coef_out_payload_0_47_21_imag = int_reg_array_47_21_imag;
  assign io_coef_out_payload_0_47_22_real = int_reg_array_47_22_real;
  assign io_coef_out_payload_0_47_22_imag = int_reg_array_47_22_imag;
  assign io_coef_out_payload_0_47_23_real = int_reg_array_47_23_real;
  assign io_coef_out_payload_0_47_23_imag = int_reg_array_47_23_imag;
  assign io_coef_out_payload_0_47_24_real = int_reg_array_47_24_real;
  assign io_coef_out_payload_0_47_24_imag = int_reg_array_47_24_imag;
  assign io_coef_out_payload_0_47_25_real = int_reg_array_47_25_real;
  assign io_coef_out_payload_0_47_25_imag = int_reg_array_47_25_imag;
  assign io_coef_out_payload_0_47_26_real = int_reg_array_47_26_real;
  assign io_coef_out_payload_0_47_26_imag = int_reg_array_47_26_imag;
  assign io_coef_out_payload_0_47_27_real = int_reg_array_47_27_real;
  assign io_coef_out_payload_0_47_27_imag = int_reg_array_47_27_imag;
  assign io_coef_out_payload_0_47_28_real = int_reg_array_47_28_real;
  assign io_coef_out_payload_0_47_28_imag = int_reg_array_47_28_imag;
  assign io_coef_out_payload_0_47_29_real = int_reg_array_47_29_real;
  assign io_coef_out_payload_0_47_29_imag = int_reg_array_47_29_imag;
  assign io_coef_out_payload_0_47_30_real = int_reg_array_47_30_real;
  assign io_coef_out_payload_0_47_30_imag = int_reg_array_47_30_imag;
  assign io_coef_out_payload_0_47_31_real = int_reg_array_47_31_real;
  assign io_coef_out_payload_0_47_31_imag = int_reg_array_47_31_imag;
  assign io_coef_out_payload_0_47_32_real = int_reg_array_47_32_real;
  assign io_coef_out_payload_0_47_32_imag = int_reg_array_47_32_imag;
  assign io_coef_out_payload_0_47_33_real = int_reg_array_47_33_real;
  assign io_coef_out_payload_0_47_33_imag = int_reg_array_47_33_imag;
  assign io_coef_out_payload_0_47_34_real = int_reg_array_47_34_real;
  assign io_coef_out_payload_0_47_34_imag = int_reg_array_47_34_imag;
  assign io_coef_out_payload_0_47_35_real = int_reg_array_47_35_real;
  assign io_coef_out_payload_0_47_35_imag = int_reg_array_47_35_imag;
  assign io_coef_out_payload_0_47_36_real = int_reg_array_47_36_real;
  assign io_coef_out_payload_0_47_36_imag = int_reg_array_47_36_imag;
  assign io_coef_out_payload_0_47_37_real = int_reg_array_47_37_real;
  assign io_coef_out_payload_0_47_37_imag = int_reg_array_47_37_imag;
  assign io_coef_out_payload_0_47_38_real = int_reg_array_47_38_real;
  assign io_coef_out_payload_0_47_38_imag = int_reg_array_47_38_imag;
  assign io_coef_out_payload_0_47_39_real = int_reg_array_47_39_real;
  assign io_coef_out_payload_0_47_39_imag = int_reg_array_47_39_imag;
  assign io_coef_out_payload_0_47_40_real = int_reg_array_47_40_real;
  assign io_coef_out_payload_0_47_40_imag = int_reg_array_47_40_imag;
  assign io_coef_out_payload_0_47_41_real = int_reg_array_47_41_real;
  assign io_coef_out_payload_0_47_41_imag = int_reg_array_47_41_imag;
  assign io_coef_out_payload_0_47_42_real = int_reg_array_47_42_real;
  assign io_coef_out_payload_0_47_42_imag = int_reg_array_47_42_imag;
  assign io_coef_out_payload_0_47_43_real = int_reg_array_47_43_real;
  assign io_coef_out_payload_0_47_43_imag = int_reg_array_47_43_imag;
  assign io_coef_out_payload_0_47_44_real = int_reg_array_47_44_real;
  assign io_coef_out_payload_0_47_44_imag = int_reg_array_47_44_imag;
  assign io_coef_out_payload_0_47_45_real = int_reg_array_47_45_real;
  assign io_coef_out_payload_0_47_45_imag = int_reg_array_47_45_imag;
  assign io_coef_out_payload_0_47_46_real = int_reg_array_47_46_real;
  assign io_coef_out_payload_0_47_46_imag = int_reg_array_47_46_imag;
  assign io_coef_out_payload_0_47_47_real = int_reg_array_47_47_real;
  assign io_coef_out_payload_0_47_47_imag = int_reg_array_47_47_imag;
  assign io_coef_out_payload_0_47_48_real = int_reg_array_47_48_real;
  assign io_coef_out_payload_0_47_48_imag = int_reg_array_47_48_imag;
  assign io_coef_out_payload_0_47_49_real = int_reg_array_47_49_real;
  assign io_coef_out_payload_0_47_49_imag = int_reg_array_47_49_imag;
  assign io_coef_out_payload_0_48_0_real = int_reg_array_48_0_real;
  assign io_coef_out_payload_0_48_0_imag = int_reg_array_48_0_imag;
  assign io_coef_out_payload_0_48_1_real = int_reg_array_48_1_real;
  assign io_coef_out_payload_0_48_1_imag = int_reg_array_48_1_imag;
  assign io_coef_out_payload_0_48_2_real = int_reg_array_48_2_real;
  assign io_coef_out_payload_0_48_2_imag = int_reg_array_48_2_imag;
  assign io_coef_out_payload_0_48_3_real = int_reg_array_48_3_real;
  assign io_coef_out_payload_0_48_3_imag = int_reg_array_48_3_imag;
  assign io_coef_out_payload_0_48_4_real = int_reg_array_48_4_real;
  assign io_coef_out_payload_0_48_4_imag = int_reg_array_48_4_imag;
  assign io_coef_out_payload_0_48_5_real = int_reg_array_48_5_real;
  assign io_coef_out_payload_0_48_5_imag = int_reg_array_48_5_imag;
  assign io_coef_out_payload_0_48_6_real = int_reg_array_48_6_real;
  assign io_coef_out_payload_0_48_6_imag = int_reg_array_48_6_imag;
  assign io_coef_out_payload_0_48_7_real = int_reg_array_48_7_real;
  assign io_coef_out_payload_0_48_7_imag = int_reg_array_48_7_imag;
  assign io_coef_out_payload_0_48_8_real = int_reg_array_48_8_real;
  assign io_coef_out_payload_0_48_8_imag = int_reg_array_48_8_imag;
  assign io_coef_out_payload_0_48_9_real = int_reg_array_48_9_real;
  assign io_coef_out_payload_0_48_9_imag = int_reg_array_48_9_imag;
  assign io_coef_out_payload_0_48_10_real = int_reg_array_48_10_real;
  assign io_coef_out_payload_0_48_10_imag = int_reg_array_48_10_imag;
  assign io_coef_out_payload_0_48_11_real = int_reg_array_48_11_real;
  assign io_coef_out_payload_0_48_11_imag = int_reg_array_48_11_imag;
  assign io_coef_out_payload_0_48_12_real = int_reg_array_48_12_real;
  assign io_coef_out_payload_0_48_12_imag = int_reg_array_48_12_imag;
  assign io_coef_out_payload_0_48_13_real = int_reg_array_48_13_real;
  assign io_coef_out_payload_0_48_13_imag = int_reg_array_48_13_imag;
  assign io_coef_out_payload_0_48_14_real = int_reg_array_48_14_real;
  assign io_coef_out_payload_0_48_14_imag = int_reg_array_48_14_imag;
  assign io_coef_out_payload_0_48_15_real = int_reg_array_48_15_real;
  assign io_coef_out_payload_0_48_15_imag = int_reg_array_48_15_imag;
  assign io_coef_out_payload_0_48_16_real = int_reg_array_48_16_real;
  assign io_coef_out_payload_0_48_16_imag = int_reg_array_48_16_imag;
  assign io_coef_out_payload_0_48_17_real = int_reg_array_48_17_real;
  assign io_coef_out_payload_0_48_17_imag = int_reg_array_48_17_imag;
  assign io_coef_out_payload_0_48_18_real = int_reg_array_48_18_real;
  assign io_coef_out_payload_0_48_18_imag = int_reg_array_48_18_imag;
  assign io_coef_out_payload_0_48_19_real = int_reg_array_48_19_real;
  assign io_coef_out_payload_0_48_19_imag = int_reg_array_48_19_imag;
  assign io_coef_out_payload_0_48_20_real = int_reg_array_48_20_real;
  assign io_coef_out_payload_0_48_20_imag = int_reg_array_48_20_imag;
  assign io_coef_out_payload_0_48_21_real = int_reg_array_48_21_real;
  assign io_coef_out_payload_0_48_21_imag = int_reg_array_48_21_imag;
  assign io_coef_out_payload_0_48_22_real = int_reg_array_48_22_real;
  assign io_coef_out_payload_0_48_22_imag = int_reg_array_48_22_imag;
  assign io_coef_out_payload_0_48_23_real = int_reg_array_48_23_real;
  assign io_coef_out_payload_0_48_23_imag = int_reg_array_48_23_imag;
  assign io_coef_out_payload_0_48_24_real = int_reg_array_48_24_real;
  assign io_coef_out_payload_0_48_24_imag = int_reg_array_48_24_imag;
  assign io_coef_out_payload_0_48_25_real = int_reg_array_48_25_real;
  assign io_coef_out_payload_0_48_25_imag = int_reg_array_48_25_imag;
  assign io_coef_out_payload_0_48_26_real = int_reg_array_48_26_real;
  assign io_coef_out_payload_0_48_26_imag = int_reg_array_48_26_imag;
  assign io_coef_out_payload_0_48_27_real = int_reg_array_48_27_real;
  assign io_coef_out_payload_0_48_27_imag = int_reg_array_48_27_imag;
  assign io_coef_out_payload_0_48_28_real = int_reg_array_48_28_real;
  assign io_coef_out_payload_0_48_28_imag = int_reg_array_48_28_imag;
  assign io_coef_out_payload_0_48_29_real = int_reg_array_48_29_real;
  assign io_coef_out_payload_0_48_29_imag = int_reg_array_48_29_imag;
  assign io_coef_out_payload_0_48_30_real = int_reg_array_48_30_real;
  assign io_coef_out_payload_0_48_30_imag = int_reg_array_48_30_imag;
  assign io_coef_out_payload_0_48_31_real = int_reg_array_48_31_real;
  assign io_coef_out_payload_0_48_31_imag = int_reg_array_48_31_imag;
  assign io_coef_out_payload_0_48_32_real = int_reg_array_48_32_real;
  assign io_coef_out_payload_0_48_32_imag = int_reg_array_48_32_imag;
  assign io_coef_out_payload_0_48_33_real = int_reg_array_48_33_real;
  assign io_coef_out_payload_0_48_33_imag = int_reg_array_48_33_imag;
  assign io_coef_out_payload_0_48_34_real = int_reg_array_48_34_real;
  assign io_coef_out_payload_0_48_34_imag = int_reg_array_48_34_imag;
  assign io_coef_out_payload_0_48_35_real = int_reg_array_48_35_real;
  assign io_coef_out_payload_0_48_35_imag = int_reg_array_48_35_imag;
  assign io_coef_out_payload_0_48_36_real = int_reg_array_48_36_real;
  assign io_coef_out_payload_0_48_36_imag = int_reg_array_48_36_imag;
  assign io_coef_out_payload_0_48_37_real = int_reg_array_48_37_real;
  assign io_coef_out_payload_0_48_37_imag = int_reg_array_48_37_imag;
  assign io_coef_out_payload_0_48_38_real = int_reg_array_48_38_real;
  assign io_coef_out_payload_0_48_38_imag = int_reg_array_48_38_imag;
  assign io_coef_out_payload_0_48_39_real = int_reg_array_48_39_real;
  assign io_coef_out_payload_0_48_39_imag = int_reg_array_48_39_imag;
  assign io_coef_out_payload_0_48_40_real = int_reg_array_48_40_real;
  assign io_coef_out_payload_0_48_40_imag = int_reg_array_48_40_imag;
  assign io_coef_out_payload_0_48_41_real = int_reg_array_48_41_real;
  assign io_coef_out_payload_0_48_41_imag = int_reg_array_48_41_imag;
  assign io_coef_out_payload_0_48_42_real = int_reg_array_48_42_real;
  assign io_coef_out_payload_0_48_42_imag = int_reg_array_48_42_imag;
  assign io_coef_out_payload_0_48_43_real = int_reg_array_48_43_real;
  assign io_coef_out_payload_0_48_43_imag = int_reg_array_48_43_imag;
  assign io_coef_out_payload_0_48_44_real = int_reg_array_48_44_real;
  assign io_coef_out_payload_0_48_44_imag = int_reg_array_48_44_imag;
  assign io_coef_out_payload_0_48_45_real = int_reg_array_48_45_real;
  assign io_coef_out_payload_0_48_45_imag = int_reg_array_48_45_imag;
  assign io_coef_out_payload_0_48_46_real = int_reg_array_48_46_real;
  assign io_coef_out_payload_0_48_46_imag = int_reg_array_48_46_imag;
  assign io_coef_out_payload_0_48_47_real = int_reg_array_48_47_real;
  assign io_coef_out_payload_0_48_47_imag = int_reg_array_48_47_imag;
  assign io_coef_out_payload_0_48_48_real = int_reg_array_48_48_real;
  assign io_coef_out_payload_0_48_48_imag = int_reg_array_48_48_imag;
  assign io_coef_out_payload_0_48_49_real = int_reg_array_48_49_real;
  assign io_coef_out_payload_0_48_49_imag = int_reg_array_48_49_imag;
  assign io_coef_out_payload_0_49_0_real = int_reg_array_49_0_real;
  assign io_coef_out_payload_0_49_0_imag = int_reg_array_49_0_imag;
  assign io_coef_out_payload_0_49_1_real = int_reg_array_49_1_real;
  assign io_coef_out_payload_0_49_1_imag = int_reg_array_49_1_imag;
  assign io_coef_out_payload_0_49_2_real = int_reg_array_49_2_real;
  assign io_coef_out_payload_0_49_2_imag = int_reg_array_49_2_imag;
  assign io_coef_out_payload_0_49_3_real = int_reg_array_49_3_real;
  assign io_coef_out_payload_0_49_3_imag = int_reg_array_49_3_imag;
  assign io_coef_out_payload_0_49_4_real = int_reg_array_49_4_real;
  assign io_coef_out_payload_0_49_4_imag = int_reg_array_49_4_imag;
  assign io_coef_out_payload_0_49_5_real = int_reg_array_49_5_real;
  assign io_coef_out_payload_0_49_5_imag = int_reg_array_49_5_imag;
  assign io_coef_out_payload_0_49_6_real = int_reg_array_49_6_real;
  assign io_coef_out_payload_0_49_6_imag = int_reg_array_49_6_imag;
  assign io_coef_out_payload_0_49_7_real = int_reg_array_49_7_real;
  assign io_coef_out_payload_0_49_7_imag = int_reg_array_49_7_imag;
  assign io_coef_out_payload_0_49_8_real = int_reg_array_49_8_real;
  assign io_coef_out_payload_0_49_8_imag = int_reg_array_49_8_imag;
  assign io_coef_out_payload_0_49_9_real = int_reg_array_49_9_real;
  assign io_coef_out_payload_0_49_9_imag = int_reg_array_49_9_imag;
  assign io_coef_out_payload_0_49_10_real = int_reg_array_49_10_real;
  assign io_coef_out_payload_0_49_10_imag = int_reg_array_49_10_imag;
  assign io_coef_out_payload_0_49_11_real = int_reg_array_49_11_real;
  assign io_coef_out_payload_0_49_11_imag = int_reg_array_49_11_imag;
  assign io_coef_out_payload_0_49_12_real = int_reg_array_49_12_real;
  assign io_coef_out_payload_0_49_12_imag = int_reg_array_49_12_imag;
  assign io_coef_out_payload_0_49_13_real = int_reg_array_49_13_real;
  assign io_coef_out_payload_0_49_13_imag = int_reg_array_49_13_imag;
  assign io_coef_out_payload_0_49_14_real = int_reg_array_49_14_real;
  assign io_coef_out_payload_0_49_14_imag = int_reg_array_49_14_imag;
  assign io_coef_out_payload_0_49_15_real = int_reg_array_49_15_real;
  assign io_coef_out_payload_0_49_15_imag = int_reg_array_49_15_imag;
  assign io_coef_out_payload_0_49_16_real = int_reg_array_49_16_real;
  assign io_coef_out_payload_0_49_16_imag = int_reg_array_49_16_imag;
  assign io_coef_out_payload_0_49_17_real = int_reg_array_49_17_real;
  assign io_coef_out_payload_0_49_17_imag = int_reg_array_49_17_imag;
  assign io_coef_out_payload_0_49_18_real = int_reg_array_49_18_real;
  assign io_coef_out_payload_0_49_18_imag = int_reg_array_49_18_imag;
  assign io_coef_out_payload_0_49_19_real = int_reg_array_49_19_real;
  assign io_coef_out_payload_0_49_19_imag = int_reg_array_49_19_imag;
  assign io_coef_out_payload_0_49_20_real = int_reg_array_49_20_real;
  assign io_coef_out_payload_0_49_20_imag = int_reg_array_49_20_imag;
  assign io_coef_out_payload_0_49_21_real = int_reg_array_49_21_real;
  assign io_coef_out_payload_0_49_21_imag = int_reg_array_49_21_imag;
  assign io_coef_out_payload_0_49_22_real = int_reg_array_49_22_real;
  assign io_coef_out_payload_0_49_22_imag = int_reg_array_49_22_imag;
  assign io_coef_out_payload_0_49_23_real = int_reg_array_49_23_real;
  assign io_coef_out_payload_0_49_23_imag = int_reg_array_49_23_imag;
  assign io_coef_out_payload_0_49_24_real = int_reg_array_49_24_real;
  assign io_coef_out_payload_0_49_24_imag = int_reg_array_49_24_imag;
  assign io_coef_out_payload_0_49_25_real = int_reg_array_49_25_real;
  assign io_coef_out_payload_0_49_25_imag = int_reg_array_49_25_imag;
  assign io_coef_out_payload_0_49_26_real = int_reg_array_49_26_real;
  assign io_coef_out_payload_0_49_26_imag = int_reg_array_49_26_imag;
  assign io_coef_out_payload_0_49_27_real = int_reg_array_49_27_real;
  assign io_coef_out_payload_0_49_27_imag = int_reg_array_49_27_imag;
  assign io_coef_out_payload_0_49_28_real = int_reg_array_49_28_real;
  assign io_coef_out_payload_0_49_28_imag = int_reg_array_49_28_imag;
  assign io_coef_out_payload_0_49_29_real = int_reg_array_49_29_real;
  assign io_coef_out_payload_0_49_29_imag = int_reg_array_49_29_imag;
  assign io_coef_out_payload_0_49_30_real = int_reg_array_49_30_real;
  assign io_coef_out_payload_0_49_30_imag = int_reg_array_49_30_imag;
  assign io_coef_out_payload_0_49_31_real = int_reg_array_49_31_real;
  assign io_coef_out_payload_0_49_31_imag = int_reg_array_49_31_imag;
  assign io_coef_out_payload_0_49_32_real = int_reg_array_49_32_real;
  assign io_coef_out_payload_0_49_32_imag = int_reg_array_49_32_imag;
  assign io_coef_out_payload_0_49_33_real = int_reg_array_49_33_real;
  assign io_coef_out_payload_0_49_33_imag = int_reg_array_49_33_imag;
  assign io_coef_out_payload_0_49_34_real = int_reg_array_49_34_real;
  assign io_coef_out_payload_0_49_34_imag = int_reg_array_49_34_imag;
  assign io_coef_out_payload_0_49_35_real = int_reg_array_49_35_real;
  assign io_coef_out_payload_0_49_35_imag = int_reg_array_49_35_imag;
  assign io_coef_out_payload_0_49_36_real = int_reg_array_49_36_real;
  assign io_coef_out_payload_0_49_36_imag = int_reg_array_49_36_imag;
  assign io_coef_out_payload_0_49_37_real = int_reg_array_49_37_real;
  assign io_coef_out_payload_0_49_37_imag = int_reg_array_49_37_imag;
  assign io_coef_out_payload_0_49_38_real = int_reg_array_49_38_real;
  assign io_coef_out_payload_0_49_38_imag = int_reg_array_49_38_imag;
  assign io_coef_out_payload_0_49_39_real = int_reg_array_49_39_real;
  assign io_coef_out_payload_0_49_39_imag = int_reg_array_49_39_imag;
  assign io_coef_out_payload_0_49_40_real = int_reg_array_49_40_real;
  assign io_coef_out_payload_0_49_40_imag = int_reg_array_49_40_imag;
  assign io_coef_out_payload_0_49_41_real = int_reg_array_49_41_real;
  assign io_coef_out_payload_0_49_41_imag = int_reg_array_49_41_imag;
  assign io_coef_out_payload_0_49_42_real = int_reg_array_49_42_real;
  assign io_coef_out_payload_0_49_42_imag = int_reg_array_49_42_imag;
  assign io_coef_out_payload_0_49_43_real = int_reg_array_49_43_real;
  assign io_coef_out_payload_0_49_43_imag = int_reg_array_49_43_imag;
  assign io_coef_out_payload_0_49_44_real = int_reg_array_49_44_real;
  assign io_coef_out_payload_0_49_44_imag = int_reg_array_49_44_imag;
  assign io_coef_out_payload_0_49_45_real = int_reg_array_49_45_real;
  assign io_coef_out_payload_0_49_45_imag = int_reg_array_49_45_imag;
  assign io_coef_out_payload_0_49_46_real = int_reg_array_49_46_real;
  assign io_coef_out_payload_0_49_46_imag = int_reg_array_49_46_imag;
  assign io_coef_out_payload_0_49_47_real = int_reg_array_49_47_real;
  assign io_coef_out_payload_0_49_47_imag = int_reg_array_49_47_imag;
  assign io_coef_out_payload_0_49_48_real = int_reg_array_49_48_real;
  assign io_coef_out_payload_0_49_48_imag = int_reg_array_49_48_imag;
  assign io_coef_out_payload_0_49_49_real = int_reg_array_49_49_real;
  assign io_coef_out_payload_0_49_49_imag = int_reg_array_49_49_imag;
  always @ (posedge clk) begin
    if(axi4_aw_valid)begin
      aw_area_awaddr_r <= axi4_aw_payload_addr;
      aw_area_awlen_r <= axi4_aw_payload_len;
      aw_area_awsize_r <= axi4_aw_payload_size;
      aw_area_awid_r <= axi4_aw_payload_id;
    end
    if(axi4_w_valid)begin
      transfer_done <= (((32'h0 <= load_data_area_current_addr) && (load_data_area_current_addr < 32'h0)) ? axi4_w_payload_data_regNext[0] : _zz_2856_[0]);
      if(_zz_4_)begin
        int_reg_array_0_0_real <= _zz_55_;
      end
      if(_zz_5_)begin
        int_reg_array_0_1_real <= _zz_55_;
      end
      if(_zz_6_)begin
        int_reg_array_0_2_real <= _zz_55_;
      end
      if(_zz_7_)begin
        int_reg_array_0_3_real <= _zz_55_;
      end
      if(_zz_8_)begin
        int_reg_array_0_4_real <= _zz_55_;
      end
      if(_zz_9_)begin
        int_reg_array_0_5_real <= _zz_55_;
      end
      if(_zz_10_)begin
        int_reg_array_0_6_real <= _zz_55_;
      end
      if(_zz_11_)begin
        int_reg_array_0_7_real <= _zz_55_;
      end
      if(_zz_12_)begin
        int_reg_array_0_8_real <= _zz_55_;
      end
      if(_zz_13_)begin
        int_reg_array_0_9_real <= _zz_55_;
      end
      if(_zz_14_)begin
        int_reg_array_0_10_real <= _zz_55_;
      end
      if(_zz_15_)begin
        int_reg_array_0_11_real <= _zz_55_;
      end
      if(_zz_16_)begin
        int_reg_array_0_12_real <= _zz_55_;
      end
      if(_zz_17_)begin
        int_reg_array_0_13_real <= _zz_55_;
      end
      if(_zz_18_)begin
        int_reg_array_0_14_real <= _zz_55_;
      end
      if(_zz_19_)begin
        int_reg_array_0_15_real <= _zz_55_;
      end
      if(_zz_20_)begin
        int_reg_array_0_16_real <= _zz_55_;
      end
      if(_zz_21_)begin
        int_reg_array_0_17_real <= _zz_55_;
      end
      if(_zz_22_)begin
        int_reg_array_0_18_real <= _zz_55_;
      end
      if(_zz_23_)begin
        int_reg_array_0_19_real <= _zz_55_;
      end
      if(_zz_24_)begin
        int_reg_array_0_20_real <= _zz_55_;
      end
      if(_zz_25_)begin
        int_reg_array_0_21_real <= _zz_55_;
      end
      if(_zz_26_)begin
        int_reg_array_0_22_real <= _zz_55_;
      end
      if(_zz_27_)begin
        int_reg_array_0_23_real <= _zz_55_;
      end
      if(_zz_28_)begin
        int_reg_array_0_24_real <= _zz_55_;
      end
      if(_zz_29_)begin
        int_reg_array_0_25_real <= _zz_55_;
      end
      if(_zz_30_)begin
        int_reg_array_0_26_real <= _zz_55_;
      end
      if(_zz_31_)begin
        int_reg_array_0_27_real <= _zz_55_;
      end
      if(_zz_32_)begin
        int_reg_array_0_28_real <= _zz_55_;
      end
      if(_zz_33_)begin
        int_reg_array_0_29_real <= _zz_55_;
      end
      if(_zz_34_)begin
        int_reg_array_0_30_real <= _zz_55_;
      end
      if(_zz_35_)begin
        int_reg_array_0_31_real <= _zz_55_;
      end
      if(_zz_36_)begin
        int_reg_array_0_32_real <= _zz_55_;
      end
      if(_zz_37_)begin
        int_reg_array_0_33_real <= _zz_55_;
      end
      if(_zz_38_)begin
        int_reg_array_0_34_real <= _zz_55_;
      end
      if(_zz_39_)begin
        int_reg_array_0_35_real <= _zz_55_;
      end
      if(_zz_40_)begin
        int_reg_array_0_36_real <= _zz_55_;
      end
      if(_zz_41_)begin
        int_reg_array_0_37_real <= _zz_55_;
      end
      if(_zz_42_)begin
        int_reg_array_0_38_real <= _zz_55_;
      end
      if(_zz_43_)begin
        int_reg_array_0_39_real <= _zz_55_;
      end
      if(_zz_44_)begin
        int_reg_array_0_40_real <= _zz_55_;
      end
      if(_zz_45_)begin
        int_reg_array_0_41_real <= _zz_55_;
      end
      if(_zz_46_)begin
        int_reg_array_0_42_real <= _zz_55_;
      end
      if(_zz_47_)begin
        int_reg_array_0_43_real <= _zz_55_;
      end
      if(_zz_48_)begin
        int_reg_array_0_44_real <= _zz_55_;
      end
      if(_zz_49_)begin
        int_reg_array_0_45_real <= _zz_55_;
      end
      if(_zz_50_)begin
        int_reg_array_0_46_real <= _zz_55_;
      end
      if(_zz_51_)begin
        int_reg_array_0_47_real <= _zz_55_;
      end
      if(_zz_52_)begin
        int_reg_array_0_48_real <= _zz_55_;
      end
      if(_zz_53_)begin
        int_reg_array_0_49_real <= _zz_55_;
      end
      if(_zz_4_)begin
        int_reg_array_0_0_imag <= _zz_56_;
      end
      if(_zz_5_)begin
        int_reg_array_0_1_imag <= _zz_56_;
      end
      if(_zz_6_)begin
        int_reg_array_0_2_imag <= _zz_56_;
      end
      if(_zz_7_)begin
        int_reg_array_0_3_imag <= _zz_56_;
      end
      if(_zz_8_)begin
        int_reg_array_0_4_imag <= _zz_56_;
      end
      if(_zz_9_)begin
        int_reg_array_0_5_imag <= _zz_56_;
      end
      if(_zz_10_)begin
        int_reg_array_0_6_imag <= _zz_56_;
      end
      if(_zz_11_)begin
        int_reg_array_0_7_imag <= _zz_56_;
      end
      if(_zz_12_)begin
        int_reg_array_0_8_imag <= _zz_56_;
      end
      if(_zz_13_)begin
        int_reg_array_0_9_imag <= _zz_56_;
      end
      if(_zz_14_)begin
        int_reg_array_0_10_imag <= _zz_56_;
      end
      if(_zz_15_)begin
        int_reg_array_0_11_imag <= _zz_56_;
      end
      if(_zz_16_)begin
        int_reg_array_0_12_imag <= _zz_56_;
      end
      if(_zz_17_)begin
        int_reg_array_0_13_imag <= _zz_56_;
      end
      if(_zz_18_)begin
        int_reg_array_0_14_imag <= _zz_56_;
      end
      if(_zz_19_)begin
        int_reg_array_0_15_imag <= _zz_56_;
      end
      if(_zz_20_)begin
        int_reg_array_0_16_imag <= _zz_56_;
      end
      if(_zz_21_)begin
        int_reg_array_0_17_imag <= _zz_56_;
      end
      if(_zz_22_)begin
        int_reg_array_0_18_imag <= _zz_56_;
      end
      if(_zz_23_)begin
        int_reg_array_0_19_imag <= _zz_56_;
      end
      if(_zz_24_)begin
        int_reg_array_0_20_imag <= _zz_56_;
      end
      if(_zz_25_)begin
        int_reg_array_0_21_imag <= _zz_56_;
      end
      if(_zz_26_)begin
        int_reg_array_0_22_imag <= _zz_56_;
      end
      if(_zz_27_)begin
        int_reg_array_0_23_imag <= _zz_56_;
      end
      if(_zz_28_)begin
        int_reg_array_0_24_imag <= _zz_56_;
      end
      if(_zz_29_)begin
        int_reg_array_0_25_imag <= _zz_56_;
      end
      if(_zz_30_)begin
        int_reg_array_0_26_imag <= _zz_56_;
      end
      if(_zz_31_)begin
        int_reg_array_0_27_imag <= _zz_56_;
      end
      if(_zz_32_)begin
        int_reg_array_0_28_imag <= _zz_56_;
      end
      if(_zz_33_)begin
        int_reg_array_0_29_imag <= _zz_56_;
      end
      if(_zz_34_)begin
        int_reg_array_0_30_imag <= _zz_56_;
      end
      if(_zz_35_)begin
        int_reg_array_0_31_imag <= _zz_56_;
      end
      if(_zz_36_)begin
        int_reg_array_0_32_imag <= _zz_56_;
      end
      if(_zz_37_)begin
        int_reg_array_0_33_imag <= _zz_56_;
      end
      if(_zz_38_)begin
        int_reg_array_0_34_imag <= _zz_56_;
      end
      if(_zz_39_)begin
        int_reg_array_0_35_imag <= _zz_56_;
      end
      if(_zz_40_)begin
        int_reg_array_0_36_imag <= _zz_56_;
      end
      if(_zz_41_)begin
        int_reg_array_0_37_imag <= _zz_56_;
      end
      if(_zz_42_)begin
        int_reg_array_0_38_imag <= _zz_56_;
      end
      if(_zz_43_)begin
        int_reg_array_0_39_imag <= _zz_56_;
      end
      if(_zz_44_)begin
        int_reg_array_0_40_imag <= _zz_56_;
      end
      if(_zz_45_)begin
        int_reg_array_0_41_imag <= _zz_56_;
      end
      if(_zz_46_)begin
        int_reg_array_0_42_imag <= _zz_56_;
      end
      if(_zz_47_)begin
        int_reg_array_0_43_imag <= _zz_56_;
      end
      if(_zz_48_)begin
        int_reg_array_0_44_imag <= _zz_56_;
      end
      if(_zz_49_)begin
        int_reg_array_0_45_imag <= _zz_56_;
      end
      if(_zz_50_)begin
        int_reg_array_0_46_imag <= _zz_56_;
      end
      if(_zz_51_)begin
        int_reg_array_0_47_imag <= _zz_56_;
      end
      if(_zz_52_)begin
        int_reg_array_0_48_imag <= _zz_56_;
      end
      if(_zz_53_)begin
        int_reg_array_0_49_imag <= _zz_56_;
      end
      if(_zz_59_)begin
        int_reg_array_1_0_real <= _zz_110_;
      end
      if(_zz_60_)begin
        int_reg_array_1_1_real <= _zz_110_;
      end
      if(_zz_61_)begin
        int_reg_array_1_2_real <= _zz_110_;
      end
      if(_zz_62_)begin
        int_reg_array_1_3_real <= _zz_110_;
      end
      if(_zz_63_)begin
        int_reg_array_1_4_real <= _zz_110_;
      end
      if(_zz_64_)begin
        int_reg_array_1_5_real <= _zz_110_;
      end
      if(_zz_65_)begin
        int_reg_array_1_6_real <= _zz_110_;
      end
      if(_zz_66_)begin
        int_reg_array_1_7_real <= _zz_110_;
      end
      if(_zz_67_)begin
        int_reg_array_1_8_real <= _zz_110_;
      end
      if(_zz_68_)begin
        int_reg_array_1_9_real <= _zz_110_;
      end
      if(_zz_69_)begin
        int_reg_array_1_10_real <= _zz_110_;
      end
      if(_zz_70_)begin
        int_reg_array_1_11_real <= _zz_110_;
      end
      if(_zz_71_)begin
        int_reg_array_1_12_real <= _zz_110_;
      end
      if(_zz_72_)begin
        int_reg_array_1_13_real <= _zz_110_;
      end
      if(_zz_73_)begin
        int_reg_array_1_14_real <= _zz_110_;
      end
      if(_zz_74_)begin
        int_reg_array_1_15_real <= _zz_110_;
      end
      if(_zz_75_)begin
        int_reg_array_1_16_real <= _zz_110_;
      end
      if(_zz_76_)begin
        int_reg_array_1_17_real <= _zz_110_;
      end
      if(_zz_77_)begin
        int_reg_array_1_18_real <= _zz_110_;
      end
      if(_zz_78_)begin
        int_reg_array_1_19_real <= _zz_110_;
      end
      if(_zz_79_)begin
        int_reg_array_1_20_real <= _zz_110_;
      end
      if(_zz_80_)begin
        int_reg_array_1_21_real <= _zz_110_;
      end
      if(_zz_81_)begin
        int_reg_array_1_22_real <= _zz_110_;
      end
      if(_zz_82_)begin
        int_reg_array_1_23_real <= _zz_110_;
      end
      if(_zz_83_)begin
        int_reg_array_1_24_real <= _zz_110_;
      end
      if(_zz_84_)begin
        int_reg_array_1_25_real <= _zz_110_;
      end
      if(_zz_85_)begin
        int_reg_array_1_26_real <= _zz_110_;
      end
      if(_zz_86_)begin
        int_reg_array_1_27_real <= _zz_110_;
      end
      if(_zz_87_)begin
        int_reg_array_1_28_real <= _zz_110_;
      end
      if(_zz_88_)begin
        int_reg_array_1_29_real <= _zz_110_;
      end
      if(_zz_89_)begin
        int_reg_array_1_30_real <= _zz_110_;
      end
      if(_zz_90_)begin
        int_reg_array_1_31_real <= _zz_110_;
      end
      if(_zz_91_)begin
        int_reg_array_1_32_real <= _zz_110_;
      end
      if(_zz_92_)begin
        int_reg_array_1_33_real <= _zz_110_;
      end
      if(_zz_93_)begin
        int_reg_array_1_34_real <= _zz_110_;
      end
      if(_zz_94_)begin
        int_reg_array_1_35_real <= _zz_110_;
      end
      if(_zz_95_)begin
        int_reg_array_1_36_real <= _zz_110_;
      end
      if(_zz_96_)begin
        int_reg_array_1_37_real <= _zz_110_;
      end
      if(_zz_97_)begin
        int_reg_array_1_38_real <= _zz_110_;
      end
      if(_zz_98_)begin
        int_reg_array_1_39_real <= _zz_110_;
      end
      if(_zz_99_)begin
        int_reg_array_1_40_real <= _zz_110_;
      end
      if(_zz_100_)begin
        int_reg_array_1_41_real <= _zz_110_;
      end
      if(_zz_101_)begin
        int_reg_array_1_42_real <= _zz_110_;
      end
      if(_zz_102_)begin
        int_reg_array_1_43_real <= _zz_110_;
      end
      if(_zz_103_)begin
        int_reg_array_1_44_real <= _zz_110_;
      end
      if(_zz_104_)begin
        int_reg_array_1_45_real <= _zz_110_;
      end
      if(_zz_105_)begin
        int_reg_array_1_46_real <= _zz_110_;
      end
      if(_zz_106_)begin
        int_reg_array_1_47_real <= _zz_110_;
      end
      if(_zz_107_)begin
        int_reg_array_1_48_real <= _zz_110_;
      end
      if(_zz_108_)begin
        int_reg_array_1_49_real <= _zz_110_;
      end
      if(_zz_59_)begin
        int_reg_array_1_0_imag <= _zz_111_;
      end
      if(_zz_60_)begin
        int_reg_array_1_1_imag <= _zz_111_;
      end
      if(_zz_61_)begin
        int_reg_array_1_2_imag <= _zz_111_;
      end
      if(_zz_62_)begin
        int_reg_array_1_3_imag <= _zz_111_;
      end
      if(_zz_63_)begin
        int_reg_array_1_4_imag <= _zz_111_;
      end
      if(_zz_64_)begin
        int_reg_array_1_5_imag <= _zz_111_;
      end
      if(_zz_65_)begin
        int_reg_array_1_6_imag <= _zz_111_;
      end
      if(_zz_66_)begin
        int_reg_array_1_7_imag <= _zz_111_;
      end
      if(_zz_67_)begin
        int_reg_array_1_8_imag <= _zz_111_;
      end
      if(_zz_68_)begin
        int_reg_array_1_9_imag <= _zz_111_;
      end
      if(_zz_69_)begin
        int_reg_array_1_10_imag <= _zz_111_;
      end
      if(_zz_70_)begin
        int_reg_array_1_11_imag <= _zz_111_;
      end
      if(_zz_71_)begin
        int_reg_array_1_12_imag <= _zz_111_;
      end
      if(_zz_72_)begin
        int_reg_array_1_13_imag <= _zz_111_;
      end
      if(_zz_73_)begin
        int_reg_array_1_14_imag <= _zz_111_;
      end
      if(_zz_74_)begin
        int_reg_array_1_15_imag <= _zz_111_;
      end
      if(_zz_75_)begin
        int_reg_array_1_16_imag <= _zz_111_;
      end
      if(_zz_76_)begin
        int_reg_array_1_17_imag <= _zz_111_;
      end
      if(_zz_77_)begin
        int_reg_array_1_18_imag <= _zz_111_;
      end
      if(_zz_78_)begin
        int_reg_array_1_19_imag <= _zz_111_;
      end
      if(_zz_79_)begin
        int_reg_array_1_20_imag <= _zz_111_;
      end
      if(_zz_80_)begin
        int_reg_array_1_21_imag <= _zz_111_;
      end
      if(_zz_81_)begin
        int_reg_array_1_22_imag <= _zz_111_;
      end
      if(_zz_82_)begin
        int_reg_array_1_23_imag <= _zz_111_;
      end
      if(_zz_83_)begin
        int_reg_array_1_24_imag <= _zz_111_;
      end
      if(_zz_84_)begin
        int_reg_array_1_25_imag <= _zz_111_;
      end
      if(_zz_85_)begin
        int_reg_array_1_26_imag <= _zz_111_;
      end
      if(_zz_86_)begin
        int_reg_array_1_27_imag <= _zz_111_;
      end
      if(_zz_87_)begin
        int_reg_array_1_28_imag <= _zz_111_;
      end
      if(_zz_88_)begin
        int_reg_array_1_29_imag <= _zz_111_;
      end
      if(_zz_89_)begin
        int_reg_array_1_30_imag <= _zz_111_;
      end
      if(_zz_90_)begin
        int_reg_array_1_31_imag <= _zz_111_;
      end
      if(_zz_91_)begin
        int_reg_array_1_32_imag <= _zz_111_;
      end
      if(_zz_92_)begin
        int_reg_array_1_33_imag <= _zz_111_;
      end
      if(_zz_93_)begin
        int_reg_array_1_34_imag <= _zz_111_;
      end
      if(_zz_94_)begin
        int_reg_array_1_35_imag <= _zz_111_;
      end
      if(_zz_95_)begin
        int_reg_array_1_36_imag <= _zz_111_;
      end
      if(_zz_96_)begin
        int_reg_array_1_37_imag <= _zz_111_;
      end
      if(_zz_97_)begin
        int_reg_array_1_38_imag <= _zz_111_;
      end
      if(_zz_98_)begin
        int_reg_array_1_39_imag <= _zz_111_;
      end
      if(_zz_99_)begin
        int_reg_array_1_40_imag <= _zz_111_;
      end
      if(_zz_100_)begin
        int_reg_array_1_41_imag <= _zz_111_;
      end
      if(_zz_101_)begin
        int_reg_array_1_42_imag <= _zz_111_;
      end
      if(_zz_102_)begin
        int_reg_array_1_43_imag <= _zz_111_;
      end
      if(_zz_103_)begin
        int_reg_array_1_44_imag <= _zz_111_;
      end
      if(_zz_104_)begin
        int_reg_array_1_45_imag <= _zz_111_;
      end
      if(_zz_105_)begin
        int_reg_array_1_46_imag <= _zz_111_;
      end
      if(_zz_106_)begin
        int_reg_array_1_47_imag <= _zz_111_;
      end
      if(_zz_107_)begin
        int_reg_array_1_48_imag <= _zz_111_;
      end
      if(_zz_108_)begin
        int_reg_array_1_49_imag <= _zz_111_;
      end
      if(_zz_114_)begin
        int_reg_array_2_0_real <= _zz_165_;
      end
      if(_zz_115_)begin
        int_reg_array_2_1_real <= _zz_165_;
      end
      if(_zz_116_)begin
        int_reg_array_2_2_real <= _zz_165_;
      end
      if(_zz_117_)begin
        int_reg_array_2_3_real <= _zz_165_;
      end
      if(_zz_118_)begin
        int_reg_array_2_4_real <= _zz_165_;
      end
      if(_zz_119_)begin
        int_reg_array_2_5_real <= _zz_165_;
      end
      if(_zz_120_)begin
        int_reg_array_2_6_real <= _zz_165_;
      end
      if(_zz_121_)begin
        int_reg_array_2_7_real <= _zz_165_;
      end
      if(_zz_122_)begin
        int_reg_array_2_8_real <= _zz_165_;
      end
      if(_zz_123_)begin
        int_reg_array_2_9_real <= _zz_165_;
      end
      if(_zz_124_)begin
        int_reg_array_2_10_real <= _zz_165_;
      end
      if(_zz_125_)begin
        int_reg_array_2_11_real <= _zz_165_;
      end
      if(_zz_126_)begin
        int_reg_array_2_12_real <= _zz_165_;
      end
      if(_zz_127_)begin
        int_reg_array_2_13_real <= _zz_165_;
      end
      if(_zz_128_)begin
        int_reg_array_2_14_real <= _zz_165_;
      end
      if(_zz_129_)begin
        int_reg_array_2_15_real <= _zz_165_;
      end
      if(_zz_130_)begin
        int_reg_array_2_16_real <= _zz_165_;
      end
      if(_zz_131_)begin
        int_reg_array_2_17_real <= _zz_165_;
      end
      if(_zz_132_)begin
        int_reg_array_2_18_real <= _zz_165_;
      end
      if(_zz_133_)begin
        int_reg_array_2_19_real <= _zz_165_;
      end
      if(_zz_134_)begin
        int_reg_array_2_20_real <= _zz_165_;
      end
      if(_zz_135_)begin
        int_reg_array_2_21_real <= _zz_165_;
      end
      if(_zz_136_)begin
        int_reg_array_2_22_real <= _zz_165_;
      end
      if(_zz_137_)begin
        int_reg_array_2_23_real <= _zz_165_;
      end
      if(_zz_138_)begin
        int_reg_array_2_24_real <= _zz_165_;
      end
      if(_zz_139_)begin
        int_reg_array_2_25_real <= _zz_165_;
      end
      if(_zz_140_)begin
        int_reg_array_2_26_real <= _zz_165_;
      end
      if(_zz_141_)begin
        int_reg_array_2_27_real <= _zz_165_;
      end
      if(_zz_142_)begin
        int_reg_array_2_28_real <= _zz_165_;
      end
      if(_zz_143_)begin
        int_reg_array_2_29_real <= _zz_165_;
      end
      if(_zz_144_)begin
        int_reg_array_2_30_real <= _zz_165_;
      end
      if(_zz_145_)begin
        int_reg_array_2_31_real <= _zz_165_;
      end
      if(_zz_146_)begin
        int_reg_array_2_32_real <= _zz_165_;
      end
      if(_zz_147_)begin
        int_reg_array_2_33_real <= _zz_165_;
      end
      if(_zz_148_)begin
        int_reg_array_2_34_real <= _zz_165_;
      end
      if(_zz_149_)begin
        int_reg_array_2_35_real <= _zz_165_;
      end
      if(_zz_150_)begin
        int_reg_array_2_36_real <= _zz_165_;
      end
      if(_zz_151_)begin
        int_reg_array_2_37_real <= _zz_165_;
      end
      if(_zz_152_)begin
        int_reg_array_2_38_real <= _zz_165_;
      end
      if(_zz_153_)begin
        int_reg_array_2_39_real <= _zz_165_;
      end
      if(_zz_154_)begin
        int_reg_array_2_40_real <= _zz_165_;
      end
      if(_zz_155_)begin
        int_reg_array_2_41_real <= _zz_165_;
      end
      if(_zz_156_)begin
        int_reg_array_2_42_real <= _zz_165_;
      end
      if(_zz_157_)begin
        int_reg_array_2_43_real <= _zz_165_;
      end
      if(_zz_158_)begin
        int_reg_array_2_44_real <= _zz_165_;
      end
      if(_zz_159_)begin
        int_reg_array_2_45_real <= _zz_165_;
      end
      if(_zz_160_)begin
        int_reg_array_2_46_real <= _zz_165_;
      end
      if(_zz_161_)begin
        int_reg_array_2_47_real <= _zz_165_;
      end
      if(_zz_162_)begin
        int_reg_array_2_48_real <= _zz_165_;
      end
      if(_zz_163_)begin
        int_reg_array_2_49_real <= _zz_165_;
      end
      if(_zz_114_)begin
        int_reg_array_2_0_imag <= _zz_166_;
      end
      if(_zz_115_)begin
        int_reg_array_2_1_imag <= _zz_166_;
      end
      if(_zz_116_)begin
        int_reg_array_2_2_imag <= _zz_166_;
      end
      if(_zz_117_)begin
        int_reg_array_2_3_imag <= _zz_166_;
      end
      if(_zz_118_)begin
        int_reg_array_2_4_imag <= _zz_166_;
      end
      if(_zz_119_)begin
        int_reg_array_2_5_imag <= _zz_166_;
      end
      if(_zz_120_)begin
        int_reg_array_2_6_imag <= _zz_166_;
      end
      if(_zz_121_)begin
        int_reg_array_2_7_imag <= _zz_166_;
      end
      if(_zz_122_)begin
        int_reg_array_2_8_imag <= _zz_166_;
      end
      if(_zz_123_)begin
        int_reg_array_2_9_imag <= _zz_166_;
      end
      if(_zz_124_)begin
        int_reg_array_2_10_imag <= _zz_166_;
      end
      if(_zz_125_)begin
        int_reg_array_2_11_imag <= _zz_166_;
      end
      if(_zz_126_)begin
        int_reg_array_2_12_imag <= _zz_166_;
      end
      if(_zz_127_)begin
        int_reg_array_2_13_imag <= _zz_166_;
      end
      if(_zz_128_)begin
        int_reg_array_2_14_imag <= _zz_166_;
      end
      if(_zz_129_)begin
        int_reg_array_2_15_imag <= _zz_166_;
      end
      if(_zz_130_)begin
        int_reg_array_2_16_imag <= _zz_166_;
      end
      if(_zz_131_)begin
        int_reg_array_2_17_imag <= _zz_166_;
      end
      if(_zz_132_)begin
        int_reg_array_2_18_imag <= _zz_166_;
      end
      if(_zz_133_)begin
        int_reg_array_2_19_imag <= _zz_166_;
      end
      if(_zz_134_)begin
        int_reg_array_2_20_imag <= _zz_166_;
      end
      if(_zz_135_)begin
        int_reg_array_2_21_imag <= _zz_166_;
      end
      if(_zz_136_)begin
        int_reg_array_2_22_imag <= _zz_166_;
      end
      if(_zz_137_)begin
        int_reg_array_2_23_imag <= _zz_166_;
      end
      if(_zz_138_)begin
        int_reg_array_2_24_imag <= _zz_166_;
      end
      if(_zz_139_)begin
        int_reg_array_2_25_imag <= _zz_166_;
      end
      if(_zz_140_)begin
        int_reg_array_2_26_imag <= _zz_166_;
      end
      if(_zz_141_)begin
        int_reg_array_2_27_imag <= _zz_166_;
      end
      if(_zz_142_)begin
        int_reg_array_2_28_imag <= _zz_166_;
      end
      if(_zz_143_)begin
        int_reg_array_2_29_imag <= _zz_166_;
      end
      if(_zz_144_)begin
        int_reg_array_2_30_imag <= _zz_166_;
      end
      if(_zz_145_)begin
        int_reg_array_2_31_imag <= _zz_166_;
      end
      if(_zz_146_)begin
        int_reg_array_2_32_imag <= _zz_166_;
      end
      if(_zz_147_)begin
        int_reg_array_2_33_imag <= _zz_166_;
      end
      if(_zz_148_)begin
        int_reg_array_2_34_imag <= _zz_166_;
      end
      if(_zz_149_)begin
        int_reg_array_2_35_imag <= _zz_166_;
      end
      if(_zz_150_)begin
        int_reg_array_2_36_imag <= _zz_166_;
      end
      if(_zz_151_)begin
        int_reg_array_2_37_imag <= _zz_166_;
      end
      if(_zz_152_)begin
        int_reg_array_2_38_imag <= _zz_166_;
      end
      if(_zz_153_)begin
        int_reg_array_2_39_imag <= _zz_166_;
      end
      if(_zz_154_)begin
        int_reg_array_2_40_imag <= _zz_166_;
      end
      if(_zz_155_)begin
        int_reg_array_2_41_imag <= _zz_166_;
      end
      if(_zz_156_)begin
        int_reg_array_2_42_imag <= _zz_166_;
      end
      if(_zz_157_)begin
        int_reg_array_2_43_imag <= _zz_166_;
      end
      if(_zz_158_)begin
        int_reg_array_2_44_imag <= _zz_166_;
      end
      if(_zz_159_)begin
        int_reg_array_2_45_imag <= _zz_166_;
      end
      if(_zz_160_)begin
        int_reg_array_2_46_imag <= _zz_166_;
      end
      if(_zz_161_)begin
        int_reg_array_2_47_imag <= _zz_166_;
      end
      if(_zz_162_)begin
        int_reg_array_2_48_imag <= _zz_166_;
      end
      if(_zz_163_)begin
        int_reg_array_2_49_imag <= _zz_166_;
      end
      if(_zz_169_)begin
        int_reg_array_3_0_real <= _zz_220_;
      end
      if(_zz_170_)begin
        int_reg_array_3_1_real <= _zz_220_;
      end
      if(_zz_171_)begin
        int_reg_array_3_2_real <= _zz_220_;
      end
      if(_zz_172_)begin
        int_reg_array_3_3_real <= _zz_220_;
      end
      if(_zz_173_)begin
        int_reg_array_3_4_real <= _zz_220_;
      end
      if(_zz_174_)begin
        int_reg_array_3_5_real <= _zz_220_;
      end
      if(_zz_175_)begin
        int_reg_array_3_6_real <= _zz_220_;
      end
      if(_zz_176_)begin
        int_reg_array_3_7_real <= _zz_220_;
      end
      if(_zz_177_)begin
        int_reg_array_3_8_real <= _zz_220_;
      end
      if(_zz_178_)begin
        int_reg_array_3_9_real <= _zz_220_;
      end
      if(_zz_179_)begin
        int_reg_array_3_10_real <= _zz_220_;
      end
      if(_zz_180_)begin
        int_reg_array_3_11_real <= _zz_220_;
      end
      if(_zz_181_)begin
        int_reg_array_3_12_real <= _zz_220_;
      end
      if(_zz_182_)begin
        int_reg_array_3_13_real <= _zz_220_;
      end
      if(_zz_183_)begin
        int_reg_array_3_14_real <= _zz_220_;
      end
      if(_zz_184_)begin
        int_reg_array_3_15_real <= _zz_220_;
      end
      if(_zz_185_)begin
        int_reg_array_3_16_real <= _zz_220_;
      end
      if(_zz_186_)begin
        int_reg_array_3_17_real <= _zz_220_;
      end
      if(_zz_187_)begin
        int_reg_array_3_18_real <= _zz_220_;
      end
      if(_zz_188_)begin
        int_reg_array_3_19_real <= _zz_220_;
      end
      if(_zz_189_)begin
        int_reg_array_3_20_real <= _zz_220_;
      end
      if(_zz_190_)begin
        int_reg_array_3_21_real <= _zz_220_;
      end
      if(_zz_191_)begin
        int_reg_array_3_22_real <= _zz_220_;
      end
      if(_zz_192_)begin
        int_reg_array_3_23_real <= _zz_220_;
      end
      if(_zz_193_)begin
        int_reg_array_3_24_real <= _zz_220_;
      end
      if(_zz_194_)begin
        int_reg_array_3_25_real <= _zz_220_;
      end
      if(_zz_195_)begin
        int_reg_array_3_26_real <= _zz_220_;
      end
      if(_zz_196_)begin
        int_reg_array_3_27_real <= _zz_220_;
      end
      if(_zz_197_)begin
        int_reg_array_3_28_real <= _zz_220_;
      end
      if(_zz_198_)begin
        int_reg_array_3_29_real <= _zz_220_;
      end
      if(_zz_199_)begin
        int_reg_array_3_30_real <= _zz_220_;
      end
      if(_zz_200_)begin
        int_reg_array_3_31_real <= _zz_220_;
      end
      if(_zz_201_)begin
        int_reg_array_3_32_real <= _zz_220_;
      end
      if(_zz_202_)begin
        int_reg_array_3_33_real <= _zz_220_;
      end
      if(_zz_203_)begin
        int_reg_array_3_34_real <= _zz_220_;
      end
      if(_zz_204_)begin
        int_reg_array_3_35_real <= _zz_220_;
      end
      if(_zz_205_)begin
        int_reg_array_3_36_real <= _zz_220_;
      end
      if(_zz_206_)begin
        int_reg_array_3_37_real <= _zz_220_;
      end
      if(_zz_207_)begin
        int_reg_array_3_38_real <= _zz_220_;
      end
      if(_zz_208_)begin
        int_reg_array_3_39_real <= _zz_220_;
      end
      if(_zz_209_)begin
        int_reg_array_3_40_real <= _zz_220_;
      end
      if(_zz_210_)begin
        int_reg_array_3_41_real <= _zz_220_;
      end
      if(_zz_211_)begin
        int_reg_array_3_42_real <= _zz_220_;
      end
      if(_zz_212_)begin
        int_reg_array_3_43_real <= _zz_220_;
      end
      if(_zz_213_)begin
        int_reg_array_3_44_real <= _zz_220_;
      end
      if(_zz_214_)begin
        int_reg_array_3_45_real <= _zz_220_;
      end
      if(_zz_215_)begin
        int_reg_array_3_46_real <= _zz_220_;
      end
      if(_zz_216_)begin
        int_reg_array_3_47_real <= _zz_220_;
      end
      if(_zz_217_)begin
        int_reg_array_3_48_real <= _zz_220_;
      end
      if(_zz_218_)begin
        int_reg_array_3_49_real <= _zz_220_;
      end
      if(_zz_169_)begin
        int_reg_array_3_0_imag <= _zz_221_;
      end
      if(_zz_170_)begin
        int_reg_array_3_1_imag <= _zz_221_;
      end
      if(_zz_171_)begin
        int_reg_array_3_2_imag <= _zz_221_;
      end
      if(_zz_172_)begin
        int_reg_array_3_3_imag <= _zz_221_;
      end
      if(_zz_173_)begin
        int_reg_array_3_4_imag <= _zz_221_;
      end
      if(_zz_174_)begin
        int_reg_array_3_5_imag <= _zz_221_;
      end
      if(_zz_175_)begin
        int_reg_array_3_6_imag <= _zz_221_;
      end
      if(_zz_176_)begin
        int_reg_array_3_7_imag <= _zz_221_;
      end
      if(_zz_177_)begin
        int_reg_array_3_8_imag <= _zz_221_;
      end
      if(_zz_178_)begin
        int_reg_array_3_9_imag <= _zz_221_;
      end
      if(_zz_179_)begin
        int_reg_array_3_10_imag <= _zz_221_;
      end
      if(_zz_180_)begin
        int_reg_array_3_11_imag <= _zz_221_;
      end
      if(_zz_181_)begin
        int_reg_array_3_12_imag <= _zz_221_;
      end
      if(_zz_182_)begin
        int_reg_array_3_13_imag <= _zz_221_;
      end
      if(_zz_183_)begin
        int_reg_array_3_14_imag <= _zz_221_;
      end
      if(_zz_184_)begin
        int_reg_array_3_15_imag <= _zz_221_;
      end
      if(_zz_185_)begin
        int_reg_array_3_16_imag <= _zz_221_;
      end
      if(_zz_186_)begin
        int_reg_array_3_17_imag <= _zz_221_;
      end
      if(_zz_187_)begin
        int_reg_array_3_18_imag <= _zz_221_;
      end
      if(_zz_188_)begin
        int_reg_array_3_19_imag <= _zz_221_;
      end
      if(_zz_189_)begin
        int_reg_array_3_20_imag <= _zz_221_;
      end
      if(_zz_190_)begin
        int_reg_array_3_21_imag <= _zz_221_;
      end
      if(_zz_191_)begin
        int_reg_array_3_22_imag <= _zz_221_;
      end
      if(_zz_192_)begin
        int_reg_array_3_23_imag <= _zz_221_;
      end
      if(_zz_193_)begin
        int_reg_array_3_24_imag <= _zz_221_;
      end
      if(_zz_194_)begin
        int_reg_array_3_25_imag <= _zz_221_;
      end
      if(_zz_195_)begin
        int_reg_array_3_26_imag <= _zz_221_;
      end
      if(_zz_196_)begin
        int_reg_array_3_27_imag <= _zz_221_;
      end
      if(_zz_197_)begin
        int_reg_array_3_28_imag <= _zz_221_;
      end
      if(_zz_198_)begin
        int_reg_array_3_29_imag <= _zz_221_;
      end
      if(_zz_199_)begin
        int_reg_array_3_30_imag <= _zz_221_;
      end
      if(_zz_200_)begin
        int_reg_array_3_31_imag <= _zz_221_;
      end
      if(_zz_201_)begin
        int_reg_array_3_32_imag <= _zz_221_;
      end
      if(_zz_202_)begin
        int_reg_array_3_33_imag <= _zz_221_;
      end
      if(_zz_203_)begin
        int_reg_array_3_34_imag <= _zz_221_;
      end
      if(_zz_204_)begin
        int_reg_array_3_35_imag <= _zz_221_;
      end
      if(_zz_205_)begin
        int_reg_array_3_36_imag <= _zz_221_;
      end
      if(_zz_206_)begin
        int_reg_array_3_37_imag <= _zz_221_;
      end
      if(_zz_207_)begin
        int_reg_array_3_38_imag <= _zz_221_;
      end
      if(_zz_208_)begin
        int_reg_array_3_39_imag <= _zz_221_;
      end
      if(_zz_209_)begin
        int_reg_array_3_40_imag <= _zz_221_;
      end
      if(_zz_210_)begin
        int_reg_array_3_41_imag <= _zz_221_;
      end
      if(_zz_211_)begin
        int_reg_array_3_42_imag <= _zz_221_;
      end
      if(_zz_212_)begin
        int_reg_array_3_43_imag <= _zz_221_;
      end
      if(_zz_213_)begin
        int_reg_array_3_44_imag <= _zz_221_;
      end
      if(_zz_214_)begin
        int_reg_array_3_45_imag <= _zz_221_;
      end
      if(_zz_215_)begin
        int_reg_array_3_46_imag <= _zz_221_;
      end
      if(_zz_216_)begin
        int_reg_array_3_47_imag <= _zz_221_;
      end
      if(_zz_217_)begin
        int_reg_array_3_48_imag <= _zz_221_;
      end
      if(_zz_218_)begin
        int_reg_array_3_49_imag <= _zz_221_;
      end
      if(_zz_224_)begin
        int_reg_array_4_0_real <= _zz_275_;
      end
      if(_zz_225_)begin
        int_reg_array_4_1_real <= _zz_275_;
      end
      if(_zz_226_)begin
        int_reg_array_4_2_real <= _zz_275_;
      end
      if(_zz_227_)begin
        int_reg_array_4_3_real <= _zz_275_;
      end
      if(_zz_228_)begin
        int_reg_array_4_4_real <= _zz_275_;
      end
      if(_zz_229_)begin
        int_reg_array_4_5_real <= _zz_275_;
      end
      if(_zz_230_)begin
        int_reg_array_4_6_real <= _zz_275_;
      end
      if(_zz_231_)begin
        int_reg_array_4_7_real <= _zz_275_;
      end
      if(_zz_232_)begin
        int_reg_array_4_8_real <= _zz_275_;
      end
      if(_zz_233_)begin
        int_reg_array_4_9_real <= _zz_275_;
      end
      if(_zz_234_)begin
        int_reg_array_4_10_real <= _zz_275_;
      end
      if(_zz_235_)begin
        int_reg_array_4_11_real <= _zz_275_;
      end
      if(_zz_236_)begin
        int_reg_array_4_12_real <= _zz_275_;
      end
      if(_zz_237_)begin
        int_reg_array_4_13_real <= _zz_275_;
      end
      if(_zz_238_)begin
        int_reg_array_4_14_real <= _zz_275_;
      end
      if(_zz_239_)begin
        int_reg_array_4_15_real <= _zz_275_;
      end
      if(_zz_240_)begin
        int_reg_array_4_16_real <= _zz_275_;
      end
      if(_zz_241_)begin
        int_reg_array_4_17_real <= _zz_275_;
      end
      if(_zz_242_)begin
        int_reg_array_4_18_real <= _zz_275_;
      end
      if(_zz_243_)begin
        int_reg_array_4_19_real <= _zz_275_;
      end
      if(_zz_244_)begin
        int_reg_array_4_20_real <= _zz_275_;
      end
      if(_zz_245_)begin
        int_reg_array_4_21_real <= _zz_275_;
      end
      if(_zz_246_)begin
        int_reg_array_4_22_real <= _zz_275_;
      end
      if(_zz_247_)begin
        int_reg_array_4_23_real <= _zz_275_;
      end
      if(_zz_248_)begin
        int_reg_array_4_24_real <= _zz_275_;
      end
      if(_zz_249_)begin
        int_reg_array_4_25_real <= _zz_275_;
      end
      if(_zz_250_)begin
        int_reg_array_4_26_real <= _zz_275_;
      end
      if(_zz_251_)begin
        int_reg_array_4_27_real <= _zz_275_;
      end
      if(_zz_252_)begin
        int_reg_array_4_28_real <= _zz_275_;
      end
      if(_zz_253_)begin
        int_reg_array_4_29_real <= _zz_275_;
      end
      if(_zz_254_)begin
        int_reg_array_4_30_real <= _zz_275_;
      end
      if(_zz_255_)begin
        int_reg_array_4_31_real <= _zz_275_;
      end
      if(_zz_256_)begin
        int_reg_array_4_32_real <= _zz_275_;
      end
      if(_zz_257_)begin
        int_reg_array_4_33_real <= _zz_275_;
      end
      if(_zz_258_)begin
        int_reg_array_4_34_real <= _zz_275_;
      end
      if(_zz_259_)begin
        int_reg_array_4_35_real <= _zz_275_;
      end
      if(_zz_260_)begin
        int_reg_array_4_36_real <= _zz_275_;
      end
      if(_zz_261_)begin
        int_reg_array_4_37_real <= _zz_275_;
      end
      if(_zz_262_)begin
        int_reg_array_4_38_real <= _zz_275_;
      end
      if(_zz_263_)begin
        int_reg_array_4_39_real <= _zz_275_;
      end
      if(_zz_264_)begin
        int_reg_array_4_40_real <= _zz_275_;
      end
      if(_zz_265_)begin
        int_reg_array_4_41_real <= _zz_275_;
      end
      if(_zz_266_)begin
        int_reg_array_4_42_real <= _zz_275_;
      end
      if(_zz_267_)begin
        int_reg_array_4_43_real <= _zz_275_;
      end
      if(_zz_268_)begin
        int_reg_array_4_44_real <= _zz_275_;
      end
      if(_zz_269_)begin
        int_reg_array_4_45_real <= _zz_275_;
      end
      if(_zz_270_)begin
        int_reg_array_4_46_real <= _zz_275_;
      end
      if(_zz_271_)begin
        int_reg_array_4_47_real <= _zz_275_;
      end
      if(_zz_272_)begin
        int_reg_array_4_48_real <= _zz_275_;
      end
      if(_zz_273_)begin
        int_reg_array_4_49_real <= _zz_275_;
      end
      if(_zz_224_)begin
        int_reg_array_4_0_imag <= _zz_276_;
      end
      if(_zz_225_)begin
        int_reg_array_4_1_imag <= _zz_276_;
      end
      if(_zz_226_)begin
        int_reg_array_4_2_imag <= _zz_276_;
      end
      if(_zz_227_)begin
        int_reg_array_4_3_imag <= _zz_276_;
      end
      if(_zz_228_)begin
        int_reg_array_4_4_imag <= _zz_276_;
      end
      if(_zz_229_)begin
        int_reg_array_4_5_imag <= _zz_276_;
      end
      if(_zz_230_)begin
        int_reg_array_4_6_imag <= _zz_276_;
      end
      if(_zz_231_)begin
        int_reg_array_4_7_imag <= _zz_276_;
      end
      if(_zz_232_)begin
        int_reg_array_4_8_imag <= _zz_276_;
      end
      if(_zz_233_)begin
        int_reg_array_4_9_imag <= _zz_276_;
      end
      if(_zz_234_)begin
        int_reg_array_4_10_imag <= _zz_276_;
      end
      if(_zz_235_)begin
        int_reg_array_4_11_imag <= _zz_276_;
      end
      if(_zz_236_)begin
        int_reg_array_4_12_imag <= _zz_276_;
      end
      if(_zz_237_)begin
        int_reg_array_4_13_imag <= _zz_276_;
      end
      if(_zz_238_)begin
        int_reg_array_4_14_imag <= _zz_276_;
      end
      if(_zz_239_)begin
        int_reg_array_4_15_imag <= _zz_276_;
      end
      if(_zz_240_)begin
        int_reg_array_4_16_imag <= _zz_276_;
      end
      if(_zz_241_)begin
        int_reg_array_4_17_imag <= _zz_276_;
      end
      if(_zz_242_)begin
        int_reg_array_4_18_imag <= _zz_276_;
      end
      if(_zz_243_)begin
        int_reg_array_4_19_imag <= _zz_276_;
      end
      if(_zz_244_)begin
        int_reg_array_4_20_imag <= _zz_276_;
      end
      if(_zz_245_)begin
        int_reg_array_4_21_imag <= _zz_276_;
      end
      if(_zz_246_)begin
        int_reg_array_4_22_imag <= _zz_276_;
      end
      if(_zz_247_)begin
        int_reg_array_4_23_imag <= _zz_276_;
      end
      if(_zz_248_)begin
        int_reg_array_4_24_imag <= _zz_276_;
      end
      if(_zz_249_)begin
        int_reg_array_4_25_imag <= _zz_276_;
      end
      if(_zz_250_)begin
        int_reg_array_4_26_imag <= _zz_276_;
      end
      if(_zz_251_)begin
        int_reg_array_4_27_imag <= _zz_276_;
      end
      if(_zz_252_)begin
        int_reg_array_4_28_imag <= _zz_276_;
      end
      if(_zz_253_)begin
        int_reg_array_4_29_imag <= _zz_276_;
      end
      if(_zz_254_)begin
        int_reg_array_4_30_imag <= _zz_276_;
      end
      if(_zz_255_)begin
        int_reg_array_4_31_imag <= _zz_276_;
      end
      if(_zz_256_)begin
        int_reg_array_4_32_imag <= _zz_276_;
      end
      if(_zz_257_)begin
        int_reg_array_4_33_imag <= _zz_276_;
      end
      if(_zz_258_)begin
        int_reg_array_4_34_imag <= _zz_276_;
      end
      if(_zz_259_)begin
        int_reg_array_4_35_imag <= _zz_276_;
      end
      if(_zz_260_)begin
        int_reg_array_4_36_imag <= _zz_276_;
      end
      if(_zz_261_)begin
        int_reg_array_4_37_imag <= _zz_276_;
      end
      if(_zz_262_)begin
        int_reg_array_4_38_imag <= _zz_276_;
      end
      if(_zz_263_)begin
        int_reg_array_4_39_imag <= _zz_276_;
      end
      if(_zz_264_)begin
        int_reg_array_4_40_imag <= _zz_276_;
      end
      if(_zz_265_)begin
        int_reg_array_4_41_imag <= _zz_276_;
      end
      if(_zz_266_)begin
        int_reg_array_4_42_imag <= _zz_276_;
      end
      if(_zz_267_)begin
        int_reg_array_4_43_imag <= _zz_276_;
      end
      if(_zz_268_)begin
        int_reg_array_4_44_imag <= _zz_276_;
      end
      if(_zz_269_)begin
        int_reg_array_4_45_imag <= _zz_276_;
      end
      if(_zz_270_)begin
        int_reg_array_4_46_imag <= _zz_276_;
      end
      if(_zz_271_)begin
        int_reg_array_4_47_imag <= _zz_276_;
      end
      if(_zz_272_)begin
        int_reg_array_4_48_imag <= _zz_276_;
      end
      if(_zz_273_)begin
        int_reg_array_4_49_imag <= _zz_276_;
      end
      if(_zz_279_)begin
        int_reg_array_5_0_real <= _zz_330_;
      end
      if(_zz_280_)begin
        int_reg_array_5_1_real <= _zz_330_;
      end
      if(_zz_281_)begin
        int_reg_array_5_2_real <= _zz_330_;
      end
      if(_zz_282_)begin
        int_reg_array_5_3_real <= _zz_330_;
      end
      if(_zz_283_)begin
        int_reg_array_5_4_real <= _zz_330_;
      end
      if(_zz_284_)begin
        int_reg_array_5_5_real <= _zz_330_;
      end
      if(_zz_285_)begin
        int_reg_array_5_6_real <= _zz_330_;
      end
      if(_zz_286_)begin
        int_reg_array_5_7_real <= _zz_330_;
      end
      if(_zz_287_)begin
        int_reg_array_5_8_real <= _zz_330_;
      end
      if(_zz_288_)begin
        int_reg_array_5_9_real <= _zz_330_;
      end
      if(_zz_289_)begin
        int_reg_array_5_10_real <= _zz_330_;
      end
      if(_zz_290_)begin
        int_reg_array_5_11_real <= _zz_330_;
      end
      if(_zz_291_)begin
        int_reg_array_5_12_real <= _zz_330_;
      end
      if(_zz_292_)begin
        int_reg_array_5_13_real <= _zz_330_;
      end
      if(_zz_293_)begin
        int_reg_array_5_14_real <= _zz_330_;
      end
      if(_zz_294_)begin
        int_reg_array_5_15_real <= _zz_330_;
      end
      if(_zz_295_)begin
        int_reg_array_5_16_real <= _zz_330_;
      end
      if(_zz_296_)begin
        int_reg_array_5_17_real <= _zz_330_;
      end
      if(_zz_297_)begin
        int_reg_array_5_18_real <= _zz_330_;
      end
      if(_zz_298_)begin
        int_reg_array_5_19_real <= _zz_330_;
      end
      if(_zz_299_)begin
        int_reg_array_5_20_real <= _zz_330_;
      end
      if(_zz_300_)begin
        int_reg_array_5_21_real <= _zz_330_;
      end
      if(_zz_301_)begin
        int_reg_array_5_22_real <= _zz_330_;
      end
      if(_zz_302_)begin
        int_reg_array_5_23_real <= _zz_330_;
      end
      if(_zz_303_)begin
        int_reg_array_5_24_real <= _zz_330_;
      end
      if(_zz_304_)begin
        int_reg_array_5_25_real <= _zz_330_;
      end
      if(_zz_305_)begin
        int_reg_array_5_26_real <= _zz_330_;
      end
      if(_zz_306_)begin
        int_reg_array_5_27_real <= _zz_330_;
      end
      if(_zz_307_)begin
        int_reg_array_5_28_real <= _zz_330_;
      end
      if(_zz_308_)begin
        int_reg_array_5_29_real <= _zz_330_;
      end
      if(_zz_309_)begin
        int_reg_array_5_30_real <= _zz_330_;
      end
      if(_zz_310_)begin
        int_reg_array_5_31_real <= _zz_330_;
      end
      if(_zz_311_)begin
        int_reg_array_5_32_real <= _zz_330_;
      end
      if(_zz_312_)begin
        int_reg_array_5_33_real <= _zz_330_;
      end
      if(_zz_313_)begin
        int_reg_array_5_34_real <= _zz_330_;
      end
      if(_zz_314_)begin
        int_reg_array_5_35_real <= _zz_330_;
      end
      if(_zz_315_)begin
        int_reg_array_5_36_real <= _zz_330_;
      end
      if(_zz_316_)begin
        int_reg_array_5_37_real <= _zz_330_;
      end
      if(_zz_317_)begin
        int_reg_array_5_38_real <= _zz_330_;
      end
      if(_zz_318_)begin
        int_reg_array_5_39_real <= _zz_330_;
      end
      if(_zz_319_)begin
        int_reg_array_5_40_real <= _zz_330_;
      end
      if(_zz_320_)begin
        int_reg_array_5_41_real <= _zz_330_;
      end
      if(_zz_321_)begin
        int_reg_array_5_42_real <= _zz_330_;
      end
      if(_zz_322_)begin
        int_reg_array_5_43_real <= _zz_330_;
      end
      if(_zz_323_)begin
        int_reg_array_5_44_real <= _zz_330_;
      end
      if(_zz_324_)begin
        int_reg_array_5_45_real <= _zz_330_;
      end
      if(_zz_325_)begin
        int_reg_array_5_46_real <= _zz_330_;
      end
      if(_zz_326_)begin
        int_reg_array_5_47_real <= _zz_330_;
      end
      if(_zz_327_)begin
        int_reg_array_5_48_real <= _zz_330_;
      end
      if(_zz_328_)begin
        int_reg_array_5_49_real <= _zz_330_;
      end
      if(_zz_279_)begin
        int_reg_array_5_0_imag <= _zz_331_;
      end
      if(_zz_280_)begin
        int_reg_array_5_1_imag <= _zz_331_;
      end
      if(_zz_281_)begin
        int_reg_array_5_2_imag <= _zz_331_;
      end
      if(_zz_282_)begin
        int_reg_array_5_3_imag <= _zz_331_;
      end
      if(_zz_283_)begin
        int_reg_array_5_4_imag <= _zz_331_;
      end
      if(_zz_284_)begin
        int_reg_array_5_5_imag <= _zz_331_;
      end
      if(_zz_285_)begin
        int_reg_array_5_6_imag <= _zz_331_;
      end
      if(_zz_286_)begin
        int_reg_array_5_7_imag <= _zz_331_;
      end
      if(_zz_287_)begin
        int_reg_array_5_8_imag <= _zz_331_;
      end
      if(_zz_288_)begin
        int_reg_array_5_9_imag <= _zz_331_;
      end
      if(_zz_289_)begin
        int_reg_array_5_10_imag <= _zz_331_;
      end
      if(_zz_290_)begin
        int_reg_array_5_11_imag <= _zz_331_;
      end
      if(_zz_291_)begin
        int_reg_array_5_12_imag <= _zz_331_;
      end
      if(_zz_292_)begin
        int_reg_array_5_13_imag <= _zz_331_;
      end
      if(_zz_293_)begin
        int_reg_array_5_14_imag <= _zz_331_;
      end
      if(_zz_294_)begin
        int_reg_array_5_15_imag <= _zz_331_;
      end
      if(_zz_295_)begin
        int_reg_array_5_16_imag <= _zz_331_;
      end
      if(_zz_296_)begin
        int_reg_array_5_17_imag <= _zz_331_;
      end
      if(_zz_297_)begin
        int_reg_array_5_18_imag <= _zz_331_;
      end
      if(_zz_298_)begin
        int_reg_array_5_19_imag <= _zz_331_;
      end
      if(_zz_299_)begin
        int_reg_array_5_20_imag <= _zz_331_;
      end
      if(_zz_300_)begin
        int_reg_array_5_21_imag <= _zz_331_;
      end
      if(_zz_301_)begin
        int_reg_array_5_22_imag <= _zz_331_;
      end
      if(_zz_302_)begin
        int_reg_array_5_23_imag <= _zz_331_;
      end
      if(_zz_303_)begin
        int_reg_array_5_24_imag <= _zz_331_;
      end
      if(_zz_304_)begin
        int_reg_array_5_25_imag <= _zz_331_;
      end
      if(_zz_305_)begin
        int_reg_array_5_26_imag <= _zz_331_;
      end
      if(_zz_306_)begin
        int_reg_array_5_27_imag <= _zz_331_;
      end
      if(_zz_307_)begin
        int_reg_array_5_28_imag <= _zz_331_;
      end
      if(_zz_308_)begin
        int_reg_array_5_29_imag <= _zz_331_;
      end
      if(_zz_309_)begin
        int_reg_array_5_30_imag <= _zz_331_;
      end
      if(_zz_310_)begin
        int_reg_array_5_31_imag <= _zz_331_;
      end
      if(_zz_311_)begin
        int_reg_array_5_32_imag <= _zz_331_;
      end
      if(_zz_312_)begin
        int_reg_array_5_33_imag <= _zz_331_;
      end
      if(_zz_313_)begin
        int_reg_array_5_34_imag <= _zz_331_;
      end
      if(_zz_314_)begin
        int_reg_array_5_35_imag <= _zz_331_;
      end
      if(_zz_315_)begin
        int_reg_array_5_36_imag <= _zz_331_;
      end
      if(_zz_316_)begin
        int_reg_array_5_37_imag <= _zz_331_;
      end
      if(_zz_317_)begin
        int_reg_array_5_38_imag <= _zz_331_;
      end
      if(_zz_318_)begin
        int_reg_array_5_39_imag <= _zz_331_;
      end
      if(_zz_319_)begin
        int_reg_array_5_40_imag <= _zz_331_;
      end
      if(_zz_320_)begin
        int_reg_array_5_41_imag <= _zz_331_;
      end
      if(_zz_321_)begin
        int_reg_array_5_42_imag <= _zz_331_;
      end
      if(_zz_322_)begin
        int_reg_array_5_43_imag <= _zz_331_;
      end
      if(_zz_323_)begin
        int_reg_array_5_44_imag <= _zz_331_;
      end
      if(_zz_324_)begin
        int_reg_array_5_45_imag <= _zz_331_;
      end
      if(_zz_325_)begin
        int_reg_array_5_46_imag <= _zz_331_;
      end
      if(_zz_326_)begin
        int_reg_array_5_47_imag <= _zz_331_;
      end
      if(_zz_327_)begin
        int_reg_array_5_48_imag <= _zz_331_;
      end
      if(_zz_328_)begin
        int_reg_array_5_49_imag <= _zz_331_;
      end
      if(_zz_334_)begin
        int_reg_array_6_0_real <= _zz_385_;
      end
      if(_zz_335_)begin
        int_reg_array_6_1_real <= _zz_385_;
      end
      if(_zz_336_)begin
        int_reg_array_6_2_real <= _zz_385_;
      end
      if(_zz_337_)begin
        int_reg_array_6_3_real <= _zz_385_;
      end
      if(_zz_338_)begin
        int_reg_array_6_4_real <= _zz_385_;
      end
      if(_zz_339_)begin
        int_reg_array_6_5_real <= _zz_385_;
      end
      if(_zz_340_)begin
        int_reg_array_6_6_real <= _zz_385_;
      end
      if(_zz_341_)begin
        int_reg_array_6_7_real <= _zz_385_;
      end
      if(_zz_342_)begin
        int_reg_array_6_8_real <= _zz_385_;
      end
      if(_zz_343_)begin
        int_reg_array_6_9_real <= _zz_385_;
      end
      if(_zz_344_)begin
        int_reg_array_6_10_real <= _zz_385_;
      end
      if(_zz_345_)begin
        int_reg_array_6_11_real <= _zz_385_;
      end
      if(_zz_346_)begin
        int_reg_array_6_12_real <= _zz_385_;
      end
      if(_zz_347_)begin
        int_reg_array_6_13_real <= _zz_385_;
      end
      if(_zz_348_)begin
        int_reg_array_6_14_real <= _zz_385_;
      end
      if(_zz_349_)begin
        int_reg_array_6_15_real <= _zz_385_;
      end
      if(_zz_350_)begin
        int_reg_array_6_16_real <= _zz_385_;
      end
      if(_zz_351_)begin
        int_reg_array_6_17_real <= _zz_385_;
      end
      if(_zz_352_)begin
        int_reg_array_6_18_real <= _zz_385_;
      end
      if(_zz_353_)begin
        int_reg_array_6_19_real <= _zz_385_;
      end
      if(_zz_354_)begin
        int_reg_array_6_20_real <= _zz_385_;
      end
      if(_zz_355_)begin
        int_reg_array_6_21_real <= _zz_385_;
      end
      if(_zz_356_)begin
        int_reg_array_6_22_real <= _zz_385_;
      end
      if(_zz_357_)begin
        int_reg_array_6_23_real <= _zz_385_;
      end
      if(_zz_358_)begin
        int_reg_array_6_24_real <= _zz_385_;
      end
      if(_zz_359_)begin
        int_reg_array_6_25_real <= _zz_385_;
      end
      if(_zz_360_)begin
        int_reg_array_6_26_real <= _zz_385_;
      end
      if(_zz_361_)begin
        int_reg_array_6_27_real <= _zz_385_;
      end
      if(_zz_362_)begin
        int_reg_array_6_28_real <= _zz_385_;
      end
      if(_zz_363_)begin
        int_reg_array_6_29_real <= _zz_385_;
      end
      if(_zz_364_)begin
        int_reg_array_6_30_real <= _zz_385_;
      end
      if(_zz_365_)begin
        int_reg_array_6_31_real <= _zz_385_;
      end
      if(_zz_366_)begin
        int_reg_array_6_32_real <= _zz_385_;
      end
      if(_zz_367_)begin
        int_reg_array_6_33_real <= _zz_385_;
      end
      if(_zz_368_)begin
        int_reg_array_6_34_real <= _zz_385_;
      end
      if(_zz_369_)begin
        int_reg_array_6_35_real <= _zz_385_;
      end
      if(_zz_370_)begin
        int_reg_array_6_36_real <= _zz_385_;
      end
      if(_zz_371_)begin
        int_reg_array_6_37_real <= _zz_385_;
      end
      if(_zz_372_)begin
        int_reg_array_6_38_real <= _zz_385_;
      end
      if(_zz_373_)begin
        int_reg_array_6_39_real <= _zz_385_;
      end
      if(_zz_374_)begin
        int_reg_array_6_40_real <= _zz_385_;
      end
      if(_zz_375_)begin
        int_reg_array_6_41_real <= _zz_385_;
      end
      if(_zz_376_)begin
        int_reg_array_6_42_real <= _zz_385_;
      end
      if(_zz_377_)begin
        int_reg_array_6_43_real <= _zz_385_;
      end
      if(_zz_378_)begin
        int_reg_array_6_44_real <= _zz_385_;
      end
      if(_zz_379_)begin
        int_reg_array_6_45_real <= _zz_385_;
      end
      if(_zz_380_)begin
        int_reg_array_6_46_real <= _zz_385_;
      end
      if(_zz_381_)begin
        int_reg_array_6_47_real <= _zz_385_;
      end
      if(_zz_382_)begin
        int_reg_array_6_48_real <= _zz_385_;
      end
      if(_zz_383_)begin
        int_reg_array_6_49_real <= _zz_385_;
      end
      if(_zz_334_)begin
        int_reg_array_6_0_imag <= _zz_386_;
      end
      if(_zz_335_)begin
        int_reg_array_6_1_imag <= _zz_386_;
      end
      if(_zz_336_)begin
        int_reg_array_6_2_imag <= _zz_386_;
      end
      if(_zz_337_)begin
        int_reg_array_6_3_imag <= _zz_386_;
      end
      if(_zz_338_)begin
        int_reg_array_6_4_imag <= _zz_386_;
      end
      if(_zz_339_)begin
        int_reg_array_6_5_imag <= _zz_386_;
      end
      if(_zz_340_)begin
        int_reg_array_6_6_imag <= _zz_386_;
      end
      if(_zz_341_)begin
        int_reg_array_6_7_imag <= _zz_386_;
      end
      if(_zz_342_)begin
        int_reg_array_6_8_imag <= _zz_386_;
      end
      if(_zz_343_)begin
        int_reg_array_6_9_imag <= _zz_386_;
      end
      if(_zz_344_)begin
        int_reg_array_6_10_imag <= _zz_386_;
      end
      if(_zz_345_)begin
        int_reg_array_6_11_imag <= _zz_386_;
      end
      if(_zz_346_)begin
        int_reg_array_6_12_imag <= _zz_386_;
      end
      if(_zz_347_)begin
        int_reg_array_6_13_imag <= _zz_386_;
      end
      if(_zz_348_)begin
        int_reg_array_6_14_imag <= _zz_386_;
      end
      if(_zz_349_)begin
        int_reg_array_6_15_imag <= _zz_386_;
      end
      if(_zz_350_)begin
        int_reg_array_6_16_imag <= _zz_386_;
      end
      if(_zz_351_)begin
        int_reg_array_6_17_imag <= _zz_386_;
      end
      if(_zz_352_)begin
        int_reg_array_6_18_imag <= _zz_386_;
      end
      if(_zz_353_)begin
        int_reg_array_6_19_imag <= _zz_386_;
      end
      if(_zz_354_)begin
        int_reg_array_6_20_imag <= _zz_386_;
      end
      if(_zz_355_)begin
        int_reg_array_6_21_imag <= _zz_386_;
      end
      if(_zz_356_)begin
        int_reg_array_6_22_imag <= _zz_386_;
      end
      if(_zz_357_)begin
        int_reg_array_6_23_imag <= _zz_386_;
      end
      if(_zz_358_)begin
        int_reg_array_6_24_imag <= _zz_386_;
      end
      if(_zz_359_)begin
        int_reg_array_6_25_imag <= _zz_386_;
      end
      if(_zz_360_)begin
        int_reg_array_6_26_imag <= _zz_386_;
      end
      if(_zz_361_)begin
        int_reg_array_6_27_imag <= _zz_386_;
      end
      if(_zz_362_)begin
        int_reg_array_6_28_imag <= _zz_386_;
      end
      if(_zz_363_)begin
        int_reg_array_6_29_imag <= _zz_386_;
      end
      if(_zz_364_)begin
        int_reg_array_6_30_imag <= _zz_386_;
      end
      if(_zz_365_)begin
        int_reg_array_6_31_imag <= _zz_386_;
      end
      if(_zz_366_)begin
        int_reg_array_6_32_imag <= _zz_386_;
      end
      if(_zz_367_)begin
        int_reg_array_6_33_imag <= _zz_386_;
      end
      if(_zz_368_)begin
        int_reg_array_6_34_imag <= _zz_386_;
      end
      if(_zz_369_)begin
        int_reg_array_6_35_imag <= _zz_386_;
      end
      if(_zz_370_)begin
        int_reg_array_6_36_imag <= _zz_386_;
      end
      if(_zz_371_)begin
        int_reg_array_6_37_imag <= _zz_386_;
      end
      if(_zz_372_)begin
        int_reg_array_6_38_imag <= _zz_386_;
      end
      if(_zz_373_)begin
        int_reg_array_6_39_imag <= _zz_386_;
      end
      if(_zz_374_)begin
        int_reg_array_6_40_imag <= _zz_386_;
      end
      if(_zz_375_)begin
        int_reg_array_6_41_imag <= _zz_386_;
      end
      if(_zz_376_)begin
        int_reg_array_6_42_imag <= _zz_386_;
      end
      if(_zz_377_)begin
        int_reg_array_6_43_imag <= _zz_386_;
      end
      if(_zz_378_)begin
        int_reg_array_6_44_imag <= _zz_386_;
      end
      if(_zz_379_)begin
        int_reg_array_6_45_imag <= _zz_386_;
      end
      if(_zz_380_)begin
        int_reg_array_6_46_imag <= _zz_386_;
      end
      if(_zz_381_)begin
        int_reg_array_6_47_imag <= _zz_386_;
      end
      if(_zz_382_)begin
        int_reg_array_6_48_imag <= _zz_386_;
      end
      if(_zz_383_)begin
        int_reg_array_6_49_imag <= _zz_386_;
      end
      if(_zz_389_)begin
        int_reg_array_7_0_real <= _zz_440_;
      end
      if(_zz_390_)begin
        int_reg_array_7_1_real <= _zz_440_;
      end
      if(_zz_391_)begin
        int_reg_array_7_2_real <= _zz_440_;
      end
      if(_zz_392_)begin
        int_reg_array_7_3_real <= _zz_440_;
      end
      if(_zz_393_)begin
        int_reg_array_7_4_real <= _zz_440_;
      end
      if(_zz_394_)begin
        int_reg_array_7_5_real <= _zz_440_;
      end
      if(_zz_395_)begin
        int_reg_array_7_6_real <= _zz_440_;
      end
      if(_zz_396_)begin
        int_reg_array_7_7_real <= _zz_440_;
      end
      if(_zz_397_)begin
        int_reg_array_7_8_real <= _zz_440_;
      end
      if(_zz_398_)begin
        int_reg_array_7_9_real <= _zz_440_;
      end
      if(_zz_399_)begin
        int_reg_array_7_10_real <= _zz_440_;
      end
      if(_zz_400_)begin
        int_reg_array_7_11_real <= _zz_440_;
      end
      if(_zz_401_)begin
        int_reg_array_7_12_real <= _zz_440_;
      end
      if(_zz_402_)begin
        int_reg_array_7_13_real <= _zz_440_;
      end
      if(_zz_403_)begin
        int_reg_array_7_14_real <= _zz_440_;
      end
      if(_zz_404_)begin
        int_reg_array_7_15_real <= _zz_440_;
      end
      if(_zz_405_)begin
        int_reg_array_7_16_real <= _zz_440_;
      end
      if(_zz_406_)begin
        int_reg_array_7_17_real <= _zz_440_;
      end
      if(_zz_407_)begin
        int_reg_array_7_18_real <= _zz_440_;
      end
      if(_zz_408_)begin
        int_reg_array_7_19_real <= _zz_440_;
      end
      if(_zz_409_)begin
        int_reg_array_7_20_real <= _zz_440_;
      end
      if(_zz_410_)begin
        int_reg_array_7_21_real <= _zz_440_;
      end
      if(_zz_411_)begin
        int_reg_array_7_22_real <= _zz_440_;
      end
      if(_zz_412_)begin
        int_reg_array_7_23_real <= _zz_440_;
      end
      if(_zz_413_)begin
        int_reg_array_7_24_real <= _zz_440_;
      end
      if(_zz_414_)begin
        int_reg_array_7_25_real <= _zz_440_;
      end
      if(_zz_415_)begin
        int_reg_array_7_26_real <= _zz_440_;
      end
      if(_zz_416_)begin
        int_reg_array_7_27_real <= _zz_440_;
      end
      if(_zz_417_)begin
        int_reg_array_7_28_real <= _zz_440_;
      end
      if(_zz_418_)begin
        int_reg_array_7_29_real <= _zz_440_;
      end
      if(_zz_419_)begin
        int_reg_array_7_30_real <= _zz_440_;
      end
      if(_zz_420_)begin
        int_reg_array_7_31_real <= _zz_440_;
      end
      if(_zz_421_)begin
        int_reg_array_7_32_real <= _zz_440_;
      end
      if(_zz_422_)begin
        int_reg_array_7_33_real <= _zz_440_;
      end
      if(_zz_423_)begin
        int_reg_array_7_34_real <= _zz_440_;
      end
      if(_zz_424_)begin
        int_reg_array_7_35_real <= _zz_440_;
      end
      if(_zz_425_)begin
        int_reg_array_7_36_real <= _zz_440_;
      end
      if(_zz_426_)begin
        int_reg_array_7_37_real <= _zz_440_;
      end
      if(_zz_427_)begin
        int_reg_array_7_38_real <= _zz_440_;
      end
      if(_zz_428_)begin
        int_reg_array_7_39_real <= _zz_440_;
      end
      if(_zz_429_)begin
        int_reg_array_7_40_real <= _zz_440_;
      end
      if(_zz_430_)begin
        int_reg_array_7_41_real <= _zz_440_;
      end
      if(_zz_431_)begin
        int_reg_array_7_42_real <= _zz_440_;
      end
      if(_zz_432_)begin
        int_reg_array_7_43_real <= _zz_440_;
      end
      if(_zz_433_)begin
        int_reg_array_7_44_real <= _zz_440_;
      end
      if(_zz_434_)begin
        int_reg_array_7_45_real <= _zz_440_;
      end
      if(_zz_435_)begin
        int_reg_array_7_46_real <= _zz_440_;
      end
      if(_zz_436_)begin
        int_reg_array_7_47_real <= _zz_440_;
      end
      if(_zz_437_)begin
        int_reg_array_7_48_real <= _zz_440_;
      end
      if(_zz_438_)begin
        int_reg_array_7_49_real <= _zz_440_;
      end
      if(_zz_389_)begin
        int_reg_array_7_0_imag <= _zz_441_;
      end
      if(_zz_390_)begin
        int_reg_array_7_1_imag <= _zz_441_;
      end
      if(_zz_391_)begin
        int_reg_array_7_2_imag <= _zz_441_;
      end
      if(_zz_392_)begin
        int_reg_array_7_3_imag <= _zz_441_;
      end
      if(_zz_393_)begin
        int_reg_array_7_4_imag <= _zz_441_;
      end
      if(_zz_394_)begin
        int_reg_array_7_5_imag <= _zz_441_;
      end
      if(_zz_395_)begin
        int_reg_array_7_6_imag <= _zz_441_;
      end
      if(_zz_396_)begin
        int_reg_array_7_7_imag <= _zz_441_;
      end
      if(_zz_397_)begin
        int_reg_array_7_8_imag <= _zz_441_;
      end
      if(_zz_398_)begin
        int_reg_array_7_9_imag <= _zz_441_;
      end
      if(_zz_399_)begin
        int_reg_array_7_10_imag <= _zz_441_;
      end
      if(_zz_400_)begin
        int_reg_array_7_11_imag <= _zz_441_;
      end
      if(_zz_401_)begin
        int_reg_array_7_12_imag <= _zz_441_;
      end
      if(_zz_402_)begin
        int_reg_array_7_13_imag <= _zz_441_;
      end
      if(_zz_403_)begin
        int_reg_array_7_14_imag <= _zz_441_;
      end
      if(_zz_404_)begin
        int_reg_array_7_15_imag <= _zz_441_;
      end
      if(_zz_405_)begin
        int_reg_array_7_16_imag <= _zz_441_;
      end
      if(_zz_406_)begin
        int_reg_array_7_17_imag <= _zz_441_;
      end
      if(_zz_407_)begin
        int_reg_array_7_18_imag <= _zz_441_;
      end
      if(_zz_408_)begin
        int_reg_array_7_19_imag <= _zz_441_;
      end
      if(_zz_409_)begin
        int_reg_array_7_20_imag <= _zz_441_;
      end
      if(_zz_410_)begin
        int_reg_array_7_21_imag <= _zz_441_;
      end
      if(_zz_411_)begin
        int_reg_array_7_22_imag <= _zz_441_;
      end
      if(_zz_412_)begin
        int_reg_array_7_23_imag <= _zz_441_;
      end
      if(_zz_413_)begin
        int_reg_array_7_24_imag <= _zz_441_;
      end
      if(_zz_414_)begin
        int_reg_array_7_25_imag <= _zz_441_;
      end
      if(_zz_415_)begin
        int_reg_array_7_26_imag <= _zz_441_;
      end
      if(_zz_416_)begin
        int_reg_array_7_27_imag <= _zz_441_;
      end
      if(_zz_417_)begin
        int_reg_array_7_28_imag <= _zz_441_;
      end
      if(_zz_418_)begin
        int_reg_array_7_29_imag <= _zz_441_;
      end
      if(_zz_419_)begin
        int_reg_array_7_30_imag <= _zz_441_;
      end
      if(_zz_420_)begin
        int_reg_array_7_31_imag <= _zz_441_;
      end
      if(_zz_421_)begin
        int_reg_array_7_32_imag <= _zz_441_;
      end
      if(_zz_422_)begin
        int_reg_array_7_33_imag <= _zz_441_;
      end
      if(_zz_423_)begin
        int_reg_array_7_34_imag <= _zz_441_;
      end
      if(_zz_424_)begin
        int_reg_array_7_35_imag <= _zz_441_;
      end
      if(_zz_425_)begin
        int_reg_array_7_36_imag <= _zz_441_;
      end
      if(_zz_426_)begin
        int_reg_array_7_37_imag <= _zz_441_;
      end
      if(_zz_427_)begin
        int_reg_array_7_38_imag <= _zz_441_;
      end
      if(_zz_428_)begin
        int_reg_array_7_39_imag <= _zz_441_;
      end
      if(_zz_429_)begin
        int_reg_array_7_40_imag <= _zz_441_;
      end
      if(_zz_430_)begin
        int_reg_array_7_41_imag <= _zz_441_;
      end
      if(_zz_431_)begin
        int_reg_array_7_42_imag <= _zz_441_;
      end
      if(_zz_432_)begin
        int_reg_array_7_43_imag <= _zz_441_;
      end
      if(_zz_433_)begin
        int_reg_array_7_44_imag <= _zz_441_;
      end
      if(_zz_434_)begin
        int_reg_array_7_45_imag <= _zz_441_;
      end
      if(_zz_435_)begin
        int_reg_array_7_46_imag <= _zz_441_;
      end
      if(_zz_436_)begin
        int_reg_array_7_47_imag <= _zz_441_;
      end
      if(_zz_437_)begin
        int_reg_array_7_48_imag <= _zz_441_;
      end
      if(_zz_438_)begin
        int_reg_array_7_49_imag <= _zz_441_;
      end
      if(_zz_444_)begin
        int_reg_array_8_0_real <= _zz_495_;
      end
      if(_zz_445_)begin
        int_reg_array_8_1_real <= _zz_495_;
      end
      if(_zz_446_)begin
        int_reg_array_8_2_real <= _zz_495_;
      end
      if(_zz_447_)begin
        int_reg_array_8_3_real <= _zz_495_;
      end
      if(_zz_448_)begin
        int_reg_array_8_4_real <= _zz_495_;
      end
      if(_zz_449_)begin
        int_reg_array_8_5_real <= _zz_495_;
      end
      if(_zz_450_)begin
        int_reg_array_8_6_real <= _zz_495_;
      end
      if(_zz_451_)begin
        int_reg_array_8_7_real <= _zz_495_;
      end
      if(_zz_452_)begin
        int_reg_array_8_8_real <= _zz_495_;
      end
      if(_zz_453_)begin
        int_reg_array_8_9_real <= _zz_495_;
      end
      if(_zz_454_)begin
        int_reg_array_8_10_real <= _zz_495_;
      end
      if(_zz_455_)begin
        int_reg_array_8_11_real <= _zz_495_;
      end
      if(_zz_456_)begin
        int_reg_array_8_12_real <= _zz_495_;
      end
      if(_zz_457_)begin
        int_reg_array_8_13_real <= _zz_495_;
      end
      if(_zz_458_)begin
        int_reg_array_8_14_real <= _zz_495_;
      end
      if(_zz_459_)begin
        int_reg_array_8_15_real <= _zz_495_;
      end
      if(_zz_460_)begin
        int_reg_array_8_16_real <= _zz_495_;
      end
      if(_zz_461_)begin
        int_reg_array_8_17_real <= _zz_495_;
      end
      if(_zz_462_)begin
        int_reg_array_8_18_real <= _zz_495_;
      end
      if(_zz_463_)begin
        int_reg_array_8_19_real <= _zz_495_;
      end
      if(_zz_464_)begin
        int_reg_array_8_20_real <= _zz_495_;
      end
      if(_zz_465_)begin
        int_reg_array_8_21_real <= _zz_495_;
      end
      if(_zz_466_)begin
        int_reg_array_8_22_real <= _zz_495_;
      end
      if(_zz_467_)begin
        int_reg_array_8_23_real <= _zz_495_;
      end
      if(_zz_468_)begin
        int_reg_array_8_24_real <= _zz_495_;
      end
      if(_zz_469_)begin
        int_reg_array_8_25_real <= _zz_495_;
      end
      if(_zz_470_)begin
        int_reg_array_8_26_real <= _zz_495_;
      end
      if(_zz_471_)begin
        int_reg_array_8_27_real <= _zz_495_;
      end
      if(_zz_472_)begin
        int_reg_array_8_28_real <= _zz_495_;
      end
      if(_zz_473_)begin
        int_reg_array_8_29_real <= _zz_495_;
      end
      if(_zz_474_)begin
        int_reg_array_8_30_real <= _zz_495_;
      end
      if(_zz_475_)begin
        int_reg_array_8_31_real <= _zz_495_;
      end
      if(_zz_476_)begin
        int_reg_array_8_32_real <= _zz_495_;
      end
      if(_zz_477_)begin
        int_reg_array_8_33_real <= _zz_495_;
      end
      if(_zz_478_)begin
        int_reg_array_8_34_real <= _zz_495_;
      end
      if(_zz_479_)begin
        int_reg_array_8_35_real <= _zz_495_;
      end
      if(_zz_480_)begin
        int_reg_array_8_36_real <= _zz_495_;
      end
      if(_zz_481_)begin
        int_reg_array_8_37_real <= _zz_495_;
      end
      if(_zz_482_)begin
        int_reg_array_8_38_real <= _zz_495_;
      end
      if(_zz_483_)begin
        int_reg_array_8_39_real <= _zz_495_;
      end
      if(_zz_484_)begin
        int_reg_array_8_40_real <= _zz_495_;
      end
      if(_zz_485_)begin
        int_reg_array_8_41_real <= _zz_495_;
      end
      if(_zz_486_)begin
        int_reg_array_8_42_real <= _zz_495_;
      end
      if(_zz_487_)begin
        int_reg_array_8_43_real <= _zz_495_;
      end
      if(_zz_488_)begin
        int_reg_array_8_44_real <= _zz_495_;
      end
      if(_zz_489_)begin
        int_reg_array_8_45_real <= _zz_495_;
      end
      if(_zz_490_)begin
        int_reg_array_8_46_real <= _zz_495_;
      end
      if(_zz_491_)begin
        int_reg_array_8_47_real <= _zz_495_;
      end
      if(_zz_492_)begin
        int_reg_array_8_48_real <= _zz_495_;
      end
      if(_zz_493_)begin
        int_reg_array_8_49_real <= _zz_495_;
      end
      if(_zz_444_)begin
        int_reg_array_8_0_imag <= _zz_496_;
      end
      if(_zz_445_)begin
        int_reg_array_8_1_imag <= _zz_496_;
      end
      if(_zz_446_)begin
        int_reg_array_8_2_imag <= _zz_496_;
      end
      if(_zz_447_)begin
        int_reg_array_8_3_imag <= _zz_496_;
      end
      if(_zz_448_)begin
        int_reg_array_8_4_imag <= _zz_496_;
      end
      if(_zz_449_)begin
        int_reg_array_8_5_imag <= _zz_496_;
      end
      if(_zz_450_)begin
        int_reg_array_8_6_imag <= _zz_496_;
      end
      if(_zz_451_)begin
        int_reg_array_8_7_imag <= _zz_496_;
      end
      if(_zz_452_)begin
        int_reg_array_8_8_imag <= _zz_496_;
      end
      if(_zz_453_)begin
        int_reg_array_8_9_imag <= _zz_496_;
      end
      if(_zz_454_)begin
        int_reg_array_8_10_imag <= _zz_496_;
      end
      if(_zz_455_)begin
        int_reg_array_8_11_imag <= _zz_496_;
      end
      if(_zz_456_)begin
        int_reg_array_8_12_imag <= _zz_496_;
      end
      if(_zz_457_)begin
        int_reg_array_8_13_imag <= _zz_496_;
      end
      if(_zz_458_)begin
        int_reg_array_8_14_imag <= _zz_496_;
      end
      if(_zz_459_)begin
        int_reg_array_8_15_imag <= _zz_496_;
      end
      if(_zz_460_)begin
        int_reg_array_8_16_imag <= _zz_496_;
      end
      if(_zz_461_)begin
        int_reg_array_8_17_imag <= _zz_496_;
      end
      if(_zz_462_)begin
        int_reg_array_8_18_imag <= _zz_496_;
      end
      if(_zz_463_)begin
        int_reg_array_8_19_imag <= _zz_496_;
      end
      if(_zz_464_)begin
        int_reg_array_8_20_imag <= _zz_496_;
      end
      if(_zz_465_)begin
        int_reg_array_8_21_imag <= _zz_496_;
      end
      if(_zz_466_)begin
        int_reg_array_8_22_imag <= _zz_496_;
      end
      if(_zz_467_)begin
        int_reg_array_8_23_imag <= _zz_496_;
      end
      if(_zz_468_)begin
        int_reg_array_8_24_imag <= _zz_496_;
      end
      if(_zz_469_)begin
        int_reg_array_8_25_imag <= _zz_496_;
      end
      if(_zz_470_)begin
        int_reg_array_8_26_imag <= _zz_496_;
      end
      if(_zz_471_)begin
        int_reg_array_8_27_imag <= _zz_496_;
      end
      if(_zz_472_)begin
        int_reg_array_8_28_imag <= _zz_496_;
      end
      if(_zz_473_)begin
        int_reg_array_8_29_imag <= _zz_496_;
      end
      if(_zz_474_)begin
        int_reg_array_8_30_imag <= _zz_496_;
      end
      if(_zz_475_)begin
        int_reg_array_8_31_imag <= _zz_496_;
      end
      if(_zz_476_)begin
        int_reg_array_8_32_imag <= _zz_496_;
      end
      if(_zz_477_)begin
        int_reg_array_8_33_imag <= _zz_496_;
      end
      if(_zz_478_)begin
        int_reg_array_8_34_imag <= _zz_496_;
      end
      if(_zz_479_)begin
        int_reg_array_8_35_imag <= _zz_496_;
      end
      if(_zz_480_)begin
        int_reg_array_8_36_imag <= _zz_496_;
      end
      if(_zz_481_)begin
        int_reg_array_8_37_imag <= _zz_496_;
      end
      if(_zz_482_)begin
        int_reg_array_8_38_imag <= _zz_496_;
      end
      if(_zz_483_)begin
        int_reg_array_8_39_imag <= _zz_496_;
      end
      if(_zz_484_)begin
        int_reg_array_8_40_imag <= _zz_496_;
      end
      if(_zz_485_)begin
        int_reg_array_8_41_imag <= _zz_496_;
      end
      if(_zz_486_)begin
        int_reg_array_8_42_imag <= _zz_496_;
      end
      if(_zz_487_)begin
        int_reg_array_8_43_imag <= _zz_496_;
      end
      if(_zz_488_)begin
        int_reg_array_8_44_imag <= _zz_496_;
      end
      if(_zz_489_)begin
        int_reg_array_8_45_imag <= _zz_496_;
      end
      if(_zz_490_)begin
        int_reg_array_8_46_imag <= _zz_496_;
      end
      if(_zz_491_)begin
        int_reg_array_8_47_imag <= _zz_496_;
      end
      if(_zz_492_)begin
        int_reg_array_8_48_imag <= _zz_496_;
      end
      if(_zz_493_)begin
        int_reg_array_8_49_imag <= _zz_496_;
      end
      if(_zz_499_)begin
        int_reg_array_9_0_real <= _zz_550_;
      end
      if(_zz_500_)begin
        int_reg_array_9_1_real <= _zz_550_;
      end
      if(_zz_501_)begin
        int_reg_array_9_2_real <= _zz_550_;
      end
      if(_zz_502_)begin
        int_reg_array_9_3_real <= _zz_550_;
      end
      if(_zz_503_)begin
        int_reg_array_9_4_real <= _zz_550_;
      end
      if(_zz_504_)begin
        int_reg_array_9_5_real <= _zz_550_;
      end
      if(_zz_505_)begin
        int_reg_array_9_6_real <= _zz_550_;
      end
      if(_zz_506_)begin
        int_reg_array_9_7_real <= _zz_550_;
      end
      if(_zz_507_)begin
        int_reg_array_9_8_real <= _zz_550_;
      end
      if(_zz_508_)begin
        int_reg_array_9_9_real <= _zz_550_;
      end
      if(_zz_509_)begin
        int_reg_array_9_10_real <= _zz_550_;
      end
      if(_zz_510_)begin
        int_reg_array_9_11_real <= _zz_550_;
      end
      if(_zz_511_)begin
        int_reg_array_9_12_real <= _zz_550_;
      end
      if(_zz_512_)begin
        int_reg_array_9_13_real <= _zz_550_;
      end
      if(_zz_513_)begin
        int_reg_array_9_14_real <= _zz_550_;
      end
      if(_zz_514_)begin
        int_reg_array_9_15_real <= _zz_550_;
      end
      if(_zz_515_)begin
        int_reg_array_9_16_real <= _zz_550_;
      end
      if(_zz_516_)begin
        int_reg_array_9_17_real <= _zz_550_;
      end
      if(_zz_517_)begin
        int_reg_array_9_18_real <= _zz_550_;
      end
      if(_zz_518_)begin
        int_reg_array_9_19_real <= _zz_550_;
      end
      if(_zz_519_)begin
        int_reg_array_9_20_real <= _zz_550_;
      end
      if(_zz_520_)begin
        int_reg_array_9_21_real <= _zz_550_;
      end
      if(_zz_521_)begin
        int_reg_array_9_22_real <= _zz_550_;
      end
      if(_zz_522_)begin
        int_reg_array_9_23_real <= _zz_550_;
      end
      if(_zz_523_)begin
        int_reg_array_9_24_real <= _zz_550_;
      end
      if(_zz_524_)begin
        int_reg_array_9_25_real <= _zz_550_;
      end
      if(_zz_525_)begin
        int_reg_array_9_26_real <= _zz_550_;
      end
      if(_zz_526_)begin
        int_reg_array_9_27_real <= _zz_550_;
      end
      if(_zz_527_)begin
        int_reg_array_9_28_real <= _zz_550_;
      end
      if(_zz_528_)begin
        int_reg_array_9_29_real <= _zz_550_;
      end
      if(_zz_529_)begin
        int_reg_array_9_30_real <= _zz_550_;
      end
      if(_zz_530_)begin
        int_reg_array_9_31_real <= _zz_550_;
      end
      if(_zz_531_)begin
        int_reg_array_9_32_real <= _zz_550_;
      end
      if(_zz_532_)begin
        int_reg_array_9_33_real <= _zz_550_;
      end
      if(_zz_533_)begin
        int_reg_array_9_34_real <= _zz_550_;
      end
      if(_zz_534_)begin
        int_reg_array_9_35_real <= _zz_550_;
      end
      if(_zz_535_)begin
        int_reg_array_9_36_real <= _zz_550_;
      end
      if(_zz_536_)begin
        int_reg_array_9_37_real <= _zz_550_;
      end
      if(_zz_537_)begin
        int_reg_array_9_38_real <= _zz_550_;
      end
      if(_zz_538_)begin
        int_reg_array_9_39_real <= _zz_550_;
      end
      if(_zz_539_)begin
        int_reg_array_9_40_real <= _zz_550_;
      end
      if(_zz_540_)begin
        int_reg_array_9_41_real <= _zz_550_;
      end
      if(_zz_541_)begin
        int_reg_array_9_42_real <= _zz_550_;
      end
      if(_zz_542_)begin
        int_reg_array_9_43_real <= _zz_550_;
      end
      if(_zz_543_)begin
        int_reg_array_9_44_real <= _zz_550_;
      end
      if(_zz_544_)begin
        int_reg_array_9_45_real <= _zz_550_;
      end
      if(_zz_545_)begin
        int_reg_array_9_46_real <= _zz_550_;
      end
      if(_zz_546_)begin
        int_reg_array_9_47_real <= _zz_550_;
      end
      if(_zz_547_)begin
        int_reg_array_9_48_real <= _zz_550_;
      end
      if(_zz_548_)begin
        int_reg_array_9_49_real <= _zz_550_;
      end
      if(_zz_499_)begin
        int_reg_array_9_0_imag <= _zz_551_;
      end
      if(_zz_500_)begin
        int_reg_array_9_1_imag <= _zz_551_;
      end
      if(_zz_501_)begin
        int_reg_array_9_2_imag <= _zz_551_;
      end
      if(_zz_502_)begin
        int_reg_array_9_3_imag <= _zz_551_;
      end
      if(_zz_503_)begin
        int_reg_array_9_4_imag <= _zz_551_;
      end
      if(_zz_504_)begin
        int_reg_array_9_5_imag <= _zz_551_;
      end
      if(_zz_505_)begin
        int_reg_array_9_6_imag <= _zz_551_;
      end
      if(_zz_506_)begin
        int_reg_array_9_7_imag <= _zz_551_;
      end
      if(_zz_507_)begin
        int_reg_array_9_8_imag <= _zz_551_;
      end
      if(_zz_508_)begin
        int_reg_array_9_9_imag <= _zz_551_;
      end
      if(_zz_509_)begin
        int_reg_array_9_10_imag <= _zz_551_;
      end
      if(_zz_510_)begin
        int_reg_array_9_11_imag <= _zz_551_;
      end
      if(_zz_511_)begin
        int_reg_array_9_12_imag <= _zz_551_;
      end
      if(_zz_512_)begin
        int_reg_array_9_13_imag <= _zz_551_;
      end
      if(_zz_513_)begin
        int_reg_array_9_14_imag <= _zz_551_;
      end
      if(_zz_514_)begin
        int_reg_array_9_15_imag <= _zz_551_;
      end
      if(_zz_515_)begin
        int_reg_array_9_16_imag <= _zz_551_;
      end
      if(_zz_516_)begin
        int_reg_array_9_17_imag <= _zz_551_;
      end
      if(_zz_517_)begin
        int_reg_array_9_18_imag <= _zz_551_;
      end
      if(_zz_518_)begin
        int_reg_array_9_19_imag <= _zz_551_;
      end
      if(_zz_519_)begin
        int_reg_array_9_20_imag <= _zz_551_;
      end
      if(_zz_520_)begin
        int_reg_array_9_21_imag <= _zz_551_;
      end
      if(_zz_521_)begin
        int_reg_array_9_22_imag <= _zz_551_;
      end
      if(_zz_522_)begin
        int_reg_array_9_23_imag <= _zz_551_;
      end
      if(_zz_523_)begin
        int_reg_array_9_24_imag <= _zz_551_;
      end
      if(_zz_524_)begin
        int_reg_array_9_25_imag <= _zz_551_;
      end
      if(_zz_525_)begin
        int_reg_array_9_26_imag <= _zz_551_;
      end
      if(_zz_526_)begin
        int_reg_array_9_27_imag <= _zz_551_;
      end
      if(_zz_527_)begin
        int_reg_array_9_28_imag <= _zz_551_;
      end
      if(_zz_528_)begin
        int_reg_array_9_29_imag <= _zz_551_;
      end
      if(_zz_529_)begin
        int_reg_array_9_30_imag <= _zz_551_;
      end
      if(_zz_530_)begin
        int_reg_array_9_31_imag <= _zz_551_;
      end
      if(_zz_531_)begin
        int_reg_array_9_32_imag <= _zz_551_;
      end
      if(_zz_532_)begin
        int_reg_array_9_33_imag <= _zz_551_;
      end
      if(_zz_533_)begin
        int_reg_array_9_34_imag <= _zz_551_;
      end
      if(_zz_534_)begin
        int_reg_array_9_35_imag <= _zz_551_;
      end
      if(_zz_535_)begin
        int_reg_array_9_36_imag <= _zz_551_;
      end
      if(_zz_536_)begin
        int_reg_array_9_37_imag <= _zz_551_;
      end
      if(_zz_537_)begin
        int_reg_array_9_38_imag <= _zz_551_;
      end
      if(_zz_538_)begin
        int_reg_array_9_39_imag <= _zz_551_;
      end
      if(_zz_539_)begin
        int_reg_array_9_40_imag <= _zz_551_;
      end
      if(_zz_540_)begin
        int_reg_array_9_41_imag <= _zz_551_;
      end
      if(_zz_541_)begin
        int_reg_array_9_42_imag <= _zz_551_;
      end
      if(_zz_542_)begin
        int_reg_array_9_43_imag <= _zz_551_;
      end
      if(_zz_543_)begin
        int_reg_array_9_44_imag <= _zz_551_;
      end
      if(_zz_544_)begin
        int_reg_array_9_45_imag <= _zz_551_;
      end
      if(_zz_545_)begin
        int_reg_array_9_46_imag <= _zz_551_;
      end
      if(_zz_546_)begin
        int_reg_array_9_47_imag <= _zz_551_;
      end
      if(_zz_547_)begin
        int_reg_array_9_48_imag <= _zz_551_;
      end
      if(_zz_548_)begin
        int_reg_array_9_49_imag <= _zz_551_;
      end
      if(_zz_554_)begin
        int_reg_array_10_0_real <= _zz_605_;
      end
      if(_zz_555_)begin
        int_reg_array_10_1_real <= _zz_605_;
      end
      if(_zz_556_)begin
        int_reg_array_10_2_real <= _zz_605_;
      end
      if(_zz_557_)begin
        int_reg_array_10_3_real <= _zz_605_;
      end
      if(_zz_558_)begin
        int_reg_array_10_4_real <= _zz_605_;
      end
      if(_zz_559_)begin
        int_reg_array_10_5_real <= _zz_605_;
      end
      if(_zz_560_)begin
        int_reg_array_10_6_real <= _zz_605_;
      end
      if(_zz_561_)begin
        int_reg_array_10_7_real <= _zz_605_;
      end
      if(_zz_562_)begin
        int_reg_array_10_8_real <= _zz_605_;
      end
      if(_zz_563_)begin
        int_reg_array_10_9_real <= _zz_605_;
      end
      if(_zz_564_)begin
        int_reg_array_10_10_real <= _zz_605_;
      end
      if(_zz_565_)begin
        int_reg_array_10_11_real <= _zz_605_;
      end
      if(_zz_566_)begin
        int_reg_array_10_12_real <= _zz_605_;
      end
      if(_zz_567_)begin
        int_reg_array_10_13_real <= _zz_605_;
      end
      if(_zz_568_)begin
        int_reg_array_10_14_real <= _zz_605_;
      end
      if(_zz_569_)begin
        int_reg_array_10_15_real <= _zz_605_;
      end
      if(_zz_570_)begin
        int_reg_array_10_16_real <= _zz_605_;
      end
      if(_zz_571_)begin
        int_reg_array_10_17_real <= _zz_605_;
      end
      if(_zz_572_)begin
        int_reg_array_10_18_real <= _zz_605_;
      end
      if(_zz_573_)begin
        int_reg_array_10_19_real <= _zz_605_;
      end
      if(_zz_574_)begin
        int_reg_array_10_20_real <= _zz_605_;
      end
      if(_zz_575_)begin
        int_reg_array_10_21_real <= _zz_605_;
      end
      if(_zz_576_)begin
        int_reg_array_10_22_real <= _zz_605_;
      end
      if(_zz_577_)begin
        int_reg_array_10_23_real <= _zz_605_;
      end
      if(_zz_578_)begin
        int_reg_array_10_24_real <= _zz_605_;
      end
      if(_zz_579_)begin
        int_reg_array_10_25_real <= _zz_605_;
      end
      if(_zz_580_)begin
        int_reg_array_10_26_real <= _zz_605_;
      end
      if(_zz_581_)begin
        int_reg_array_10_27_real <= _zz_605_;
      end
      if(_zz_582_)begin
        int_reg_array_10_28_real <= _zz_605_;
      end
      if(_zz_583_)begin
        int_reg_array_10_29_real <= _zz_605_;
      end
      if(_zz_584_)begin
        int_reg_array_10_30_real <= _zz_605_;
      end
      if(_zz_585_)begin
        int_reg_array_10_31_real <= _zz_605_;
      end
      if(_zz_586_)begin
        int_reg_array_10_32_real <= _zz_605_;
      end
      if(_zz_587_)begin
        int_reg_array_10_33_real <= _zz_605_;
      end
      if(_zz_588_)begin
        int_reg_array_10_34_real <= _zz_605_;
      end
      if(_zz_589_)begin
        int_reg_array_10_35_real <= _zz_605_;
      end
      if(_zz_590_)begin
        int_reg_array_10_36_real <= _zz_605_;
      end
      if(_zz_591_)begin
        int_reg_array_10_37_real <= _zz_605_;
      end
      if(_zz_592_)begin
        int_reg_array_10_38_real <= _zz_605_;
      end
      if(_zz_593_)begin
        int_reg_array_10_39_real <= _zz_605_;
      end
      if(_zz_594_)begin
        int_reg_array_10_40_real <= _zz_605_;
      end
      if(_zz_595_)begin
        int_reg_array_10_41_real <= _zz_605_;
      end
      if(_zz_596_)begin
        int_reg_array_10_42_real <= _zz_605_;
      end
      if(_zz_597_)begin
        int_reg_array_10_43_real <= _zz_605_;
      end
      if(_zz_598_)begin
        int_reg_array_10_44_real <= _zz_605_;
      end
      if(_zz_599_)begin
        int_reg_array_10_45_real <= _zz_605_;
      end
      if(_zz_600_)begin
        int_reg_array_10_46_real <= _zz_605_;
      end
      if(_zz_601_)begin
        int_reg_array_10_47_real <= _zz_605_;
      end
      if(_zz_602_)begin
        int_reg_array_10_48_real <= _zz_605_;
      end
      if(_zz_603_)begin
        int_reg_array_10_49_real <= _zz_605_;
      end
      if(_zz_554_)begin
        int_reg_array_10_0_imag <= _zz_606_;
      end
      if(_zz_555_)begin
        int_reg_array_10_1_imag <= _zz_606_;
      end
      if(_zz_556_)begin
        int_reg_array_10_2_imag <= _zz_606_;
      end
      if(_zz_557_)begin
        int_reg_array_10_3_imag <= _zz_606_;
      end
      if(_zz_558_)begin
        int_reg_array_10_4_imag <= _zz_606_;
      end
      if(_zz_559_)begin
        int_reg_array_10_5_imag <= _zz_606_;
      end
      if(_zz_560_)begin
        int_reg_array_10_6_imag <= _zz_606_;
      end
      if(_zz_561_)begin
        int_reg_array_10_7_imag <= _zz_606_;
      end
      if(_zz_562_)begin
        int_reg_array_10_8_imag <= _zz_606_;
      end
      if(_zz_563_)begin
        int_reg_array_10_9_imag <= _zz_606_;
      end
      if(_zz_564_)begin
        int_reg_array_10_10_imag <= _zz_606_;
      end
      if(_zz_565_)begin
        int_reg_array_10_11_imag <= _zz_606_;
      end
      if(_zz_566_)begin
        int_reg_array_10_12_imag <= _zz_606_;
      end
      if(_zz_567_)begin
        int_reg_array_10_13_imag <= _zz_606_;
      end
      if(_zz_568_)begin
        int_reg_array_10_14_imag <= _zz_606_;
      end
      if(_zz_569_)begin
        int_reg_array_10_15_imag <= _zz_606_;
      end
      if(_zz_570_)begin
        int_reg_array_10_16_imag <= _zz_606_;
      end
      if(_zz_571_)begin
        int_reg_array_10_17_imag <= _zz_606_;
      end
      if(_zz_572_)begin
        int_reg_array_10_18_imag <= _zz_606_;
      end
      if(_zz_573_)begin
        int_reg_array_10_19_imag <= _zz_606_;
      end
      if(_zz_574_)begin
        int_reg_array_10_20_imag <= _zz_606_;
      end
      if(_zz_575_)begin
        int_reg_array_10_21_imag <= _zz_606_;
      end
      if(_zz_576_)begin
        int_reg_array_10_22_imag <= _zz_606_;
      end
      if(_zz_577_)begin
        int_reg_array_10_23_imag <= _zz_606_;
      end
      if(_zz_578_)begin
        int_reg_array_10_24_imag <= _zz_606_;
      end
      if(_zz_579_)begin
        int_reg_array_10_25_imag <= _zz_606_;
      end
      if(_zz_580_)begin
        int_reg_array_10_26_imag <= _zz_606_;
      end
      if(_zz_581_)begin
        int_reg_array_10_27_imag <= _zz_606_;
      end
      if(_zz_582_)begin
        int_reg_array_10_28_imag <= _zz_606_;
      end
      if(_zz_583_)begin
        int_reg_array_10_29_imag <= _zz_606_;
      end
      if(_zz_584_)begin
        int_reg_array_10_30_imag <= _zz_606_;
      end
      if(_zz_585_)begin
        int_reg_array_10_31_imag <= _zz_606_;
      end
      if(_zz_586_)begin
        int_reg_array_10_32_imag <= _zz_606_;
      end
      if(_zz_587_)begin
        int_reg_array_10_33_imag <= _zz_606_;
      end
      if(_zz_588_)begin
        int_reg_array_10_34_imag <= _zz_606_;
      end
      if(_zz_589_)begin
        int_reg_array_10_35_imag <= _zz_606_;
      end
      if(_zz_590_)begin
        int_reg_array_10_36_imag <= _zz_606_;
      end
      if(_zz_591_)begin
        int_reg_array_10_37_imag <= _zz_606_;
      end
      if(_zz_592_)begin
        int_reg_array_10_38_imag <= _zz_606_;
      end
      if(_zz_593_)begin
        int_reg_array_10_39_imag <= _zz_606_;
      end
      if(_zz_594_)begin
        int_reg_array_10_40_imag <= _zz_606_;
      end
      if(_zz_595_)begin
        int_reg_array_10_41_imag <= _zz_606_;
      end
      if(_zz_596_)begin
        int_reg_array_10_42_imag <= _zz_606_;
      end
      if(_zz_597_)begin
        int_reg_array_10_43_imag <= _zz_606_;
      end
      if(_zz_598_)begin
        int_reg_array_10_44_imag <= _zz_606_;
      end
      if(_zz_599_)begin
        int_reg_array_10_45_imag <= _zz_606_;
      end
      if(_zz_600_)begin
        int_reg_array_10_46_imag <= _zz_606_;
      end
      if(_zz_601_)begin
        int_reg_array_10_47_imag <= _zz_606_;
      end
      if(_zz_602_)begin
        int_reg_array_10_48_imag <= _zz_606_;
      end
      if(_zz_603_)begin
        int_reg_array_10_49_imag <= _zz_606_;
      end
      if(_zz_609_)begin
        int_reg_array_11_0_real <= _zz_660_;
      end
      if(_zz_610_)begin
        int_reg_array_11_1_real <= _zz_660_;
      end
      if(_zz_611_)begin
        int_reg_array_11_2_real <= _zz_660_;
      end
      if(_zz_612_)begin
        int_reg_array_11_3_real <= _zz_660_;
      end
      if(_zz_613_)begin
        int_reg_array_11_4_real <= _zz_660_;
      end
      if(_zz_614_)begin
        int_reg_array_11_5_real <= _zz_660_;
      end
      if(_zz_615_)begin
        int_reg_array_11_6_real <= _zz_660_;
      end
      if(_zz_616_)begin
        int_reg_array_11_7_real <= _zz_660_;
      end
      if(_zz_617_)begin
        int_reg_array_11_8_real <= _zz_660_;
      end
      if(_zz_618_)begin
        int_reg_array_11_9_real <= _zz_660_;
      end
      if(_zz_619_)begin
        int_reg_array_11_10_real <= _zz_660_;
      end
      if(_zz_620_)begin
        int_reg_array_11_11_real <= _zz_660_;
      end
      if(_zz_621_)begin
        int_reg_array_11_12_real <= _zz_660_;
      end
      if(_zz_622_)begin
        int_reg_array_11_13_real <= _zz_660_;
      end
      if(_zz_623_)begin
        int_reg_array_11_14_real <= _zz_660_;
      end
      if(_zz_624_)begin
        int_reg_array_11_15_real <= _zz_660_;
      end
      if(_zz_625_)begin
        int_reg_array_11_16_real <= _zz_660_;
      end
      if(_zz_626_)begin
        int_reg_array_11_17_real <= _zz_660_;
      end
      if(_zz_627_)begin
        int_reg_array_11_18_real <= _zz_660_;
      end
      if(_zz_628_)begin
        int_reg_array_11_19_real <= _zz_660_;
      end
      if(_zz_629_)begin
        int_reg_array_11_20_real <= _zz_660_;
      end
      if(_zz_630_)begin
        int_reg_array_11_21_real <= _zz_660_;
      end
      if(_zz_631_)begin
        int_reg_array_11_22_real <= _zz_660_;
      end
      if(_zz_632_)begin
        int_reg_array_11_23_real <= _zz_660_;
      end
      if(_zz_633_)begin
        int_reg_array_11_24_real <= _zz_660_;
      end
      if(_zz_634_)begin
        int_reg_array_11_25_real <= _zz_660_;
      end
      if(_zz_635_)begin
        int_reg_array_11_26_real <= _zz_660_;
      end
      if(_zz_636_)begin
        int_reg_array_11_27_real <= _zz_660_;
      end
      if(_zz_637_)begin
        int_reg_array_11_28_real <= _zz_660_;
      end
      if(_zz_638_)begin
        int_reg_array_11_29_real <= _zz_660_;
      end
      if(_zz_639_)begin
        int_reg_array_11_30_real <= _zz_660_;
      end
      if(_zz_640_)begin
        int_reg_array_11_31_real <= _zz_660_;
      end
      if(_zz_641_)begin
        int_reg_array_11_32_real <= _zz_660_;
      end
      if(_zz_642_)begin
        int_reg_array_11_33_real <= _zz_660_;
      end
      if(_zz_643_)begin
        int_reg_array_11_34_real <= _zz_660_;
      end
      if(_zz_644_)begin
        int_reg_array_11_35_real <= _zz_660_;
      end
      if(_zz_645_)begin
        int_reg_array_11_36_real <= _zz_660_;
      end
      if(_zz_646_)begin
        int_reg_array_11_37_real <= _zz_660_;
      end
      if(_zz_647_)begin
        int_reg_array_11_38_real <= _zz_660_;
      end
      if(_zz_648_)begin
        int_reg_array_11_39_real <= _zz_660_;
      end
      if(_zz_649_)begin
        int_reg_array_11_40_real <= _zz_660_;
      end
      if(_zz_650_)begin
        int_reg_array_11_41_real <= _zz_660_;
      end
      if(_zz_651_)begin
        int_reg_array_11_42_real <= _zz_660_;
      end
      if(_zz_652_)begin
        int_reg_array_11_43_real <= _zz_660_;
      end
      if(_zz_653_)begin
        int_reg_array_11_44_real <= _zz_660_;
      end
      if(_zz_654_)begin
        int_reg_array_11_45_real <= _zz_660_;
      end
      if(_zz_655_)begin
        int_reg_array_11_46_real <= _zz_660_;
      end
      if(_zz_656_)begin
        int_reg_array_11_47_real <= _zz_660_;
      end
      if(_zz_657_)begin
        int_reg_array_11_48_real <= _zz_660_;
      end
      if(_zz_658_)begin
        int_reg_array_11_49_real <= _zz_660_;
      end
      if(_zz_609_)begin
        int_reg_array_11_0_imag <= _zz_661_;
      end
      if(_zz_610_)begin
        int_reg_array_11_1_imag <= _zz_661_;
      end
      if(_zz_611_)begin
        int_reg_array_11_2_imag <= _zz_661_;
      end
      if(_zz_612_)begin
        int_reg_array_11_3_imag <= _zz_661_;
      end
      if(_zz_613_)begin
        int_reg_array_11_4_imag <= _zz_661_;
      end
      if(_zz_614_)begin
        int_reg_array_11_5_imag <= _zz_661_;
      end
      if(_zz_615_)begin
        int_reg_array_11_6_imag <= _zz_661_;
      end
      if(_zz_616_)begin
        int_reg_array_11_7_imag <= _zz_661_;
      end
      if(_zz_617_)begin
        int_reg_array_11_8_imag <= _zz_661_;
      end
      if(_zz_618_)begin
        int_reg_array_11_9_imag <= _zz_661_;
      end
      if(_zz_619_)begin
        int_reg_array_11_10_imag <= _zz_661_;
      end
      if(_zz_620_)begin
        int_reg_array_11_11_imag <= _zz_661_;
      end
      if(_zz_621_)begin
        int_reg_array_11_12_imag <= _zz_661_;
      end
      if(_zz_622_)begin
        int_reg_array_11_13_imag <= _zz_661_;
      end
      if(_zz_623_)begin
        int_reg_array_11_14_imag <= _zz_661_;
      end
      if(_zz_624_)begin
        int_reg_array_11_15_imag <= _zz_661_;
      end
      if(_zz_625_)begin
        int_reg_array_11_16_imag <= _zz_661_;
      end
      if(_zz_626_)begin
        int_reg_array_11_17_imag <= _zz_661_;
      end
      if(_zz_627_)begin
        int_reg_array_11_18_imag <= _zz_661_;
      end
      if(_zz_628_)begin
        int_reg_array_11_19_imag <= _zz_661_;
      end
      if(_zz_629_)begin
        int_reg_array_11_20_imag <= _zz_661_;
      end
      if(_zz_630_)begin
        int_reg_array_11_21_imag <= _zz_661_;
      end
      if(_zz_631_)begin
        int_reg_array_11_22_imag <= _zz_661_;
      end
      if(_zz_632_)begin
        int_reg_array_11_23_imag <= _zz_661_;
      end
      if(_zz_633_)begin
        int_reg_array_11_24_imag <= _zz_661_;
      end
      if(_zz_634_)begin
        int_reg_array_11_25_imag <= _zz_661_;
      end
      if(_zz_635_)begin
        int_reg_array_11_26_imag <= _zz_661_;
      end
      if(_zz_636_)begin
        int_reg_array_11_27_imag <= _zz_661_;
      end
      if(_zz_637_)begin
        int_reg_array_11_28_imag <= _zz_661_;
      end
      if(_zz_638_)begin
        int_reg_array_11_29_imag <= _zz_661_;
      end
      if(_zz_639_)begin
        int_reg_array_11_30_imag <= _zz_661_;
      end
      if(_zz_640_)begin
        int_reg_array_11_31_imag <= _zz_661_;
      end
      if(_zz_641_)begin
        int_reg_array_11_32_imag <= _zz_661_;
      end
      if(_zz_642_)begin
        int_reg_array_11_33_imag <= _zz_661_;
      end
      if(_zz_643_)begin
        int_reg_array_11_34_imag <= _zz_661_;
      end
      if(_zz_644_)begin
        int_reg_array_11_35_imag <= _zz_661_;
      end
      if(_zz_645_)begin
        int_reg_array_11_36_imag <= _zz_661_;
      end
      if(_zz_646_)begin
        int_reg_array_11_37_imag <= _zz_661_;
      end
      if(_zz_647_)begin
        int_reg_array_11_38_imag <= _zz_661_;
      end
      if(_zz_648_)begin
        int_reg_array_11_39_imag <= _zz_661_;
      end
      if(_zz_649_)begin
        int_reg_array_11_40_imag <= _zz_661_;
      end
      if(_zz_650_)begin
        int_reg_array_11_41_imag <= _zz_661_;
      end
      if(_zz_651_)begin
        int_reg_array_11_42_imag <= _zz_661_;
      end
      if(_zz_652_)begin
        int_reg_array_11_43_imag <= _zz_661_;
      end
      if(_zz_653_)begin
        int_reg_array_11_44_imag <= _zz_661_;
      end
      if(_zz_654_)begin
        int_reg_array_11_45_imag <= _zz_661_;
      end
      if(_zz_655_)begin
        int_reg_array_11_46_imag <= _zz_661_;
      end
      if(_zz_656_)begin
        int_reg_array_11_47_imag <= _zz_661_;
      end
      if(_zz_657_)begin
        int_reg_array_11_48_imag <= _zz_661_;
      end
      if(_zz_658_)begin
        int_reg_array_11_49_imag <= _zz_661_;
      end
      if(_zz_664_)begin
        int_reg_array_12_0_real <= _zz_715_;
      end
      if(_zz_665_)begin
        int_reg_array_12_1_real <= _zz_715_;
      end
      if(_zz_666_)begin
        int_reg_array_12_2_real <= _zz_715_;
      end
      if(_zz_667_)begin
        int_reg_array_12_3_real <= _zz_715_;
      end
      if(_zz_668_)begin
        int_reg_array_12_4_real <= _zz_715_;
      end
      if(_zz_669_)begin
        int_reg_array_12_5_real <= _zz_715_;
      end
      if(_zz_670_)begin
        int_reg_array_12_6_real <= _zz_715_;
      end
      if(_zz_671_)begin
        int_reg_array_12_7_real <= _zz_715_;
      end
      if(_zz_672_)begin
        int_reg_array_12_8_real <= _zz_715_;
      end
      if(_zz_673_)begin
        int_reg_array_12_9_real <= _zz_715_;
      end
      if(_zz_674_)begin
        int_reg_array_12_10_real <= _zz_715_;
      end
      if(_zz_675_)begin
        int_reg_array_12_11_real <= _zz_715_;
      end
      if(_zz_676_)begin
        int_reg_array_12_12_real <= _zz_715_;
      end
      if(_zz_677_)begin
        int_reg_array_12_13_real <= _zz_715_;
      end
      if(_zz_678_)begin
        int_reg_array_12_14_real <= _zz_715_;
      end
      if(_zz_679_)begin
        int_reg_array_12_15_real <= _zz_715_;
      end
      if(_zz_680_)begin
        int_reg_array_12_16_real <= _zz_715_;
      end
      if(_zz_681_)begin
        int_reg_array_12_17_real <= _zz_715_;
      end
      if(_zz_682_)begin
        int_reg_array_12_18_real <= _zz_715_;
      end
      if(_zz_683_)begin
        int_reg_array_12_19_real <= _zz_715_;
      end
      if(_zz_684_)begin
        int_reg_array_12_20_real <= _zz_715_;
      end
      if(_zz_685_)begin
        int_reg_array_12_21_real <= _zz_715_;
      end
      if(_zz_686_)begin
        int_reg_array_12_22_real <= _zz_715_;
      end
      if(_zz_687_)begin
        int_reg_array_12_23_real <= _zz_715_;
      end
      if(_zz_688_)begin
        int_reg_array_12_24_real <= _zz_715_;
      end
      if(_zz_689_)begin
        int_reg_array_12_25_real <= _zz_715_;
      end
      if(_zz_690_)begin
        int_reg_array_12_26_real <= _zz_715_;
      end
      if(_zz_691_)begin
        int_reg_array_12_27_real <= _zz_715_;
      end
      if(_zz_692_)begin
        int_reg_array_12_28_real <= _zz_715_;
      end
      if(_zz_693_)begin
        int_reg_array_12_29_real <= _zz_715_;
      end
      if(_zz_694_)begin
        int_reg_array_12_30_real <= _zz_715_;
      end
      if(_zz_695_)begin
        int_reg_array_12_31_real <= _zz_715_;
      end
      if(_zz_696_)begin
        int_reg_array_12_32_real <= _zz_715_;
      end
      if(_zz_697_)begin
        int_reg_array_12_33_real <= _zz_715_;
      end
      if(_zz_698_)begin
        int_reg_array_12_34_real <= _zz_715_;
      end
      if(_zz_699_)begin
        int_reg_array_12_35_real <= _zz_715_;
      end
      if(_zz_700_)begin
        int_reg_array_12_36_real <= _zz_715_;
      end
      if(_zz_701_)begin
        int_reg_array_12_37_real <= _zz_715_;
      end
      if(_zz_702_)begin
        int_reg_array_12_38_real <= _zz_715_;
      end
      if(_zz_703_)begin
        int_reg_array_12_39_real <= _zz_715_;
      end
      if(_zz_704_)begin
        int_reg_array_12_40_real <= _zz_715_;
      end
      if(_zz_705_)begin
        int_reg_array_12_41_real <= _zz_715_;
      end
      if(_zz_706_)begin
        int_reg_array_12_42_real <= _zz_715_;
      end
      if(_zz_707_)begin
        int_reg_array_12_43_real <= _zz_715_;
      end
      if(_zz_708_)begin
        int_reg_array_12_44_real <= _zz_715_;
      end
      if(_zz_709_)begin
        int_reg_array_12_45_real <= _zz_715_;
      end
      if(_zz_710_)begin
        int_reg_array_12_46_real <= _zz_715_;
      end
      if(_zz_711_)begin
        int_reg_array_12_47_real <= _zz_715_;
      end
      if(_zz_712_)begin
        int_reg_array_12_48_real <= _zz_715_;
      end
      if(_zz_713_)begin
        int_reg_array_12_49_real <= _zz_715_;
      end
      if(_zz_664_)begin
        int_reg_array_12_0_imag <= _zz_716_;
      end
      if(_zz_665_)begin
        int_reg_array_12_1_imag <= _zz_716_;
      end
      if(_zz_666_)begin
        int_reg_array_12_2_imag <= _zz_716_;
      end
      if(_zz_667_)begin
        int_reg_array_12_3_imag <= _zz_716_;
      end
      if(_zz_668_)begin
        int_reg_array_12_4_imag <= _zz_716_;
      end
      if(_zz_669_)begin
        int_reg_array_12_5_imag <= _zz_716_;
      end
      if(_zz_670_)begin
        int_reg_array_12_6_imag <= _zz_716_;
      end
      if(_zz_671_)begin
        int_reg_array_12_7_imag <= _zz_716_;
      end
      if(_zz_672_)begin
        int_reg_array_12_8_imag <= _zz_716_;
      end
      if(_zz_673_)begin
        int_reg_array_12_9_imag <= _zz_716_;
      end
      if(_zz_674_)begin
        int_reg_array_12_10_imag <= _zz_716_;
      end
      if(_zz_675_)begin
        int_reg_array_12_11_imag <= _zz_716_;
      end
      if(_zz_676_)begin
        int_reg_array_12_12_imag <= _zz_716_;
      end
      if(_zz_677_)begin
        int_reg_array_12_13_imag <= _zz_716_;
      end
      if(_zz_678_)begin
        int_reg_array_12_14_imag <= _zz_716_;
      end
      if(_zz_679_)begin
        int_reg_array_12_15_imag <= _zz_716_;
      end
      if(_zz_680_)begin
        int_reg_array_12_16_imag <= _zz_716_;
      end
      if(_zz_681_)begin
        int_reg_array_12_17_imag <= _zz_716_;
      end
      if(_zz_682_)begin
        int_reg_array_12_18_imag <= _zz_716_;
      end
      if(_zz_683_)begin
        int_reg_array_12_19_imag <= _zz_716_;
      end
      if(_zz_684_)begin
        int_reg_array_12_20_imag <= _zz_716_;
      end
      if(_zz_685_)begin
        int_reg_array_12_21_imag <= _zz_716_;
      end
      if(_zz_686_)begin
        int_reg_array_12_22_imag <= _zz_716_;
      end
      if(_zz_687_)begin
        int_reg_array_12_23_imag <= _zz_716_;
      end
      if(_zz_688_)begin
        int_reg_array_12_24_imag <= _zz_716_;
      end
      if(_zz_689_)begin
        int_reg_array_12_25_imag <= _zz_716_;
      end
      if(_zz_690_)begin
        int_reg_array_12_26_imag <= _zz_716_;
      end
      if(_zz_691_)begin
        int_reg_array_12_27_imag <= _zz_716_;
      end
      if(_zz_692_)begin
        int_reg_array_12_28_imag <= _zz_716_;
      end
      if(_zz_693_)begin
        int_reg_array_12_29_imag <= _zz_716_;
      end
      if(_zz_694_)begin
        int_reg_array_12_30_imag <= _zz_716_;
      end
      if(_zz_695_)begin
        int_reg_array_12_31_imag <= _zz_716_;
      end
      if(_zz_696_)begin
        int_reg_array_12_32_imag <= _zz_716_;
      end
      if(_zz_697_)begin
        int_reg_array_12_33_imag <= _zz_716_;
      end
      if(_zz_698_)begin
        int_reg_array_12_34_imag <= _zz_716_;
      end
      if(_zz_699_)begin
        int_reg_array_12_35_imag <= _zz_716_;
      end
      if(_zz_700_)begin
        int_reg_array_12_36_imag <= _zz_716_;
      end
      if(_zz_701_)begin
        int_reg_array_12_37_imag <= _zz_716_;
      end
      if(_zz_702_)begin
        int_reg_array_12_38_imag <= _zz_716_;
      end
      if(_zz_703_)begin
        int_reg_array_12_39_imag <= _zz_716_;
      end
      if(_zz_704_)begin
        int_reg_array_12_40_imag <= _zz_716_;
      end
      if(_zz_705_)begin
        int_reg_array_12_41_imag <= _zz_716_;
      end
      if(_zz_706_)begin
        int_reg_array_12_42_imag <= _zz_716_;
      end
      if(_zz_707_)begin
        int_reg_array_12_43_imag <= _zz_716_;
      end
      if(_zz_708_)begin
        int_reg_array_12_44_imag <= _zz_716_;
      end
      if(_zz_709_)begin
        int_reg_array_12_45_imag <= _zz_716_;
      end
      if(_zz_710_)begin
        int_reg_array_12_46_imag <= _zz_716_;
      end
      if(_zz_711_)begin
        int_reg_array_12_47_imag <= _zz_716_;
      end
      if(_zz_712_)begin
        int_reg_array_12_48_imag <= _zz_716_;
      end
      if(_zz_713_)begin
        int_reg_array_12_49_imag <= _zz_716_;
      end
      if(_zz_719_)begin
        int_reg_array_13_0_real <= _zz_770_;
      end
      if(_zz_720_)begin
        int_reg_array_13_1_real <= _zz_770_;
      end
      if(_zz_721_)begin
        int_reg_array_13_2_real <= _zz_770_;
      end
      if(_zz_722_)begin
        int_reg_array_13_3_real <= _zz_770_;
      end
      if(_zz_723_)begin
        int_reg_array_13_4_real <= _zz_770_;
      end
      if(_zz_724_)begin
        int_reg_array_13_5_real <= _zz_770_;
      end
      if(_zz_725_)begin
        int_reg_array_13_6_real <= _zz_770_;
      end
      if(_zz_726_)begin
        int_reg_array_13_7_real <= _zz_770_;
      end
      if(_zz_727_)begin
        int_reg_array_13_8_real <= _zz_770_;
      end
      if(_zz_728_)begin
        int_reg_array_13_9_real <= _zz_770_;
      end
      if(_zz_729_)begin
        int_reg_array_13_10_real <= _zz_770_;
      end
      if(_zz_730_)begin
        int_reg_array_13_11_real <= _zz_770_;
      end
      if(_zz_731_)begin
        int_reg_array_13_12_real <= _zz_770_;
      end
      if(_zz_732_)begin
        int_reg_array_13_13_real <= _zz_770_;
      end
      if(_zz_733_)begin
        int_reg_array_13_14_real <= _zz_770_;
      end
      if(_zz_734_)begin
        int_reg_array_13_15_real <= _zz_770_;
      end
      if(_zz_735_)begin
        int_reg_array_13_16_real <= _zz_770_;
      end
      if(_zz_736_)begin
        int_reg_array_13_17_real <= _zz_770_;
      end
      if(_zz_737_)begin
        int_reg_array_13_18_real <= _zz_770_;
      end
      if(_zz_738_)begin
        int_reg_array_13_19_real <= _zz_770_;
      end
      if(_zz_739_)begin
        int_reg_array_13_20_real <= _zz_770_;
      end
      if(_zz_740_)begin
        int_reg_array_13_21_real <= _zz_770_;
      end
      if(_zz_741_)begin
        int_reg_array_13_22_real <= _zz_770_;
      end
      if(_zz_742_)begin
        int_reg_array_13_23_real <= _zz_770_;
      end
      if(_zz_743_)begin
        int_reg_array_13_24_real <= _zz_770_;
      end
      if(_zz_744_)begin
        int_reg_array_13_25_real <= _zz_770_;
      end
      if(_zz_745_)begin
        int_reg_array_13_26_real <= _zz_770_;
      end
      if(_zz_746_)begin
        int_reg_array_13_27_real <= _zz_770_;
      end
      if(_zz_747_)begin
        int_reg_array_13_28_real <= _zz_770_;
      end
      if(_zz_748_)begin
        int_reg_array_13_29_real <= _zz_770_;
      end
      if(_zz_749_)begin
        int_reg_array_13_30_real <= _zz_770_;
      end
      if(_zz_750_)begin
        int_reg_array_13_31_real <= _zz_770_;
      end
      if(_zz_751_)begin
        int_reg_array_13_32_real <= _zz_770_;
      end
      if(_zz_752_)begin
        int_reg_array_13_33_real <= _zz_770_;
      end
      if(_zz_753_)begin
        int_reg_array_13_34_real <= _zz_770_;
      end
      if(_zz_754_)begin
        int_reg_array_13_35_real <= _zz_770_;
      end
      if(_zz_755_)begin
        int_reg_array_13_36_real <= _zz_770_;
      end
      if(_zz_756_)begin
        int_reg_array_13_37_real <= _zz_770_;
      end
      if(_zz_757_)begin
        int_reg_array_13_38_real <= _zz_770_;
      end
      if(_zz_758_)begin
        int_reg_array_13_39_real <= _zz_770_;
      end
      if(_zz_759_)begin
        int_reg_array_13_40_real <= _zz_770_;
      end
      if(_zz_760_)begin
        int_reg_array_13_41_real <= _zz_770_;
      end
      if(_zz_761_)begin
        int_reg_array_13_42_real <= _zz_770_;
      end
      if(_zz_762_)begin
        int_reg_array_13_43_real <= _zz_770_;
      end
      if(_zz_763_)begin
        int_reg_array_13_44_real <= _zz_770_;
      end
      if(_zz_764_)begin
        int_reg_array_13_45_real <= _zz_770_;
      end
      if(_zz_765_)begin
        int_reg_array_13_46_real <= _zz_770_;
      end
      if(_zz_766_)begin
        int_reg_array_13_47_real <= _zz_770_;
      end
      if(_zz_767_)begin
        int_reg_array_13_48_real <= _zz_770_;
      end
      if(_zz_768_)begin
        int_reg_array_13_49_real <= _zz_770_;
      end
      if(_zz_719_)begin
        int_reg_array_13_0_imag <= _zz_771_;
      end
      if(_zz_720_)begin
        int_reg_array_13_1_imag <= _zz_771_;
      end
      if(_zz_721_)begin
        int_reg_array_13_2_imag <= _zz_771_;
      end
      if(_zz_722_)begin
        int_reg_array_13_3_imag <= _zz_771_;
      end
      if(_zz_723_)begin
        int_reg_array_13_4_imag <= _zz_771_;
      end
      if(_zz_724_)begin
        int_reg_array_13_5_imag <= _zz_771_;
      end
      if(_zz_725_)begin
        int_reg_array_13_6_imag <= _zz_771_;
      end
      if(_zz_726_)begin
        int_reg_array_13_7_imag <= _zz_771_;
      end
      if(_zz_727_)begin
        int_reg_array_13_8_imag <= _zz_771_;
      end
      if(_zz_728_)begin
        int_reg_array_13_9_imag <= _zz_771_;
      end
      if(_zz_729_)begin
        int_reg_array_13_10_imag <= _zz_771_;
      end
      if(_zz_730_)begin
        int_reg_array_13_11_imag <= _zz_771_;
      end
      if(_zz_731_)begin
        int_reg_array_13_12_imag <= _zz_771_;
      end
      if(_zz_732_)begin
        int_reg_array_13_13_imag <= _zz_771_;
      end
      if(_zz_733_)begin
        int_reg_array_13_14_imag <= _zz_771_;
      end
      if(_zz_734_)begin
        int_reg_array_13_15_imag <= _zz_771_;
      end
      if(_zz_735_)begin
        int_reg_array_13_16_imag <= _zz_771_;
      end
      if(_zz_736_)begin
        int_reg_array_13_17_imag <= _zz_771_;
      end
      if(_zz_737_)begin
        int_reg_array_13_18_imag <= _zz_771_;
      end
      if(_zz_738_)begin
        int_reg_array_13_19_imag <= _zz_771_;
      end
      if(_zz_739_)begin
        int_reg_array_13_20_imag <= _zz_771_;
      end
      if(_zz_740_)begin
        int_reg_array_13_21_imag <= _zz_771_;
      end
      if(_zz_741_)begin
        int_reg_array_13_22_imag <= _zz_771_;
      end
      if(_zz_742_)begin
        int_reg_array_13_23_imag <= _zz_771_;
      end
      if(_zz_743_)begin
        int_reg_array_13_24_imag <= _zz_771_;
      end
      if(_zz_744_)begin
        int_reg_array_13_25_imag <= _zz_771_;
      end
      if(_zz_745_)begin
        int_reg_array_13_26_imag <= _zz_771_;
      end
      if(_zz_746_)begin
        int_reg_array_13_27_imag <= _zz_771_;
      end
      if(_zz_747_)begin
        int_reg_array_13_28_imag <= _zz_771_;
      end
      if(_zz_748_)begin
        int_reg_array_13_29_imag <= _zz_771_;
      end
      if(_zz_749_)begin
        int_reg_array_13_30_imag <= _zz_771_;
      end
      if(_zz_750_)begin
        int_reg_array_13_31_imag <= _zz_771_;
      end
      if(_zz_751_)begin
        int_reg_array_13_32_imag <= _zz_771_;
      end
      if(_zz_752_)begin
        int_reg_array_13_33_imag <= _zz_771_;
      end
      if(_zz_753_)begin
        int_reg_array_13_34_imag <= _zz_771_;
      end
      if(_zz_754_)begin
        int_reg_array_13_35_imag <= _zz_771_;
      end
      if(_zz_755_)begin
        int_reg_array_13_36_imag <= _zz_771_;
      end
      if(_zz_756_)begin
        int_reg_array_13_37_imag <= _zz_771_;
      end
      if(_zz_757_)begin
        int_reg_array_13_38_imag <= _zz_771_;
      end
      if(_zz_758_)begin
        int_reg_array_13_39_imag <= _zz_771_;
      end
      if(_zz_759_)begin
        int_reg_array_13_40_imag <= _zz_771_;
      end
      if(_zz_760_)begin
        int_reg_array_13_41_imag <= _zz_771_;
      end
      if(_zz_761_)begin
        int_reg_array_13_42_imag <= _zz_771_;
      end
      if(_zz_762_)begin
        int_reg_array_13_43_imag <= _zz_771_;
      end
      if(_zz_763_)begin
        int_reg_array_13_44_imag <= _zz_771_;
      end
      if(_zz_764_)begin
        int_reg_array_13_45_imag <= _zz_771_;
      end
      if(_zz_765_)begin
        int_reg_array_13_46_imag <= _zz_771_;
      end
      if(_zz_766_)begin
        int_reg_array_13_47_imag <= _zz_771_;
      end
      if(_zz_767_)begin
        int_reg_array_13_48_imag <= _zz_771_;
      end
      if(_zz_768_)begin
        int_reg_array_13_49_imag <= _zz_771_;
      end
      if(_zz_774_)begin
        int_reg_array_14_0_real <= _zz_825_;
      end
      if(_zz_775_)begin
        int_reg_array_14_1_real <= _zz_825_;
      end
      if(_zz_776_)begin
        int_reg_array_14_2_real <= _zz_825_;
      end
      if(_zz_777_)begin
        int_reg_array_14_3_real <= _zz_825_;
      end
      if(_zz_778_)begin
        int_reg_array_14_4_real <= _zz_825_;
      end
      if(_zz_779_)begin
        int_reg_array_14_5_real <= _zz_825_;
      end
      if(_zz_780_)begin
        int_reg_array_14_6_real <= _zz_825_;
      end
      if(_zz_781_)begin
        int_reg_array_14_7_real <= _zz_825_;
      end
      if(_zz_782_)begin
        int_reg_array_14_8_real <= _zz_825_;
      end
      if(_zz_783_)begin
        int_reg_array_14_9_real <= _zz_825_;
      end
      if(_zz_784_)begin
        int_reg_array_14_10_real <= _zz_825_;
      end
      if(_zz_785_)begin
        int_reg_array_14_11_real <= _zz_825_;
      end
      if(_zz_786_)begin
        int_reg_array_14_12_real <= _zz_825_;
      end
      if(_zz_787_)begin
        int_reg_array_14_13_real <= _zz_825_;
      end
      if(_zz_788_)begin
        int_reg_array_14_14_real <= _zz_825_;
      end
      if(_zz_789_)begin
        int_reg_array_14_15_real <= _zz_825_;
      end
      if(_zz_790_)begin
        int_reg_array_14_16_real <= _zz_825_;
      end
      if(_zz_791_)begin
        int_reg_array_14_17_real <= _zz_825_;
      end
      if(_zz_792_)begin
        int_reg_array_14_18_real <= _zz_825_;
      end
      if(_zz_793_)begin
        int_reg_array_14_19_real <= _zz_825_;
      end
      if(_zz_794_)begin
        int_reg_array_14_20_real <= _zz_825_;
      end
      if(_zz_795_)begin
        int_reg_array_14_21_real <= _zz_825_;
      end
      if(_zz_796_)begin
        int_reg_array_14_22_real <= _zz_825_;
      end
      if(_zz_797_)begin
        int_reg_array_14_23_real <= _zz_825_;
      end
      if(_zz_798_)begin
        int_reg_array_14_24_real <= _zz_825_;
      end
      if(_zz_799_)begin
        int_reg_array_14_25_real <= _zz_825_;
      end
      if(_zz_800_)begin
        int_reg_array_14_26_real <= _zz_825_;
      end
      if(_zz_801_)begin
        int_reg_array_14_27_real <= _zz_825_;
      end
      if(_zz_802_)begin
        int_reg_array_14_28_real <= _zz_825_;
      end
      if(_zz_803_)begin
        int_reg_array_14_29_real <= _zz_825_;
      end
      if(_zz_804_)begin
        int_reg_array_14_30_real <= _zz_825_;
      end
      if(_zz_805_)begin
        int_reg_array_14_31_real <= _zz_825_;
      end
      if(_zz_806_)begin
        int_reg_array_14_32_real <= _zz_825_;
      end
      if(_zz_807_)begin
        int_reg_array_14_33_real <= _zz_825_;
      end
      if(_zz_808_)begin
        int_reg_array_14_34_real <= _zz_825_;
      end
      if(_zz_809_)begin
        int_reg_array_14_35_real <= _zz_825_;
      end
      if(_zz_810_)begin
        int_reg_array_14_36_real <= _zz_825_;
      end
      if(_zz_811_)begin
        int_reg_array_14_37_real <= _zz_825_;
      end
      if(_zz_812_)begin
        int_reg_array_14_38_real <= _zz_825_;
      end
      if(_zz_813_)begin
        int_reg_array_14_39_real <= _zz_825_;
      end
      if(_zz_814_)begin
        int_reg_array_14_40_real <= _zz_825_;
      end
      if(_zz_815_)begin
        int_reg_array_14_41_real <= _zz_825_;
      end
      if(_zz_816_)begin
        int_reg_array_14_42_real <= _zz_825_;
      end
      if(_zz_817_)begin
        int_reg_array_14_43_real <= _zz_825_;
      end
      if(_zz_818_)begin
        int_reg_array_14_44_real <= _zz_825_;
      end
      if(_zz_819_)begin
        int_reg_array_14_45_real <= _zz_825_;
      end
      if(_zz_820_)begin
        int_reg_array_14_46_real <= _zz_825_;
      end
      if(_zz_821_)begin
        int_reg_array_14_47_real <= _zz_825_;
      end
      if(_zz_822_)begin
        int_reg_array_14_48_real <= _zz_825_;
      end
      if(_zz_823_)begin
        int_reg_array_14_49_real <= _zz_825_;
      end
      if(_zz_774_)begin
        int_reg_array_14_0_imag <= _zz_826_;
      end
      if(_zz_775_)begin
        int_reg_array_14_1_imag <= _zz_826_;
      end
      if(_zz_776_)begin
        int_reg_array_14_2_imag <= _zz_826_;
      end
      if(_zz_777_)begin
        int_reg_array_14_3_imag <= _zz_826_;
      end
      if(_zz_778_)begin
        int_reg_array_14_4_imag <= _zz_826_;
      end
      if(_zz_779_)begin
        int_reg_array_14_5_imag <= _zz_826_;
      end
      if(_zz_780_)begin
        int_reg_array_14_6_imag <= _zz_826_;
      end
      if(_zz_781_)begin
        int_reg_array_14_7_imag <= _zz_826_;
      end
      if(_zz_782_)begin
        int_reg_array_14_8_imag <= _zz_826_;
      end
      if(_zz_783_)begin
        int_reg_array_14_9_imag <= _zz_826_;
      end
      if(_zz_784_)begin
        int_reg_array_14_10_imag <= _zz_826_;
      end
      if(_zz_785_)begin
        int_reg_array_14_11_imag <= _zz_826_;
      end
      if(_zz_786_)begin
        int_reg_array_14_12_imag <= _zz_826_;
      end
      if(_zz_787_)begin
        int_reg_array_14_13_imag <= _zz_826_;
      end
      if(_zz_788_)begin
        int_reg_array_14_14_imag <= _zz_826_;
      end
      if(_zz_789_)begin
        int_reg_array_14_15_imag <= _zz_826_;
      end
      if(_zz_790_)begin
        int_reg_array_14_16_imag <= _zz_826_;
      end
      if(_zz_791_)begin
        int_reg_array_14_17_imag <= _zz_826_;
      end
      if(_zz_792_)begin
        int_reg_array_14_18_imag <= _zz_826_;
      end
      if(_zz_793_)begin
        int_reg_array_14_19_imag <= _zz_826_;
      end
      if(_zz_794_)begin
        int_reg_array_14_20_imag <= _zz_826_;
      end
      if(_zz_795_)begin
        int_reg_array_14_21_imag <= _zz_826_;
      end
      if(_zz_796_)begin
        int_reg_array_14_22_imag <= _zz_826_;
      end
      if(_zz_797_)begin
        int_reg_array_14_23_imag <= _zz_826_;
      end
      if(_zz_798_)begin
        int_reg_array_14_24_imag <= _zz_826_;
      end
      if(_zz_799_)begin
        int_reg_array_14_25_imag <= _zz_826_;
      end
      if(_zz_800_)begin
        int_reg_array_14_26_imag <= _zz_826_;
      end
      if(_zz_801_)begin
        int_reg_array_14_27_imag <= _zz_826_;
      end
      if(_zz_802_)begin
        int_reg_array_14_28_imag <= _zz_826_;
      end
      if(_zz_803_)begin
        int_reg_array_14_29_imag <= _zz_826_;
      end
      if(_zz_804_)begin
        int_reg_array_14_30_imag <= _zz_826_;
      end
      if(_zz_805_)begin
        int_reg_array_14_31_imag <= _zz_826_;
      end
      if(_zz_806_)begin
        int_reg_array_14_32_imag <= _zz_826_;
      end
      if(_zz_807_)begin
        int_reg_array_14_33_imag <= _zz_826_;
      end
      if(_zz_808_)begin
        int_reg_array_14_34_imag <= _zz_826_;
      end
      if(_zz_809_)begin
        int_reg_array_14_35_imag <= _zz_826_;
      end
      if(_zz_810_)begin
        int_reg_array_14_36_imag <= _zz_826_;
      end
      if(_zz_811_)begin
        int_reg_array_14_37_imag <= _zz_826_;
      end
      if(_zz_812_)begin
        int_reg_array_14_38_imag <= _zz_826_;
      end
      if(_zz_813_)begin
        int_reg_array_14_39_imag <= _zz_826_;
      end
      if(_zz_814_)begin
        int_reg_array_14_40_imag <= _zz_826_;
      end
      if(_zz_815_)begin
        int_reg_array_14_41_imag <= _zz_826_;
      end
      if(_zz_816_)begin
        int_reg_array_14_42_imag <= _zz_826_;
      end
      if(_zz_817_)begin
        int_reg_array_14_43_imag <= _zz_826_;
      end
      if(_zz_818_)begin
        int_reg_array_14_44_imag <= _zz_826_;
      end
      if(_zz_819_)begin
        int_reg_array_14_45_imag <= _zz_826_;
      end
      if(_zz_820_)begin
        int_reg_array_14_46_imag <= _zz_826_;
      end
      if(_zz_821_)begin
        int_reg_array_14_47_imag <= _zz_826_;
      end
      if(_zz_822_)begin
        int_reg_array_14_48_imag <= _zz_826_;
      end
      if(_zz_823_)begin
        int_reg_array_14_49_imag <= _zz_826_;
      end
      if(_zz_829_)begin
        int_reg_array_15_0_real <= _zz_880_;
      end
      if(_zz_830_)begin
        int_reg_array_15_1_real <= _zz_880_;
      end
      if(_zz_831_)begin
        int_reg_array_15_2_real <= _zz_880_;
      end
      if(_zz_832_)begin
        int_reg_array_15_3_real <= _zz_880_;
      end
      if(_zz_833_)begin
        int_reg_array_15_4_real <= _zz_880_;
      end
      if(_zz_834_)begin
        int_reg_array_15_5_real <= _zz_880_;
      end
      if(_zz_835_)begin
        int_reg_array_15_6_real <= _zz_880_;
      end
      if(_zz_836_)begin
        int_reg_array_15_7_real <= _zz_880_;
      end
      if(_zz_837_)begin
        int_reg_array_15_8_real <= _zz_880_;
      end
      if(_zz_838_)begin
        int_reg_array_15_9_real <= _zz_880_;
      end
      if(_zz_839_)begin
        int_reg_array_15_10_real <= _zz_880_;
      end
      if(_zz_840_)begin
        int_reg_array_15_11_real <= _zz_880_;
      end
      if(_zz_841_)begin
        int_reg_array_15_12_real <= _zz_880_;
      end
      if(_zz_842_)begin
        int_reg_array_15_13_real <= _zz_880_;
      end
      if(_zz_843_)begin
        int_reg_array_15_14_real <= _zz_880_;
      end
      if(_zz_844_)begin
        int_reg_array_15_15_real <= _zz_880_;
      end
      if(_zz_845_)begin
        int_reg_array_15_16_real <= _zz_880_;
      end
      if(_zz_846_)begin
        int_reg_array_15_17_real <= _zz_880_;
      end
      if(_zz_847_)begin
        int_reg_array_15_18_real <= _zz_880_;
      end
      if(_zz_848_)begin
        int_reg_array_15_19_real <= _zz_880_;
      end
      if(_zz_849_)begin
        int_reg_array_15_20_real <= _zz_880_;
      end
      if(_zz_850_)begin
        int_reg_array_15_21_real <= _zz_880_;
      end
      if(_zz_851_)begin
        int_reg_array_15_22_real <= _zz_880_;
      end
      if(_zz_852_)begin
        int_reg_array_15_23_real <= _zz_880_;
      end
      if(_zz_853_)begin
        int_reg_array_15_24_real <= _zz_880_;
      end
      if(_zz_854_)begin
        int_reg_array_15_25_real <= _zz_880_;
      end
      if(_zz_855_)begin
        int_reg_array_15_26_real <= _zz_880_;
      end
      if(_zz_856_)begin
        int_reg_array_15_27_real <= _zz_880_;
      end
      if(_zz_857_)begin
        int_reg_array_15_28_real <= _zz_880_;
      end
      if(_zz_858_)begin
        int_reg_array_15_29_real <= _zz_880_;
      end
      if(_zz_859_)begin
        int_reg_array_15_30_real <= _zz_880_;
      end
      if(_zz_860_)begin
        int_reg_array_15_31_real <= _zz_880_;
      end
      if(_zz_861_)begin
        int_reg_array_15_32_real <= _zz_880_;
      end
      if(_zz_862_)begin
        int_reg_array_15_33_real <= _zz_880_;
      end
      if(_zz_863_)begin
        int_reg_array_15_34_real <= _zz_880_;
      end
      if(_zz_864_)begin
        int_reg_array_15_35_real <= _zz_880_;
      end
      if(_zz_865_)begin
        int_reg_array_15_36_real <= _zz_880_;
      end
      if(_zz_866_)begin
        int_reg_array_15_37_real <= _zz_880_;
      end
      if(_zz_867_)begin
        int_reg_array_15_38_real <= _zz_880_;
      end
      if(_zz_868_)begin
        int_reg_array_15_39_real <= _zz_880_;
      end
      if(_zz_869_)begin
        int_reg_array_15_40_real <= _zz_880_;
      end
      if(_zz_870_)begin
        int_reg_array_15_41_real <= _zz_880_;
      end
      if(_zz_871_)begin
        int_reg_array_15_42_real <= _zz_880_;
      end
      if(_zz_872_)begin
        int_reg_array_15_43_real <= _zz_880_;
      end
      if(_zz_873_)begin
        int_reg_array_15_44_real <= _zz_880_;
      end
      if(_zz_874_)begin
        int_reg_array_15_45_real <= _zz_880_;
      end
      if(_zz_875_)begin
        int_reg_array_15_46_real <= _zz_880_;
      end
      if(_zz_876_)begin
        int_reg_array_15_47_real <= _zz_880_;
      end
      if(_zz_877_)begin
        int_reg_array_15_48_real <= _zz_880_;
      end
      if(_zz_878_)begin
        int_reg_array_15_49_real <= _zz_880_;
      end
      if(_zz_829_)begin
        int_reg_array_15_0_imag <= _zz_881_;
      end
      if(_zz_830_)begin
        int_reg_array_15_1_imag <= _zz_881_;
      end
      if(_zz_831_)begin
        int_reg_array_15_2_imag <= _zz_881_;
      end
      if(_zz_832_)begin
        int_reg_array_15_3_imag <= _zz_881_;
      end
      if(_zz_833_)begin
        int_reg_array_15_4_imag <= _zz_881_;
      end
      if(_zz_834_)begin
        int_reg_array_15_5_imag <= _zz_881_;
      end
      if(_zz_835_)begin
        int_reg_array_15_6_imag <= _zz_881_;
      end
      if(_zz_836_)begin
        int_reg_array_15_7_imag <= _zz_881_;
      end
      if(_zz_837_)begin
        int_reg_array_15_8_imag <= _zz_881_;
      end
      if(_zz_838_)begin
        int_reg_array_15_9_imag <= _zz_881_;
      end
      if(_zz_839_)begin
        int_reg_array_15_10_imag <= _zz_881_;
      end
      if(_zz_840_)begin
        int_reg_array_15_11_imag <= _zz_881_;
      end
      if(_zz_841_)begin
        int_reg_array_15_12_imag <= _zz_881_;
      end
      if(_zz_842_)begin
        int_reg_array_15_13_imag <= _zz_881_;
      end
      if(_zz_843_)begin
        int_reg_array_15_14_imag <= _zz_881_;
      end
      if(_zz_844_)begin
        int_reg_array_15_15_imag <= _zz_881_;
      end
      if(_zz_845_)begin
        int_reg_array_15_16_imag <= _zz_881_;
      end
      if(_zz_846_)begin
        int_reg_array_15_17_imag <= _zz_881_;
      end
      if(_zz_847_)begin
        int_reg_array_15_18_imag <= _zz_881_;
      end
      if(_zz_848_)begin
        int_reg_array_15_19_imag <= _zz_881_;
      end
      if(_zz_849_)begin
        int_reg_array_15_20_imag <= _zz_881_;
      end
      if(_zz_850_)begin
        int_reg_array_15_21_imag <= _zz_881_;
      end
      if(_zz_851_)begin
        int_reg_array_15_22_imag <= _zz_881_;
      end
      if(_zz_852_)begin
        int_reg_array_15_23_imag <= _zz_881_;
      end
      if(_zz_853_)begin
        int_reg_array_15_24_imag <= _zz_881_;
      end
      if(_zz_854_)begin
        int_reg_array_15_25_imag <= _zz_881_;
      end
      if(_zz_855_)begin
        int_reg_array_15_26_imag <= _zz_881_;
      end
      if(_zz_856_)begin
        int_reg_array_15_27_imag <= _zz_881_;
      end
      if(_zz_857_)begin
        int_reg_array_15_28_imag <= _zz_881_;
      end
      if(_zz_858_)begin
        int_reg_array_15_29_imag <= _zz_881_;
      end
      if(_zz_859_)begin
        int_reg_array_15_30_imag <= _zz_881_;
      end
      if(_zz_860_)begin
        int_reg_array_15_31_imag <= _zz_881_;
      end
      if(_zz_861_)begin
        int_reg_array_15_32_imag <= _zz_881_;
      end
      if(_zz_862_)begin
        int_reg_array_15_33_imag <= _zz_881_;
      end
      if(_zz_863_)begin
        int_reg_array_15_34_imag <= _zz_881_;
      end
      if(_zz_864_)begin
        int_reg_array_15_35_imag <= _zz_881_;
      end
      if(_zz_865_)begin
        int_reg_array_15_36_imag <= _zz_881_;
      end
      if(_zz_866_)begin
        int_reg_array_15_37_imag <= _zz_881_;
      end
      if(_zz_867_)begin
        int_reg_array_15_38_imag <= _zz_881_;
      end
      if(_zz_868_)begin
        int_reg_array_15_39_imag <= _zz_881_;
      end
      if(_zz_869_)begin
        int_reg_array_15_40_imag <= _zz_881_;
      end
      if(_zz_870_)begin
        int_reg_array_15_41_imag <= _zz_881_;
      end
      if(_zz_871_)begin
        int_reg_array_15_42_imag <= _zz_881_;
      end
      if(_zz_872_)begin
        int_reg_array_15_43_imag <= _zz_881_;
      end
      if(_zz_873_)begin
        int_reg_array_15_44_imag <= _zz_881_;
      end
      if(_zz_874_)begin
        int_reg_array_15_45_imag <= _zz_881_;
      end
      if(_zz_875_)begin
        int_reg_array_15_46_imag <= _zz_881_;
      end
      if(_zz_876_)begin
        int_reg_array_15_47_imag <= _zz_881_;
      end
      if(_zz_877_)begin
        int_reg_array_15_48_imag <= _zz_881_;
      end
      if(_zz_878_)begin
        int_reg_array_15_49_imag <= _zz_881_;
      end
      if(_zz_884_)begin
        int_reg_array_16_0_real <= _zz_935_;
      end
      if(_zz_885_)begin
        int_reg_array_16_1_real <= _zz_935_;
      end
      if(_zz_886_)begin
        int_reg_array_16_2_real <= _zz_935_;
      end
      if(_zz_887_)begin
        int_reg_array_16_3_real <= _zz_935_;
      end
      if(_zz_888_)begin
        int_reg_array_16_4_real <= _zz_935_;
      end
      if(_zz_889_)begin
        int_reg_array_16_5_real <= _zz_935_;
      end
      if(_zz_890_)begin
        int_reg_array_16_6_real <= _zz_935_;
      end
      if(_zz_891_)begin
        int_reg_array_16_7_real <= _zz_935_;
      end
      if(_zz_892_)begin
        int_reg_array_16_8_real <= _zz_935_;
      end
      if(_zz_893_)begin
        int_reg_array_16_9_real <= _zz_935_;
      end
      if(_zz_894_)begin
        int_reg_array_16_10_real <= _zz_935_;
      end
      if(_zz_895_)begin
        int_reg_array_16_11_real <= _zz_935_;
      end
      if(_zz_896_)begin
        int_reg_array_16_12_real <= _zz_935_;
      end
      if(_zz_897_)begin
        int_reg_array_16_13_real <= _zz_935_;
      end
      if(_zz_898_)begin
        int_reg_array_16_14_real <= _zz_935_;
      end
      if(_zz_899_)begin
        int_reg_array_16_15_real <= _zz_935_;
      end
      if(_zz_900_)begin
        int_reg_array_16_16_real <= _zz_935_;
      end
      if(_zz_901_)begin
        int_reg_array_16_17_real <= _zz_935_;
      end
      if(_zz_902_)begin
        int_reg_array_16_18_real <= _zz_935_;
      end
      if(_zz_903_)begin
        int_reg_array_16_19_real <= _zz_935_;
      end
      if(_zz_904_)begin
        int_reg_array_16_20_real <= _zz_935_;
      end
      if(_zz_905_)begin
        int_reg_array_16_21_real <= _zz_935_;
      end
      if(_zz_906_)begin
        int_reg_array_16_22_real <= _zz_935_;
      end
      if(_zz_907_)begin
        int_reg_array_16_23_real <= _zz_935_;
      end
      if(_zz_908_)begin
        int_reg_array_16_24_real <= _zz_935_;
      end
      if(_zz_909_)begin
        int_reg_array_16_25_real <= _zz_935_;
      end
      if(_zz_910_)begin
        int_reg_array_16_26_real <= _zz_935_;
      end
      if(_zz_911_)begin
        int_reg_array_16_27_real <= _zz_935_;
      end
      if(_zz_912_)begin
        int_reg_array_16_28_real <= _zz_935_;
      end
      if(_zz_913_)begin
        int_reg_array_16_29_real <= _zz_935_;
      end
      if(_zz_914_)begin
        int_reg_array_16_30_real <= _zz_935_;
      end
      if(_zz_915_)begin
        int_reg_array_16_31_real <= _zz_935_;
      end
      if(_zz_916_)begin
        int_reg_array_16_32_real <= _zz_935_;
      end
      if(_zz_917_)begin
        int_reg_array_16_33_real <= _zz_935_;
      end
      if(_zz_918_)begin
        int_reg_array_16_34_real <= _zz_935_;
      end
      if(_zz_919_)begin
        int_reg_array_16_35_real <= _zz_935_;
      end
      if(_zz_920_)begin
        int_reg_array_16_36_real <= _zz_935_;
      end
      if(_zz_921_)begin
        int_reg_array_16_37_real <= _zz_935_;
      end
      if(_zz_922_)begin
        int_reg_array_16_38_real <= _zz_935_;
      end
      if(_zz_923_)begin
        int_reg_array_16_39_real <= _zz_935_;
      end
      if(_zz_924_)begin
        int_reg_array_16_40_real <= _zz_935_;
      end
      if(_zz_925_)begin
        int_reg_array_16_41_real <= _zz_935_;
      end
      if(_zz_926_)begin
        int_reg_array_16_42_real <= _zz_935_;
      end
      if(_zz_927_)begin
        int_reg_array_16_43_real <= _zz_935_;
      end
      if(_zz_928_)begin
        int_reg_array_16_44_real <= _zz_935_;
      end
      if(_zz_929_)begin
        int_reg_array_16_45_real <= _zz_935_;
      end
      if(_zz_930_)begin
        int_reg_array_16_46_real <= _zz_935_;
      end
      if(_zz_931_)begin
        int_reg_array_16_47_real <= _zz_935_;
      end
      if(_zz_932_)begin
        int_reg_array_16_48_real <= _zz_935_;
      end
      if(_zz_933_)begin
        int_reg_array_16_49_real <= _zz_935_;
      end
      if(_zz_884_)begin
        int_reg_array_16_0_imag <= _zz_936_;
      end
      if(_zz_885_)begin
        int_reg_array_16_1_imag <= _zz_936_;
      end
      if(_zz_886_)begin
        int_reg_array_16_2_imag <= _zz_936_;
      end
      if(_zz_887_)begin
        int_reg_array_16_3_imag <= _zz_936_;
      end
      if(_zz_888_)begin
        int_reg_array_16_4_imag <= _zz_936_;
      end
      if(_zz_889_)begin
        int_reg_array_16_5_imag <= _zz_936_;
      end
      if(_zz_890_)begin
        int_reg_array_16_6_imag <= _zz_936_;
      end
      if(_zz_891_)begin
        int_reg_array_16_7_imag <= _zz_936_;
      end
      if(_zz_892_)begin
        int_reg_array_16_8_imag <= _zz_936_;
      end
      if(_zz_893_)begin
        int_reg_array_16_9_imag <= _zz_936_;
      end
      if(_zz_894_)begin
        int_reg_array_16_10_imag <= _zz_936_;
      end
      if(_zz_895_)begin
        int_reg_array_16_11_imag <= _zz_936_;
      end
      if(_zz_896_)begin
        int_reg_array_16_12_imag <= _zz_936_;
      end
      if(_zz_897_)begin
        int_reg_array_16_13_imag <= _zz_936_;
      end
      if(_zz_898_)begin
        int_reg_array_16_14_imag <= _zz_936_;
      end
      if(_zz_899_)begin
        int_reg_array_16_15_imag <= _zz_936_;
      end
      if(_zz_900_)begin
        int_reg_array_16_16_imag <= _zz_936_;
      end
      if(_zz_901_)begin
        int_reg_array_16_17_imag <= _zz_936_;
      end
      if(_zz_902_)begin
        int_reg_array_16_18_imag <= _zz_936_;
      end
      if(_zz_903_)begin
        int_reg_array_16_19_imag <= _zz_936_;
      end
      if(_zz_904_)begin
        int_reg_array_16_20_imag <= _zz_936_;
      end
      if(_zz_905_)begin
        int_reg_array_16_21_imag <= _zz_936_;
      end
      if(_zz_906_)begin
        int_reg_array_16_22_imag <= _zz_936_;
      end
      if(_zz_907_)begin
        int_reg_array_16_23_imag <= _zz_936_;
      end
      if(_zz_908_)begin
        int_reg_array_16_24_imag <= _zz_936_;
      end
      if(_zz_909_)begin
        int_reg_array_16_25_imag <= _zz_936_;
      end
      if(_zz_910_)begin
        int_reg_array_16_26_imag <= _zz_936_;
      end
      if(_zz_911_)begin
        int_reg_array_16_27_imag <= _zz_936_;
      end
      if(_zz_912_)begin
        int_reg_array_16_28_imag <= _zz_936_;
      end
      if(_zz_913_)begin
        int_reg_array_16_29_imag <= _zz_936_;
      end
      if(_zz_914_)begin
        int_reg_array_16_30_imag <= _zz_936_;
      end
      if(_zz_915_)begin
        int_reg_array_16_31_imag <= _zz_936_;
      end
      if(_zz_916_)begin
        int_reg_array_16_32_imag <= _zz_936_;
      end
      if(_zz_917_)begin
        int_reg_array_16_33_imag <= _zz_936_;
      end
      if(_zz_918_)begin
        int_reg_array_16_34_imag <= _zz_936_;
      end
      if(_zz_919_)begin
        int_reg_array_16_35_imag <= _zz_936_;
      end
      if(_zz_920_)begin
        int_reg_array_16_36_imag <= _zz_936_;
      end
      if(_zz_921_)begin
        int_reg_array_16_37_imag <= _zz_936_;
      end
      if(_zz_922_)begin
        int_reg_array_16_38_imag <= _zz_936_;
      end
      if(_zz_923_)begin
        int_reg_array_16_39_imag <= _zz_936_;
      end
      if(_zz_924_)begin
        int_reg_array_16_40_imag <= _zz_936_;
      end
      if(_zz_925_)begin
        int_reg_array_16_41_imag <= _zz_936_;
      end
      if(_zz_926_)begin
        int_reg_array_16_42_imag <= _zz_936_;
      end
      if(_zz_927_)begin
        int_reg_array_16_43_imag <= _zz_936_;
      end
      if(_zz_928_)begin
        int_reg_array_16_44_imag <= _zz_936_;
      end
      if(_zz_929_)begin
        int_reg_array_16_45_imag <= _zz_936_;
      end
      if(_zz_930_)begin
        int_reg_array_16_46_imag <= _zz_936_;
      end
      if(_zz_931_)begin
        int_reg_array_16_47_imag <= _zz_936_;
      end
      if(_zz_932_)begin
        int_reg_array_16_48_imag <= _zz_936_;
      end
      if(_zz_933_)begin
        int_reg_array_16_49_imag <= _zz_936_;
      end
      if(_zz_939_)begin
        int_reg_array_17_0_real <= _zz_990_;
      end
      if(_zz_940_)begin
        int_reg_array_17_1_real <= _zz_990_;
      end
      if(_zz_941_)begin
        int_reg_array_17_2_real <= _zz_990_;
      end
      if(_zz_942_)begin
        int_reg_array_17_3_real <= _zz_990_;
      end
      if(_zz_943_)begin
        int_reg_array_17_4_real <= _zz_990_;
      end
      if(_zz_944_)begin
        int_reg_array_17_5_real <= _zz_990_;
      end
      if(_zz_945_)begin
        int_reg_array_17_6_real <= _zz_990_;
      end
      if(_zz_946_)begin
        int_reg_array_17_7_real <= _zz_990_;
      end
      if(_zz_947_)begin
        int_reg_array_17_8_real <= _zz_990_;
      end
      if(_zz_948_)begin
        int_reg_array_17_9_real <= _zz_990_;
      end
      if(_zz_949_)begin
        int_reg_array_17_10_real <= _zz_990_;
      end
      if(_zz_950_)begin
        int_reg_array_17_11_real <= _zz_990_;
      end
      if(_zz_951_)begin
        int_reg_array_17_12_real <= _zz_990_;
      end
      if(_zz_952_)begin
        int_reg_array_17_13_real <= _zz_990_;
      end
      if(_zz_953_)begin
        int_reg_array_17_14_real <= _zz_990_;
      end
      if(_zz_954_)begin
        int_reg_array_17_15_real <= _zz_990_;
      end
      if(_zz_955_)begin
        int_reg_array_17_16_real <= _zz_990_;
      end
      if(_zz_956_)begin
        int_reg_array_17_17_real <= _zz_990_;
      end
      if(_zz_957_)begin
        int_reg_array_17_18_real <= _zz_990_;
      end
      if(_zz_958_)begin
        int_reg_array_17_19_real <= _zz_990_;
      end
      if(_zz_959_)begin
        int_reg_array_17_20_real <= _zz_990_;
      end
      if(_zz_960_)begin
        int_reg_array_17_21_real <= _zz_990_;
      end
      if(_zz_961_)begin
        int_reg_array_17_22_real <= _zz_990_;
      end
      if(_zz_962_)begin
        int_reg_array_17_23_real <= _zz_990_;
      end
      if(_zz_963_)begin
        int_reg_array_17_24_real <= _zz_990_;
      end
      if(_zz_964_)begin
        int_reg_array_17_25_real <= _zz_990_;
      end
      if(_zz_965_)begin
        int_reg_array_17_26_real <= _zz_990_;
      end
      if(_zz_966_)begin
        int_reg_array_17_27_real <= _zz_990_;
      end
      if(_zz_967_)begin
        int_reg_array_17_28_real <= _zz_990_;
      end
      if(_zz_968_)begin
        int_reg_array_17_29_real <= _zz_990_;
      end
      if(_zz_969_)begin
        int_reg_array_17_30_real <= _zz_990_;
      end
      if(_zz_970_)begin
        int_reg_array_17_31_real <= _zz_990_;
      end
      if(_zz_971_)begin
        int_reg_array_17_32_real <= _zz_990_;
      end
      if(_zz_972_)begin
        int_reg_array_17_33_real <= _zz_990_;
      end
      if(_zz_973_)begin
        int_reg_array_17_34_real <= _zz_990_;
      end
      if(_zz_974_)begin
        int_reg_array_17_35_real <= _zz_990_;
      end
      if(_zz_975_)begin
        int_reg_array_17_36_real <= _zz_990_;
      end
      if(_zz_976_)begin
        int_reg_array_17_37_real <= _zz_990_;
      end
      if(_zz_977_)begin
        int_reg_array_17_38_real <= _zz_990_;
      end
      if(_zz_978_)begin
        int_reg_array_17_39_real <= _zz_990_;
      end
      if(_zz_979_)begin
        int_reg_array_17_40_real <= _zz_990_;
      end
      if(_zz_980_)begin
        int_reg_array_17_41_real <= _zz_990_;
      end
      if(_zz_981_)begin
        int_reg_array_17_42_real <= _zz_990_;
      end
      if(_zz_982_)begin
        int_reg_array_17_43_real <= _zz_990_;
      end
      if(_zz_983_)begin
        int_reg_array_17_44_real <= _zz_990_;
      end
      if(_zz_984_)begin
        int_reg_array_17_45_real <= _zz_990_;
      end
      if(_zz_985_)begin
        int_reg_array_17_46_real <= _zz_990_;
      end
      if(_zz_986_)begin
        int_reg_array_17_47_real <= _zz_990_;
      end
      if(_zz_987_)begin
        int_reg_array_17_48_real <= _zz_990_;
      end
      if(_zz_988_)begin
        int_reg_array_17_49_real <= _zz_990_;
      end
      if(_zz_939_)begin
        int_reg_array_17_0_imag <= _zz_991_;
      end
      if(_zz_940_)begin
        int_reg_array_17_1_imag <= _zz_991_;
      end
      if(_zz_941_)begin
        int_reg_array_17_2_imag <= _zz_991_;
      end
      if(_zz_942_)begin
        int_reg_array_17_3_imag <= _zz_991_;
      end
      if(_zz_943_)begin
        int_reg_array_17_4_imag <= _zz_991_;
      end
      if(_zz_944_)begin
        int_reg_array_17_5_imag <= _zz_991_;
      end
      if(_zz_945_)begin
        int_reg_array_17_6_imag <= _zz_991_;
      end
      if(_zz_946_)begin
        int_reg_array_17_7_imag <= _zz_991_;
      end
      if(_zz_947_)begin
        int_reg_array_17_8_imag <= _zz_991_;
      end
      if(_zz_948_)begin
        int_reg_array_17_9_imag <= _zz_991_;
      end
      if(_zz_949_)begin
        int_reg_array_17_10_imag <= _zz_991_;
      end
      if(_zz_950_)begin
        int_reg_array_17_11_imag <= _zz_991_;
      end
      if(_zz_951_)begin
        int_reg_array_17_12_imag <= _zz_991_;
      end
      if(_zz_952_)begin
        int_reg_array_17_13_imag <= _zz_991_;
      end
      if(_zz_953_)begin
        int_reg_array_17_14_imag <= _zz_991_;
      end
      if(_zz_954_)begin
        int_reg_array_17_15_imag <= _zz_991_;
      end
      if(_zz_955_)begin
        int_reg_array_17_16_imag <= _zz_991_;
      end
      if(_zz_956_)begin
        int_reg_array_17_17_imag <= _zz_991_;
      end
      if(_zz_957_)begin
        int_reg_array_17_18_imag <= _zz_991_;
      end
      if(_zz_958_)begin
        int_reg_array_17_19_imag <= _zz_991_;
      end
      if(_zz_959_)begin
        int_reg_array_17_20_imag <= _zz_991_;
      end
      if(_zz_960_)begin
        int_reg_array_17_21_imag <= _zz_991_;
      end
      if(_zz_961_)begin
        int_reg_array_17_22_imag <= _zz_991_;
      end
      if(_zz_962_)begin
        int_reg_array_17_23_imag <= _zz_991_;
      end
      if(_zz_963_)begin
        int_reg_array_17_24_imag <= _zz_991_;
      end
      if(_zz_964_)begin
        int_reg_array_17_25_imag <= _zz_991_;
      end
      if(_zz_965_)begin
        int_reg_array_17_26_imag <= _zz_991_;
      end
      if(_zz_966_)begin
        int_reg_array_17_27_imag <= _zz_991_;
      end
      if(_zz_967_)begin
        int_reg_array_17_28_imag <= _zz_991_;
      end
      if(_zz_968_)begin
        int_reg_array_17_29_imag <= _zz_991_;
      end
      if(_zz_969_)begin
        int_reg_array_17_30_imag <= _zz_991_;
      end
      if(_zz_970_)begin
        int_reg_array_17_31_imag <= _zz_991_;
      end
      if(_zz_971_)begin
        int_reg_array_17_32_imag <= _zz_991_;
      end
      if(_zz_972_)begin
        int_reg_array_17_33_imag <= _zz_991_;
      end
      if(_zz_973_)begin
        int_reg_array_17_34_imag <= _zz_991_;
      end
      if(_zz_974_)begin
        int_reg_array_17_35_imag <= _zz_991_;
      end
      if(_zz_975_)begin
        int_reg_array_17_36_imag <= _zz_991_;
      end
      if(_zz_976_)begin
        int_reg_array_17_37_imag <= _zz_991_;
      end
      if(_zz_977_)begin
        int_reg_array_17_38_imag <= _zz_991_;
      end
      if(_zz_978_)begin
        int_reg_array_17_39_imag <= _zz_991_;
      end
      if(_zz_979_)begin
        int_reg_array_17_40_imag <= _zz_991_;
      end
      if(_zz_980_)begin
        int_reg_array_17_41_imag <= _zz_991_;
      end
      if(_zz_981_)begin
        int_reg_array_17_42_imag <= _zz_991_;
      end
      if(_zz_982_)begin
        int_reg_array_17_43_imag <= _zz_991_;
      end
      if(_zz_983_)begin
        int_reg_array_17_44_imag <= _zz_991_;
      end
      if(_zz_984_)begin
        int_reg_array_17_45_imag <= _zz_991_;
      end
      if(_zz_985_)begin
        int_reg_array_17_46_imag <= _zz_991_;
      end
      if(_zz_986_)begin
        int_reg_array_17_47_imag <= _zz_991_;
      end
      if(_zz_987_)begin
        int_reg_array_17_48_imag <= _zz_991_;
      end
      if(_zz_988_)begin
        int_reg_array_17_49_imag <= _zz_991_;
      end
      if(_zz_994_)begin
        int_reg_array_18_0_real <= _zz_1045_;
      end
      if(_zz_995_)begin
        int_reg_array_18_1_real <= _zz_1045_;
      end
      if(_zz_996_)begin
        int_reg_array_18_2_real <= _zz_1045_;
      end
      if(_zz_997_)begin
        int_reg_array_18_3_real <= _zz_1045_;
      end
      if(_zz_998_)begin
        int_reg_array_18_4_real <= _zz_1045_;
      end
      if(_zz_999_)begin
        int_reg_array_18_5_real <= _zz_1045_;
      end
      if(_zz_1000_)begin
        int_reg_array_18_6_real <= _zz_1045_;
      end
      if(_zz_1001_)begin
        int_reg_array_18_7_real <= _zz_1045_;
      end
      if(_zz_1002_)begin
        int_reg_array_18_8_real <= _zz_1045_;
      end
      if(_zz_1003_)begin
        int_reg_array_18_9_real <= _zz_1045_;
      end
      if(_zz_1004_)begin
        int_reg_array_18_10_real <= _zz_1045_;
      end
      if(_zz_1005_)begin
        int_reg_array_18_11_real <= _zz_1045_;
      end
      if(_zz_1006_)begin
        int_reg_array_18_12_real <= _zz_1045_;
      end
      if(_zz_1007_)begin
        int_reg_array_18_13_real <= _zz_1045_;
      end
      if(_zz_1008_)begin
        int_reg_array_18_14_real <= _zz_1045_;
      end
      if(_zz_1009_)begin
        int_reg_array_18_15_real <= _zz_1045_;
      end
      if(_zz_1010_)begin
        int_reg_array_18_16_real <= _zz_1045_;
      end
      if(_zz_1011_)begin
        int_reg_array_18_17_real <= _zz_1045_;
      end
      if(_zz_1012_)begin
        int_reg_array_18_18_real <= _zz_1045_;
      end
      if(_zz_1013_)begin
        int_reg_array_18_19_real <= _zz_1045_;
      end
      if(_zz_1014_)begin
        int_reg_array_18_20_real <= _zz_1045_;
      end
      if(_zz_1015_)begin
        int_reg_array_18_21_real <= _zz_1045_;
      end
      if(_zz_1016_)begin
        int_reg_array_18_22_real <= _zz_1045_;
      end
      if(_zz_1017_)begin
        int_reg_array_18_23_real <= _zz_1045_;
      end
      if(_zz_1018_)begin
        int_reg_array_18_24_real <= _zz_1045_;
      end
      if(_zz_1019_)begin
        int_reg_array_18_25_real <= _zz_1045_;
      end
      if(_zz_1020_)begin
        int_reg_array_18_26_real <= _zz_1045_;
      end
      if(_zz_1021_)begin
        int_reg_array_18_27_real <= _zz_1045_;
      end
      if(_zz_1022_)begin
        int_reg_array_18_28_real <= _zz_1045_;
      end
      if(_zz_1023_)begin
        int_reg_array_18_29_real <= _zz_1045_;
      end
      if(_zz_1024_)begin
        int_reg_array_18_30_real <= _zz_1045_;
      end
      if(_zz_1025_)begin
        int_reg_array_18_31_real <= _zz_1045_;
      end
      if(_zz_1026_)begin
        int_reg_array_18_32_real <= _zz_1045_;
      end
      if(_zz_1027_)begin
        int_reg_array_18_33_real <= _zz_1045_;
      end
      if(_zz_1028_)begin
        int_reg_array_18_34_real <= _zz_1045_;
      end
      if(_zz_1029_)begin
        int_reg_array_18_35_real <= _zz_1045_;
      end
      if(_zz_1030_)begin
        int_reg_array_18_36_real <= _zz_1045_;
      end
      if(_zz_1031_)begin
        int_reg_array_18_37_real <= _zz_1045_;
      end
      if(_zz_1032_)begin
        int_reg_array_18_38_real <= _zz_1045_;
      end
      if(_zz_1033_)begin
        int_reg_array_18_39_real <= _zz_1045_;
      end
      if(_zz_1034_)begin
        int_reg_array_18_40_real <= _zz_1045_;
      end
      if(_zz_1035_)begin
        int_reg_array_18_41_real <= _zz_1045_;
      end
      if(_zz_1036_)begin
        int_reg_array_18_42_real <= _zz_1045_;
      end
      if(_zz_1037_)begin
        int_reg_array_18_43_real <= _zz_1045_;
      end
      if(_zz_1038_)begin
        int_reg_array_18_44_real <= _zz_1045_;
      end
      if(_zz_1039_)begin
        int_reg_array_18_45_real <= _zz_1045_;
      end
      if(_zz_1040_)begin
        int_reg_array_18_46_real <= _zz_1045_;
      end
      if(_zz_1041_)begin
        int_reg_array_18_47_real <= _zz_1045_;
      end
      if(_zz_1042_)begin
        int_reg_array_18_48_real <= _zz_1045_;
      end
      if(_zz_1043_)begin
        int_reg_array_18_49_real <= _zz_1045_;
      end
      if(_zz_994_)begin
        int_reg_array_18_0_imag <= _zz_1046_;
      end
      if(_zz_995_)begin
        int_reg_array_18_1_imag <= _zz_1046_;
      end
      if(_zz_996_)begin
        int_reg_array_18_2_imag <= _zz_1046_;
      end
      if(_zz_997_)begin
        int_reg_array_18_3_imag <= _zz_1046_;
      end
      if(_zz_998_)begin
        int_reg_array_18_4_imag <= _zz_1046_;
      end
      if(_zz_999_)begin
        int_reg_array_18_5_imag <= _zz_1046_;
      end
      if(_zz_1000_)begin
        int_reg_array_18_6_imag <= _zz_1046_;
      end
      if(_zz_1001_)begin
        int_reg_array_18_7_imag <= _zz_1046_;
      end
      if(_zz_1002_)begin
        int_reg_array_18_8_imag <= _zz_1046_;
      end
      if(_zz_1003_)begin
        int_reg_array_18_9_imag <= _zz_1046_;
      end
      if(_zz_1004_)begin
        int_reg_array_18_10_imag <= _zz_1046_;
      end
      if(_zz_1005_)begin
        int_reg_array_18_11_imag <= _zz_1046_;
      end
      if(_zz_1006_)begin
        int_reg_array_18_12_imag <= _zz_1046_;
      end
      if(_zz_1007_)begin
        int_reg_array_18_13_imag <= _zz_1046_;
      end
      if(_zz_1008_)begin
        int_reg_array_18_14_imag <= _zz_1046_;
      end
      if(_zz_1009_)begin
        int_reg_array_18_15_imag <= _zz_1046_;
      end
      if(_zz_1010_)begin
        int_reg_array_18_16_imag <= _zz_1046_;
      end
      if(_zz_1011_)begin
        int_reg_array_18_17_imag <= _zz_1046_;
      end
      if(_zz_1012_)begin
        int_reg_array_18_18_imag <= _zz_1046_;
      end
      if(_zz_1013_)begin
        int_reg_array_18_19_imag <= _zz_1046_;
      end
      if(_zz_1014_)begin
        int_reg_array_18_20_imag <= _zz_1046_;
      end
      if(_zz_1015_)begin
        int_reg_array_18_21_imag <= _zz_1046_;
      end
      if(_zz_1016_)begin
        int_reg_array_18_22_imag <= _zz_1046_;
      end
      if(_zz_1017_)begin
        int_reg_array_18_23_imag <= _zz_1046_;
      end
      if(_zz_1018_)begin
        int_reg_array_18_24_imag <= _zz_1046_;
      end
      if(_zz_1019_)begin
        int_reg_array_18_25_imag <= _zz_1046_;
      end
      if(_zz_1020_)begin
        int_reg_array_18_26_imag <= _zz_1046_;
      end
      if(_zz_1021_)begin
        int_reg_array_18_27_imag <= _zz_1046_;
      end
      if(_zz_1022_)begin
        int_reg_array_18_28_imag <= _zz_1046_;
      end
      if(_zz_1023_)begin
        int_reg_array_18_29_imag <= _zz_1046_;
      end
      if(_zz_1024_)begin
        int_reg_array_18_30_imag <= _zz_1046_;
      end
      if(_zz_1025_)begin
        int_reg_array_18_31_imag <= _zz_1046_;
      end
      if(_zz_1026_)begin
        int_reg_array_18_32_imag <= _zz_1046_;
      end
      if(_zz_1027_)begin
        int_reg_array_18_33_imag <= _zz_1046_;
      end
      if(_zz_1028_)begin
        int_reg_array_18_34_imag <= _zz_1046_;
      end
      if(_zz_1029_)begin
        int_reg_array_18_35_imag <= _zz_1046_;
      end
      if(_zz_1030_)begin
        int_reg_array_18_36_imag <= _zz_1046_;
      end
      if(_zz_1031_)begin
        int_reg_array_18_37_imag <= _zz_1046_;
      end
      if(_zz_1032_)begin
        int_reg_array_18_38_imag <= _zz_1046_;
      end
      if(_zz_1033_)begin
        int_reg_array_18_39_imag <= _zz_1046_;
      end
      if(_zz_1034_)begin
        int_reg_array_18_40_imag <= _zz_1046_;
      end
      if(_zz_1035_)begin
        int_reg_array_18_41_imag <= _zz_1046_;
      end
      if(_zz_1036_)begin
        int_reg_array_18_42_imag <= _zz_1046_;
      end
      if(_zz_1037_)begin
        int_reg_array_18_43_imag <= _zz_1046_;
      end
      if(_zz_1038_)begin
        int_reg_array_18_44_imag <= _zz_1046_;
      end
      if(_zz_1039_)begin
        int_reg_array_18_45_imag <= _zz_1046_;
      end
      if(_zz_1040_)begin
        int_reg_array_18_46_imag <= _zz_1046_;
      end
      if(_zz_1041_)begin
        int_reg_array_18_47_imag <= _zz_1046_;
      end
      if(_zz_1042_)begin
        int_reg_array_18_48_imag <= _zz_1046_;
      end
      if(_zz_1043_)begin
        int_reg_array_18_49_imag <= _zz_1046_;
      end
      if(_zz_1049_)begin
        int_reg_array_19_0_real <= _zz_1100_;
      end
      if(_zz_1050_)begin
        int_reg_array_19_1_real <= _zz_1100_;
      end
      if(_zz_1051_)begin
        int_reg_array_19_2_real <= _zz_1100_;
      end
      if(_zz_1052_)begin
        int_reg_array_19_3_real <= _zz_1100_;
      end
      if(_zz_1053_)begin
        int_reg_array_19_4_real <= _zz_1100_;
      end
      if(_zz_1054_)begin
        int_reg_array_19_5_real <= _zz_1100_;
      end
      if(_zz_1055_)begin
        int_reg_array_19_6_real <= _zz_1100_;
      end
      if(_zz_1056_)begin
        int_reg_array_19_7_real <= _zz_1100_;
      end
      if(_zz_1057_)begin
        int_reg_array_19_8_real <= _zz_1100_;
      end
      if(_zz_1058_)begin
        int_reg_array_19_9_real <= _zz_1100_;
      end
      if(_zz_1059_)begin
        int_reg_array_19_10_real <= _zz_1100_;
      end
      if(_zz_1060_)begin
        int_reg_array_19_11_real <= _zz_1100_;
      end
      if(_zz_1061_)begin
        int_reg_array_19_12_real <= _zz_1100_;
      end
      if(_zz_1062_)begin
        int_reg_array_19_13_real <= _zz_1100_;
      end
      if(_zz_1063_)begin
        int_reg_array_19_14_real <= _zz_1100_;
      end
      if(_zz_1064_)begin
        int_reg_array_19_15_real <= _zz_1100_;
      end
      if(_zz_1065_)begin
        int_reg_array_19_16_real <= _zz_1100_;
      end
      if(_zz_1066_)begin
        int_reg_array_19_17_real <= _zz_1100_;
      end
      if(_zz_1067_)begin
        int_reg_array_19_18_real <= _zz_1100_;
      end
      if(_zz_1068_)begin
        int_reg_array_19_19_real <= _zz_1100_;
      end
      if(_zz_1069_)begin
        int_reg_array_19_20_real <= _zz_1100_;
      end
      if(_zz_1070_)begin
        int_reg_array_19_21_real <= _zz_1100_;
      end
      if(_zz_1071_)begin
        int_reg_array_19_22_real <= _zz_1100_;
      end
      if(_zz_1072_)begin
        int_reg_array_19_23_real <= _zz_1100_;
      end
      if(_zz_1073_)begin
        int_reg_array_19_24_real <= _zz_1100_;
      end
      if(_zz_1074_)begin
        int_reg_array_19_25_real <= _zz_1100_;
      end
      if(_zz_1075_)begin
        int_reg_array_19_26_real <= _zz_1100_;
      end
      if(_zz_1076_)begin
        int_reg_array_19_27_real <= _zz_1100_;
      end
      if(_zz_1077_)begin
        int_reg_array_19_28_real <= _zz_1100_;
      end
      if(_zz_1078_)begin
        int_reg_array_19_29_real <= _zz_1100_;
      end
      if(_zz_1079_)begin
        int_reg_array_19_30_real <= _zz_1100_;
      end
      if(_zz_1080_)begin
        int_reg_array_19_31_real <= _zz_1100_;
      end
      if(_zz_1081_)begin
        int_reg_array_19_32_real <= _zz_1100_;
      end
      if(_zz_1082_)begin
        int_reg_array_19_33_real <= _zz_1100_;
      end
      if(_zz_1083_)begin
        int_reg_array_19_34_real <= _zz_1100_;
      end
      if(_zz_1084_)begin
        int_reg_array_19_35_real <= _zz_1100_;
      end
      if(_zz_1085_)begin
        int_reg_array_19_36_real <= _zz_1100_;
      end
      if(_zz_1086_)begin
        int_reg_array_19_37_real <= _zz_1100_;
      end
      if(_zz_1087_)begin
        int_reg_array_19_38_real <= _zz_1100_;
      end
      if(_zz_1088_)begin
        int_reg_array_19_39_real <= _zz_1100_;
      end
      if(_zz_1089_)begin
        int_reg_array_19_40_real <= _zz_1100_;
      end
      if(_zz_1090_)begin
        int_reg_array_19_41_real <= _zz_1100_;
      end
      if(_zz_1091_)begin
        int_reg_array_19_42_real <= _zz_1100_;
      end
      if(_zz_1092_)begin
        int_reg_array_19_43_real <= _zz_1100_;
      end
      if(_zz_1093_)begin
        int_reg_array_19_44_real <= _zz_1100_;
      end
      if(_zz_1094_)begin
        int_reg_array_19_45_real <= _zz_1100_;
      end
      if(_zz_1095_)begin
        int_reg_array_19_46_real <= _zz_1100_;
      end
      if(_zz_1096_)begin
        int_reg_array_19_47_real <= _zz_1100_;
      end
      if(_zz_1097_)begin
        int_reg_array_19_48_real <= _zz_1100_;
      end
      if(_zz_1098_)begin
        int_reg_array_19_49_real <= _zz_1100_;
      end
      if(_zz_1049_)begin
        int_reg_array_19_0_imag <= _zz_1101_;
      end
      if(_zz_1050_)begin
        int_reg_array_19_1_imag <= _zz_1101_;
      end
      if(_zz_1051_)begin
        int_reg_array_19_2_imag <= _zz_1101_;
      end
      if(_zz_1052_)begin
        int_reg_array_19_3_imag <= _zz_1101_;
      end
      if(_zz_1053_)begin
        int_reg_array_19_4_imag <= _zz_1101_;
      end
      if(_zz_1054_)begin
        int_reg_array_19_5_imag <= _zz_1101_;
      end
      if(_zz_1055_)begin
        int_reg_array_19_6_imag <= _zz_1101_;
      end
      if(_zz_1056_)begin
        int_reg_array_19_7_imag <= _zz_1101_;
      end
      if(_zz_1057_)begin
        int_reg_array_19_8_imag <= _zz_1101_;
      end
      if(_zz_1058_)begin
        int_reg_array_19_9_imag <= _zz_1101_;
      end
      if(_zz_1059_)begin
        int_reg_array_19_10_imag <= _zz_1101_;
      end
      if(_zz_1060_)begin
        int_reg_array_19_11_imag <= _zz_1101_;
      end
      if(_zz_1061_)begin
        int_reg_array_19_12_imag <= _zz_1101_;
      end
      if(_zz_1062_)begin
        int_reg_array_19_13_imag <= _zz_1101_;
      end
      if(_zz_1063_)begin
        int_reg_array_19_14_imag <= _zz_1101_;
      end
      if(_zz_1064_)begin
        int_reg_array_19_15_imag <= _zz_1101_;
      end
      if(_zz_1065_)begin
        int_reg_array_19_16_imag <= _zz_1101_;
      end
      if(_zz_1066_)begin
        int_reg_array_19_17_imag <= _zz_1101_;
      end
      if(_zz_1067_)begin
        int_reg_array_19_18_imag <= _zz_1101_;
      end
      if(_zz_1068_)begin
        int_reg_array_19_19_imag <= _zz_1101_;
      end
      if(_zz_1069_)begin
        int_reg_array_19_20_imag <= _zz_1101_;
      end
      if(_zz_1070_)begin
        int_reg_array_19_21_imag <= _zz_1101_;
      end
      if(_zz_1071_)begin
        int_reg_array_19_22_imag <= _zz_1101_;
      end
      if(_zz_1072_)begin
        int_reg_array_19_23_imag <= _zz_1101_;
      end
      if(_zz_1073_)begin
        int_reg_array_19_24_imag <= _zz_1101_;
      end
      if(_zz_1074_)begin
        int_reg_array_19_25_imag <= _zz_1101_;
      end
      if(_zz_1075_)begin
        int_reg_array_19_26_imag <= _zz_1101_;
      end
      if(_zz_1076_)begin
        int_reg_array_19_27_imag <= _zz_1101_;
      end
      if(_zz_1077_)begin
        int_reg_array_19_28_imag <= _zz_1101_;
      end
      if(_zz_1078_)begin
        int_reg_array_19_29_imag <= _zz_1101_;
      end
      if(_zz_1079_)begin
        int_reg_array_19_30_imag <= _zz_1101_;
      end
      if(_zz_1080_)begin
        int_reg_array_19_31_imag <= _zz_1101_;
      end
      if(_zz_1081_)begin
        int_reg_array_19_32_imag <= _zz_1101_;
      end
      if(_zz_1082_)begin
        int_reg_array_19_33_imag <= _zz_1101_;
      end
      if(_zz_1083_)begin
        int_reg_array_19_34_imag <= _zz_1101_;
      end
      if(_zz_1084_)begin
        int_reg_array_19_35_imag <= _zz_1101_;
      end
      if(_zz_1085_)begin
        int_reg_array_19_36_imag <= _zz_1101_;
      end
      if(_zz_1086_)begin
        int_reg_array_19_37_imag <= _zz_1101_;
      end
      if(_zz_1087_)begin
        int_reg_array_19_38_imag <= _zz_1101_;
      end
      if(_zz_1088_)begin
        int_reg_array_19_39_imag <= _zz_1101_;
      end
      if(_zz_1089_)begin
        int_reg_array_19_40_imag <= _zz_1101_;
      end
      if(_zz_1090_)begin
        int_reg_array_19_41_imag <= _zz_1101_;
      end
      if(_zz_1091_)begin
        int_reg_array_19_42_imag <= _zz_1101_;
      end
      if(_zz_1092_)begin
        int_reg_array_19_43_imag <= _zz_1101_;
      end
      if(_zz_1093_)begin
        int_reg_array_19_44_imag <= _zz_1101_;
      end
      if(_zz_1094_)begin
        int_reg_array_19_45_imag <= _zz_1101_;
      end
      if(_zz_1095_)begin
        int_reg_array_19_46_imag <= _zz_1101_;
      end
      if(_zz_1096_)begin
        int_reg_array_19_47_imag <= _zz_1101_;
      end
      if(_zz_1097_)begin
        int_reg_array_19_48_imag <= _zz_1101_;
      end
      if(_zz_1098_)begin
        int_reg_array_19_49_imag <= _zz_1101_;
      end
      if(_zz_1104_)begin
        int_reg_array_20_0_real <= _zz_1155_;
      end
      if(_zz_1105_)begin
        int_reg_array_20_1_real <= _zz_1155_;
      end
      if(_zz_1106_)begin
        int_reg_array_20_2_real <= _zz_1155_;
      end
      if(_zz_1107_)begin
        int_reg_array_20_3_real <= _zz_1155_;
      end
      if(_zz_1108_)begin
        int_reg_array_20_4_real <= _zz_1155_;
      end
      if(_zz_1109_)begin
        int_reg_array_20_5_real <= _zz_1155_;
      end
      if(_zz_1110_)begin
        int_reg_array_20_6_real <= _zz_1155_;
      end
      if(_zz_1111_)begin
        int_reg_array_20_7_real <= _zz_1155_;
      end
      if(_zz_1112_)begin
        int_reg_array_20_8_real <= _zz_1155_;
      end
      if(_zz_1113_)begin
        int_reg_array_20_9_real <= _zz_1155_;
      end
      if(_zz_1114_)begin
        int_reg_array_20_10_real <= _zz_1155_;
      end
      if(_zz_1115_)begin
        int_reg_array_20_11_real <= _zz_1155_;
      end
      if(_zz_1116_)begin
        int_reg_array_20_12_real <= _zz_1155_;
      end
      if(_zz_1117_)begin
        int_reg_array_20_13_real <= _zz_1155_;
      end
      if(_zz_1118_)begin
        int_reg_array_20_14_real <= _zz_1155_;
      end
      if(_zz_1119_)begin
        int_reg_array_20_15_real <= _zz_1155_;
      end
      if(_zz_1120_)begin
        int_reg_array_20_16_real <= _zz_1155_;
      end
      if(_zz_1121_)begin
        int_reg_array_20_17_real <= _zz_1155_;
      end
      if(_zz_1122_)begin
        int_reg_array_20_18_real <= _zz_1155_;
      end
      if(_zz_1123_)begin
        int_reg_array_20_19_real <= _zz_1155_;
      end
      if(_zz_1124_)begin
        int_reg_array_20_20_real <= _zz_1155_;
      end
      if(_zz_1125_)begin
        int_reg_array_20_21_real <= _zz_1155_;
      end
      if(_zz_1126_)begin
        int_reg_array_20_22_real <= _zz_1155_;
      end
      if(_zz_1127_)begin
        int_reg_array_20_23_real <= _zz_1155_;
      end
      if(_zz_1128_)begin
        int_reg_array_20_24_real <= _zz_1155_;
      end
      if(_zz_1129_)begin
        int_reg_array_20_25_real <= _zz_1155_;
      end
      if(_zz_1130_)begin
        int_reg_array_20_26_real <= _zz_1155_;
      end
      if(_zz_1131_)begin
        int_reg_array_20_27_real <= _zz_1155_;
      end
      if(_zz_1132_)begin
        int_reg_array_20_28_real <= _zz_1155_;
      end
      if(_zz_1133_)begin
        int_reg_array_20_29_real <= _zz_1155_;
      end
      if(_zz_1134_)begin
        int_reg_array_20_30_real <= _zz_1155_;
      end
      if(_zz_1135_)begin
        int_reg_array_20_31_real <= _zz_1155_;
      end
      if(_zz_1136_)begin
        int_reg_array_20_32_real <= _zz_1155_;
      end
      if(_zz_1137_)begin
        int_reg_array_20_33_real <= _zz_1155_;
      end
      if(_zz_1138_)begin
        int_reg_array_20_34_real <= _zz_1155_;
      end
      if(_zz_1139_)begin
        int_reg_array_20_35_real <= _zz_1155_;
      end
      if(_zz_1140_)begin
        int_reg_array_20_36_real <= _zz_1155_;
      end
      if(_zz_1141_)begin
        int_reg_array_20_37_real <= _zz_1155_;
      end
      if(_zz_1142_)begin
        int_reg_array_20_38_real <= _zz_1155_;
      end
      if(_zz_1143_)begin
        int_reg_array_20_39_real <= _zz_1155_;
      end
      if(_zz_1144_)begin
        int_reg_array_20_40_real <= _zz_1155_;
      end
      if(_zz_1145_)begin
        int_reg_array_20_41_real <= _zz_1155_;
      end
      if(_zz_1146_)begin
        int_reg_array_20_42_real <= _zz_1155_;
      end
      if(_zz_1147_)begin
        int_reg_array_20_43_real <= _zz_1155_;
      end
      if(_zz_1148_)begin
        int_reg_array_20_44_real <= _zz_1155_;
      end
      if(_zz_1149_)begin
        int_reg_array_20_45_real <= _zz_1155_;
      end
      if(_zz_1150_)begin
        int_reg_array_20_46_real <= _zz_1155_;
      end
      if(_zz_1151_)begin
        int_reg_array_20_47_real <= _zz_1155_;
      end
      if(_zz_1152_)begin
        int_reg_array_20_48_real <= _zz_1155_;
      end
      if(_zz_1153_)begin
        int_reg_array_20_49_real <= _zz_1155_;
      end
      if(_zz_1104_)begin
        int_reg_array_20_0_imag <= _zz_1156_;
      end
      if(_zz_1105_)begin
        int_reg_array_20_1_imag <= _zz_1156_;
      end
      if(_zz_1106_)begin
        int_reg_array_20_2_imag <= _zz_1156_;
      end
      if(_zz_1107_)begin
        int_reg_array_20_3_imag <= _zz_1156_;
      end
      if(_zz_1108_)begin
        int_reg_array_20_4_imag <= _zz_1156_;
      end
      if(_zz_1109_)begin
        int_reg_array_20_5_imag <= _zz_1156_;
      end
      if(_zz_1110_)begin
        int_reg_array_20_6_imag <= _zz_1156_;
      end
      if(_zz_1111_)begin
        int_reg_array_20_7_imag <= _zz_1156_;
      end
      if(_zz_1112_)begin
        int_reg_array_20_8_imag <= _zz_1156_;
      end
      if(_zz_1113_)begin
        int_reg_array_20_9_imag <= _zz_1156_;
      end
      if(_zz_1114_)begin
        int_reg_array_20_10_imag <= _zz_1156_;
      end
      if(_zz_1115_)begin
        int_reg_array_20_11_imag <= _zz_1156_;
      end
      if(_zz_1116_)begin
        int_reg_array_20_12_imag <= _zz_1156_;
      end
      if(_zz_1117_)begin
        int_reg_array_20_13_imag <= _zz_1156_;
      end
      if(_zz_1118_)begin
        int_reg_array_20_14_imag <= _zz_1156_;
      end
      if(_zz_1119_)begin
        int_reg_array_20_15_imag <= _zz_1156_;
      end
      if(_zz_1120_)begin
        int_reg_array_20_16_imag <= _zz_1156_;
      end
      if(_zz_1121_)begin
        int_reg_array_20_17_imag <= _zz_1156_;
      end
      if(_zz_1122_)begin
        int_reg_array_20_18_imag <= _zz_1156_;
      end
      if(_zz_1123_)begin
        int_reg_array_20_19_imag <= _zz_1156_;
      end
      if(_zz_1124_)begin
        int_reg_array_20_20_imag <= _zz_1156_;
      end
      if(_zz_1125_)begin
        int_reg_array_20_21_imag <= _zz_1156_;
      end
      if(_zz_1126_)begin
        int_reg_array_20_22_imag <= _zz_1156_;
      end
      if(_zz_1127_)begin
        int_reg_array_20_23_imag <= _zz_1156_;
      end
      if(_zz_1128_)begin
        int_reg_array_20_24_imag <= _zz_1156_;
      end
      if(_zz_1129_)begin
        int_reg_array_20_25_imag <= _zz_1156_;
      end
      if(_zz_1130_)begin
        int_reg_array_20_26_imag <= _zz_1156_;
      end
      if(_zz_1131_)begin
        int_reg_array_20_27_imag <= _zz_1156_;
      end
      if(_zz_1132_)begin
        int_reg_array_20_28_imag <= _zz_1156_;
      end
      if(_zz_1133_)begin
        int_reg_array_20_29_imag <= _zz_1156_;
      end
      if(_zz_1134_)begin
        int_reg_array_20_30_imag <= _zz_1156_;
      end
      if(_zz_1135_)begin
        int_reg_array_20_31_imag <= _zz_1156_;
      end
      if(_zz_1136_)begin
        int_reg_array_20_32_imag <= _zz_1156_;
      end
      if(_zz_1137_)begin
        int_reg_array_20_33_imag <= _zz_1156_;
      end
      if(_zz_1138_)begin
        int_reg_array_20_34_imag <= _zz_1156_;
      end
      if(_zz_1139_)begin
        int_reg_array_20_35_imag <= _zz_1156_;
      end
      if(_zz_1140_)begin
        int_reg_array_20_36_imag <= _zz_1156_;
      end
      if(_zz_1141_)begin
        int_reg_array_20_37_imag <= _zz_1156_;
      end
      if(_zz_1142_)begin
        int_reg_array_20_38_imag <= _zz_1156_;
      end
      if(_zz_1143_)begin
        int_reg_array_20_39_imag <= _zz_1156_;
      end
      if(_zz_1144_)begin
        int_reg_array_20_40_imag <= _zz_1156_;
      end
      if(_zz_1145_)begin
        int_reg_array_20_41_imag <= _zz_1156_;
      end
      if(_zz_1146_)begin
        int_reg_array_20_42_imag <= _zz_1156_;
      end
      if(_zz_1147_)begin
        int_reg_array_20_43_imag <= _zz_1156_;
      end
      if(_zz_1148_)begin
        int_reg_array_20_44_imag <= _zz_1156_;
      end
      if(_zz_1149_)begin
        int_reg_array_20_45_imag <= _zz_1156_;
      end
      if(_zz_1150_)begin
        int_reg_array_20_46_imag <= _zz_1156_;
      end
      if(_zz_1151_)begin
        int_reg_array_20_47_imag <= _zz_1156_;
      end
      if(_zz_1152_)begin
        int_reg_array_20_48_imag <= _zz_1156_;
      end
      if(_zz_1153_)begin
        int_reg_array_20_49_imag <= _zz_1156_;
      end
      if(_zz_1159_)begin
        int_reg_array_21_0_real <= _zz_1210_;
      end
      if(_zz_1160_)begin
        int_reg_array_21_1_real <= _zz_1210_;
      end
      if(_zz_1161_)begin
        int_reg_array_21_2_real <= _zz_1210_;
      end
      if(_zz_1162_)begin
        int_reg_array_21_3_real <= _zz_1210_;
      end
      if(_zz_1163_)begin
        int_reg_array_21_4_real <= _zz_1210_;
      end
      if(_zz_1164_)begin
        int_reg_array_21_5_real <= _zz_1210_;
      end
      if(_zz_1165_)begin
        int_reg_array_21_6_real <= _zz_1210_;
      end
      if(_zz_1166_)begin
        int_reg_array_21_7_real <= _zz_1210_;
      end
      if(_zz_1167_)begin
        int_reg_array_21_8_real <= _zz_1210_;
      end
      if(_zz_1168_)begin
        int_reg_array_21_9_real <= _zz_1210_;
      end
      if(_zz_1169_)begin
        int_reg_array_21_10_real <= _zz_1210_;
      end
      if(_zz_1170_)begin
        int_reg_array_21_11_real <= _zz_1210_;
      end
      if(_zz_1171_)begin
        int_reg_array_21_12_real <= _zz_1210_;
      end
      if(_zz_1172_)begin
        int_reg_array_21_13_real <= _zz_1210_;
      end
      if(_zz_1173_)begin
        int_reg_array_21_14_real <= _zz_1210_;
      end
      if(_zz_1174_)begin
        int_reg_array_21_15_real <= _zz_1210_;
      end
      if(_zz_1175_)begin
        int_reg_array_21_16_real <= _zz_1210_;
      end
      if(_zz_1176_)begin
        int_reg_array_21_17_real <= _zz_1210_;
      end
      if(_zz_1177_)begin
        int_reg_array_21_18_real <= _zz_1210_;
      end
      if(_zz_1178_)begin
        int_reg_array_21_19_real <= _zz_1210_;
      end
      if(_zz_1179_)begin
        int_reg_array_21_20_real <= _zz_1210_;
      end
      if(_zz_1180_)begin
        int_reg_array_21_21_real <= _zz_1210_;
      end
      if(_zz_1181_)begin
        int_reg_array_21_22_real <= _zz_1210_;
      end
      if(_zz_1182_)begin
        int_reg_array_21_23_real <= _zz_1210_;
      end
      if(_zz_1183_)begin
        int_reg_array_21_24_real <= _zz_1210_;
      end
      if(_zz_1184_)begin
        int_reg_array_21_25_real <= _zz_1210_;
      end
      if(_zz_1185_)begin
        int_reg_array_21_26_real <= _zz_1210_;
      end
      if(_zz_1186_)begin
        int_reg_array_21_27_real <= _zz_1210_;
      end
      if(_zz_1187_)begin
        int_reg_array_21_28_real <= _zz_1210_;
      end
      if(_zz_1188_)begin
        int_reg_array_21_29_real <= _zz_1210_;
      end
      if(_zz_1189_)begin
        int_reg_array_21_30_real <= _zz_1210_;
      end
      if(_zz_1190_)begin
        int_reg_array_21_31_real <= _zz_1210_;
      end
      if(_zz_1191_)begin
        int_reg_array_21_32_real <= _zz_1210_;
      end
      if(_zz_1192_)begin
        int_reg_array_21_33_real <= _zz_1210_;
      end
      if(_zz_1193_)begin
        int_reg_array_21_34_real <= _zz_1210_;
      end
      if(_zz_1194_)begin
        int_reg_array_21_35_real <= _zz_1210_;
      end
      if(_zz_1195_)begin
        int_reg_array_21_36_real <= _zz_1210_;
      end
      if(_zz_1196_)begin
        int_reg_array_21_37_real <= _zz_1210_;
      end
      if(_zz_1197_)begin
        int_reg_array_21_38_real <= _zz_1210_;
      end
      if(_zz_1198_)begin
        int_reg_array_21_39_real <= _zz_1210_;
      end
      if(_zz_1199_)begin
        int_reg_array_21_40_real <= _zz_1210_;
      end
      if(_zz_1200_)begin
        int_reg_array_21_41_real <= _zz_1210_;
      end
      if(_zz_1201_)begin
        int_reg_array_21_42_real <= _zz_1210_;
      end
      if(_zz_1202_)begin
        int_reg_array_21_43_real <= _zz_1210_;
      end
      if(_zz_1203_)begin
        int_reg_array_21_44_real <= _zz_1210_;
      end
      if(_zz_1204_)begin
        int_reg_array_21_45_real <= _zz_1210_;
      end
      if(_zz_1205_)begin
        int_reg_array_21_46_real <= _zz_1210_;
      end
      if(_zz_1206_)begin
        int_reg_array_21_47_real <= _zz_1210_;
      end
      if(_zz_1207_)begin
        int_reg_array_21_48_real <= _zz_1210_;
      end
      if(_zz_1208_)begin
        int_reg_array_21_49_real <= _zz_1210_;
      end
      if(_zz_1159_)begin
        int_reg_array_21_0_imag <= _zz_1211_;
      end
      if(_zz_1160_)begin
        int_reg_array_21_1_imag <= _zz_1211_;
      end
      if(_zz_1161_)begin
        int_reg_array_21_2_imag <= _zz_1211_;
      end
      if(_zz_1162_)begin
        int_reg_array_21_3_imag <= _zz_1211_;
      end
      if(_zz_1163_)begin
        int_reg_array_21_4_imag <= _zz_1211_;
      end
      if(_zz_1164_)begin
        int_reg_array_21_5_imag <= _zz_1211_;
      end
      if(_zz_1165_)begin
        int_reg_array_21_6_imag <= _zz_1211_;
      end
      if(_zz_1166_)begin
        int_reg_array_21_7_imag <= _zz_1211_;
      end
      if(_zz_1167_)begin
        int_reg_array_21_8_imag <= _zz_1211_;
      end
      if(_zz_1168_)begin
        int_reg_array_21_9_imag <= _zz_1211_;
      end
      if(_zz_1169_)begin
        int_reg_array_21_10_imag <= _zz_1211_;
      end
      if(_zz_1170_)begin
        int_reg_array_21_11_imag <= _zz_1211_;
      end
      if(_zz_1171_)begin
        int_reg_array_21_12_imag <= _zz_1211_;
      end
      if(_zz_1172_)begin
        int_reg_array_21_13_imag <= _zz_1211_;
      end
      if(_zz_1173_)begin
        int_reg_array_21_14_imag <= _zz_1211_;
      end
      if(_zz_1174_)begin
        int_reg_array_21_15_imag <= _zz_1211_;
      end
      if(_zz_1175_)begin
        int_reg_array_21_16_imag <= _zz_1211_;
      end
      if(_zz_1176_)begin
        int_reg_array_21_17_imag <= _zz_1211_;
      end
      if(_zz_1177_)begin
        int_reg_array_21_18_imag <= _zz_1211_;
      end
      if(_zz_1178_)begin
        int_reg_array_21_19_imag <= _zz_1211_;
      end
      if(_zz_1179_)begin
        int_reg_array_21_20_imag <= _zz_1211_;
      end
      if(_zz_1180_)begin
        int_reg_array_21_21_imag <= _zz_1211_;
      end
      if(_zz_1181_)begin
        int_reg_array_21_22_imag <= _zz_1211_;
      end
      if(_zz_1182_)begin
        int_reg_array_21_23_imag <= _zz_1211_;
      end
      if(_zz_1183_)begin
        int_reg_array_21_24_imag <= _zz_1211_;
      end
      if(_zz_1184_)begin
        int_reg_array_21_25_imag <= _zz_1211_;
      end
      if(_zz_1185_)begin
        int_reg_array_21_26_imag <= _zz_1211_;
      end
      if(_zz_1186_)begin
        int_reg_array_21_27_imag <= _zz_1211_;
      end
      if(_zz_1187_)begin
        int_reg_array_21_28_imag <= _zz_1211_;
      end
      if(_zz_1188_)begin
        int_reg_array_21_29_imag <= _zz_1211_;
      end
      if(_zz_1189_)begin
        int_reg_array_21_30_imag <= _zz_1211_;
      end
      if(_zz_1190_)begin
        int_reg_array_21_31_imag <= _zz_1211_;
      end
      if(_zz_1191_)begin
        int_reg_array_21_32_imag <= _zz_1211_;
      end
      if(_zz_1192_)begin
        int_reg_array_21_33_imag <= _zz_1211_;
      end
      if(_zz_1193_)begin
        int_reg_array_21_34_imag <= _zz_1211_;
      end
      if(_zz_1194_)begin
        int_reg_array_21_35_imag <= _zz_1211_;
      end
      if(_zz_1195_)begin
        int_reg_array_21_36_imag <= _zz_1211_;
      end
      if(_zz_1196_)begin
        int_reg_array_21_37_imag <= _zz_1211_;
      end
      if(_zz_1197_)begin
        int_reg_array_21_38_imag <= _zz_1211_;
      end
      if(_zz_1198_)begin
        int_reg_array_21_39_imag <= _zz_1211_;
      end
      if(_zz_1199_)begin
        int_reg_array_21_40_imag <= _zz_1211_;
      end
      if(_zz_1200_)begin
        int_reg_array_21_41_imag <= _zz_1211_;
      end
      if(_zz_1201_)begin
        int_reg_array_21_42_imag <= _zz_1211_;
      end
      if(_zz_1202_)begin
        int_reg_array_21_43_imag <= _zz_1211_;
      end
      if(_zz_1203_)begin
        int_reg_array_21_44_imag <= _zz_1211_;
      end
      if(_zz_1204_)begin
        int_reg_array_21_45_imag <= _zz_1211_;
      end
      if(_zz_1205_)begin
        int_reg_array_21_46_imag <= _zz_1211_;
      end
      if(_zz_1206_)begin
        int_reg_array_21_47_imag <= _zz_1211_;
      end
      if(_zz_1207_)begin
        int_reg_array_21_48_imag <= _zz_1211_;
      end
      if(_zz_1208_)begin
        int_reg_array_21_49_imag <= _zz_1211_;
      end
      if(_zz_1214_)begin
        int_reg_array_22_0_real <= _zz_1265_;
      end
      if(_zz_1215_)begin
        int_reg_array_22_1_real <= _zz_1265_;
      end
      if(_zz_1216_)begin
        int_reg_array_22_2_real <= _zz_1265_;
      end
      if(_zz_1217_)begin
        int_reg_array_22_3_real <= _zz_1265_;
      end
      if(_zz_1218_)begin
        int_reg_array_22_4_real <= _zz_1265_;
      end
      if(_zz_1219_)begin
        int_reg_array_22_5_real <= _zz_1265_;
      end
      if(_zz_1220_)begin
        int_reg_array_22_6_real <= _zz_1265_;
      end
      if(_zz_1221_)begin
        int_reg_array_22_7_real <= _zz_1265_;
      end
      if(_zz_1222_)begin
        int_reg_array_22_8_real <= _zz_1265_;
      end
      if(_zz_1223_)begin
        int_reg_array_22_9_real <= _zz_1265_;
      end
      if(_zz_1224_)begin
        int_reg_array_22_10_real <= _zz_1265_;
      end
      if(_zz_1225_)begin
        int_reg_array_22_11_real <= _zz_1265_;
      end
      if(_zz_1226_)begin
        int_reg_array_22_12_real <= _zz_1265_;
      end
      if(_zz_1227_)begin
        int_reg_array_22_13_real <= _zz_1265_;
      end
      if(_zz_1228_)begin
        int_reg_array_22_14_real <= _zz_1265_;
      end
      if(_zz_1229_)begin
        int_reg_array_22_15_real <= _zz_1265_;
      end
      if(_zz_1230_)begin
        int_reg_array_22_16_real <= _zz_1265_;
      end
      if(_zz_1231_)begin
        int_reg_array_22_17_real <= _zz_1265_;
      end
      if(_zz_1232_)begin
        int_reg_array_22_18_real <= _zz_1265_;
      end
      if(_zz_1233_)begin
        int_reg_array_22_19_real <= _zz_1265_;
      end
      if(_zz_1234_)begin
        int_reg_array_22_20_real <= _zz_1265_;
      end
      if(_zz_1235_)begin
        int_reg_array_22_21_real <= _zz_1265_;
      end
      if(_zz_1236_)begin
        int_reg_array_22_22_real <= _zz_1265_;
      end
      if(_zz_1237_)begin
        int_reg_array_22_23_real <= _zz_1265_;
      end
      if(_zz_1238_)begin
        int_reg_array_22_24_real <= _zz_1265_;
      end
      if(_zz_1239_)begin
        int_reg_array_22_25_real <= _zz_1265_;
      end
      if(_zz_1240_)begin
        int_reg_array_22_26_real <= _zz_1265_;
      end
      if(_zz_1241_)begin
        int_reg_array_22_27_real <= _zz_1265_;
      end
      if(_zz_1242_)begin
        int_reg_array_22_28_real <= _zz_1265_;
      end
      if(_zz_1243_)begin
        int_reg_array_22_29_real <= _zz_1265_;
      end
      if(_zz_1244_)begin
        int_reg_array_22_30_real <= _zz_1265_;
      end
      if(_zz_1245_)begin
        int_reg_array_22_31_real <= _zz_1265_;
      end
      if(_zz_1246_)begin
        int_reg_array_22_32_real <= _zz_1265_;
      end
      if(_zz_1247_)begin
        int_reg_array_22_33_real <= _zz_1265_;
      end
      if(_zz_1248_)begin
        int_reg_array_22_34_real <= _zz_1265_;
      end
      if(_zz_1249_)begin
        int_reg_array_22_35_real <= _zz_1265_;
      end
      if(_zz_1250_)begin
        int_reg_array_22_36_real <= _zz_1265_;
      end
      if(_zz_1251_)begin
        int_reg_array_22_37_real <= _zz_1265_;
      end
      if(_zz_1252_)begin
        int_reg_array_22_38_real <= _zz_1265_;
      end
      if(_zz_1253_)begin
        int_reg_array_22_39_real <= _zz_1265_;
      end
      if(_zz_1254_)begin
        int_reg_array_22_40_real <= _zz_1265_;
      end
      if(_zz_1255_)begin
        int_reg_array_22_41_real <= _zz_1265_;
      end
      if(_zz_1256_)begin
        int_reg_array_22_42_real <= _zz_1265_;
      end
      if(_zz_1257_)begin
        int_reg_array_22_43_real <= _zz_1265_;
      end
      if(_zz_1258_)begin
        int_reg_array_22_44_real <= _zz_1265_;
      end
      if(_zz_1259_)begin
        int_reg_array_22_45_real <= _zz_1265_;
      end
      if(_zz_1260_)begin
        int_reg_array_22_46_real <= _zz_1265_;
      end
      if(_zz_1261_)begin
        int_reg_array_22_47_real <= _zz_1265_;
      end
      if(_zz_1262_)begin
        int_reg_array_22_48_real <= _zz_1265_;
      end
      if(_zz_1263_)begin
        int_reg_array_22_49_real <= _zz_1265_;
      end
      if(_zz_1214_)begin
        int_reg_array_22_0_imag <= _zz_1266_;
      end
      if(_zz_1215_)begin
        int_reg_array_22_1_imag <= _zz_1266_;
      end
      if(_zz_1216_)begin
        int_reg_array_22_2_imag <= _zz_1266_;
      end
      if(_zz_1217_)begin
        int_reg_array_22_3_imag <= _zz_1266_;
      end
      if(_zz_1218_)begin
        int_reg_array_22_4_imag <= _zz_1266_;
      end
      if(_zz_1219_)begin
        int_reg_array_22_5_imag <= _zz_1266_;
      end
      if(_zz_1220_)begin
        int_reg_array_22_6_imag <= _zz_1266_;
      end
      if(_zz_1221_)begin
        int_reg_array_22_7_imag <= _zz_1266_;
      end
      if(_zz_1222_)begin
        int_reg_array_22_8_imag <= _zz_1266_;
      end
      if(_zz_1223_)begin
        int_reg_array_22_9_imag <= _zz_1266_;
      end
      if(_zz_1224_)begin
        int_reg_array_22_10_imag <= _zz_1266_;
      end
      if(_zz_1225_)begin
        int_reg_array_22_11_imag <= _zz_1266_;
      end
      if(_zz_1226_)begin
        int_reg_array_22_12_imag <= _zz_1266_;
      end
      if(_zz_1227_)begin
        int_reg_array_22_13_imag <= _zz_1266_;
      end
      if(_zz_1228_)begin
        int_reg_array_22_14_imag <= _zz_1266_;
      end
      if(_zz_1229_)begin
        int_reg_array_22_15_imag <= _zz_1266_;
      end
      if(_zz_1230_)begin
        int_reg_array_22_16_imag <= _zz_1266_;
      end
      if(_zz_1231_)begin
        int_reg_array_22_17_imag <= _zz_1266_;
      end
      if(_zz_1232_)begin
        int_reg_array_22_18_imag <= _zz_1266_;
      end
      if(_zz_1233_)begin
        int_reg_array_22_19_imag <= _zz_1266_;
      end
      if(_zz_1234_)begin
        int_reg_array_22_20_imag <= _zz_1266_;
      end
      if(_zz_1235_)begin
        int_reg_array_22_21_imag <= _zz_1266_;
      end
      if(_zz_1236_)begin
        int_reg_array_22_22_imag <= _zz_1266_;
      end
      if(_zz_1237_)begin
        int_reg_array_22_23_imag <= _zz_1266_;
      end
      if(_zz_1238_)begin
        int_reg_array_22_24_imag <= _zz_1266_;
      end
      if(_zz_1239_)begin
        int_reg_array_22_25_imag <= _zz_1266_;
      end
      if(_zz_1240_)begin
        int_reg_array_22_26_imag <= _zz_1266_;
      end
      if(_zz_1241_)begin
        int_reg_array_22_27_imag <= _zz_1266_;
      end
      if(_zz_1242_)begin
        int_reg_array_22_28_imag <= _zz_1266_;
      end
      if(_zz_1243_)begin
        int_reg_array_22_29_imag <= _zz_1266_;
      end
      if(_zz_1244_)begin
        int_reg_array_22_30_imag <= _zz_1266_;
      end
      if(_zz_1245_)begin
        int_reg_array_22_31_imag <= _zz_1266_;
      end
      if(_zz_1246_)begin
        int_reg_array_22_32_imag <= _zz_1266_;
      end
      if(_zz_1247_)begin
        int_reg_array_22_33_imag <= _zz_1266_;
      end
      if(_zz_1248_)begin
        int_reg_array_22_34_imag <= _zz_1266_;
      end
      if(_zz_1249_)begin
        int_reg_array_22_35_imag <= _zz_1266_;
      end
      if(_zz_1250_)begin
        int_reg_array_22_36_imag <= _zz_1266_;
      end
      if(_zz_1251_)begin
        int_reg_array_22_37_imag <= _zz_1266_;
      end
      if(_zz_1252_)begin
        int_reg_array_22_38_imag <= _zz_1266_;
      end
      if(_zz_1253_)begin
        int_reg_array_22_39_imag <= _zz_1266_;
      end
      if(_zz_1254_)begin
        int_reg_array_22_40_imag <= _zz_1266_;
      end
      if(_zz_1255_)begin
        int_reg_array_22_41_imag <= _zz_1266_;
      end
      if(_zz_1256_)begin
        int_reg_array_22_42_imag <= _zz_1266_;
      end
      if(_zz_1257_)begin
        int_reg_array_22_43_imag <= _zz_1266_;
      end
      if(_zz_1258_)begin
        int_reg_array_22_44_imag <= _zz_1266_;
      end
      if(_zz_1259_)begin
        int_reg_array_22_45_imag <= _zz_1266_;
      end
      if(_zz_1260_)begin
        int_reg_array_22_46_imag <= _zz_1266_;
      end
      if(_zz_1261_)begin
        int_reg_array_22_47_imag <= _zz_1266_;
      end
      if(_zz_1262_)begin
        int_reg_array_22_48_imag <= _zz_1266_;
      end
      if(_zz_1263_)begin
        int_reg_array_22_49_imag <= _zz_1266_;
      end
      if(_zz_1269_)begin
        int_reg_array_23_0_real <= _zz_1320_;
      end
      if(_zz_1270_)begin
        int_reg_array_23_1_real <= _zz_1320_;
      end
      if(_zz_1271_)begin
        int_reg_array_23_2_real <= _zz_1320_;
      end
      if(_zz_1272_)begin
        int_reg_array_23_3_real <= _zz_1320_;
      end
      if(_zz_1273_)begin
        int_reg_array_23_4_real <= _zz_1320_;
      end
      if(_zz_1274_)begin
        int_reg_array_23_5_real <= _zz_1320_;
      end
      if(_zz_1275_)begin
        int_reg_array_23_6_real <= _zz_1320_;
      end
      if(_zz_1276_)begin
        int_reg_array_23_7_real <= _zz_1320_;
      end
      if(_zz_1277_)begin
        int_reg_array_23_8_real <= _zz_1320_;
      end
      if(_zz_1278_)begin
        int_reg_array_23_9_real <= _zz_1320_;
      end
      if(_zz_1279_)begin
        int_reg_array_23_10_real <= _zz_1320_;
      end
      if(_zz_1280_)begin
        int_reg_array_23_11_real <= _zz_1320_;
      end
      if(_zz_1281_)begin
        int_reg_array_23_12_real <= _zz_1320_;
      end
      if(_zz_1282_)begin
        int_reg_array_23_13_real <= _zz_1320_;
      end
      if(_zz_1283_)begin
        int_reg_array_23_14_real <= _zz_1320_;
      end
      if(_zz_1284_)begin
        int_reg_array_23_15_real <= _zz_1320_;
      end
      if(_zz_1285_)begin
        int_reg_array_23_16_real <= _zz_1320_;
      end
      if(_zz_1286_)begin
        int_reg_array_23_17_real <= _zz_1320_;
      end
      if(_zz_1287_)begin
        int_reg_array_23_18_real <= _zz_1320_;
      end
      if(_zz_1288_)begin
        int_reg_array_23_19_real <= _zz_1320_;
      end
      if(_zz_1289_)begin
        int_reg_array_23_20_real <= _zz_1320_;
      end
      if(_zz_1290_)begin
        int_reg_array_23_21_real <= _zz_1320_;
      end
      if(_zz_1291_)begin
        int_reg_array_23_22_real <= _zz_1320_;
      end
      if(_zz_1292_)begin
        int_reg_array_23_23_real <= _zz_1320_;
      end
      if(_zz_1293_)begin
        int_reg_array_23_24_real <= _zz_1320_;
      end
      if(_zz_1294_)begin
        int_reg_array_23_25_real <= _zz_1320_;
      end
      if(_zz_1295_)begin
        int_reg_array_23_26_real <= _zz_1320_;
      end
      if(_zz_1296_)begin
        int_reg_array_23_27_real <= _zz_1320_;
      end
      if(_zz_1297_)begin
        int_reg_array_23_28_real <= _zz_1320_;
      end
      if(_zz_1298_)begin
        int_reg_array_23_29_real <= _zz_1320_;
      end
      if(_zz_1299_)begin
        int_reg_array_23_30_real <= _zz_1320_;
      end
      if(_zz_1300_)begin
        int_reg_array_23_31_real <= _zz_1320_;
      end
      if(_zz_1301_)begin
        int_reg_array_23_32_real <= _zz_1320_;
      end
      if(_zz_1302_)begin
        int_reg_array_23_33_real <= _zz_1320_;
      end
      if(_zz_1303_)begin
        int_reg_array_23_34_real <= _zz_1320_;
      end
      if(_zz_1304_)begin
        int_reg_array_23_35_real <= _zz_1320_;
      end
      if(_zz_1305_)begin
        int_reg_array_23_36_real <= _zz_1320_;
      end
      if(_zz_1306_)begin
        int_reg_array_23_37_real <= _zz_1320_;
      end
      if(_zz_1307_)begin
        int_reg_array_23_38_real <= _zz_1320_;
      end
      if(_zz_1308_)begin
        int_reg_array_23_39_real <= _zz_1320_;
      end
      if(_zz_1309_)begin
        int_reg_array_23_40_real <= _zz_1320_;
      end
      if(_zz_1310_)begin
        int_reg_array_23_41_real <= _zz_1320_;
      end
      if(_zz_1311_)begin
        int_reg_array_23_42_real <= _zz_1320_;
      end
      if(_zz_1312_)begin
        int_reg_array_23_43_real <= _zz_1320_;
      end
      if(_zz_1313_)begin
        int_reg_array_23_44_real <= _zz_1320_;
      end
      if(_zz_1314_)begin
        int_reg_array_23_45_real <= _zz_1320_;
      end
      if(_zz_1315_)begin
        int_reg_array_23_46_real <= _zz_1320_;
      end
      if(_zz_1316_)begin
        int_reg_array_23_47_real <= _zz_1320_;
      end
      if(_zz_1317_)begin
        int_reg_array_23_48_real <= _zz_1320_;
      end
      if(_zz_1318_)begin
        int_reg_array_23_49_real <= _zz_1320_;
      end
      if(_zz_1269_)begin
        int_reg_array_23_0_imag <= _zz_1321_;
      end
      if(_zz_1270_)begin
        int_reg_array_23_1_imag <= _zz_1321_;
      end
      if(_zz_1271_)begin
        int_reg_array_23_2_imag <= _zz_1321_;
      end
      if(_zz_1272_)begin
        int_reg_array_23_3_imag <= _zz_1321_;
      end
      if(_zz_1273_)begin
        int_reg_array_23_4_imag <= _zz_1321_;
      end
      if(_zz_1274_)begin
        int_reg_array_23_5_imag <= _zz_1321_;
      end
      if(_zz_1275_)begin
        int_reg_array_23_6_imag <= _zz_1321_;
      end
      if(_zz_1276_)begin
        int_reg_array_23_7_imag <= _zz_1321_;
      end
      if(_zz_1277_)begin
        int_reg_array_23_8_imag <= _zz_1321_;
      end
      if(_zz_1278_)begin
        int_reg_array_23_9_imag <= _zz_1321_;
      end
      if(_zz_1279_)begin
        int_reg_array_23_10_imag <= _zz_1321_;
      end
      if(_zz_1280_)begin
        int_reg_array_23_11_imag <= _zz_1321_;
      end
      if(_zz_1281_)begin
        int_reg_array_23_12_imag <= _zz_1321_;
      end
      if(_zz_1282_)begin
        int_reg_array_23_13_imag <= _zz_1321_;
      end
      if(_zz_1283_)begin
        int_reg_array_23_14_imag <= _zz_1321_;
      end
      if(_zz_1284_)begin
        int_reg_array_23_15_imag <= _zz_1321_;
      end
      if(_zz_1285_)begin
        int_reg_array_23_16_imag <= _zz_1321_;
      end
      if(_zz_1286_)begin
        int_reg_array_23_17_imag <= _zz_1321_;
      end
      if(_zz_1287_)begin
        int_reg_array_23_18_imag <= _zz_1321_;
      end
      if(_zz_1288_)begin
        int_reg_array_23_19_imag <= _zz_1321_;
      end
      if(_zz_1289_)begin
        int_reg_array_23_20_imag <= _zz_1321_;
      end
      if(_zz_1290_)begin
        int_reg_array_23_21_imag <= _zz_1321_;
      end
      if(_zz_1291_)begin
        int_reg_array_23_22_imag <= _zz_1321_;
      end
      if(_zz_1292_)begin
        int_reg_array_23_23_imag <= _zz_1321_;
      end
      if(_zz_1293_)begin
        int_reg_array_23_24_imag <= _zz_1321_;
      end
      if(_zz_1294_)begin
        int_reg_array_23_25_imag <= _zz_1321_;
      end
      if(_zz_1295_)begin
        int_reg_array_23_26_imag <= _zz_1321_;
      end
      if(_zz_1296_)begin
        int_reg_array_23_27_imag <= _zz_1321_;
      end
      if(_zz_1297_)begin
        int_reg_array_23_28_imag <= _zz_1321_;
      end
      if(_zz_1298_)begin
        int_reg_array_23_29_imag <= _zz_1321_;
      end
      if(_zz_1299_)begin
        int_reg_array_23_30_imag <= _zz_1321_;
      end
      if(_zz_1300_)begin
        int_reg_array_23_31_imag <= _zz_1321_;
      end
      if(_zz_1301_)begin
        int_reg_array_23_32_imag <= _zz_1321_;
      end
      if(_zz_1302_)begin
        int_reg_array_23_33_imag <= _zz_1321_;
      end
      if(_zz_1303_)begin
        int_reg_array_23_34_imag <= _zz_1321_;
      end
      if(_zz_1304_)begin
        int_reg_array_23_35_imag <= _zz_1321_;
      end
      if(_zz_1305_)begin
        int_reg_array_23_36_imag <= _zz_1321_;
      end
      if(_zz_1306_)begin
        int_reg_array_23_37_imag <= _zz_1321_;
      end
      if(_zz_1307_)begin
        int_reg_array_23_38_imag <= _zz_1321_;
      end
      if(_zz_1308_)begin
        int_reg_array_23_39_imag <= _zz_1321_;
      end
      if(_zz_1309_)begin
        int_reg_array_23_40_imag <= _zz_1321_;
      end
      if(_zz_1310_)begin
        int_reg_array_23_41_imag <= _zz_1321_;
      end
      if(_zz_1311_)begin
        int_reg_array_23_42_imag <= _zz_1321_;
      end
      if(_zz_1312_)begin
        int_reg_array_23_43_imag <= _zz_1321_;
      end
      if(_zz_1313_)begin
        int_reg_array_23_44_imag <= _zz_1321_;
      end
      if(_zz_1314_)begin
        int_reg_array_23_45_imag <= _zz_1321_;
      end
      if(_zz_1315_)begin
        int_reg_array_23_46_imag <= _zz_1321_;
      end
      if(_zz_1316_)begin
        int_reg_array_23_47_imag <= _zz_1321_;
      end
      if(_zz_1317_)begin
        int_reg_array_23_48_imag <= _zz_1321_;
      end
      if(_zz_1318_)begin
        int_reg_array_23_49_imag <= _zz_1321_;
      end
      if(_zz_1324_)begin
        int_reg_array_24_0_real <= _zz_1375_;
      end
      if(_zz_1325_)begin
        int_reg_array_24_1_real <= _zz_1375_;
      end
      if(_zz_1326_)begin
        int_reg_array_24_2_real <= _zz_1375_;
      end
      if(_zz_1327_)begin
        int_reg_array_24_3_real <= _zz_1375_;
      end
      if(_zz_1328_)begin
        int_reg_array_24_4_real <= _zz_1375_;
      end
      if(_zz_1329_)begin
        int_reg_array_24_5_real <= _zz_1375_;
      end
      if(_zz_1330_)begin
        int_reg_array_24_6_real <= _zz_1375_;
      end
      if(_zz_1331_)begin
        int_reg_array_24_7_real <= _zz_1375_;
      end
      if(_zz_1332_)begin
        int_reg_array_24_8_real <= _zz_1375_;
      end
      if(_zz_1333_)begin
        int_reg_array_24_9_real <= _zz_1375_;
      end
      if(_zz_1334_)begin
        int_reg_array_24_10_real <= _zz_1375_;
      end
      if(_zz_1335_)begin
        int_reg_array_24_11_real <= _zz_1375_;
      end
      if(_zz_1336_)begin
        int_reg_array_24_12_real <= _zz_1375_;
      end
      if(_zz_1337_)begin
        int_reg_array_24_13_real <= _zz_1375_;
      end
      if(_zz_1338_)begin
        int_reg_array_24_14_real <= _zz_1375_;
      end
      if(_zz_1339_)begin
        int_reg_array_24_15_real <= _zz_1375_;
      end
      if(_zz_1340_)begin
        int_reg_array_24_16_real <= _zz_1375_;
      end
      if(_zz_1341_)begin
        int_reg_array_24_17_real <= _zz_1375_;
      end
      if(_zz_1342_)begin
        int_reg_array_24_18_real <= _zz_1375_;
      end
      if(_zz_1343_)begin
        int_reg_array_24_19_real <= _zz_1375_;
      end
      if(_zz_1344_)begin
        int_reg_array_24_20_real <= _zz_1375_;
      end
      if(_zz_1345_)begin
        int_reg_array_24_21_real <= _zz_1375_;
      end
      if(_zz_1346_)begin
        int_reg_array_24_22_real <= _zz_1375_;
      end
      if(_zz_1347_)begin
        int_reg_array_24_23_real <= _zz_1375_;
      end
      if(_zz_1348_)begin
        int_reg_array_24_24_real <= _zz_1375_;
      end
      if(_zz_1349_)begin
        int_reg_array_24_25_real <= _zz_1375_;
      end
      if(_zz_1350_)begin
        int_reg_array_24_26_real <= _zz_1375_;
      end
      if(_zz_1351_)begin
        int_reg_array_24_27_real <= _zz_1375_;
      end
      if(_zz_1352_)begin
        int_reg_array_24_28_real <= _zz_1375_;
      end
      if(_zz_1353_)begin
        int_reg_array_24_29_real <= _zz_1375_;
      end
      if(_zz_1354_)begin
        int_reg_array_24_30_real <= _zz_1375_;
      end
      if(_zz_1355_)begin
        int_reg_array_24_31_real <= _zz_1375_;
      end
      if(_zz_1356_)begin
        int_reg_array_24_32_real <= _zz_1375_;
      end
      if(_zz_1357_)begin
        int_reg_array_24_33_real <= _zz_1375_;
      end
      if(_zz_1358_)begin
        int_reg_array_24_34_real <= _zz_1375_;
      end
      if(_zz_1359_)begin
        int_reg_array_24_35_real <= _zz_1375_;
      end
      if(_zz_1360_)begin
        int_reg_array_24_36_real <= _zz_1375_;
      end
      if(_zz_1361_)begin
        int_reg_array_24_37_real <= _zz_1375_;
      end
      if(_zz_1362_)begin
        int_reg_array_24_38_real <= _zz_1375_;
      end
      if(_zz_1363_)begin
        int_reg_array_24_39_real <= _zz_1375_;
      end
      if(_zz_1364_)begin
        int_reg_array_24_40_real <= _zz_1375_;
      end
      if(_zz_1365_)begin
        int_reg_array_24_41_real <= _zz_1375_;
      end
      if(_zz_1366_)begin
        int_reg_array_24_42_real <= _zz_1375_;
      end
      if(_zz_1367_)begin
        int_reg_array_24_43_real <= _zz_1375_;
      end
      if(_zz_1368_)begin
        int_reg_array_24_44_real <= _zz_1375_;
      end
      if(_zz_1369_)begin
        int_reg_array_24_45_real <= _zz_1375_;
      end
      if(_zz_1370_)begin
        int_reg_array_24_46_real <= _zz_1375_;
      end
      if(_zz_1371_)begin
        int_reg_array_24_47_real <= _zz_1375_;
      end
      if(_zz_1372_)begin
        int_reg_array_24_48_real <= _zz_1375_;
      end
      if(_zz_1373_)begin
        int_reg_array_24_49_real <= _zz_1375_;
      end
      if(_zz_1324_)begin
        int_reg_array_24_0_imag <= _zz_1376_;
      end
      if(_zz_1325_)begin
        int_reg_array_24_1_imag <= _zz_1376_;
      end
      if(_zz_1326_)begin
        int_reg_array_24_2_imag <= _zz_1376_;
      end
      if(_zz_1327_)begin
        int_reg_array_24_3_imag <= _zz_1376_;
      end
      if(_zz_1328_)begin
        int_reg_array_24_4_imag <= _zz_1376_;
      end
      if(_zz_1329_)begin
        int_reg_array_24_5_imag <= _zz_1376_;
      end
      if(_zz_1330_)begin
        int_reg_array_24_6_imag <= _zz_1376_;
      end
      if(_zz_1331_)begin
        int_reg_array_24_7_imag <= _zz_1376_;
      end
      if(_zz_1332_)begin
        int_reg_array_24_8_imag <= _zz_1376_;
      end
      if(_zz_1333_)begin
        int_reg_array_24_9_imag <= _zz_1376_;
      end
      if(_zz_1334_)begin
        int_reg_array_24_10_imag <= _zz_1376_;
      end
      if(_zz_1335_)begin
        int_reg_array_24_11_imag <= _zz_1376_;
      end
      if(_zz_1336_)begin
        int_reg_array_24_12_imag <= _zz_1376_;
      end
      if(_zz_1337_)begin
        int_reg_array_24_13_imag <= _zz_1376_;
      end
      if(_zz_1338_)begin
        int_reg_array_24_14_imag <= _zz_1376_;
      end
      if(_zz_1339_)begin
        int_reg_array_24_15_imag <= _zz_1376_;
      end
      if(_zz_1340_)begin
        int_reg_array_24_16_imag <= _zz_1376_;
      end
      if(_zz_1341_)begin
        int_reg_array_24_17_imag <= _zz_1376_;
      end
      if(_zz_1342_)begin
        int_reg_array_24_18_imag <= _zz_1376_;
      end
      if(_zz_1343_)begin
        int_reg_array_24_19_imag <= _zz_1376_;
      end
      if(_zz_1344_)begin
        int_reg_array_24_20_imag <= _zz_1376_;
      end
      if(_zz_1345_)begin
        int_reg_array_24_21_imag <= _zz_1376_;
      end
      if(_zz_1346_)begin
        int_reg_array_24_22_imag <= _zz_1376_;
      end
      if(_zz_1347_)begin
        int_reg_array_24_23_imag <= _zz_1376_;
      end
      if(_zz_1348_)begin
        int_reg_array_24_24_imag <= _zz_1376_;
      end
      if(_zz_1349_)begin
        int_reg_array_24_25_imag <= _zz_1376_;
      end
      if(_zz_1350_)begin
        int_reg_array_24_26_imag <= _zz_1376_;
      end
      if(_zz_1351_)begin
        int_reg_array_24_27_imag <= _zz_1376_;
      end
      if(_zz_1352_)begin
        int_reg_array_24_28_imag <= _zz_1376_;
      end
      if(_zz_1353_)begin
        int_reg_array_24_29_imag <= _zz_1376_;
      end
      if(_zz_1354_)begin
        int_reg_array_24_30_imag <= _zz_1376_;
      end
      if(_zz_1355_)begin
        int_reg_array_24_31_imag <= _zz_1376_;
      end
      if(_zz_1356_)begin
        int_reg_array_24_32_imag <= _zz_1376_;
      end
      if(_zz_1357_)begin
        int_reg_array_24_33_imag <= _zz_1376_;
      end
      if(_zz_1358_)begin
        int_reg_array_24_34_imag <= _zz_1376_;
      end
      if(_zz_1359_)begin
        int_reg_array_24_35_imag <= _zz_1376_;
      end
      if(_zz_1360_)begin
        int_reg_array_24_36_imag <= _zz_1376_;
      end
      if(_zz_1361_)begin
        int_reg_array_24_37_imag <= _zz_1376_;
      end
      if(_zz_1362_)begin
        int_reg_array_24_38_imag <= _zz_1376_;
      end
      if(_zz_1363_)begin
        int_reg_array_24_39_imag <= _zz_1376_;
      end
      if(_zz_1364_)begin
        int_reg_array_24_40_imag <= _zz_1376_;
      end
      if(_zz_1365_)begin
        int_reg_array_24_41_imag <= _zz_1376_;
      end
      if(_zz_1366_)begin
        int_reg_array_24_42_imag <= _zz_1376_;
      end
      if(_zz_1367_)begin
        int_reg_array_24_43_imag <= _zz_1376_;
      end
      if(_zz_1368_)begin
        int_reg_array_24_44_imag <= _zz_1376_;
      end
      if(_zz_1369_)begin
        int_reg_array_24_45_imag <= _zz_1376_;
      end
      if(_zz_1370_)begin
        int_reg_array_24_46_imag <= _zz_1376_;
      end
      if(_zz_1371_)begin
        int_reg_array_24_47_imag <= _zz_1376_;
      end
      if(_zz_1372_)begin
        int_reg_array_24_48_imag <= _zz_1376_;
      end
      if(_zz_1373_)begin
        int_reg_array_24_49_imag <= _zz_1376_;
      end
      if(_zz_1379_)begin
        int_reg_array_25_0_real <= _zz_1430_;
      end
      if(_zz_1380_)begin
        int_reg_array_25_1_real <= _zz_1430_;
      end
      if(_zz_1381_)begin
        int_reg_array_25_2_real <= _zz_1430_;
      end
      if(_zz_1382_)begin
        int_reg_array_25_3_real <= _zz_1430_;
      end
      if(_zz_1383_)begin
        int_reg_array_25_4_real <= _zz_1430_;
      end
      if(_zz_1384_)begin
        int_reg_array_25_5_real <= _zz_1430_;
      end
      if(_zz_1385_)begin
        int_reg_array_25_6_real <= _zz_1430_;
      end
      if(_zz_1386_)begin
        int_reg_array_25_7_real <= _zz_1430_;
      end
      if(_zz_1387_)begin
        int_reg_array_25_8_real <= _zz_1430_;
      end
      if(_zz_1388_)begin
        int_reg_array_25_9_real <= _zz_1430_;
      end
      if(_zz_1389_)begin
        int_reg_array_25_10_real <= _zz_1430_;
      end
      if(_zz_1390_)begin
        int_reg_array_25_11_real <= _zz_1430_;
      end
      if(_zz_1391_)begin
        int_reg_array_25_12_real <= _zz_1430_;
      end
      if(_zz_1392_)begin
        int_reg_array_25_13_real <= _zz_1430_;
      end
      if(_zz_1393_)begin
        int_reg_array_25_14_real <= _zz_1430_;
      end
      if(_zz_1394_)begin
        int_reg_array_25_15_real <= _zz_1430_;
      end
      if(_zz_1395_)begin
        int_reg_array_25_16_real <= _zz_1430_;
      end
      if(_zz_1396_)begin
        int_reg_array_25_17_real <= _zz_1430_;
      end
      if(_zz_1397_)begin
        int_reg_array_25_18_real <= _zz_1430_;
      end
      if(_zz_1398_)begin
        int_reg_array_25_19_real <= _zz_1430_;
      end
      if(_zz_1399_)begin
        int_reg_array_25_20_real <= _zz_1430_;
      end
      if(_zz_1400_)begin
        int_reg_array_25_21_real <= _zz_1430_;
      end
      if(_zz_1401_)begin
        int_reg_array_25_22_real <= _zz_1430_;
      end
      if(_zz_1402_)begin
        int_reg_array_25_23_real <= _zz_1430_;
      end
      if(_zz_1403_)begin
        int_reg_array_25_24_real <= _zz_1430_;
      end
      if(_zz_1404_)begin
        int_reg_array_25_25_real <= _zz_1430_;
      end
      if(_zz_1405_)begin
        int_reg_array_25_26_real <= _zz_1430_;
      end
      if(_zz_1406_)begin
        int_reg_array_25_27_real <= _zz_1430_;
      end
      if(_zz_1407_)begin
        int_reg_array_25_28_real <= _zz_1430_;
      end
      if(_zz_1408_)begin
        int_reg_array_25_29_real <= _zz_1430_;
      end
      if(_zz_1409_)begin
        int_reg_array_25_30_real <= _zz_1430_;
      end
      if(_zz_1410_)begin
        int_reg_array_25_31_real <= _zz_1430_;
      end
      if(_zz_1411_)begin
        int_reg_array_25_32_real <= _zz_1430_;
      end
      if(_zz_1412_)begin
        int_reg_array_25_33_real <= _zz_1430_;
      end
      if(_zz_1413_)begin
        int_reg_array_25_34_real <= _zz_1430_;
      end
      if(_zz_1414_)begin
        int_reg_array_25_35_real <= _zz_1430_;
      end
      if(_zz_1415_)begin
        int_reg_array_25_36_real <= _zz_1430_;
      end
      if(_zz_1416_)begin
        int_reg_array_25_37_real <= _zz_1430_;
      end
      if(_zz_1417_)begin
        int_reg_array_25_38_real <= _zz_1430_;
      end
      if(_zz_1418_)begin
        int_reg_array_25_39_real <= _zz_1430_;
      end
      if(_zz_1419_)begin
        int_reg_array_25_40_real <= _zz_1430_;
      end
      if(_zz_1420_)begin
        int_reg_array_25_41_real <= _zz_1430_;
      end
      if(_zz_1421_)begin
        int_reg_array_25_42_real <= _zz_1430_;
      end
      if(_zz_1422_)begin
        int_reg_array_25_43_real <= _zz_1430_;
      end
      if(_zz_1423_)begin
        int_reg_array_25_44_real <= _zz_1430_;
      end
      if(_zz_1424_)begin
        int_reg_array_25_45_real <= _zz_1430_;
      end
      if(_zz_1425_)begin
        int_reg_array_25_46_real <= _zz_1430_;
      end
      if(_zz_1426_)begin
        int_reg_array_25_47_real <= _zz_1430_;
      end
      if(_zz_1427_)begin
        int_reg_array_25_48_real <= _zz_1430_;
      end
      if(_zz_1428_)begin
        int_reg_array_25_49_real <= _zz_1430_;
      end
      if(_zz_1379_)begin
        int_reg_array_25_0_imag <= _zz_1431_;
      end
      if(_zz_1380_)begin
        int_reg_array_25_1_imag <= _zz_1431_;
      end
      if(_zz_1381_)begin
        int_reg_array_25_2_imag <= _zz_1431_;
      end
      if(_zz_1382_)begin
        int_reg_array_25_3_imag <= _zz_1431_;
      end
      if(_zz_1383_)begin
        int_reg_array_25_4_imag <= _zz_1431_;
      end
      if(_zz_1384_)begin
        int_reg_array_25_5_imag <= _zz_1431_;
      end
      if(_zz_1385_)begin
        int_reg_array_25_6_imag <= _zz_1431_;
      end
      if(_zz_1386_)begin
        int_reg_array_25_7_imag <= _zz_1431_;
      end
      if(_zz_1387_)begin
        int_reg_array_25_8_imag <= _zz_1431_;
      end
      if(_zz_1388_)begin
        int_reg_array_25_9_imag <= _zz_1431_;
      end
      if(_zz_1389_)begin
        int_reg_array_25_10_imag <= _zz_1431_;
      end
      if(_zz_1390_)begin
        int_reg_array_25_11_imag <= _zz_1431_;
      end
      if(_zz_1391_)begin
        int_reg_array_25_12_imag <= _zz_1431_;
      end
      if(_zz_1392_)begin
        int_reg_array_25_13_imag <= _zz_1431_;
      end
      if(_zz_1393_)begin
        int_reg_array_25_14_imag <= _zz_1431_;
      end
      if(_zz_1394_)begin
        int_reg_array_25_15_imag <= _zz_1431_;
      end
      if(_zz_1395_)begin
        int_reg_array_25_16_imag <= _zz_1431_;
      end
      if(_zz_1396_)begin
        int_reg_array_25_17_imag <= _zz_1431_;
      end
      if(_zz_1397_)begin
        int_reg_array_25_18_imag <= _zz_1431_;
      end
      if(_zz_1398_)begin
        int_reg_array_25_19_imag <= _zz_1431_;
      end
      if(_zz_1399_)begin
        int_reg_array_25_20_imag <= _zz_1431_;
      end
      if(_zz_1400_)begin
        int_reg_array_25_21_imag <= _zz_1431_;
      end
      if(_zz_1401_)begin
        int_reg_array_25_22_imag <= _zz_1431_;
      end
      if(_zz_1402_)begin
        int_reg_array_25_23_imag <= _zz_1431_;
      end
      if(_zz_1403_)begin
        int_reg_array_25_24_imag <= _zz_1431_;
      end
      if(_zz_1404_)begin
        int_reg_array_25_25_imag <= _zz_1431_;
      end
      if(_zz_1405_)begin
        int_reg_array_25_26_imag <= _zz_1431_;
      end
      if(_zz_1406_)begin
        int_reg_array_25_27_imag <= _zz_1431_;
      end
      if(_zz_1407_)begin
        int_reg_array_25_28_imag <= _zz_1431_;
      end
      if(_zz_1408_)begin
        int_reg_array_25_29_imag <= _zz_1431_;
      end
      if(_zz_1409_)begin
        int_reg_array_25_30_imag <= _zz_1431_;
      end
      if(_zz_1410_)begin
        int_reg_array_25_31_imag <= _zz_1431_;
      end
      if(_zz_1411_)begin
        int_reg_array_25_32_imag <= _zz_1431_;
      end
      if(_zz_1412_)begin
        int_reg_array_25_33_imag <= _zz_1431_;
      end
      if(_zz_1413_)begin
        int_reg_array_25_34_imag <= _zz_1431_;
      end
      if(_zz_1414_)begin
        int_reg_array_25_35_imag <= _zz_1431_;
      end
      if(_zz_1415_)begin
        int_reg_array_25_36_imag <= _zz_1431_;
      end
      if(_zz_1416_)begin
        int_reg_array_25_37_imag <= _zz_1431_;
      end
      if(_zz_1417_)begin
        int_reg_array_25_38_imag <= _zz_1431_;
      end
      if(_zz_1418_)begin
        int_reg_array_25_39_imag <= _zz_1431_;
      end
      if(_zz_1419_)begin
        int_reg_array_25_40_imag <= _zz_1431_;
      end
      if(_zz_1420_)begin
        int_reg_array_25_41_imag <= _zz_1431_;
      end
      if(_zz_1421_)begin
        int_reg_array_25_42_imag <= _zz_1431_;
      end
      if(_zz_1422_)begin
        int_reg_array_25_43_imag <= _zz_1431_;
      end
      if(_zz_1423_)begin
        int_reg_array_25_44_imag <= _zz_1431_;
      end
      if(_zz_1424_)begin
        int_reg_array_25_45_imag <= _zz_1431_;
      end
      if(_zz_1425_)begin
        int_reg_array_25_46_imag <= _zz_1431_;
      end
      if(_zz_1426_)begin
        int_reg_array_25_47_imag <= _zz_1431_;
      end
      if(_zz_1427_)begin
        int_reg_array_25_48_imag <= _zz_1431_;
      end
      if(_zz_1428_)begin
        int_reg_array_25_49_imag <= _zz_1431_;
      end
      if(_zz_1434_)begin
        int_reg_array_26_0_real <= _zz_1485_;
      end
      if(_zz_1435_)begin
        int_reg_array_26_1_real <= _zz_1485_;
      end
      if(_zz_1436_)begin
        int_reg_array_26_2_real <= _zz_1485_;
      end
      if(_zz_1437_)begin
        int_reg_array_26_3_real <= _zz_1485_;
      end
      if(_zz_1438_)begin
        int_reg_array_26_4_real <= _zz_1485_;
      end
      if(_zz_1439_)begin
        int_reg_array_26_5_real <= _zz_1485_;
      end
      if(_zz_1440_)begin
        int_reg_array_26_6_real <= _zz_1485_;
      end
      if(_zz_1441_)begin
        int_reg_array_26_7_real <= _zz_1485_;
      end
      if(_zz_1442_)begin
        int_reg_array_26_8_real <= _zz_1485_;
      end
      if(_zz_1443_)begin
        int_reg_array_26_9_real <= _zz_1485_;
      end
      if(_zz_1444_)begin
        int_reg_array_26_10_real <= _zz_1485_;
      end
      if(_zz_1445_)begin
        int_reg_array_26_11_real <= _zz_1485_;
      end
      if(_zz_1446_)begin
        int_reg_array_26_12_real <= _zz_1485_;
      end
      if(_zz_1447_)begin
        int_reg_array_26_13_real <= _zz_1485_;
      end
      if(_zz_1448_)begin
        int_reg_array_26_14_real <= _zz_1485_;
      end
      if(_zz_1449_)begin
        int_reg_array_26_15_real <= _zz_1485_;
      end
      if(_zz_1450_)begin
        int_reg_array_26_16_real <= _zz_1485_;
      end
      if(_zz_1451_)begin
        int_reg_array_26_17_real <= _zz_1485_;
      end
      if(_zz_1452_)begin
        int_reg_array_26_18_real <= _zz_1485_;
      end
      if(_zz_1453_)begin
        int_reg_array_26_19_real <= _zz_1485_;
      end
      if(_zz_1454_)begin
        int_reg_array_26_20_real <= _zz_1485_;
      end
      if(_zz_1455_)begin
        int_reg_array_26_21_real <= _zz_1485_;
      end
      if(_zz_1456_)begin
        int_reg_array_26_22_real <= _zz_1485_;
      end
      if(_zz_1457_)begin
        int_reg_array_26_23_real <= _zz_1485_;
      end
      if(_zz_1458_)begin
        int_reg_array_26_24_real <= _zz_1485_;
      end
      if(_zz_1459_)begin
        int_reg_array_26_25_real <= _zz_1485_;
      end
      if(_zz_1460_)begin
        int_reg_array_26_26_real <= _zz_1485_;
      end
      if(_zz_1461_)begin
        int_reg_array_26_27_real <= _zz_1485_;
      end
      if(_zz_1462_)begin
        int_reg_array_26_28_real <= _zz_1485_;
      end
      if(_zz_1463_)begin
        int_reg_array_26_29_real <= _zz_1485_;
      end
      if(_zz_1464_)begin
        int_reg_array_26_30_real <= _zz_1485_;
      end
      if(_zz_1465_)begin
        int_reg_array_26_31_real <= _zz_1485_;
      end
      if(_zz_1466_)begin
        int_reg_array_26_32_real <= _zz_1485_;
      end
      if(_zz_1467_)begin
        int_reg_array_26_33_real <= _zz_1485_;
      end
      if(_zz_1468_)begin
        int_reg_array_26_34_real <= _zz_1485_;
      end
      if(_zz_1469_)begin
        int_reg_array_26_35_real <= _zz_1485_;
      end
      if(_zz_1470_)begin
        int_reg_array_26_36_real <= _zz_1485_;
      end
      if(_zz_1471_)begin
        int_reg_array_26_37_real <= _zz_1485_;
      end
      if(_zz_1472_)begin
        int_reg_array_26_38_real <= _zz_1485_;
      end
      if(_zz_1473_)begin
        int_reg_array_26_39_real <= _zz_1485_;
      end
      if(_zz_1474_)begin
        int_reg_array_26_40_real <= _zz_1485_;
      end
      if(_zz_1475_)begin
        int_reg_array_26_41_real <= _zz_1485_;
      end
      if(_zz_1476_)begin
        int_reg_array_26_42_real <= _zz_1485_;
      end
      if(_zz_1477_)begin
        int_reg_array_26_43_real <= _zz_1485_;
      end
      if(_zz_1478_)begin
        int_reg_array_26_44_real <= _zz_1485_;
      end
      if(_zz_1479_)begin
        int_reg_array_26_45_real <= _zz_1485_;
      end
      if(_zz_1480_)begin
        int_reg_array_26_46_real <= _zz_1485_;
      end
      if(_zz_1481_)begin
        int_reg_array_26_47_real <= _zz_1485_;
      end
      if(_zz_1482_)begin
        int_reg_array_26_48_real <= _zz_1485_;
      end
      if(_zz_1483_)begin
        int_reg_array_26_49_real <= _zz_1485_;
      end
      if(_zz_1434_)begin
        int_reg_array_26_0_imag <= _zz_1486_;
      end
      if(_zz_1435_)begin
        int_reg_array_26_1_imag <= _zz_1486_;
      end
      if(_zz_1436_)begin
        int_reg_array_26_2_imag <= _zz_1486_;
      end
      if(_zz_1437_)begin
        int_reg_array_26_3_imag <= _zz_1486_;
      end
      if(_zz_1438_)begin
        int_reg_array_26_4_imag <= _zz_1486_;
      end
      if(_zz_1439_)begin
        int_reg_array_26_5_imag <= _zz_1486_;
      end
      if(_zz_1440_)begin
        int_reg_array_26_6_imag <= _zz_1486_;
      end
      if(_zz_1441_)begin
        int_reg_array_26_7_imag <= _zz_1486_;
      end
      if(_zz_1442_)begin
        int_reg_array_26_8_imag <= _zz_1486_;
      end
      if(_zz_1443_)begin
        int_reg_array_26_9_imag <= _zz_1486_;
      end
      if(_zz_1444_)begin
        int_reg_array_26_10_imag <= _zz_1486_;
      end
      if(_zz_1445_)begin
        int_reg_array_26_11_imag <= _zz_1486_;
      end
      if(_zz_1446_)begin
        int_reg_array_26_12_imag <= _zz_1486_;
      end
      if(_zz_1447_)begin
        int_reg_array_26_13_imag <= _zz_1486_;
      end
      if(_zz_1448_)begin
        int_reg_array_26_14_imag <= _zz_1486_;
      end
      if(_zz_1449_)begin
        int_reg_array_26_15_imag <= _zz_1486_;
      end
      if(_zz_1450_)begin
        int_reg_array_26_16_imag <= _zz_1486_;
      end
      if(_zz_1451_)begin
        int_reg_array_26_17_imag <= _zz_1486_;
      end
      if(_zz_1452_)begin
        int_reg_array_26_18_imag <= _zz_1486_;
      end
      if(_zz_1453_)begin
        int_reg_array_26_19_imag <= _zz_1486_;
      end
      if(_zz_1454_)begin
        int_reg_array_26_20_imag <= _zz_1486_;
      end
      if(_zz_1455_)begin
        int_reg_array_26_21_imag <= _zz_1486_;
      end
      if(_zz_1456_)begin
        int_reg_array_26_22_imag <= _zz_1486_;
      end
      if(_zz_1457_)begin
        int_reg_array_26_23_imag <= _zz_1486_;
      end
      if(_zz_1458_)begin
        int_reg_array_26_24_imag <= _zz_1486_;
      end
      if(_zz_1459_)begin
        int_reg_array_26_25_imag <= _zz_1486_;
      end
      if(_zz_1460_)begin
        int_reg_array_26_26_imag <= _zz_1486_;
      end
      if(_zz_1461_)begin
        int_reg_array_26_27_imag <= _zz_1486_;
      end
      if(_zz_1462_)begin
        int_reg_array_26_28_imag <= _zz_1486_;
      end
      if(_zz_1463_)begin
        int_reg_array_26_29_imag <= _zz_1486_;
      end
      if(_zz_1464_)begin
        int_reg_array_26_30_imag <= _zz_1486_;
      end
      if(_zz_1465_)begin
        int_reg_array_26_31_imag <= _zz_1486_;
      end
      if(_zz_1466_)begin
        int_reg_array_26_32_imag <= _zz_1486_;
      end
      if(_zz_1467_)begin
        int_reg_array_26_33_imag <= _zz_1486_;
      end
      if(_zz_1468_)begin
        int_reg_array_26_34_imag <= _zz_1486_;
      end
      if(_zz_1469_)begin
        int_reg_array_26_35_imag <= _zz_1486_;
      end
      if(_zz_1470_)begin
        int_reg_array_26_36_imag <= _zz_1486_;
      end
      if(_zz_1471_)begin
        int_reg_array_26_37_imag <= _zz_1486_;
      end
      if(_zz_1472_)begin
        int_reg_array_26_38_imag <= _zz_1486_;
      end
      if(_zz_1473_)begin
        int_reg_array_26_39_imag <= _zz_1486_;
      end
      if(_zz_1474_)begin
        int_reg_array_26_40_imag <= _zz_1486_;
      end
      if(_zz_1475_)begin
        int_reg_array_26_41_imag <= _zz_1486_;
      end
      if(_zz_1476_)begin
        int_reg_array_26_42_imag <= _zz_1486_;
      end
      if(_zz_1477_)begin
        int_reg_array_26_43_imag <= _zz_1486_;
      end
      if(_zz_1478_)begin
        int_reg_array_26_44_imag <= _zz_1486_;
      end
      if(_zz_1479_)begin
        int_reg_array_26_45_imag <= _zz_1486_;
      end
      if(_zz_1480_)begin
        int_reg_array_26_46_imag <= _zz_1486_;
      end
      if(_zz_1481_)begin
        int_reg_array_26_47_imag <= _zz_1486_;
      end
      if(_zz_1482_)begin
        int_reg_array_26_48_imag <= _zz_1486_;
      end
      if(_zz_1483_)begin
        int_reg_array_26_49_imag <= _zz_1486_;
      end
      if(_zz_1489_)begin
        int_reg_array_27_0_real <= _zz_1540_;
      end
      if(_zz_1490_)begin
        int_reg_array_27_1_real <= _zz_1540_;
      end
      if(_zz_1491_)begin
        int_reg_array_27_2_real <= _zz_1540_;
      end
      if(_zz_1492_)begin
        int_reg_array_27_3_real <= _zz_1540_;
      end
      if(_zz_1493_)begin
        int_reg_array_27_4_real <= _zz_1540_;
      end
      if(_zz_1494_)begin
        int_reg_array_27_5_real <= _zz_1540_;
      end
      if(_zz_1495_)begin
        int_reg_array_27_6_real <= _zz_1540_;
      end
      if(_zz_1496_)begin
        int_reg_array_27_7_real <= _zz_1540_;
      end
      if(_zz_1497_)begin
        int_reg_array_27_8_real <= _zz_1540_;
      end
      if(_zz_1498_)begin
        int_reg_array_27_9_real <= _zz_1540_;
      end
      if(_zz_1499_)begin
        int_reg_array_27_10_real <= _zz_1540_;
      end
      if(_zz_1500_)begin
        int_reg_array_27_11_real <= _zz_1540_;
      end
      if(_zz_1501_)begin
        int_reg_array_27_12_real <= _zz_1540_;
      end
      if(_zz_1502_)begin
        int_reg_array_27_13_real <= _zz_1540_;
      end
      if(_zz_1503_)begin
        int_reg_array_27_14_real <= _zz_1540_;
      end
      if(_zz_1504_)begin
        int_reg_array_27_15_real <= _zz_1540_;
      end
      if(_zz_1505_)begin
        int_reg_array_27_16_real <= _zz_1540_;
      end
      if(_zz_1506_)begin
        int_reg_array_27_17_real <= _zz_1540_;
      end
      if(_zz_1507_)begin
        int_reg_array_27_18_real <= _zz_1540_;
      end
      if(_zz_1508_)begin
        int_reg_array_27_19_real <= _zz_1540_;
      end
      if(_zz_1509_)begin
        int_reg_array_27_20_real <= _zz_1540_;
      end
      if(_zz_1510_)begin
        int_reg_array_27_21_real <= _zz_1540_;
      end
      if(_zz_1511_)begin
        int_reg_array_27_22_real <= _zz_1540_;
      end
      if(_zz_1512_)begin
        int_reg_array_27_23_real <= _zz_1540_;
      end
      if(_zz_1513_)begin
        int_reg_array_27_24_real <= _zz_1540_;
      end
      if(_zz_1514_)begin
        int_reg_array_27_25_real <= _zz_1540_;
      end
      if(_zz_1515_)begin
        int_reg_array_27_26_real <= _zz_1540_;
      end
      if(_zz_1516_)begin
        int_reg_array_27_27_real <= _zz_1540_;
      end
      if(_zz_1517_)begin
        int_reg_array_27_28_real <= _zz_1540_;
      end
      if(_zz_1518_)begin
        int_reg_array_27_29_real <= _zz_1540_;
      end
      if(_zz_1519_)begin
        int_reg_array_27_30_real <= _zz_1540_;
      end
      if(_zz_1520_)begin
        int_reg_array_27_31_real <= _zz_1540_;
      end
      if(_zz_1521_)begin
        int_reg_array_27_32_real <= _zz_1540_;
      end
      if(_zz_1522_)begin
        int_reg_array_27_33_real <= _zz_1540_;
      end
      if(_zz_1523_)begin
        int_reg_array_27_34_real <= _zz_1540_;
      end
      if(_zz_1524_)begin
        int_reg_array_27_35_real <= _zz_1540_;
      end
      if(_zz_1525_)begin
        int_reg_array_27_36_real <= _zz_1540_;
      end
      if(_zz_1526_)begin
        int_reg_array_27_37_real <= _zz_1540_;
      end
      if(_zz_1527_)begin
        int_reg_array_27_38_real <= _zz_1540_;
      end
      if(_zz_1528_)begin
        int_reg_array_27_39_real <= _zz_1540_;
      end
      if(_zz_1529_)begin
        int_reg_array_27_40_real <= _zz_1540_;
      end
      if(_zz_1530_)begin
        int_reg_array_27_41_real <= _zz_1540_;
      end
      if(_zz_1531_)begin
        int_reg_array_27_42_real <= _zz_1540_;
      end
      if(_zz_1532_)begin
        int_reg_array_27_43_real <= _zz_1540_;
      end
      if(_zz_1533_)begin
        int_reg_array_27_44_real <= _zz_1540_;
      end
      if(_zz_1534_)begin
        int_reg_array_27_45_real <= _zz_1540_;
      end
      if(_zz_1535_)begin
        int_reg_array_27_46_real <= _zz_1540_;
      end
      if(_zz_1536_)begin
        int_reg_array_27_47_real <= _zz_1540_;
      end
      if(_zz_1537_)begin
        int_reg_array_27_48_real <= _zz_1540_;
      end
      if(_zz_1538_)begin
        int_reg_array_27_49_real <= _zz_1540_;
      end
      if(_zz_1489_)begin
        int_reg_array_27_0_imag <= _zz_1541_;
      end
      if(_zz_1490_)begin
        int_reg_array_27_1_imag <= _zz_1541_;
      end
      if(_zz_1491_)begin
        int_reg_array_27_2_imag <= _zz_1541_;
      end
      if(_zz_1492_)begin
        int_reg_array_27_3_imag <= _zz_1541_;
      end
      if(_zz_1493_)begin
        int_reg_array_27_4_imag <= _zz_1541_;
      end
      if(_zz_1494_)begin
        int_reg_array_27_5_imag <= _zz_1541_;
      end
      if(_zz_1495_)begin
        int_reg_array_27_6_imag <= _zz_1541_;
      end
      if(_zz_1496_)begin
        int_reg_array_27_7_imag <= _zz_1541_;
      end
      if(_zz_1497_)begin
        int_reg_array_27_8_imag <= _zz_1541_;
      end
      if(_zz_1498_)begin
        int_reg_array_27_9_imag <= _zz_1541_;
      end
      if(_zz_1499_)begin
        int_reg_array_27_10_imag <= _zz_1541_;
      end
      if(_zz_1500_)begin
        int_reg_array_27_11_imag <= _zz_1541_;
      end
      if(_zz_1501_)begin
        int_reg_array_27_12_imag <= _zz_1541_;
      end
      if(_zz_1502_)begin
        int_reg_array_27_13_imag <= _zz_1541_;
      end
      if(_zz_1503_)begin
        int_reg_array_27_14_imag <= _zz_1541_;
      end
      if(_zz_1504_)begin
        int_reg_array_27_15_imag <= _zz_1541_;
      end
      if(_zz_1505_)begin
        int_reg_array_27_16_imag <= _zz_1541_;
      end
      if(_zz_1506_)begin
        int_reg_array_27_17_imag <= _zz_1541_;
      end
      if(_zz_1507_)begin
        int_reg_array_27_18_imag <= _zz_1541_;
      end
      if(_zz_1508_)begin
        int_reg_array_27_19_imag <= _zz_1541_;
      end
      if(_zz_1509_)begin
        int_reg_array_27_20_imag <= _zz_1541_;
      end
      if(_zz_1510_)begin
        int_reg_array_27_21_imag <= _zz_1541_;
      end
      if(_zz_1511_)begin
        int_reg_array_27_22_imag <= _zz_1541_;
      end
      if(_zz_1512_)begin
        int_reg_array_27_23_imag <= _zz_1541_;
      end
      if(_zz_1513_)begin
        int_reg_array_27_24_imag <= _zz_1541_;
      end
      if(_zz_1514_)begin
        int_reg_array_27_25_imag <= _zz_1541_;
      end
      if(_zz_1515_)begin
        int_reg_array_27_26_imag <= _zz_1541_;
      end
      if(_zz_1516_)begin
        int_reg_array_27_27_imag <= _zz_1541_;
      end
      if(_zz_1517_)begin
        int_reg_array_27_28_imag <= _zz_1541_;
      end
      if(_zz_1518_)begin
        int_reg_array_27_29_imag <= _zz_1541_;
      end
      if(_zz_1519_)begin
        int_reg_array_27_30_imag <= _zz_1541_;
      end
      if(_zz_1520_)begin
        int_reg_array_27_31_imag <= _zz_1541_;
      end
      if(_zz_1521_)begin
        int_reg_array_27_32_imag <= _zz_1541_;
      end
      if(_zz_1522_)begin
        int_reg_array_27_33_imag <= _zz_1541_;
      end
      if(_zz_1523_)begin
        int_reg_array_27_34_imag <= _zz_1541_;
      end
      if(_zz_1524_)begin
        int_reg_array_27_35_imag <= _zz_1541_;
      end
      if(_zz_1525_)begin
        int_reg_array_27_36_imag <= _zz_1541_;
      end
      if(_zz_1526_)begin
        int_reg_array_27_37_imag <= _zz_1541_;
      end
      if(_zz_1527_)begin
        int_reg_array_27_38_imag <= _zz_1541_;
      end
      if(_zz_1528_)begin
        int_reg_array_27_39_imag <= _zz_1541_;
      end
      if(_zz_1529_)begin
        int_reg_array_27_40_imag <= _zz_1541_;
      end
      if(_zz_1530_)begin
        int_reg_array_27_41_imag <= _zz_1541_;
      end
      if(_zz_1531_)begin
        int_reg_array_27_42_imag <= _zz_1541_;
      end
      if(_zz_1532_)begin
        int_reg_array_27_43_imag <= _zz_1541_;
      end
      if(_zz_1533_)begin
        int_reg_array_27_44_imag <= _zz_1541_;
      end
      if(_zz_1534_)begin
        int_reg_array_27_45_imag <= _zz_1541_;
      end
      if(_zz_1535_)begin
        int_reg_array_27_46_imag <= _zz_1541_;
      end
      if(_zz_1536_)begin
        int_reg_array_27_47_imag <= _zz_1541_;
      end
      if(_zz_1537_)begin
        int_reg_array_27_48_imag <= _zz_1541_;
      end
      if(_zz_1538_)begin
        int_reg_array_27_49_imag <= _zz_1541_;
      end
      if(_zz_1544_)begin
        int_reg_array_28_0_real <= _zz_1595_;
      end
      if(_zz_1545_)begin
        int_reg_array_28_1_real <= _zz_1595_;
      end
      if(_zz_1546_)begin
        int_reg_array_28_2_real <= _zz_1595_;
      end
      if(_zz_1547_)begin
        int_reg_array_28_3_real <= _zz_1595_;
      end
      if(_zz_1548_)begin
        int_reg_array_28_4_real <= _zz_1595_;
      end
      if(_zz_1549_)begin
        int_reg_array_28_5_real <= _zz_1595_;
      end
      if(_zz_1550_)begin
        int_reg_array_28_6_real <= _zz_1595_;
      end
      if(_zz_1551_)begin
        int_reg_array_28_7_real <= _zz_1595_;
      end
      if(_zz_1552_)begin
        int_reg_array_28_8_real <= _zz_1595_;
      end
      if(_zz_1553_)begin
        int_reg_array_28_9_real <= _zz_1595_;
      end
      if(_zz_1554_)begin
        int_reg_array_28_10_real <= _zz_1595_;
      end
      if(_zz_1555_)begin
        int_reg_array_28_11_real <= _zz_1595_;
      end
      if(_zz_1556_)begin
        int_reg_array_28_12_real <= _zz_1595_;
      end
      if(_zz_1557_)begin
        int_reg_array_28_13_real <= _zz_1595_;
      end
      if(_zz_1558_)begin
        int_reg_array_28_14_real <= _zz_1595_;
      end
      if(_zz_1559_)begin
        int_reg_array_28_15_real <= _zz_1595_;
      end
      if(_zz_1560_)begin
        int_reg_array_28_16_real <= _zz_1595_;
      end
      if(_zz_1561_)begin
        int_reg_array_28_17_real <= _zz_1595_;
      end
      if(_zz_1562_)begin
        int_reg_array_28_18_real <= _zz_1595_;
      end
      if(_zz_1563_)begin
        int_reg_array_28_19_real <= _zz_1595_;
      end
      if(_zz_1564_)begin
        int_reg_array_28_20_real <= _zz_1595_;
      end
      if(_zz_1565_)begin
        int_reg_array_28_21_real <= _zz_1595_;
      end
      if(_zz_1566_)begin
        int_reg_array_28_22_real <= _zz_1595_;
      end
      if(_zz_1567_)begin
        int_reg_array_28_23_real <= _zz_1595_;
      end
      if(_zz_1568_)begin
        int_reg_array_28_24_real <= _zz_1595_;
      end
      if(_zz_1569_)begin
        int_reg_array_28_25_real <= _zz_1595_;
      end
      if(_zz_1570_)begin
        int_reg_array_28_26_real <= _zz_1595_;
      end
      if(_zz_1571_)begin
        int_reg_array_28_27_real <= _zz_1595_;
      end
      if(_zz_1572_)begin
        int_reg_array_28_28_real <= _zz_1595_;
      end
      if(_zz_1573_)begin
        int_reg_array_28_29_real <= _zz_1595_;
      end
      if(_zz_1574_)begin
        int_reg_array_28_30_real <= _zz_1595_;
      end
      if(_zz_1575_)begin
        int_reg_array_28_31_real <= _zz_1595_;
      end
      if(_zz_1576_)begin
        int_reg_array_28_32_real <= _zz_1595_;
      end
      if(_zz_1577_)begin
        int_reg_array_28_33_real <= _zz_1595_;
      end
      if(_zz_1578_)begin
        int_reg_array_28_34_real <= _zz_1595_;
      end
      if(_zz_1579_)begin
        int_reg_array_28_35_real <= _zz_1595_;
      end
      if(_zz_1580_)begin
        int_reg_array_28_36_real <= _zz_1595_;
      end
      if(_zz_1581_)begin
        int_reg_array_28_37_real <= _zz_1595_;
      end
      if(_zz_1582_)begin
        int_reg_array_28_38_real <= _zz_1595_;
      end
      if(_zz_1583_)begin
        int_reg_array_28_39_real <= _zz_1595_;
      end
      if(_zz_1584_)begin
        int_reg_array_28_40_real <= _zz_1595_;
      end
      if(_zz_1585_)begin
        int_reg_array_28_41_real <= _zz_1595_;
      end
      if(_zz_1586_)begin
        int_reg_array_28_42_real <= _zz_1595_;
      end
      if(_zz_1587_)begin
        int_reg_array_28_43_real <= _zz_1595_;
      end
      if(_zz_1588_)begin
        int_reg_array_28_44_real <= _zz_1595_;
      end
      if(_zz_1589_)begin
        int_reg_array_28_45_real <= _zz_1595_;
      end
      if(_zz_1590_)begin
        int_reg_array_28_46_real <= _zz_1595_;
      end
      if(_zz_1591_)begin
        int_reg_array_28_47_real <= _zz_1595_;
      end
      if(_zz_1592_)begin
        int_reg_array_28_48_real <= _zz_1595_;
      end
      if(_zz_1593_)begin
        int_reg_array_28_49_real <= _zz_1595_;
      end
      if(_zz_1544_)begin
        int_reg_array_28_0_imag <= _zz_1596_;
      end
      if(_zz_1545_)begin
        int_reg_array_28_1_imag <= _zz_1596_;
      end
      if(_zz_1546_)begin
        int_reg_array_28_2_imag <= _zz_1596_;
      end
      if(_zz_1547_)begin
        int_reg_array_28_3_imag <= _zz_1596_;
      end
      if(_zz_1548_)begin
        int_reg_array_28_4_imag <= _zz_1596_;
      end
      if(_zz_1549_)begin
        int_reg_array_28_5_imag <= _zz_1596_;
      end
      if(_zz_1550_)begin
        int_reg_array_28_6_imag <= _zz_1596_;
      end
      if(_zz_1551_)begin
        int_reg_array_28_7_imag <= _zz_1596_;
      end
      if(_zz_1552_)begin
        int_reg_array_28_8_imag <= _zz_1596_;
      end
      if(_zz_1553_)begin
        int_reg_array_28_9_imag <= _zz_1596_;
      end
      if(_zz_1554_)begin
        int_reg_array_28_10_imag <= _zz_1596_;
      end
      if(_zz_1555_)begin
        int_reg_array_28_11_imag <= _zz_1596_;
      end
      if(_zz_1556_)begin
        int_reg_array_28_12_imag <= _zz_1596_;
      end
      if(_zz_1557_)begin
        int_reg_array_28_13_imag <= _zz_1596_;
      end
      if(_zz_1558_)begin
        int_reg_array_28_14_imag <= _zz_1596_;
      end
      if(_zz_1559_)begin
        int_reg_array_28_15_imag <= _zz_1596_;
      end
      if(_zz_1560_)begin
        int_reg_array_28_16_imag <= _zz_1596_;
      end
      if(_zz_1561_)begin
        int_reg_array_28_17_imag <= _zz_1596_;
      end
      if(_zz_1562_)begin
        int_reg_array_28_18_imag <= _zz_1596_;
      end
      if(_zz_1563_)begin
        int_reg_array_28_19_imag <= _zz_1596_;
      end
      if(_zz_1564_)begin
        int_reg_array_28_20_imag <= _zz_1596_;
      end
      if(_zz_1565_)begin
        int_reg_array_28_21_imag <= _zz_1596_;
      end
      if(_zz_1566_)begin
        int_reg_array_28_22_imag <= _zz_1596_;
      end
      if(_zz_1567_)begin
        int_reg_array_28_23_imag <= _zz_1596_;
      end
      if(_zz_1568_)begin
        int_reg_array_28_24_imag <= _zz_1596_;
      end
      if(_zz_1569_)begin
        int_reg_array_28_25_imag <= _zz_1596_;
      end
      if(_zz_1570_)begin
        int_reg_array_28_26_imag <= _zz_1596_;
      end
      if(_zz_1571_)begin
        int_reg_array_28_27_imag <= _zz_1596_;
      end
      if(_zz_1572_)begin
        int_reg_array_28_28_imag <= _zz_1596_;
      end
      if(_zz_1573_)begin
        int_reg_array_28_29_imag <= _zz_1596_;
      end
      if(_zz_1574_)begin
        int_reg_array_28_30_imag <= _zz_1596_;
      end
      if(_zz_1575_)begin
        int_reg_array_28_31_imag <= _zz_1596_;
      end
      if(_zz_1576_)begin
        int_reg_array_28_32_imag <= _zz_1596_;
      end
      if(_zz_1577_)begin
        int_reg_array_28_33_imag <= _zz_1596_;
      end
      if(_zz_1578_)begin
        int_reg_array_28_34_imag <= _zz_1596_;
      end
      if(_zz_1579_)begin
        int_reg_array_28_35_imag <= _zz_1596_;
      end
      if(_zz_1580_)begin
        int_reg_array_28_36_imag <= _zz_1596_;
      end
      if(_zz_1581_)begin
        int_reg_array_28_37_imag <= _zz_1596_;
      end
      if(_zz_1582_)begin
        int_reg_array_28_38_imag <= _zz_1596_;
      end
      if(_zz_1583_)begin
        int_reg_array_28_39_imag <= _zz_1596_;
      end
      if(_zz_1584_)begin
        int_reg_array_28_40_imag <= _zz_1596_;
      end
      if(_zz_1585_)begin
        int_reg_array_28_41_imag <= _zz_1596_;
      end
      if(_zz_1586_)begin
        int_reg_array_28_42_imag <= _zz_1596_;
      end
      if(_zz_1587_)begin
        int_reg_array_28_43_imag <= _zz_1596_;
      end
      if(_zz_1588_)begin
        int_reg_array_28_44_imag <= _zz_1596_;
      end
      if(_zz_1589_)begin
        int_reg_array_28_45_imag <= _zz_1596_;
      end
      if(_zz_1590_)begin
        int_reg_array_28_46_imag <= _zz_1596_;
      end
      if(_zz_1591_)begin
        int_reg_array_28_47_imag <= _zz_1596_;
      end
      if(_zz_1592_)begin
        int_reg_array_28_48_imag <= _zz_1596_;
      end
      if(_zz_1593_)begin
        int_reg_array_28_49_imag <= _zz_1596_;
      end
      if(_zz_1599_)begin
        int_reg_array_29_0_real <= _zz_1650_;
      end
      if(_zz_1600_)begin
        int_reg_array_29_1_real <= _zz_1650_;
      end
      if(_zz_1601_)begin
        int_reg_array_29_2_real <= _zz_1650_;
      end
      if(_zz_1602_)begin
        int_reg_array_29_3_real <= _zz_1650_;
      end
      if(_zz_1603_)begin
        int_reg_array_29_4_real <= _zz_1650_;
      end
      if(_zz_1604_)begin
        int_reg_array_29_5_real <= _zz_1650_;
      end
      if(_zz_1605_)begin
        int_reg_array_29_6_real <= _zz_1650_;
      end
      if(_zz_1606_)begin
        int_reg_array_29_7_real <= _zz_1650_;
      end
      if(_zz_1607_)begin
        int_reg_array_29_8_real <= _zz_1650_;
      end
      if(_zz_1608_)begin
        int_reg_array_29_9_real <= _zz_1650_;
      end
      if(_zz_1609_)begin
        int_reg_array_29_10_real <= _zz_1650_;
      end
      if(_zz_1610_)begin
        int_reg_array_29_11_real <= _zz_1650_;
      end
      if(_zz_1611_)begin
        int_reg_array_29_12_real <= _zz_1650_;
      end
      if(_zz_1612_)begin
        int_reg_array_29_13_real <= _zz_1650_;
      end
      if(_zz_1613_)begin
        int_reg_array_29_14_real <= _zz_1650_;
      end
      if(_zz_1614_)begin
        int_reg_array_29_15_real <= _zz_1650_;
      end
      if(_zz_1615_)begin
        int_reg_array_29_16_real <= _zz_1650_;
      end
      if(_zz_1616_)begin
        int_reg_array_29_17_real <= _zz_1650_;
      end
      if(_zz_1617_)begin
        int_reg_array_29_18_real <= _zz_1650_;
      end
      if(_zz_1618_)begin
        int_reg_array_29_19_real <= _zz_1650_;
      end
      if(_zz_1619_)begin
        int_reg_array_29_20_real <= _zz_1650_;
      end
      if(_zz_1620_)begin
        int_reg_array_29_21_real <= _zz_1650_;
      end
      if(_zz_1621_)begin
        int_reg_array_29_22_real <= _zz_1650_;
      end
      if(_zz_1622_)begin
        int_reg_array_29_23_real <= _zz_1650_;
      end
      if(_zz_1623_)begin
        int_reg_array_29_24_real <= _zz_1650_;
      end
      if(_zz_1624_)begin
        int_reg_array_29_25_real <= _zz_1650_;
      end
      if(_zz_1625_)begin
        int_reg_array_29_26_real <= _zz_1650_;
      end
      if(_zz_1626_)begin
        int_reg_array_29_27_real <= _zz_1650_;
      end
      if(_zz_1627_)begin
        int_reg_array_29_28_real <= _zz_1650_;
      end
      if(_zz_1628_)begin
        int_reg_array_29_29_real <= _zz_1650_;
      end
      if(_zz_1629_)begin
        int_reg_array_29_30_real <= _zz_1650_;
      end
      if(_zz_1630_)begin
        int_reg_array_29_31_real <= _zz_1650_;
      end
      if(_zz_1631_)begin
        int_reg_array_29_32_real <= _zz_1650_;
      end
      if(_zz_1632_)begin
        int_reg_array_29_33_real <= _zz_1650_;
      end
      if(_zz_1633_)begin
        int_reg_array_29_34_real <= _zz_1650_;
      end
      if(_zz_1634_)begin
        int_reg_array_29_35_real <= _zz_1650_;
      end
      if(_zz_1635_)begin
        int_reg_array_29_36_real <= _zz_1650_;
      end
      if(_zz_1636_)begin
        int_reg_array_29_37_real <= _zz_1650_;
      end
      if(_zz_1637_)begin
        int_reg_array_29_38_real <= _zz_1650_;
      end
      if(_zz_1638_)begin
        int_reg_array_29_39_real <= _zz_1650_;
      end
      if(_zz_1639_)begin
        int_reg_array_29_40_real <= _zz_1650_;
      end
      if(_zz_1640_)begin
        int_reg_array_29_41_real <= _zz_1650_;
      end
      if(_zz_1641_)begin
        int_reg_array_29_42_real <= _zz_1650_;
      end
      if(_zz_1642_)begin
        int_reg_array_29_43_real <= _zz_1650_;
      end
      if(_zz_1643_)begin
        int_reg_array_29_44_real <= _zz_1650_;
      end
      if(_zz_1644_)begin
        int_reg_array_29_45_real <= _zz_1650_;
      end
      if(_zz_1645_)begin
        int_reg_array_29_46_real <= _zz_1650_;
      end
      if(_zz_1646_)begin
        int_reg_array_29_47_real <= _zz_1650_;
      end
      if(_zz_1647_)begin
        int_reg_array_29_48_real <= _zz_1650_;
      end
      if(_zz_1648_)begin
        int_reg_array_29_49_real <= _zz_1650_;
      end
      if(_zz_1599_)begin
        int_reg_array_29_0_imag <= _zz_1651_;
      end
      if(_zz_1600_)begin
        int_reg_array_29_1_imag <= _zz_1651_;
      end
      if(_zz_1601_)begin
        int_reg_array_29_2_imag <= _zz_1651_;
      end
      if(_zz_1602_)begin
        int_reg_array_29_3_imag <= _zz_1651_;
      end
      if(_zz_1603_)begin
        int_reg_array_29_4_imag <= _zz_1651_;
      end
      if(_zz_1604_)begin
        int_reg_array_29_5_imag <= _zz_1651_;
      end
      if(_zz_1605_)begin
        int_reg_array_29_6_imag <= _zz_1651_;
      end
      if(_zz_1606_)begin
        int_reg_array_29_7_imag <= _zz_1651_;
      end
      if(_zz_1607_)begin
        int_reg_array_29_8_imag <= _zz_1651_;
      end
      if(_zz_1608_)begin
        int_reg_array_29_9_imag <= _zz_1651_;
      end
      if(_zz_1609_)begin
        int_reg_array_29_10_imag <= _zz_1651_;
      end
      if(_zz_1610_)begin
        int_reg_array_29_11_imag <= _zz_1651_;
      end
      if(_zz_1611_)begin
        int_reg_array_29_12_imag <= _zz_1651_;
      end
      if(_zz_1612_)begin
        int_reg_array_29_13_imag <= _zz_1651_;
      end
      if(_zz_1613_)begin
        int_reg_array_29_14_imag <= _zz_1651_;
      end
      if(_zz_1614_)begin
        int_reg_array_29_15_imag <= _zz_1651_;
      end
      if(_zz_1615_)begin
        int_reg_array_29_16_imag <= _zz_1651_;
      end
      if(_zz_1616_)begin
        int_reg_array_29_17_imag <= _zz_1651_;
      end
      if(_zz_1617_)begin
        int_reg_array_29_18_imag <= _zz_1651_;
      end
      if(_zz_1618_)begin
        int_reg_array_29_19_imag <= _zz_1651_;
      end
      if(_zz_1619_)begin
        int_reg_array_29_20_imag <= _zz_1651_;
      end
      if(_zz_1620_)begin
        int_reg_array_29_21_imag <= _zz_1651_;
      end
      if(_zz_1621_)begin
        int_reg_array_29_22_imag <= _zz_1651_;
      end
      if(_zz_1622_)begin
        int_reg_array_29_23_imag <= _zz_1651_;
      end
      if(_zz_1623_)begin
        int_reg_array_29_24_imag <= _zz_1651_;
      end
      if(_zz_1624_)begin
        int_reg_array_29_25_imag <= _zz_1651_;
      end
      if(_zz_1625_)begin
        int_reg_array_29_26_imag <= _zz_1651_;
      end
      if(_zz_1626_)begin
        int_reg_array_29_27_imag <= _zz_1651_;
      end
      if(_zz_1627_)begin
        int_reg_array_29_28_imag <= _zz_1651_;
      end
      if(_zz_1628_)begin
        int_reg_array_29_29_imag <= _zz_1651_;
      end
      if(_zz_1629_)begin
        int_reg_array_29_30_imag <= _zz_1651_;
      end
      if(_zz_1630_)begin
        int_reg_array_29_31_imag <= _zz_1651_;
      end
      if(_zz_1631_)begin
        int_reg_array_29_32_imag <= _zz_1651_;
      end
      if(_zz_1632_)begin
        int_reg_array_29_33_imag <= _zz_1651_;
      end
      if(_zz_1633_)begin
        int_reg_array_29_34_imag <= _zz_1651_;
      end
      if(_zz_1634_)begin
        int_reg_array_29_35_imag <= _zz_1651_;
      end
      if(_zz_1635_)begin
        int_reg_array_29_36_imag <= _zz_1651_;
      end
      if(_zz_1636_)begin
        int_reg_array_29_37_imag <= _zz_1651_;
      end
      if(_zz_1637_)begin
        int_reg_array_29_38_imag <= _zz_1651_;
      end
      if(_zz_1638_)begin
        int_reg_array_29_39_imag <= _zz_1651_;
      end
      if(_zz_1639_)begin
        int_reg_array_29_40_imag <= _zz_1651_;
      end
      if(_zz_1640_)begin
        int_reg_array_29_41_imag <= _zz_1651_;
      end
      if(_zz_1641_)begin
        int_reg_array_29_42_imag <= _zz_1651_;
      end
      if(_zz_1642_)begin
        int_reg_array_29_43_imag <= _zz_1651_;
      end
      if(_zz_1643_)begin
        int_reg_array_29_44_imag <= _zz_1651_;
      end
      if(_zz_1644_)begin
        int_reg_array_29_45_imag <= _zz_1651_;
      end
      if(_zz_1645_)begin
        int_reg_array_29_46_imag <= _zz_1651_;
      end
      if(_zz_1646_)begin
        int_reg_array_29_47_imag <= _zz_1651_;
      end
      if(_zz_1647_)begin
        int_reg_array_29_48_imag <= _zz_1651_;
      end
      if(_zz_1648_)begin
        int_reg_array_29_49_imag <= _zz_1651_;
      end
      if(_zz_1654_)begin
        int_reg_array_30_0_real <= _zz_1705_;
      end
      if(_zz_1655_)begin
        int_reg_array_30_1_real <= _zz_1705_;
      end
      if(_zz_1656_)begin
        int_reg_array_30_2_real <= _zz_1705_;
      end
      if(_zz_1657_)begin
        int_reg_array_30_3_real <= _zz_1705_;
      end
      if(_zz_1658_)begin
        int_reg_array_30_4_real <= _zz_1705_;
      end
      if(_zz_1659_)begin
        int_reg_array_30_5_real <= _zz_1705_;
      end
      if(_zz_1660_)begin
        int_reg_array_30_6_real <= _zz_1705_;
      end
      if(_zz_1661_)begin
        int_reg_array_30_7_real <= _zz_1705_;
      end
      if(_zz_1662_)begin
        int_reg_array_30_8_real <= _zz_1705_;
      end
      if(_zz_1663_)begin
        int_reg_array_30_9_real <= _zz_1705_;
      end
      if(_zz_1664_)begin
        int_reg_array_30_10_real <= _zz_1705_;
      end
      if(_zz_1665_)begin
        int_reg_array_30_11_real <= _zz_1705_;
      end
      if(_zz_1666_)begin
        int_reg_array_30_12_real <= _zz_1705_;
      end
      if(_zz_1667_)begin
        int_reg_array_30_13_real <= _zz_1705_;
      end
      if(_zz_1668_)begin
        int_reg_array_30_14_real <= _zz_1705_;
      end
      if(_zz_1669_)begin
        int_reg_array_30_15_real <= _zz_1705_;
      end
      if(_zz_1670_)begin
        int_reg_array_30_16_real <= _zz_1705_;
      end
      if(_zz_1671_)begin
        int_reg_array_30_17_real <= _zz_1705_;
      end
      if(_zz_1672_)begin
        int_reg_array_30_18_real <= _zz_1705_;
      end
      if(_zz_1673_)begin
        int_reg_array_30_19_real <= _zz_1705_;
      end
      if(_zz_1674_)begin
        int_reg_array_30_20_real <= _zz_1705_;
      end
      if(_zz_1675_)begin
        int_reg_array_30_21_real <= _zz_1705_;
      end
      if(_zz_1676_)begin
        int_reg_array_30_22_real <= _zz_1705_;
      end
      if(_zz_1677_)begin
        int_reg_array_30_23_real <= _zz_1705_;
      end
      if(_zz_1678_)begin
        int_reg_array_30_24_real <= _zz_1705_;
      end
      if(_zz_1679_)begin
        int_reg_array_30_25_real <= _zz_1705_;
      end
      if(_zz_1680_)begin
        int_reg_array_30_26_real <= _zz_1705_;
      end
      if(_zz_1681_)begin
        int_reg_array_30_27_real <= _zz_1705_;
      end
      if(_zz_1682_)begin
        int_reg_array_30_28_real <= _zz_1705_;
      end
      if(_zz_1683_)begin
        int_reg_array_30_29_real <= _zz_1705_;
      end
      if(_zz_1684_)begin
        int_reg_array_30_30_real <= _zz_1705_;
      end
      if(_zz_1685_)begin
        int_reg_array_30_31_real <= _zz_1705_;
      end
      if(_zz_1686_)begin
        int_reg_array_30_32_real <= _zz_1705_;
      end
      if(_zz_1687_)begin
        int_reg_array_30_33_real <= _zz_1705_;
      end
      if(_zz_1688_)begin
        int_reg_array_30_34_real <= _zz_1705_;
      end
      if(_zz_1689_)begin
        int_reg_array_30_35_real <= _zz_1705_;
      end
      if(_zz_1690_)begin
        int_reg_array_30_36_real <= _zz_1705_;
      end
      if(_zz_1691_)begin
        int_reg_array_30_37_real <= _zz_1705_;
      end
      if(_zz_1692_)begin
        int_reg_array_30_38_real <= _zz_1705_;
      end
      if(_zz_1693_)begin
        int_reg_array_30_39_real <= _zz_1705_;
      end
      if(_zz_1694_)begin
        int_reg_array_30_40_real <= _zz_1705_;
      end
      if(_zz_1695_)begin
        int_reg_array_30_41_real <= _zz_1705_;
      end
      if(_zz_1696_)begin
        int_reg_array_30_42_real <= _zz_1705_;
      end
      if(_zz_1697_)begin
        int_reg_array_30_43_real <= _zz_1705_;
      end
      if(_zz_1698_)begin
        int_reg_array_30_44_real <= _zz_1705_;
      end
      if(_zz_1699_)begin
        int_reg_array_30_45_real <= _zz_1705_;
      end
      if(_zz_1700_)begin
        int_reg_array_30_46_real <= _zz_1705_;
      end
      if(_zz_1701_)begin
        int_reg_array_30_47_real <= _zz_1705_;
      end
      if(_zz_1702_)begin
        int_reg_array_30_48_real <= _zz_1705_;
      end
      if(_zz_1703_)begin
        int_reg_array_30_49_real <= _zz_1705_;
      end
      if(_zz_1654_)begin
        int_reg_array_30_0_imag <= _zz_1706_;
      end
      if(_zz_1655_)begin
        int_reg_array_30_1_imag <= _zz_1706_;
      end
      if(_zz_1656_)begin
        int_reg_array_30_2_imag <= _zz_1706_;
      end
      if(_zz_1657_)begin
        int_reg_array_30_3_imag <= _zz_1706_;
      end
      if(_zz_1658_)begin
        int_reg_array_30_4_imag <= _zz_1706_;
      end
      if(_zz_1659_)begin
        int_reg_array_30_5_imag <= _zz_1706_;
      end
      if(_zz_1660_)begin
        int_reg_array_30_6_imag <= _zz_1706_;
      end
      if(_zz_1661_)begin
        int_reg_array_30_7_imag <= _zz_1706_;
      end
      if(_zz_1662_)begin
        int_reg_array_30_8_imag <= _zz_1706_;
      end
      if(_zz_1663_)begin
        int_reg_array_30_9_imag <= _zz_1706_;
      end
      if(_zz_1664_)begin
        int_reg_array_30_10_imag <= _zz_1706_;
      end
      if(_zz_1665_)begin
        int_reg_array_30_11_imag <= _zz_1706_;
      end
      if(_zz_1666_)begin
        int_reg_array_30_12_imag <= _zz_1706_;
      end
      if(_zz_1667_)begin
        int_reg_array_30_13_imag <= _zz_1706_;
      end
      if(_zz_1668_)begin
        int_reg_array_30_14_imag <= _zz_1706_;
      end
      if(_zz_1669_)begin
        int_reg_array_30_15_imag <= _zz_1706_;
      end
      if(_zz_1670_)begin
        int_reg_array_30_16_imag <= _zz_1706_;
      end
      if(_zz_1671_)begin
        int_reg_array_30_17_imag <= _zz_1706_;
      end
      if(_zz_1672_)begin
        int_reg_array_30_18_imag <= _zz_1706_;
      end
      if(_zz_1673_)begin
        int_reg_array_30_19_imag <= _zz_1706_;
      end
      if(_zz_1674_)begin
        int_reg_array_30_20_imag <= _zz_1706_;
      end
      if(_zz_1675_)begin
        int_reg_array_30_21_imag <= _zz_1706_;
      end
      if(_zz_1676_)begin
        int_reg_array_30_22_imag <= _zz_1706_;
      end
      if(_zz_1677_)begin
        int_reg_array_30_23_imag <= _zz_1706_;
      end
      if(_zz_1678_)begin
        int_reg_array_30_24_imag <= _zz_1706_;
      end
      if(_zz_1679_)begin
        int_reg_array_30_25_imag <= _zz_1706_;
      end
      if(_zz_1680_)begin
        int_reg_array_30_26_imag <= _zz_1706_;
      end
      if(_zz_1681_)begin
        int_reg_array_30_27_imag <= _zz_1706_;
      end
      if(_zz_1682_)begin
        int_reg_array_30_28_imag <= _zz_1706_;
      end
      if(_zz_1683_)begin
        int_reg_array_30_29_imag <= _zz_1706_;
      end
      if(_zz_1684_)begin
        int_reg_array_30_30_imag <= _zz_1706_;
      end
      if(_zz_1685_)begin
        int_reg_array_30_31_imag <= _zz_1706_;
      end
      if(_zz_1686_)begin
        int_reg_array_30_32_imag <= _zz_1706_;
      end
      if(_zz_1687_)begin
        int_reg_array_30_33_imag <= _zz_1706_;
      end
      if(_zz_1688_)begin
        int_reg_array_30_34_imag <= _zz_1706_;
      end
      if(_zz_1689_)begin
        int_reg_array_30_35_imag <= _zz_1706_;
      end
      if(_zz_1690_)begin
        int_reg_array_30_36_imag <= _zz_1706_;
      end
      if(_zz_1691_)begin
        int_reg_array_30_37_imag <= _zz_1706_;
      end
      if(_zz_1692_)begin
        int_reg_array_30_38_imag <= _zz_1706_;
      end
      if(_zz_1693_)begin
        int_reg_array_30_39_imag <= _zz_1706_;
      end
      if(_zz_1694_)begin
        int_reg_array_30_40_imag <= _zz_1706_;
      end
      if(_zz_1695_)begin
        int_reg_array_30_41_imag <= _zz_1706_;
      end
      if(_zz_1696_)begin
        int_reg_array_30_42_imag <= _zz_1706_;
      end
      if(_zz_1697_)begin
        int_reg_array_30_43_imag <= _zz_1706_;
      end
      if(_zz_1698_)begin
        int_reg_array_30_44_imag <= _zz_1706_;
      end
      if(_zz_1699_)begin
        int_reg_array_30_45_imag <= _zz_1706_;
      end
      if(_zz_1700_)begin
        int_reg_array_30_46_imag <= _zz_1706_;
      end
      if(_zz_1701_)begin
        int_reg_array_30_47_imag <= _zz_1706_;
      end
      if(_zz_1702_)begin
        int_reg_array_30_48_imag <= _zz_1706_;
      end
      if(_zz_1703_)begin
        int_reg_array_30_49_imag <= _zz_1706_;
      end
      if(_zz_1709_)begin
        int_reg_array_31_0_real <= _zz_1760_;
      end
      if(_zz_1710_)begin
        int_reg_array_31_1_real <= _zz_1760_;
      end
      if(_zz_1711_)begin
        int_reg_array_31_2_real <= _zz_1760_;
      end
      if(_zz_1712_)begin
        int_reg_array_31_3_real <= _zz_1760_;
      end
      if(_zz_1713_)begin
        int_reg_array_31_4_real <= _zz_1760_;
      end
      if(_zz_1714_)begin
        int_reg_array_31_5_real <= _zz_1760_;
      end
      if(_zz_1715_)begin
        int_reg_array_31_6_real <= _zz_1760_;
      end
      if(_zz_1716_)begin
        int_reg_array_31_7_real <= _zz_1760_;
      end
      if(_zz_1717_)begin
        int_reg_array_31_8_real <= _zz_1760_;
      end
      if(_zz_1718_)begin
        int_reg_array_31_9_real <= _zz_1760_;
      end
      if(_zz_1719_)begin
        int_reg_array_31_10_real <= _zz_1760_;
      end
      if(_zz_1720_)begin
        int_reg_array_31_11_real <= _zz_1760_;
      end
      if(_zz_1721_)begin
        int_reg_array_31_12_real <= _zz_1760_;
      end
      if(_zz_1722_)begin
        int_reg_array_31_13_real <= _zz_1760_;
      end
      if(_zz_1723_)begin
        int_reg_array_31_14_real <= _zz_1760_;
      end
      if(_zz_1724_)begin
        int_reg_array_31_15_real <= _zz_1760_;
      end
      if(_zz_1725_)begin
        int_reg_array_31_16_real <= _zz_1760_;
      end
      if(_zz_1726_)begin
        int_reg_array_31_17_real <= _zz_1760_;
      end
      if(_zz_1727_)begin
        int_reg_array_31_18_real <= _zz_1760_;
      end
      if(_zz_1728_)begin
        int_reg_array_31_19_real <= _zz_1760_;
      end
      if(_zz_1729_)begin
        int_reg_array_31_20_real <= _zz_1760_;
      end
      if(_zz_1730_)begin
        int_reg_array_31_21_real <= _zz_1760_;
      end
      if(_zz_1731_)begin
        int_reg_array_31_22_real <= _zz_1760_;
      end
      if(_zz_1732_)begin
        int_reg_array_31_23_real <= _zz_1760_;
      end
      if(_zz_1733_)begin
        int_reg_array_31_24_real <= _zz_1760_;
      end
      if(_zz_1734_)begin
        int_reg_array_31_25_real <= _zz_1760_;
      end
      if(_zz_1735_)begin
        int_reg_array_31_26_real <= _zz_1760_;
      end
      if(_zz_1736_)begin
        int_reg_array_31_27_real <= _zz_1760_;
      end
      if(_zz_1737_)begin
        int_reg_array_31_28_real <= _zz_1760_;
      end
      if(_zz_1738_)begin
        int_reg_array_31_29_real <= _zz_1760_;
      end
      if(_zz_1739_)begin
        int_reg_array_31_30_real <= _zz_1760_;
      end
      if(_zz_1740_)begin
        int_reg_array_31_31_real <= _zz_1760_;
      end
      if(_zz_1741_)begin
        int_reg_array_31_32_real <= _zz_1760_;
      end
      if(_zz_1742_)begin
        int_reg_array_31_33_real <= _zz_1760_;
      end
      if(_zz_1743_)begin
        int_reg_array_31_34_real <= _zz_1760_;
      end
      if(_zz_1744_)begin
        int_reg_array_31_35_real <= _zz_1760_;
      end
      if(_zz_1745_)begin
        int_reg_array_31_36_real <= _zz_1760_;
      end
      if(_zz_1746_)begin
        int_reg_array_31_37_real <= _zz_1760_;
      end
      if(_zz_1747_)begin
        int_reg_array_31_38_real <= _zz_1760_;
      end
      if(_zz_1748_)begin
        int_reg_array_31_39_real <= _zz_1760_;
      end
      if(_zz_1749_)begin
        int_reg_array_31_40_real <= _zz_1760_;
      end
      if(_zz_1750_)begin
        int_reg_array_31_41_real <= _zz_1760_;
      end
      if(_zz_1751_)begin
        int_reg_array_31_42_real <= _zz_1760_;
      end
      if(_zz_1752_)begin
        int_reg_array_31_43_real <= _zz_1760_;
      end
      if(_zz_1753_)begin
        int_reg_array_31_44_real <= _zz_1760_;
      end
      if(_zz_1754_)begin
        int_reg_array_31_45_real <= _zz_1760_;
      end
      if(_zz_1755_)begin
        int_reg_array_31_46_real <= _zz_1760_;
      end
      if(_zz_1756_)begin
        int_reg_array_31_47_real <= _zz_1760_;
      end
      if(_zz_1757_)begin
        int_reg_array_31_48_real <= _zz_1760_;
      end
      if(_zz_1758_)begin
        int_reg_array_31_49_real <= _zz_1760_;
      end
      if(_zz_1709_)begin
        int_reg_array_31_0_imag <= _zz_1761_;
      end
      if(_zz_1710_)begin
        int_reg_array_31_1_imag <= _zz_1761_;
      end
      if(_zz_1711_)begin
        int_reg_array_31_2_imag <= _zz_1761_;
      end
      if(_zz_1712_)begin
        int_reg_array_31_3_imag <= _zz_1761_;
      end
      if(_zz_1713_)begin
        int_reg_array_31_4_imag <= _zz_1761_;
      end
      if(_zz_1714_)begin
        int_reg_array_31_5_imag <= _zz_1761_;
      end
      if(_zz_1715_)begin
        int_reg_array_31_6_imag <= _zz_1761_;
      end
      if(_zz_1716_)begin
        int_reg_array_31_7_imag <= _zz_1761_;
      end
      if(_zz_1717_)begin
        int_reg_array_31_8_imag <= _zz_1761_;
      end
      if(_zz_1718_)begin
        int_reg_array_31_9_imag <= _zz_1761_;
      end
      if(_zz_1719_)begin
        int_reg_array_31_10_imag <= _zz_1761_;
      end
      if(_zz_1720_)begin
        int_reg_array_31_11_imag <= _zz_1761_;
      end
      if(_zz_1721_)begin
        int_reg_array_31_12_imag <= _zz_1761_;
      end
      if(_zz_1722_)begin
        int_reg_array_31_13_imag <= _zz_1761_;
      end
      if(_zz_1723_)begin
        int_reg_array_31_14_imag <= _zz_1761_;
      end
      if(_zz_1724_)begin
        int_reg_array_31_15_imag <= _zz_1761_;
      end
      if(_zz_1725_)begin
        int_reg_array_31_16_imag <= _zz_1761_;
      end
      if(_zz_1726_)begin
        int_reg_array_31_17_imag <= _zz_1761_;
      end
      if(_zz_1727_)begin
        int_reg_array_31_18_imag <= _zz_1761_;
      end
      if(_zz_1728_)begin
        int_reg_array_31_19_imag <= _zz_1761_;
      end
      if(_zz_1729_)begin
        int_reg_array_31_20_imag <= _zz_1761_;
      end
      if(_zz_1730_)begin
        int_reg_array_31_21_imag <= _zz_1761_;
      end
      if(_zz_1731_)begin
        int_reg_array_31_22_imag <= _zz_1761_;
      end
      if(_zz_1732_)begin
        int_reg_array_31_23_imag <= _zz_1761_;
      end
      if(_zz_1733_)begin
        int_reg_array_31_24_imag <= _zz_1761_;
      end
      if(_zz_1734_)begin
        int_reg_array_31_25_imag <= _zz_1761_;
      end
      if(_zz_1735_)begin
        int_reg_array_31_26_imag <= _zz_1761_;
      end
      if(_zz_1736_)begin
        int_reg_array_31_27_imag <= _zz_1761_;
      end
      if(_zz_1737_)begin
        int_reg_array_31_28_imag <= _zz_1761_;
      end
      if(_zz_1738_)begin
        int_reg_array_31_29_imag <= _zz_1761_;
      end
      if(_zz_1739_)begin
        int_reg_array_31_30_imag <= _zz_1761_;
      end
      if(_zz_1740_)begin
        int_reg_array_31_31_imag <= _zz_1761_;
      end
      if(_zz_1741_)begin
        int_reg_array_31_32_imag <= _zz_1761_;
      end
      if(_zz_1742_)begin
        int_reg_array_31_33_imag <= _zz_1761_;
      end
      if(_zz_1743_)begin
        int_reg_array_31_34_imag <= _zz_1761_;
      end
      if(_zz_1744_)begin
        int_reg_array_31_35_imag <= _zz_1761_;
      end
      if(_zz_1745_)begin
        int_reg_array_31_36_imag <= _zz_1761_;
      end
      if(_zz_1746_)begin
        int_reg_array_31_37_imag <= _zz_1761_;
      end
      if(_zz_1747_)begin
        int_reg_array_31_38_imag <= _zz_1761_;
      end
      if(_zz_1748_)begin
        int_reg_array_31_39_imag <= _zz_1761_;
      end
      if(_zz_1749_)begin
        int_reg_array_31_40_imag <= _zz_1761_;
      end
      if(_zz_1750_)begin
        int_reg_array_31_41_imag <= _zz_1761_;
      end
      if(_zz_1751_)begin
        int_reg_array_31_42_imag <= _zz_1761_;
      end
      if(_zz_1752_)begin
        int_reg_array_31_43_imag <= _zz_1761_;
      end
      if(_zz_1753_)begin
        int_reg_array_31_44_imag <= _zz_1761_;
      end
      if(_zz_1754_)begin
        int_reg_array_31_45_imag <= _zz_1761_;
      end
      if(_zz_1755_)begin
        int_reg_array_31_46_imag <= _zz_1761_;
      end
      if(_zz_1756_)begin
        int_reg_array_31_47_imag <= _zz_1761_;
      end
      if(_zz_1757_)begin
        int_reg_array_31_48_imag <= _zz_1761_;
      end
      if(_zz_1758_)begin
        int_reg_array_31_49_imag <= _zz_1761_;
      end
      if(_zz_1764_)begin
        int_reg_array_32_0_real <= _zz_1815_;
      end
      if(_zz_1765_)begin
        int_reg_array_32_1_real <= _zz_1815_;
      end
      if(_zz_1766_)begin
        int_reg_array_32_2_real <= _zz_1815_;
      end
      if(_zz_1767_)begin
        int_reg_array_32_3_real <= _zz_1815_;
      end
      if(_zz_1768_)begin
        int_reg_array_32_4_real <= _zz_1815_;
      end
      if(_zz_1769_)begin
        int_reg_array_32_5_real <= _zz_1815_;
      end
      if(_zz_1770_)begin
        int_reg_array_32_6_real <= _zz_1815_;
      end
      if(_zz_1771_)begin
        int_reg_array_32_7_real <= _zz_1815_;
      end
      if(_zz_1772_)begin
        int_reg_array_32_8_real <= _zz_1815_;
      end
      if(_zz_1773_)begin
        int_reg_array_32_9_real <= _zz_1815_;
      end
      if(_zz_1774_)begin
        int_reg_array_32_10_real <= _zz_1815_;
      end
      if(_zz_1775_)begin
        int_reg_array_32_11_real <= _zz_1815_;
      end
      if(_zz_1776_)begin
        int_reg_array_32_12_real <= _zz_1815_;
      end
      if(_zz_1777_)begin
        int_reg_array_32_13_real <= _zz_1815_;
      end
      if(_zz_1778_)begin
        int_reg_array_32_14_real <= _zz_1815_;
      end
      if(_zz_1779_)begin
        int_reg_array_32_15_real <= _zz_1815_;
      end
      if(_zz_1780_)begin
        int_reg_array_32_16_real <= _zz_1815_;
      end
      if(_zz_1781_)begin
        int_reg_array_32_17_real <= _zz_1815_;
      end
      if(_zz_1782_)begin
        int_reg_array_32_18_real <= _zz_1815_;
      end
      if(_zz_1783_)begin
        int_reg_array_32_19_real <= _zz_1815_;
      end
      if(_zz_1784_)begin
        int_reg_array_32_20_real <= _zz_1815_;
      end
      if(_zz_1785_)begin
        int_reg_array_32_21_real <= _zz_1815_;
      end
      if(_zz_1786_)begin
        int_reg_array_32_22_real <= _zz_1815_;
      end
      if(_zz_1787_)begin
        int_reg_array_32_23_real <= _zz_1815_;
      end
      if(_zz_1788_)begin
        int_reg_array_32_24_real <= _zz_1815_;
      end
      if(_zz_1789_)begin
        int_reg_array_32_25_real <= _zz_1815_;
      end
      if(_zz_1790_)begin
        int_reg_array_32_26_real <= _zz_1815_;
      end
      if(_zz_1791_)begin
        int_reg_array_32_27_real <= _zz_1815_;
      end
      if(_zz_1792_)begin
        int_reg_array_32_28_real <= _zz_1815_;
      end
      if(_zz_1793_)begin
        int_reg_array_32_29_real <= _zz_1815_;
      end
      if(_zz_1794_)begin
        int_reg_array_32_30_real <= _zz_1815_;
      end
      if(_zz_1795_)begin
        int_reg_array_32_31_real <= _zz_1815_;
      end
      if(_zz_1796_)begin
        int_reg_array_32_32_real <= _zz_1815_;
      end
      if(_zz_1797_)begin
        int_reg_array_32_33_real <= _zz_1815_;
      end
      if(_zz_1798_)begin
        int_reg_array_32_34_real <= _zz_1815_;
      end
      if(_zz_1799_)begin
        int_reg_array_32_35_real <= _zz_1815_;
      end
      if(_zz_1800_)begin
        int_reg_array_32_36_real <= _zz_1815_;
      end
      if(_zz_1801_)begin
        int_reg_array_32_37_real <= _zz_1815_;
      end
      if(_zz_1802_)begin
        int_reg_array_32_38_real <= _zz_1815_;
      end
      if(_zz_1803_)begin
        int_reg_array_32_39_real <= _zz_1815_;
      end
      if(_zz_1804_)begin
        int_reg_array_32_40_real <= _zz_1815_;
      end
      if(_zz_1805_)begin
        int_reg_array_32_41_real <= _zz_1815_;
      end
      if(_zz_1806_)begin
        int_reg_array_32_42_real <= _zz_1815_;
      end
      if(_zz_1807_)begin
        int_reg_array_32_43_real <= _zz_1815_;
      end
      if(_zz_1808_)begin
        int_reg_array_32_44_real <= _zz_1815_;
      end
      if(_zz_1809_)begin
        int_reg_array_32_45_real <= _zz_1815_;
      end
      if(_zz_1810_)begin
        int_reg_array_32_46_real <= _zz_1815_;
      end
      if(_zz_1811_)begin
        int_reg_array_32_47_real <= _zz_1815_;
      end
      if(_zz_1812_)begin
        int_reg_array_32_48_real <= _zz_1815_;
      end
      if(_zz_1813_)begin
        int_reg_array_32_49_real <= _zz_1815_;
      end
      if(_zz_1764_)begin
        int_reg_array_32_0_imag <= _zz_1816_;
      end
      if(_zz_1765_)begin
        int_reg_array_32_1_imag <= _zz_1816_;
      end
      if(_zz_1766_)begin
        int_reg_array_32_2_imag <= _zz_1816_;
      end
      if(_zz_1767_)begin
        int_reg_array_32_3_imag <= _zz_1816_;
      end
      if(_zz_1768_)begin
        int_reg_array_32_4_imag <= _zz_1816_;
      end
      if(_zz_1769_)begin
        int_reg_array_32_5_imag <= _zz_1816_;
      end
      if(_zz_1770_)begin
        int_reg_array_32_6_imag <= _zz_1816_;
      end
      if(_zz_1771_)begin
        int_reg_array_32_7_imag <= _zz_1816_;
      end
      if(_zz_1772_)begin
        int_reg_array_32_8_imag <= _zz_1816_;
      end
      if(_zz_1773_)begin
        int_reg_array_32_9_imag <= _zz_1816_;
      end
      if(_zz_1774_)begin
        int_reg_array_32_10_imag <= _zz_1816_;
      end
      if(_zz_1775_)begin
        int_reg_array_32_11_imag <= _zz_1816_;
      end
      if(_zz_1776_)begin
        int_reg_array_32_12_imag <= _zz_1816_;
      end
      if(_zz_1777_)begin
        int_reg_array_32_13_imag <= _zz_1816_;
      end
      if(_zz_1778_)begin
        int_reg_array_32_14_imag <= _zz_1816_;
      end
      if(_zz_1779_)begin
        int_reg_array_32_15_imag <= _zz_1816_;
      end
      if(_zz_1780_)begin
        int_reg_array_32_16_imag <= _zz_1816_;
      end
      if(_zz_1781_)begin
        int_reg_array_32_17_imag <= _zz_1816_;
      end
      if(_zz_1782_)begin
        int_reg_array_32_18_imag <= _zz_1816_;
      end
      if(_zz_1783_)begin
        int_reg_array_32_19_imag <= _zz_1816_;
      end
      if(_zz_1784_)begin
        int_reg_array_32_20_imag <= _zz_1816_;
      end
      if(_zz_1785_)begin
        int_reg_array_32_21_imag <= _zz_1816_;
      end
      if(_zz_1786_)begin
        int_reg_array_32_22_imag <= _zz_1816_;
      end
      if(_zz_1787_)begin
        int_reg_array_32_23_imag <= _zz_1816_;
      end
      if(_zz_1788_)begin
        int_reg_array_32_24_imag <= _zz_1816_;
      end
      if(_zz_1789_)begin
        int_reg_array_32_25_imag <= _zz_1816_;
      end
      if(_zz_1790_)begin
        int_reg_array_32_26_imag <= _zz_1816_;
      end
      if(_zz_1791_)begin
        int_reg_array_32_27_imag <= _zz_1816_;
      end
      if(_zz_1792_)begin
        int_reg_array_32_28_imag <= _zz_1816_;
      end
      if(_zz_1793_)begin
        int_reg_array_32_29_imag <= _zz_1816_;
      end
      if(_zz_1794_)begin
        int_reg_array_32_30_imag <= _zz_1816_;
      end
      if(_zz_1795_)begin
        int_reg_array_32_31_imag <= _zz_1816_;
      end
      if(_zz_1796_)begin
        int_reg_array_32_32_imag <= _zz_1816_;
      end
      if(_zz_1797_)begin
        int_reg_array_32_33_imag <= _zz_1816_;
      end
      if(_zz_1798_)begin
        int_reg_array_32_34_imag <= _zz_1816_;
      end
      if(_zz_1799_)begin
        int_reg_array_32_35_imag <= _zz_1816_;
      end
      if(_zz_1800_)begin
        int_reg_array_32_36_imag <= _zz_1816_;
      end
      if(_zz_1801_)begin
        int_reg_array_32_37_imag <= _zz_1816_;
      end
      if(_zz_1802_)begin
        int_reg_array_32_38_imag <= _zz_1816_;
      end
      if(_zz_1803_)begin
        int_reg_array_32_39_imag <= _zz_1816_;
      end
      if(_zz_1804_)begin
        int_reg_array_32_40_imag <= _zz_1816_;
      end
      if(_zz_1805_)begin
        int_reg_array_32_41_imag <= _zz_1816_;
      end
      if(_zz_1806_)begin
        int_reg_array_32_42_imag <= _zz_1816_;
      end
      if(_zz_1807_)begin
        int_reg_array_32_43_imag <= _zz_1816_;
      end
      if(_zz_1808_)begin
        int_reg_array_32_44_imag <= _zz_1816_;
      end
      if(_zz_1809_)begin
        int_reg_array_32_45_imag <= _zz_1816_;
      end
      if(_zz_1810_)begin
        int_reg_array_32_46_imag <= _zz_1816_;
      end
      if(_zz_1811_)begin
        int_reg_array_32_47_imag <= _zz_1816_;
      end
      if(_zz_1812_)begin
        int_reg_array_32_48_imag <= _zz_1816_;
      end
      if(_zz_1813_)begin
        int_reg_array_32_49_imag <= _zz_1816_;
      end
      if(_zz_1819_)begin
        int_reg_array_33_0_real <= _zz_1870_;
      end
      if(_zz_1820_)begin
        int_reg_array_33_1_real <= _zz_1870_;
      end
      if(_zz_1821_)begin
        int_reg_array_33_2_real <= _zz_1870_;
      end
      if(_zz_1822_)begin
        int_reg_array_33_3_real <= _zz_1870_;
      end
      if(_zz_1823_)begin
        int_reg_array_33_4_real <= _zz_1870_;
      end
      if(_zz_1824_)begin
        int_reg_array_33_5_real <= _zz_1870_;
      end
      if(_zz_1825_)begin
        int_reg_array_33_6_real <= _zz_1870_;
      end
      if(_zz_1826_)begin
        int_reg_array_33_7_real <= _zz_1870_;
      end
      if(_zz_1827_)begin
        int_reg_array_33_8_real <= _zz_1870_;
      end
      if(_zz_1828_)begin
        int_reg_array_33_9_real <= _zz_1870_;
      end
      if(_zz_1829_)begin
        int_reg_array_33_10_real <= _zz_1870_;
      end
      if(_zz_1830_)begin
        int_reg_array_33_11_real <= _zz_1870_;
      end
      if(_zz_1831_)begin
        int_reg_array_33_12_real <= _zz_1870_;
      end
      if(_zz_1832_)begin
        int_reg_array_33_13_real <= _zz_1870_;
      end
      if(_zz_1833_)begin
        int_reg_array_33_14_real <= _zz_1870_;
      end
      if(_zz_1834_)begin
        int_reg_array_33_15_real <= _zz_1870_;
      end
      if(_zz_1835_)begin
        int_reg_array_33_16_real <= _zz_1870_;
      end
      if(_zz_1836_)begin
        int_reg_array_33_17_real <= _zz_1870_;
      end
      if(_zz_1837_)begin
        int_reg_array_33_18_real <= _zz_1870_;
      end
      if(_zz_1838_)begin
        int_reg_array_33_19_real <= _zz_1870_;
      end
      if(_zz_1839_)begin
        int_reg_array_33_20_real <= _zz_1870_;
      end
      if(_zz_1840_)begin
        int_reg_array_33_21_real <= _zz_1870_;
      end
      if(_zz_1841_)begin
        int_reg_array_33_22_real <= _zz_1870_;
      end
      if(_zz_1842_)begin
        int_reg_array_33_23_real <= _zz_1870_;
      end
      if(_zz_1843_)begin
        int_reg_array_33_24_real <= _zz_1870_;
      end
      if(_zz_1844_)begin
        int_reg_array_33_25_real <= _zz_1870_;
      end
      if(_zz_1845_)begin
        int_reg_array_33_26_real <= _zz_1870_;
      end
      if(_zz_1846_)begin
        int_reg_array_33_27_real <= _zz_1870_;
      end
      if(_zz_1847_)begin
        int_reg_array_33_28_real <= _zz_1870_;
      end
      if(_zz_1848_)begin
        int_reg_array_33_29_real <= _zz_1870_;
      end
      if(_zz_1849_)begin
        int_reg_array_33_30_real <= _zz_1870_;
      end
      if(_zz_1850_)begin
        int_reg_array_33_31_real <= _zz_1870_;
      end
      if(_zz_1851_)begin
        int_reg_array_33_32_real <= _zz_1870_;
      end
      if(_zz_1852_)begin
        int_reg_array_33_33_real <= _zz_1870_;
      end
      if(_zz_1853_)begin
        int_reg_array_33_34_real <= _zz_1870_;
      end
      if(_zz_1854_)begin
        int_reg_array_33_35_real <= _zz_1870_;
      end
      if(_zz_1855_)begin
        int_reg_array_33_36_real <= _zz_1870_;
      end
      if(_zz_1856_)begin
        int_reg_array_33_37_real <= _zz_1870_;
      end
      if(_zz_1857_)begin
        int_reg_array_33_38_real <= _zz_1870_;
      end
      if(_zz_1858_)begin
        int_reg_array_33_39_real <= _zz_1870_;
      end
      if(_zz_1859_)begin
        int_reg_array_33_40_real <= _zz_1870_;
      end
      if(_zz_1860_)begin
        int_reg_array_33_41_real <= _zz_1870_;
      end
      if(_zz_1861_)begin
        int_reg_array_33_42_real <= _zz_1870_;
      end
      if(_zz_1862_)begin
        int_reg_array_33_43_real <= _zz_1870_;
      end
      if(_zz_1863_)begin
        int_reg_array_33_44_real <= _zz_1870_;
      end
      if(_zz_1864_)begin
        int_reg_array_33_45_real <= _zz_1870_;
      end
      if(_zz_1865_)begin
        int_reg_array_33_46_real <= _zz_1870_;
      end
      if(_zz_1866_)begin
        int_reg_array_33_47_real <= _zz_1870_;
      end
      if(_zz_1867_)begin
        int_reg_array_33_48_real <= _zz_1870_;
      end
      if(_zz_1868_)begin
        int_reg_array_33_49_real <= _zz_1870_;
      end
      if(_zz_1819_)begin
        int_reg_array_33_0_imag <= _zz_1871_;
      end
      if(_zz_1820_)begin
        int_reg_array_33_1_imag <= _zz_1871_;
      end
      if(_zz_1821_)begin
        int_reg_array_33_2_imag <= _zz_1871_;
      end
      if(_zz_1822_)begin
        int_reg_array_33_3_imag <= _zz_1871_;
      end
      if(_zz_1823_)begin
        int_reg_array_33_4_imag <= _zz_1871_;
      end
      if(_zz_1824_)begin
        int_reg_array_33_5_imag <= _zz_1871_;
      end
      if(_zz_1825_)begin
        int_reg_array_33_6_imag <= _zz_1871_;
      end
      if(_zz_1826_)begin
        int_reg_array_33_7_imag <= _zz_1871_;
      end
      if(_zz_1827_)begin
        int_reg_array_33_8_imag <= _zz_1871_;
      end
      if(_zz_1828_)begin
        int_reg_array_33_9_imag <= _zz_1871_;
      end
      if(_zz_1829_)begin
        int_reg_array_33_10_imag <= _zz_1871_;
      end
      if(_zz_1830_)begin
        int_reg_array_33_11_imag <= _zz_1871_;
      end
      if(_zz_1831_)begin
        int_reg_array_33_12_imag <= _zz_1871_;
      end
      if(_zz_1832_)begin
        int_reg_array_33_13_imag <= _zz_1871_;
      end
      if(_zz_1833_)begin
        int_reg_array_33_14_imag <= _zz_1871_;
      end
      if(_zz_1834_)begin
        int_reg_array_33_15_imag <= _zz_1871_;
      end
      if(_zz_1835_)begin
        int_reg_array_33_16_imag <= _zz_1871_;
      end
      if(_zz_1836_)begin
        int_reg_array_33_17_imag <= _zz_1871_;
      end
      if(_zz_1837_)begin
        int_reg_array_33_18_imag <= _zz_1871_;
      end
      if(_zz_1838_)begin
        int_reg_array_33_19_imag <= _zz_1871_;
      end
      if(_zz_1839_)begin
        int_reg_array_33_20_imag <= _zz_1871_;
      end
      if(_zz_1840_)begin
        int_reg_array_33_21_imag <= _zz_1871_;
      end
      if(_zz_1841_)begin
        int_reg_array_33_22_imag <= _zz_1871_;
      end
      if(_zz_1842_)begin
        int_reg_array_33_23_imag <= _zz_1871_;
      end
      if(_zz_1843_)begin
        int_reg_array_33_24_imag <= _zz_1871_;
      end
      if(_zz_1844_)begin
        int_reg_array_33_25_imag <= _zz_1871_;
      end
      if(_zz_1845_)begin
        int_reg_array_33_26_imag <= _zz_1871_;
      end
      if(_zz_1846_)begin
        int_reg_array_33_27_imag <= _zz_1871_;
      end
      if(_zz_1847_)begin
        int_reg_array_33_28_imag <= _zz_1871_;
      end
      if(_zz_1848_)begin
        int_reg_array_33_29_imag <= _zz_1871_;
      end
      if(_zz_1849_)begin
        int_reg_array_33_30_imag <= _zz_1871_;
      end
      if(_zz_1850_)begin
        int_reg_array_33_31_imag <= _zz_1871_;
      end
      if(_zz_1851_)begin
        int_reg_array_33_32_imag <= _zz_1871_;
      end
      if(_zz_1852_)begin
        int_reg_array_33_33_imag <= _zz_1871_;
      end
      if(_zz_1853_)begin
        int_reg_array_33_34_imag <= _zz_1871_;
      end
      if(_zz_1854_)begin
        int_reg_array_33_35_imag <= _zz_1871_;
      end
      if(_zz_1855_)begin
        int_reg_array_33_36_imag <= _zz_1871_;
      end
      if(_zz_1856_)begin
        int_reg_array_33_37_imag <= _zz_1871_;
      end
      if(_zz_1857_)begin
        int_reg_array_33_38_imag <= _zz_1871_;
      end
      if(_zz_1858_)begin
        int_reg_array_33_39_imag <= _zz_1871_;
      end
      if(_zz_1859_)begin
        int_reg_array_33_40_imag <= _zz_1871_;
      end
      if(_zz_1860_)begin
        int_reg_array_33_41_imag <= _zz_1871_;
      end
      if(_zz_1861_)begin
        int_reg_array_33_42_imag <= _zz_1871_;
      end
      if(_zz_1862_)begin
        int_reg_array_33_43_imag <= _zz_1871_;
      end
      if(_zz_1863_)begin
        int_reg_array_33_44_imag <= _zz_1871_;
      end
      if(_zz_1864_)begin
        int_reg_array_33_45_imag <= _zz_1871_;
      end
      if(_zz_1865_)begin
        int_reg_array_33_46_imag <= _zz_1871_;
      end
      if(_zz_1866_)begin
        int_reg_array_33_47_imag <= _zz_1871_;
      end
      if(_zz_1867_)begin
        int_reg_array_33_48_imag <= _zz_1871_;
      end
      if(_zz_1868_)begin
        int_reg_array_33_49_imag <= _zz_1871_;
      end
      if(_zz_1874_)begin
        int_reg_array_34_0_real <= _zz_1925_;
      end
      if(_zz_1875_)begin
        int_reg_array_34_1_real <= _zz_1925_;
      end
      if(_zz_1876_)begin
        int_reg_array_34_2_real <= _zz_1925_;
      end
      if(_zz_1877_)begin
        int_reg_array_34_3_real <= _zz_1925_;
      end
      if(_zz_1878_)begin
        int_reg_array_34_4_real <= _zz_1925_;
      end
      if(_zz_1879_)begin
        int_reg_array_34_5_real <= _zz_1925_;
      end
      if(_zz_1880_)begin
        int_reg_array_34_6_real <= _zz_1925_;
      end
      if(_zz_1881_)begin
        int_reg_array_34_7_real <= _zz_1925_;
      end
      if(_zz_1882_)begin
        int_reg_array_34_8_real <= _zz_1925_;
      end
      if(_zz_1883_)begin
        int_reg_array_34_9_real <= _zz_1925_;
      end
      if(_zz_1884_)begin
        int_reg_array_34_10_real <= _zz_1925_;
      end
      if(_zz_1885_)begin
        int_reg_array_34_11_real <= _zz_1925_;
      end
      if(_zz_1886_)begin
        int_reg_array_34_12_real <= _zz_1925_;
      end
      if(_zz_1887_)begin
        int_reg_array_34_13_real <= _zz_1925_;
      end
      if(_zz_1888_)begin
        int_reg_array_34_14_real <= _zz_1925_;
      end
      if(_zz_1889_)begin
        int_reg_array_34_15_real <= _zz_1925_;
      end
      if(_zz_1890_)begin
        int_reg_array_34_16_real <= _zz_1925_;
      end
      if(_zz_1891_)begin
        int_reg_array_34_17_real <= _zz_1925_;
      end
      if(_zz_1892_)begin
        int_reg_array_34_18_real <= _zz_1925_;
      end
      if(_zz_1893_)begin
        int_reg_array_34_19_real <= _zz_1925_;
      end
      if(_zz_1894_)begin
        int_reg_array_34_20_real <= _zz_1925_;
      end
      if(_zz_1895_)begin
        int_reg_array_34_21_real <= _zz_1925_;
      end
      if(_zz_1896_)begin
        int_reg_array_34_22_real <= _zz_1925_;
      end
      if(_zz_1897_)begin
        int_reg_array_34_23_real <= _zz_1925_;
      end
      if(_zz_1898_)begin
        int_reg_array_34_24_real <= _zz_1925_;
      end
      if(_zz_1899_)begin
        int_reg_array_34_25_real <= _zz_1925_;
      end
      if(_zz_1900_)begin
        int_reg_array_34_26_real <= _zz_1925_;
      end
      if(_zz_1901_)begin
        int_reg_array_34_27_real <= _zz_1925_;
      end
      if(_zz_1902_)begin
        int_reg_array_34_28_real <= _zz_1925_;
      end
      if(_zz_1903_)begin
        int_reg_array_34_29_real <= _zz_1925_;
      end
      if(_zz_1904_)begin
        int_reg_array_34_30_real <= _zz_1925_;
      end
      if(_zz_1905_)begin
        int_reg_array_34_31_real <= _zz_1925_;
      end
      if(_zz_1906_)begin
        int_reg_array_34_32_real <= _zz_1925_;
      end
      if(_zz_1907_)begin
        int_reg_array_34_33_real <= _zz_1925_;
      end
      if(_zz_1908_)begin
        int_reg_array_34_34_real <= _zz_1925_;
      end
      if(_zz_1909_)begin
        int_reg_array_34_35_real <= _zz_1925_;
      end
      if(_zz_1910_)begin
        int_reg_array_34_36_real <= _zz_1925_;
      end
      if(_zz_1911_)begin
        int_reg_array_34_37_real <= _zz_1925_;
      end
      if(_zz_1912_)begin
        int_reg_array_34_38_real <= _zz_1925_;
      end
      if(_zz_1913_)begin
        int_reg_array_34_39_real <= _zz_1925_;
      end
      if(_zz_1914_)begin
        int_reg_array_34_40_real <= _zz_1925_;
      end
      if(_zz_1915_)begin
        int_reg_array_34_41_real <= _zz_1925_;
      end
      if(_zz_1916_)begin
        int_reg_array_34_42_real <= _zz_1925_;
      end
      if(_zz_1917_)begin
        int_reg_array_34_43_real <= _zz_1925_;
      end
      if(_zz_1918_)begin
        int_reg_array_34_44_real <= _zz_1925_;
      end
      if(_zz_1919_)begin
        int_reg_array_34_45_real <= _zz_1925_;
      end
      if(_zz_1920_)begin
        int_reg_array_34_46_real <= _zz_1925_;
      end
      if(_zz_1921_)begin
        int_reg_array_34_47_real <= _zz_1925_;
      end
      if(_zz_1922_)begin
        int_reg_array_34_48_real <= _zz_1925_;
      end
      if(_zz_1923_)begin
        int_reg_array_34_49_real <= _zz_1925_;
      end
      if(_zz_1874_)begin
        int_reg_array_34_0_imag <= _zz_1926_;
      end
      if(_zz_1875_)begin
        int_reg_array_34_1_imag <= _zz_1926_;
      end
      if(_zz_1876_)begin
        int_reg_array_34_2_imag <= _zz_1926_;
      end
      if(_zz_1877_)begin
        int_reg_array_34_3_imag <= _zz_1926_;
      end
      if(_zz_1878_)begin
        int_reg_array_34_4_imag <= _zz_1926_;
      end
      if(_zz_1879_)begin
        int_reg_array_34_5_imag <= _zz_1926_;
      end
      if(_zz_1880_)begin
        int_reg_array_34_6_imag <= _zz_1926_;
      end
      if(_zz_1881_)begin
        int_reg_array_34_7_imag <= _zz_1926_;
      end
      if(_zz_1882_)begin
        int_reg_array_34_8_imag <= _zz_1926_;
      end
      if(_zz_1883_)begin
        int_reg_array_34_9_imag <= _zz_1926_;
      end
      if(_zz_1884_)begin
        int_reg_array_34_10_imag <= _zz_1926_;
      end
      if(_zz_1885_)begin
        int_reg_array_34_11_imag <= _zz_1926_;
      end
      if(_zz_1886_)begin
        int_reg_array_34_12_imag <= _zz_1926_;
      end
      if(_zz_1887_)begin
        int_reg_array_34_13_imag <= _zz_1926_;
      end
      if(_zz_1888_)begin
        int_reg_array_34_14_imag <= _zz_1926_;
      end
      if(_zz_1889_)begin
        int_reg_array_34_15_imag <= _zz_1926_;
      end
      if(_zz_1890_)begin
        int_reg_array_34_16_imag <= _zz_1926_;
      end
      if(_zz_1891_)begin
        int_reg_array_34_17_imag <= _zz_1926_;
      end
      if(_zz_1892_)begin
        int_reg_array_34_18_imag <= _zz_1926_;
      end
      if(_zz_1893_)begin
        int_reg_array_34_19_imag <= _zz_1926_;
      end
      if(_zz_1894_)begin
        int_reg_array_34_20_imag <= _zz_1926_;
      end
      if(_zz_1895_)begin
        int_reg_array_34_21_imag <= _zz_1926_;
      end
      if(_zz_1896_)begin
        int_reg_array_34_22_imag <= _zz_1926_;
      end
      if(_zz_1897_)begin
        int_reg_array_34_23_imag <= _zz_1926_;
      end
      if(_zz_1898_)begin
        int_reg_array_34_24_imag <= _zz_1926_;
      end
      if(_zz_1899_)begin
        int_reg_array_34_25_imag <= _zz_1926_;
      end
      if(_zz_1900_)begin
        int_reg_array_34_26_imag <= _zz_1926_;
      end
      if(_zz_1901_)begin
        int_reg_array_34_27_imag <= _zz_1926_;
      end
      if(_zz_1902_)begin
        int_reg_array_34_28_imag <= _zz_1926_;
      end
      if(_zz_1903_)begin
        int_reg_array_34_29_imag <= _zz_1926_;
      end
      if(_zz_1904_)begin
        int_reg_array_34_30_imag <= _zz_1926_;
      end
      if(_zz_1905_)begin
        int_reg_array_34_31_imag <= _zz_1926_;
      end
      if(_zz_1906_)begin
        int_reg_array_34_32_imag <= _zz_1926_;
      end
      if(_zz_1907_)begin
        int_reg_array_34_33_imag <= _zz_1926_;
      end
      if(_zz_1908_)begin
        int_reg_array_34_34_imag <= _zz_1926_;
      end
      if(_zz_1909_)begin
        int_reg_array_34_35_imag <= _zz_1926_;
      end
      if(_zz_1910_)begin
        int_reg_array_34_36_imag <= _zz_1926_;
      end
      if(_zz_1911_)begin
        int_reg_array_34_37_imag <= _zz_1926_;
      end
      if(_zz_1912_)begin
        int_reg_array_34_38_imag <= _zz_1926_;
      end
      if(_zz_1913_)begin
        int_reg_array_34_39_imag <= _zz_1926_;
      end
      if(_zz_1914_)begin
        int_reg_array_34_40_imag <= _zz_1926_;
      end
      if(_zz_1915_)begin
        int_reg_array_34_41_imag <= _zz_1926_;
      end
      if(_zz_1916_)begin
        int_reg_array_34_42_imag <= _zz_1926_;
      end
      if(_zz_1917_)begin
        int_reg_array_34_43_imag <= _zz_1926_;
      end
      if(_zz_1918_)begin
        int_reg_array_34_44_imag <= _zz_1926_;
      end
      if(_zz_1919_)begin
        int_reg_array_34_45_imag <= _zz_1926_;
      end
      if(_zz_1920_)begin
        int_reg_array_34_46_imag <= _zz_1926_;
      end
      if(_zz_1921_)begin
        int_reg_array_34_47_imag <= _zz_1926_;
      end
      if(_zz_1922_)begin
        int_reg_array_34_48_imag <= _zz_1926_;
      end
      if(_zz_1923_)begin
        int_reg_array_34_49_imag <= _zz_1926_;
      end
      if(_zz_1929_)begin
        int_reg_array_35_0_real <= _zz_1980_;
      end
      if(_zz_1930_)begin
        int_reg_array_35_1_real <= _zz_1980_;
      end
      if(_zz_1931_)begin
        int_reg_array_35_2_real <= _zz_1980_;
      end
      if(_zz_1932_)begin
        int_reg_array_35_3_real <= _zz_1980_;
      end
      if(_zz_1933_)begin
        int_reg_array_35_4_real <= _zz_1980_;
      end
      if(_zz_1934_)begin
        int_reg_array_35_5_real <= _zz_1980_;
      end
      if(_zz_1935_)begin
        int_reg_array_35_6_real <= _zz_1980_;
      end
      if(_zz_1936_)begin
        int_reg_array_35_7_real <= _zz_1980_;
      end
      if(_zz_1937_)begin
        int_reg_array_35_8_real <= _zz_1980_;
      end
      if(_zz_1938_)begin
        int_reg_array_35_9_real <= _zz_1980_;
      end
      if(_zz_1939_)begin
        int_reg_array_35_10_real <= _zz_1980_;
      end
      if(_zz_1940_)begin
        int_reg_array_35_11_real <= _zz_1980_;
      end
      if(_zz_1941_)begin
        int_reg_array_35_12_real <= _zz_1980_;
      end
      if(_zz_1942_)begin
        int_reg_array_35_13_real <= _zz_1980_;
      end
      if(_zz_1943_)begin
        int_reg_array_35_14_real <= _zz_1980_;
      end
      if(_zz_1944_)begin
        int_reg_array_35_15_real <= _zz_1980_;
      end
      if(_zz_1945_)begin
        int_reg_array_35_16_real <= _zz_1980_;
      end
      if(_zz_1946_)begin
        int_reg_array_35_17_real <= _zz_1980_;
      end
      if(_zz_1947_)begin
        int_reg_array_35_18_real <= _zz_1980_;
      end
      if(_zz_1948_)begin
        int_reg_array_35_19_real <= _zz_1980_;
      end
      if(_zz_1949_)begin
        int_reg_array_35_20_real <= _zz_1980_;
      end
      if(_zz_1950_)begin
        int_reg_array_35_21_real <= _zz_1980_;
      end
      if(_zz_1951_)begin
        int_reg_array_35_22_real <= _zz_1980_;
      end
      if(_zz_1952_)begin
        int_reg_array_35_23_real <= _zz_1980_;
      end
      if(_zz_1953_)begin
        int_reg_array_35_24_real <= _zz_1980_;
      end
      if(_zz_1954_)begin
        int_reg_array_35_25_real <= _zz_1980_;
      end
      if(_zz_1955_)begin
        int_reg_array_35_26_real <= _zz_1980_;
      end
      if(_zz_1956_)begin
        int_reg_array_35_27_real <= _zz_1980_;
      end
      if(_zz_1957_)begin
        int_reg_array_35_28_real <= _zz_1980_;
      end
      if(_zz_1958_)begin
        int_reg_array_35_29_real <= _zz_1980_;
      end
      if(_zz_1959_)begin
        int_reg_array_35_30_real <= _zz_1980_;
      end
      if(_zz_1960_)begin
        int_reg_array_35_31_real <= _zz_1980_;
      end
      if(_zz_1961_)begin
        int_reg_array_35_32_real <= _zz_1980_;
      end
      if(_zz_1962_)begin
        int_reg_array_35_33_real <= _zz_1980_;
      end
      if(_zz_1963_)begin
        int_reg_array_35_34_real <= _zz_1980_;
      end
      if(_zz_1964_)begin
        int_reg_array_35_35_real <= _zz_1980_;
      end
      if(_zz_1965_)begin
        int_reg_array_35_36_real <= _zz_1980_;
      end
      if(_zz_1966_)begin
        int_reg_array_35_37_real <= _zz_1980_;
      end
      if(_zz_1967_)begin
        int_reg_array_35_38_real <= _zz_1980_;
      end
      if(_zz_1968_)begin
        int_reg_array_35_39_real <= _zz_1980_;
      end
      if(_zz_1969_)begin
        int_reg_array_35_40_real <= _zz_1980_;
      end
      if(_zz_1970_)begin
        int_reg_array_35_41_real <= _zz_1980_;
      end
      if(_zz_1971_)begin
        int_reg_array_35_42_real <= _zz_1980_;
      end
      if(_zz_1972_)begin
        int_reg_array_35_43_real <= _zz_1980_;
      end
      if(_zz_1973_)begin
        int_reg_array_35_44_real <= _zz_1980_;
      end
      if(_zz_1974_)begin
        int_reg_array_35_45_real <= _zz_1980_;
      end
      if(_zz_1975_)begin
        int_reg_array_35_46_real <= _zz_1980_;
      end
      if(_zz_1976_)begin
        int_reg_array_35_47_real <= _zz_1980_;
      end
      if(_zz_1977_)begin
        int_reg_array_35_48_real <= _zz_1980_;
      end
      if(_zz_1978_)begin
        int_reg_array_35_49_real <= _zz_1980_;
      end
      if(_zz_1929_)begin
        int_reg_array_35_0_imag <= _zz_1981_;
      end
      if(_zz_1930_)begin
        int_reg_array_35_1_imag <= _zz_1981_;
      end
      if(_zz_1931_)begin
        int_reg_array_35_2_imag <= _zz_1981_;
      end
      if(_zz_1932_)begin
        int_reg_array_35_3_imag <= _zz_1981_;
      end
      if(_zz_1933_)begin
        int_reg_array_35_4_imag <= _zz_1981_;
      end
      if(_zz_1934_)begin
        int_reg_array_35_5_imag <= _zz_1981_;
      end
      if(_zz_1935_)begin
        int_reg_array_35_6_imag <= _zz_1981_;
      end
      if(_zz_1936_)begin
        int_reg_array_35_7_imag <= _zz_1981_;
      end
      if(_zz_1937_)begin
        int_reg_array_35_8_imag <= _zz_1981_;
      end
      if(_zz_1938_)begin
        int_reg_array_35_9_imag <= _zz_1981_;
      end
      if(_zz_1939_)begin
        int_reg_array_35_10_imag <= _zz_1981_;
      end
      if(_zz_1940_)begin
        int_reg_array_35_11_imag <= _zz_1981_;
      end
      if(_zz_1941_)begin
        int_reg_array_35_12_imag <= _zz_1981_;
      end
      if(_zz_1942_)begin
        int_reg_array_35_13_imag <= _zz_1981_;
      end
      if(_zz_1943_)begin
        int_reg_array_35_14_imag <= _zz_1981_;
      end
      if(_zz_1944_)begin
        int_reg_array_35_15_imag <= _zz_1981_;
      end
      if(_zz_1945_)begin
        int_reg_array_35_16_imag <= _zz_1981_;
      end
      if(_zz_1946_)begin
        int_reg_array_35_17_imag <= _zz_1981_;
      end
      if(_zz_1947_)begin
        int_reg_array_35_18_imag <= _zz_1981_;
      end
      if(_zz_1948_)begin
        int_reg_array_35_19_imag <= _zz_1981_;
      end
      if(_zz_1949_)begin
        int_reg_array_35_20_imag <= _zz_1981_;
      end
      if(_zz_1950_)begin
        int_reg_array_35_21_imag <= _zz_1981_;
      end
      if(_zz_1951_)begin
        int_reg_array_35_22_imag <= _zz_1981_;
      end
      if(_zz_1952_)begin
        int_reg_array_35_23_imag <= _zz_1981_;
      end
      if(_zz_1953_)begin
        int_reg_array_35_24_imag <= _zz_1981_;
      end
      if(_zz_1954_)begin
        int_reg_array_35_25_imag <= _zz_1981_;
      end
      if(_zz_1955_)begin
        int_reg_array_35_26_imag <= _zz_1981_;
      end
      if(_zz_1956_)begin
        int_reg_array_35_27_imag <= _zz_1981_;
      end
      if(_zz_1957_)begin
        int_reg_array_35_28_imag <= _zz_1981_;
      end
      if(_zz_1958_)begin
        int_reg_array_35_29_imag <= _zz_1981_;
      end
      if(_zz_1959_)begin
        int_reg_array_35_30_imag <= _zz_1981_;
      end
      if(_zz_1960_)begin
        int_reg_array_35_31_imag <= _zz_1981_;
      end
      if(_zz_1961_)begin
        int_reg_array_35_32_imag <= _zz_1981_;
      end
      if(_zz_1962_)begin
        int_reg_array_35_33_imag <= _zz_1981_;
      end
      if(_zz_1963_)begin
        int_reg_array_35_34_imag <= _zz_1981_;
      end
      if(_zz_1964_)begin
        int_reg_array_35_35_imag <= _zz_1981_;
      end
      if(_zz_1965_)begin
        int_reg_array_35_36_imag <= _zz_1981_;
      end
      if(_zz_1966_)begin
        int_reg_array_35_37_imag <= _zz_1981_;
      end
      if(_zz_1967_)begin
        int_reg_array_35_38_imag <= _zz_1981_;
      end
      if(_zz_1968_)begin
        int_reg_array_35_39_imag <= _zz_1981_;
      end
      if(_zz_1969_)begin
        int_reg_array_35_40_imag <= _zz_1981_;
      end
      if(_zz_1970_)begin
        int_reg_array_35_41_imag <= _zz_1981_;
      end
      if(_zz_1971_)begin
        int_reg_array_35_42_imag <= _zz_1981_;
      end
      if(_zz_1972_)begin
        int_reg_array_35_43_imag <= _zz_1981_;
      end
      if(_zz_1973_)begin
        int_reg_array_35_44_imag <= _zz_1981_;
      end
      if(_zz_1974_)begin
        int_reg_array_35_45_imag <= _zz_1981_;
      end
      if(_zz_1975_)begin
        int_reg_array_35_46_imag <= _zz_1981_;
      end
      if(_zz_1976_)begin
        int_reg_array_35_47_imag <= _zz_1981_;
      end
      if(_zz_1977_)begin
        int_reg_array_35_48_imag <= _zz_1981_;
      end
      if(_zz_1978_)begin
        int_reg_array_35_49_imag <= _zz_1981_;
      end
      if(_zz_1984_)begin
        int_reg_array_36_0_real <= _zz_2035_;
      end
      if(_zz_1985_)begin
        int_reg_array_36_1_real <= _zz_2035_;
      end
      if(_zz_1986_)begin
        int_reg_array_36_2_real <= _zz_2035_;
      end
      if(_zz_1987_)begin
        int_reg_array_36_3_real <= _zz_2035_;
      end
      if(_zz_1988_)begin
        int_reg_array_36_4_real <= _zz_2035_;
      end
      if(_zz_1989_)begin
        int_reg_array_36_5_real <= _zz_2035_;
      end
      if(_zz_1990_)begin
        int_reg_array_36_6_real <= _zz_2035_;
      end
      if(_zz_1991_)begin
        int_reg_array_36_7_real <= _zz_2035_;
      end
      if(_zz_1992_)begin
        int_reg_array_36_8_real <= _zz_2035_;
      end
      if(_zz_1993_)begin
        int_reg_array_36_9_real <= _zz_2035_;
      end
      if(_zz_1994_)begin
        int_reg_array_36_10_real <= _zz_2035_;
      end
      if(_zz_1995_)begin
        int_reg_array_36_11_real <= _zz_2035_;
      end
      if(_zz_1996_)begin
        int_reg_array_36_12_real <= _zz_2035_;
      end
      if(_zz_1997_)begin
        int_reg_array_36_13_real <= _zz_2035_;
      end
      if(_zz_1998_)begin
        int_reg_array_36_14_real <= _zz_2035_;
      end
      if(_zz_1999_)begin
        int_reg_array_36_15_real <= _zz_2035_;
      end
      if(_zz_2000_)begin
        int_reg_array_36_16_real <= _zz_2035_;
      end
      if(_zz_2001_)begin
        int_reg_array_36_17_real <= _zz_2035_;
      end
      if(_zz_2002_)begin
        int_reg_array_36_18_real <= _zz_2035_;
      end
      if(_zz_2003_)begin
        int_reg_array_36_19_real <= _zz_2035_;
      end
      if(_zz_2004_)begin
        int_reg_array_36_20_real <= _zz_2035_;
      end
      if(_zz_2005_)begin
        int_reg_array_36_21_real <= _zz_2035_;
      end
      if(_zz_2006_)begin
        int_reg_array_36_22_real <= _zz_2035_;
      end
      if(_zz_2007_)begin
        int_reg_array_36_23_real <= _zz_2035_;
      end
      if(_zz_2008_)begin
        int_reg_array_36_24_real <= _zz_2035_;
      end
      if(_zz_2009_)begin
        int_reg_array_36_25_real <= _zz_2035_;
      end
      if(_zz_2010_)begin
        int_reg_array_36_26_real <= _zz_2035_;
      end
      if(_zz_2011_)begin
        int_reg_array_36_27_real <= _zz_2035_;
      end
      if(_zz_2012_)begin
        int_reg_array_36_28_real <= _zz_2035_;
      end
      if(_zz_2013_)begin
        int_reg_array_36_29_real <= _zz_2035_;
      end
      if(_zz_2014_)begin
        int_reg_array_36_30_real <= _zz_2035_;
      end
      if(_zz_2015_)begin
        int_reg_array_36_31_real <= _zz_2035_;
      end
      if(_zz_2016_)begin
        int_reg_array_36_32_real <= _zz_2035_;
      end
      if(_zz_2017_)begin
        int_reg_array_36_33_real <= _zz_2035_;
      end
      if(_zz_2018_)begin
        int_reg_array_36_34_real <= _zz_2035_;
      end
      if(_zz_2019_)begin
        int_reg_array_36_35_real <= _zz_2035_;
      end
      if(_zz_2020_)begin
        int_reg_array_36_36_real <= _zz_2035_;
      end
      if(_zz_2021_)begin
        int_reg_array_36_37_real <= _zz_2035_;
      end
      if(_zz_2022_)begin
        int_reg_array_36_38_real <= _zz_2035_;
      end
      if(_zz_2023_)begin
        int_reg_array_36_39_real <= _zz_2035_;
      end
      if(_zz_2024_)begin
        int_reg_array_36_40_real <= _zz_2035_;
      end
      if(_zz_2025_)begin
        int_reg_array_36_41_real <= _zz_2035_;
      end
      if(_zz_2026_)begin
        int_reg_array_36_42_real <= _zz_2035_;
      end
      if(_zz_2027_)begin
        int_reg_array_36_43_real <= _zz_2035_;
      end
      if(_zz_2028_)begin
        int_reg_array_36_44_real <= _zz_2035_;
      end
      if(_zz_2029_)begin
        int_reg_array_36_45_real <= _zz_2035_;
      end
      if(_zz_2030_)begin
        int_reg_array_36_46_real <= _zz_2035_;
      end
      if(_zz_2031_)begin
        int_reg_array_36_47_real <= _zz_2035_;
      end
      if(_zz_2032_)begin
        int_reg_array_36_48_real <= _zz_2035_;
      end
      if(_zz_2033_)begin
        int_reg_array_36_49_real <= _zz_2035_;
      end
      if(_zz_1984_)begin
        int_reg_array_36_0_imag <= _zz_2036_;
      end
      if(_zz_1985_)begin
        int_reg_array_36_1_imag <= _zz_2036_;
      end
      if(_zz_1986_)begin
        int_reg_array_36_2_imag <= _zz_2036_;
      end
      if(_zz_1987_)begin
        int_reg_array_36_3_imag <= _zz_2036_;
      end
      if(_zz_1988_)begin
        int_reg_array_36_4_imag <= _zz_2036_;
      end
      if(_zz_1989_)begin
        int_reg_array_36_5_imag <= _zz_2036_;
      end
      if(_zz_1990_)begin
        int_reg_array_36_6_imag <= _zz_2036_;
      end
      if(_zz_1991_)begin
        int_reg_array_36_7_imag <= _zz_2036_;
      end
      if(_zz_1992_)begin
        int_reg_array_36_8_imag <= _zz_2036_;
      end
      if(_zz_1993_)begin
        int_reg_array_36_9_imag <= _zz_2036_;
      end
      if(_zz_1994_)begin
        int_reg_array_36_10_imag <= _zz_2036_;
      end
      if(_zz_1995_)begin
        int_reg_array_36_11_imag <= _zz_2036_;
      end
      if(_zz_1996_)begin
        int_reg_array_36_12_imag <= _zz_2036_;
      end
      if(_zz_1997_)begin
        int_reg_array_36_13_imag <= _zz_2036_;
      end
      if(_zz_1998_)begin
        int_reg_array_36_14_imag <= _zz_2036_;
      end
      if(_zz_1999_)begin
        int_reg_array_36_15_imag <= _zz_2036_;
      end
      if(_zz_2000_)begin
        int_reg_array_36_16_imag <= _zz_2036_;
      end
      if(_zz_2001_)begin
        int_reg_array_36_17_imag <= _zz_2036_;
      end
      if(_zz_2002_)begin
        int_reg_array_36_18_imag <= _zz_2036_;
      end
      if(_zz_2003_)begin
        int_reg_array_36_19_imag <= _zz_2036_;
      end
      if(_zz_2004_)begin
        int_reg_array_36_20_imag <= _zz_2036_;
      end
      if(_zz_2005_)begin
        int_reg_array_36_21_imag <= _zz_2036_;
      end
      if(_zz_2006_)begin
        int_reg_array_36_22_imag <= _zz_2036_;
      end
      if(_zz_2007_)begin
        int_reg_array_36_23_imag <= _zz_2036_;
      end
      if(_zz_2008_)begin
        int_reg_array_36_24_imag <= _zz_2036_;
      end
      if(_zz_2009_)begin
        int_reg_array_36_25_imag <= _zz_2036_;
      end
      if(_zz_2010_)begin
        int_reg_array_36_26_imag <= _zz_2036_;
      end
      if(_zz_2011_)begin
        int_reg_array_36_27_imag <= _zz_2036_;
      end
      if(_zz_2012_)begin
        int_reg_array_36_28_imag <= _zz_2036_;
      end
      if(_zz_2013_)begin
        int_reg_array_36_29_imag <= _zz_2036_;
      end
      if(_zz_2014_)begin
        int_reg_array_36_30_imag <= _zz_2036_;
      end
      if(_zz_2015_)begin
        int_reg_array_36_31_imag <= _zz_2036_;
      end
      if(_zz_2016_)begin
        int_reg_array_36_32_imag <= _zz_2036_;
      end
      if(_zz_2017_)begin
        int_reg_array_36_33_imag <= _zz_2036_;
      end
      if(_zz_2018_)begin
        int_reg_array_36_34_imag <= _zz_2036_;
      end
      if(_zz_2019_)begin
        int_reg_array_36_35_imag <= _zz_2036_;
      end
      if(_zz_2020_)begin
        int_reg_array_36_36_imag <= _zz_2036_;
      end
      if(_zz_2021_)begin
        int_reg_array_36_37_imag <= _zz_2036_;
      end
      if(_zz_2022_)begin
        int_reg_array_36_38_imag <= _zz_2036_;
      end
      if(_zz_2023_)begin
        int_reg_array_36_39_imag <= _zz_2036_;
      end
      if(_zz_2024_)begin
        int_reg_array_36_40_imag <= _zz_2036_;
      end
      if(_zz_2025_)begin
        int_reg_array_36_41_imag <= _zz_2036_;
      end
      if(_zz_2026_)begin
        int_reg_array_36_42_imag <= _zz_2036_;
      end
      if(_zz_2027_)begin
        int_reg_array_36_43_imag <= _zz_2036_;
      end
      if(_zz_2028_)begin
        int_reg_array_36_44_imag <= _zz_2036_;
      end
      if(_zz_2029_)begin
        int_reg_array_36_45_imag <= _zz_2036_;
      end
      if(_zz_2030_)begin
        int_reg_array_36_46_imag <= _zz_2036_;
      end
      if(_zz_2031_)begin
        int_reg_array_36_47_imag <= _zz_2036_;
      end
      if(_zz_2032_)begin
        int_reg_array_36_48_imag <= _zz_2036_;
      end
      if(_zz_2033_)begin
        int_reg_array_36_49_imag <= _zz_2036_;
      end
      if(_zz_2039_)begin
        int_reg_array_37_0_real <= _zz_2090_;
      end
      if(_zz_2040_)begin
        int_reg_array_37_1_real <= _zz_2090_;
      end
      if(_zz_2041_)begin
        int_reg_array_37_2_real <= _zz_2090_;
      end
      if(_zz_2042_)begin
        int_reg_array_37_3_real <= _zz_2090_;
      end
      if(_zz_2043_)begin
        int_reg_array_37_4_real <= _zz_2090_;
      end
      if(_zz_2044_)begin
        int_reg_array_37_5_real <= _zz_2090_;
      end
      if(_zz_2045_)begin
        int_reg_array_37_6_real <= _zz_2090_;
      end
      if(_zz_2046_)begin
        int_reg_array_37_7_real <= _zz_2090_;
      end
      if(_zz_2047_)begin
        int_reg_array_37_8_real <= _zz_2090_;
      end
      if(_zz_2048_)begin
        int_reg_array_37_9_real <= _zz_2090_;
      end
      if(_zz_2049_)begin
        int_reg_array_37_10_real <= _zz_2090_;
      end
      if(_zz_2050_)begin
        int_reg_array_37_11_real <= _zz_2090_;
      end
      if(_zz_2051_)begin
        int_reg_array_37_12_real <= _zz_2090_;
      end
      if(_zz_2052_)begin
        int_reg_array_37_13_real <= _zz_2090_;
      end
      if(_zz_2053_)begin
        int_reg_array_37_14_real <= _zz_2090_;
      end
      if(_zz_2054_)begin
        int_reg_array_37_15_real <= _zz_2090_;
      end
      if(_zz_2055_)begin
        int_reg_array_37_16_real <= _zz_2090_;
      end
      if(_zz_2056_)begin
        int_reg_array_37_17_real <= _zz_2090_;
      end
      if(_zz_2057_)begin
        int_reg_array_37_18_real <= _zz_2090_;
      end
      if(_zz_2058_)begin
        int_reg_array_37_19_real <= _zz_2090_;
      end
      if(_zz_2059_)begin
        int_reg_array_37_20_real <= _zz_2090_;
      end
      if(_zz_2060_)begin
        int_reg_array_37_21_real <= _zz_2090_;
      end
      if(_zz_2061_)begin
        int_reg_array_37_22_real <= _zz_2090_;
      end
      if(_zz_2062_)begin
        int_reg_array_37_23_real <= _zz_2090_;
      end
      if(_zz_2063_)begin
        int_reg_array_37_24_real <= _zz_2090_;
      end
      if(_zz_2064_)begin
        int_reg_array_37_25_real <= _zz_2090_;
      end
      if(_zz_2065_)begin
        int_reg_array_37_26_real <= _zz_2090_;
      end
      if(_zz_2066_)begin
        int_reg_array_37_27_real <= _zz_2090_;
      end
      if(_zz_2067_)begin
        int_reg_array_37_28_real <= _zz_2090_;
      end
      if(_zz_2068_)begin
        int_reg_array_37_29_real <= _zz_2090_;
      end
      if(_zz_2069_)begin
        int_reg_array_37_30_real <= _zz_2090_;
      end
      if(_zz_2070_)begin
        int_reg_array_37_31_real <= _zz_2090_;
      end
      if(_zz_2071_)begin
        int_reg_array_37_32_real <= _zz_2090_;
      end
      if(_zz_2072_)begin
        int_reg_array_37_33_real <= _zz_2090_;
      end
      if(_zz_2073_)begin
        int_reg_array_37_34_real <= _zz_2090_;
      end
      if(_zz_2074_)begin
        int_reg_array_37_35_real <= _zz_2090_;
      end
      if(_zz_2075_)begin
        int_reg_array_37_36_real <= _zz_2090_;
      end
      if(_zz_2076_)begin
        int_reg_array_37_37_real <= _zz_2090_;
      end
      if(_zz_2077_)begin
        int_reg_array_37_38_real <= _zz_2090_;
      end
      if(_zz_2078_)begin
        int_reg_array_37_39_real <= _zz_2090_;
      end
      if(_zz_2079_)begin
        int_reg_array_37_40_real <= _zz_2090_;
      end
      if(_zz_2080_)begin
        int_reg_array_37_41_real <= _zz_2090_;
      end
      if(_zz_2081_)begin
        int_reg_array_37_42_real <= _zz_2090_;
      end
      if(_zz_2082_)begin
        int_reg_array_37_43_real <= _zz_2090_;
      end
      if(_zz_2083_)begin
        int_reg_array_37_44_real <= _zz_2090_;
      end
      if(_zz_2084_)begin
        int_reg_array_37_45_real <= _zz_2090_;
      end
      if(_zz_2085_)begin
        int_reg_array_37_46_real <= _zz_2090_;
      end
      if(_zz_2086_)begin
        int_reg_array_37_47_real <= _zz_2090_;
      end
      if(_zz_2087_)begin
        int_reg_array_37_48_real <= _zz_2090_;
      end
      if(_zz_2088_)begin
        int_reg_array_37_49_real <= _zz_2090_;
      end
      if(_zz_2039_)begin
        int_reg_array_37_0_imag <= _zz_2091_;
      end
      if(_zz_2040_)begin
        int_reg_array_37_1_imag <= _zz_2091_;
      end
      if(_zz_2041_)begin
        int_reg_array_37_2_imag <= _zz_2091_;
      end
      if(_zz_2042_)begin
        int_reg_array_37_3_imag <= _zz_2091_;
      end
      if(_zz_2043_)begin
        int_reg_array_37_4_imag <= _zz_2091_;
      end
      if(_zz_2044_)begin
        int_reg_array_37_5_imag <= _zz_2091_;
      end
      if(_zz_2045_)begin
        int_reg_array_37_6_imag <= _zz_2091_;
      end
      if(_zz_2046_)begin
        int_reg_array_37_7_imag <= _zz_2091_;
      end
      if(_zz_2047_)begin
        int_reg_array_37_8_imag <= _zz_2091_;
      end
      if(_zz_2048_)begin
        int_reg_array_37_9_imag <= _zz_2091_;
      end
      if(_zz_2049_)begin
        int_reg_array_37_10_imag <= _zz_2091_;
      end
      if(_zz_2050_)begin
        int_reg_array_37_11_imag <= _zz_2091_;
      end
      if(_zz_2051_)begin
        int_reg_array_37_12_imag <= _zz_2091_;
      end
      if(_zz_2052_)begin
        int_reg_array_37_13_imag <= _zz_2091_;
      end
      if(_zz_2053_)begin
        int_reg_array_37_14_imag <= _zz_2091_;
      end
      if(_zz_2054_)begin
        int_reg_array_37_15_imag <= _zz_2091_;
      end
      if(_zz_2055_)begin
        int_reg_array_37_16_imag <= _zz_2091_;
      end
      if(_zz_2056_)begin
        int_reg_array_37_17_imag <= _zz_2091_;
      end
      if(_zz_2057_)begin
        int_reg_array_37_18_imag <= _zz_2091_;
      end
      if(_zz_2058_)begin
        int_reg_array_37_19_imag <= _zz_2091_;
      end
      if(_zz_2059_)begin
        int_reg_array_37_20_imag <= _zz_2091_;
      end
      if(_zz_2060_)begin
        int_reg_array_37_21_imag <= _zz_2091_;
      end
      if(_zz_2061_)begin
        int_reg_array_37_22_imag <= _zz_2091_;
      end
      if(_zz_2062_)begin
        int_reg_array_37_23_imag <= _zz_2091_;
      end
      if(_zz_2063_)begin
        int_reg_array_37_24_imag <= _zz_2091_;
      end
      if(_zz_2064_)begin
        int_reg_array_37_25_imag <= _zz_2091_;
      end
      if(_zz_2065_)begin
        int_reg_array_37_26_imag <= _zz_2091_;
      end
      if(_zz_2066_)begin
        int_reg_array_37_27_imag <= _zz_2091_;
      end
      if(_zz_2067_)begin
        int_reg_array_37_28_imag <= _zz_2091_;
      end
      if(_zz_2068_)begin
        int_reg_array_37_29_imag <= _zz_2091_;
      end
      if(_zz_2069_)begin
        int_reg_array_37_30_imag <= _zz_2091_;
      end
      if(_zz_2070_)begin
        int_reg_array_37_31_imag <= _zz_2091_;
      end
      if(_zz_2071_)begin
        int_reg_array_37_32_imag <= _zz_2091_;
      end
      if(_zz_2072_)begin
        int_reg_array_37_33_imag <= _zz_2091_;
      end
      if(_zz_2073_)begin
        int_reg_array_37_34_imag <= _zz_2091_;
      end
      if(_zz_2074_)begin
        int_reg_array_37_35_imag <= _zz_2091_;
      end
      if(_zz_2075_)begin
        int_reg_array_37_36_imag <= _zz_2091_;
      end
      if(_zz_2076_)begin
        int_reg_array_37_37_imag <= _zz_2091_;
      end
      if(_zz_2077_)begin
        int_reg_array_37_38_imag <= _zz_2091_;
      end
      if(_zz_2078_)begin
        int_reg_array_37_39_imag <= _zz_2091_;
      end
      if(_zz_2079_)begin
        int_reg_array_37_40_imag <= _zz_2091_;
      end
      if(_zz_2080_)begin
        int_reg_array_37_41_imag <= _zz_2091_;
      end
      if(_zz_2081_)begin
        int_reg_array_37_42_imag <= _zz_2091_;
      end
      if(_zz_2082_)begin
        int_reg_array_37_43_imag <= _zz_2091_;
      end
      if(_zz_2083_)begin
        int_reg_array_37_44_imag <= _zz_2091_;
      end
      if(_zz_2084_)begin
        int_reg_array_37_45_imag <= _zz_2091_;
      end
      if(_zz_2085_)begin
        int_reg_array_37_46_imag <= _zz_2091_;
      end
      if(_zz_2086_)begin
        int_reg_array_37_47_imag <= _zz_2091_;
      end
      if(_zz_2087_)begin
        int_reg_array_37_48_imag <= _zz_2091_;
      end
      if(_zz_2088_)begin
        int_reg_array_37_49_imag <= _zz_2091_;
      end
      if(_zz_2094_)begin
        int_reg_array_38_0_real <= _zz_2145_;
      end
      if(_zz_2095_)begin
        int_reg_array_38_1_real <= _zz_2145_;
      end
      if(_zz_2096_)begin
        int_reg_array_38_2_real <= _zz_2145_;
      end
      if(_zz_2097_)begin
        int_reg_array_38_3_real <= _zz_2145_;
      end
      if(_zz_2098_)begin
        int_reg_array_38_4_real <= _zz_2145_;
      end
      if(_zz_2099_)begin
        int_reg_array_38_5_real <= _zz_2145_;
      end
      if(_zz_2100_)begin
        int_reg_array_38_6_real <= _zz_2145_;
      end
      if(_zz_2101_)begin
        int_reg_array_38_7_real <= _zz_2145_;
      end
      if(_zz_2102_)begin
        int_reg_array_38_8_real <= _zz_2145_;
      end
      if(_zz_2103_)begin
        int_reg_array_38_9_real <= _zz_2145_;
      end
      if(_zz_2104_)begin
        int_reg_array_38_10_real <= _zz_2145_;
      end
      if(_zz_2105_)begin
        int_reg_array_38_11_real <= _zz_2145_;
      end
      if(_zz_2106_)begin
        int_reg_array_38_12_real <= _zz_2145_;
      end
      if(_zz_2107_)begin
        int_reg_array_38_13_real <= _zz_2145_;
      end
      if(_zz_2108_)begin
        int_reg_array_38_14_real <= _zz_2145_;
      end
      if(_zz_2109_)begin
        int_reg_array_38_15_real <= _zz_2145_;
      end
      if(_zz_2110_)begin
        int_reg_array_38_16_real <= _zz_2145_;
      end
      if(_zz_2111_)begin
        int_reg_array_38_17_real <= _zz_2145_;
      end
      if(_zz_2112_)begin
        int_reg_array_38_18_real <= _zz_2145_;
      end
      if(_zz_2113_)begin
        int_reg_array_38_19_real <= _zz_2145_;
      end
      if(_zz_2114_)begin
        int_reg_array_38_20_real <= _zz_2145_;
      end
      if(_zz_2115_)begin
        int_reg_array_38_21_real <= _zz_2145_;
      end
      if(_zz_2116_)begin
        int_reg_array_38_22_real <= _zz_2145_;
      end
      if(_zz_2117_)begin
        int_reg_array_38_23_real <= _zz_2145_;
      end
      if(_zz_2118_)begin
        int_reg_array_38_24_real <= _zz_2145_;
      end
      if(_zz_2119_)begin
        int_reg_array_38_25_real <= _zz_2145_;
      end
      if(_zz_2120_)begin
        int_reg_array_38_26_real <= _zz_2145_;
      end
      if(_zz_2121_)begin
        int_reg_array_38_27_real <= _zz_2145_;
      end
      if(_zz_2122_)begin
        int_reg_array_38_28_real <= _zz_2145_;
      end
      if(_zz_2123_)begin
        int_reg_array_38_29_real <= _zz_2145_;
      end
      if(_zz_2124_)begin
        int_reg_array_38_30_real <= _zz_2145_;
      end
      if(_zz_2125_)begin
        int_reg_array_38_31_real <= _zz_2145_;
      end
      if(_zz_2126_)begin
        int_reg_array_38_32_real <= _zz_2145_;
      end
      if(_zz_2127_)begin
        int_reg_array_38_33_real <= _zz_2145_;
      end
      if(_zz_2128_)begin
        int_reg_array_38_34_real <= _zz_2145_;
      end
      if(_zz_2129_)begin
        int_reg_array_38_35_real <= _zz_2145_;
      end
      if(_zz_2130_)begin
        int_reg_array_38_36_real <= _zz_2145_;
      end
      if(_zz_2131_)begin
        int_reg_array_38_37_real <= _zz_2145_;
      end
      if(_zz_2132_)begin
        int_reg_array_38_38_real <= _zz_2145_;
      end
      if(_zz_2133_)begin
        int_reg_array_38_39_real <= _zz_2145_;
      end
      if(_zz_2134_)begin
        int_reg_array_38_40_real <= _zz_2145_;
      end
      if(_zz_2135_)begin
        int_reg_array_38_41_real <= _zz_2145_;
      end
      if(_zz_2136_)begin
        int_reg_array_38_42_real <= _zz_2145_;
      end
      if(_zz_2137_)begin
        int_reg_array_38_43_real <= _zz_2145_;
      end
      if(_zz_2138_)begin
        int_reg_array_38_44_real <= _zz_2145_;
      end
      if(_zz_2139_)begin
        int_reg_array_38_45_real <= _zz_2145_;
      end
      if(_zz_2140_)begin
        int_reg_array_38_46_real <= _zz_2145_;
      end
      if(_zz_2141_)begin
        int_reg_array_38_47_real <= _zz_2145_;
      end
      if(_zz_2142_)begin
        int_reg_array_38_48_real <= _zz_2145_;
      end
      if(_zz_2143_)begin
        int_reg_array_38_49_real <= _zz_2145_;
      end
      if(_zz_2094_)begin
        int_reg_array_38_0_imag <= _zz_2146_;
      end
      if(_zz_2095_)begin
        int_reg_array_38_1_imag <= _zz_2146_;
      end
      if(_zz_2096_)begin
        int_reg_array_38_2_imag <= _zz_2146_;
      end
      if(_zz_2097_)begin
        int_reg_array_38_3_imag <= _zz_2146_;
      end
      if(_zz_2098_)begin
        int_reg_array_38_4_imag <= _zz_2146_;
      end
      if(_zz_2099_)begin
        int_reg_array_38_5_imag <= _zz_2146_;
      end
      if(_zz_2100_)begin
        int_reg_array_38_6_imag <= _zz_2146_;
      end
      if(_zz_2101_)begin
        int_reg_array_38_7_imag <= _zz_2146_;
      end
      if(_zz_2102_)begin
        int_reg_array_38_8_imag <= _zz_2146_;
      end
      if(_zz_2103_)begin
        int_reg_array_38_9_imag <= _zz_2146_;
      end
      if(_zz_2104_)begin
        int_reg_array_38_10_imag <= _zz_2146_;
      end
      if(_zz_2105_)begin
        int_reg_array_38_11_imag <= _zz_2146_;
      end
      if(_zz_2106_)begin
        int_reg_array_38_12_imag <= _zz_2146_;
      end
      if(_zz_2107_)begin
        int_reg_array_38_13_imag <= _zz_2146_;
      end
      if(_zz_2108_)begin
        int_reg_array_38_14_imag <= _zz_2146_;
      end
      if(_zz_2109_)begin
        int_reg_array_38_15_imag <= _zz_2146_;
      end
      if(_zz_2110_)begin
        int_reg_array_38_16_imag <= _zz_2146_;
      end
      if(_zz_2111_)begin
        int_reg_array_38_17_imag <= _zz_2146_;
      end
      if(_zz_2112_)begin
        int_reg_array_38_18_imag <= _zz_2146_;
      end
      if(_zz_2113_)begin
        int_reg_array_38_19_imag <= _zz_2146_;
      end
      if(_zz_2114_)begin
        int_reg_array_38_20_imag <= _zz_2146_;
      end
      if(_zz_2115_)begin
        int_reg_array_38_21_imag <= _zz_2146_;
      end
      if(_zz_2116_)begin
        int_reg_array_38_22_imag <= _zz_2146_;
      end
      if(_zz_2117_)begin
        int_reg_array_38_23_imag <= _zz_2146_;
      end
      if(_zz_2118_)begin
        int_reg_array_38_24_imag <= _zz_2146_;
      end
      if(_zz_2119_)begin
        int_reg_array_38_25_imag <= _zz_2146_;
      end
      if(_zz_2120_)begin
        int_reg_array_38_26_imag <= _zz_2146_;
      end
      if(_zz_2121_)begin
        int_reg_array_38_27_imag <= _zz_2146_;
      end
      if(_zz_2122_)begin
        int_reg_array_38_28_imag <= _zz_2146_;
      end
      if(_zz_2123_)begin
        int_reg_array_38_29_imag <= _zz_2146_;
      end
      if(_zz_2124_)begin
        int_reg_array_38_30_imag <= _zz_2146_;
      end
      if(_zz_2125_)begin
        int_reg_array_38_31_imag <= _zz_2146_;
      end
      if(_zz_2126_)begin
        int_reg_array_38_32_imag <= _zz_2146_;
      end
      if(_zz_2127_)begin
        int_reg_array_38_33_imag <= _zz_2146_;
      end
      if(_zz_2128_)begin
        int_reg_array_38_34_imag <= _zz_2146_;
      end
      if(_zz_2129_)begin
        int_reg_array_38_35_imag <= _zz_2146_;
      end
      if(_zz_2130_)begin
        int_reg_array_38_36_imag <= _zz_2146_;
      end
      if(_zz_2131_)begin
        int_reg_array_38_37_imag <= _zz_2146_;
      end
      if(_zz_2132_)begin
        int_reg_array_38_38_imag <= _zz_2146_;
      end
      if(_zz_2133_)begin
        int_reg_array_38_39_imag <= _zz_2146_;
      end
      if(_zz_2134_)begin
        int_reg_array_38_40_imag <= _zz_2146_;
      end
      if(_zz_2135_)begin
        int_reg_array_38_41_imag <= _zz_2146_;
      end
      if(_zz_2136_)begin
        int_reg_array_38_42_imag <= _zz_2146_;
      end
      if(_zz_2137_)begin
        int_reg_array_38_43_imag <= _zz_2146_;
      end
      if(_zz_2138_)begin
        int_reg_array_38_44_imag <= _zz_2146_;
      end
      if(_zz_2139_)begin
        int_reg_array_38_45_imag <= _zz_2146_;
      end
      if(_zz_2140_)begin
        int_reg_array_38_46_imag <= _zz_2146_;
      end
      if(_zz_2141_)begin
        int_reg_array_38_47_imag <= _zz_2146_;
      end
      if(_zz_2142_)begin
        int_reg_array_38_48_imag <= _zz_2146_;
      end
      if(_zz_2143_)begin
        int_reg_array_38_49_imag <= _zz_2146_;
      end
      if(_zz_2149_)begin
        int_reg_array_39_0_real <= _zz_2200_;
      end
      if(_zz_2150_)begin
        int_reg_array_39_1_real <= _zz_2200_;
      end
      if(_zz_2151_)begin
        int_reg_array_39_2_real <= _zz_2200_;
      end
      if(_zz_2152_)begin
        int_reg_array_39_3_real <= _zz_2200_;
      end
      if(_zz_2153_)begin
        int_reg_array_39_4_real <= _zz_2200_;
      end
      if(_zz_2154_)begin
        int_reg_array_39_5_real <= _zz_2200_;
      end
      if(_zz_2155_)begin
        int_reg_array_39_6_real <= _zz_2200_;
      end
      if(_zz_2156_)begin
        int_reg_array_39_7_real <= _zz_2200_;
      end
      if(_zz_2157_)begin
        int_reg_array_39_8_real <= _zz_2200_;
      end
      if(_zz_2158_)begin
        int_reg_array_39_9_real <= _zz_2200_;
      end
      if(_zz_2159_)begin
        int_reg_array_39_10_real <= _zz_2200_;
      end
      if(_zz_2160_)begin
        int_reg_array_39_11_real <= _zz_2200_;
      end
      if(_zz_2161_)begin
        int_reg_array_39_12_real <= _zz_2200_;
      end
      if(_zz_2162_)begin
        int_reg_array_39_13_real <= _zz_2200_;
      end
      if(_zz_2163_)begin
        int_reg_array_39_14_real <= _zz_2200_;
      end
      if(_zz_2164_)begin
        int_reg_array_39_15_real <= _zz_2200_;
      end
      if(_zz_2165_)begin
        int_reg_array_39_16_real <= _zz_2200_;
      end
      if(_zz_2166_)begin
        int_reg_array_39_17_real <= _zz_2200_;
      end
      if(_zz_2167_)begin
        int_reg_array_39_18_real <= _zz_2200_;
      end
      if(_zz_2168_)begin
        int_reg_array_39_19_real <= _zz_2200_;
      end
      if(_zz_2169_)begin
        int_reg_array_39_20_real <= _zz_2200_;
      end
      if(_zz_2170_)begin
        int_reg_array_39_21_real <= _zz_2200_;
      end
      if(_zz_2171_)begin
        int_reg_array_39_22_real <= _zz_2200_;
      end
      if(_zz_2172_)begin
        int_reg_array_39_23_real <= _zz_2200_;
      end
      if(_zz_2173_)begin
        int_reg_array_39_24_real <= _zz_2200_;
      end
      if(_zz_2174_)begin
        int_reg_array_39_25_real <= _zz_2200_;
      end
      if(_zz_2175_)begin
        int_reg_array_39_26_real <= _zz_2200_;
      end
      if(_zz_2176_)begin
        int_reg_array_39_27_real <= _zz_2200_;
      end
      if(_zz_2177_)begin
        int_reg_array_39_28_real <= _zz_2200_;
      end
      if(_zz_2178_)begin
        int_reg_array_39_29_real <= _zz_2200_;
      end
      if(_zz_2179_)begin
        int_reg_array_39_30_real <= _zz_2200_;
      end
      if(_zz_2180_)begin
        int_reg_array_39_31_real <= _zz_2200_;
      end
      if(_zz_2181_)begin
        int_reg_array_39_32_real <= _zz_2200_;
      end
      if(_zz_2182_)begin
        int_reg_array_39_33_real <= _zz_2200_;
      end
      if(_zz_2183_)begin
        int_reg_array_39_34_real <= _zz_2200_;
      end
      if(_zz_2184_)begin
        int_reg_array_39_35_real <= _zz_2200_;
      end
      if(_zz_2185_)begin
        int_reg_array_39_36_real <= _zz_2200_;
      end
      if(_zz_2186_)begin
        int_reg_array_39_37_real <= _zz_2200_;
      end
      if(_zz_2187_)begin
        int_reg_array_39_38_real <= _zz_2200_;
      end
      if(_zz_2188_)begin
        int_reg_array_39_39_real <= _zz_2200_;
      end
      if(_zz_2189_)begin
        int_reg_array_39_40_real <= _zz_2200_;
      end
      if(_zz_2190_)begin
        int_reg_array_39_41_real <= _zz_2200_;
      end
      if(_zz_2191_)begin
        int_reg_array_39_42_real <= _zz_2200_;
      end
      if(_zz_2192_)begin
        int_reg_array_39_43_real <= _zz_2200_;
      end
      if(_zz_2193_)begin
        int_reg_array_39_44_real <= _zz_2200_;
      end
      if(_zz_2194_)begin
        int_reg_array_39_45_real <= _zz_2200_;
      end
      if(_zz_2195_)begin
        int_reg_array_39_46_real <= _zz_2200_;
      end
      if(_zz_2196_)begin
        int_reg_array_39_47_real <= _zz_2200_;
      end
      if(_zz_2197_)begin
        int_reg_array_39_48_real <= _zz_2200_;
      end
      if(_zz_2198_)begin
        int_reg_array_39_49_real <= _zz_2200_;
      end
      if(_zz_2149_)begin
        int_reg_array_39_0_imag <= _zz_2201_;
      end
      if(_zz_2150_)begin
        int_reg_array_39_1_imag <= _zz_2201_;
      end
      if(_zz_2151_)begin
        int_reg_array_39_2_imag <= _zz_2201_;
      end
      if(_zz_2152_)begin
        int_reg_array_39_3_imag <= _zz_2201_;
      end
      if(_zz_2153_)begin
        int_reg_array_39_4_imag <= _zz_2201_;
      end
      if(_zz_2154_)begin
        int_reg_array_39_5_imag <= _zz_2201_;
      end
      if(_zz_2155_)begin
        int_reg_array_39_6_imag <= _zz_2201_;
      end
      if(_zz_2156_)begin
        int_reg_array_39_7_imag <= _zz_2201_;
      end
      if(_zz_2157_)begin
        int_reg_array_39_8_imag <= _zz_2201_;
      end
      if(_zz_2158_)begin
        int_reg_array_39_9_imag <= _zz_2201_;
      end
      if(_zz_2159_)begin
        int_reg_array_39_10_imag <= _zz_2201_;
      end
      if(_zz_2160_)begin
        int_reg_array_39_11_imag <= _zz_2201_;
      end
      if(_zz_2161_)begin
        int_reg_array_39_12_imag <= _zz_2201_;
      end
      if(_zz_2162_)begin
        int_reg_array_39_13_imag <= _zz_2201_;
      end
      if(_zz_2163_)begin
        int_reg_array_39_14_imag <= _zz_2201_;
      end
      if(_zz_2164_)begin
        int_reg_array_39_15_imag <= _zz_2201_;
      end
      if(_zz_2165_)begin
        int_reg_array_39_16_imag <= _zz_2201_;
      end
      if(_zz_2166_)begin
        int_reg_array_39_17_imag <= _zz_2201_;
      end
      if(_zz_2167_)begin
        int_reg_array_39_18_imag <= _zz_2201_;
      end
      if(_zz_2168_)begin
        int_reg_array_39_19_imag <= _zz_2201_;
      end
      if(_zz_2169_)begin
        int_reg_array_39_20_imag <= _zz_2201_;
      end
      if(_zz_2170_)begin
        int_reg_array_39_21_imag <= _zz_2201_;
      end
      if(_zz_2171_)begin
        int_reg_array_39_22_imag <= _zz_2201_;
      end
      if(_zz_2172_)begin
        int_reg_array_39_23_imag <= _zz_2201_;
      end
      if(_zz_2173_)begin
        int_reg_array_39_24_imag <= _zz_2201_;
      end
      if(_zz_2174_)begin
        int_reg_array_39_25_imag <= _zz_2201_;
      end
      if(_zz_2175_)begin
        int_reg_array_39_26_imag <= _zz_2201_;
      end
      if(_zz_2176_)begin
        int_reg_array_39_27_imag <= _zz_2201_;
      end
      if(_zz_2177_)begin
        int_reg_array_39_28_imag <= _zz_2201_;
      end
      if(_zz_2178_)begin
        int_reg_array_39_29_imag <= _zz_2201_;
      end
      if(_zz_2179_)begin
        int_reg_array_39_30_imag <= _zz_2201_;
      end
      if(_zz_2180_)begin
        int_reg_array_39_31_imag <= _zz_2201_;
      end
      if(_zz_2181_)begin
        int_reg_array_39_32_imag <= _zz_2201_;
      end
      if(_zz_2182_)begin
        int_reg_array_39_33_imag <= _zz_2201_;
      end
      if(_zz_2183_)begin
        int_reg_array_39_34_imag <= _zz_2201_;
      end
      if(_zz_2184_)begin
        int_reg_array_39_35_imag <= _zz_2201_;
      end
      if(_zz_2185_)begin
        int_reg_array_39_36_imag <= _zz_2201_;
      end
      if(_zz_2186_)begin
        int_reg_array_39_37_imag <= _zz_2201_;
      end
      if(_zz_2187_)begin
        int_reg_array_39_38_imag <= _zz_2201_;
      end
      if(_zz_2188_)begin
        int_reg_array_39_39_imag <= _zz_2201_;
      end
      if(_zz_2189_)begin
        int_reg_array_39_40_imag <= _zz_2201_;
      end
      if(_zz_2190_)begin
        int_reg_array_39_41_imag <= _zz_2201_;
      end
      if(_zz_2191_)begin
        int_reg_array_39_42_imag <= _zz_2201_;
      end
      if(_zz_2192_)begin
        int_reg_array_39_43_imag <= _zz_2201_;
      end
      if(_zz_2193_)begin
        int_reg_array_39_44_imag <= _zz_2201_;
      end
      if(_zz_2194_)begin
        int_reg_array_39_45_imag <= _zz_2201_;
      end
      if(_zz_2195_)begin
        int_reg_array_39_46_imag <= _zz_2201_;
      end
      if(_zz_2196_)begin
        int_reg_array_39_47_imag <= _zz_2201_;
      end
      if(_zz_2197_)begin
        int_reg_array_39_48_imag <= _zz_2201_;
      end
      if(_zz_2198_)begin
        int_reg_array_39_49_imag <= _zz_2201_;
      end
      if(_zz_2204_)begin
        int_reg_array_40_0_real <= _zz_2255_;
      end
      if(_zz_2205_)begin
        int_reg_array_40_1_real <= _zz_2255_;
      end
      if(_zz_2206_)begin
        int_reg_array_40_2_real <= _zz_2255_;
      end
      if(_zz_2207_)begin
        int_reg_array_40_3_real <= _zz_2255_;
      end
      if(_zz_2208_)begin
        int_reg_array_40_4_real <= _zz_2255_;
      end
      if(_zz_2209_)begin
        int_reg_array_40_5_real <= _zz_2255_;
      end
      if(_zz_2210_)begin
        int_reg_array_40_6_real <= _zz_2255_;
      end
      if(_zz_2211_)begin
        int_reg_array_40_7_real <= _zz_2255_;
      end
      if(_zz_2212_)begin
        int_reg_array_40_8_real <= _zz_2255_;
      end
      if(_zz_2213_)begin
        int_reg_array_40_9_real <= _zz_2255_;
      end
      if(_zz_2214_)begin
        int_reg_array_40_10_real <= _zz_2255_;
      end
      if(_zz_2215_)begin
        int_reg_array_40_11_real <= _zz_2255_;
      end
      if(_zz_2216_)begin
        int_reg_array_40_12_real <= _zz_2255_;
      end
      if(_zz_2217_)begin
        int_reg_array_40_13_real <= _zz_2255_;
      end
      if(_zz_2218_)begin
        int_reg_array_40_14_real <= _zz_2255_;
      end
      if(_zz_2219_)begin
        int_reg_array_40_15_real <= _zz_2255_;
      end
      if(_zz_2220_)begin
        int_reg_array_40_16_real <= _zz_2255_;
      end
      if(_zz_2221_)begin
        int_reg_array_40_17_real <= _zz_2255_;
      end
      if(_zz_2222_)begin
        int_reg_array_40_18_real <= _zz_2255_;
      end
      if(_zz_2223_)begin
        int_reg_array_40_19_real <= _zz_2255_;
      end
      if(_zz_2224_)begin
        int_reg_array_40_20_real <= _zz_2255_;
      end
      if(_zz_2225_)begin
        int_reg_array_40_21_real <= _zz_2255_;
      end
      if(_zz_2226_)begin
        int_reg_array_40_22_real <= _zz_2255_;
      end
      if(_zz_2227_)begin
        int_reg_array_40_23_real <= _zz_2255_;
      end
      if(_zz_2228_)begin
        int_reg_array_40_24_real <= _zz_2255_;
      end
      if(_zz_2229_)begin
        int_reg_array_40_25_real <= _zz_2255_;
      end
      if(_zz_2230_)begin
        int_reg_array_40_26_real <= _zz_2255_;
      end
      if(_zz_2231_)begin
        int_reg_array_40_27_real <= _zz_2255_;
      end
      if(_zz_2232_)begin
        int_reg_array_40_28_real <= _zz_2255_;
      end
      if(_zz_2233_)begin
        int_reg_array_40_29_real <= _zz_2255_;
      end
      if(_zz_2234_)begin
        int_reg_array_40_30_real <= _zz_2255_;
      end
      if(_zz_2235_)begin
        int_reg_array_40_31_real <= _zz_2255_;
      end
      if(_zz_2236_)begin
        int_reg_array_40_32_real <= _zz_2255_;
      end
      if(_zz_2237_)begin
        int_reg_array_40_33_real <= _zz_2255_;
      end
      if(_zz_2238_)begin
        int_reg_array_40_34_real <= _zz_2255_;
      end
      if(_zz_2239_)begin
        int_reg_array_40_35_real <= _zz_2255_;
      end
      if(_zz_2240_)begin
        int_reg_array_40_36_real <= _zz_2255_;
      end
      if(_zz_2241_)begin
        int_reg_array_40_37_real <= _zz_2255_;
      end
      if(_zz_2242_)begin
        int_reg_array_40_38_real <= _zz_2255_;
      end
      if(_zz_2243_)begin
        int_reg_array_40_39_real <= _zz_2255_;
      end
      if(_zz_2244_)begin
        int_reg_array_40_40_real <= _zz_2255_;
      end
      if(_zz_2245_)begin
        int_reg_array_40_41_real <= _zz_2255_;
      end
      if(_zz_2246_)begin
        int_reg_array_40_42_real <= _zz_2255_;
      end
      if(_zz_2247_)begin
        int_reg_array_40_43_real <= _zz_2255_;
      end
      if(_zz_2248_)begin
        int_reg_array_40_44_real <= _zz_2255_;
      end
      if(_zz_2249_)begin
        int_reg_array_40_45_real <= _zz_2255_;
      end
      if(_zz_2250_)begin
        int_reg_array_40_46_real <= _zz_2255_;
      end
      if(_zz_2251_)begin
        int_reg_array_40_47_real <= _zz_2255_;
      end
      if(_zz_2252_)begin
        int_reg_array_40_48_real <= _zz_2255_;
      end
      if(_zz_2253_)begin
        int_reg_array_40_49_real <= _zz_2255_;
      end
      if(_zz_2204_)begin
        int_reg_array_40_0_imag <= _zz_2256_;
      end
      if(_zz_2205_)begin
        int_reg_array_40_1_imag <= _zz_2256_;
      end
      if(_zz_2206_)begin
        int_reg_array_40_2_imag <= _zz_2256_;
      end
      if(_zz_2207_)begin
        int_reg_array_40_3_imag <= _zz_2256_;
      end
      if(_zz_2208_)begin
        int_reg_array_40_4_imag <= _zz_2256_;
      end
      if(_zz_2209_)begin
        int_reg_array_40_5_imag <= _zz_2256_;
      end
      if(_zz_2210_)begin
        int_reg_array_40_6_imag <= _zz_2256_;
      end
      if(_zz_2211_)begin
        int_reg_array_40_7_imag <= _zz_2256_;
      end
      if(_zz_2212_)begin
        int_reg_array_40_8_imag <= _zz_2256_;
      end
      if(_zz_2213_)begin
        int_reg_array_40_9_imag <= _zz_2256_;
      end
      if(_zz_2214_)begin
        int_reg_array_40_10_imag <= _zz_2256_;
      end
      if(_zz_2215_)begin
        int_reg_array_40_11_imag <= _zz_2256_;
      end
      if(_zz_2216_)begin
        int_reg_array_40_12_imag <= _zz_2256_;
      end
      if(_zz_2217_)begin
        int_reg_array_40_13_imag <= _zz_2256_;
      end
      if(_zz_2218_)begin
        int_reg_array_40_14_imag <= _zz_2256_;
      end
      if(_zz_2219_)begin
        int_reg_array_40_15_imag <= _zz_2256_;
      end
      if(_zz_2220_)begin
        int_reg_array_40_16_imag <= _zz_2256_;
      end
      if(_zz_2221_)begin
        int_reg_array_40_17_imag <= _zz_2256_;
      end
      if(_zz_2222_)begin
        int_reg_array_40_18_imag <= _zz_2256_;
      end
      if(_zz_2223_)begin
        int_reg_array_40_19_imag <= _zz_2256_;
      end
      if(_zz_2224_)begin
        int_reg_array_40_20_imag <= _zz_2256_;
      end
      if(_zz_2225_)begin
        int_reg_array_40_21_imag <= _zz_2256_;
      end
      if(_zz_2226_)begin
        int_reg_array_40_22_imag <= _zz_2256_;
      end
      if(_zz_2227_)begin
        int_reg_array_40_23_imag <= _zz_2256_;
      end
      if(_zz_2228_)begin
        int_reg_array_40_24_imag <= _zz_2256_;
      end
      if(_zz_2229_)begin
        int_reg_array_40_25_imag <= _zz_2256_;
      end
      if(_zz_2230_)begin
        int_reg_array_40_26_imag <= _zz_2256_;
      end
      if(_zz_2231_)begin
        int_reg_array_40_27_imag <= _zz_2256_;
      end
      if(_zz_2232_)begin
        int_reg_array_40_28_imag <= _zz_2256_;
      end
      if(_zz_2233_)begin
        int_reg_array_40_29_imag <= _zz_2256_;
      end
      if(_zz_2234_)begin
        int_reg_array_40_30_imag <= _zz_2256_;
      end
      if(_zz_2235_)begin
        int_reg_array_40_31_imag <= _zz_2256_;
      end
      if(_zz_2236_)begin
        int_reg_array_40_32_imag <= _zz_2256_;
      end
      if(_zz_2237_)begin
        int_reg_array_40_33_imag <= _zz_2256_;
      end
      if(_zz_2238_)begin
        int_reg_array_40_34_imag <= _zz_2256_;
      end
      if(_zz_2239_)begin
        int_reg_array_40_35_imag <= _zz_2256_;
      end
      if(_zz_2240_)begin
        int_reg_array_40_36_imag <= _zz_2256_;
      end
      if(_zz_2241_)begin
        int_reg_array_40_37_imag <= _zz_2256_;
      end
      if(_zz_2242_)begin
        int_reg_array_40_38_imag <= _zz_2256_;
      end
      if(_zz_2243_)begin
        int_reg_array_40_39_imag <= _zz_2256_;
      end
      if(_zz_2244_)begin
        int_reg_array_40_40_imag <= _zz_2256_;
      end
      if(_zz_2245_)begin
        int_reg_array_40_41_imag <= _zz_2256_;
      end
      if(_zz_2246_)begin
        int_reg_array_40_42_imag <= _zz_2256_;
      end
      if(_zz_2247_)begin
        int_reg_array_40_43_imag <= _zz_2256_;
      end
      if(_zz_2248_)begin
        int_reg_array_40_44_imag <= _zz_2256_;
      end
      if(_zz_2249_)begin
        int_reg_array_40_45_imag <= _zz_2256_;
      end
      if(_zz_2250_)begin
        int_reg_array_40_46_imag <= _zz_2256_;
      end
      if(_zz_2251_)begin
        int_reg_array_40_47_imag <= _zz_2256_;
      end
      if(_zz_2252_)begin
        int_reg_array_40_48_imag <= _zz_2256_;
      end
      if(_zz_2253_)begin
        int_reg_array_40_49_imag <= _zz_2256_;
      end
      if(_zz_2259_)begin
        int_reg_array_41_0_real <= _zz_2310_;
      end
      if(_zz_2260_)begin
        int_reg_array_41_1_real <= _zz_2310_;
      end
      if(_zz_2261_)begin
        int_reg_array_41_2_real <= _zz_2310_;
      end
      if(_zz_2262_)begin
        int_reg_array_41_3_real <= _zz_2310_;
      end
      if(_zz_2263_)begin
        int_reg_array_41_4_real <= _zz_2310_;
      end
      if(_zz_2264_)begin
        int_reg_array_41_5_real <= _zz_2310_;
      end
      if(_zz_2265_)begin
        int_reg_array_41_6_real <= _zz_2310_;
      end
      if(_zz_2266_)begin
        int_reg_array_41_7_real <= _zz_2310_;
      end
      if(_zz_2267_)begin
        int_reg_array_41_8_real <= _zz_2310_;
      end
      if(_zz_2268_)begin
        int_reg_array_41_9_real <= _zz_2310_;
      end
      if(_zz_2269_)begin
        int_reg_array_41_10_real <= _zz_2310_;
      end
      if(_zz_2270_)begin
        int_reg_array_41_11_real <= _zz_2310_;
      end
      if(_zz_2271_)begin
        int_reg_array_41_12_real <= _zz_2310_;
      end
      if(_zz_2272_)begin
        int_reg_array_41_13_real <= _zz_2310_;
      end
      if(_zz_2273_)begin
        int_reg_array_41_14_real <= _zz_2310_;
      end
      if(_zz_2274_)begin
        int_reg_array_41_15_real <= _zz_2310_;
      end
      if(_zz_2275_)begin
        int_reg_array_41_16_real <= _zz_2310_;
      end
      if(_zz_2276_)begin
        int_reg_array_41_17_real <= _zz_2310_;
      end
      if(_zz_2277_)begin
        int_reg_array_41_18_real <= _zz_2310_;
      end
      if(_zz_2278_)begin
        int_reg_array_41_19_real <= _zz_2310_;
      end
      if(_zz_2279_)begin
        int_reg_array_41_20_real <= _zz_2310_;
      end
      if(_zz_2280_)begin
        int_reg_array_41_21_real <= _zz_2310_;
      end
      if(_zz_2281_)begin
        int_reg_array_41_22_real <= _zz_2310_;
      end
      if(_zz_2282_)begin
        int_reg_array_41_23_real <= _zz_2310_;
      end
      if(_zz_2283_)begin
        int_reg_array_41_24_real <= _zz_2310_;
      end
      if(_zz_2284_)begin
        int_reg_array_41_25_real <= _zz_2310_;
      end
      if(_zz_2285_)begin
        int_reg_array_41_26_real <= _zz_2310_;
      end
      if(_zz_2286_)begin
        int_reg_array_41_27_real <= _zz_2310_;
      end
      if(_zz_2287_)begin
        int_reg_array_41_28_real <= _zz_2310_;
      end
      if(_zz_2288_)begin
        int_reg_array_41_29_real <= _zz_2310_;
      end
      if(_zz_2289_)begin
        int_reg_array_41_30_real <= _zz_2310_;
      end
      if(_zz_2290_)begin
        int_reg_array_41_31_real <= _zz_2310_;
      end
      if(_zz_2291_)begin
        int_reg_array_41_32_real <= _zz_2310_;
      end
      if(_zz_2292_)begin
        int_reg_array_41_33_real <= _zz_2310_;
      end
      if(_zz_2293_)begin
        int_reg_array_41_34_real <= _zz_2310_;
      end
      if(_zz_2294_)begin
        int_reg_array_41_35_real <= _zz_2310_;
      end
      if(_zz_2295_)begin
        int_reg_array_41_36_real <= _zz_2310_;
      end
      if(_zz_2296_)begin
        int_reg_array_41_37_real <= _zz_2310_;
      end
      if(_zz_2297_)begin
        int_reg_array_41_38_real <= _zz_2310_;
      end
      if(_zz_2298_)begin
        int_reg_array_41_39_real <= _zz_2310_;
      end
      if(_zz_2299_)begin
        int_reg_array_41_40_real <= _zz_2310_;
      end
      if(_zz_2300_)begin
        int_reg_array_41_41_real <= _zz_2310_;
      end
      if(_zz_2301_)begin
        int_reg_array_41_42_real <= _zz_2310_;
      end
      if(_zz_2302_)begin
        int_reg_array_41_43_real <= _zz_2310_;
      end
      if(_zz_2303_)begin
        int_reg_array_41_44_real <= _zz_2310_;
      end
      if(_zz_2304_)begin
        int_reg_array_41_45_real <= _zz_2310_;
      end
      if(_zz_2305_)begin
        int_reg_array_41_46_real <= _zz_2310_;
      end
      if(_zz_2306_)begin
        int_reg_array_41_47_real <= _zz_2310_;
      end
      if(_zz_2307_)begin
        int_reg_array_41_48_real <= _zz_2310_;
      end
      if(_zz_2308_)begin
        int_reg_array_41_49_real <= _zz_2310_;
      end
      if(_zz_2259_)begin
        int_reg_array_41_0_imag <= _zz_2311_;
      end
      if(_zz_2260_)begin
        int_reg_array_41_1_imag <= _zz_2311_;
      end
      if(_zz_2261_)begin
        int_reg_array_41_2_imag <= _zz_2311_;
      end
      if(_zz_2262_)begin
        int_reg_array_41_3_imag <= _zz_2311_;
      end
      if(_zz_2263_)begin
        int_reg_array_41_4_imag <= _zz_2311_;
      end
      if(_zz_2264_)begin
        int_reg_array_41_5_imag <= _zz_2311_;
      end
      if(_zz_2265_)begin
        int_reg_array_41_6_imag <= _zz_2311_;
      end
      if(_zz_2266_)begin
        int_reg_array_41_7_imag <= _zz_2311_;
      end
      if(_zz_2267_)begin
        int_reg_array_41_8_imag <= _zz_2311_;
      end
      if(_zz_2268_)begin
        int_reg_array_41_9_imag <= _zz_2311_;
      end
      if(_zz_2269_)begin
        int_reg_array_41_10_imag <= _zz_2311_;
      end
      if(_zz_2270_)begin
        int_reg_array_41_11_imag <= _zz_2311_;
      end
      if(_zz_2271_)begin
        int_reg_array_41_12_imag <= _zz_2311_;
      end
      if(_zz_2272_)begin
        int_reg_array_41_13_imag <= _zz_2311_;
      end
      if(_zz_2273_)begin
        int_reg_array_41_14_imag <= _zz_2311_;
      end
      if(_zz_2274_)begin
        int_reg_array_41_15_imag <= _zz_2311_;
      end
      if(_zz_2275_)begin
        int_reg_array_41_16_imag <= _zz_2311_;
      end
      if(_zz_2276_)begin
        int_reg_array_41_17_imag <= _zz_2311_;
      end
      if(_zz_2277_)begin
        int_reg_array_41_18_imag <= _zz_2311_;
      end
      if(_zz_2278_)begin
        int_reg_array_41_19_imag <= _zz_2311_;
      end
      if(_zz_2279_)begin
        int_reg_array_41_20_imag <= _zz_2311_;
      end
      if(_zz_2280_)begin
        int_reg_array_41_21_imag <= _zz_2311_;
      end
      if(_zz_2281_)begin
        int_reg_array_41_22_imag <= _zz_2311_;
      end
      if(_zz_2282_)begin
        int_reg_array_41_23_imag <= _zz_2311_;
      end
      if(_zz_2283_)begin
        int_reg_array_41_24_imag <= _zz_2311_;
      end
      if(_zz_2284_)begin
        int_reg_array_41_25_imag <= _zz_2311_;
      end
      if(_zz_2285_)begin
        int_reg_array_41_26_imag <= _zz_2311_;
      end
      if(_zz_2286_)begin
        int_reg_array_41_27_imag <= _zz_2311_;
      end
      if(_zz_2287_)begin
        int_reg_array_41_28_imag <= _zz_2311_;
      end
      if(_zz_2288_)begin
        int_reg_array_41_29_imag <= _zz_2311_;
      end
      if(_zz_2289_)begin
        int_reg_array_41_30_imag <= _zz_2311_;
      end
      if(_zz_2290_)begin
        int_reg_array_41_31_imag <= _zz_2311_;
      end
      if(_zz_2291_)begin
        int_reg_array_41_32_imag <= _zz_2311_;
      end
      if(_zz_2292_)begin
        int_reg_array_41_33_imag <= _zz_2311_;
      end
      if(_zz_2293_)begin
        int_reg_array_41_34_imag <= _zz_2311_;
      end
      if(_zz_2294_)begin
        int_reg_array_41_35_imag <= _zz_2311_;
      end
      if(_zz_2295_)begin
        int_reg_array_41_36_imag <= _zz_2311_;
      end
      if(_zz_2296_)begin
        int_reg_array_41_37_imag <= _zz_2311_;
      end
      if(_zz_2297_)begin
        int_reg_array_41_38_imag <= _zz_2311_;
      end
      if(_zz_2298_)begin
        int_reg_array_41_39_imag <= _zz_2311_;
      end
      if(_zz_2299_)begin
        int_reg_array_41_40_imag <= _zz_2311_;
      end
      if(_zz_2300_)begin
        int_reg_array_41_41_imag <= _zz_2311_;
      end
      if(_zz_2301_)begin
        int_reg_array_41_42_imag <= _zz_2311_;
      end
      if(_zz_2302_)begin
        int_reg_array_41_43_imag <= _zz_2311_;
      end
      if(_zz_2303_)begin
        int_reg_array_41_44_imag <= _zz_2311_;
      end
      if(_zz_2304_)begin
        int_reg_array_41_45_imag <= _zz_2311_;
      end
      if(_zz_2305_)begin
        int_reg_array_41_46_imag <= _zz_2311_;
      end
      if(_zz_2306_)begin
        int_reg_array_41_47_imag <= _zz_2311_;
      end
      if(_zz_2307_)begin
        int_reg_array_41_48_imag <= _zz_2311_;
      end
      if(_zz_2308_)begin
        int_reg_array_41_49_imag <= _zz_2311_;
      end
      if(_zz_2314_)begin
        int_reg_array_42_0_real <= _zz_2365_;
      end
      if(_zz_2315_)begin
        int_reg_array_42_1_real <= _zz_2365_;
      end
      if(_zz_2316_)begin
        int_reg_array_42_2_real <= _zz_2365_;
      end
      if(_zz_2317_)begin
        int_reg_array_42_3_real <= _zz_2365_;
      end
      if(_zz_2318_)begin
        int_reg_array_42_4_real <= _zz_2365_;
      end
      if(_zz_2319_)begin
        int_reg_array_42_5_real <= _zz_2365_;
      end
      if(_zz_2320_)begin
        int_reg_array_42_6_real <= _zz_2365_;
      end
      if(_zz_2321_)begin
        int_reg_array_42_7_real <= _zz_2365_;
      end
      if(_zz_2322_)begin
        int_reg_array_42_8_real <= _zz_2365_;
      end
      if(_zz_2323_)begin
        int_reg_array_42_9_real <= _zz_2365_;
      end
      if(_zz_2324_)begin
        int_reg_array_42_10_real <= _zz_2365_;
      end
      if(_zz_2325_)begin
        int_reg_array_42_11_real <= _zz_2365_;
      end
      if(_zz_2326_)begin
        int_reg_array_42_12_real <= _zz_2365_;
      end
      if(_zz_2327_)begin
        int_reg_array_42_13_real <= _zz_2365_;
      end
      if(_zz_2328_)begin
        int_reg_array_42_14_real <= _zz_2365_;
      end
      if(_zz_2329_)begin
        int_reg_array_42_15_real <= _zz_2365_;
      end
      if(_zz_2330_)begin
        int_reg_array_42_16_real <= _zz_2365_;
      end
      if(_zz_2331_)begin
        int_reg_array_42_17_real <= _zz_2365_;
      end
      if(_zz_2332_)begin
        int_reg_array_42_18_real <= _zz_2365_;
      end
      if(_zz_2333_)begin
        int_reg_array_42_19_real <= _zz_2365_;
      end
      if(_zz_2334_)begin
        int_reg_array_42_20_real <= _zz_2365_;
      end
      if(_zz_2335_)begin
        int_reg_array_42_21_real <= _zz_2365_;
      end
      if(_zz_2336_)begin
        int_reg_array_42_22_real <= _zz_2365_;
      end
      if(_zz_2337_)begin
        int_reg_array_42_23_real <= _zz_2365_;
      end
      if(_zz_2338_)begin
        int_reg_array_42_24_real <= _zz_2365_;
      end
      if(_zz_2339_)begin
        int_reg_array_42_25_real <= _zz_2365_;
      end
      if(_zz_2340_)begin
        int_reg_array_42_26_real <= _zz_2365_;
      end
      if(_zz_2341_)begin
        int_reg_array_42_27_real <= _zz_2365_;
      end
      if(_zz_2342_)begin
        int_reg_array_42_28_real <= _zz_2365_;
      end
      if(_zz_2343_)begin
        int_reg_array_42_29_real <= _zz_2365_;
      end
      if(_zz_2344_)begin
        int_reg_array_42_30_real <= _zz_2365_;
      end
      if(_zz_2345_)begin
        int_reg_array_42_31_real <= _zz_2365_;
      end
      if(_zz_2346_)begin
        int_reg_array_42_32_real <= _zz_2365_;
      end
      if(_zz_2347_)begin
        int_reg_array_42_33_real <= _zz_2365_;
      end
      if(_zz_2348_)begin
        int_reg_array_42_34_real <= _zz_2365_;
      end
      if(_zz_2349_)begin
        int_reg_array_42_35_real <= _zz_2365_;
      end
      if(_zz_2350_)begin
        int_reg_array_42_36_real <= _zz_2365_;
      end
      if(_zz_2351_)begin
        int_reg_array_42_37_real <= _zz_2365_;
      end
      if(_zz_2352_)begin
        int_reg_array_42_38_real <= _zz_2365_;
      end
      if(_zz_2353_)begin
        int_reg_array_42_39_real <= _zz_2365_;
      end
      if(_zz_2354_)begin
        int_reg_array_42_40_real <= _zz_2365_;
      end
      if(_zz_2355_)begin
        int_reg_array_42_41_real <= _zz_2365_;
      end
      if(_zz_2356_)begin
        int_reg_array_42_42_real <= _zz_2365_;
      end
      if(_zz_2357_)begin
        int_reg_array_42_43_real <= _zz_2365_;
      end
      if(_zz_2358_)begin
        int_reg_array_42_44_real <= _zz_2365_;
      end
      if(_zz_2359_)begin
        int_reg_array_42_45_real <= _zz_2365_;
      end
      if(_zz_2360_)begin
        int_reg_array_42_46_real <= _zz_2365_;
      end
      if(_zz_2361_)begin
        int_reg_array_42_47_real <= _zz_2365_;
      end
      if(_zz_2362_)begin
        int_reg_array_42_48_real <= _zz_2365_;
      end
      if(_zz_2363_)begin
        int_reg_array_42_49_real <= _zz_2365_;
      end
      if(_zz_2314_)begin
        int_reg_array_42_0_imag <= _zz_2366_;
      end
      if(_zz_2315_)begin
        int_reg_array_42_1_imag <= _zz_2366_;
      end
      if(_zz_2316_)begin
        int_reg_array_42_2_imag <= _zz_2366_;
      end
      if(_zz_2317_)begin
        int_reg_array_42_3_imag <= _zz_2366_;
      end
      if(_zz_2318_)begin
        int_reg_array_42_4_imag <= _zz_2366_;
      end
      if(_zz_2319_)begin
        int_reg_array_42_5_imag <= _zz_2366_;
      end
      if(_zz_2320_)begin
        int_reg_array_42_6_imag <= _zz_2366_;
      end
      if(_zz_2321_)begin
        int_reg_array_42_7_imag <= _zz_2366_;
      end
      if(_zz_2322_)begin
        int_reg_array_42_8_imag <= _zz_2366_;
      end
      if(_zz_2323_)begin
        int_reg_array_42_9_imag <= _zz_2366_;
      end
      if(_zz_2324_)begin
        int_reg_array_42_10_imag <= _zz_2366_;
      end
      if(_zz_2325_)begin
        int_reg_array_42_11_imag <= _zz_2366_;
      end
      if(_zz_2326_)begin
        int_reg_array_42_12_imag <= _zz_2366_;
      end
      if(_zz_2327_)begin
        int_reg_array_42_13_imag <= _zz_2366_;
      end
      if(_zz_2328_)begin
        int_reg_array_42_14_imag <= _zz_2366_;
      end
      if(_zz_2329_)begin
        int_reg_array_42_15_imag <= _zz_2366_;
      end
      if(_zz_2330_)begin
        int_reg_array_42_16_imag <= _zz_2366_;
      end
      if(_zz_2331_)begin
        int_reg_array_42_17_imag <= _zz_2366_;
      end
      if(_zz_2332_)begin
        int_reg_array_42_18_imag <= _zz_2366_;
      end
      if(_zz_2333_)begin
        int_reg_array_42_19_imag <= _zz_2366_;
      end
      if(_zz_2334_)begin
        int_reg_array_42_20_imag <= _zz_2366_;
      end
      if(_zz_2335_)begin
        int_reg_array_42_21_imag <= _zz_2366_;
      end
      if(_zz_2336_)begin
        int_reg_array_42_22_imag <= _zz_2366_;
      end
      if(_zz_2337_)begin
        int_reg_array_42_23_imag <= _zz_2366_;
      end
      if(_zz_2338_)begin
        int_reg_array_42_24_imag <= _zz_2366_;
      end
      if(_zz_2339_)begin
        int_reg_array_42_25_imag <= _zz_2366_;
      end
      if(_zz_2340_)begin
        int_reg_array_42_26_imag <= _zz_2366_;
      end
      if(_zz_2341_)begin
        int_reg_array_42_27_imag <= _zz_2366_;
      end
      if(_zz_2342_)begin
        int_reg_array_42_28_imag <= _zz_2366_;
      end
      if(_zz_2343_)begin
        int_reg_array_42_29_imag <= _zz_2366_;
      end
      if(_zz_2344_)begin
        int_reg_array_42_30_imag <= _zz_2366_;
      end
      if(_zz_2345_)begin
        int_reg_array_42_31_imag <= _zz_2366_;
      end
      if(_zz_2346_)begin
        int_reg_array_42_32_imag <= _zz_2366_;
      end
      if(_zz_2347_)begin
        int_reg_array_42_33_imag <= _zz_2366_;
      end
      if(_zz_2348_)begin
        int_reg_array_42_34_imag <= _zz_2366_;
      end
      if(_zz_2349_)begin
        int_reg_array_42_35_imag <= _zz_2366_;
      end
      if(_zz_2350_)begin
        int_reg_array_42_36_imag <= _zz_2366_;
      end
      if(_zz_2351_)begin
        int_reg_array_42_37_imag <= _zz_2366_;
      end
      if(_zz_2352_)begin
        int_reg_array_42_38_imag <= _zz_2366_;
      end
      if(_zz_2353_)begin
        int_reg_array_42_39_imag <= _zz_2366_;
      end
      if(_zz_2354_)begin
        int_reg_array_42_40_imag <= _zz_2366_;
      end
      if(_zz_2355_)begin
        int_reg_array_42_41_imag <= _zz_2366_;
      end
      if(_zz_2356_)begin
        int_reg_array_42_42_imag <= _zz_2366_;
      end
      if(_zz_2357_)begin
        int_reg_array_42_43_imag <= _zz_2366_;
      end
      if(_zz_2358_)begin
        int_reg_array_42_44_imag <= _zz_2366_;
      end
      if(_zz_2359_)begin
        int_reg_array_42_45_imag <= _zz_2366_;
      end
      if(_zz_2360_)begin
        int_reg_array_42_46_imag <= _zz_2366_;
      end
      if(_zz_2361_)begin
        int_reg_array_42_47_imag <= _zz_2366_;
      end
      if(_zz_2362_)begin
        int_reg_array_42_48_imag <= _zz_2366_;
      end
      if(_zz_2363_)begin
        int_reg_array_42_49_imag <= _zz_2366_;
      end
      if(_zz_2369_)begin
        int_reg_array_43_0_real <= _zz_2420_;
      end
      if(_zz_2370_)begin
        int_reg_array_43_1_real <= _zz_2420_;
      end
      if(_zz_2371_)begin
        int_reg_array_43_2_real <= _zz_2420_;
      end
      if(_zz_2372_)begin
        int_reg_array_43_3_real <= _zz_2420_;
      end
      if(_zz_2373_)begin
        int_reg_array_43_4_real <= _zz_2420_;
      end
      if(_zz_2374_)begin
        int_reg_array_43_5_real <= _zz_2420_;
      end
      if(_zz_2375_)begin
        int_reg_array_43_6_real <= _zz_2420_;
      end
      if(_zz_2376_)begin
        int_reg_array_43_7_real <= _zz_2420_;
      end
      if(_zz_2377_)begin
        int_reg_array_43_8_real <= _zz_2420_;
      end
      if(_zz_2378_)begin
        int_reg_array_43_9_real <= _zz_2420_;
      end
      if(_zz_2379_)begin
        int_reg_array_43_10_real <= _zz_2420_;
      end
      if(_zz_2380_)begin
        int_reg_array_43_11_real <= _zz_2420_;
      end
      if(_zz_2381_)begin
        int_reg_array_43_12_real <= _zz_2420_;
      end
      if(_zz_2382_)begin
        int_reg_array_43_13_real <= _zz_2420_;
      end
      if(_zz_2383_)begin
        int_reg_array_43_14_real <= _zz_2420_;
      end
      if(_zz_2384_)begin
        int_reg_array_43_15_real <= _zz_2420_;
      end
      if(_zz_2385_)begin
        int_reg_array_43_16_real <= _zz_2420_;
      end
      if(_zz_2386_)begin
        int_reg_array_43_17_real <= _zz_2420_;
      end
      if(_zz_2387_)begin
        int_reg_array_43_18_real <= _zz_2420_;
      end
      if(_zz_2388_)begin
        int_reg_array_43_19_real <= _zz_2420_;
      end
      if(_zz_2389_)begin
        int_reg_array_43_20_real <= _zz_2420_;
      end
      if(_zz_2390_)begin
        int_reg_array_43_21_real <= _zz_2420_;
      end
      if(_zz_2391_)begin
        int_reg_array_43_22_real <= _zz_2420_;
      end
      if(_zz_2392_)begin
        int_reg_array_43_23_real <= _zz_2420_;
      end
      if(_zz_2393_)begin
        int_reg_array_43_24_real <= _zz_2420_;
      end
      if(_zz_2394_)begin
        int_reg_array_43_25_real <= _zz_2420_;
      end
      if(_zz_2395_)begin
        int_reg_array_43_26_real <= _zz_2420_;
      end
      if(_zz_2396_)begin
        int_reg_array_43_27_real <= _zz_2420_;
      end
      if(_zz_2397_)begin
        int_reg_array_43_28_real <= _zz_2420_;
      end
      if(_zz_2398_)begin
        int_reg_array_43_29_real <= _zz_2420_;
      end
      if(_zz_2399_)begin
        int_reg_array_43_30_real <= _zz_2420_;
      end
      if(_zz_2400_)begin
        int_reg_array_43_31_real <= _zz_2420_;
      end
      if(_zz_2401_)begin
        int_reg_array_43_32_real <= _zz_2420_;
      end
      if(_zz_2402_)begin
        int_reg_array_43_33_real <= _zz_2420_;
      end
      if(_zz_2403_)begin
        int_reg_array_43_34_real <= _zz_2420_;
      end
      if(_zz_2404_)begin
        int_reg_array_43_35_real <= _zz_2420_;
      end
      if(_zz_2405_)begin
        int_reg_array_43_36_real <= _zz_2420_;
      end
      if(_zz_2406_)begin
        int_reg_array_43_37_real <= _zz_2420_;
      end
      if(_zz_2407_)begin
        int_reg_array_43_38_real <= _zz_2420_;
      end
      if(_zz_2408_)begin
        int_reg_array_43_39_real <= _zz_2420_;
      end
      if(_zz_2409_)begin
        int_reg_array_43_40_real <= _zz_2420_;
      end
      if(_zz_2410_)begin
        int_reg_array_43_41_real <= _zz_2420_;
      end
      if(_zz_2411_)begin
        int_reg_array_43_42_real <= _zz_2420_;
      end
      if(_zz_2412_)begin
        int_reg_array_43_43_real <= _zz_2420_;
      end
      if(_zz_2413_)begin
        int_reg_array_43_44_real <= _zz_2420_;
      end
      if(_zz_2414_)begin
        int_reg_array_43_45_real <= _zz_2420_;
      end
      if(_zz_2415_)begin
        int_reg_array_43_46_real <= _zz_2420_;
      end
      if(_zz_2416_)begin
        int_reg_array_43_47_real <= _zz_2420_;
      end
      if(_zz_2417_)begin
        int_reg_array_43_48_real <= _zz_2420_;
      end
      if(_zz_2418_)begin
        int_reg_array_43_49_real <= _zz_2420_;
      end
      if(_zz_2369_)begin
        int_reg_array_43_0_imag <= _zz_2421_;
      end
      if(_zz_2370_)begin
        int_reg_array_43_1_imag <= _zz_2421_;
      end
      if(_zz_2371_)begin
        int_reg_array_43_2_imag <= _zz_2421_;
      end
      if(_zz_2372_)begin
        int_reg_array_43_3_imag <= _zz_2421_;
      end
      if(_zz_2373_)begin
        int_reg_array_43_4_imag <= _zz_2421_;
      end
      if(_zz_2374_)begin
        int_reg_array_43_5_imag <= _zz_2421_;
      end
      if(_zz_2375_)begin
        int_reg_array_43_6_imag <= _zz_2421_;
      end
      if(_zz_2376_)begin
        int_reg_array_43_7_imag <= _zz_2421_;
      end
      if(_zz_2377_)begin
        int_reg_array_43_8_imag <= _zz_2421_;
      end
      if(_zz_2378_)begin
        int_reg_array_43_9_imag <= _zz_2421_;
      end
      if(_zz_2379_)begin
        int_reg_array_43_10_imag <= _zz_2421_;
      end
      if(_zz_2380_)begin
        int_reg_array_43_11_imag <= _zz_2421_;
      end
      if(_zz_2381_)begin
        int_reg_array_43_12_imag <= _zz_2421_;
      end
      if(_zz_2382_)begin
        int_reg_array_43_13_imag <= _zz_2421_;
      end
      if(_zz_2383_)begin
        int_reg_array_43_14_imag <= _zz_2421_;
      end
      if(_zz_2384_)begin
        int_reg_array_43_15_imag <= _zz_2421_;
      end
      if(_zz_2385_)begin
        int_reg_array_43_16_imag <= _zz_2421_;
      end
      if(_zz_2386_)begin
        int_reg_array_43_17_imag <= _zz_2421_;
      end
      if(_zz_2387_)begin
        int_reg_array_43_18_imag <= _zz_2421_;
      end
      if(_zz_2388_)begin
        int_reg_array_43_19_imag <= _zz_2421_;
      end
      if(_zz_2389_)begin
        int_reg_array_43_20_imag <= _zz_2421_;
      end
      if(_zz_2390_)begin
        int_reg_array_43_21_imag <= _zz_2421_;
      end
      if(_zz_2391_)begin
        int_reg_array_43_22_imag <= _zz_2421_;
      end
      if(_zz_2392_)begin
        int_reg_array_43_23_imag <= _zz_2421_;
      end
      if(_zz_2393_)begin
        int_reg_array_43_24_imag <= _zz_2421_;
      end
      if(_zz_2394_)begin
        int_reg_array_43_25_imag <= _zz_2421_;
      end
      if(_zz_2395_)begin
        int_reg_array_43_26_imag <= _zz_2421_;
      end
      if(_zz_2396_)begin
        int_reg_array_43_27_imag <= _zz_2421_;
      end
      if(_zz_2397_)begin
        int_reg_array_43_28_imag <= _zz_2421_;
      end
      if(_zz_2398_)begin
        int_reg_array_43_29_imag <= _zz_2421_;
      end
      if(_zz_2399_)begin
        int_reg_array_43_30_imag <= _zz_2421_;
      end
      if(_zz_2400_)begin
        int_reg_array_43_31_imag <= _zz_2421_;
      end
      if(_zz_2401_)begin
        int_reg_array_43_32_imag <= _zz_2421_;
      end
      if(_zz_2402_)begin
        int_reg_array_43_33_imag <= _zz_2421_;
      end
      if(_zz_2403_)begin
        int_reg_array_43_34_imag <= _zz_2421_;
      end
      if(_zz_2404_)begin
        int_reg_array_43_35_imag <= _zz_2421_;
      end
      if(_zz_2405_)begin
        int_reg_array_43_36_imag <= _zz_2421_;
      end
      if(_zz_2406_)begin
        int_reg_array_43_37_imag <= _zz_2421_;
      end
      if(_zz_2407_)begin
        int_reg_array_43_38_imag <= _zz_2421_;
      end
      if(_zz_2408_)begin
        int_reg_array_43_39_imag <= _zz_2421_;
      end
      if(_zz_2409_)begin
        int_reg_array_43_40_imag <= _zz_2421_;
      end
      if(_zz_2410_)begin
        int_reg_array_43_41_imag <= _zz_2421_;
      end
      if(_zz_2411_)begin
        int_reg_array_43_42_imag <= _zz_2421_;
      end
      if(_zz_2412_)begin
        int_reg_array_43_43_imag <= _zz_2421_;
      end
      if(_zz_2413_)begin
        int_reg_array_43_44_imag <= _zz_2421_;
      end
      if(_zz_2414_)begin
        int_reg_array_43_45_imag <= _zz_2421_;
      end
      if(_zz_2415_)begin
        int_reg_array_43_46_imag <= _zz_2421_;
      end
      if(_zz_2416_)begin
        int_reg_array_43_47_imag <= _zz_2421_;
      end
      if(_zz_2417_)begin
        int_reg_array_43_48_imag <= _zz_2421_;
      end
      if(_zz_2418_)begin
        int_reg_array_43_49_imag <= _zz_2421_;
      end
      if(_zz_2424_)begin
        int_reg_array_44_0_real <= _zz_2475_;
      end
      if(_zz_2425_)begin
        int_reg_array_44_1_real <= _zz_2475_;
      end
      if(_zz_2426_)begin
        int_reg_array_44_2_real <= _zz_2475_;
      end
      if(_zz_2427_)begin
        int_reg_array_44_3_real <= _zz_2475_;
      end
      if(_zz_2428_)begin
        int_reg_array_44_4_real <= _zz_2475_;
      end
      if(_zz_2429_)begin
        int_reg_array_44_5_real <= _zz_2475_;
      end
      if(_zz_2430_)begin
        int_reg_array_44_6_real <= _zz_2475_;
      end
      if(_zz_2431_)begin
        int_reg_array_44_7_real <= _zz_2475_;
      end
      if(_zz_2432_)begin
        int_reg_array_44_8_real <= _zz_2475_;
      end
      if(_zz_2433_)begin
        int_reg_array_44_9_real <= _zz_2475_;
      end
      if(_zz_2434_)begin
        int_reg_array_44_10_real <= _zz_2475_;
      end
      if(_zz_2435_)begin
        int_reg_array_44_11_real <= _zz_2475_;
      end
      if(_zz_2436_)begin
        int_reg_array_44_12_real <= _zz_2475_;
      end
      if(_zz_2437_)begin
        int_reg_array_44_13_real <= _zz_2475_;
      end
      if(_zz_2438_)begin
        int_reg_array_44_14_real <= _zz_2475_;
      end
      if(_zz_2439_)begin
        int_reg_array_44_15_real <= _zz_2475_;
      end
      if(_zz_2440_)begin
        int_reg_array_44_16_real <= _zz_2475_;
      end
      if(_zz_2441_)begin
        int_reg_array_44_17_real <= _zz_2475_;
      end
      if(_zz_2442_)begin
        int_reg_array_44_18_real <= _zz_2475_;
      end
      if(_zz_2443_)begin
        int_reg_array_44_19_real <= _zz_2475_;
      end
      if(_zz_2444_)begin
        int_reg_array_44_20_real <= _zz_2475_;
      end
      if(_zz_2445_)begin
        int_reg_array_44_21_real <= _zz_2475_;
      end
      if(_zz_2446_)begin
        int_reg_array_44_22_real <= _zz_2475_;
      end
      if(_zz_2447_)begin
        int_reg_array_44_23_real <= _zz_2475_;
      end
      if(_zz_2448_)begin
        int_reg_array_44_24_real <= _zz_2475_;
      end
      if(_zz_2449_)begin
        int_reg_array_44_25_real <= _zz_2475_;
      end
      if(_zz_2450_)begin
        int_reg_array_44_26_real <= _zz_2475_;
      end
      if(_zz_2451_)begin
        int_reg_array_44_27_real <= _zz_2475_;
      end
      if(_zz_2452_)begin
        int_reg_array_44_28_real <= _zz_2475_;
      end
      if(_zz_2453_)begin
        int_reg_array_44_29_real <= _zz_2475_;
      end
      if(_zz_2454_)begin
        int_reg_array_44_30_real <= _zz_2475_;
      end
      if(_zz_2455_)begin
        int_reg_array_44_31_real <= _zz_2475_;
      end
      if(_zz_2456_)begin
        int_reg_array_44_32_real <= _zz_2475_;
      end
      if(_zz_2457_)begin
        int_reg_array_44_33_real <= _zz_2475_;
      end
      if(_zz_2458_)begin
        int_reg_array_44_34_real <= _zz_2475_;
      end
      if(_zz_2459_)begin
        int_reg_array_44_35_real <= _zz_2475_;
      end
      if(_zz_2460_)begin
        int_reg_array_44_36_real <= _zz_2475_;
      end
      if(_zz_2461_)begin
        int_reg_array_44_37_real <= _zz_2475_;
      end
      if(_zz_2462_)begin
        int_reg_array_44_38_real <= _zz_2475_;
      end
      if(_zz_2463_)begin
        int_reg_array_44_39_real <= _zz_2475_;
      end
      if(_zz_2464_)begin
        int_reg_array_44_40_real <= _zz_2475_;
      end
      if(_zz_2465_)begin
        int_reg_array_44_41_real <= _zz_2475_;
      end
      if(_zz_2466_)begin
        int_reg_array_44_42_real <= _zz_2475_;
      end
      if(_zz_2467_)begin
        int_reg_array_44_43_real <= _zz_2475_;
      end
      if(_zz_2468_)begin
        int_reg_array_44_44_real <= _zz_2475_;
      end
      if(_zz_2469_)begin
        int_reg_array_44_45_real <= _zz_2475_;
      end
      if(_zz_2470_)begin
        int_reg_array_44_46_real <= _zz_2475_;
      end
      if(_zz_2471_)begin
        int_reg_array_44_47_real <= _zz_2475_;
      end
      if(_zz_2472_)begin
        int_reg_array_44_48_real <= _zz_2475_;
      end
      if(_zz_2473_)begin
        int_reg_array_44_49_real <= _zz_2475_;
      end
      if(_zz_2424_)begin
        int_reg_array_44_0_imag <= _zz_2476_;
      end
      if(_zz_2425_)begin
        int_reg_array_44_1_imag <= _zz_2476_;
      end
      if(_zz_2426_)begin
        int_reg_array_44_2_imag <= _zz_2476_;
      end
      if(_zz_2427_)begin
        int_reg_array_44_3_imag <= _zz_2476_;
      end
      if(_zz_2428_)begin
        int_reg_array_44_4_imag <= _zz_2476_;
      end
      if(_zz_2429_)begin
        int_reg_array_44_5_imag <= _zz_2476_;
      end
      if(_zz_2430_)begin
        int_reg_array_44_6_imag <= _zz_2476_;
      end
      if(_zz_2431_)begin
        int_reg_array_44_7_imag <= _zz_2476_;
      end
      if(_zz_2432_)begin
        int_reg_array_44_8_imag <= _zz_2476_;
      end
      if(_zz_2433_)begin
        int_reg_array_44_9_imag <= _zz_2476_;
      end
      if(_zz_2434_)begin
        int_reg_array_44_10_imag <= _zz_2476_;
      end
      if(_zz_2435_)begin
        int_reg_array_44_11_imag <= _zz_2476_;
      end
      if(_zz_2436_)begin
        int_reg_array_44_12_imag <= _zz_2476_;
      end
      if(_zz_2437_)begin
        int_reg_array_44_13_imag <= _zz_2476_;
      end
      if(_zz_2438_)begin
        int_reg_array_44_14_imag <= _zz_2476_;
      end
      if(_zz_2439_)begin
        int_reg_array_44_15_imag <= _zz_2476_;
      end
      if(_zz_2440_)begin
        int_reg_array_44_16_imag <= _zz_2476_;
      end
      if(_zz_2441_)begin
        int_reg_array_44_17_imag <= _zz_2476_;
      end
      if(_zz_2442_)begin
        int_reg_array_44_18_imag <= _zz_2476_;
      end
      if(_zz_2443_)begin
        int_reg_array_44_19_imag <= _zz_2476_;
      end
      if(_zz_2444_)begin
        int_reg_array_44_20_imag <= _zz_2476_;
      end
      if(_zz_2445_)begin
        int_reg_array_44_21_imag <= _zz_2476_;
      end
      if(_zz_2446_)begin
        int_reg_array_44_22_imag <= _zz_2476_;
      end
      if(_zz_2447_)begin
        int_reg_array_44_23_imag <= _zz_2476_;
      end
      if(_zz_2448_)begin
        int_reg_array_44_24_imag <= _zz_2476_;
      end
      if(_zz_2449_)begin
        int_reg_array_44_25_imag <= _zz_2476_;
      end
      if(_zz_2450_)begin
        int_reg_array_44_26_imag <= _zz_2476_;
      end
      if(_zz_2451_)begin
        int_reg_array_44_27_imag <= _zz_2476_;
      end
      if(_zz_2452_)begin
        int_reg_array_44_28_imag <= _zz_2476_;
      end
      if(_zz_2453_)begin
        int_reg_array_44_29_imag <= _zz_2476_;
      end
      if(_zz_2454_)begin
        int_reg_array_44_30_imag <= _zz_2476_;
      end
      if(_zz_2455_)begin
        int_reg_array_44_31_imag <= _zz_2476_;
      end
      if(_zz_2456_)begin
        int_reg_array_44_32_imag <= _zz_2476_;
      end
      if(_zz_2457_)begin
        int_reg_array_44_33_imag <= _zz_2476_;
      end
      if(_zz_2458_)begin
        int_reg_array_44_34_imag <= _zz_2476_;
      end
      if(_zz_2459_)begin
        int_reg_array_44_35_imag <= _zz_2476_;
      end
      if(_zz_2460_)begin
        int_reg_array_44_36_imag <= _zz_2476_;
      end
      if(_zz_2461_)begin
        int_reg_array_44_37_imag <= _zz_2476_;
      end
      if(_zz_2462_)begin
        int_reg_array_44_38_imag <= _zz_2476_;
      end
      if(_zz_2463_)begin
        int_reg_array_44_39_imag <= _zz_2476_;
      end
      if(_zz_2464_)begin
        int_reg_array_44_40_imag <= _zz_2476_;
      end
      if(_zz_2465_)begin
        int_reg_array_44_41_imag <= _zz_2476_;
      end
      if(_zz_2466_)begin
        int_reg_array_44_42_imag <= _zz_2476_;
      end
      if(_zz_2467_)begin
        int_reg_array_44_43_imag <= _zz_2476_;
      end
      if(_zz_2468_)begin
        int_reg_array_44_44_imag <= _zz_2476_;
      end
      if(_zz_2469_)begin
        int_reg_array_44_45_imag <= _zz_2476_;
      end
      if(_zz_2470_)begin
        int_reg_array_44_46_imag <= _zz_2476_;
      end
      if(_zz_2471_)begin
        int_reg_array_44_47_imag <= _zz_2476_;
      end
      if(_zz_2472_)begin
        int_reg_array_44_48_imag <= _zz_2476_;
      end
      if(_zz_2473_)begin
        int_reg_array_44_49_imag <= _zz_2476_;
      end
      if(_zz_2479_)begin
        int_reg_array_45_0_real <= _zz_2530_;
      end
      if(_zz_2480_)begin
        int_reg_array_45_1_real <= _zz_2530_;
      end
      if(_zz_2481_)begin
        int_reg_array_45_2_real <= _zz_2530_;
      end
      if(_zz_2482_)begin
        int_reg_array_45_3_real <= _zz_2530_;
      end
      if(_zz_2483_)begin
        int_reg_array_45_4_real <= _zz_2530_;
      end
      if(_zz_2484_)begin
        int_reg_array_45_5_real <= _zz_2530_;
      end
      if(_zz_2485_)begin
        int_reg_array_45_6_real <= _zz_2530_;
      end
      if(_zz_2486_)begin
        int_reg_array_45_7_real <= _zz_2530_;
      end
      if(_zz_2487_)begin
        int_reg_array_45_8_real <= _zz_2530_;
      end
      if(_zz_2488_)begin
        int_reg_array_45_9_real <= _zz_2530_;
      end
      if(_zz_2489_)begin
        int_reg_array_45_10_real <= _zz_2530_;
      end
      if(_zz_2490_)begin
        int_reg_array_45_11_real <= _zz_2530_;
      end
      if(_zz_2491_)begin
        int_reg_array_45_12_real <= _zz_2530_;
      end
      if(_zz_2492_)begin
        int_reg_array_45_13_real <= _zz_2530_;
      end
      if(_zz_2493_)begin
        int_reg_array_45_14_real <= _zz_2530_;
      end
      if(_zz_2494_)begin
        int_reg_array_45_15_real <= _zz_2530_;
      end
      if(_zz_2495_)begin
        int_reg_array_45_16_real <= _zz_2530_;
      end
      if(_zz_2496_)begin
        int_reg_array_45_17_real <= _zz_2530_;
      end
      if(_zz_2497_)begin
        int_reg_array_45_18_real <= _zz_2530_;
      end
      if(_zz_2498_)begin
        int_reg_array_45_19_real <= _zz_2530_;
      end
      if(_zz_2499_)begin
        int_reg_array_45_20_real <= _zz_2530_;
      end
      if(_zz_2500_)begin
        int_reg_array_45_21_real <= _zz_2530_;
      end
      if(_zz_2501_)begin
        int_reg_array_45_22_real <= _zz_2530_;
      end
      if(_zz_2502_)begin
        int_reg_array_45_23_real <= _zz_2530_;
      end
      if(_zz_2503_)begin
        int_reg_array_45_24_real <= _zz_2530_;
      end
      if(_zz_2504_)begin
        int_reg_array_45_25_real <= _zz_2530_;
      end
      if(_zz_2505_)begin
        int_reg_array_45_26_real <= _zz_2530_;
      end
      if(_zz_2506_)begin
        int_reg_array_45_27_real <= _zz_2530_;
      end
      if(_zz_2507_)begin
        int_reg_array_45_28_real <= _zz_2530_;
      end
      if(_zz_2508_)begin
        int_reg_array_45_29_real <= _zz_2530_;
      end
      if(_zz_2509_)begin
        int_reg_array_45_30_real <= _zz_2530_;
      end
      if(_zz_2510_)begin
        int_reg_array_45_31_real <= _zz_2530_;
      end
      if(_zz_2511_)begin
        int_reg_array_45_32_real <= _zz_2530_;
      end
      if(_zz_2512_)begin
        int_reg_array_45_33_real <= _zz_2530_;
      end
      if(_zz_2513_)begin
        int_reg_array_45_34_real <= _zz_2530_;
      end
      if(_zz_2514_)begin
        int_reg_array_45_35_real <= _zz_2530_;
      end
      if(_zz_2515_)begin
        int_reg_array_45_36_real <= _zz_2530_;
      end
      if(_zz_2516_)begin
        int_reg_array_45_37_real <= _zz_2530_;
      end
      if(_zz_2517_)begin
        int_reg_array_45_38_real <= _zz_2530_;
      end
      if(_zz_2518_)begin
        int_reg_array_45_39_real <= _zz_2530_;
      end
      if(_zz_2519_)begin
        int_reg_array_45_40_real <= _zz_2530_;
      end
      if(_zz_2520_)begin
        int_reg_array_45_41_real <= _zz_2530_;
      end
      if(_zz_2521_)begin
        int_reg_array_45_42_real <= _zz_2530_;
      end
      if(_zz_2522_)begin
        int_reg_array_45_43_real <= _zz_2530_;
      end
      if(_zz_2523_)begin
        int_reg_array_45_44_real <= _zz_2530_;
      end
      if(_zz_2524_)begin
        int_reg_array_45_45_real <= _zz_2530_;
      end
      if(_zz_2525_)begin
        int_reg_array_45_46_real <= _zz_2530_;
      end
      if(_zz_2526_)begin
        int_reg_array_45_47_real <= _zz_2530_;
      end
      if(_zz_2527_)begin
        int_reg_array_45_48_real <= _zz_2530_;
      end
      if(_zz_2528_)begin
        int_reg_array_45_49_real <= _zz_2530_;
      end
      if(_zz_2479_)begin
        int_reg_array_45_0_imag <= _zz_2531_;
      end
      if(_zz_2480_)begin
        int_reg_array_45_1_imag <= _zz_2531_;
      end
      if(_zz_2481_)begin
        int_reg_array_45_2_imag <= _zz_2531_;
      end
      if(_zz_2482_)begin
        int_reg_array_45_3_imag <= _zz_2531_;
      end
      if(_zz_2483_)begin
        int_reg_array_45_4_imag <= _zz_2531_;
      end
      if(_zz_2484_)begin
        int_reg_array_45_5_imag <= _zz_2531_;
      end
      if(_zz_2485_)begin
        int_reg_array_45_6_imag <= _zz_2531_;
      end
      if(_zz_2486_)begin
        int_reg_array_45_7_imag <= _zz_2531_;
      end
      if(_zz_2487_)begin
        int_reg_array_45_8_imag <= _zz_2531_;
      end
      if(_zz_2488_)begin
        int_reg_array_45_9_imag <= _zz_2531_;
      end
      if(_zz_2489_)begin
        int_reg_array_45_10_imag <= _zz_2531_;
      end
      if(_zz_2490_)begin
        int_reg_array_45_11_imag <= _zz_2531_;
      end
      if(_zz_2491_)begin
        int_reg_array_45_12_imag <= _zz_2531_;
      end
      if(_zz_2492_)begin
        int_reg_array_45_13_imag <= _zz_2531_;
      end
      if(_zz_2493_)begin
        int_reg_array_45_14_imag <= _zz_2531_;
      end
      if(_zz_2494_)begin
        int_reg_array_45_15_imag <= _zz_2531_;
      end
      if(_zz_2495_)begin
        int_reg_array_45_16_imag <= _zz_2531_;
      end
      if(_zz_2496_)begin
        int_reg_array_45_17_imag <= _zz_2531_;
      end
      if(_zz_2497_)begin
        int_reg_array_45_18_imag <= _zz_2531_;
      end
      if(_zz_2498_)begin
        int_reg_array_45_19_imag <= _zz_2531_;
      end
      if(_zz_2499_)begin
        int_reg_array_45_20_imag <= _zz_2531_;
      end
      if(_zz_2500_)begin
        int_reg_array_45_21_imag <= _zz_2531_;
      end
      if(_zz_2501_)begin
        int_reg_array_45_22_imag <= _zz_2531_;
      end
      if(_zz_2502_)begin
        int_reg_array_45_23_imag <= _zz_2531_;
      end
      if(_zz_2503_)begin
        int_reg_array_45_24_imag <= _zz_2531_;
      end
      if(_zz_2504_)begin
        int_reg_array_45_25_imag <= _zz_2531_;
      end
      if(_zz_2505_)begin
        int_reg_array_45_26_imag <= _zz_2531_;
      end
      if(_zz_2506_)begin
        int_reg_array_45_27_imag <= _zz_2531_;
      end
      if(_zz_2507_)begin
        int_reg_array_45_28_imag <= _zz_2531_;
      end
      if(_zz_2508_)begin
        int_reg_array_45_29_imag <= _zz_2531_;
      end
      if(_zz_2509_)begin
        int_reg_array_45_30_imag <= _zz_2531_;
      end
      if(_zz_2510_)begin
        int_reg_array_45_31_imag <= _zz_2531_;
      end
      if(_zz_2511_)begin
        int_reg_array_45_32_imag <= _zz_2531_;
      end
      if(_zz_2512_)begin
        int_reg_array_45_33_imag <= _zz_2531_;
      end
      if(_zz_2513_)begin
        int_reg_array_45_34_imag <= _zz_2531_;
      end
      if(_zz_2514_)begin
        int_reg_array_45_35_imag <= _zz_2531_;
      end
      if(_zz_2515_)begin
        int_reg_array_45_36_imag <= _zz_2531_;
      end
      if(_zz_2516_)begin
        int_reg_array_45_37_imag <= _zz_2531_;
      end
      if(_zz_2517_)begin
        int_reg_array_45_38_imag <= _zz_2531_;
      end
      if(_zz_2518_)begin
        int_reg_array_45_39_imag <= _zz_2531_;
      end
      if(_zz_2519_)begin
        int_reg_array_45_40_imag <= _zz_2531_;
      end
      if(_zz_2520_)begin
        int_reg_array_45_41_imag <= _zz_2531_;
      end
      if(_zz_2521_)begin
        int_reg_array_45_42_imag <= _zz_2531_;
      end
      if(_zz_2522_)begin
        int_reg_array_45_43_imag <= _zz_2531_;
      end
      if(_zz_2523_)begin
        int_reg_array_45_44_imag <= _zz_2531_;
      end
      if(_zz_2524_)begin
        int_reg_array_45_45_imag <= _zz_2531_;
      end
      if(_zz_2525_)begin
        int_reg_array_45_46_imag <= _zz_2531_;
      end
      if(_zz_2526_)begin
        int_reg_array_45_47_imag <= _zz_2531_;
      end
      if(_zz_2527_)begin
        int_reg_array_45_48_imag <= _zz_2531_;
      end
      if(_zz_2528_)begin
        int_reg_array_45_49_imag <= _zz_2531_;
      end
      if(_zz_2534_)begin
        int_reg_array_46_0_real <= _zz_2585_;
      end
      if(_zz_2535_)begin
        int_reg_array_46_1_real <= _zz_2585_;
      end
      if(_zz_2536_)begin
        int_reg_array_46_2_real <= _zz_2585_;
      end
      if(_zz_2537_)begin
        int_reg_array_46_3_real <= _zz_2585_;
      end
      if(_zz_2538_)begin
        int_reg_array_46_4_real <= _zz_2585_;
      end
      if(_zz_2539_)begin
        int_reg_array_46_5_real <= _zz_2585_;
      end
      if(_zz_2540_)begin
        int_reg_array_46_6_real <= _zz_2585_;
      end
      if(_zz_2541_)begin
        int_reg_array_46_7_real <= _zz_2585_;
      end
      if(_zz_2542_)begin
        int_reg_array_46_8_real <= _zz_2585_;
      end
      if(_zz_2543_)begin
        int_reg_array_46_9_real <= _zz_2585_;
      end
      if(_zz_2544_)begin
        int_reg_array_46_10_real <= _zz_2585_;
      end
      if(_zz_2545_)begin
        int_reg_array_46_11_real <= _zz_2585_;
      end
      if(_zz_2546_)begin
        int_reg_array_46_12_real <= _zz_2585_;
      end
      if(_zz_2547_)begin
        int_reg_array_46_13_real <= _zz_2585_;
      end
      if(_zz_2548_)begin
        int_reg_array_46_14_real <= _zz_2585_;
      end
      if(_zz_2549_)begin
        int_reg_array_46_15_real <= _zz_2585_;
      end
      if(_zz_2550_)begin
        int_reg_array_46_16_real <= _zz_2585_;
      end
      if(_zz_2551_)begin
        int_reg_array_46_17_real <= _zz_2585_;
      end
      if(_zz_2552_)begin
        int_reg_array_46_18_real <= _zz_2585_;
      end
      if(_zz_2553_)begin
        int_reg_array_46_19_real <= _zz_2585_;
      end
      if(_zz_2554_)begin
        int_reg_array_46_20_real <= _zz_2585_;
      end
      if(_zz_2555_)begin
        int_reg_array_46_21_real <= _zz_2585_;
      end
      if(_zz_2556_)begin
        int_reg_array_46_22_real <= _zz_2585_;
      end
      if(_zz_2557_)begin
        int_reg_array_46_23_real <= _zz_2585_;
      end
      if(_zz_2558_)begin
        int_reg_array_46_24_real <= _zz_2585_;
      end
      if(_zz_2559_)begin
        int_reg_array_46_25_real <= _zz_2585_;
      end
      if(_zz_2560_)begin
        int_reg_array_46_26_real <= _zz_2585_;
      end
      if(_zz_2561_)begin
        int_reg_array_46_27_real <= _zz_2585_;
      end
      if(_zz_2562_)begin
        int_reg_array_46_28_real <= _zz_2585_;
      end
      if(_zz_2563_)begin
        int_reg_array_46_29_real <= _zz_2585_;
      end
      if(_zz_2564_)begin
        int_reg_array_46_30_real <= _zz_2585_;
      end
      if(_zz_2565_)begin
        int_reg_array_46_31_real <= _zz_2585_;
      end
      if(_zz_2566_)begin
        int_reg_array_46_32_real <= _zz_2585_;
      end
      if(_zz_2567_)begin
        int_reg_array_46_33_real <= _zz_2585_;
      end
      if(_zz_2568_)begin
        int_reg_array_46_34_real <= _zz_2585_;
      end
      if(_zz_2569_)begin
        int_reg_array_46_35_real <= _zz_2585_;
      end
      if(_zz_2570_)begin
        int_reg_array_46_36_real <= _zz_2585_;
      end
      if(_zz_2571_)begin
        int_reg_array_46_37_real <= _zz_2585_;
      end
      if(_zz_2572_)begin
        int_reg_array_46_38_real <= _zz_2585_;
      end
      if(_zz_2573_)begin
        int_reg_array_46_39_real <= _zz_2585_;
      end
      if(_zz_2574_)begin
        int_reg_array_46_40_real <= _zz_2585_;
      end
      if(_zz_2575_)begin
        int_reg_array_46_41_real <= _zz_2585_;
      end
      if(_zz_2576_)begin
        int_reg_array_46_42_real <= _zz_2585_;
      end
      if(_zz_2577_)begin
        int_reg_array_46_43_real <= _zz_2585_;
      end
      if(_zz_2578_)begin
        int_reg_array_46_44_real <= _zz_2585_;
      end
      if(_zz_2579_)begin
        int_reg_array_46_45_real <= _zz_2585_;
      end
      if(_zz_2580_)begin
        int_reg_array_46_46_real <= _zz_2585_;
      end
      if(_zz_2581_)begin
        int_reg_array_46_47_real <= _zz_2585_;
      end
      if(_zz_2582_)begin
        int_reg_array_46_48_real <= _zz_2585_;
      end
      if(_zz_2583_)begin
        int_reg_array_46_49_real <= _zz_2585_;
      end
      if(_zz_2534_)begin
        int_reg_array_46_0_imag <= _zz_2586_;
      end
      if(_zz_2535_)begin
        int_reg_array_46_1_imag <= _zz_2586_;
      end
      if(_zz_2536_)begin
        int_reg_array_46_2_imag <= _zz_2586_;
      end
      if(_zz_2537_)begin
        int_reg_array_46_3_imag <= _zz_2586_;
      end
      if(_zz_2538_)begin
        int_reg_array_46_4_imag <= _zz_2586_;
      end
      if(_zz_2539_)begin
        int_reg_array_46_5_imag <= _zz_2586_;
      end
      if(_zz_2540_)begin
        int_reg_array_46_6_imag <= _zz_2586_;
      end
      if(_zz_2541_)begin
        int_reg_array_46_7_imag <= _zz_2586_;
      end
      if(_zz_2542_)begin
        int_reg_array_46_8_imag <= _zz_2586_;
      end
      if(_zz_2543_)begin
        int_reg_array_46_9_imag <= _zz_2586_;
      end
      if(_zz_2544_)begin
        int_reg_array_46_10_imag <= _zz_2586_;
      end
      if(_zz_2545_)begin
        int_reg_array_46_11_imag <= _zz_2586_;
      end
      if(_zz_2546_)begin
        int_reg_array_46_12_imag <= _zz_2586_;
      end
      if(_zz_2547_)begin
        int_reg_array_46_13_imag <= _zz_2586_;
      end
      if(_zz_2548_)begin
        int_reg_array_46_14_imag <= _zz_2586_;
      end
      if(_zz_2549_)begin
        int_reg_array_46_15_imag <= _zz_2586_;
      end
      if(_zz_2550_)begin
        int_reg_array_46_16_imag <= _zz_2586_;
      end
      if(_zz_2551_)begin
        int_reg_array_46_17_imag <= _zz_2586_;
      end
      if(_zz_2552_)begin
        int_reg_array_46_18_imag <= _zz_2586_;
      end
      if(_zz_2553_)begin
        int_reg_array_46_19_imag <= _zz_2586_;
      end
      if(_zz_2554_)begin
        int_reg_array_46_20_imag <= _zz_2586_;
      end
      if(_zz_2555_)begin
        int_reg_array_46_21_imag <= _zz_2586_;
      end
      if(_zz_2556_)begin
        int_reg_array_46_22_imag <= _zz_2586_;
      end
      if(_zz_2557_)begin
        int_reg_array_46_23_imag <= _zz_2586_;
      end
      if(_zz_2558_)begin
        int_reg_array_46_24_imag <= _zz_2586_;
      end
      if(_zz_2559_)begin
        int_reg_array_46_25_imag <= _zz_2586_;
      end
      if(_zz_2560_)begin
        int_reg_array_46_26_imag <= _zz_2586_;
      end
      if(_zz_2561_)begin
        int_reg_array_46_27_imag <= _zz_2586_;
      end
      if(_zz_2562_)begin
        int_reg_array_46_28_imag <= _zz_2586_;
      end
      if(_zz_2563_)begin
        int_reg_array_46_29_imag <= _zz_2586_;
      end
      if(_zz_2564_)begin
        int_reg_array_46_30_imag <= _zz_2586_;
      end
      if(_zz_2565_)begin
        int_reg_array_46_31_imag <= _zz_2586_;
      end
      if(_zz_2566_)begin
        int_reg_array_46_32_imag <= _zz_2586_;
      end
      if(_zz_2567_)begin
        int_reg_array_46_33_imag <= _zz_2586_;
      end
      if(_zz_2568_)begin
        int_reg_array_46_34_imag <= _zz_2586_;
      end
      if(_zz_2569_)begin
        int_reg_array_46_35_imag <= _zz_2586_;
      end
      if(_zz_2570_)begin
        int_reg_array_46_36_imag <= _zz_2586_;
      end
      if(_zz_2571_)begin
        int_reg_array_46_37_imag <= _zz_2586_;
      end
      if(_zz_2572_)begin
        int_reg_array_46_38_imag <= _zz_2586_;
      end
      if(_zz_2573_)begin
        int_reg_array_46_39_imag <= _zz_2586_;
      end
      if(_zz_2574_)begin
        int_reg_array_46_40_imag <= _zz_2586_;
      end
      if(_zz_2575_)begin
        int_reg_array_46_41_imag <= _zz_2586_;
      end
      if(_zz_2576_)begin
        int_reg_array_46_42_imag <= _zz_2586_;
      end
      if(_zz_2577_)begin
        int_reg_array_46_43_imag <= _zz_2586_;
      end
      if(_zz_2578_)begin
        int_reg_array_46_44_imag <= _zz_2586_;
      end
      if(_zz_2579_)begin
        int_reg_array_46_45_imag <= _zz_2586_;
      end
      if(_zz_2580_)begin
        int_reg_array_46_46_imag <= _zz_2586_;
      end
      if(_zz_2581_)begin
        int_reg_array_46_47_imag <= _zz_2586_;
      end
      if(_zz_2582_)begin
        int_reg_array_46_48_imag <= _zz_2586_;
      end
      if(_zz_2583_)begin
        int_reg_array_46_49_imag <= _zz_2586_;
      end
      if(_zz_2589_)begin
        int_reg_array_47_0_real <= _zz_2640_;
      end
      if(_zz_2590_)begin
        int_reg_array_47_1_real <= _zz_2640_;
      end
      if(_zz_2591_)begin
        int_reg_array_47_2_real <= _zz_2640_;
      end
      if(_zz_2592_)begin
        int_reg_array_47_3_real <= _zz_2640_;
      end
      if(_zz_2593_)begin
        int_reg_array_47_4_real <= _zz_2640_;
      end
      if(_zz_2594_)begin
        int_reg_array_47_5_real <= _zz_2640_;
      end
      if(_zz_2595_)begin
        int_reg_array_47_6_real <= _zz_2640_;
      end
      if(_zz_2596_)begin
        int_reg_array_47_7_real <= _zz_2640_;
      end
      if(_zz_2597_)begin
        int_reg_array_47_8_real <= _zz_2640_;
      end
      if(_zz_2598_)begin
        int_reg_array_47_9_real <= _zz_2640_;
      end
      if(_zz_2599_)begin
        int_reg_array_47_10_real <= _zz_2640_;
      end
      if(_zz_2600_)begin
        int_reg_array_47_11_real <= _zz_2640_;
      end
      if(_zz_2601_)begin
        int_reg_array_47_12_real <= _zz_2640_;
      end
      if(_zz_2602_)begin
        int_reg_array_47_13_real <= _zz_2640_;
      end
      if(_zz_2603_)begin
        int_reg_array_47_14_real <= _zz_2640_;
      end
      if(_zz_2604_)begin
        int_reg_array_47_15_real <= _zz_2640_;
      end
      if(_zz_2605_)begin
        int_reg_array_47_16_real <= _zz_2640_;
      end
      if(_zz_2606_)begin
        int_reg_array_47_17_real <= _zz_2640_;
      end
      if(_zz_2607_)begin
        int_reg_array_47_18_real <= _zz_2640_;
      end
      if(_zz_2608_)begin
        int_reg_array_47_19_real <= _zz_2640_;
      end
      if(_zz_2609_)begin
        int_reg_array_47_20_real <= _zz_2640_;
      end
      if(_zz_2610_)begin
        int_reg_array_47_21_real <= _zz_2640_;
      end
      if(_zz_2611_)begin
        int_reg_array_47_22_real <= _zz_2640_;
      end
      if(_zz_2612_)begin
        int_reg_array_47_23_real <= _zz_2640_;
      end
      if(_zz_2613_)begin
        int_reg_array_47_24_real <= _zz_2640_;
      end
      if(_zz_2614_)begin
        int_reg_array_47_25_real <= _zz_2640_;
      end
      if(_zz_2615_)begin
        int_reg_array_47_26_real <= _zz_2640_;
      end
      if(_zz_2616_)begin
        int_reg_array_47_27_real <= _zz_2640_;
      end
      if(_zz_2617_)begin
        int_reg_array_47_28_real <= _zz_2640_;
      end
      if(_zz_2618_)begin
        int_reg_array_47_29_real <= _zz_2640_;
      end
      if(_zz_2619_)begin
        int_reg_array_47_30_real <= _zz_2640_;
      end
      if(_zz_2620_)begin
        int_reg_array_47_31_real <= _zz_2640_;
      end
      if(_zz_2621_)begin
        int_reg_array_47_32_real <= _zz_2640_;
      end
      if(_zz_2622_)begin
        int_reg_array_47_33_real <= _zz_2640_;
      end
      if(_zz_2623_)begin
        int_reg_array_47_34_real <= _zz_2640_;
      end
      if(_zz_2624_)begin
        int_reg_array_47_35_real <= _zz_2640_;
      end
      if(_zz_2625_)begin
        int_reg_array_47_36_real <= _zz_2640_;
      end
      if(_zz_2626_)begin
        int_reg_array_47_37_real <= _zz_2640_;
      end
      if(_zz_2627_)begin
        int_reg_array_47_38_real <= _zz_2640_;
      end
      if(_zz_2628_)begin
        int_reg_array_47_39_real <= _zz_2640_;
      end
      if(_zz_2629_)begin
        int_reg_array_47_40_real <= _zz_2640_;
      end
      if(_zz_2630_)begin
        int_reg_array_47_41_real <= _zz_2640_;
      end
      if(_zz_2631_)begin
        int_reg_array_47_42_real <= _zz_2640_;
      end
      if(_zz_2632_)begin
        int_reg_array_47_43_real <= _zz_2640_;
      end
      if(_zz_2633_)begin
        int_reg_array_47_44_real <= _zz_2640_;
      end
      if(_zz_2634_)begin
        int_reg_array_47_45_real <= _zz_2640_;
      end
      if(_zz_2635_)begin
        int_reg_array_47_46_real <= _zz_2640_;
      end
      if(_zz_2636_)begin
        int_reg_array_47_47_real <= _zz_2640_;
      end
      if(_zz_2637_)begin
        int_reg_array_47_48_real <= _zz_2640_;
      end
      if(_zz_2638_)begin
        int_reg_array_47_49_real <= _zz_2640_;
      end
      if(_zz_2589_)begin
        int_reg_array_47_0_imag <= _zz_2641_;
      end
      if(_zz_2590_)begin
        int_reg_array_47_1_imag <= _zz_2641_;
      end
      if(_zz_2591_)begin
        int_reg_array_47_2_imag <= _zz_2641_;
      end
      if(_zz_2592_)begin
        int_reg_array_47_3_imag <= _zz_2641_;
      end
      if(_zz_2593_)begin
        int_reg_array_47_4_imag <= _zz_2641_;
      end
      if(_zz_2594_)begin
        int_reg_array_47_5_imag <= _zz_2641_;
      end
      if(_zz_2595_)begin
        int_reg_array_47_6_imag <= _zz_2641_;
      end
      if(_zz_2596_)begin
        int_reg_array_47_7_imag <= _zz_2641_;
      end
      if(_zz_2597_)begin
        int_reg_array_47_8_imag <= _zz_2641_;
      end
      if(_zz_2598_)begin
        int_reg_array_47_9_imag <= _zz_2641_;
      end
      if(_zz_2599_)begin
        int_reg_array_47_10_imag <= _zz_2641_;
      end
      if(_zz_2600_)begin
        int_reg_array_47_11_imag <= _zz_2641_;
      end
      if(_zz_2601_)begin
        int_reg_array_47_12_imag <= _zz_2641_;
      end
      if(_zz_2602_)begin
        int_reg_array_47_13_imag <= _zz_2641_;
      end
      if(_zz_2603_)begin
        int_reg_array_47_14_imag <= _zz_2641_;
      end
      if(_zz_2604_)begin
        int_reg_array_47_15_imag <= _zz_2641_;
      end
      if(_zz_2605_)begin
        int_reg_array_47_16_imag <= _zz_2641_;
      end
      if(_zz_2606_)begin
        int_reg_array_47_17_imag <= _zz_2641_;
      end
      if(_zz_2607_)begin
        int_reg_array_47_18_imag <= _zz_2641_;
      end
      if(_zz_2608_)begin
        int_reg_array_47_19_imag <= _zz_2641_;
      end
      if(_zz_2609_)begin
        int_reg_array_47_20_imag <= _zz_2641_;
      end
      if(_zz_2610_)begin
        int_reg_array_47_21_imag <= _zz_2641_;
      end
      if(_zz_2611_)begin
        int_reg_array_47_22_imag <= _zz_2641_;
      end
      if(_zz_2612_)begin
        int_reg_array_47_23_imag <= _zz_2641_;
      end
      if(_zz_2613_)begin
        int_reg_array_47_24_imag <= _zz_2641_;
      end
      if(_zz_2614_)begin
        int_reg_array_47_25_imag <= _zz_2641_;
      end
      if(_zz_2615_)begin
        int_reg_array_47_26_imag <= _zz_2641_;
      end
      if(_zz_2616_)begin
        int_reg_array_47_27_imag <= _zz_2641_;
      end
      if(_zz_2617_)begin
        int_reg_array_47_28_imag <= _zz_2641_;
      end
      if(_zz_2618_)begin
        int_reg_array_47_29_imag <= _zz_2641_;
      end
      if(_zz_2619_)begin
        int_reg_array_47_30_imag <= _zz_2641_;
      end
      if(_zz_2620_)begin
        int_reg_array_47_31_imag <= _zz_2641_;
      end
      if(_zz_2621_)begin
        int_reg_array_47_32_imag <= _zz_2641_;
      end
      if(_zz_2622_)begin
        int_reg_array_47_33_imag <= _zz_2641_;
      end
      if(_zz_2623_)begin
        int_reg_array_47_34_imag <= _zz_2641_;
      end
      if(_zz_2624_)begin
        int_reg_array_47_35_imag <= _zz_2641_;
      end
      if(_zz_2625_)begin
        int_reg_array_47_36_imag <= _zz_2641_;
      end
      if(_zz_2626_)begin
        int_reg_array_47_37_imag <= _zz_2641_;
      end
      if(_zz_2627_)begin
        int_reg_array_47_38_imag <= _zz_2641_;
      end
      if(_zz_2628_)begin
        int_reg_array_47_39_imag <= _zz_2641_;
      end
      if(_zz_2629_)begin
        int_reg_array_47_40_imag <= _zz_2641_;
      end
      if(_zz_2630_)begin
        int_reg_array_47_41_imag <= _zz_2641_;
      end
      if(_zz_2631_)begin
        int_reg_array_47_42_imag <= _zz_2641_;
      end
      if(_zz_2632_)begin
        int_reg_array_47_43_imag <= _zz_2641_;
      end
      if(_zz_2633_)begin
        int_reg_array_47_44_imag <= _zz_2641_;
      end
      if(_zz_2634_)begin
        int_reg_array_47_45_imag <= _zz_2641_;
      end
      if(_zz_2635_)begin
        int_reg_array_47_46_imag <= _zz_2641_;
      end
      if(_zz_2636_)begin
        int_reg_array_47_47_imag <= _zz_2641_;
      end
      if(_zz_2637_)begin
        int_reg_array_47_48_imag <= _zz_2641_;
      end
      if(_zz_2638_)begin
        int_reg_array_47_49_imag <= _zz_2641_;
      end
      if(_zz_2644_)begin
        int_reg_array_48_0_real <= _zz_2695_;
      end
      if(_zz_2645_)begin
        int_reg_array_48_1_real <= _zz_2695_;
      end
      if(_zz_2646_)begin
        int_reg_array_48_2_real <= _zz_2695_;
      end
      if(_zz_2647_)begin
        int_reg_array_48_3_real <= _zz_2695_;
      end
      if(_zz_2648_)begin
        int_reg_array_48_4_real <= _zz_2695_;
      end
      if(_zz_2649_)begin
        int_reg_array_48_5_real <= _zz_2695_;
      end
      if(_zz_2650_)begin
        int_reg_array_48_6_real <= _zz_2695_;
      end
      if(_zz_2651_)begin
        int_reg_array_48_7_real <= _zz_2695_;
      end
      if(_zz_2652_)begin
        int_reg_array_48_8_real <= _zz_2695_;
      end
      if(_zz_2653_)begin
        int_reg_array_48_9_real <= _zz_2695_;
      end
      if(_zz_2654_)begin
        int_reg_array_48_10_real <= _zz_2695_;
      end
      if(_zz_2655_)begin
        int_reg_array_48_11_real <= _zz_2695_;
      end
      if(_zz_2656_)begin
        int_reg_array_48_12_real <= _zz_2695_;
      end
      if(_zz_2657_)begin
        int_reg_array_48_13_real <= _zz_2695_;
      end
      if(_zz_2658_)begin
        int_reg_array_48_14_real <= _zz_2695_;
      end
      if(_zz_2659_)begin
        int_reg_array_48_15_real <= _zz_2695_;
      end
      if(_zz_2660_)begin
        int_reg_array_48_16_real <= _zz_2695_;
      end
      if(_zz_2661_)begin
        int_reg_array_48_17_real <= _zz_2695_;
      end
      if(_zz_2662_)begin
        int_reg_array_48_18_real <= _zz_2695_;
      end
      if(_zz_2663_)begin
        int_reg_array_48_19_real <= _zz_2695_;
      end
      if(_zz_2664_)begin
        int_reg_array_48_20_real <= _zz_2695_;
      end
      if(_zz_2665_)begin
        int_reg_array_48_21_real <= _zz_2695_;
      end
      if(_zz_2666_)begin
        int_reg_array_48_22_real <= _zz_2695_;
      end
      if(_zz_2667_)begin
        int_reg_array_48_23_real <= _zz_2695_;
      end
      if(_zz_2668_)begin
        int_reg_array_48_24_real <= _zz_2695_;
      end
      if(_zz_2669_)begin
        int_reg_array_48_25_real <= _zz_2695_;
      end
      if(_zz_2670_)begin
        int_reg_array_48_26_real <= _zz_2695_;
      end
      if(_zz_2671_)begin
        int_reg_array_48_27_real <= _zz_2695_;
      end
      if(_zz_2672_)begin
        int_reg_array_48_28_real <= _zz_2695_;
      end
      if(_zz_2673_)begin
        int_reg_array_48_29_real <= _zz_2695_;
      end
      if(_zz_2674_)begin
        int_reg_array_48_30_real <= _zz_2695_;
      end
      if(_zz_2675_)begin
        int_reg_array_48_31_real <= _zz_2695_;
      end
      if(_zz_2676_)begin
        int_reg_array_48_32_real <= _zz_2695_;
      end
      if(_zz_2677_)begin
        int_reg_array_48_33_real <= _zz_2695_;
      end
      if(_zz_2678_)begin
        int_reg_array_48_34_real <= _zz_2695_;
      end
      if(_zz_2679_)begin
        int_reg_array_48_35_real <= _zz_2695_;
      end
      if(_zz_2680_)begin
        int_reg_array_48_36_real <= _zz_2695_;
      end
      if(_zz_2681_)begin
        int_reg_array_48_37_real <= _zz_2695_;
      end
      if(_zz_2682_)begin
        int_reg_array_48_38_real <= _zz_2695_;
      end
      if(_zz_2683_)begin
        int_reg_array_48_39_real <= _zz_2695_;
      end
      if(_zz_2684_)begin
        int_reg_array_48_40_real <= _zz_2695_;
      end
      if(_zz_2685_)begin
        int_reg_array_48_41_real <= _zz_2695_;
      end
      if(_zz_2686_)begin
        int_reg_array_48_42_real <= _zz_2695_;
      end
      if(_zz_2687_)begin
        int_reg_array_48_43_real <= _zz_2695_;
      end
      if(_zz_2688_)begin
        int_reg_array_48_44_real <= _zz_2695_;
      end
      if(_zz_2689_)begin
        int_reg_array_48_45_real <= _zz_2695_;
      end
      if(_zz_2690_)begin
        int_reg_array_48_46_real <= _zz_2695_;
      end
      if(_zz_2691_)begin
        int_reg_array_48_47_real <= _zz_2695_;
      end
      if(_zz_2692_)begin
        int_reg_array_48_48_real <= _zz_2695_;
      end
      if(_zz_2693_)begin
        int_reg_array_48_49_real <= _zz_2695_;
      end
      if(_zz_2644_)begin
        int_reg_array_48_0_imag <= _zz_2696_;
      end
      if(_zz_2645_)begin
        int_reg_array_48_1_imag <= _zz_2696_;
      end
      if(_zz_2646_)begin
        int_reg_array_48_2_imag <= _zz_2696_;
      end
      if(_zz_2647_)begin
        int_reg_array_48_3_imag <= _zz_2696_;
      end
      if(_zz_2648_)begin
        int_reg_array_48_4_imag <= _zz_2696_;
      end
      if(_zz_2649_)begin
        int_reg_array_48_5_imag <= _zz_2696_;
      end
      if(_zz_2650_)begin
        int_reg_array_48_6_imag <= _zz_2696_;
      end
      if(_zz_2651_)begin
        int_reg_array_48_7_imag <= _zz_2696_;
      end
      if(_zz_2652_)begin
        int_reg_array_48_8_imag <= _zz_2696_;
      end
      if(_zz_2653_)begin
        int_reg_array_48_9_imag <= _zz_2696_;
      end
      if(_zz_2654_)begin
        int_reg_array_48_10_imag <= _zz_2696_;
      end
      if(_zz_2655_)begin
        int_reg_array_48_11_imag <= _zz_2696_;
      end
      if(_zz_2656_)begin
        int_reg_array_48_12_imag <= _zz_2696_;
      end
      if(_zz_2657_)begin
        int_reg_array_48_13_imag <= _zz_2696_;
      end
      if(_zz_2658_)begin
        int_reg_array_48_14_imag <= _zz_2696_;
      end
      if(_zz_2659_)begin
        int_reg_array_48_15_imag <= _zz_2696_;
      end
      if(_zz_2660_)begin
        int_reg_array_48_16_imag <= _zz_2696_;
      end
      if(_zz_2661_)begin
        int_reg_array_48_17_imag <= _zz_2696_;
      end
      if(_zz_2662_)begin
        int_reg_array_48_18_imag <= _zz_2696_;
      end
      if(_zz_2663_)begin
        int_reg_array_48_19_imag <= _zz_2696_;
      end
      if(_zz_2664_)begin
        int_reg_array_48_20_imag <= _zz_2696_;
      end
      if(_zz_2665_)begin
        int_reg_array_48_21_imag <= _zz_2696_;
      end
      if(_zz_2666_)begin
        int_reg_array_48_22_imag <= _zz_2696_;
      end
      if(_zz_2667_)begin
        int_reg_array_48_23_imag <= _zz_2696_;
      end
      if(_zz_2668_)begin
        int_reg_array_48_24_imag <= _zz_2696_;
      end
      if(_zz_2669_)begin
        int_reg_array_48_25_imag <= _zz_2696_;
      end
      if(_zz_2670_)begin
        int_reg_array_48_26_imag <= _zz_2696_;
      end
      if(_zz_2671_)begin
        int_reg_array_48_27_imag <= _zz_2696_;
      end
      if(_zz_2672_)begin
        int_reg_array_48_28_imag <= _zz_2696_;
      end
      if(_zz_2673_)begin
        int_reg_array_48_29_imag <= _zz_2696_;
      end
      if(_zz_2674_)begin
        int_reg_array_48_30_imag <= _zz_2696_;
      end
      if(_zz_2675_)begin
        int_reg_array_48_31_imag <= _zz_2696_;
      end
      if(_zz_2676_)begin
        int_reg_array_48_32_imag <= _zz_2696_;
      end
      if(_zz_2677_)begin
        int_reg_array_48_33_imag <= _zz_2696_;
      end
      if(_zz_2678_)begin
        int_reg_array_48_34_imag <= _zz_2696_;
      end
      if(_zz_2679_)begin
        int_reg_array_48_35_imag <= _zz_2696_;
      end
      if(_zz_2680_)begin
        int_reg_array_48_36_imag <= _zz_2696_;
      end
      if(_zz_2681_)begin
        int_reg_array_48_37_imag <= _zz_2696_;
      end
      if(_zz_2682_)begin
        int_reg_array_48_38_imag <= _zz_2696_;
      end
      if(_zz_2683_)begin
        int_reg_array_48_39_imag <= _zz_2696_;
      end
      if(_zz_2684_)begin
        int_reg_array_48_40_imag <= _zz_2696_;
      end
      if(_zz_2685_)begin
        int_reg_array_48_41_imag <= _zz_2696_;
      end
      if(_zz_2686_)begin
        int_reg_array_48_42_imag <= _zz_2696_;
      end
      if(_zz_2687_)begin
        int_reg_array_48_43_imag <= _zz_2696_;
      end
      if(_zz_2688_)begin
        int_reg_array_48_44_imag <= _zz_2696_;
      end
      if(_zz_2689_)begin
        int_reg_array_48_45_imag <= _zz_2696_;
      end
      if(_zz_2690_)begin
        int_reg_array_48_46_imag <= _zz_2696_;
      end
      if(_zz_2691_)begin
        int_reg_array_48_47_imag <= _zz_2696_;
      end
      if(_zz_2692_)begin
        int_reg_array_48_48_imag <= _zz_2696_;
      end
      if(_zz_2693_)begin
        int_reg_array_48_49_imag <= _zz_2696_;
      end
      if(_zz_2699_)begin
        int_reg_array_49_0_real <= _zz_2750_;
      end
      if(_zz_2700_)begin
        int_reg_array_49_1_real <= _zz_2750_;
      end
      if(_zz_2701_)begin
        int_reg_array_49_2_real <= _zz_2750_;
      end
      if(_zz_2702_)begin
        int_reg_array_49_3_real <= _zz_2750_;
      end
      if(_zz_2703_)begin
        int_reg_array_49_4_real <= _zz_2750_;
      end
      if(_zz_2704_)begin
        int_reg_array_49_5_real <= _zz_2750_;
      end
      if(_zz_2705_)begin
        int_reg_array_49_6_real <= _zz_2750_;
      end
      if(_zz_2706_)begin
        int_reg_array_49_7_real <= _zz_2750_;
      end
      if(_zz_2707_)begin
        int_reg_array_49_8_real <= _zz_2750_;
      end
      if(_zz_2708_)begin
        int_reg_array_49_9_real <= _zz_2750_;
      end
      if(_zz_2709_)begin
        int_reg_array_49_10_real <= _zz_2750_;
      end
      if(_zz_2710_)begin
        int_reg_array_49_11_real <= _zz_2750_;
      end
      if(_zz_2711_)begin
        int_reg_array_49_12_real <= _zz_2750_;
      end
      if(_zz_2712_)begin
        int_reg_array_49_13_real <= _zz_2750_;
      end
      if(_zz_2713_)begin
        int_reg_array_49_14_real <= _zz_2750_;
      end
      if(_zz_2714_)begin
        int_reg_array_49_15_real <= _zz_2750_;
      end
      if(_zz_2715_)begin
        int_reg_array_49_16_real <= _zz_2750_;
      end
      if(_zz_2716_)begin
        int_reg_array_49_17_real <= _zz_2750_;
      end
      if(_zz_2717_)begin
        int_reg_array_49_18_real <= _zz_2750_;
      end
      if(_zz_2718_)begin
        int_reg_array_49_19_real <= _zz_2750_;
      end
      if(_zz_2719_)begin
        int_reg_array_49_20_real <= _zz_2750_;
      end
      if(_zz_2720_)begin
        int_reg_array_49_21_real <= _zz_2750_;
      end
      if(_zz_2721_)begin
        int_reg_array_49_22_real <= _zz_2750_;
      end
      if(_zz_2722_)begin
        int_reg_array_49_23_real <= _zz_2750_;
      end
      if(_zz_2723_)begin
        int_reg_array_49_24_real <= _zz_2750_;
      end
      if(_zz_2724_)begin
        int_reg_array_49_25_real <= _zz_2750_;
      end
      if(_zz_2725_)begin
        int_reg_array_49_26_real <= _zz_2750_;
      end
      if(_zz_2726_)begin
        int_reg_array_49_27_real <= _zz_2750_;
      end
      if(_zz_2727_)begin
        int_reg_array_49_28_real <= _zz_2750_;
      end
      if(_zz_2728_)begin
        int_reg_array_49_29_real <= _zz_2750_;
      end
      if(_zz_2729_)begin
        int_reg_array_49_30_real <= _zz_2750_;
      end
      if(_zz_2730_)begin
        int_reg_array_49_31_real <= _zz_2750_;
      end
      if(_zz_2731_)begin
        int_reg_array_49_32_real <= _zz_2750_;
      end
      if(_zz_2732_)begin
        int_reg_array_49_33_real <= _zz_2750_;
      end
      if(_zz_2733_)begin
        int_reg_array_49_34_real <= _zz_2750_;
      end
      if(_zz_2734_)begin
        int_reg_array_49_35_real <= _zz_2750_;
      end
      if(_zz_2735_)begin
        int_reg_array_49_36_real <= _zz_2750_;
      end
      if(_zz_2736_)begin
        int_reg_array_49_37_real <= _zz_2750_;
      end
      if(_zz_2737_)begin
        int_reg_array_49_38_real <= _zz_2750_;
      end
      if(_zz_2738_)begin
        int_reg_array_49_39_real <= _zz_2750_;
      end
      if(_zz_2739_)begin
        int_reg_array_49_40_real <= _zz_2750_;
      end
      if(_zz_2740_)begin
        int_reg_array_49_41_real <= _zz_2750_;
      end
      if(_zz_2741_)begin
        int_reg_array_49_42_real <= _zz_2750_;
      end
      if(_zz_2742_)begin
        int_reg_array_49_43_real <= _zz_2750_;
      end
      if(_zz_2743_)begin
        int_reg_array_49_44_real <= _zz_2750_;
      end
      if(_zz_2744_)begin
        int_reg_array_49_45_real <= _zz_2750_;
      end
      if(_zz_2745_)begin
        int_reg_array_49_46_real <= _zz_2750_;
      end
      if(_zz_2746_)begin
        int_reg_array_49_47_real <= _zz_2750_;
      end
      if(_zz_2747_)begin
        int_reg_array_49_48_real <= _zz_2750_;
      end
      if(_zz_2748_)begin
        int_reg_array_49_49_real <= _zz_2750_;
      end
      if(_zz_2699_)begin
        int_reg_array_49_0_imag <= _zz_2751_;
      end
      if(_zz_2700_)begin
        int_reg_array_49_1_imag <= _zz_2751_;
      end
      if(_zz_2701_)begin
        int_reg_array_49_2_imag <= _zz_2751_;
      end
      if(_zz_2702_)begin
        int_reg_array_49_3_imag <= _zz_2751_;
      end
      if(_zz_2703_)begin
        int_reg_array_49_4_imag <= _zz_2751_;
      end
      if(_zz_2704_)begin
        int_reg_array_49_5_imag <= _zz_2751_;
      end
      if(_zz_2705_)begin
        int_reg_array_49_6_imag <= _zz_2751_;
      end
      if(_zz_2706_)begin
        int_reg_array_49_7_imag <= _zz_2751_;
      end
      if(_zz_2707_)begin
        int_reg_array_49_8_imag <= _zz_2751_;
      end
      if(_zz_2708_)begin
        int_reg_array_49_9_imag <= _zz_2751_;
      end
      if(_zz_2709_)begin
        int_reg_array_49_10_imag <= _zz_2751_;
      end
      if(_zz_2710_)begin
        int_reg_array_49_11_imag <= _zz_2751_;
      end
      if(_zz_2711_)begin
        int_reg_array_49_12_imag <= _zz_2751_;
      end
      if(_zz_2712_)begin
        int_reg_array_49_13_imag <= _zz_2751_;
      end
      if(_zz_2713_)begin
        int_reg_array_49_14_imag <= _zz_2751_;
      end
      if(_zz_2714_)begin
        int_reg_array_49_15_imag <= _zz_2751_;
      end
      if(_zz_2715_)begin
        int_reg_array_49_16_imag <= _zz_2751_;
      end
      if(_zz_2716_)begin
        int_reg_array_49_17_imag <= _zz_2751_;
      end
      if(_zz_2717_)begin
        int_reg_array_49_18_imag <= _zz_2751_;
      end
      if(_zz_2718_)begin
        int_reg_array_49_19_imag <= _zz_2751_;
      end
      if(_zz_2719_)begin
        int_reg_array_49_20_imag <= _zz_2751_;
      end
      if(_zz_2720_)begin
        int_reg_array_49_21_imag <= _zz_2751_;
      end
      if(_zz_2721_)begin
        int_reg_array_49_22_imag <= _zz_2751_;
      end
      if(_zz_2722_)begin
        int_reg_array_49_23_imag <= _zz_2751_;
      end
      if(_zz_2723_)begin
        int_reg_array_49_24_imag <= _zz_2751_;
      end
      if(_zz_2724_)begin
        int_reg_array_49_25_imag <= _zz_2751_;
      end
      if(_zz_2725_)begin
        int_reg_array_49_26_imag <= _zz_2751_;
      end
      if(_zz_2726_)begin
        int_reg_array_49_27_imag <= _zz_2751_;
      end
      if(_zz_2727_)begin
        int_reg_array_49_28_imag <= _zz_2751_;
      end
      if(_zz_2728_)begin
        int_reg_array_49_29_imag <= _zz_2751_;
      end
      if(_zz_2729_)begin
        int_reg_array_49_30_imag <= _zz_2751_;
      end
      if(_zz_2730_)begin
        int_reg_array_49_31_imag <= _zz_2751_;
      end
      if(_zz_2731_)begin
        int_reg_array_49_32_imag <= _zz_2751_;
      end
      if(_zz_2732_)begin
        int_reg_array_49_33_imag <= _zz_2751_;
      end
      if(_zz_2733_)begin
        int_reg_array_49_34_imag <= _zz_2751_;
      end
      if(_zz_2734_)begin
        int_reg_array_49_35_imag <= _zz_2751_;
      end
      if(_zz_2735_)begin
        int_reg_array_49_36_imag <= _zz_2751_;
      end
      if(_zz_2736_)begin
        int_reg_array_49_37_imag <= _zz_2751_;
      end
      if(_zz_2737_)begin
        int_reg_array_49_38_imag <= _zz_2751_;
      end
      if(_zz_2738_)begin
        int_reg_array_49_39_imag <= _zz_2751_;
      end
      if(_zz_2739_)begin
        int_reg_array_49_40_imag <= _zz_2751_;
      end
      if(_zz_2740_)begin
        int_reg_array_49_41_imag <= _zz_2751_;
      end
      if(_zz_2741_)begin
        int_reg_array_49_42_imag <= _zz_2751_;
      end
      if(_zz_2742_)begin
        int_reg_array_49_43_imag <= _zz_2751_;
      end
      if(_zz_2743_)begin
        int_reg_array_49_44_imag <= _zz_2751_;
      end
      if(_zz_2744_)begin
        int_reg_array_49_45_imag <= _zz_2751_;
      end
      if(_zz_2745_)begin
        int_reg_array_49_46_imag <= _zz_2751_;
      end
      if(_zz_2746_)begin
        int_reg_array_49_47_imag <= _zz_2751_;
      end
      if(_zz_2747_)begin
        int_reg_array_49_48_imag <= _zz_2751_;
      end
      if(_zz_2748_)begin
        int_reg_array_49_49_imag <= _zz_2751_;
      end
    end
  end

  always @ (posedge clk or posedge reset) begin
    if (reset) begin
      load_data_area_current_addr <= 32'h0;
    end else begin
      if(axi4_w_valid)begin
        load_data_area_current_addr <= Axi4Incr_result;
      end
    end
  end

  always @ (posedge clk) begin
    axi4_w_payload_data_regNext <= axi4_w_payload_data;
  end


endmodule
